module basic_2000_20000_2500_25_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1912,In_205);
or U1 (N_1,In_495,In_317);
xor U2 (N_2,In_1160,In_530);
or U3 (N_3,In_1837,In_1044);
xor U4 (N_4,In_411,In_1388);
nand U5 (N_5,In_519,In_840);
or U6 (N_6,In_1868,In_731);
and U7 (N_7,In_1309,In_136);
or U8 (N_8,In_646,In_36);
xnor U9 (N_9,In_717,In_1575);
nor U10 (N_10,In_71,In_595);
nand U11 (N_11,In_603,In_1719);
nand U12 (N_12,In_1104,In_358);
nor U13 (N_13,In_851,In_1282);
and U14 (N_14,In_1821,In_1188);
and U15 (N_15,In_1470,In_765);
or U16 (N_16,In_1169,In_927);
and U17 (N_17,In_1720,In_1899);
nand U18 (N_18,In_876,In_874);
xor U19 (N_19,In_1963,In_941);
or U20 (N_20,In_648,In_284);
or U21 (N_21,In_1448,In_1469);
and U22 (N_22,In_1123,In_84);
and U23 (N_23,In_700,In_797);
or U24 (N_24,In_1498,In_1763);
and U25 (N_25,In_50,In_1144);
or U26 (N_26,In_1019,In_1693);
and U27 (N_27,In_1096,In_747);
xnor U28 (N_28,In_100,In_1822);
nand U29 (N_29,In_526,In_327);
or U30 (N_30,In_107,In_1924);
nor U31 (N_31,In_1077,In_393);
nor U32 (N_32,In_1460,In_1292);
nand U33 (N_33,In_1039,In_764);
or U34 (N_34,In_1185,In_65);
xnor U35 (N_35,In_249,In_506);
or U36 (N_36,In_1653,In_846);
nor U37 (N_37,In_1259,In_493);
nand U38 (N_38,In_273,In_268);
or U39 (N_39,In_342,In_1594);
nand U40 (N_40,In_1327,In_1948);
and U41 (N_41,In_948,In_966);
and U42 (N_42,In_908,In_1084);
or U43 (N_43,In_191,In_1781);
nor U44 (N_44,In_1983,In_281);
nor U45 (N_45,In_68,In_1136);
xor U46 (N_46,In_839,In_1848);
and U47 (N_47,In_684,In_716);
xnor U48 (N_48,In_1744,In_993);
nor U49 (N_49,In_135,In_954);
nand U50 (N_50,In_338,In_254);
nand U51 (N_51,In_1794,In_287);
xor U52 (N_52,In_1145,In_1355);
nand U53 (N_53,In_1254,In_1587);
nor U54 (N_54,In_726,In_1263);
nor U55 (N_55,In_178,In_473);
nor U56 (N_56,In_538,In_776);
or U57 (N_57,In_1181,In_15);
nor U58 (N_58,In_924,In_1844);
nor U59 (N_59,In_313,In_1356);
and U60 (N_60,In_754,In_1116);
and U61 (N_61,In_322,In_44);
and U62 (N_62,In_1676,In_1289);
or U63 (N_63,In_520,In_1729);
nand U64 (N_64,In_374,In_1885);
nor U65 (N_65,In_1688,In_1463);
and U66 (N_66,In_918,In_718);
xnor U67 (N_67,In_1101,In_184);
nand U68 (N_68,In_1870,In_1256);
nor U69 (N_69,In_768,In_219);
nor U70 (N_70,In_841,In_1206);
and U71 (N_71,In_577,In_1678);
nand U72 (N_72,In_1775,In_827);
nor U73 (N_73,In_1212,In_1863);
nor U74 (N_74,In_451,In_467);
nand U75 (N_75,In_1825,In_1590);
nand U76 (N_76,In_1417,In_1467);
or U77 (N_77,In_346,In_759);
xnor U78 (N_78,In_807,In_1666);
xor U79 (N_79,In_1051,In_1006);
nand U80 (N_80,In_1357,In_1619);
or U81 (N_81,In_898,In_814);
or U82 (N_82,In_1570,In_1758);
nor U83 (N_83,In_537,In_750);
nor U84 (N_84,In_240,In_864);
and U85 (N_85,In_1397,In_1779);
nor U86 (N_86,In_945,In_366);
nor U87 (N_87,In_1815,In_1886);
and U88 (N_88,In_891,In_434);
or U89 (N_89,In_630,In_1050);
or U90 (N_90,In_19,In_328);
xor U91 (N_91,In_1313,In_562);
nor U92 (N_92,In_799,In_1090);
or U93 (N_93,In_1344,In_126);
or U94 (N_94,In_1632,In_1927);
xor U95 (N_95,In_987,In_1195);
and U96 (N_96,In_1211,In_881);
or U97 (N_97,In_984,In_410);
nand U98 (N_98,In_431,In_792);
xor U99 (N_99,In_31,In_1841);
nor U100 (N_100,In_246,In_504);
and U101 (N_101,In_1478,In_1119);
and U102 (N_102,In_942,In_962);
nor U103 (N_103,In_1319,In_277);
and U104 (N_104,In_999,In_594);
nand U105 (N_105,In_1706,In_415);
nor U106 (N_106,In_173,In_632);
and U107 (N_107,In_1163,In_1329);
or U108 (N_108,In_832,In_967);
or U109 (N_109,In_816,In_1400);
nand U110 (N_110,In_748,In_1554);
or U111 (N_111,In_472,In_1147);
nor U112 (N_112,In_509,In_1129);
nand U113 (N_113,In_800,In_1081);
or U114 (N_114,In_705,In_521);
xnor U115 (N_115,In_1975,In_271);
nand U116 (N_116,In_1978,In_805);
nor U117 (N_117,In_1384,In_818);
xnor U118 (N_118,In_917,In_586);
and U119 (N_119,In_546,In_713);
nor U120 (N_120,In_1152,In_87);
or U121 (N_121,In_911,In_1450);
and U122 (N_122,In_306,In_1777);
and U123 (N_123,In_496,In_1043);
xnor U124 (N_124,In_1317,In_784);
or U125 (N_125,In_949,In_261);
or U126 (N_126,In_398,In_760);
or U127 (N_127,In_1243,In_310);
nand U128 (N_128,In_1035,In_875);
or U129 (N_129,In_1511,In_1331);
and U130 (N_130,In_1823,In_968);
nand U131 (N_131,In_117,In_1860);
and U132 (N_132,In_303,In_953);
xnor U133 (N_133,In_1003,In_873);
nor U134 (N_134,In_1434,In_605);
xor U135 (N_135,In_479,In_1293);
nand U136 (N_136,In_588,In_1800);
or U137 (N_137,In_1962,In_1440);
nand U138 (N_138,In_1459,In_266);
or U139 (N_139,In_934,In_34);
nand U140 (N_140,In_1454,In_659);
and U141 (N_141,In_1974,In_1651);
or U142 (N_142,In_1894,In_429);
and U143 (N_143,In_1342,In_815);
xnor U144 (N_144,In_1114,In_762);
nand U145 (N_145,In_318,In_123);
nand U146 (N_146,In_641,In_1407);
nor U147 (N_147,In_1674,In_1445);
and U148 (N_148,In_323,In_1545);
nand U149 (N_149,In_1071,In_693);
nor U150 (N_150,In_1449,In_572);
nand U151 (N_151,In_1190,In_1656);
nand U152 (N_152,In_1154,In_1032);
nor U153 (N_153,In_1618,In_143);
and U154 (N_154,In_735,In_1170);
xor U155 (N_155,In_1739,In_1857);
xor U156 (N_156,In_1380,In_212);
nand U157 (N_157,In_264,In_1913);
xor U158 (N_158,In_1178,In_1245);
xnor U159 (N_159,In_1012,In_1193);
and U160 (N_160,In_217,In_1923);
xnor U161 (N_161,In_608,In_964);
nor U162 (N_162,In_391,In_1695);
nand U163 (N_163,In_1146,In_1661);
xnor U164 (N_164,In_422,In_542);
or U165 (N_165,In_475,In_1063);
and U166 (N_166,In_940,In_1864);
xor U167 (N_167,In_1303,In_892);
nand U168 (N_168,In_298,In_1166);
nor U169 (N_169,In_179,In_823);
or U170 (N_170,In_516,In_1061);
nand U171 (N_171,In_348,In_335);
nand U172 (N_172,In_736,In_1062);
nand U173 (N_173,In_1403,In_1711);
nand U174 (N_174,In_1861,In_373);
nand U175 (N_175,In_150,In_216);
or U176 (N_176,In_1369,In_947);
xnor U177 (N_177,In_1031,In_1872);
nor U178 (N_178,In_1907,In_337);
or U179 (N_179,In_1422,In_1785);
nor U180 (N_180,In_1892,In_676);
and U181 (N_181,In_1811,In_529);
nand U182 (N_182,In_231,In_969);
and U183 (N_183,In_1205,In_1843);
and U184 (N_184,In_704,In_424);
and U185 (N_185,In_963,In_1073);
xnor U186 (N_186,In_1749,In_1559);
xnor U187 (N_187,In_372,In_1672);
nor U188 (N_188,In_1348,In_336);
and U189 (N_189,In_35,In_1476);
nand U190 (N_190,In_1566,In_1360);
and U191 (N_191,In_1829,In_1471);
nor U192 (N_192,In_796,In_1772);
or U193 (N_193,In_541,In_213);
nor U194 (N_194,In_75,In_1065);
xnor U195 (N_195,In_1228,In_1932);
nand U196 (N_196,In_1396,In_331);
and U197 (N_197,In_210,In_1548);
and U198 (N_198,In_1067,In_1410);
or U199 (N_199,In_1778,In_972);
and U200 (N_200,In_142,In_1328);
nand U201 (N_201,In_1516,In_1472);
and U202 (N_202,In_152,In_952);
xnor U203 (N_203,In_308,In_1041);
or U204 (N_204,In_1350,In_879);
nor U205 (N_205,In_958,In_442);
and U206 (N_206,In_364,In_1072);
nor U207 (N_207,In_1264,In_1918);
nor U208 (N_208,In_1036,In_1806);
and U209 (N_209,In_767,In_1338);
xor U210 (N_210,In_181,In_443);
xor U211 (N_211,In_33,In_503);
or U212 (N_212,In_1708,In_1173);
or U213 (N_213,In_1855,In_1761);
or U214 (N_214,In_1372,In_1518);
or U215 (N_215,In_1808,In_302);
and U216 (N_216,In_1877,In_689);
or U217 (N_217,In_1294,In_1724);
nand U218 (N_218,In_761,In_1268);
nor U219 (N_219,In_105,In_709);
xnor U220 (N_220,In_359,In_1972);
nor U221 (N_221,In_356,In_779);
nor U222 (N_222,In_230,In_899);
and U223 (N_223,In_532,In_853);
xnor U224 (N_224,In_719,In_1311);
or U225 (N_225,In_885,In_108);
or U226 (N_226,In_1520,In_666);
or U227 (N_227,In_1222,In_599);
and U228 (N_228,In_852,In_24);
xnor U229 (N_229,In_1611,In_703);
or U230 (N_230,In_1934,In_1588);
or U231 (N_231,In_1537,In_1412);
and U232 (N_232,In_1982,In_1842);
and U233 (N_233,In_1510,In_1846);
or U234 (N_234,In_817,In_724);
or U235 (N_235,In_580,In_1789);
or U236 (N_236,In_1964,In_1229);
nand U237 (N_237,In_1603,In_569);
or U238 (N_238,In_174,In_843);
nand U239 (N_239,In_1503,In_1179);
or U240 (N_240,In_482,In_1701);
xor U241 (N_241,In_511,In_560);
and U242 (N_242,In_534,In_1379);
nor U243 (N_243,In_1158,In_1394);
xnor U244 (N_244,In_1240,In_1607);
or U245 (N_245,In_417,In_1917);
or U246 (N_246,In_1446,In_1456);
nand U247 (N_247,In_1272,In_1307);
and U248 (N_248,In_1895,In_830);
and U249 (N_249,In_1536,In_1954);
or U250 (N_250,In_1896,In_1792);
or U251 (N_251,In_1585,In_771);
and U252 (N_252,In_674,In_187);
xnor U253 (N_253,In_444,In_494);
nand U254 (N_254,In_665,In_1906);
or U255 (N_255,In_638,In_315);
nor U256 (N_256,In_1491,In_1699);
and U257 (N_257,In_725,In_1018);
nand U258 (N_258,In_656,In_1248);
xnor U259 (N_259,In_1143,In_1713);
nand U260 (N_260,In_1984,In_1453);
nor U261 (N_261,In_286,In_1740);
xor U262 (N_262,In_1312,In_921);
or U263 (N_263,In_1920,In_757);
xor U264 (N_264,In_76,In_1552);
or U265 (N_265,In_402,In_1052);
nor U266 (N_266,In_545,In_606);
nor U267 (N_267,In_1675,In_118);
nand U268 (N_268,In_939,In_1636);
nor U269 (N_269,In_1564,In_722);
nor U270 (N_270,In_125,In_1217);
xor U271 (N_271,In_1945,In_8);
nand U272 (N_272,In_414,In_396);
xnor U273 (N_273,In_986,In_379);
nand U274 (N_274,In_407,In_73);
nand U275 (N_275,In_675,In_1939);
and U276 (N_276,In_1582,In_25);
nand U277 (N_277,In_865,In_1308);
or U278 (N_278,In_980,In_45);
xor U279 (N_279,In_289,In_883);
xnor U280 (N_280,In_1990,In_459);
nand U281 (N_281,In_806,In_637);
nand U282 (N_282,In_1743,In_32);
and U283 (N_283,In_772,In_1659);
nor U284 (N_284,In_1466,In_733);
nor U285 (N_285,In_103,In_824);
nor U286 (N_286,In_37,In_0);
nor U287 (N_287,In_1302,In_1483);
xnor U288 (N_288,In_995,In_1133);
or U289 (N_289,In_826,In_1057);
and U290 (N_290,In_894,In_753);
or U291 (N_291,In_1754,In_1058);
and U292 (N_292,In_1405,In_1223);
nand U293 (N_293,In_460,In_1782);
nor U294 (N_294,In_621,In_1813);
and U295 (N_295,In_1458,In_845);
nand U296 (N_296,In_1647,In_1315);
nand U297 (N_297,In_682,In_1845);
xnor U298 (N_298,In_1935,In_701);
xor U299 (N_299,In_5,In_1122);
and U300 (N_300,In_868,In_1669);
nand U301 (N_301,In_1325,In_1128);
or U302 (N_302,In_1125,In_470);
and U303 (N_303,In_250,In_644);
nand U304 (N_304,In_354,In_1411);
nor U305 (N_305,In_1183,In_1241);
or U306 (N_306,In_159,In_1750);
xnor U307 (N_307,In_651,In_1488);
xor U308 (N_308,In_279,In_56);
nor U309 (N_309,In_1765,In_1343);
nor U310 (N_310,In_1149,In_309);
xor U311 (N_311,In_1883,In_307);
nand U312 (N_312,In_1658,In_1650);
nand U313 (N_313,In_631,In_887);
nor U314 (N_314,In_766,In_893);
xnor U315 (N_315,In_1504,In_12);
nand U316 (N_316,In_1056,In_1363);
and U317 (N_317,In_1465,In_1105);
and U318 (N_318,In_614,In_928);
xor U319 (N_319,In_1118,In_1595);
or U320 (N_320,In_1768,In_755);
nor U321 (N_321,In_1722,In_344);
xnor U322 (N_322,In_668,In_1486);
xor U323 (N_323,In_1887,In_1297);
or U324 (N_324,In_1989,In_1383);
nand U325 (N_325,In_1871,In_869);
nor U326 (N_326,In_828,In_332);
or U327 (N_327,In_1649,In_794);
and U328 (N_328,In_1578,In_1340);
and U329 (N_329,In_262,In_488);
nor U330 (N_330,In_1783,In_996);
nand U331 (N_331,In_1210,In_1539);
xor U332 (N_332,In_1878,In_1828);
nor U333 (N_333,In_1555,In_1421);
and U334 (N_334,In_1902,In_1291);
or U335 (N_335,In_923,In_58);
nor U336 (N_336,In_1691,In_448);
or U337 (N_337,In_413,In_1441);
xnor U338 (N_338,In_28,In_1477);
xnor U339 (N_339,In_990,In_1452);
nand U340 (N_340,In_522,In_485);
nand U341 (N_341,In_1176,In_1365);
nor U342 (N_342,In_1506,In_1958);
nor U343 (N_343,In_1787,In_1544);
nor U344 (N_344,In_1267,In_1873);
nor U345 (N_345,In_533,In_1533);
nand U346 (N_346,In_1599,In_1574);
xnor U347 (N_347,In_1694,In_1189);
and U348 (N_348,In_1199,In_738);
nor U349 (N_349,In_1606,In_188);
and U350 (N_350,In_175,In_549);
xor U351 (N_351,In_1364,In_801);
nor U352 (N_352,In_1943,In_343);
nor U353 (N_353,In_1604,In_206);
or U354 (N_354,In_1629,In_1089);
and U355 (N_355,In_955,In_436);
or U356 (N_356,In_1735,In_1583);
nand U357 (N_357,In_746,In_1076);
nand U358 (N_358,In_1002,In_296);
xnor U359 (N_359,In_938,In_1856);
nor U360 (N_360,In_1086,In_1203);
nand U361 (N_361,In_1126,In_1091);
nand U362 (N_362,In_1697,In_10);
xnor U363 (N_363,In_1234,In_395);
nor U364 (N_364,In_1623,In_388);
or U365 (N_365,In_320,In_1786);
and U366 (N_366,In_1026,In_769);
nand U367 (N_367,In_1078,In_554);
nand U368 (N_368,In_355,In_678);
nand U369 (N_369,In_23,In_1534);
and U370 (N_370,In_1949,In_548);
nor U371 (N_371,In_507,In_596);
or U372 (N_372,In_1529,In_1700);
and U373 (N_373,In_1151,In_426);
xnor U374 (N_374,In_1517,In_6);
xor U375 (N_375,In_1579,In_790);
or U376 (N_376,In_812,In_362);
nand U377 (N_377,In_706,In_186);
and U378 (N_378,In_134,In_177);
or U379 (N_379,In_1771,In_502);
xor U380 (N_380,In_1580,In_285);
nand U381 (N_381,In_745,In_360);
and U382 (N_382,In_994,In_381);
nor U383 (N_383,In_438,In_565);
xor U384 (N_384,In_930,In_623);
and U385 (N_385,In_581,In_1029);
and U386 (N_386,In_804,In_1762);
or U387 (N_387,In_1351,In_825);
xnor U388 (N_388,In_1148,In_1074);
or U389 (N_389,In_1398,In_1279);
and U390 (N_390,In_74,In_446);
or U391 (N_391,In_243,In_1326);
or U392 (N_392,In_242,In_1462);
or U393 (N_393,In_1741,In_1847);
and U394 (N_394,In_855,In_627);
xor U395 (N_395,In_1998,In_1499);
and U396 (N_396,In_283,In_1936);
nor U397 (N_397,In_829,In_1484);
nand U398 (N_398,In_1435,In_385);
xor U399 (N_399,In_1959,In_1247);
or U400 (N_400,In_1494,In_867);
nor U401 (N_401,In_456,In_18);
xor U402 (N_402,In_1730,In_1481);
and U403 (N_403,In_1752,In_1374);
xor U404 (N_404,In_180,In_214);
nor U405 (N_405,In_1736,In_933);
or U406 (N_406,In_278,In_1625);
nand U407 (N_407,In_1733,In_365);
and U408 (N_408,In_1524,In_93);
xnor U409 (N_409,In_575,In_1055);
xor U410 (N_410,In_1005,In_1634);
and U411 (N_411,In_113,In_418);
or U412 (N_412,In_1513,In_428);
nor U413 (N_413,In_1921,In_793);
or U414 (N_414,In_808,In_1996);
nand U415 (N_415,In_1010,In_591);
nor U416 (N_416,In_1541,In_232);
xnor U417 (N_417,In_1406,In_1956);
nor U418 (N_418,In_1341,In_1371);
nor U419 (N_419,In_880,In_1770);
xor U420 (N_420,In_587,In_333);
xor U421 (N_421,In_66,In_1621);
xor U422 (N_422,In_1930,In_325);
and U423 (N_423,In_169,In_1358);
or U424 (N_424,In_1682,In_1137);
and U425 (N_425,In_492,In_201);
nor U426 (N_426,In_1523,In_1285);
or U427 (N_427,In_405,In_256);
and U428 (N_428,In_1776,In_461);
xor U429 (N_429,In_836,In_609);
xnor U430 (N_430,In_61,In_1260);
nor U431 (N_431,In_1393,In_1816);
and U432 (N_432,In_1352,In_854);
or U433 (N_433,In_1028,In_1284);
nand U434 (N_434,In_1437,In_1495);
and U435 (N_435,In_1880,In_1296);
xnor U436 (N_436,In_137,In_389);
nand U437 (N_437,In_960,In_208);
nor U438 (N_438,In_1530,In_280);
xnor U439 (N_439,In_406,In_168);
nor U440 (N_440,In_267,In_165);
or U441 (N_441,In_1251,In_1278);
and U442 (N_442,In_1953,In_1696);
nand U443 (N_443,In_1280,In_1095);
nand U444 (N_444,In_985,In_1760);
nor U445 (N_445,In_314,In_1527);
and U446 (N_446,In_153,In_1947);
and U447 (N_447,In_1689,In_1631);
xnor U448 (N_448,In_895,In_345);
nand U449 (N_449,In_1994,In_1097);
nor U450 (N_450,In_1037,In_1270);
or U451 (N_451,In_1102,In_601);
nand U452 (N_452,In_774,In_1187);
nor U453 (N_453,In_1017,In_62);
or U454 (N_454,In_1444,In_570);
xor U455 (N_455,In_913,In_878);
and U456 (N_456,In_163,In_1392);
nand U457 (N_457,In_1370,In_1753);
and U458 (N_458,In_510,In_300);
and U459 (N_459,In_1904,In_896);
xor U460 (N_460,In_1550,In_1404);
and U461 (N_461,In_99,In_54);
nand U462 (N_462,In_721,In_1424);
nor U463 (N_463,In_1246,In_110);
and U464 (N_464,In_425,In_1113);
xnor U465 (N_465,In_781,In_1721);
and U466 (N_466,In_1426,In_1798);
and U467 (N_467,In_539,In_584);
and U468 (N_468,In_1926,In_129);
nor U469 (N_469,In_1347,In_1184);
nor U470 (N_470,In_162,In_900);
or U471 (N_471,In_600,In_88);
nor U472 (N_472,In_140,In_192);
or U473 (N_473,In_305,In_1299);
nor U474 (N_474,In_1960,In_859);
and U475 (N_475,In_920,In_1004);
nand U476 (N_476,In_775,In_399);
nand U477 (N_477,In_926,In_1138);
or U478 (N_478,In_612,In_1734);
xnor U479 (N_479,In_1409,In_1216);
and U480 (N_480,In_1723,In_1961);
xor U481 (N_481,In_639,In_525);
nand U482 (N_482,In_932,In_866);
and U483 (N_483,In_903,In_1117);
xnor U484 (N_484,In_288,In_518);
xor U485 (N_485,In_847,In_86);
and U486 (N_486,In_1318,In_1316);
and U487 (N_487,In_89,In_1876);
nand U488 (N_488,In_1718,In_291);
xnor U489 (N_489,In_401,In_1979);
nor U490 (N_490,In_1748,In_469);
and U491 (N_491,In_1509,In_732);
nand U492 (N_492,In_687,In_1690);
or U493 (N_493,In_1556,In_400);
and U494 (N_494,In_1232,In_710);
nor U495 (N_495,In_1333,In_1429);
and U496 (N_496,In_1009,In_1991);
xnor U497 (N_497,In_1637,In_904);
or U498 (N_498,In_340,In_311);
or U499 (N_499,In_1455,In_235);
nand U500 (N_500,In_189,In_1981);
and U501 (N_501,In_1221,In_578);
nor U502 (N_502,In_1571,In_369);
nand U503 (N_503,In_1253,In_1952);
or U504 (N_504,In_477,In_272);
nor U505 (N_505,In_1186,In_55);
nand U506 (N_506,In_1258,In_1747);
xor U507 (N_507,In_190,In_1999);
xor U508 (N_508,In_1985,In_1266);
and U509 (N_509,In_1769,In_301);
or U510 (N_510,In_367,In_1099);
xor U511 (N_511,In_218,In_1290);
nor U512 (N_512,In_615,In_649);
nor U513 (N_513,In_1764,In_1851);
or U514 (N_514,In_1933,In_421);
nor U515 (N_515,In_1614,In_1702);
and U516 (N_516,In_1395,In_81);
and U517 (N_517,In_773,In_1528);
or U518 (N_518,In_49,In_613);
or U519 (N_519,In_624,In_524);
and U520 (N_520,In_1168,In_1835);
or U521 (N_521,In_1814,In_112);
xor U522 (N_522,In_1602,In_514);
nor U523 (N_523,In_1336,In_171);
nand U524 (N_524,In_1859,In_59);
and U525 (N_525,In_1208,In_909);
xor U526 (N_526,In_1865,In_1833);
xnor U527 (N_527,In_798,In_1362);
xnor U528 (N_528,In_1642,In_47);
nand U529 (N_529,In_1480,In_1202);
nor U530 (N_530,In_1827,In_1834);
nor U531 (N_531,In_1738,In_1644);
nor U532 (N_532,In_63,In_590);
nand U533 (N_533,In_85,In_1218);
or U534 (N_534,In_1558,In_1755);
and U535 (N_535,In_116,In_41);
and U536 (N_536,In_622,In_239);
nor U537 (N_537,In_959,In_1977);
nor U538 (N_538,In_38,In_1773);
nand U539 (N_539,In_269,In_378);
nor U540 (N_540,In_1940,In_1922);
nand U541 (N_541,In_685,In_1387);
and U542 (N_542,In_1655,In_1714);
nand U543 (N_543,In_789,In_741);
nor U544 (N_544,In_1626,In_1354);
nand U545 (N_545,In_708,In_1283);
and U546 (N_546,In_863,In_1881);
nand U547 (N_547,In_1925,In_1732);
nor U548 (N_548,In_294,In_1505);
xor U549 (N_549,In_1201,In_1810);
nand U550 (N_550,In_1609,In_956);
nor U551 (N_551,In_777,In_274);
or U552 (N_552,In_1451,In_1322);
and U553 (N_553,In_1442,In_616);
nor U554 (N_554,In_1596,In_1492);
or U555 (N_555,In_40,In_363);
or U556 (N_556,In_1597,In_423);
and U557 (N_557,In_1898,In_1225);
nand U558 (N_558,In_453,In_77);
or U559 (N_559,In_559,In_371);
or U560 (N_560,In_445,In_645);
or U561 (N_561,In_1024,In_844);
nand U562 (N_562,In_53,In_1103);
nand U563 (N_563,In_1269,In_403);
xor U564 (N_564,In_1159,In_540);
and U565 (N_565,In_234,In_57);
nand U566 (N_566,In_1879,In_1633);
nand U567 (N_567,In_1993,In_94);
nand U568 (N_568,In_683,In_1054);
nand U569 (N_569,In_1500,In_1046);
xnor U570 (N_570,In_1986,In_1359);
nand U571 (N_571,In_1335,In_1542);
or U572 (N_572,In_199,In_1301);
and U573 (N_573,In_22,In_133);
xor U574 (N_574,In_1645,In_597);
and U575 (N_575,In_147,In_729);
xnor U576 (N_576,In_329,In_1903);
xnor U577 (N_577,In_1557,In_1261);
xor U578 (N_578,In_394,In_951);
or U579 (N_579,In_1436,In_463);
nor U580 (N_580,In_1973,In_1698);
xor U581 (N_581,In_929,In_919);
and U582 (N_582,In_1522,In_292);
or U583 (N_583,In_211,In_1592);
and U584 (N_584,In_669,In_711);
and U585 (N_585,In_1941,In_299);
nand U586 (N_586,In_1840,In_1124);
nor U587 (N_587,In_330,In_223);
and U588 (N_588,In_247,In_215);
xor U589 (N_589,In_770,In_43);
nand U590 (N_590,In_9,In_1938);
or U591 (N_591,In_1784,In_1164);
and U592 (N_592,In_1901,In_1382);
nand U593 (N_593,In_257,In_1802);
nor U594 (N_594,In_1438,In_447);
nor U595 (N_595,In_1155,In_1910);
xnor U596 (N_596,In_1000,In_1809);
and U597 (N_597,In_1546,In_1728);
or U598 (N_598,In_1069,In_936);
and U599 (N_599,In_1108,In_1858);
nand U600 (N_600,In_3,In_1106);
and U601 (N_601,In_1501,In_1635);
or U602 (N_602,In_1929,In_1390);
or U603 (N_603,In_751,In_244);
nand U604 (N_604,In_1230,In_409);
nand U605 (N_605,In_452,In_1415);
nand U606 (N_606,In_430,In_1161);
nand U607 (N_607,In_691,In_1746);
xnor U608 (N_608,In_149,In_1657);
or U609 (N_609,In_260,In_70);
nand U610 (N_610,In_988,In_566);
and U611 (N_611,In_1600,In_16);
nor U612 (N_612,In_1831,In_970);
xnor U613 (N_613,In_1027,In_1015);
nor U614 (N_614,In_1427,In_464);
nor U615 (N_615,In_1705,In_1153);
or U616 (N_616,In_1367,In_154);
nand U617 (N_617,In_1710,In_957);
xnor U618 (N_618,In_712,In_1021);
xor U619 (N_619,In_420,In_109);
nor U620 (N_620,In_1854,In_527);
or U621 (N_621,In_1820,In_1830);
or U622 (N_622,In_1897,In_120);
xor U623 (N_623,In_155,In_1496);
or U624 (N_624,In_48,In_1610);
or U625 (N_625,In_756,In_1332);
nor U626 (N_626,In_543,In_387);
xnor U627 (N_627,In_1167,In_1514);
nand U628 (N_628,In_1013,In_156);
xor U629 (N_629,In_1643,In_1493);
and U630 (N_630,In_1684,In_2);
and U631 (N_631,In_758,In_458);
xnor U632 (N_632,In_1969,In_151);
nor U633 (N_633,In_419,In_160);
or U634 (N_634,In_1242,In_647);
or U635 (N_635,In_650,In_1366);
nor U636 (N_636,In_1968,In_1692);
xnor U637 (N_637,In_640,In_227);
or U638 (N_638,In_324,In_1023);
nand U639 (N_639,In_450,In_1196);
or U640 (N_640,In_860,In_914);
nand U641 (N_641,In_1716,In_654);
or U642 (N_642,In_505,In_592);
or U643 (N_643,In_702,In_556);
or U644 (N_644,In_1804,In_204);
xor U645 (N_645,In_1014,In_658);
xor U646 (N_646,In_164,In_1497);
xnor U647 (N_647,In_1059,In_1172);
xor U648 (N_648,In_1572,In_1955);
nand U649 (N_649,In_500,In_1867);
nor U650 (N_650,In_1641,In_981);
or U651 (N_651,In_1121,In_241);
or U652 (N_652,In_558,In_1330);
or U653 (N_653,In_1717,In_1937);
or U654 (N_654,In_1640,In_1060);
and U655 (N_655,In_1034,In_350);
and U656 (N_656,In_697,In_1361);
and U657 (N_657,In_1432,In_1092);
or U658 (N_658,In_1219,In_1045);
or U659 (N_659,In_1304,In_1030);
or U660 (N_660,In_1737,In_297);
nor U661 (N_661,In_655,In_476);
or U662 (N_662,In_997,In_728);
xor U663 (N_663,In_78,In_1064);
xnor U664 (N_664,In_170,In_1679);
and U665 (N_665,In_1068,In_618);
or U666 (N_666,In_680,In_1378);
nand U667 (N_667,In_1731,In_907);
or U668 (N_668,In_1141,In_576);
nor U669 (N_669,In_1589,In_528);
and U670 (N_670,In_998,In_1345);
nand U671 (N_671,In_838,In_1563);
and U672 (N_672,In_782,In_316);
or U673 (N_673,In_925,In_730);
xor U674 (N_674,In_652,In_490);
nand U675 (N_675,In_304,In_635);
xnor U676 (N_676,In_1487,In_589);
or U677 (N_677,In_571,In_408);
or U678 (N_678,In_902,In_831);
xnor U679 (N_679,In_749,In_226);
xnor U680 (N_680,In_1997,In_1617);
nor U681 (N_681,In_837,In_435);
nand U682 (N_682,In_141,In_671);
or U683 (N_683,In_821,In_744);
nand U684 (N_684,In_157,In_1882);
xor U685 (N_685,In_1112,In_1812);
nor U686 (N_686,In_1414,In_1274);
and U687 (N_687,In_1224,In_1337);
or U688 (N_688,In_1875,In_1461);
xor U689 (N_689,In_4,In_198);
xnor U690 (N_690,In_811,In_579);
xor U691 (N_691,In_1826,In_585);
nand U692 (N_692,In_91,In_1408);
nand U693 (N_693,In_1852,In_1306);
nand U694 (N_694,In_229,In_1080);
or U695 (N_695,In_1215,In_1194);
or U696 (N_696,In_203,In_1681);
xor U697 (N_697,In_1134,In_1805);
xor U698 (N_698,In_1976,In_978);
xor U699 (N_699,In_848,In_568);
xor U700 (N_700,In_686,In_1667);
nor U701 (N_701,In_384,In_1321);
xor U702 (N_702,In_1376,In_194);
nand U703 (N_703,In_583,In_1853);
xnor U704 (N_704,In_1767,In_1418);
nor U705 (N_705,In_80,In_1389);
xor U706 (N_706,In_1704,In_1165);
nor U707 (N_707,In_1156,In_695);
nor U708 (N_708,In_1531,In_870);
and U709 (N_709,In_1756,In_1703);
and U710 (N_710,In_114,In_1443);
and U711 (N_711,In_146,In_861);
xor U712 (N_712,In_1946,In_433);
nand U713 (N_713,In_1475,In_1803);
or U714 (N_714,In_122,In_353);
xor U715 (N_715,In_1662,In_1576);
xnor U716 (N_716,In_386,In_484);
nand U717 (N_717,In_97,In_1900);
and U718 (N_718,In_1573,In_1638);
or U719 (N_719,In_17,In_523);
nor U720 (N_720,In_21,In_1271);
nor U721 (N_721,In_1162,In_1725);
nand U722 (N_722,In_803,In_1066);
or U723 (N_723,In_1048,In_788);
and U724 (N_724,In_1286,In_1265);
xor U725 (N_725,In_1323,In_357);
nor U726 (N_726,In_1416,In_1150);
and U727 (N_727,In_1560,In_1687);
nor U728 (N_728,In_1479,In_1233);
nor U729 (N_729,In_1001,In_1107);
nand U730 (N_730,In_101,In_563);
or U731 (N_731,In_46,In_1608);
or U732 (N_732,In_265,In_321);
xor U733 (N_733,In_167,In_255);
and U734 (N_734,In_822,In_481);
and U735 (N_735,In_193,In_633);
nand U736 (N_736,In_351,In_341);
xnor U737 (N_737,In_1909,In_1489);
nor U738 (N_738,In_1115,In_1276);
and U739 (N_739,In_857,In_1889);
nand U740 (N_740,In_1175,In_1673);
or U741 (N_741,In_884,In_1120);
xor U742 (N_742,In_380,In_1111);
xnor U743 (N_743,In_1180,In_1519);
or U744 (N_744,In_1569,In_1944);
xor U745 (N_745,In_1287,In_1049);
xor U746 (N_746,In_182,In_1818);
nor U747 (N_747,In_1807,In_1098);
nor U748 (N_748,In_973,In_1774);
xor U749 (N_749,In_787,In_1581);
and U750 (N_750,In_1796,In_1275);
or U751 (N_751,In_1238,In_1174);
xor U752 (N_752,In_282,In_468);
and U753 (N_753,In_1249,In_574);
or U754 (N_754,In_1433,In_83);
or U755 (N_755,In_1381,In_564);
xnor U756 (N_756,In_1237,In_1553);
or U757 (N_757,In_196,In_7);
xor U758 (N_758,In_145,In_517);
nand U759 (N_759,In_127,In_1866);
nor U760 (N_760,In_478,In_185);
nand U761 (N_761,In_780,In_1988);
nand U762 (N_762,In_901,In_849);
and U763 (N_763,In_1157,In_547);
nand U764 (N_764,In_30,In_222);
nand U765 (N_765,In_39,In_111);
xnor U766 (N_766,In_660,In_440);
xnor U767 (N_767,In_412,In_259);
nor U768 (N_768,In_1685,In_263);
xor U769 (N_769,In_989,In_290);
and U770 (N_770,In_1349,In_1874);
nor U771 (N_771,In_1093,In_1670);
nor U772 (N_772,In_1314,In_130);
nor U773 (N_773,In_1430,In_498);
or U774 (N_774,In_465,In_1965);
nand U775 (N_775,In_1742,In_915);
nand U776 (N_776,In_1709,In_166);
and U777 (N_777,In_626,In_392);
nor U778 (N_778,In_723,In_1082);
and U779 (N_779,In_742,In_1007);
xnor U780 (N_780,In_270,In_1135);
and U781 (N_781,In_119,In_661);
nand U782 (N_782,In_236,In_1227);
or U783 (N_783,In_20,In_1473);
or U784 (N_784,In_1040,In_1428);
nand U785 (N_785,In_1759,In_1368);
nand U786 (N_786,In_1915,In_739);
xor U787 (N_787,In_1891,In_376);
and U788 (N_788,In_1916,In_1817);
xor U789 (N_789,In_501,In_1987);
xor U790 (N_790,In_95,In_1131);
or U791 (N_791,In_1079,In_679);
or U792 (N_792,In_607,In_474);
nand U793 (N_793,In_1281,In_752);
nand U794 (N_794,In_727,In_1420);
nor U795 (N_795,In_833,In_276);
nand U796 (N_796,In_375,In_877);
nand U797 (N_797,In_1928,In_489);
and U798 (N_798,In_1235,In_245);
xnor U799 (N_799,In_416,In_1521);
nand U800 (N_800,In_1966,N_290);
nand U801 (N_801,In_1100,N_470);
nand U802 (N_802,N_696,In_1277);
nor U803 (N_803,In_544,N_710);
xnor U804 (N_804,N_468,N_549);
and U805 (N_805,In_383,N_294);
nor U806 (N_806,In_512,N_538);
xnor U807 (N_807,N_409,N_364);
and U808 (N_808,N_403,N_46);
or U809 (N_809,N_429,In_1593);
nor U810 (N_810,In_1132,N_720);
or U811 (N_811,In_1791,N_497);
nand U812 (N_812,N_207,In_937);
or U813 (N_813,In_582,N_231);
nor U814 (N_814,N_413,N_214);
xor U815 (N_815,N_41,N_483);
nor U816 (N_816,In_1950,N_487);
nor U817 (N_817,N_192,N_414);
or U818 (N_818,N_446,In_1239);
xnor U819 (N_819,N_285,N_713);
nand U820 (N_820,N_779,N_97);
and U821 (N_821,N_389,N_62);
and U822 (N_822,N_254,N_755);
nor U823 (N_823,N_501,N_114);
nand U824 (N_824,In_121,N_343);
xnor U825 (N_825,In_11,N_621);
xnor U826 (N_826,N_158,N_649);
nand U827 (N_827,N_173,In_890);
nand U828 (N_828,N_616,N_243);
nand U829 (N_829,N_111,N_208);
or U830 (N_830,N_126,In_1464);
xnor U831 (N_831,N_560,N_740);
nor U832 (N_832,N_84,N_175);
and U833 (N_833,N_204,N_199);
nand U834 (N_834,N_225,N_556);
or U835 (N_835,In_1712,In_251);
or U836 (N_836,In_791,N_319);
and U837 (N_837,N_259,In_221);
nand U838 (N_838,In_1905,N_261);
and U839 (N_839,N_421,N_190);
and U840 (N_840,In_1385,N_42);
nor U841 (N_841,In_491,N_134);
nand U842 (N_842,N_291,N_110);
nand U843 (N_843,N_39,N_671);
xor U844 (N_844,In_629,N_411);
xor U845 (N_845,N_642,N_360);
xor U846 (N_846,N_433,In_42);
xor U847 (N_847,In_27,N_639);
or U848 (N_848,In_611,In_1795);
nand U849 (N_849,N_734,In_1677);
or U850 (N_850,N_438,N_26);
and U851 (N_851,N_528,N_416);
xor U852 (N_852,N_310,N_187);
or U853 (N_853,N_99,N_792);
nor U854 (N_854,N_33,In_916);
nor U855 (N_855,N_386,N_732);
xnor U856 (N_856,N_674,In_377);
nand U857 (N_857,N_542,In_1020);
and U858 (N_858,N_11,N_377);
nand U859 (N_859,N_257,In_1538);
nand U860 (N_860,N_506,N_241);
nand U861 (N_861,In_1660,In_535);
nor U862 (N_862,N_85,In_1757);
xnor U863 (N_863,N_338,N_320);
and U864 (N_864,N_10,N_215);
or U865 (N_865,In_361,N_605);
and U866 (N_866,N_183,N_361);
xor U867 (N_867,N_584,In_912);
nand U868 (N_868,N_171,N_43);
or U869 (N_869,N_131,N_741);
nand U870 (N_870,N_434,In_1967);
nor U871 (N_871,N_680,N_169);
xnor U872 (N_872,In_1022,In_1310);
xor U873 (N_873,N_572,In_1042);
nor U874 (N_874,N_17,N_25);
nor U875 (N_875,N_238,In_1110);
or U876 (N_876,N_602,N_252);
or U877 (N_877,In_1515,N_188);
nor U878 (N_878,N_176,In_26);
nand U879 (N_879,N_758,In_1648);
and U880 (N_880,N_38,N_718);
nand U881 (N_881,In_1586,N_767);
nand U882 (N_882,N_725,In_228);
nand U883 (N_883,N_676,In_14);
xor U884 (N_884,N_482,In_1793);
xnor U885 (N_885,N_568,N_61);
and U886 (N_886,In_1008,In_1726);
xor U887 (N_887,In_195,N_559);
or U888 (N_888,N_461,N_406);
and U889 (N_889,N_390,N_366);
nor U890 (N_890,N_673,In_483);
xor U891 (N_891,N_128,N_628);
and U892 (N_892,In_220,N_139);
xor U893 (N_893,N_724,N_784);
xnor U894 (N_894,N_666,N_145);
nand U895 (N_895,N_711,N_473);
or U896 (N_896,In_1431,N_148);
nor U897 (N_897,In_1620,N_198);
nand U898 (N_898,N_441,In_778);
nand U899 (N_899,N_304,In_1549);
or U900 (N_900,In_551,N_562);
or U901 (N_901,In_397,In_92);
nor U902 (N_902,In_1033,N_194);
xnor U903 (N_903,N_200,In_610);
or U904 (N_904,N_702,In_1707);
nor U905 (N_905,N_342,In_720);
or U906 (N_906,In_1177,N_74);
and U907 (N_907,In_1577,N_532);
and U908 (N_908,In_1888,N_270);
or U909 (N_909,N_393,N_443);
xor U910 (N_910,N_459,In_82);
nand U911 (N_911,N_216,N_355);
nand U912 (N_912,N_112,In_977);
nor U913 (N_913,N_174,N_184);
nor U914 (N_914,N_729,N_60);
nor U915 (N_915,N_348,N_465);
nor U916 (N_916,N_689,N_777);
and U917 (N_917,In_486,In_698);
or U918 (N_918,N_283,N_594);
nor U919 (N_919,In_1680,N_653);
nor U920 (N_920,N_89,N_44);
and U921 (N_921,In_161,N_95);
xor U922 (N_922,N_239,N_159);
nor U923 (N_923,In_1083,N_12);
nand U924 (N_924,In_1334,N_205);
xnor U925 (N_925,In_1715,In_1127);
xor U926 (N_926,N_115,In_871);
or U927 (N_927,N_144,In_974);
and U928 (N_928,N_775,In_1914);
nor U929 (N_929,N_161,N_54);
nand U930 (N_930,N_504,In_382);
nor U931 (N_931,N_684,N_604);
nor U932 (N_932,N_519,In_850);
nor U933 (N_933,In_1839,N_73);
xnor U934 (N_934,N_18,In_834);
and U935 (N_935,N_796,In_1543);
or U936 (N_936,N_349,In_1788);
and U937 (N_937,N_742,N_731);
and U938 (N_938,In_1893,In_1038);
and U939 (N_939,N_109,N_596);
nand U940 (N_940,N_353,N_599);
nor U941 (N_941,N_472,N_375);
or U942 (N_942,N_24,N_764);
and U943 (N_943,In_72,In_785);
or U944 (N_944,N_481,N_307);
and U945 (N_945,N_629,N_3);
nor U946 (N_946,In_1598,In_1236);
nor U947 (N_947,In_664,N_747);
nand U948 (N_948,N_224,N_510);
nand U949 (N_949,N_799,N_659);
nor U950 (N_950,N_250,N_681);
nand U951 (N_951,In_813,In_1353);
and U952 (N_952,In_1207,N_242);
nor U953 (N_953,In_992,In_1204);
xnor U954 (N_954,N_790,In_1862);
nand U955 (N_955,N_72,N_769);
or U956 (N_956,N_645,N_576);
nand U957 (N_957,In_922,N_227);
nor U958 (N_958,N_683,In_238);
xor U959 (N_959,N_603,N_193);
nand U960 (N_960,N_778,N_401);
xnor U961 (N_961,N_70,N_571);
or U962 (N_962,In_439,N_670);
nand U963 (N_963,N_454,N_511);
nand U964 (N_964,N_419,In_743);
nand U965 (N_965,In_690,N_756);
nor U966 (N_966,N_655,In_1836);
nor U967 (N_967,N_35,In_1209);
nand U968 (N_968,In_1295,N_716);
nor U969 (N_969,N_768,N_247);
or U970 (N_970,N_658,N_578);
or U971 (N_971,N_773,N_369);
nand U972 (N_972,N_440,N_7);
nor U973 (N_973,N_782,In_872);
or U974 (N_974,N_631,N_293);
or U975 (N_975,N_395,In_508);
nor U976 (N_976,In_991,N_337);
xnor U977 (N_977,N_630,N_228);
nand U978 (N_978,In_1799,N_739);
and U979 (N_979,In_1562,N_494);
nor U980 (N_980,N_700,N_67);
and U981 (N_981,N_396,In_1273);
nor U982 (N_982,N_704,In_1257);
nor U983 (N_983,In_1262,N_332);
xor U984 (N_984,N_679,N_140);
xor U985 (N_985,N_68,N_592);
nand U986 (N_986,In_225,N_690);
or U987 (N_987,In_1613,In_906);
nand U988 (N_988,N_484,N_493);
and U989 (N_989,N_408,N_6);
and U990 (N_990,In_29,In_233);
xnor U991 (N_991,N_305,In_888);
nor U992 (N_992,N_55,N_554);
xnor U993 (N_993,N_398,In_138);
and U994 (N_994,N_500,N_453);
and U995 (N_995,In_449,N_723);
xnor U996 (N_996,N_597,In_531);
xor U997 (N_997,N_379,N_191);
or U998 (N_998,N_490,In_856);
nand U999 (N_999,In_694,N_514);
and U1000 (N_1000,N_668,N_708);
xnor U1001 (N_1001,N_794,In_593);
nor U1002 (N_1002,In_982,N_302);
xnor U1003 (N_1003,In_628,In_965);
or U1004 (N_1004,N_646,In_404);
nand U1005 (N_1005,In_1627,In_1951);
nand U1006 (N_1006,In_1616,N_2);
nor U1007 (N_1007,N_410,N_321);
and U1008 (N_1008,In_51,N_424);
nand U1009 (N_1009,N_116,In_1971);
nand U1010 (N_1010,N_518,N_287);
xor U1011 (N_1011,N_373,N_632);
nor U1012 (N_1012,N_164,In_515);
nand U1013 (N_1013,N_157,In_795);
or U1014 (N_1014,In_148,In_1457);
or U1015 (N_1015,N_317,In_202);
nand U1016 (N_1016,In_104,In_295);
nand U1017 (N_1017,N_617,N_600);
nor U1018 (N_1018,N_464,In_802);
nor U1019 (N_1019,In_1654,In_497);
nand U1020 (N_1020,In_253,N_533);
xor U1021 (N_1021,In_555,N_327);
xnor U1022 (N_1022,N_267,N_495);
or U1023 (N_1023,N_524,N_580);
or U1024 (N_1024,In_499,In_1512);
nand U1025 (N_1025,N_212,In_672);
or U1026 (N_1026,N_652,N_455);
nand U1027 (N_1027,N_475,N_167);
nand U1028 (N_1028,N_362,N_130);
or U1029 (N_1029,N_430,N_397);
nand U1030 (N_1030,In_96,In_1850);
and U1031 (N_1031,N_27,N_548);
nand U1032 (N_1032,In_1819,N_611);
nor U1033 (N_1033,N_147,N_480);
and U1034 (N_1034,In_1797,N_31);
nor U1035 (N_1035,N_78,N_313);
nand U1036 (N_1036,N_260,In_1751);
xor U1037 (N_1037,N_686,N_467);
nor U1038 (N_1038,In_1088,In_557);
nor U1039 (N_1039,In_139,N_712);
nor U1040 (N_1040,In_1869,N_20);
or U1041 (N_1041,N_491,In_1423);
nor U1042 (N_1042,N_347,N_69);
nor U1043 (N_1043,In_487,N_358);
xor U1044 (N_1044,In_1624,In_124);
or U1045 (N_1045,N_195,N_182);
nor U1046 (N_1046,N_656,N_16);
nor U1047 (N_1047,In_740,In_1567);
nand U1048 (N_1048,N_474,In_1214);
nand U1049 (N_1049,N_160,N_19);
xnor U1050 (N_1050,In_897,In_975);
xor U1051 (N_1051,N_330,In_1526);
nand U1052 (N_1052,N_774,N_382);
nor U1053 (N_1053,N_48,N_757);
and U1054 (N_1054,In_567,In_714);
or U1055 (N_1055,N_795,N_350);
xnor U1056 (N_1056,N_743,N_255);
xnor U1057 (N_1057,N_730,N_280);
and U1058 (N_1058,In_670,N_100);
or U1059 (N_1059,N_626,In_158);
and U1060 (N_1060,N_289,In_454);
or U1061 (N_1061,N_122,N_277);
or U1062 (N_1062,N_625,In_1671);
and U1063 (N_1063,N_266,In_1630);
nor U1064 (N_1064,N_240,N_751);
or U1065 (N_1065,N_117,In_248);
nand U1066 (N_1066,In_1551,N_123);
nand U1067 (N_1067,In_90,N_47);
or U1068 (N_1068,N_335,N_318);
and U1069 (N_1069,N_551,N_9);
nor U1070 (N_1070,In_1565,N_93);
and U1071 (N_1071,N_460,N_13);
nor U1072 (N_1072,In_882,N_218);
nor U1073 (N_1073,In_79,N_202);
nor U1074 (N_1074,N_81,N_64);
nor U1075 (N_1075,In_1525,In_1663);
and U1076 (N_1076,N_770,N_181);
and U1077 (N_1077,In_1646,In_1485);
and U1078 (N_1078,N_550,N_448);
nand U1079 (N_1079,In_1490,N_113);
or U1080 (N_1080,N_451,N_508);
xor U1081 (N_1081,N_384,N_780);
nand U1082 (N_1082,N_376,N_404);
or U1083 (N_1083,In_1849,N_575);
or U1084 (N_1084,N_91,N_154);
nor U1085 (N_1085,In_1373,N_590);
xnor U1086 (N_1086,N_14,N_103);
and U1087 (N_1087,In_944,N_721);
nor U1088 (N_1088,N_71,In_657);
xnor U1089 (N_1089,N_311,N_598);
nor U1090 (N_1090,In_513,N_537);
and U1091 (N_1091,N_633,N_80);
or U1092 (N_1092,In_1727,In_352);
nand U1093 (N_1093,In_1931,In_620);
nor U1094 (N_1094,N_563,N_138);
and U1095 (N_1095,N_223,N_788);
xor U1096 (N_1096,N_776,N_336);
xor U1097 (N_1097,In_1605,In_1085);
or U1098 (N_1098,N_541,In_1919);
and U1099 (N_1099,N_682,N_463);
or U1100 (N_1100,N_163,N_477);
or U1101 (N_1101,N_220,In_636);
xor U1102 (N_1102,N_346,N_614);
or U1103 (N_1103,In_858,In_971);
and U1104 (N_1104,In_480,In_1568);
or U1105 (N_1105,N_286,N_698);
nor U1106 (N_1106,In_1502,N_135);
xor U1107 (N_1107,N_388,In_1200);
xor U1108 (N_1108,N_418,In_835);
nor U1109 (N_1109,N_5,N_149);
xor U1110 (N_1110,In_1139,In_809);
and U1111 (N_1111,N_420,N_663);
nand U1112 (N_1112,N_785,N_101);
nand U1113 (N_1113,N_707,N_86);
or U1114 (N_1114,In_1130,In_820);
nor U1115 (N_1115,In_1288,N_762);
nor U1116 (N_1116,In_662,N_771);
nor U1117 (N_1117,In_1346,In_783);
nand U1118 (N_1118,N_322,N_744);
and U1119 (N_1119,In_573,N_251);
nor U1120 (N_1120,N_76,In_128);
xnor U1121 (N_1121,In_1339,N_507);
or U1122 (N_1122,N_341,N_565);
nor U1123 (N_1123,N_301,In_561);
and U1124 (N_1124,In_1,N_564);
nand U1125 (N_1125,N_634,In_1252);
nor U1126 (N_1126,N_735,N_539);
and U1127 (N_1127,N_657,N_423);
nand U1128 (N_1128,In_1197,In_1980);
nor U1129 (N_1129,In_69,N_90);
xnor U1130 (N_1130,In_1970,N_79);
nand U1131 (N_1131,N_469,In_617);
xnor U1132 (N_1132,N_180,N_763);
nand U1133 (N_1133,N_63,N_210);
xnor U1134 (N_1134,N_272,N_75);
or U1135 (N_1135,In_1391,N_219);
and U1136 (N_1136,N_344,N_249);
and U1137 (N_1137,In_224,N_526);
nand U1138 (N_1138,N_331,N_766);
and U1139 (N_1139,In_67,N_352);
or U1140 (N_1140,N_498,N_426);
nor U1141 (N_1141,In_810,N_125);
and U1142 (N_1142,In_1995,N_77);
nand U1143 (N_1143,N_797,In_950);
and U1144 (N_1144,N_40,N_165);
and U1145 (N_1145,In_98,N_236);
xnor U1146 (N_1146,In_1824,N_701);
or U1147 (N_1147,N_489,N_87);
xor U1148 (N_1148,N_749,In_1087);
xor U1149 (N_1149,N_107,N_595);
and U1150 (N_1150,N_717,N_356);
nand U1151 (N_1151,N_442,In_1561);
and U1152 (N_1152,N_363,In_1838);
nor U1153 (N_1153,N_641,N_781);
xor U1154 (N_1154,N_136,N_714);
and U1155 (N_1155,In_862,N_613);
xor U1156 (N_1156,In_1884,N_4);
and U1157 (N_1157,N_333,N_405);
xor U1158 (N_1158,N_523,N_156);
and U1159 (N_1159,N_694,N_525);
nor U1160 (N_1160,N_316,N_479);
or U1161 (N_1161,N_509,N_23);
or U1162 (N_1162,N_1,N_692);
and U1163 (N_1163,N_650,N_326);
or U1164 (N_1164,N_253,N_521);
xnor U1165 (N_1165,In_1053,N_662);
or U1166 (N_1166,N_697,N_715);
nand U1167 (N_1167,N_234,N_120);
and U1168 (N_1168,N_561,In_200);
and U1169 (N_1169,N_417,In_1482);
and U1170 (N_1170,N_471,In_1399);
and U1171 (N_1171,N_624,N_719);
or U1172 (N_1172,N_585,N_705);
and U1173 (N_1173,N_328,N_142);
or U1174 (N_1174,N_371,N_299);
nand U1175 (N_1175,In_326,N_750);
nor U1176 (N_1176,In_1447,In_1070);
nand U1177 (N_1177,N_789,N_601);
or U1178 (N_1178,N_759,N_284);
and U1179 (N_1179,N_351,N_593);
and U1180 (N_1180,N_637,In_349);
or U1181 (N_1181,In_1639,N_209);
nor U1182 (N_1182,N_37,N_582);
or U1183 (N_1183,In_1686,In_550);
nor U1184 (N_1184,N_738,N_693);
or U1185 (N_1185,N_28,In_1192);
xnor U1186 (N_1186,N_664,N_235);
and U1187 (N_1187,In_1298,N_573);
nor U1188 (N_1188,N_258,In_598);
and U1189 (N_1189,N_295,N_606);
nand U1190 (N_1190,N_237,In_1305);
or U1191 (N_1191,In_688,N_450);
xor U1192 (N_1192,N_196,N_581);
xnor U1193 (N_1193,N_137,N_0);
nand U1194 (N_1194,N_226,N_667);
nand U1195 (N_1195,N_98,N_245);
and U1196 (N_1196,N_189,In_1324);
nor U1197 (N_1197,N_452,In_643);
nor U1198 (N_1198,In_935,N_688);
or U1199 (N_1199,N_669,N_323);
nor U1200 (N_1200,In_1226,N_798);
and U1201 (N_1201,In_1745,In_172);
or U1202 (N_1202,In_441,N_643);
nor U1203 (N_1203,In_819,N_619);
or U1204 (N_1204,In_466,N_88);
and U1205 (N_1205,In_737,N_399);
nand U1206 (N_1206,N_282,In_1016);
or U1207 (N_1207,In_1250,N_52);
xor U1208 (N_1208,N_558,In_1198);
xor U1209 (N_1209,N_791,N_248);
and U1210 (N_1210,N_50,N_8);
and U1211 (N_1211,N_622,N_269);
or U1212 (N_1212,In_734,In_462);
and U1213 (N_1213,In_1386,N_288);
nand U1214 (N_1214,N_30,In_1402);
nand U1215 (N_1215,N_172,In_910);
nor U1216 (N_1216,N_124,N_203);
or U1217 (N_1217,N_665,N_213);
nand U1218 (N_1218,N_66,N_623);
or U1219 (N_1219,N_325,N_703);
or U1220 (N_1220,N_340,N_612);
nand U1221 (N_1221,N_345,N_579);
nand U1222 (N_1222,N_422,N_589);
or U1223 (N_1223,N_133,In_943);
nor U1224 (N_1224,In_237,N_534);
nand U1225 (N_1225,N_503,In_1439);
and U1226 (N_1226,N_515,N_748);
nor U1227 (N_1227,N_427,In_258);
nor U1228 (N_1228,In_1244,N_211);
and U1229 (N_1229,N_380,N_569);
or U1230 (N_1230,N_635,N_392);
nor U1231 (N_1231,N_531,In_536);
nor U1232 (N_1232,N_82,N_737);
or U1233 (N_1233,In_1628,In_625);
or U1234 (N_1234,N_677,N_687);
xnor U1235 (N_1235,N_752,In_1507);
xor U1236 (N_1236,N_162,N_309);
and U1237 (N_1237,N_496,In_293);
or U1238 (N_1238,In_1142,In_1075);
or U1239 (N_1239,In_390,N_276);
or U1240 (N_1240,N_92,N_647);
or U1241 (N_1241,N_651,N_312);
or U1242 (N_1242,N_793,N_458);
xnor U1243 (N_1243,In_106,N_547);
nor U1244 (N_1244,N_383,In_1413);
nor U1245 (N_1245,N_273,N_615);
and U1246 (N_1246,N_709,N_56);
nor U1247 (N_1247,N_178,N_21);
and U1248 (N_1248,N_546,N_765);
and U1249 (N_1249,In_1320,N_706);
nor U1250 (N_1250,In_889,In_1890);
nor U1251 (N_1251,In_1908,N_278);
nor U1252 (N_1252,N_772,In_886);
and U1253 (N_1253,N_185,In_1171);
nand U1254 (N_1254,In_1532,N_535);
and U1255 (N_1255,N_447,N_292);
and U1256 (N_1256,N_233,In_1652);
or U1257 (N_1257,N_609,In_52);
xnor U1258 (N_1258,In_471,In_667);
nor U1259 (N_1259,N_520,N_587);
nand U1260 (N_1260,N_436,In_1683);
or U1261 (N_1261,In_1140,N_588);
or U1262 (N_1262,N_466,N_206);
nand U1263 (N_1263,N_372,In_1540);
nor U1264 (N_1264,N_296,In_1109);
nand U1265 (N_1265,N_726,N_150);
nor U1266 (N_1266,N_699,N_83);
xor U1267 (N_1267,N_230,In_1584);
xor U1268 (N_1268,N_146,In_604);
or U1269 (N_1269,N_733,N_691);
or U1270 (N_1270,N_728,N_675);
or U1271 (N_1271,In_699,N_627);
nor U1272 (N_1272,N_264,N_29);
xor U1273 (N_1273,In_786,N_229);
and U1274 (N_1274,In_976,In_552);
nor U1275 (N_1275,N_654,N_530);
nand U1276 (N_1276,In_979,In_692);
and U1277 (N_1277,N_502,N_499);
xor U1278 (N_1278,N_640,N_127);
and U1279 (N_1279,N_512,In_1047);
or U1280 (N_1280,N_660,N_119);
and U1281 (N_1281,N_608,N_308);
nor U1282 (N_1282,N_306,N_179);
nand U1283 (N_1283,In_1231,N_722);
or U1284 (N_1284,N_517,N_552);
nand U1285 (N_1285,N_170,In_1419);
nor U1286 (N_1286,N_141,In_553);
xnor U1287 (N_1287,N_232,N_437);
and U1288 (N_1288,In_1790,In_1377);
nand U1289 (N_1289,In_1401,N_607);
nor U1290 (N_1290,N_152,N_129);
and U1291 (N_1291,In_102,N_104);
xnor U1292 (N_1292,N_536,N_186);
xnor U1293 (N_1293,N_678,In_673);
or U1294 (N_1294,In_983,In_64);
and U1295 (N_1295,N_387,N_314);
and U1296 (N_1296,N_745,N_391);
xnor U1297 (N_1297,In_1182,N_586);
and U1298 (N_1298,In_931,N_168);
xnor U1299 (N_1299,In_1957,In_1220);
nand U1300 (N_1300,In_455,N_407);
and U1301 (N_1301,N_583,N_108);
nor U1302 (N_1302,In_677,N_754);
and U1303 (N_1303,N_354,In_437);
and U1304 (N_1304,N_428,In_1612);
nor U1305 (N_1305,N_370,In_1992);
and U1306 (N_1306,N_58,N_394);
nand U1307 (N_1307,N_201,N_610);
xnor U1308 (N_1308,In_1942,In_207);
or U1309 (N_1309,In_252,In_642);
nand U1310 (N_1310,In_60,N_275);
nand U1311 (N_1311,N_177,In_334);
and U1312 (N_1312,N_102,N_315);
xor U1313 (N_1313,N_412,N_367);
xnor U1314 (N_1314,In_1468,N_271);
nor U1315 (N_1315,N_297,N_486);
nor U1316 (N_1316,N_505,N_118);
or U1317 (N_1317,In_115,N_431);
and U1318 (N_1318,N_15,N_476);
nand U1319 (N_1319,N_761,N_553);
and U1320 (N_1320,N_22,N_522);
or U1321 (N_1321,N_544,N_262);
xor U1322 (N_1322,N_263,In_1011);
nor U1323 (N_1323,N_105,N_197);
xor U1324 (N_1324,In_1547,N_155);
nand U1325 (N_1325,In_1591,In_1615);
and U1326 (N_1326,N_478,N_620);
and U1327 (N_1327,N_279,N_488);
and U1328 (N_1328,In_1601,N_516);
and U1329 (N_1329,N_644,N_648);
nand U1330 (N_1330,N_132,In_1425);
nor U1331 (N_1331,N_435,N_746);
xnor U1332 (N_1332,In_432,N_34);
xnor U1333 (N_1333,N_381,N_727);
nand U1334 (N_1334,N_557,N_638);
or U1335 (N_1335,In_1622,In_1535);
nor U1336 (N_1336,In_144,N_222);
or U1337 (N_1337,In_176,In_1474);
and U1338 (N_1338,N_415,N_378);
or U1339 (N_1339,N_529,N_368);
or U1340 (N_1340,N_217,In_427);
xnor U1341 (N_1341,N_303,N_540);
nor U1342 (N_1342,N_329,N_385);
xnor U1343 (N_1343,N_153,N_736);
and U1344 (N_1344,In_131,N_485);
xor U1345 (N_1345,N_324,In_1094);
and U1346 (N_1346,In_275,In_132);
or U1347 (N_1347,In_696,N_268);
and U1348 (N_1348,N_166,N_57);
or U1349 (N_1349,N_365,N_432);
and U1350 (N_1350,N_298,N_244);
or U1351 (N_1351,N_374,N_53);
xnor U1352 (N_1352,N_513,N_492);
nor U1353 (N_1353,N_753,In_368);
or U1354 (N_1354,N_151,In_1375);
xor U1355 (N_1355,N_334,In_1255);
nor U1356 (N_1356,N_636,In_1213);
xnor U1357 (N_1357,In_1665,N_457);
xor U1358 (N_1358,In_209,In_1911);
and U1359 (N_1359,N_339,In_347);
and U1360 (N_1360,N_425,In_763);
nor U1361 (N_1361,N_685,N_577);
nand U1362 (N_1362,N_445,In_619);
and U1363 (N_1363,N_786,In_1664);
xor U1364 (N_1364,In_1025,N_545);
and U1365 (N_1365,In_842,N_672);
xnor U1366 (N_1366,N_221,N_256);
nand U1367 (N_1367,N_357,N_543);
and U1368 (N_1368,In_370,N_462);
xnor U1369 (N_1369,N_591,N_661);
nor U1370 (N_1370,In_715,In_1780);
nor U1371 (N_1371,In_339,In_1801);
xor U1372 (N_1372,N_566,N_94);
or U1373 (N_1373,N_400,In_1191);
and U1374 (N_1374,N_32,In_602);
nand U1375 (N_1375,N_402,N_36);
nand U1376 (N_1376,N_45,N_51);
nand U1377 (N_1377,In_707,In_1832);
nor U1378 (N_1378,N_265,N_787);
nor U1379 (N_1379,N_760,N_527);
xor U1380 (N_1380,N_359,In_946);
nor U1381 (N_1381,In_961,In_634);
and U1382 (N_1382,N_618,N_59);
or U1383 (N_1383,N_555,N_281);
or U1384 (N_1384,N_449,N_121);
or U1385 (N_1385,N_570,In_653);
or U1386 (N_1386,N_444,In_13);
or U1387 (N_1387,In_1668,In_319);
or U1388 (N_1388,N_49,N_439);
and U1389 (N_1389,N_65,In_681);
and U1390 (N_1390,In_1300,In_457);
nor U1391 (N_1391,N_96,N_695);
and U1392 (N_1392,In_905,In_1508);
nand U1393 (N_1393,N_783,N_143);
xor U1394 (N_1394,N_456,N_567);
and U1395 (N_1395,In_197,N_246);
xnor U1396 (N_1396,N_574,In_312);
or U1397 (N_1397,In_663,In_1766);
or U1398 (N_1398,In_183,N_106);
nand U1399 (N_1399,N_274,N_300);
nand U1400 (N_1400,N_350,N_283);
or U1401 (N_1401,N_94,N_354);
or U1402 (N_1402,N_13,In_96);
or U1403 (N_1403,In_370,N_88);
nand U1404 (N_1404,N_645,N_725);
xor U1405 (N_1405,In_1586,N_390);
and U1406 (N_1406,N_611,N_510);
and U1407 (N_1407,N_364,N_58);
or U1408 (N_1408,N_342,N_490);
nand U1409 (N_1409,N_764,In_642);
or U1410 (N_1410,N_411,N_735);
xor U1411 (N_1411,N_417,In_1385);
or U1412 (N_1412,In_1686,N_748);
and U1413 (N_1413,N_687,N_333);
nor U1414 (N_1414,In_1565,N_471);
or U1415 (N_1415,In_604,N_735);
nor U1416 (N_1416,In_497,N_397);
nand U1417 (N_1417,N_660,N_495);
nor U1418 (N_1418,N_250,N_391);
and U1419 (N_1419,In_1613,N_402);
and U1420 (N_1420,N_62,N_185);
or U1421 (N_1421,In_1593,In_1919);
and U1422 (N_1422,In_1198,In_1862);
or U1423 (N_1423,In_383,In_1838);
xor U1424 (N_1424,N_676,In_714);
nor U1425 (N_1425,N_644,N_194);
nand U1426 (N_1426,N_695,In_90);
and U1427 (N_1427,In_1665,N_362);
nand U1428 (N_1428,N_339,In_349);
or U1429 (N_1429,N_557,N_446);
or U1430 (N_1430,N_531,N_243);
xnor U1431 (N_1431,In_293,In_1797);
xnor U1432 (N_1432,In_69,N_156);
nand U1433 (N_1433,In_1839,N_435);
nand U1434 (N_1434,N_348,N_512);
nor U1435 (N_1435,N_575,N_694);
nand U1436 (N_1436,N_497,N_396);
xor U1437 (N_1437,N_620,N_475);
nand U1438 (N_1438,N_758,In_1712);
or U1439 (N_1439,In_1401,N_299);
or U1440 (N_1440,N_385,N_670);
xor U1441 (N_1441,N_487,N_767);
nand U1442 (N_1442,N_426,In_1011);
xor U1443 (N_1443,N_256,In_1507);
nand U1444 (N_1444,N_182,In_1257);
xor U1445 (N_1445,N_223,N_127);
nand U1446 (N_1446,N_81,N_495);
nand U1447 (N_1447,N_690,In_462);
nand U1448 (N_1448,N_500,N_198);
or U1449 (N_1449,In_275,In_326);
or U1450 (N_1450,N_124,N_799);
xnor U1451 (N_1451,N_382,N_283);
nand U1452 (N_1452,N_694,In_1791);
nor U1453 (N_1453,In_1324,N_45);
xnor U1454 (N_1454,N_771,In_1757);
xor U1455 (N_1455,N_583,N_546);
and U1456 (N_1456,In_653,In_1339);
and U1457 (N_1457,N_650,N_193);
or U1458 (N_1458,N_773,N_574);
and U1459 (N_1459,In_1025,N_162);
nor U1460 (N_1460,N_237,N_788);
and U1461 (N_1461,N_174,N_469);
xnor U1462 (N_1462,N_415,N_604);
nand U1463 (N_1463,In_1627,N_289);
or U1464 (N_1464,N_103,N_380);
nand U1465 (N_1465,N_417,N_324);
nor U1466 (N_1466,In_888,In_1911);
nand U1467 (N_1467,In_906,In_471);
or U1468 (N_1468,In_672,N_21);
and U1469 (N_1469,N_67,In_1745);
xor U1470 (N_1470,N_569,In_148);
nand U1471 (N_1471,N_441,In_427);
xor U1472 (N_1472,In_1799,N_202);
nand U1473 (N_1473,N_54,N_53);
xnor U1474 (N_1474,N_304,In_946);
and U1475 (N_1475,N_246,N_700);
or U1476 (N_1476,N_470,In_1022);
nor U1477 (N_1477,N_194,N_540);
xnor U1478 (N_1478,N_315,N_769);
nand U1479 (N_1479,N_384,In_1801);
nor U1480 (N_1480,N_650,In_1320);
and U1481 (N_1481,In_931,N_605);
and U1482 (N_1482,N_46,N_113);
nand U1483 (N_1483,N_562,N_778);
nand U1484 (N_1484,N_520,In_943);
xor U1485 (N_1485,N_365,In_1707);
nand U1486 (N_1486,In_1801,N_246);
nand U1487 (N_1487,N_551,N_290);
xnor U1488 (N_1488,In_383,N_128);
nand U1489 (N_1489,N_794,N_70);
or U1490 (N_1490,N_705,N_0);
xor U1491 (N_1491,N_133,In_1790);
xnor U1492 (N_1492,In_1525,N_610);
and U1493 (N_1493,In_439,N_157);
xnor U1494 (N_1494,In_1011,N_349);
or U1495 (N_1495,N_452,N_631);
or U1496 (N_1496,N_591,In_620);
xnor U1497 (N_1497,In_1914,In_1033);
and U1498 (N_1498,N_778,N_44);
and U1499 (N_1499,N_541,N_281);
nand U1500 (N_1500,N_660,N_792);
nor U1501 (N_1501,N_418,N_57);
and U1502 (N_1502,N_429,N_387);
nor U1503 (N_1503,N_603,In_544);
xor U1504 (N_1504,In_1485,N_645);
and U1505 (N_1505,In_1584,N_32);
nor U1506 (N_1506,N_351,N_142);
and U1507 (N_1507,In_1957,In_1605);
or U1508 (N_1508,N_677,N_421);
or U1509 (N_1509,N_271,N_454);
or U1510 (N_1510,In_1334,N_311);
nand U1511 (N_1511,In_491,N_399);
nor U1512 (N_1512,N_402,N_296);
xnor U1513 (N_1513,N_760,In_992);
and U1514 (N_1514,N_179,N_405);
xor U1515 (N_1515,In_1008,N_629);
or U1516 (N_1516,In_248,In_550);
or U1517 (N_1517,In_1401,N_55);
nor U1518 (N_1518,N_272,N_646);
nor U1519 (N_1519,N_527,N_337);
and U1520 (N_1520,N_53,N_311);
and U1521 (N_1521,In_432,In_1893);
xor U1522 (N_1522,In_922,N_659);
nand U1523 (N_1523,N_93,In_1680);
nand U1524 (N_1524,N_193,In_1226);
nand U1525 (N_1525,N_37,N_359);
or U1526 (N_1526,N_574,N_625);
nor U1527 (N_1527,N_2,N_499);
xor U1528 (N_1528,In_819,In_1033);
nor U1529 (N_1529,N_754,N_500);
nand U1530 (N_1530,N_433,N_186);
xnor U1531 (N_1531,N_502,N_336);
and U1532 (N_1532,N_429,In_1766);
xnor U1533 (N_1533,In_176,N_626);
nand U1534 (N_1534,N_136,N_396);
xnor U1535 (N_1535,N_304,N_397);
nand U1536 (N_1536,N_25,N_210);
or U1537 (N_1537,N_119,N_747);
or U1538 (N_1538,N_142,N_474);
nand U1539 (N_1539,N_119,N_438);
and U1540 (N_1540,N_364,N_85);
nand U1541 (N_1541,N_612,In_1908);
xor U1542 (N_1542,In_971,N_501);
nand U1543 (N_1543,N_371,N_556);
nand U1544 (N_1544,In_72,N_718);
nor U1545 (N_1545,In_763,N_3);
xor U1546 (N_1546,N_70,N_237);
nand U1547 (N_1547,N_680,N_195);
or U1548 (N_1548,In_692,N_128);
or U1549 (N_1549,In_237,N_265);
or U1550 (N_1550,In_13,N_496);
or U1551 (N_1551,N_618,N_653);
nand U1552 (N_1552,N_472,N_730);
nand U1553 (N_1553,In_1127,In_1413);
nor U1554 (N_1554,In_634,N_353);
nor U1555 (N_1555,N_616,N_385);
or U1556 (N_1556,In_200,N_491);
and U1557 (N_1557,N_114,N_37);
xnor U1558 (N_1558,N_83,N_454);
nor U1559 (N_1559,N_194,N_179);
and U1560 (N_1560,N_420,N_683);
or U1561 (N_1561,N_416,In_462);
nand U1562 (N_1562,N_549,In_1565);
or U1563 (N_1563,N_139,In_991);
xnor U1564 (N_1564,N_360,N_645);
nor U1565 (N_1565,N_736,N_740);
nand U1566 (N_1566,In_842,N_784);
nand U1567 (N_1567,N_421,N_714);
and U1568 (N_1568,N_612,N_519);
nand U1569 (N_1569,In_842,N_321);
nor U1570 (N_1570,N_679,N_629);
or U1571 (N_1571,N_496,N_312);
nand U1572 (N_1572,In_1244,N_129);
and U1573 (N_1573,N_217,N_297);
and U1574 (N_1574,N_191,In_653);
nor U1575 (N_1575,N_578,N_369);
nand U1576 (N_1576,In_1970,N_613);
nor U1577 (N_1577,In_1707,N_614);
xor U1578 (N_1578,N_788,N_58);
and U1579 (N_1579,N_776,N_376);
xor U1580 (N_1580,N_266,In_1305);
xor U1581 (N_1581,In_98,N_83);
or U1582 (N_1582,N_214,N_784);
nand U1583 (N_1583,N_784,N_735);
and U1584 (N_1584,N_322,In_677);
nor U1585 (N_1585,N_6,In_102);
xor U1586 (N_1586,N_665,N_74);
or U1587 (N_1587,In_1262,In_1646);
nand U1588 (N_1588,In_326,N_169);
nor U1589 (N_1589,N_344,N_74);
xor U1590 (N_1590,In_557,N_476);
and U1591 (N_1591,In_888,In_1584);
nor U1592 (N_1592,In_783,In_439);
nand U1593 (N_1593,N_756,N_28);
nor U1594 (N_1594,In_946,N_412);
and U1595 (N_1595,N_351,N_330);
and U1596 (N_1596,N_661,In_1715);
and U1597 (N_1597,N_134,In_1020);
nand U1598 (N_1598,N_777,In_228);
or U1599 (N_1599,N_232,N_678);
and U1600 (N_1600,N_1039,N_835);
nand U1601 (N_1601,N_1420,N_1129);
nand U1602 (N_1602,N_1574,N_1109);
xnor U1603 (N_1603,N_1245,N_1440);
or U1604 (N_1604,N_1230,N_963);
nand U1605 (N_1605,N_1155,N_1032);
nand U1606 (N_1606,N_810,N_1120);
or U1607 (N_1607,N_1392,N_1436);
xor U1608 (N_1608,N_1591,N_1412);
nor U1609 (N_1609,N_813,N_1215);
xor U1610 (N_1610,N_1486,N_1240);
or U1611 (N_1611,N_1564,N_1006);
and U1612 (N_1612,N_1345,N_1449);
nand U1613 (N_1613,N_1547,N_1121);
xor U1614 (N_1614,N_1361,N_1333);
nand U1615 (N_1615,N_816,N_1551);
xor U1616 (N_1616,N_1188,N_1369);
nor U1617 (N_1617,N_1115,N_1335);
nand U1618 (N_1618,N_1183,N_979);
nand U1619 (N_1619,N_968,N_971);
nand U1620 (N_1620,N_1062,N_1445);
or U1621 (N_1621,N_966,N_931);
or U1622 (N_1622,N_1527,N_1171);
xor U1623 (N_1623,N_826,N_887);
xnor U1624 (N_1624,N_1516,N_1057);
and U1625 (N_1625,N_1279,N_1541);
xor U1626 (N_1626,N_1487,N_1016);
nor U1627 (N_1627,N_1566,N_1572);
and U1628 (N_1628,N_881,N_1110);
xnor U1629 (N_1629,N_1242,N_877);
or U1630 (N_1630,N_1148,N_1071);
nor U1631 (N_1631,N_1139,N_1151);
nand U1632 (N_1632,N_883,N_875);
nor U1633 (N_1633,N_1145,N_1446);
nor U1634 (N_1634,N_1315,N_1273);
nand U1635 (N_1635,N_1167,N_1508);
xnor U1636 (N_1636,N_1521,N_1176);
and U1637 (N_1637,N_1321,N_822);
or U1638 (N_1638,N_1237,N_1530);
nand U1639 (N_1639,N_1403,N_1316);
xnor U1640 (N_1640,N_1443,N_1222);
or U1641 (N_1641,N_1178,N_1571);
or U1642 (N_1642,N_1543,N_1209);
or U1643 (N_1643,N_1568,N_1424);
xnor U1644 (N_1644,N_1320,N_1428);
and U1645 (N_1645,N_1563,N_1134);
or U1646 (N_1646,N_1448,N_1002);
and U1647 (N_1647,N_1219,N_1042);
xnor U1648 (N_1648,N_1096,N_836);
nand U1649 (N_1649,N_871,N_969);
nand U1650 (N_1650,N_1437,N_1444);
nand U1651 (N_1651,N_1341,N_950);
or U1652 (N_1652,N_1282,N_806);
xnor U1653 (N_1653,N_1373,N_874);
xor U1654 (N_1654,N_1101,N_956);
and U1655 (N_1655,N_1291,N_1138);
nor U1656 (N_1656,N_1463,N_891);
or U1657 (N_1657,N_1146,N_1290);
nand U1658 (N_1658,N_1498,N_833);
xnor U1659 (N_1659,N_1458,N_909);
xor U1660 (N_1660,N_985,N_1575);
nor U1661 (N_1661,N_1475,N_1493);
nor U1662 (N_1662,N_1308,N_1106);
and U1663 (N_1663,N_890,N_1506);
and U1664 (N_1664,N_1413,N_1131);
xor U1665 (N_1665,N_975,N_1266);
xor U1666 (N_1666,N_1218,N_1092);
and U1667 (N_1667,N_1348,N_1077);
nor U1668 (N_1668,N_869,N_1268);
and U1669 (N_1669,N_1388,N_1525);
nand U1670 (N_1670,N_1011,N_1267);
nor U1671 (N_1671,N_1081,N_1231);
nor U1672 (N_1672,N_957,N_999);
or U1673 (N_1673,N_866,N_862);
and U1674 (N_1674,N_937,N_953);
and U1675 (N_1675,N_1075,N_1037);
nor U1676 (N_1676,N_853,N_1358);
nand U1677 (N_1677,N_1125,N_1089);
nand U1678 (N_1678,N_1597,N_1422);
nand U1679 (N_1679,N_1326,N_807);
and U1680 (N_1680,N_1269,N_1324);
nor U1681 (N_1681,N_1022,N_1073);
xnor U1682 (N_1682,N_1334,N_1226);
nand U1683 (N_1683,N_1085,N_834);
nand U1684 (N_1684,N_1154,N_1312);
nor U1685 (N_1685,N_1189,N_818);
and U1686 (N_1686,N_1123,N_908);
xnor U1687 (N_1687,N_1492,N_1586);
and U1688 (N_1688,N_1205,N_947);
and U1689 (N_1689,N_1452,N_1046);
nand U1690 (N_1690,N_1313,N_828);
nand U1691 (N_1691,N_1397,N_1304);
nand U1692 (N_1692,N_839,N_885);
xnor U1693 (N_1693,N_965,N_1009);
nor U1694 (N_1694,N_815,N_1410);
and U1695 (N_1695,N_1459,N_1367);
xnor U1696 (N_1696,N_1052,N_1264);
or U1697 (N_1697,N_1191,N_1133);
xnor U1698 (N_1698,N_992,N_1441);
and U1699 (N_1699,N_1224,N_1434);
or U1700 (N_1700,N_1284,N_1535);
nand U1701 (N_1701,N_1285,N_1514);
nand U1702 (N_1702,N_1490,N_990);
or U1703 (N_1703,N_1466,N_867);
or U1704 (N_1704,N_1108,N_856);
or U1705 (N_1705,N_1587,N_1599);
and U1706 (N_1706,N_811,N_1309);
and U1707 (N_1707,N_872,N_1534);
nor U1708 (N_1708,N_1286,N_1462);
or U1709 (N_1709,N_1461,N_1589);
nand U1710 (N_1710,N_1518,N_1233);
or U1711 (N_1711,N_1501,N_1254);
nand U1712 (N_1712,N_1540,N_845);
nand U1713 (N_1713,N_805,N_1318);
nor U1714 (N_1714,N_1287,N_1142);
or U1715 (N_1715,N_1064,N_944);
nor U1716 (N_1716,N_1179,N_889);
nand U1717 (N_1717,N_1225,N_1074);
nand U1718 (N_1718,N_1280,N_1206);
xor U1719 (N_1719,N_1132,N_1387);
nor U1720 (N_1720,N_1402,N_951);
or U1721 (N_1721,N_1473,N_1031);
nand U1722 (N_1722,N_972,N_1447);
nand U1723 (N_1723,N_1578,N_1338);
and U1724 (N_1724,N_1210,N_840);
nor U1725 (N_1725,N_1303,N_1430);
xor U1726 (N_1726,N_1033,N_1378);
or U1727 (N_1727,N_838,N_1519);
or U1728 (N_1728,N_1433,N_981);
xor U1729 (N_1729,N_1295,N_1281);
nor U1730 (N_1730,N_893,N_1405);
nor U1731 (N_1731,N_1349,N_1272);
xnor U1732 (N_1732,N_913,N_1474);
or U1733 (N_1733,N_1024,N_1152);
or U1734 (N_1734,N_1255,N_857);
xor U1735 (N_1735,N_1160,N_1478);
or U1736 (N_1736,N_1013,N_1066);
xnor U1737 (N_1737,N_1329,N_1300);
and U1738 (N_1738,N_939,N_1485);
nor U1739 (N_1739,N_1552,N_1336);
nand U1740 (N_1740,N_1107,N_960);
xnor U1741 (N_1741,N_1330,N_1112);
nor U1742 (N_1742,N_932,N_1435);
xnor U1743 (N_1743,N_1021,N_1292);
nor U1744 (N_1744,N_922,N_1169);
nand U1745 (N_1745,N_830,N_1327);
and U1746 (N_1746,N_1213,N_1034);
xnor U1747 (N_1747,N_1208,N_1400);
nor U1748 (N_1748,N_1418,N_1542);
xor U1749 (N_1749,N_1298,N_1451);
or U1750 (N_1750,N_1407,N_1078);
and U1751 (N_1751,N_1510,N_1256);
or U1752 (N_1752,N_1122,N_1027);
nor U1753 (N_1753,N_912,N_1584);
xnor U1754 (N_1754,N_1246,N_850);
xor U1755 (N_1755,N_1372,N_1271);
xnor U1756 (N_1756,N_879,N_829);
nand U1757 (N_1757,N_858,N_1135);
or U1758 (N_1758,N_911,N_1425);
nor U1759 (N_1759,N_1035,N_1211);
or U1760 (N_1760,N_1481,N_1217);
and U1761 (N_1761,N_1414,N_1576);
nand U1762 (N_1762,N_846,N_1140);
and U1763 (N_1763,N_1194,N_1370);
and U1764 (N_1764,N_1340,N_1590);
xor U1765 (N_1765,N_855,N_1374);
and U1766 (N_1766,N_1247,N_1323);
nor U1767 (N_1767,N_1043,N_989);
nand U1768 (N_1768,N_832,N_1394);
nor U1769 (N_1769,N_1366,N_1343);
or U1770 (N_1770,N_914,N_1162);
and U1771 (N_1771,N_986,N_1310);
xor U1772 (N_1772,N_1117,N_1150);
xnor U1773 (N_1773,N_1427,N_1297);
nand U1774 (N_1774,N_1362,N_1003);
or U1775 (N_1775,N_928,N_1393);
nor U1776 (N_1776,N_1357,N_1221);
nor U1777 (N_1777,N_1328,N_1149);
and U1778 (N_1778,N_1235,N_1517);
nand U1779 (N_1779,N_1509,N_1168);
and U1780 (N_1780,N_1356,N_924);
and U1781 (N_1781,N_1382,N_854);
nand U1782 (N_1782,N_1099,N_1229);
or U1783 (N_1783,N_895,N_1293);
and U1784 (N_1784,N_1124,N_1248);
nor U1785 (N_1785,N_994,N_1094);
nand U1786 (N_1786,N_1082,N_1198);
and U1787 (N_1787,N_842,N_1084);
nor U1788 (N_1788,N_1128,N_1539);
nand U1789 (N_1789,N_1594,N_852);
or U1790 (N_1790,N_1438,N_1396);
nand U1791 (N_1791,N_1456,N_1522);
or U1792 (N_1792,N_925,N_970);
or U1793 (N_1793,N_1265,N_1197);
and U1794 (N_1794,N_917,N_1192);
and U1795 (N_1795,N_1018,N_1243);
or U1796 (N_1796,N_915,N_1331);
and U1797 (N_1797,N_1058,N_1214);
nand U1798 (N_1798,N_1137,N_896);
and U1799 (N_1799,N_1536,N_1172);
xnor U1800 (N_1800,N_1480,N_1008);
and U1801 (N_1801,N_906,N_1180);
or U1802 (N_1802,N_1274,N_1581);
xor U1803 (N_1803,N_1143,N_1283);
xnor U1804 (N_1804,N_1000,N_1472);
xnor U1805 (N_1805,N_1431,N_1147);
or U1806 (N_1806,N_1070,N_1524);
or U1807 (N_1807,N_1098,N_1439);
and U1808 (N_1808,N_1177,N_1296);
and U1809 (N_1809,N_821,N_1464);
and U1810 (N_1810,N_997,N_1352);
and U1811 (N_1811,N_1558,N_907);
nand U1812 (N_1812,N_802,N_1004);
and U1813 (N_1813,N_1093,N_1241);
xor U1814 (N_1814,N_1411,N_897);
and U1815 (N_1815,N_1158,N_940);
xor U1816 (N_1816,N_894,N_809);
and U1817 (N_1817,N_1555,N_942);
and U1818 (N_1818,N_1068,N_935);
and U1819 (N_1819,N_1363,N_1546);
xnor U1820 (N_1820,N_1409,N_1469);
nor U1821 (N_1821,N_1565,N_886);
or U1822 (N_1822,N_1127,N_949);
and U1823 (N_1823,N_1398,N_1442);
nand U1824 (N_1824,N_1550,N_1342);
and U1825 (N_1825,N_1100,N_1570);
xor U1826 (N_1826,N_1041,N_977);
or U1827 (N_1827,N_1030,N_1025);
nor U1828 (N_1828,N_1216,N_1561);
xor U1829 (N_1829,N_1260,N_870);
xnor U1830 (N_1830,N_1088,N_1061);
nand U1831 (N_1831,N_1259,N_1454);
xnor U1832 (N_1832,N_982,N_878);
and U1833 (N_1833,N_1317,N_976);
or U1834 (N_1834,N_1090,N_921);
or U1835 (N_1835,N_1505,N_1429);
nand U1836 (N_1836,N_1353,N_1588);
xor U1837 (N_1837,N_1484,N_1060);
nand U1838 (N_1838,N_988,N_1116);
or U1839 (N_1839,N_1250,N_1212);
nand U1840 (N_1840,N_927,N_1350);
or U1841 (N_1841,N_1175,N_843);
nor U1842 (N_1842,N_1419,N_1306);
xnor U1843 (N_1843,N_1360,N_800);
or U1844 (N_1844,N_801,N_1028);
or U1845 (N_1845,N_959,N_1499);
or U1846 (N_1846,N_1063,N_1562);
nand U1847 (N_1847,N_1095,N_1253);
xor U1848 (N_1848,N_1347,N_1174);
xnor U1849 (N_1849,N_1488,N_1423);
and U1850 (N_1850,N_903,N_861);
nand U1851 (N_1851,N_1526,N_945);
or U1852 (N_1852,N_868,N_1453);
or U1853 (N_1853,N_1497,N_1079);
and U1854 (N_1854,N_1513,N_923);
nand U1855 (N_1855,N_1426,N_1165);
xor U1856 (N_1856,N_1386,N_1007);
nor U1857 (N_1857,N_1126,N_1119);
or U1858 (N_1858,N_1585,N_1166);
nor U1859 (N_1859,N_1005,N_1163);
or U1860 (N_1860,N_978,N_1053);
nand U1861 (N_1861,N_1252,N_1385);
nor U1862 (N_1862,N_1406,N_1470);
nor U1863 (N_1863,N_1038,N_1118);
and U1864 (N_1864,N_991,N_948);
nand U1865 (N_1865,N_1170,N_902);
xor U1866 (N_1866,N_1544,N_1311);
xor U1867 (N_1867,N_1579,N_1153);
nor U1868 (N_1868,N_1500,N_1019);
xor U1869 (N_1869,N_1346,N_1087);
or U1870 (N_1870,N_954,N_920);
or U1871 (N_1871,N_955,N_933);
nor U1872 (N_1872,N_1190,N_1036);
or U1873 (N_1873,N_1220,N_1261);
or U1874 (N_1874,N_1054,N_1528);
nor U1875 (N_1875,N_1389,N_1538);
xor U1876 (N_1876,N_1263,N_1047);
nor U1877 (N_1877,N_1258,N_1017);
nand U1878 (N_1878,N_1379,N_1023);
nor U1879 (N_1879,N_1332,N_1489);
nor U1880 (N_1880,N_930,N_1529);
nor U1881 (N_1881,N_1593,N_1399);
xor U1882 (N_1882,N_1104,N_1365);
xnor U1883 (N_1883,N_1111,N_1202);
xnor U1884 (N_1884,N_1548,N_863);
nor U1885 (N_1885,N_888,N_1523);
and U1886 (N_1886,N_1020,N_1583);
xor U1887 (N_1887,N_1236,N_827);
xnor U1888 (N_1888,N_1314,N_1598);
nand U1889 (N_1889,N_1344,N_1181);
xor U1890 (N_1890,N_1432,N_1200);
nor U1891 (N_1891,N_803,N_1204);
and U1892 (N_1892,N_980,N_1199);
and U1893 (N_1893,N_1503,N_1299);
or U1894 (N_1894,N_1375,N_1460);
or U1895 (N_1895,N_1537,N_1186);
nor U1896 (N_1896,N_1161,N_1390);
nor U1897 (N_1897,N_1069,N_1185);
nand U1898 (N_1898,N_824,N_1187);
nor U1899 (N_1899,N_814,N_831);
xnor U1900 (N_1900,N_1026,N_819);
xor U1901 (N_1901,N_1065,N_918);
nor U1902 (N_1902,N_1559,N_1319);
xnor U1903 (N_1903,N_1351,N_1195);
xnor U1904 (N_1904,N_967,N_926);
and U1905 (N_1905,N_1048,N_1322);
xor U1906 (N_1906,N_1483,N_1244);
and U1907 (N_1907,N_1278,N_973);
nand U1908 (N_1908,N_958,N_983);
or U1909 (N_1909,N_1288,N_1238);
nor U1910 (N_1910,N_1044,N_1495);
or U1911 (N_1911,N_1228,N_880);
and U1912 (N_1912,N_1595,N_864);
and U1913 (N_1913,N_1376,N_820);
nand U1914 (N_1914,N_892,N_1457);
nand U1915 (N_1915,N_1086,N_808);
nor U1916 (N_1916,N_1339,N_905);
nor U1917 (N_1917,N_1049,N_812);
nand U1918 (N_1918,N_1029,N_1182);
and U1919 (N_1919,N_1582,N_1476);
xnor U1920 (N_1920,N_1479,N_1533);
and U1921 (N_1921,N_1381,N_901);
nor U1922 (N_1922,N_1289,N_1553);
nor U1923 (N_1923,N_1421,N_1203);
or U1924 (N_1924,N_1091,N_882);
and U1925 (N_1925,N_938,N_1196);
and U1926 (N_1926,N_1257,N_1223);
nor U1927 (N_1927,N_1144,N_1383);
or U1928 (N_1928,N_847,N_865);
and U1929 (N_1929,N_1502,N_946);
xnor U1930 (N_1930,N_876,N_1251);
nor U1931 (N_1931,N_1401,N_984);
xor U1932 (N_1932,N_1141,N_1051);
nand U1933 (N_1933,N_987,N_1468);
or U1934 (N_1934,N_929,N_1371);
xor U1935 (N_1935,N_1416,N_1294);
or U1936 (N_1936,N_1249,N_1050);
and U1937 (N_1937,N_1159,N_995);
nor U1938 (N_1938,N_1477,N_1384);
and U1939 (N_1939,N_1055,N_898);
nor U1940 (N_1940,N_934,N_1368);
xnor U1941 (N_1941,N_1302,N_1105);
or U1942 (N_1942,N_1201,N_1377);
xnor U1943 (N_1943,N_1232,N_1515);
nor U1944 (N_1944,N_1337,N_1450);
nor U1945 (N_1945,N_1262,N_1097);
nor U1946 (N_1946,N_1395,N_1560);
nand U1947 (N_1947,N_1083,N_1415);
and U1948 (N_1948,N_1270,N_1080);
and U1949 (N_1949,N_1404,N_1102);
nand U1950 (N_1950,N_1072,N_1482);
xnor U1951 (N_1951,N_1059,N_859);
or U1952 (N_1952,N_1491,N_1554);
nor U1953 (N_1953,N_1157,N_996);
nor U1954 (N_1954,N_1355,N_1040);
or U1955 (N_1955,N_1354,N_1234);
and U1956 (N_1956,N_1001,N_1227);
nor U1957 (N_1957,N_998,N_1207);
xnor U1958 (N_1958,N_1015,N_900);
and U1959 (N_1959,N_1596,N_943);
and U1960 (N_1960,N_1184,N_860);
nor U1961 (N_1961,N_1504,N_1545);
nor U1962 (N_1962,N_884,N_1577);
nand U1963 (N_1963,N_1408,N_825);
nor U1964 (N_1964,N_1494,N_1364);
and U1965 (N_1965,N_841,N_910);
nand U1966 (N_1966,N_851,N_1276);
nand U1967 (N_1967,N_1193,N_1056);
nor U1968 (N_1968,N_1592,N_1173);
and U1969 (N_1969,N_899,N_1531);
nand U1970 (N_1970,N_1467,N_1567);
and U1971 (N_1971,N_1012,N_844);
xor U1972 (N_1972,N_916,N_1532);
or U1973 (N_1973,N_1391,N_936);
or U1974 (N_1974,N_993,N_1275);
or U1975 (N_1975,N_1010,N_1507);
xnor U1976 (N_1976,N_1239,N_1014);
nand U1977 (N_1977,N_837,N_848);
and U1978 (N_1978,N_1164,N_1136);
nand U1979 (N_1979,N_1301,N_964);
nor U1980 (N_1980,N_974,N_961);
xor U1981 (N_1981,N_1556,N_1156);
and U1982 (N_1982,N_1455,N_1305);
nand U1983 (N_1983,N_1573,N_1130);
and U1984 (N_1984,N_1512,N_817);
or U1985 (N_1985,N_952,N_1045);
xor U1986 (N_1986,N_1569,N_1113);
and U1987 (N_1987,N_1067,N_1471);
xnor U1988 (N_1988,N_1557,N_823);
nor U1989 (N_1989,N_1307,N_1465);
and U1990 (N_1990,N_1417,N_1496);
or U1991 (N_1991,N_849,N_1520);
nand U1992 (N_1992,N_904,N_1076);
nor U1993 (N_1993,N_804,N_962);
xor U1994 (N_1994,N_1580,N_1277);
xnor U1995 (N_1995,N_873,N_1549);
nand U1996 (N_1996,N_919,N_1325);
and U1997 (N_1997,N_1103,N_1380);
nand U1998 (N_1998,N_941,N_1114);
or U1999 (N_1999,N_1511,N_1359);
nand U2000 (N_2000,N_1354,N_1072);
and U2001 (N_2001,N_1027,N_1081);
and U2002 (N_2002,N_930,N_1486);
or U2003 (N_2003,N_888,N_1072);
nor U2004 (N_2004,N_1026,N_1528);
or U2005 (N_2005,N_1449,N_1208);
and U2006 (N_2006,N_1184,N_1334);
nor U2007 (N_2007,N_1454,N_1060);
nand U2008 (N_2008,N_1333,N_1095);
nand U2009 (N_2009,N_806,N_946);
or U2010 (N_2010,N_1531,N_1114);
and U2011 (N_2011,N_1051,N_1599);
xnor U2012 (N_2012,N_1393,N_1444);
nor U2013 (N_2013,N_1110,N_1239);
nor U2014 (N_2014,N_846,N_1544);
xor U2015 (N_2015,N_1269,N_922);
xor U2016 (N_2016,N_1562,N_848);
xor U2017 (N_2017,N_1061,N_1562);
or U2018 (N_2018,N_966,N_1555);
xor U2019 (N_2019,N_1557,N_850);
xor U2020 (N_2020,N_1383,N_1559);
nor U2021 (N_2021,N_1395,N_912);
xnor U2022 (N_2022,N_844,N_906);
nor U2023 (N_2023,N_1102,N_1226);
or U2024 (N_2024,N_1124,N_1299);
nand U2025 (N_2025,N_1593,N_1151);
and U2026 (N_2026,N_838,N_1046);
and U2027 (N_2027,N_1380,N_1467);
and U2028 (N_2028,N_1331,N_1388);
and U2029 (N_2029,N_1178,N_1430);
or U2030 (N_2030,N_870,N_1087);
and U2031 (N_2031,N_953,N_1057);
xor U2032 (N_2032,N_1201,N_929);
xnor U2033 (N_2033,N_1200,N_1184);
nand U2034 (N_2034,N_1554,N_865);
or U2035 (N_2035,N_1250,N_1106);
nor U2036 (N_2036,N_1558,N_1319);
xnor U2037 (N_2037,N_1256,N_1159);
or U2038 (N_2038,N_1564,N_1409);
nand U2039 (N_2039,N_1089,N_1265);
or U2040 (N_2040,N_1305,N_1147);
or U2041 (N_2041,N_1155,N_1197);
nor U2042 (N_2042,N_869,N_1028);
xnor U2043 (N_2043,N_1120,N_1172);
nand U2044 (N_2044,N_839,N_1057);
or U2045 (N_2045,N_800,N_1168);
or U2046 (N_2046,N_1135,N_1161);
or U2047 (N_2047,N_1227,N_1437);
nand U2048 (N_2048,N_852,N_922);
nor U2049 (N_2049,N_1381,N_1201);
nand U2050 (N_2050,N_1506,N_1231);
xor U2051 (N_2051,N_898,N_1172);
and U2052 (N_2052,N_1363,N_1088);
nor U2053 (N_2053,N_904,N_1255);
nand U2054 (N_2054,N_958,N_1214);
or U2055 (N_2055,N_1383,N_1235);
or U2056 (N_2056,N_1540,N_1265);
or U2057 (N_2057,N_987,N_1103);
and U2058 (N_2058,N_1074,N_1538);
nor U2059 (N_2059,N_1303,N_1367);
and U2060 (N_2060,N_1424,N_1282);
nand U2061 (N_2061,N_1405,N_1181);
or U2062 (N_2062,N_981,N_1005);
nor U2063 (N_2063,N_977,N_1334);
nor U2064 (N_2064,N_1568,N_1060);
and U2065 (N_2065,N_1417,N_1091);
xnor U2066 (N_2066,N_1439,N_1163);
or U2067 (N_2067,N_1497,N_1358);
xor U2068 (N_2068,N_1149,N_1407);
nor U2069 (N_2069,N_871,N_1283);
nor U2070 (N_2070,N_1547,N_861);
nand U2071 (N_2071,N_1414,N_897);
and U2072 (N_2072,N_1245,N_1307);
xnor U2073 (N_2073,N_1167,N_1289);
and U2074 (N_2074,N_1221,N_878);
xnor U2075 (N_2075,N_1243,N_1333);
nand U2076 (N_2076,N_1137,N_1525);
nor U2077 (N_2077,N_1053,N_1526);
xor U2078 (N_2078,N_1028,N_1471);
or U2079 (N_2079,N_1190,N_1260);
xnor U2080 (N_2080,N_1064,N_835);
nor U2081 (N_2081,N_1599,N_896);
nand U2082 (N_2082,N_1421,N_1353);
nor U2083 (N_2083,N_1199,N_1278);
and U2084 (N_2084,N_1139,N_943);
nor U2085 (N_2085,N_1324,N_826);
or U2086 (N_2086,N_800,N_1364);
nand U2087 (N_2087,N_1107,N_1280);
and U2088 (N_2088,N_1119,N_1309);
and U2089 (N_2089,N_1146,N_1066);
xor U2090 (N_2090,N_1278,N_1237);
and U2091 (N_2091,N_1262,N_837);
and U2092 (N_2092,N_1382,N_1218);
xor U2093 (N_2093,N_1327,N_875);
or U2094 (N_2094,N_1131,N_1568);
and U2095 (N_2095,N_1460,N_1068);
nand U2096 (N_2096,N_1190,N_960);
nand U2097 (N_2097,N_1030,N_1447);
nand U2098 (N_2098,N_949,N_1558);
and U2099 (N_2099,N_1329,N_990);
or U2100 (N_2100,N_1204,N_873);
nand U2101 (N_2101,N_1486,N_1403);
and U2102 (N_2102,N_1346,N_1218);
nand U2103 (N_2103,N_1483,N_1242);
or U2104 (N_2104,N_1133,N_1138);
xnor U2105 (N_2105,N_823,N_887);
xnor U2106 (N_2106,N_1490,N_1046);
nor U2107 (N_2107,N_860,N_1230);
nand U2108 (N_2108,N_1498,N_1558);
or U2109 (N_2109,N_939,N_1348);
and U2110 (N_2110,N_1069,N_904);
or U2111 (N_2111,N_884,N_828);
and U2112 (N_2112,N_1146,N_869);
or U2113 (N_2113,N_802,N_984);
nand U2114 (N_2114,N_1247,N_950);
nand U2115 (N_2115,N_850,N_1136);
nand U2116 (N_2116,N_1171,N_1320);
nand U2117 (N_2117,N_1239,N_1418);
or U2118 (N_2118,N_1089,N_1019);
nor U2119 (N_2119,N_818,N_1246);
or U2120 (N_2120,N_1018,N_1236);
nor U2121 (N_2121,N_1351,N_852);
xor U2122 (N_2122,N_1425,N_1056);
or U2123 (N_2123,N_1356,N_1507);
or U2124 (N_2124,N_938,N_1565);
or U2125 (N_2125,N_1257,N_1224);
nor U2126 (N_2126,N_1147,N_1531);
or U2127 (N_2127,N_1385,N_1582);
and U2128 (N_2128,N_1121,N_1162);
nand U2129 (N_2129,N_1324,N_1516);
xnor U2130 (N_2130,N_830,N_1414);
or U2131 (N_2131,N_1304,N_1401);
nor U2132 (N_2132,N_869,N_878);
and U2133 (N_2133,N_1255,N_1132);
nor U2134 (N_2134,N_811,N_1383);
or U2135 (N_2135,N_1016,N_1544);
and U2136 (N_2136,N_1089,N_1544);
xor U2137 (N_2137,N_1255,N_1599);
xnor U2138 (N_2138,N_1447,N_1427);
xnor U2139 (N_2139,N_1537,N_1319);
nand U2140 (N_2140,N_1146,N_1407);
nor U2141 (N_2141,N_1342,N_904);
xnor U2142 (N_2142,N_1326,N_1103);
xor U2143 (N_2143,N_1137,N_1514);
and U2144 (N_2144,N_989,N_1275);
and U2145 (N_2145,N_1596,N_1313);
or U2146 (N_2146,N_1048,N_1413);
and U2147 (N_2147,N_846,N_910);
xnor U2148 (N_2148,N_1538,N_1494);
xnor U2149 (N_2149,N_1208,N_1375);
or U2150 (N_2150,N_1170,N_1339);
xnor U2151 (N_2151,N_1124,N_1332);
or U2152 (N_2152,N_905,N_1077);
nor U2153 (N_2153,N_1531,N_1591);
nand U2154 (N_2154,N_1369,N_1297);
xnor U2155 (N_2155,N_1030,N_1169);
xor U2156 (N_2156,N_1311,N_943);
nor U2157 (N_2157,N_1087,N_1059);
and U2158 (N_2158,N_1023,N_1544);
xor U2159 (N_2159,N_1246,N_1069);
and U2160 (N_2160,N_1413,N_1557);
and U2161 (N_2161,N_1574,N_1186);
and U2162 (N_2162,N_849,N_1080);
xnor U2163 (N_2163,N_1301,N_1024);
xnor U2164 (N_2164,N_910,N_838);
xnor U2165 (N_2165,N_853,N_1262);
xor U2166 (N_2166,N_1536,N_1365);
nand U2167 (N_2167,N_1088,N_1238);
xnor U2168 (N_2168,N_1531,N_1117);
xnor U2169 (N_2169,N_1128,N_1041);
nand U2170 (N_2170,N_1021,N_1172);
nor U2171 (N_2171,N_1350,N_1240);
nand U2172 (N_2172,N_926,N_1580);
nand U2173 (N_2173,N_823,N_952);
nor U2174 (N_2174,N_899,N_1561);
nor U2175 (N_2175,N_1168,N_1048);
nand U2176 (N_2176,N_1073,N_1334);
and U2177 (N_2177,N_959,N_1012);
nor U2178 (N_2178,N_1511,N_978);
xnor U2179 (N_2179,N_809,N_816);
and U2180 (N_2180,N_1500,N_1370);
xor U2181 (N_2181,N_1138,N_1112);
nand U2182 (N_2182,N_1055,N_1297);
or U2183 (N_2183,N_870,N_1042);
nor U2184 (N_2184,N_1558,N_1006);
nand U2185 (N_2185,N_1330,N_1126);
xor U2186 (N_2186,N_1042,N_1034);
nand U2187 (N_2187,N_1058,N_1270);
nor U2188 (N_2188,N_1347,N_1582);
nand U2189 (N_2189,N_911,N_1014);
nand U2190 (N_2190,N_1589,N_1299);
nand U2191 (N_2191,N_1361,N_1272);
and U2192 (N_2192,N_907,N_1414);
and U2193 (N_2193,N_1194,N_1524);
nor U2194 (N_2194,N_890,N_863);
xor U2195 (N_2195,N_1438,N_1009);
nand U2196 (N_2196,N_1181,N_954);
or U2197 (N_2197,N_1036,N_1207);
xnor U2198 (N_2198,N_1362,N_1234);
nand U2199 (N_2199,N_888,N_1169);
or U2200 (N_2200,N_1119,N_824);
nand U2201 (N_2201,N_1009,N_1211);
nor U2202 (N_2202,N_1499,N_1297);
nor U2203 (N_2203,N_1515,N_1021);
and U2204 (N_2204,N_1341,N_1488);
or U2205 (N_2205,N_1254,N_813);
and U2206 (N_2206,N_932,N_1083);
nand U2207 (N_2207,N_1468,N_843);
and U2208 (N_2208,N_971,N_964);
or U2209 (N_2209,N_1193,N_1130);
and U2210 (N_2210,N_896,N_1525);
xnor U2211 (N_2211,N_1189,N_854);
nand U2212 (N_2212,N_1193,N_1302);
and U2213 (N_2213,N_874,N_1546);
nor U2214 (N_2214,N_1130,N_980);
or U2215 (N_2215,N_972,N_829);
nor U2216 (N_2216,N_1558,N_1399);
or U2217 (N_2217,N_907,N_1362);
and U2218 (N_2218,N_1009,N_1566);
nor U2219 (N_2219,N_1004,N_1504);
nand U2220 (N_2220,N_1353,N_1199);
and U2221 (N_2221,N_847,N_1290);
nand U2222 (N_2222,N_1534,N_1544);
and U2223 (N_2223,N_1384,N_1216);
nand U2224 (N_2224,N_1055,N_1520);
nor U2225 (N_2225,N_1225,N_1412);
or U2226 (N_2226,N_1372,N_1105);
and U2227 (N_2227,N_1146,N_822);
nand U2228 (N_2228,N_1389,N_951);
or U2229 (N_2229,N_1268,N_991);
xnor U2230 (N_2230,N_896,N_838);
nand U2231 (N_2231,N_1033,N_1552);
nor U2232 (N_2232,N_1097,N_1104);
or U2233 (N_2233,N_1492,N_1444);
nand U2234 (N_2234,N_947,N_1367);
and U2235 (N_2235,N_1230,N_809);
nor U2236 (N_2236,N_1530,N_1484);
or U2237 (N_2237,N_1496,N_1015);
or U2238 (N_2238,N_945,N_1437);
nand U2239 (N_2239,N_809,N_1365);
or U2240 (N_2240,N_1350,N_1134);
nand U2241 (N_2241,N_1176,N_854);
or U2242 (N_2242,N_1072,N_1102);
xor U2243 (N_2243,N_812,N_821);
or U2244 (N_2244,N_1159,N_1285);
nand U2245 (N_2245,N_980,N_1553);
nor U2246 (N_2246,N_1305,N_812);
nor U2247 (N_2247,N_1592,N_939);
nand U2248 (N_2248,N_868,N_1404);
or U2249 (N_2249,N_1034,N_1312);
xnor U2250 (N_2250,N_980,N_1264);
or U2251 (N_2251,N_1599,N_1458);
xnor U2252 (N_2252,N_1582,N_1545);
or U2253 (N_2253,N_1462,N_1093);
or U2254 (N_2254,N_949,N_1547);
nor U2255 (N_2255,N_990,N_1456);
xnor U2256 (N_2256,N_1393,N_1029);
xnor U2257 (N_2257,N_1530,N_1251);
xor U2258 (N_2258,N_889,N_926);
xor U2259 (N_2259,N_860,N_1267);
nor U2260 (N_2260,N_1441,N_951);
or U2261 (N_2261,N_800,N_1196);
nor U2262 (N_2262,N_888,N_801);
xnor U2263 (N_2263,N_1366,N_1490);
or U2264 (N_2264,N_1002,N_826);
or U2265 (N_2265,N_1160,N_1549);
nor U2266 (N_2266,N_1058,N_971);
xor U2267 (N_2267,N_837,N_1205);
and U2268 (N_2268,N_1297,N_1166);
and U2269 (N_2269,N_1426,N_931);
and U2270 (N_2270,N_1384,N_1549);
nand U2271 (N_2271,N_1308,N_1591);
nor U2272 (N_2272,N_1180,N_1592);
or U2273 (N_2273,N_1148,N_867);
and U2274 (N_2274,N_1322,N_950);
or U2275 (N_2275,N_1405,N_1424);
xor U2276 (N_2276,N_1200,N_1018);
and U2277 (N_2277,N_953,N_1567);
nand U2278 (N_2278,N_814,N_1226);
xnor U2279 (N_2279,N_1080,N_1372);
nor U2280 (N_2280,N_903,N_930);
xnor U2281 (N_2281,N_1405,N_1275);
nand U2282 (N_2282,N_891,N_1209);
and U2283 (N_2283,N_953,N_1232);
nor U2284 (N_2284,N_1157,N_1435);
or U2285 (N_2285,N_1593,N_1590);
xor U2286 (N_2286,N_1117,N_1121);
and U2287 (N_2287,N_1074,N_1263);
nand U2288 (N_2288,N_1181,N_1029);
nor U2289 (N_2289,N_1487,N_910);
and U2290 (N_2290,N_1080,N_1358);
and U2291 (N_2291,N_939,N_1138);
nand U2292 (N_2292,N_1407,N_1127);
xnor U2293 (N_2293,N_1217,N_965);
nor U2294 (N_2294,N_882,N_1233);
xnor U2295 (N_2295,N_1378,N_1472);
xnor U2296 (N_2296,N_831,N_1525);
nor U2297 (N_2297,N_1072,N_1099);
nand U2298 (N_2298,N_1408,N_1565);
or U2299 (N_2299,N_961,N_1241);
and U2300 (N_2300,N_974,N_827);
nand U2301 (N_2301,N_1207,N_867);
and U2302 (N_2302,N_1049,N_1292);
nand U2303 (N_2303,N_946,N_801);
nor U2304 (N_2304,N_1444,N_1323);
and U2305 (N_2305,N_1092,N_1545);
nand U2306 (N_2306,N_958,N_1445);
nor U2307 (N_2307,N_1431,N_1117);
nor U2308 (N_2308,N_1321,N_1463);
nor U2309 (N_2309,N_1024,N_820);
nand U2310 (N_2310,N_1187,N_911);
nand U2311 (N_2311,N_868,N_911);
xnor U2312 (N_2312,N_1111,N_1470);
xor U2313 (N_2313,N_981,N_1299);
and U2314 (N_2314,N_1331,N_1290);
nand U2315 (N_2315,N_1127,N_958);
nand U2316 (N_2316,N_1323,N_1372);
and U2317 (N_2317,N_1238,N_882);
or U2318 (N_2318,N_1165,N_814);
nor U2319 (N_2319,N_1371,N_1098);
and U2320 (N_2320,N_1228,N_1267);
and U2321 (N_2321,N_1235,N_1286);
or U2322 (N_2322,N_819,N_1349);
or U2323 (N_2323,N_1178,N_1132);
nand U2324 (N_2324,N_1422,N_852);
nand U2325 (N_2325,N_1203,N_988);
xnor U2326 (N_2326,N_1529,N_1006);
and U2327 (N_2327,N_1046,N_1528);
nor U2328 (N_2328,N_1234,N_1439);
or U2329 (N_2329,N_838,N_1006);
or U2330 (N_2330,N_1322,N_1268);
xor U2331 (N_2331,N_888,N_1343);
and U2332 (N_2332,N_1455,N_1416);
and U2333 (N_2333,N_1110,N_1467);
nor U2334 (N_2334,N_1247,N_935);
and U2335 (N_2335,N_996,N_816);
or U2336 (N_2336,N_1392,N_1263);
or U2337 (N_2337,N_1406,N_1090);
or U2338 (N_2338,N_1372,N_1368);
or U2339 (N_2339,N_1308,N_1186);
xnor U2340 (N_2340,N_918,N_1537);
or U2341 (N_2341,N_1079,N_1407);
nor U2342 (N_2342,N_871,N_1382);
or U2343 (N_2343,N_1115,N_1562);
or U2344 (N_2344,N_1354,N_1012);
nand U2345 (N_2345,N_971,N_914);
nor U2346 (N_2346,N_1546,N_1152);
nand U2347 (N_2347,N_1315,N_923);
and U2348 (N_2348,N_1297,N_1505);
or U2349 (N_2349,N_1143,N_1101);
nor U2350 (N_2350,N_1032,N_1263);
xor U2351 (N_2351,N_961,N_898);
nand U2352 (N_2352,N_826,N_1147);
nor U2353 (N_2353,N_1467,N_1051);
xor U2354 (N_2354,N_1374,N_1406);
nand U2355 (N_2355,N_1444,N_1130);
xnor U2356 (N_2356,N_888,N_853);
nand U2357 (N_2357,N_1431,N_1335);
and U2358 (N_2358,N_986,N_977);
and U2359 (N_2359,N_1454,N_1111);
or U2360 (N_2360,N_1243,N_1586);
or U2361 (N_2361,N_1085,N_1265);
and U2362 (N_2362,N_1437,N_1057);
xor U2363 (N_2363,N_1005,N_974);
and U2364 (N_2364,N_1049,N_1564);
or U2365 (N_2365,N_1574,N_1047);
and U2366 (N_2366,N_975,N_1278);
xnor U2367 (N_2367,N_979,N_867);
nor U2368 (N_2368,N_1420,N_1213);
or U2369 (N_2369,N_1202,N_1340);
nand U2370 (N_2370,N_1128,N_1030);
and U2371 (N_2371,N_1218,N_1329);
and U2372 (N_2372,N_1478,N_998);
xnor U2373 (N_2373,N_1559,N_1307);
xnor U2374 (N_2374,N_1128,N_1519);
xor U2375 (N_2375,N_853,N_1177);
nand U2376 (N_2376,N_1422,N_1598);
and U2377 (N_2377,N_810,N_1262);
or U2378 (N_2378,N_1253,N_1458);
xor U2379 (N_2379,N_1551,N_1070);
or U2380 (N_2380,N_1040,N_837);
xor U2381 (N_2381,N_985,N_888);
nand U2382 (N_2382,N_1163,N_1482);
nor U2383 (N_2383,N_920,N_1256);
or U2384 (N_2384,N_1487,N_1343);
or U2385 (N_2385,N_1553,N_1178);
nor U2386 (N_2386,N_1354,N_1342);
and U2387 (N_2387,N_970,N_1426);
and U2388 (N_2388,N_1449,N_1429);
nor U2389 (N_2389,N_1239,N_1248);
nor U2390 (N_2390,N_1460,N_1583);
nor U2391 (N_2391,N_1416,N_1548);
or U2392 (N_2392,N_1543,N_1557);
nand U2393 (N_2393,N_1221,N_1244);
xnor U2394 (N_2394,N_1248,N_1595);
nand U2395 (N_2395,N_1043,N_936);
nand U2396 (N_2396,N_1388,N_1546);
or U2397 (N_2397,N_969,N_1586);
and U2398 (N_2398,N_900,N_1585);
or U2399 (N_2399,N_1016,N_1429);
and U2400 (N_2400,N_2242,N_2295);
nor U2401 (N_2401,N_1937,N_1951);
xor U2402 (N_2402,N_2397,N_1991);
nand U2403 (N_2403,N_1875,N_2247);
nand U2404 (N_2404,N_1810,N_2148);
nand U2405 (N_2405,N_2332,N_2105);
nand U2406 (N_2406,N_1739,N_2134);
and U2407 (N_2407,N_2157,N_1908);
and U2408 (N_2408,N_1858,N_2354);
or U2409 (N_2409,N_1837,N_2051);
nand U2410 (N_2410,N_2233,N_1771);
xor U2411 (N_2411,N_2282,N_2097);
nor U2412 (N_2412,N_1987,N_1948);
nor U2413 (N_2413,N_1836,N_2151);
nand U2414 (N_2414,N_2228,N_2240);
or U2415 (N_2415,N_1890,N_1746);
nand U2416 (N_2416,N_1902,N_2376);
and U2417 (N_2417,N_1792,N_1927);
nand U2418 (N_2418,N_2081,N_2175);
xor U2419 (N_2419,N_2079,N_1730);
nand U2420 (N_2420,N_2275,N_1964);
nor U2421 (N_2421,N_2193,N_1852);
xor U2422 (N_2422,N_2230,N_2319);
or U2423 (N_2423,N_1826,N_1667);
or U2424 (N_2424,N_1957,N_1777);
and U2425 (N_2425,N_2351,N_1726);
or U2426 (N_2426,N_1863,N_1648);
nand U2427 (N_2427,N_2125,N_2205);
nand U2428 (N_2428,N_1738,N_2025);
and U2429 (N_2429,N_2234,N_2321);
nor U2430 (N_2430,N_2024,N_1926);
and U2431 (N_2431,N_2216,N_1924);
nand U2432 (N_2432,N_2209,N_2269);
nand U2433 (N_2433,N_2019,N_1815);
xor U2434 (N_2434,N_2217,N_2342);
nor U2435 (N_2435,N_1664,N_2244);
and U2436 (N_2436,N_1958,N_2361);
nand U2437 (N_2437,N_1993,N_1687);
nor U2438 (N_2438,N_1805,N_1950);
nand U2439 (N_2439,N_1692,N_2178);
or U2440 (N_2440,N_2281,N_1772);
xor U2441 (N_2441,N_2182,N_2374);
xnor U2442 (N_2442,N_1980,N_1702);
or U2443 (N_2443,N_2325,N_1780);
or U2444 (N_2444,N_1804,N_2044);
nand U2445 (N_2445,N_2150,N_2066);
or U2446 (N_2446,N_2312,N_2252);
nor U2447 (N_2447,N_2398,N_1939);
and U2448 (N_2448,N_1838,N_1713);
xor U2449 (N_2449,N_2337,N_1676);
xnor U2450 (N_2450,N_2388,N_1659);
and U2451 (N_2451,N_2339,N_1775);
or U2452 (N_2452,N_2259,N_2028);
xor U2453 (N_2453,N_2063,N_2095);
and U2454 (N_2454,N_1982,N_2224);
nand U2455 (N_2455,N_2147,N_2001);
xnor U2456 (N_2456,N_1936,N_1685);
or U2457 (N_2457,N_1720,N_1967);
or U2458 (N_2458,N_2219,N_2049);
nand U2459 (N_2459,N_1707,N_1921);
nand U2460 (N_2460,N_2386,N_1671);
nand U2461 (N_2461,N_2077,N_2393);
nor U2462 (N_2462,N_2304,N_1626);
nand U2463 (N_2463,N_1873,N_1829);
and U2464 (N_2464,N_2368,N_2174);
or U2465 (N_2465,N_2061,N_2099);
xor U2466 (N_2466,N_1725,N_1963);
nor U2467 (N_2467,N_1846,N_2006);
xnor U2468 (N_2468,N_1680,N_1642);
nor U2469 (N_2469,N_2267,N_2322);
or U2470 (N_2470,N_2221,N_2232);
or U2471 (N_2471,N_2262,N_2017);
and U2472 (N_2472,N_1818,N_2199);
xnor U2473 (N_2473,N_1768,N_2004);
and U2474 (N_2474,N_1920,N_2293);
and U2475 (N_2475,N_1828,N_2067);
xor U2476 (N_2476,N_2359,N_2333);
xor U2477 (N_2477,N_1946,N_2071);
nor U2478 (N_2478,N_2083,N_2016);
nor U2479 (N_2479,N_1744,N_1691);
xor U2480 (N_2480,N_1990,N_1756);
xnor U2481 (N_2481,N_1679,N_1786);
and U2482 (N_2482,N_1952,N_2029);
and U2483 (N_2483,N_2085,N_1623);
and U2484 (N_2484,N_1645,N_1953);
and U2485 (N_2485,N_2270,N_2145);
xor U2486 (N_2486,N_1827,N_1715);
nand U2487 (N_2487,N_1968,N_1822);
and U2488 (N_2488,N_2377,N_1718);
nand U2489 (N_2489,N_1974,N_2180);
nand U2490 (N_2490,N_2363,N_1997);
or U2491 (N_2491,N_1811,N_1901);
nor U2492 (N_2492,N_2346,N_2208);
xnor U2493 (N_2493,N_1868,N_2265);
nand U2494 (N_2494,N_1847,N_2106);
nand U2495 (N_2495,N_2204,N_2033);
nand U2496 (N_2496,N_1985,N_1918);
nand U2497 (N_2497,N_1959,N_2306);
xor U2498 (N_2498,N_2311,N_1857);
or U2499 (N_2499,N_2328,N_2168);
nor U2500 (N_2500,N_1923,N_1840);
nand U2501 (N_2501,N_2301,N_2197);
and U2502 (N_2502,N_1612,N_2039);
nand U2503 (N_2503,N_2349,N_2202);
nor U2504 (N_2504,N_2384,N_2036);
xnor U2505 (N_2505,N_2280,N_2268);
nand U2506 (N_2506,N_1709,N_1930);
nand U2507 (N_2507,N_1661,N_1844);
nor U2508 (N_2508,N_2241,N_2166);
or U2509 (N_2509,N_2188,N_1616);
or U2510 (N_2510,N_2082,N_1611);
xor U2511 (N_2511,N_2052,N_1878);
nor U2512 (N_2512,N_1871,N_2013);
and U2513 (N_2513,N_2096,N_1719);
nor U2514 (N_2514,N_2191,N_1755);
and U2515 (N_2515,N_2394,N_2130);
xnor U2516 (N_2516,N_2399,N_2264);
xor U2517 (N_2517,N_2245,N_2355);
xor U2518 (N_2518,N_2032,N_2250);
or U2519 (N_2519,N_2173,N_1798);
and U2520 (N_2520,N_2059,N_1977);
nor U2521 (N_2521,N_2334,N_2313);
or U2522 (N_2522,N_1649,N_2222);
xnor U2523 (N_2523,N_1657,N_2225);
nor U2524 (N_2524,N_1619,N_1861);
nand U2525 (N_2525,N_2088,N_1915);
xor U2526 (N_2526,N_2366,N_1632);
xor U2527 (N_2527,N_2251,N_1885);
nor U2528 (N_2528,N_1891,N_1678);
or U2529 (N_2529,N_2046,N_1637);
or U2530 (N_2530,N_2102,N_2153);
nor U2531 (N_2531,N_2220,N_2119);
and U2532 (N_2532,N_2315,N_1866);
xnor U2533 (N_2533,N_1631,N_1943);
nand U2534 (N_2534,N_1621,N_1851);
nor U2535 (N_2535,N_1893,N_2190);
nor U2536 (N_2536,N_1620,N_2296);
xnor U2537 (N_2537,N_2141,N_2135);
and U2538 (N_2538,N_1938,N_1874);
and U2539 (N_2539,N_2164,N_1971);
xor U2540 (N_2540,N_2327,N_2292);
nor U2541 (N_2541,N_1770,N_1865);
or U2542 (N_2542,N_1710,N_1842);
nor U2543 (N_2543,N_2114,N_2323);
nor U2544 (N_2544,N_2158,N_1763);
or U2545 (N_2545,N_1869,N_1684);
nor U2546 (N_2546,N_1793,N_1655);
nor U2547 (N_2547,N_2189,N_2035);
and U2548 (N_2548,N_1894,N_2116);
xor U2549 (N_2549,N_2131,N_2239);
nor U2550 (N_2550,N_1622,N_2162);
and U2551 (N_2551,N_1727,N_1643);
or U2552 (N_2552,N_1724,N_1774);
nor U2553 (N_2553,N_2179,N_1779);
or U2554 (N_2554,N_1813,N_2196);
nor U2555 (N_2555,N_1625,N_1834);
nor U2556 (N_2556,N_2139,N_2258);
or U2557 (N_2557,N_1624,N_1797);
nor U2558 (N_2558,N_1633,N_1759);
xor U2559 (N_2559,N_1748,N_2290);
and U2560 (N_2560,N_1884,N_1652);
and U2561 (N_2561,N_1758,N_1882);
nand U2562 (N_2562,N_1799,N_2299);
and U2563 (N_2563,N_1636,N_2211);
nor U2564 (N_2564,N_2177,N_2243);
nand U2565 (N_2565,N_1752,N_2195);
nor U2566 (N_2566,N_2170,N_1658);
or U2567 (N_2567,N_1925,N_1881);
or U2568 (N_2568,N_1654,N_2201);
and U2569 (N_2569,N_1911,N_2038);
or U2570 (N_2570,N_2065,N_2331);
nand U2571 (N_2571,N_1895,N_2068);
and U2572 (N_2572,N_2031,N_1954);
nand U2573 (N_2573,N_1751,N_1864);
nand U2574 (N_2574,N_2317,N_1618);
and U2575 (N_2575,N_1870,N_2336);
and U2576 (N_2576,N_2003,N_2060);
nand U2577 (N_2577,N_2020,N_2372);
nor U2578 (N_2578,N_1802,N_2272);
xnor U2579 (N_2579,N_1635,N_2340);
nand U2580 (N_2580,N_1975,N_2070);
and U2581 (N_2581,N_1883,N_1704);
and U2582 (N_2582,N_2030,N_1711);
nand U2583 (N_2583,N_2045,N_1675);
and U2584 (N_2584,N_1877,N_2360);
nand U2585 (N_2585,N_2223,N_2380);
nor U2586 (N_2586,N_1969,N_2379);
nor U2587 (N_2587,N_2218,N_1889);
or U2588 (N_2588,N_1809,N_2192);
xnor U2589 (N_2589,N_2200,N_1742);
and U2590 (N_2590,N_1766,N_2140);
nor U2591 (N_2591,N_1694,N_2289);
nor U2592 (N_2592,N_1686,N_2369);
nor U2593 (N_2593,N_2255,N_2329);
xor U2594 (N_2594,N_1830,N_1919);
or U2595 (N_2595,N_2002,N_1849);
xnor U2596 (N_2596,N_1788,N_2365);
and U2597 (N_2597,N_2261,N_1860);
nor U2598 (N_2598,N_2136,N_1929);
nor U2599 (N_2599,N_1723,N_1613);
nand U2600 (N_2600,N_1634,N_2187);
nor U2601 (N_2601,N_2287,N_2142);
xnor U2602 (N_2602,N_2027,N_1972);
nor U2603 (N_2603,N_1647,N_1761);
nor U2604 (N_2604,N_2344,N_1888);
and U2605 (N_2605,N_1955,N_2310);
and U2606 (N_2606,N_1904,N_2056);
nand U2607 (N_2607,N_2010,N_1845);
or U2608 (N_2608,N_2260,N_1690);
nand U2609 (N_2609,N_2214,N_2037);
or U2610 (N_2610,N_1970,N_1716);
or U2611 (N_2611,N_2152,N_1862);
nor U2612 (N_2612,N_2090,N_2364);
nand U2613 (N_2613,N_1749,N_1731);
nor U2614 (N_2614,N_2098,N_1941);
nor U2615 (N_2615,N_2091,N_2387);
and U2616 (N_2616,N_1767,N_1602);
nand U2617 (N_2617,N_1850,N_2254);
or U2618 (N_2618,N_2129,N_2236);
nand U2619 (N_2619,N_1764,N_1745);
xor U2620 (N_2620,N_1714,N_2383);
nand U2621 (N_2621,N_1614,N_1601);
xnor U2622 (N_2622,N_2127,N_2103);
or U2623 (N_2623,N_1996,N_2078);
and U2624 (N_2624,N_1898,N_1892);
and U2625 (N_2625,N_1922,N_1728);
nor U2626 (N_2626,N_2367,N_2335);
and U2627 (N_2627,N_1722,N_1703);
or U2628 (N_2628,N_2318,N_1905);
nand U2629 (N_2629,N_1769,N_2207);
nand U2630 (N_2630,N_2014,N_2326);
xor U2631 (N_2631,N_2283,N_1670);
nand U2632 (N_2632,N_1747,N_2146);
nand U2633 (N_2633,N_2396,N_1897);
xor U2634 (N_2634,N_1833,N_2277);
xnor U2635 (N_2635,N_1785,N_2171);
nand U2636 (N_2636,N_2133,N_1832);
or U2637 (N_2637,N_1914,N_1665);
nor U2638 (N_2638,N_2165,N_2298);
nor U2639 (N_2639,N_2348,N_2279);
nand U2640 (N_2640,N_1879,N_2297);
nand U2641 (N_2641,N_1773,N_1700);
or U2642 (N_2642,N_1663,N_1682);
nand U2643 (N_2643,N_2112,N_2084);
xnor U2644 (N_2644,N_1956,N_2314);
xnor U2645 (N_2645,N_1672,N_2062);
or U2646 (N_2646,N_2212,N_2373);
or U2647 (N_2647,N_1896,N_1988);
nor U2648 (N_2648,N_2235,N_2138);
and U2649 (N_2649,N_2213,N_2149);
and U2650 (N_2650,N_2385,N_1949);
nor U2651 (N_2651,N_2113,N_1812);
xor U2652 (N_2652,N_2126,N_2155);
xor U2653 (N_2653,N_2302,N_2352);
nand U2654 (N_2654,N_1853,N_2276);
nand U2655 (N_2655,N_2163,N_2054);
or U2656 (N_2656,N_2042,N_2238);
nor U2657 (N_2657,N_2274,N_2072);
xor U2658 (N_2658,N_1604,N_2172);
nor U2659 (N_2659,N_2012,N_1708);
or U2660 (N_2660,N_2023,N_1706);
or U2661 (N_2661,N_2058,N_1617);
nor U2662 (N_2662,N_2169,N_2167);
or U2663 (N_2663,N_2215,N_1754);
nand U2664 (N_2664,N_2055,N_1784);
and U2665 (N_2665,N_2249,N_2370);
and U2666 (N_2666,N_2076,N_1629);
xnor U2667 (N_2667,N_2294,N_2330);
nor U2668 (N_2668,N_2176,N_2338);
xnor U2669 (N_2669,N_1807,N_1666);
xor U2670 (N_2670,N_1765,N_2007);
or U2671 (N_2671,N_1732,N_2288);
xor U2672 (N_2672,N_1683,N_2390);
nand U2673 (N_2673,N_1992,N_1856);
nor U2674 (N_2674,N_2362,N_1935);
xnor U2675 (N_2675,N_1729,N_1867);
and U2676 (N_2676,N_2256,N_2389);
and U2677 (N_2677,N_2104,N_1907);
xnor U2678 (N_2678,N_1932,N_1933);
or U2679 (N_2679,N_2011,N_1942);
nor U2680 (N_2680,N_1825,N_2266);
or U2681 (N_2681,N_1790,N_2120);
and U2682 (N_2682,N_2381,N_2021);
nand U2683 (N_2683,N_2307,N_1615);
or U2684 (N_2684,N_2047,N_1880);
or U2685 (N_2685,N_1931,N_2137);
and U2686 (N_2686,N_2350,N_1848);
nor U2687 (N_2687,N_1795,N_1721);
nand U2688 (N_2688,N_2353,N_1843);
nor U2689 (N_2689,N_1839,N_2206);
nand U2690 (N_2690,N_2073,N_1787);
or U2691 (N_2691,N_2356,N_2237);
and U2692 (N_2692,N_1859,N_1876);
and U2693 (N_2693,N_1688,N_2053);
nand U2694 (N_2694,N_1960,N_1803);
nor U2695 (N_2695,N_1651,N_1757);
nor U2696 (N_2696,N_2111,N_1824);
xor U2697 (N_2697,N_2101,N_1650);
nand U2698 (N_2698,N_2375,N_1947);
nor U2699 (N_2699,N_2253,N_1607);
and U2700 (N_2700,N_1854,N_2194);
nand U2701 (N_2701,N_2122,N_1609);
or U2702 (N_2702,N_1979,N_1981);
or U2703 (N_2703,N_2286,N_1821);
or U2704 (N_2704,N_2395,N_2022);
nand U2705 (N_2705,N_2303,N_2278);
xor U2706 (N_2706,N_1741,N_2285);
or U2707 (N_2707,N_1961,N_1791);
or U2708 (N_2708,N_1762,N_2005);
or U2709 (N_2709,N_1989,N_2392);
nor U2710 (N_2710,N_1886,N_1872);
or U2711 (N_2711,N_1934,N_2305);
nor U2712 (N_2712,N_2093,N_1819);
nand U2713 (N_2713,N_2057,N_2124);
nand U2714 (N_2714,N_2118,N_1630);
and U2715 (N_2715,N_2161,N_1794);
nor U2716 (N_2716,N_1734,N_2257);
or U2717 (N_2717,N_1928,N_1668);
or U2718 (N_2718,N_1945,N_1962);
and U2719 (N_2719,N_1900,N_2358);
xnor U2720 (N_2720,N_1778,N_1660);
xor U2721 (N_2721,N_2271,N_1673);
and U2722 (N_2722,N_1628,N_2080);
xnor U2723 (N_2723,N_1760,N_1603);
and U2724 (N_2724,N_1646,N_1699);
nand U2725 (N_2725,N_2391,N_1677);
nor U2726 (N_2726,N_1823,N_2086);
and U2727 (N_2727,N_1750,N_2229);
and U2728 (N_2728,N_2026,N_1717);
nor U2729 (N_2729,N_1627,N_1712);
and U2730 (N_2730,N_2343,N_2040);
xor U2731 (N_2731,N_2308,N_1965);
xor U2732 (N_2732,N_1817,N_1831);
or U2733 (N_2733,N_2227,N_1806);
nor U2734 (N_2734,N_2341,N_2345);
nor U2735 (N_2735,N_2092,N_1662);
or U2736 (N_2736,N_1693,N_2089);
xor U2737 (N_2737,N_1973,N_1743);
xnor U2738 (N_2738,N_1841,N_2132);
nor U2739 (N_2739,N_2121,N_1610);
nor U2740 (N_2740,N_2094,N_2231);
nand U2741 (N_2741,N_2009,N_2316);
or U2742 (N_2742,N_1800,N_2123);
nand U2743 (N_2743,N_2246,N_2110);
and U2744 (N_2744,N_2357,N_1966);
or U2745 (N_2745,N_2226,N_1753);
nand U2746 (N_2746,N_2160,N_2186);
xnor U2747 (N_2747,N_2382,N_1909);
xnor U2748 (N_2748,N_2185,N_1600);
nor U2749 (N_2749,N_1940,N_1814);
and U2750 (N_2750,N_2371,N_2156);
and U2751 (N_2751,N_1776,N_2159);
nor U2752 (N_2752,N_1994,N_1820);
nand U2753 (N_2753,N_1608,N_1783);
nand U2754 (N_2754,N_1782,N_2074);
nand U2755 (N_2755,N_1835,N_2210);
or U2756 (N_2756,N_1735,N_1605);
nor U2757 (N_2757,N_1789,N_2043);
or U2758 (N_2758,N_1669,N_2109);
nand U2759 (N_2759,N_2181,N_1917);
or U2760 (N_2760,N_2075,N_2263);
and U2761 (N_2761,N_1695,N_1903);
nor U2762 (N_2762,N_2184,N_1698);
nand U2763 (N_2763,N_2018,N_2107);
or U2764 (N_2764,N_2273,N_1640);
nor U2765 (N_2765,N_1606,N_2320);
nor U2766 (N_2766,N_1740,N_1906);
and U2767 (N_2767,N_1705,N_2034);
and U2768 (N_2768,N_1781,N_2008);
nand U2769 (N_2769,N_2284,N_2108);
nor U2770 (N_2770,N_1639,N_2378);
or U2771 (N_2771,N_1816,N_2015);
nand U2772 (N_2772,N_2154,N_1701);
nand U2773 (N_2773,N_1656,N_1983);
nand U2774 (N_2774,N_2198,N_1986);
xnor U2775 (N_2775,N_2100,N_2291);
nand U2776 (N_2776,N_1737,N_2143);
xnor U2777 (N_2777,N_2128,N_1855);
or U2778 (N_2778,N_1995,N_2050);
nor U2779 (N_2779,N_1733,N_1913);
and U2780 (N_2780,N_1978,N_1674);
nand U2781 (N_2781,N_1689,N_2144);
or U2782 (N_2782,N_1999,N_1808);
nor U2783 (N_2783,N_2309,N_2183);
nor U2784 (N_2784,N_2064,N_1887);
and U2785 (N_2785,N_2000,N_2117);
xnor U2786 (N_2786,N_1998,N_2300);
and U2787 (N_2787,N_1916,N_2041);
nor U2788 (N_2788,N_1976,N_1912);
or U2789 (N_2789,N_1736,N_1910);
or U2790 (N_2790,N_1796,N_2115);
or U2791 (N_2791,N_1644,N_1641);
or U2792 (N_2792,N_2087,N_1944);
nand U2793 (N_2793,N_1697,N_1638);
or U2794 (N_2794,N_1696,N_2203);
xnor U2795 (N_2795,N_1801,N_2248);
or U2796 (N_2796,N_2347,N_1681);
or U2797 (N_2797,N_2324,N_1653);
and U2798 (N_2798,N_2069,N_1899);
or U2799 (N_2799,N_1984,N_2048);
or U2800 (N_2800,N_2090,N_2180);
and U2801 (N_2801,N_2341,N_1890);
nand U2802 (N_2802,N_2041,N_2390);
and U2803 (N_2803,N_2184,N_2129);
or U2804 (N_2804,N_2336,N_1855);
xnor U2805 (N_2805,N_1781,N_1810);
and U2806 (N_2806,N_1848,N_2201);
xnor U2807 (N_2807,N_1718,N_1678);
nand U2808 (N_2808,N_2223,N_1602);
nand U2809 (N_2809,N_2212,N_1810);
and U2810 (N_2810,N_2329,N_2344);
nand U2811 (N_2811,N_1624,N_2081);
or U2812 (N_2812,N_2173,N_1811);
and U2813 (N_2813,N_1858,N_1922);
or U2814 (N_2814,N_1810,N_2105);
nand U2815 (N_2815,N_1621,N_1853);
nand U2816 (N_2816,N_1883,N_1958);
and U2817 (N_2817,N_2395,N_2137);
and U2818 (N_2818,N_2044,N_1744);
nand U2819 (N_2819,N_2221,N_1647);
nand U2820 (N_2820,N_2259,N_1953);
or U2821 (N_2821,N_1909,N_2034);
nor U2822 (N_2822,N_1664,N_1989);
or U2823 (N_2823,N_2266,N_2340);
and U2824 (N_2824,N_2269,N_2266);
nor U2825 (N_2825,N_1612,N_2167);
or U2826 (N_2826,N_2275,N_2025);
and U2827 (N_2827,N_2315,N_2196);
or U2828 (N_2828,N_1689,N_2213);
nand U2829 (N_2829,N_2267,N_1787);
and U2830 (N_2830,N_2011,N_2199);
nand U2831 (N_2831,N_2229,N_2140);
nand U2832 (N_2832,N_1830,N_2150);
nand U2833 (N_2833,N_1683,N_1975);
nor U2834 (N_2834,N_2309,N_1793);
nand U2835 (N_2835,N_1871,N_1737);
xor U2836 (N_2836,N_1795,N_2373);
xor U2837 (N_2837,N_1971,N_1702);
nand U2838 (N_2838,N_2181,N_1877);
nor U2839 (N_2839,N_2364,N_1987);
and U2840 (N_2840,N_1703,N_2321);
or U2841 (N_2841,N_1963,N_2022);
or U2842 (N_2842,N_2038,N_2151);
nand U2843 (N_2843,N_1665,N_1677);
nor U2844 (N_2844,N_2119,N_1727);
xor U2845 (N_2845,N_1645,N_2396);
nor U2846 (N_2846,N_2136,N_1824);
or U2847 (N_2847,N_2329,N_1611);
or U2848 (N_2848,N_1903,N_1970);
or U2849 (N_2849,N_2290,N_2208);
nor U2850 (N_2850,N_1791,N_1747);
xor U2851 (N_2851,N_1723,N_1786);
and U2852 (N_2852,N_2217,N_2091);
xnor U2853 (N_2853,N_1706,N_2015);
or U2854 (N_2854,N_2224,N_2380);
or U2855 (N_2855,N_2144,N_2170);
and U2856 (N_2856,N_2252,N_1657);
or U2857 (N_2857,N_2097,N_2320);
nand U2858 (N_2858,N_2366,N_2105);
nor U2859 (N_2859,N_2098,N_1881);
nor U2860 (N_2860,N_2120,N_2154);
or U2861 (N_2861,N_1938,N_1609);
and U2862 (N_2862,N_2310,N_1854);
nand U2863 (N_2863,N_1720,N_1753);
and U2864 (N_2864,N_2281,N_2245);
xor U2865 (N_2865,N_2393,N_1651);
xor U2866 (N_2866,N_1845,N_2262);
and U2867 (N_2867,N_1716,N_2135);
nand U2868 (N_2868,N_2082,N_1687);
and U2869 (N_2869,N_1786,N_1662);
and U2870 (N_2870,N_1836,N_2290);
nor U2871 (N_2871,N_1866,N_2269);
xor U2872 (N_2872,N_2020,N_2150);
xnor U2873 (N_2873,N_2133,N_1911);
nor U2874 (N_2874,N_1719,N_1928);
and U2875 (N_2875,N_1659,N_2065);
nor U2876 (N_2876,N_2316,N_1651);
nor U2877 (N_2877,N_1699,N_2103);
xor U2878 (N_2878,N_2131,N_2257);
nor U2879 (N_2879,N_2218,N_2372);
nand U2880 (N_2880,N_1611,N_1924);
and U2881 (N_2881,N_1857,N_2369);
or U2882 (N_2882,N_2159,N_2227);
xor U2883 (N_2883,N_2004,N_2315);
or U2884 (N_2884,N_2158,N_2380);
nand U2885 (N_2885,N_1979,N_1982);
or U2886 (N_2886,N_1770,N_2262);
nand U2887 (N_2887,N_1756,N_1614);
xor U2888 (N_2888,N_1806,N_2151);
or U2889 (N_2889,N_2163,N_2191);
nand U2890 (N_2890,N_1989,N_2386);
and U2891 (N_2891,N_1896,N_1880);
xor U2892 (N_2892,N_1942,N_1997);
nand U2893 (N_2893,N_1726,N_1996);
xor U2894 (N_2894,N_2293,N_2217);
or U2895 (N_2895,N_1748,N_2317);
and U2896 (N_2896,N_1734,N_1976);
nand U2897 (N_2897,N_1916,N_2332);
xor U2898 (N_2898,N_1802,N_1990);
nor U2899 (N_2899,N_1666,N_2066);
nor U2900 (N_2900,N_2022,N_1866);
nor U2901 (N_2901,N_2231,N_2296);
nand U2902 (N_2902,N_2287,N_2032);
nand U2903 (N_2903,N_1697,N_2263);
xor U2904 (N_2904,N_1644,N_1979);
nor U2905 (N_2905,N_2129,N_1707);
nand U2906 (N_2906,N_2181,N_2245);
and U2907 (N_2907,N_1935,N_1661);
nor U2908 (N_2908,N_2347,N_1628);
nand U2909 (N_2909,N_2376,N_2287);
nand U2910 (N_2910,N_2103,N_2362);
xor U2911 (N_2911,N_1979,N_1868);
nand U2912 (N_2912,N_2344,N_2185);
xnor U2913 (N_2913,N_1956,N_2120);
nor U2914 (N_2914,N_2208,N_1675);
and U2915 (N_2915,N_1851,N_2305);
and U2916 (N_2916,N_1906,N_2330);
or U2917 (N_2917,N_1828,N_1901);
and U2918 (N_2918,N_2261,N_2227);
nand U2919 (N_2919,N_2371,N_1825);
xnor U2920 (N_2920,N_1906,N_1600);
nor U2921 (N_2921,N_2263,N_1710);
and U2922 (N_2922,N_1639,N_2070);
nand U2923 (N_2923,N_1995,N_1761);
nor U2924 (N_2924,N_1941,N_1656);
nand U2925 (N_2925,N_2228,N_1627);
nand U2926 (N_2926,N_1989,N_1928);
nand U2927 (N_2927,N_2102,N_1967);
xor U2928 (N_2928,N_2243,N_2344);
and U2929 (N_2929,N_1622,N_1766);
and U2930 (N_2930,N_2044,N_1716);
nor U2931 (N_2931,N_1964,N_1616);
nor U2932 (N_2932,N_1910,N_1662);
nor U2933 (N_2933,N_2294,N_1682);
and U2934 (N_2934,N_1857,N_1850);
nor U2935 (N_2935,N_2081,N_1714);
or U2936 (N_2936,N_2327,N_2306);
nor U2937 (N_2937,N_1718,N_1873);
or U2938 (N_2938,N_2323,N_1692);
or U2939 (N_2939,N_1790,N_2071);
nand U2940 (N_2940,N_2347,N_1651);
nand U2941 (N_2941,N_2292,N_2379);
or U2942 (N_2942,N_2220,N_2240);
and U2943 (N_2943,N_2066,N_1678);
or U2944 (N_2944,N_1660,N_2295);
xor U2945 (N_2945,N_1611,N_2262);
and U2946 (N_2946,N_1806,N_2251);
and U2947 (N_2947,N_1689,N_2316);
or U2948 (N_2948,N_2336,N_1644);
and U2949 (N_2949,N_2159,N_2031);
nand U2950 (N_2950,N_2227,N_1744);
xnor U2951 (N_2951,N_1854,N_2106);
xor U2952 (N_2952,N_1994,N_1997);
nand U2953 (N_2953,N_2339,N_1956);
nor U2954 (N_2954,N_1877,N_2227);
and U2955 (N_2955,N_1812,N_1966);
nor U2956 (N_2956,N_1705,N_1647);
and U2957 (N_2957,N_2198,N_1901);
or U2958 (N_2958,N_2395,N_2104);
nand U2959 (N_2959,N_2266,N_2229);
nand U2960 (N_2960,N_1959,N_2058);
nor U2961 (N_2961,N_2020,N_1700);
or U2962 (N_2962,N_1849,N_1603);
nor U2963 (N_2963,N_2154,N_1734);
or U2964 (N_2964,N_2198,N_2229);
nand U2965 (N_2965,N_2336,N_1770);
nand U2966 (N_2966,N_1644,N_2069);
and U2967 (N_2967,N_1826,N_1954);
nand U2968 (N_2968,N_1961,N_2126);
nor U2969 (N_2969,N_1622,N_2370);
or U2970 (N_2970,N_1916,N_1680);
nor U2971 (N_2971,N_2394,N_2259);
xor U2972 (N_2972,N_1867,N_2002);
or U2973 (N_2973,N_1675,N_2323);
xnor U2974 (N_2974,N_1670,N_1684);
and U2975 (N_2975,N_1839,N_2279);
and U2976 (N_2976,N_1990,N_1997);
nand U2977 (N_2977,N_1677,N_1737);
or U2978 (N_2978,N_1757,N_1677);
xnor U2979 (N_2979,N_2015,N_1700);
nand U2980 (N_2980,N_2248,N_2053);
or U2981 (N_2981,N_2177,N_2385);
and U2982 (N_2982,N_1962,N_2225);
and U2983 (N_2983,N_1984,N_2314);
nand U2984 (N_2984,N_2048,N_2233);
or U2985 (N_2985,N_1951,N_1939);
or U2986 (N_2986,N_2358,N_1819);
or U2987 (N_2987,N_1697,N_1691);
nand U2988 (N_2988,N_2117,N_2327);
nand U2989 (N_2989,N_2140,N_1663);
and U2990 (N_2990,N_1609,N_1728);
nor U2991 (N_2991,N_1656,N_2140);
nand U2992 (N_2992,N_2148,N_1987);
nor U2993 (N_2993,N_1850,N_2075);
nand U2994 (N_2994,N_2328,N_2233);
or U2995 (N_2995,N_1733,N_1828);
nand U2996 (N_2996,N_2009,N_2211);
xor U2997 (N_2997,N_2166,N_2331);
nor U2998 (N_2998,N_2280,N_1841);
xnor U2999 (N_2999,N_1897,N_1837);
nand U3000 (N_3000,N_1625,N_2215);
xnor U3001 (N_3001,N_1959,N_2366);
nand U3002 (N_3002,N_1664,N_1822);
xor U3003 (N_3003,N_1785,N_1670);
xnor U3004 (N_3004,N_1898,N_1693);
nand U3005 (N_3005,N_2351,N_2018);
nand U3006 (N_3006,N_1840,N_1714);
and U3007 (N_3007,N_2087,N_1763);
or U3008 (N_3008,N_1951,N_1878);
and U3009 (N_3009,N_1836,N_2308);
and U3010 (N_3010,N_2311,N_2009);
nor U3011 (N_3011,N_1922,N_1766);
nand U3012 (N_3012,N_2196,N_1669);
nor U3013 (N_3013,N_2300,N_1621);
and U3014 (N_3014,N_1796,N_2216);
nand U3015 (N_3015,N_1941,N_1951);
nor U3016 (N_3016,N_1754,N_1802);
nand U3017 (N_3017,N_2330,N_2107);
and U3018 (N_3018,N_2089,N_2357);
nand U3019 (N_3019,N_1959,N_1891);
or U3020 (N_3020,N_1630,N_1610);
or U3021 (N_3021,N_2360,N_1770);
and U3022 (N_3022,N_1755,N_2182);
xnor U3023 (N_3023,N_1757,N_2180);
or U3024 (N_3024,N_2058,N_1717);
xor U3025 (N_3025,N_2174,N_1854);
nor U3026 (N_3026,N_2181,N_2103);
nand U3027 (N_3027,N_2287,N_2295);
nand U3028 (N_3028,N_1622,N_1656);
nand U3029 (N_3029,N_2366,N_1931);
nor U3030 (N_3030,N_1812,N_2025);
nand U3031 (N_3031,N_2328,N_1935);
and U3032 (N_3032,N_2394,N_2111);
xnor U3033 (N_3033,N_2387,N_2374);
or U3034 (N_3034,N_2062,N_2143);
nor U3035 (N_3035,N_2203,N_1863);
or U3036 (N_3036,N_2041,N_2130);
xor U3037 (N_3037,N_2194,N_1662);
xnor U3038 (N_3038,N_2200,N_2304);
and U3039 (N_3039,N_2164,N_2332);
nor U3040 (N_3040,N_2356,N_1715);
and U3041 (N_3041,N_1991,N_1862);
or U3042 (N_3042,N_1866,N_1801);
nor U3043 (N_3043,N_1975,N_1636);
or U3044 (N_3044,N_1748,N_1694);
nor U3045 (N_3045,N_1703,N_1976);
nor U3046 (N_3046,N_2200,N_2156);
xnor U3047 (N_3047,N_1844,N_1962);
xor U3048 (N_3048,N_2250,N_2396);
or U3049 (N_3049,N_2286,N_1973);
nand U3050 (N_3050,N_2053,N_1818);
nor U3051 (N_3051,N_2241,N_2030);
and U3052 (N_3052,N_1819,N_2056);
or U3053 (N_3053,N_1604,N_1680);
nand U3054 (N_3054,N_1689,N_1894);
nand U3055 (N_3055,N_1841,N_2304);
nand U3056 (N_3056,N_2219,N_1746);
nand U3057 (N_3057,N_1946,N_2357);
nand U3058 (N_3058,N_1795,N_1898);
nand U3059 (N_3059,N_1634,N_1820);
nor U3060 (N_3060,N_2059,N_2351);
and U3061 (N_3061,N_2332,N_2292);
and U3062 (N_3062,N_2078,N_2135);
nand U3063 (N_3063,N_2257,N_1922);
and U3064 (N_3064,N_2399,N_1695);
nand U3065 (N_3065,N_2325,N_1709);
or U3066 (N_3066,N_1887,N_2166);
or U3067 (N_3067,N_2020,N_2247);
or U3068 (N_3068,N_1948,N_1795);
nor U3069 (N_3069,N_1622,N_2060);
or U3070 (N_3070,N_2284,N_1804);
or U3071 (N_3071,N_1619,N_2238);
or U3072 (N_3072,N_1882,N_2316);
nor U3073 (N_3073,N_2037,N_2032);
or U3074 (N_3074,N_1840,N_2154);
and U3075 (N_3075,N_2206,N_1761);
or U3076 (N_3076,N_2348,N_2031);
or U3077 (N_3077,N_2070,N_1628);
nand U3078 (N_3078,N_1911,N_1671);
nand U3079 (N_3079,N_2150,N_1805);
and U3080 (N_3080,N_2031,N_2324);
nand U3081 (N_3081,N_2356,N_2258);
nand U3082 (N_3082,N_1842,N_1933);
nor U3083 (N_3083,N_1734,N_2393);
nand U3084 (N_3084,N_1684,N_1997);
xnor U3085 (N_3085,N_2191,N_1991);
nor U3086 (N_3086,N_1707,N_2081);
nor U3087 (N_3087,N_2055,N_1765);
or U3088 (N_3088,N_2134,N_2278);
xnor U3089 (N_3089,N_1822,N_2262);
or U3090 (N_3090,N_1816,N_1831);
and U3091 (N_3091,N_1836,N_2334);
or U3092 (N_3092,N_1908,N_2150);
nor U3093 (N_3093,N_2223,N_1719);
and U3094 (N_3094,N_1950,N_1670);
nor U3095 (N_3095,N_1699,N_2055);
nand U3096 (N_3096,N_2358,N_2179);
nand U3097 (N_3097,N_2137,N_1941);
xor U3098 (N_3098,N_2303,N_1913);
and U3099 (N_3099,N_2057,N_1773);
and U3100 (N_3100,N_1785,N_2140);
and U3101 (N_3101,N_2203,N_2129);
and U3102 (N_3102,N_2220,N_1676);
xor U3103 (N_3103,N_2155,N_1642);
nor U3104 (N_3104,N_2140,N_1727);
nor U3105 (N_3105,N_2299,N_2111);
or U3106 (N_3106,N_2395,N_1875);
nand U3107 (N_3107,N_1947,N_1689);
nand U3108 (N_3108,N_2383,N_2282);
and U3109 (N_3109,N_1643,N_1717);
xnor U3110 (N_3110,N_2311,N_1826);
nor U3111 (N_3111,N_1808,N_2270);
xor U3112 (N_3112,N_1614,N_2297);
and U3113 (N_3113,N_2116,N_1611);
nor U3114 (N_3114,N_2075,N_1625);
nor U3115 (N_3115,N_2166,N_1708);
or U3116 (N_3116,N_2344,N_1867);
and U3117 (N_3117,N_2053,N_2111);
nand U3118 (N_3118,N_2110,N_1992);
nand U3119 (N_3119,N_1813,N_2335);
and U3120 (N_3120,N_2158,N_2379);
nand U3121 (N_3121,N_2386,N_2034);
or U3122 (N_3122,N_1936,N_1764);
nor U3123 (N_3123,N_2332,N_2318);
or U3124 (N_3124,N_2244,N_2086);
nand U3125 (N_3125,N_2391,N_2235);
nor U3126 (N_3126,N_2090,N_1653);
nor U3127 (N_3127,N_1854,N_1610);
xnor U3128 (N_3128,N_1679,N_1693);
xnor U3129 (N_3129,N_2078,N_1677);
or U3130 (N_3130,N_2120,N_2231);
or U3131 (N_3131,N_2046,N_2160);
or U3132 (N_3132,N_2386,N_2330);
and U3133 (N_3133,N_1805,N_2246);
and U3134 (N_3134,N_1705,N_2120);
nor U3135 (N_3135,N_1752,N_1833);
nor U3136 (N_3136,N_2085,N_2106);
and U3137 (N_3137,N_2163,N_2320);
and U3138 (N_3138,N_2240,N_2221);
nor U3139 (N_3139,N_2011,N_1851);
and U3140 (N_3140,N_2222,N_1986);
or U3141 (N_3141,N_2107,N_2317);
xor U3142 (N_3142,N_2000,N_1631);
nand U3143 (N_3143,N_1783,N_1772);
xnor U3144 (N_3144,N_1716,N_1893);
nand U3145 (N_3145,N_1772,N_1856);
xnor U3146 (N_3146,N_1786,N_2345);
or U3147 (N_3147,N_2110,N_1635);
nand U3148 (N_3148,N_1963,N_1845);
nand U3149 (N_3149,N_2025,N_2282);
nand U3150 (N_3150,N_2156,N_2242);
and U3151 (N_3151,N_2059,N_2335);
nand U3152 (N_3152,N_1967,N_2059);
xor U3153 (N_3153,N_1651,N_1870);
nor U3154 (N_3154,N_2220,N_1698);
nor U3155 (N_3155,N_1604,N_1972);
nor U3156 (N_3156,N_2217,N_1915);
and U3157 (N_3157,N_1725,N_2036);
nor U3158 (N_3158,N_1696,N_1704);
and U3159 (N_3159,N_2222,N_1991);
and U3160 (N_3160,N_2332,N_1727);
xor U3161 (N_3161,N_2087,N_2309);
and U3162 (N_3162,N_1825,N_2242);
and U3163 (N_3163,N_2032,N_2281);
or U3164 (N_3164,N_1990,N_2207);
and U3165 (N_3165,N_2128,N_2286);
or U3166 (N_3166,N_1686,N_1892);
nand U3167 (N_3167,N_2230,N_2217);
nor U3168 (N_3168,N_1608,N_1872);
nor U3169 (N_3169,N_2146,N_1894);
or U3170 (N_3170,N_2340,N_1688);
or U3171 (N_3171,N_2245,N_2356);
nor U3172 (N_3172,N_2294,N_2068);
nand U3173 (N_3173,N_2084,N_2310);
xnor U3174 (N_3174,N_2366,N_2195);
and U3175 (N_3175,N_1755,N_1611);
nor U3176 (N_3176,N_1724,N_1934);
nand U3177 (N_3177,N_1650,N_2392);
nor U3178 (N_3178,N_2268,N_2023);
nand U3179 (N_3179,N_1764,N_2262);
nor U3180 (N_3180,N_2042,N_2131);
or U3181 (N_3181,N_1681,N_2278);
or U3182 (N_3182,N_1836,N_1669);
nor U3183 (N_3183,N_1751,N_1697);
nor U3184 (N_3184,N_1910,N_2102);
xor U3185 (N_3185,N_1821,N_1979);
or U3186 (N_3186,N_2380,N_2391);
and U3187 (N_3187,N_2191,N_1880);
or U3188 (N_3188,N_1946,N_1827);
and U3189 (N_3189,N_2245,N_1638);
nor U3190 (N_3190,N_2187,N_2073);
nor U3191 (N_3191,N_2086,N_2135);
or U3192 (N_3192,N_2172,N_1701);
and U3193 (N_3193,N_2245,N_1929);
nor U3194 (N_3194,N_2083,N_2354);
nor U3195 (N_3195,N_2097,N_1827);
xnor U3196 (N_3196,N_2126,N_1801);
and U3197 (N_3197,N_2375,N_1862);
xnor U3198 (N_3198,N_2305,N_2035);
nand U3199 (N_3199,N_1612,N_2002);
xnor U3200 (N_3200,N_3026,N_2516);
nand U3201 (N_3201,N_3064,N_2881);
or U3202 (N_3202,N_2483,N_3023);
xnor U3203 (N_3203,N_2811,N_2755);
nand U3204 (N_3204,N_2757,N_2707);
nand U3205 (N_3205,N_3028,N_3097);
nor U3206 (N_3206,N_2851,N_2688);
or U3207 (N_3207,N_2526,N_2415);
xor U3208 (N_3208,N_3124,N_2865);
and U3209 (N_3209,N_2775,N_2787);
nand U3210 (N_3210,N_2424,N_2654);
and U3211 (N_3211,N_2511,N_3132);
or U3212 (N_3212,N_2763,N_3082);
and U3213 (N_3213,N_2978,N_2842);
and U3214 (N_3214,N_2721,N_2886);
nor U3215 (N_3215,N_3025,N_2653);
nor U3216 (N_3216,N_2670,N_2446);
xnor U3217 (N_3217,N_3105,N_3162);
and U3218 (N_3218,N_2910,N_2841);
or U3219 (N_3219,N_2783,N_3004);
or U3220 (N_3220,N_2436,N_3088);
nand U3221 (N_3221,N_2805,N_3080);
and U3222 (N_3222,N_2590,N_2856);
and U3223 (N_3223,N_2903,N_2835);
and U3224 (N_3224,N_2573,N_2403);
and U3225 (N_3225,N_2990,N_3012);
nand U3226 (N_3226,N_2419,N_2955);
nand U3227 (N_3227,N_2433,N_2826);
or U3228 (N_3228,N_3065,N_3079);
or U3229 (N_3229,N_2977,N_2912);
xnor U3230 (N_3230,N_2494,N_2488);
xnor U3231 (N_3231,N_2742,N_2777);
and U3232 (N_3232,N_3147,N_2413);
nor U3233 (N_3233,N_2497,N_2411);
or U3234 (N_3234,N_2523,N_2578);
and U3235 (N_3235,N_2723,N_2822);
and U3236 (N_3236,N_3129,N_2678);
and U3237 (N_3237,N_2510,N_2830);
xor U3238 (N_3238,N_2458,N_3145);
xnor U3239 (N_3239,N_2999,N_2871);
xnor U3240 (N_3240,N_3178,N_3019);
and U3241 (N_3241,N_2480,N_3030);
nor U3242 (N_3242,N_3165,N_2652);
nand U3243 (N_3243,N_2496,N_2529);
or U3244 (N_3244,N_2569,N_2612);
nor U3245 (N_3245,N_2854,N_2767);
or U3246 (N_3246,N_2741,N_3137);
nor U3247 (N_3247,N_3160,N_2878);
and U3248 (N_3248,N_2768,N_3052);
or U3249 (N_3249,N_2486,N_2710);
xnor U3250 (N_3250,N_3094,N_2778);
xor U3251 (N_3251,N_3121,N_3152);
xor U3252 (N_3252,N_3133,N_2400);
nor U3253 (N_3253,N_2925,N_3143);
and U3254 (N_3254,N_2607,N_3078);
xor U3255 (N_3255,N_2979,N_2543);
or U3256 (N_3256,N_2490,N_2837);
or U3257 (N_3257,N_3157,N_2535);
nor U3258 (N_3258,N_3060,N_2551);
and U3259 (N_3259,N_3135,N_2662);
nor U3260 (N_3260,N_2565,N_2816);
nand U3261 (N_3261,N_2439,N_2421);
nand U3262 (N_3262,N_3044,N_2997);
nand U3263 (N_3263,N_3081,N_2457);
or U3264 (N_3264,N_2725,N_2857);
xor U3265 (N_3265,N_2638,N_2471);
or U3266 (N_3266,N_2584,N_3122);
xor U3267 (N_3267,N_2926,N_2795);
nor U3268 (N_3268,N_3182,N_3036);
and U3269 (N_3269,N_2452,N_3013);
nand U3270 (N_3270,N_2771,N_3130);
nor U3271 (N_3271,N_2624,N_3051);
or U3272 (N_3272,N_2530,N_2637);
xnor U3273 (N_3273,N_2639,N_3144);
or U3274 (N_3274,N_2834,N_3022);
or U3275 (N_3275,N_3155,N_2736);
nand U3276 (N_3276,N_2524,N_2823);
nor U3277 (N_3277,N_2727,N_2579);
or U3278 (N_3278,N_2924,N_2769);
or U3279 (N_3279,N_2527,N_2459);
or U3280 (N_3280,N_3008,N_2525);
or U3281 (N_3281,N_2939,N_2897);
or U3282 (N_3282,N_2713,N_2942);
xor U3283 (N_3283,N_2562,N_2934);
xor U3284 (N_3284,N_2809,N_3007);
xnor U3285 (N_3285,N_3168,N_3126);
nand U3286 (N_3286,N_2532,N_2405);
xnor U3287 (N_3287,N_3016,N_2738);
nor U3288 (N_3288,N_2862,N_3125);
or U3289 (N_3289,N_2583,N_3164);
and U3290 (N_3290,N_2460,N_2949);
nand U3291 (N_3291,N_2882,N_2784);
nand U3292 (N_3292,N_2967,N_2613);
nand U3293 (N_3293,N_2920,N_3106);
or U3294 (N_3294,N_2689,N_2675);
nor U3295 (N_3295,N_2941,N_2981);
xor U3296 (N_3296,N_2517,N_3111);
xnor U3297 (N_3297,N_3173,N_3046);
and U3298 (N_3298,N_3110,N_2895);
nand U3299 (N_3299,N_2695,N_3159);
and U3300 (N_3300,N_2616,N_2976);
or U3301 (N_3301,N_2799,N_2476);
and U3302 (N_3302,N_2699,N_2968);
and U3303 (N_3303,N_2776,N_3090);
nor U3304 (N_3304,N_2683,N_2940);
nand U3305 (N_3305,N_3139,N_2748);
and U3306 (N_3306,N_2863,N_3072);
nor U3307 (N_3307,N_2916,N_2921);
or U3308 (N_3308,N_2845,N_3181);
and U3309 (N_3309,N_2447,N_2853);
and U3310 (N_3310,N_2847,N_2644);
or U3311 (N_3311,N_3043,N_2404);
and U3312 (N_3312,N_2720,N_2745);
xor U3313 (N_3313,N_2900,N_2766);
and U3314 (N_3314,N_2450,N_2765);
nand U3315 (N_3315,N_2614,N_2697);
nor U3316 (N_3316,N_3010,N_2541);
or U3317 (N_3317,N_2883,N_2589);
xnor U3318 (N_3318,N_3116,N_3069);
xor U3319 (N_3319,N_2866,N_2894);
xor U3320 (N_3320,N_2849,N_2819);
and U3321 (N_3321,N_2455,N_2625);
nor U3322 (N_3322,N_3154,N_2434);
and U3323 (N_3323,N_2761,N_3120);
nor U3324 (N_3324,N_2576,N_3141);
or U3325 (N_3325,N_3179,N_2571);
nor U3326 (N_3326,N_2703,N_2575);
nand U3327 (N_3327,N_2509,N_2864);
nor U3328 (N_3328,N_2453,N_2566);
xor U3329 (N_3329,N_3146,N_2500);
xnor U3330 (N_3330,N_2982,N_2658);
nor U3331 (N_3331,N_2611,N_2595);
nand U3332 (N_3332,N_2706,N_2915);
xnor U3333 (N_3333,N_2868,N_2686);
nand U3334 (N_3334,N_2779,N_3188);
nor U3335 (N_3335,N_2892,N_2615);
xnor U3336 (N_3336,N_2513,N_3114);
nor U3337 (N_3337,N_2563,N_3033);
nand U3338 (N_3338,N_3180,N_2512);
or U3339 (N_3339,N_2508,N_2520);
xor U3340 (N_3340,N_2759,N_2729);
nand U3341 (N_3341,N_3005,N_2793);
and U3342 (N_3342,N_2893,N_2665);
or U3343 (N_3343,N_2993,N_3170);
or U3344 (N_3344,N_2591,N_3134);
and U3345 (N_3345,N_3039,N_2682);
or U3346 (N_3346,N_2609,N_2429);
nor U3347 (N_3347,N_2917,N_2632);
nand U3348 (N_3348,N_2617,N_2998);
nor U3349 (N_3349,N_2598,N_2904);
nand U3350 (N_3350,N_2676,N_3193);
or U3351 (N_3351,N_2531,N_2971);
and U3352 (N_3352,N_2909,N_2807);
nor U3353 (N_3353,N_2600,N_3042);
nor U3354 (N_3354,N_2561,N_2974);
xor U3355 (N_3355,N_2740,N_2972);
nand U3356 (N_3356,N_2728,N_3040);
nand U3357 (N_3357,N_3045,N_2827);
nand U3358 (N_3358,N_2786,N_2908);
nand U3359 (N_3359,N_2973,N_2604);
nand U3360 (N_3360,N_3186,N_3057);
nor U3361 (N_3361,N_2952,N_2664);
xnor U3362 (N_3362,N_3029,N_3108);
nand U3363 (N_3363,N_3015,N_3076);
nor U3364 (N_3364,N_2933,N_2691);
and U3365 (N_3365,N_3075,N_2495);
xor U3366 (N_3366,N_2582,N_2422);
xor U3367 (N_3367,N_3190,N_2431);
and U3368 (N_3368,N_2770,N_3103);
or U3369 (N_3369,N_3068,N_3021);
nand U3370 (N_3370,N_2409,N_2420);
and U3371 (N_3371,N_2680,N_3092);
or U3372 (N_3372,N_2712,N_3140);
xnor U3373 (N_3373,N_2923,N_2645);
nand U3374 (N_3374,N_2959,N_2461);
nand U3375 (N_3375,N_2482,N_2756);
nor U3376 (N_3376,N_3037,N_2467);
nand U3377 (N_3377,N_2626,N_2760);
nand U3378 (N_3378,N_2628,N_2839);
and U3379 (N_3379,N_2465,N_3171);
nand U3380 (N_3380,N_3095,N_2487);
nor U3381 (N_3381,N_2618,N_3032);
or U3382 (N_3382,N_2679,N_2674);
and U3383 (N_3383,N_2430,N_3050);
and U3384 (N_3384,N_2666,N_2550);
xor U3385 (N_3385,N_2965,N_2634);
or U3386 (N_3386,N_2648,N_2454);
or U3387 (N_3387,N_2813,N_3070);
xnor U3388 (N_3388,N_2717,N_2947);
or U3389 (N_3389,N_2463,N_3098);
or U3390 (N_3390,N_2521,N_2891);
and U3391 (N_3391,N_2899,N_2432);
nor U3392 (N_3392,N_3198,N_2929);
xnor U3393 (N_3393,N_2410,N_2928);
and U3394 (N_3394,N_2859,N_2623);
xor U3395 (N_3395,N_3011,N_3151);
xnor U3396 (N_3396,N_3192,N_3018);
xnor U3397 (N_3397,N_2522,N_2715);
xnor U3398 (N_3398,N_2440,N_2414);
and U3399 (N_3399,N_2696,N_2442);
xnor U3400 (N_3400,N_2806,N_3074);
and U3401 (N_3401,N_2661,N_2448);
nand U3402 (N_3402,N_2983,N_2681);
xor U3403 (N_3403,N_2630,N_2518);
or U3404 (N_3404,N_2962,N_2451);
and U3405 (N_3405,N_2547,N_2602);
nor U3406 (N_3406,N_2701,N_3194);
and U3407 (N_3407,N_2650,N_2427);
nand U3408 (N_3408,N_2796,N_2758);
nand U3409 (N_3409,N_3142,N_3183);
nand U3410 (N_3410,N_3104,N_2629);
nor U3411 (N_3411,N_2441,N_2633);
and U3412 (N_3412,N_2656,N_2764);
nand U3413 (N_3413,N_2491,N_2534);
nand U3414 (N_3414,N_2836,N_2533);
xor U3415 (N_3415,N_2724,N_2426);
and U3416 (N_3416,N_2594,N_2911);
xor U3417 (N_3417,N_2961,N_2515);
xnor U3418 (N_3418,N_3002,N_3112);
nor U3419 (N_3419,N_3077,N_2671);
nand U3420 (N_3420,N_2672,N_2705);
and U3421 (N_3421,N_2870,N_2580);
nor U3422 (N_3422,N_2744,N_2821);
nor U3423 (N_3423,N_2781,N_2660);
and U3424 (N_3424,N_2466,N_2558);
and U3425 (N_3425,N_2931,N_2810);
nor U3426 (N_3426,N_2732,N_3009);
and U3427 (N_3427,N_2860,N_3163);
xnor U3428 (N_3428,N_2873,N_2640);
nand U3429 (N_3429,N_3199,N_2889);
nor U3430 (N_3430,N_2932,N_2984);
nor U3431 (N_3431,N_2473,N_2647);
nand U3432 (N_3432,N_2872,N_2840);
nor U3433 (N_3433,N_3059,N_2946);
nor U3434 (N_3434,N_2754,N_2995);
nor U3435 (N_3435,N_2449,N_2970);
or U3436 (N_3436,N_2443,N_2407);
and U3437 (N_3437,N_2479,N_2601);
or U3438 (N_3438,N_2782,N_2503);
and U3439 (N_3439,N_2791,N_3093);
nand U3440 (N_3440,N_2416,N_2985);
nor U3441 (N_3441,N_3066,N_2966);
and U3442 (N_3442,N_2850,N_2504);
nor U3443 (N_3443,N_2627,N_2673);
nor U3444 (N_3444,N_2846,N_2991);
nand U3445 (N_3445,N_2867,N_3071);
and U3446 (N_3446,N_3156,N_2798);
nand U3447 (N_3447,N_3020,N_3117);
xnor U3448 (N_3448,N_2668,N_2501);
nor U3449 (N_3449,N_2914,N_2718);
nand U3450 (N_3450,N_2749,N_2557);
xnor U3451 (N_3451,N_3027,N_2560);
xnor U3452 (N_3452,N_2708,N_2852);
xor U3453 (N_3453,N_3035,N_3102);
and U3454 (N_3454,N_3091,N_2938);
nand U3455 (N_3455,N_2577,N_2554);
and U3456 (N_3456,N_2989,N_2537);
and U3457 (N_3457,N_3172,N_2963);
nand U3458 (N_3458,N_2772,N_3089);
nand U3459 (N_3459,N_3197,N_2622);
and U3460 (N_3460,N_2502,N_2901);
and U3461 (N_3461,N_2536,N_2519);
nand U3462 (N_3462,N_3148,N_2722);
or U3463 (N_3463,N_2499,N_2657);
and U3464 (N_3464,N_2437,N_2975);
and U3465 (N_3465,N_3149,N_2788);
xor U3466 (N_3466,N_2667,N_2472);
or U3467 (N_3467,N_2631,N_3085);
nand U3468 (N_3468,N_2737,N_2980);
xnor U3469 (N_3469,N_2542,N_2719);
and U3470 (N_3470,N_2743,N_3123);
nand U3471 (N_3471,N_2789,N_2462);
xor U3472 (N_3472,N_2954,N_3115);
nor U3473 (N_3473,N_3061,N_3100);
and U3474 (N_3474,N_2879,N_3166);
xor U3475 (N_3475,N_3063,N_2877);
and U3476 (N_3476,N_2762,N_2858);
and U3477 (N_3477,N_2774,N_2956);
nand U3478 (N_3478,N_2960,N_2545);
nand U3479 (N_3479,N_2444,N_2481);
xor U3480 (N_3480,N_2651,N_2876);
xor U3481 (N_3481,N_3196,N_2478);
xor U3482 (N_3482,N_2733,N_3056);
nand U3483 (N_3483,N_2425,N_2548);
nand U3484 (N_3484,N_2546,N_2553);
or U3485 (N_3485,N_2825,N_2555);
and U3486 (N_3486,N_2552,N_2890);
nor U3487 (N_3487,N_3048,N_2418);
nor U3488 (N_3488,N_2669,N_2913);
and U3489 (N_3489,N_2572,N_2642);
or U3490 (N_3490,N_2731,N_2606);
nor U3491 (N_3491,N_2935,N_3049);
and U3492 (N_3492,N_2588,N_2704);
or U3493 (N_3493,N_2636,N_2474);
or U3494 (N_3494,N_3158,N_3189);
xnor U3495 (N_3495,N_2988,N_3001);
nand U3496 (N_3496,N_2953,N_2401);
or U3497 (N_3497,N_2655,N_2423);
nor U3498 (N_3498,N_2620,N_3054);
xnor U3499 (N_3499,N_2898,N_2659);
nor U3500 (N_3500,N_2752,N_3161);
xnor U3501 (N_3501,N_3119,N_2751);
nand U3502 (N_3502,N_2726,N_2937);
and U3503 (N_3503,N_2568,N_2570);
xnor U3504 (N_3504,N_2693,N_2801);
or U3505 (N_3505,N_2790,N_2700);
nand U3506 (N_3506,N_3041,N_2994);
nand U3507 (N_3507,N_2874,N_2567);
or U3508 (N_3508,N_2484,N_3138);
and U3509 (N_3509,N_2498,N_3169);
nand U3510 (N_3510,N_3031,N_2702);
nor U3511 (N_3511,N_3003,N_2599);
nand U3512 (N_3512,N_2564,N_2435);
nor U3513 (N_3513,N_2730,N_2818);
nor U3514 (N_3514,N_2875,N_2944);
xor U3515 (N_3515,N_2888,N_3109);
nand U3516 (N_3516,N_2586,N_2957);
and U3517 (N_3517,N_3127,N_2687);
nand U3518 (N_3518,N_3017,N_2986);
nor U3519 (N_3519,N_3167,N_3086);
or U3520 (N_3520,N_3153,N_2469);
or U3521 (N_3521,N_2643,N_2677);
nor U3522 (N_3522,N_3038,N_2815);
or U3523 (N_3523,N_2750,N_3174);
nor U3524 (N_3524,N_3024,N_2848);
nor U3525 (N_3525,N_2597,N_2906);
nor U3526 (N_3526,N_3073,N_2663);
nor U3527 (N_3527,N_3101,N_2907);
nand U3528 (N_3528,N_2538,N_2896);
nor U3529 (N_3529,N_2649,N_2549);
and U3530 (N_3530,N_2887,N_3176);
and U3531 (N_3531,N_3083,N_2610);
nor U3532 (N_3532,N_2746,N_2605);
and U3533 (N_3533,N_3087,N_2804);
or U3534 (N_3534,N_2950,N_2685);
nor U3535 (N_3535,N_2641,N_2922);
nor U3536 (N_3536,N_2540,N_3184);
and U3537 (N_3537,N_2714,N_2800);
nor U3538 (N_3538,N_2902,N_2918);
nand U3539 (N_3539,N_2817,N_2820);
or U3540 (N_3540,N_3000,N_2945);
nor U3541 (N_3541,N_2838,N_2828);
nand U3542 (N_3542,N_2844,N_2785);
and U3543 (N_3543,N_2507,N_2843);
nand U3544 (N_3544,N_2803,N_2646);
or U3545 (N_3545,N_2698,N_2797);
or U3546 (N_3546,N_3113,N_3128);
xor U3547 (N_3547,N_2936,N_3185);
and U3548 (N_3548,N_2402,N_2574);
xnor U3549 (N_3549,N_2445,N_2927);
or U3550 (N_3550,N_2493,N_2996);
and U3551 (N_3551,N_2587,N_2619);
nor U3552 (N_3552,N_2506,N_2794);
or U3553 (N_3553,N_2880,N_2930);
nand U3554 (N_3554,N_2958,N_2884);
and U3555 (N_3555,N_3187,N_2753);
nand U3556 (N_3556,N_2919,N_2855);
xor U3557 (N_3557,N_2814,N_2829);
and U3558 (N_3558,N_2812,N_3195);
and U3559 (N_3559,N_2709,N_2694);
and U3560 (N_3560,N_3096,N_2869);
nor U3561 (N_3561,N_2581,N_2585);
nor U3562 (N_3562,N_2539,N_2690);
nand U3563 (N_3563,N_2477,N_2831);
xor U3564 (N_3564,N_2734,N_3191);
or U3565 (N_3565,N_2492,N_2559);
and U3566 (N_3566,N_2684,N_3055);
or U3567 (N_3567,N_3062,N_2438);
nand U3568 (N_3568,N_2861,N_2408);
nor U3569 (N_3569,N_2468,N_2635);
and U3570 (N_3570,N_2808,N_2987);
xor U3571 (N_3571,N_2528,N_2802);
xnor U3572 (N_3572,N_2711,N_2475);
nor U3573 (N_3573,N_2832,N_2792);
or U3574 (N_3574,N_2692,N_3058);
and U3575 (N_3575,N_2948,N_2964);
and U3576 (N_3576,N_3107,N_2992);
xnor U3577 (N_3577,N_3067,N_2505);
nand U3578 (N_3578,N_2406,N_3084);
xnor U3579 (N_3579,N_2470,N_2905);
and U3580 (N_3580,N_2621,N_2544);
nor U3581 (N_3581,N_3175,N_3177);
nor U3582 (N_3582,N_3053,N_2456);
and U3583 (N_3583,N_3099,N_2780);
or U3584 (N_3584,N_3150,N_2951);
or U3585 (N_3585,N_2417,N_2739);
nor U3586 (N_3586,N_3006,N_2824);
and U3587 (N_3587,N_2943,N_2833);
xnor U3588 (N_3588,N_2735,N_2464);
or U3589 (N_3589,N_2556,N_2593);
xor U3590 (N_3590,N_2596,N_2773);
nor U3591 (N_3591,N_2514,N_3014);
nor U3592 (N_3592,N_2485,N_2603);
xnor U3593 (N_3593,N_2592,N_2885);
xnor U3594 (N_3594,N_2747,N_3118);
or U3595 (N_3595,N_3131,N_2716);
or U3596 (N_3596,N_3136,N_2489);
or U3597 (N_3597,N_2969,N_3034);
nand U3598 (N_3598,N_2608,N_2412);
nand U3599 (N_3599,N_2428,N_3047);
xor U3600 (N_3600,N_2649,N_2599);
and U3601 (N_3601,N_2664,N_3043);
xor U3602 (N_3602,N_2411,N_2814);
or U3603 (N_3603,N_2472,N_2440);
and U3604 (N_3604,N_2735,N_2406);
nand U3605 (N_3605,N_2570,N_2734);
and U3606 (N_3606,N_2867,N_2633);
nor U3607 (N_3607,N_2417,N_2643);
nor U3608 (N_3608,N_3120,N_2864);
nor U3609 (N_3609,N_2992,N_2872);
nand U3610 (N_3610,N_3188,N_2903);
nand U3611 (N_3611,N_2972,N_3044);
xnor U3612 (N_3612,N_2917,N_2599);
xor U3613 (N_3613,N_2514,N_2841);
and U3614 (N_3614,N_2879,N_2443);
nor U3615 (N_3615,N_2595,N_3163);
and U3616 (N_3616,N_2451,N_2475);
nand U3617 (N_3617,N_2675,N_3174);
nor U3618 (N_3618,N_2648,N_2626);
xor U3619 (N_3619,N_2902,N_3140);
nand U3620 (N_3620,N_2445,N_2853);
nor U3621 (N_3621,N_3146,N_2557);
xnor U3622 (N_3622,N_2873,N_2912);
xnor U3623 (N_3623,N_2430,N_2435);
or U3624 (N_3624,N_3079,N_3160);
nor U3625 (N_3625,N_2606,N_2406);
nor U3626 (N_3626,N_2421,N_2772);
xnor U3627 (N_3627,N_2611,N_3148);
nand U3628 (N_3628,N_2524,N_3098);
nand U3629 (N_3629,N_2987,N_2761);
or U3630 (N_3630,N_2699,N_2881);
or U3631 (N_3631,N_2419,N_2655);
and U3632 (N_3632,N_2860,N_2649);
xnor U3633 (N_3633,N_2870,N_2897);
or U3634 (N_3634,N_2566,N_2685);
or U3635 (N_3635,N_2839,N_2444);
and U3636 (N_3636,N_3083,N_2582);
or U3637 (N_3637,N_3153,N_2513);
nor U3638 (N_3638,N_2436,N_3075);
and U3639 (N_3639,N_2745,N_2724);
xnor U3640 (N_3640,N_2906,N_2998);
and U3641 (N_3641,N_2855,N_2470);
or U3642 (N_3642,N_3010,N_3097);
xor U3643 (N_3643,N_2971,N_2918);
or U3644 (N_3644,N_3132,N_2986);
nor U3645 (N_3645,N_2986,N_3045);
and U3646 (N_3646,N_3021,N_2403);
nand U3647 (N_3647,N_2472,N_2607);
or U3648 (N_3648,N_2894,N_2427);
or U3649 (N_3649,N_2490,N_2986);
or U3650 (N_3650,N_3198,N_2476);
nand U3651 (N_3651,N_2987,N_3027);
nand U3652 (N_3652,N_2811,N_2628);
or U3653 (N_3653,N_2664,N_3110);
xnor U3654 (N_3654,N_3084,N_2773);
and U3655 (N_3655,N_3192,N_2437);
or U3656 (N_3656,N_2553,N_2472);
and U3657 (N_3657,N_2872,N_2490);
xor U3658 (N_3658,N_2670,N_2918);
and U3659 (N_3659,N_2463,N_2781);
or U3660 (N_3660,N_2696,N_2990);
and U3661 (N_3661,N_2618,N_3144);
or U3662 (N_3662,N_2930,N_2459);
nand U3663 (N_3663,N_2657,N_2787);
nor U3664 (N_3664,N_2847,N_3080);
or U3665 (N_3665,N_2945,N_3122);
nor U3666 (N_3666,N_3192,N_2834);
xnor U3667 (N_3667,N_2979,N_2498);
or U3668 (N_3668,N_2610,N_2674);
or U3669 (N_3669,N_3156,N_2989);
xor U3670 (N_3670,N_2547,N_2509);
nand U3671 (N_3671,N_3006,N_2849);
xor U3672 (N_3672,N_2906,N_2444);
or U3673 (N_3673,N_2861,N_2959);
nor U3674 (N_3674,N_3176,N_3112);
and U3675 (N_3675,N_3105,N_2630);
and U3676 (N_3676,N_2519,N_3019);
nand U3677 (N_3677,N_2426,N_3150);
or U3678 (N_3678,N_2414,N_3149);
or U3679 (N_3679,N_2406,N_2533);
or U3680 (N_3680,N_2841,N_2622);
xor U3681 (N_3681,N_2929,N_2640);
or U3682 (N_3682,N_3052,N_2463);
nor U3683 (N_3683,N_2810,N_3120);
nand U3684 (N_3684,N_3199,N_2725);
or U3685 (N_3685,N_2927,N_2577);
xor U3686 (N_3686,N_2857,N_2411);
nor U3687 (N_3687,N_2822,N_2695);
xor U3688 (N_3688,N_2499,N_2956);
nand U3689 (N_3689,N_3164,N_2535);
and U3690 (N_3690,N_2709,N_2505);
and U3691 (N_3691,N_2554,N_2645);
nand U3692 (N_3692,N_2515,N_2527);
nand U3693 (N_3693,N_2746,N_2618);
xor U3694 (N_3694,N_3147,N_2434);
nand U3695 (N_3695,N_2574,N_2842);
nor U3696 (N_3696,N_2756,N_2713);
or U3697 (N_3697,N_2453,N_2451);
xnor U3698 (N_3698,N_2430,N_2547);
xnor U3699 (N_3699,N_2759,N_2438);
nand U3700 (N_3700,N_2902,N_2947);
and U3701 (N_3701,N_3050,N_2894);
or U3702 (N_3702,N_2412,N_2803);
or U3703 (N_3703,N_3075,N_2910);
nor U3704 (N_3704,N_2784,N_3010);
nor U3705 (N_3705,N_2401,N_3190);
nor U3706 (N_3706,N_2571,N_3122);
or U3707 (N_3707,N_2958,N_2957);
and U3708 (N_3708,N_2573,N_2879);
or U3709 (N_3709,N_2562,N_2511);
nand U3710 (N_3710,N_3198,N_2723);
and U3711 (N_3711,N_2840,N_2903);
or U3712 (N_3712,N_2589,N_2515);
nor U3713 (N_3713,N_2634,N_2801);
xor U3714 (N_3714,N_2608,N_2889);
xnor U3715 (N_3715,N_2437,N_2608);
nand U3716 (N_3716,N_2460,N_2921);
xnor U3717 (N_3717,N_2864,N_2896);
nor U3718 (N_3718,N_3117,N_2756);
nor U3719 (N_3719,N_2471,N_3053);
and U3720 (N_3720,N_2632,N_2424);
xor U3721 (N_3721,N_2718,N_2408);
nor U3722 (N_3722,N_2821,N_2954);
or U3723 (N_3723,N_2985,N_2549);
and U3724 (N_3724,N_2566,N_2861);
or U3725 (N_3725,N_2443,N_2572);
or U3726 (N_3726,N_3156,N_3132);
nand U3727 (N_3727,N_2867,N_3019);
nand U3728 (N_3728,N_2524,N_3018);
or U3729 (N_3729,N_2710,N_3075);
or U3730 (N_3730,N_2981,N_3048);
xnor U3731 (N_3731,N_2587,N_2747);
nand U3732 (N_3732,N_2787,N_3189);
or U3733 (N_3733,N_2828,N_2657);
nor U3734 (N_3734,N_2709,N_2581);
and U3735 (N_3735,N_3094,N_2499);
nand U3736 (N_3736,N_2559,N_2512);
or U3737 (N_3737,N_2744,N_2747);
nor U3738 (N_3738,N_2839,N_2529);
nand U3739 (N_3739,N_2965,N_2787);
nor U3740 (N_3740,N_2884,N_2580);
nor U3741 (N_3741,N_3145,N_2941);
xor U3742 (N_3742,N_2506,N_3178);
and U3743 (N_3743,N_3023,N_2460);
or U3744 (N_3744,N_2565,N_2856);
or U3745 (N_3745,N_2718,N_3085);
xnor U3746 (N_3746,N_3111,N_2897);
and U3747 (N_3747,N_2534,N_2863);
or U3748 (N_3748,N_2423,N_2525);
nor U3749 (N_3749,N_2406,N_2604);
xor U3750 (N_3750,N_2536,N_2849);
nor U3751 (N_3751,N_2731,N_2710);
nor U3752 (N_3752,N_3070,N_2639);
nand U3753 (N_3753,N_3053,N_2715);
xnor U3754 (N_3754,N_2521,N_3159);
nor U3755 (N_3755,N_2585,N_2441);
nand U3756 (N_3756,N_2547,N_2919);
nor U3757 (N_3757,N_2870,N_2670);
xnor U3758 (N_3758,N_2643,N_2759);
and U3759 (N_3759,N_3079,N_2890);
xnor U3760 (N_3760,N_3142,N_2973);
nor U3761 (N_3761,N_2683,N_2976);
nand U3762 (N_3762,N_3173,N_2576);
or U3763 (N_3763,N_2695,N_2436);
and U3764 (N_3764,N_2460,N_3035);
nand U3765 (N_3765,N_2695,N_2612);
nand U3766 (N_3766,N_3161,N_2705);
nor U3767 (N_3767,N_2805,N_2682);
and U3768 (N_3768,N_3056,N_3156);
and U3769 (N_3769,N_2974,N_3135);
nand U3770 (N_3770,N_2963,N_2766);
and U3771 (N_3771,N_2870,N_2853);
nand U3772 (N_3772,N_3099,N_3127);
and U3773 (N_3773,N_2578,N_3014);
and U3774 (N_3774,N_2892,N_2759);
nor U3775 (N_3775,N_2494,N_2803);
nand U3776 (N_3776,N_2834,N_2809);
or U3777 (N_3777,N_3110,N_2536);
nand U3778 (N_3778,N_2553,N_3132);
nor U3779 (N_3779,N_2667,N_2808);
xor U3780 (N_3780,N_3194,N_2599);
nand U3781 (N_3781,N_2502,N_3175);
or U3782 (N_3782,N_2439,N_2514);
or U3783 (N_3783,N_3073,N_2744);
and U3784 (N_3784,N_3083,N_2420);
nor U3785 (N_3785,N_2737,N_3129);
nand U3786 (N_3786,N_2410,N_3097);
or U3787 (N_3787,N_2615,N_2680);
or U3788 (N_3788,N_2625,N_2468);
or U3789 (N_3789,N_2471,N_2456);
nor U3790 (N_3790,N_2685,N_2440);
nand U3791 (N_3791,N_2652,N_2592);
nor U3792 (N_3792,N_3055,N_2635);
and U3793 (N_3793,N_2414,N_2868);
and U3794 (N_3794,N_2925,N_3183);
xnor U3795 (N_3795,N_3008,N_2545);
or U3796 (N_3796,N_2729,N_3122);
and U3797 (N_3797,N_3016,N_2460);
xnor U3798 (N_3798,N_2440,N_2805);
nand U3799 (N_3799,N_3042,N_2572);
xnor U3800 (N_3800,N_2894,N_2586);
nand U3801 (N_3801,N_2619,N_3140);
nand U3802 (N_3802,N_2722,N_2638);
or U3803 (N_3803,N_2671,N_2555);
nor U3804 (N_3804,N_2572,N_3020);
nor U3805 (N_3805,N_2446,N_3181);
and U3806 (N_3806,N_2923,N_3135);
nand U3807 (N_3807,N_3144,N_3086);
nand U3808 (N_3808,N_2545,N_3048);
xor U3809 (N_3809,N_2912,N_2416);
nor U3810 (N_3810,N_3089,N_2719);
nor U3811 (N_3811,N_3114,N_2697);
and U3812 (N_3812,N_2804,N_3135);
nor U3813 (N_3813,N_2853,N_3046);
xnor U3814 (N_3814,N_2934,N_2642);
nand U3815 (N_3815,N_2448,N_2878);
and U3816 (N_3816,N_2557,N_2567);
nor U3817 (N_3817,N_3072,N_2816);
xnor U3818 (N_3818,N_2571,N_2784);
nor U3819 (N_3819,N_3071,N_2964);
or U3820 (N_3820,N_2798,N_2672);
nor U3821 (N_3821,N_3115,N_2950);
and U3822 (N_3822,N_2657,N_3185);
and U3823 (N_3823,N_2568,N_2820);
nor U3824 (N_3824,N_2846,N_2857);
nor U3825 (N_3825,N_2895,N_2465);
nand U3826 (N_3826,N_2472,N_2934);
nand U3827 (N_3827,N_2502,N_2691);
xnor U3828 (N_3828,N_2717,N_2540);
xnor U3829 (N_3829,N_2825,N_2837);
nor U3830 (N_3830,N_2988,N_2985);
nand U3831 (N_3831,N_2528,N_2940);
nor U3832 (N_3832,N_2754,N_2776);
or U3833 (N_3833,N_2703,N_2701);
xnor U3834 (N_3834,N_2631,N_2786);
nor U3835 (N_3835,N_2915,N_2975);
nor U3836 (N_3836,N_3052,N_2989);
nor U3837 (N_3837,N_2524,N_3183);
or U3838 (N_3838,N_2710,N_2820);
and U3839 (N_3839,N_2720,N_2670);
or U3840 (N_3840,N_2406,N_2912);
nor U3841 (N_3841,N_3165,N_2519);
or U3842 (N_3842,N_3085,N_2650);
nand U3843 (N_3843,N_3044,N_2697);
nor U3844 (N_3844,N_2543,N_2911);
nor U3845 (N_3845,N_2619,N_3154);
nand U3846 (N_3846,N_2469,N_2479);
xnor U3847 (N_3847,N_2979,N_3110);
xnor U3848 (N_3848,N_2551,N_2905);
xor U3849 (N_3849,N_2429,N_2967);
or U3850 (N_3850,N_3020,N_3083);
and U3851 (N_3851,N_2677,N_2438);
xnor U3852 (N_3852,N_3121,N_2506);
nand U3853 (N_3853,N_3169,N_2481);
nand U3854 (N_3854,N_3077,N_2410);
and U3855 (N_3855,N_2613,N_2437);
nor U3856 (N_3856,N_2568,N_2430);
or U3857 (N_3857,N_2836,N_2797);
nor U3858 (N_3858,N_2410,N_2972);
and U3859 (N_3859,N_3116,N_2709);
xnor U3860 (N_3860,N_3023,N_2886);
and U3861 (N_3861,N_2739,N_3076);
and U3862 (N_3862,N_3063,N_3029);
nand U3863 (N_3863,N_2885,N_2558);
nand U3864 (N_3864,N_2657,N_2582);
nor U3865 (N_3865,N_2454,N_2811);
xnor U3866 (N_3866,N_2739,N_3069);
and U3867 (N_3867,N_2572,N_2915);
or U3868 (N_3868,N_3078,N_2430);
nor U3869 (N_3869,N_3074,N_2724);
xnor U3870 (N_3870,N_3190,N_2807);
nand U3871 (N_3871,N_2752,N_2876);
nor U3872 (N_3872,N_3070,N_2858);
and U3873 (N_3873,N_3014,N_2411);
and U3874 (N_3874,N_2507,N_2876);
xnor U3875 (N_3875,N_3001,N_2931);
nor U3876 (N_3876,N_3066,N_3121);
and U3877 (N_3877,N_2539,N_2686);
or U3878 (N_3878,N_3046,N_3135);
or U3879 (N_3879,N_2514,N_2696);
and U3880 (N_3880,N_2786,N_3198);
nand U3881 (N_3881,N_2791,N_2841);
nand U3882 (N_3882,N_2945,N_2935);
nor U3883 (N_3883,N_2770,N_2738);
nand U3884 (N_3884,N_2625,N_2900);
or U3885 (N_3885,N_2833,N_2907);
and U3886 (N_3886,N_2526,N_2782);
or U3887 (N_3887,N_2462,N_2995);
nand U3888 (N_3888,N_2950,N_3194);
nor U3889 (N_3889,N_3040,N_3088);
nor U3890 (N_3890,N_2448,N_3106);
and U3891 (N_3891,N_2779,N_3016);
and U3892 (N_3892,N_2663,N_2809);
and U3893 (N_3893,N_2533,N_2587);
nor U3894 (N_3894,N_2413,N_3172);
nor U3895 (N_3895,N_2817,N_2915);
and U3896 (N_3896,N_2537,N_2419);
xor U3897 (N_3897,N_2590,N_2981);
nor U3898 (N_3898,N_2903,N_2901);
or U3899 (N_3899,N_3035,N_3080);
and U3900 (N_3900,N_3155,N_2420);
nand U3901 (N_3901,N_3096,N_2523);
or U3902 (N_3902,N_2928,N_2913);
and U3903 (N_3903,N_2815,N_2637);
or U3904 (N_3904,N_2463,N_3122);
xor U3905 (N_3905,N_2589,N_3119);
xor U3906 (N_3906,N_2496,N_2556);
and U3907 (N_3907,N_2432,N_2598);
xnor U3908 (N_3908,N_2858,N_2749);
nand U3909 (N_3909,N_3156,N_2620);
nand U3910 (N_3910,N_3182,N_3165);
and U3911 (N_3911,N_3064,N_3123);
nand U3912 (N_3912,N_2738,N_2647);
or U3913 (N_3913,N_2648,N_2610);
and U3914 (N_3914,N_2577,N_2836);
xnor U3915 (N_3915,N_2600,N_2711);
nor U3916 (N_3916,N_3164,N_2412);
xor U3917 (N_3917,N_2615,N_2922);
or U3918 (N_3918,N_3094,N_2991);
xor U3919 (N_3919,N_2972,N_3016);
nor U3920 (N_3920,N_2760,N_3174);
or U3921 (N_3921,N_2846,N_2602);
and U3922 (N_3922,N_3089,N_2480);
or U3923 (N_3923,N_2820,N_2405);
nand U3924 (N_3924,N_2892,N_2503);
and U3925 (N_3925,N_2507,N_2870);
nand U3926 (N_3926,N_2906,N_2449);
and U3927 (N_3927,N_2716,N_3146);
nand U3928 (N_3928,N_2549,N_2928);
or U3929 (N_3929,N_3169,N_2539);
nor U3930 (N_3930,N_3057,N_2713);
nand U3931 (N_3931,N_2757,N_2589);
nand U3932 (N_3932,N_2822,N_3139);
nand U3933 (N_3933,N_2606,N_2668);
and U3934 (N_3934,N_2633,N_2809);
nand U3935 (N_3935,N_2877,N_2780);
xnor U3936 (N_3936,N_2983,N_2663);
nor U3937 (N_3937,N_2712,N_3031);
or U3938 (N_3938,N_3176,N_2789);
and U3939 (N_3939,N_2804,N_2988);
xor U3940 (N_3940,N_2692,N_2855);
nor U3941 (N_3941,N_3177,N_2754);
or U3942 (N_3942,N_3088,N_3109);
nor U3943 (N_3943,N_2411,N_2517);
or U3944 (N_3944,N_2720,N_3020);
and U3945 (N_3945,N_2747,N_2489);
and U3946 (N_3946,N_2728,N_3066);
and U3947 (N_3947,N_2722,N_2975);
nand U3948 (N_3948,N_3158,N_2471);
xnor U3949 (N_3949,N_2720,N_2739);
nand U3950 (N_3950,N_2685,N_2571);
nor U3951 (N_3951,N_2476,N_3016);
nor U3952 (N_3952,N_2479,N_2691);
or U3953 (N_3953,N_3052,N_3045);
and U3954 (N_3954,N_3181,N_2799);
xnor U3955 (N_3955,N_3167,N_2715);
and U3956 (N_3956,N_2963,N_3117);
and U3957 (N_3957,N_2752,N_3185);
or U3958 (N_3958,N_2875,N_2552);
or U3959 (N_3959,N_3003,N_2979);
nor U3960 (N_3960,N_2443,N_3172);
nor U3961 (N_3961,N_2702,N_2942);
and U3962 (N_3962,N_3021,N_3093);
and U3963 (N_3963,N_3159,N_2702);
or U3964 (N_3964,N_2872,N_2663);
and U3965 (N_3965,N_2932,N_2963);
and U3966 (N_3966,N_3040,N_2682);
and U3967 (N_3967,N_2620,N_2695);
xnor U3968 (N_3968,N_2637,N_2837);
xnor U3969 (N_3969,N_3037,N_2572);
and U3970 (N_3970,N_2693,N_2411);
or U3971 (N_3971,N_2618,N_2801);
nand U3972 (N_3972,N_2965,N_3150);
nand U3973 (N_3973,N_3043,N_2543);
xnor U3974 (N_3974,N_2433,N_2622);
nor U3975 (N_3975,N_3097,N_2734);
xnor U3976 (N_3976,N_2778,N_2699);
nand U3977 (N_3977,N_3058,N_2853);
or U3978 (N_3978,N_3089,N_2431);
or U3979 (N_3979,N_3093,N_2428);
and U3980 (N_3980,N_3098,N_2918);
or U3981 (N_3981,N_3101,N_2573);
nor U3982 (N_3982,N_2543,N_2753);
or U3983 (N_3983,N_2444,N_2627);
or U3984 (N_3984,N_2411,N_3135);
and U3985 (N_3985,N_3121,N_3069);
or U3986 (N_3986,N_3161,N_2610);
or U3987 (N_3987,N_2965,N_2709);
xor U3988 (N_3988,N_2590,N_3120);
or U3989 (N_3989,N_2847,N_3087);
or U3990 (N_3990,N_2921,N_2563);
nand U3991 (N_3991,N_3159,N_2856);
and U3992 (N_3992,N_2848,N_2776);
and U3993 (N_3993,N_3141,N_2828);
or U3994 (N_3994,N_2765,N_2934);
or U3995 (N_3995,N_2429,N_2891);
and U3996 (N_3996,N_2768,N_2514);
nand U3997 (N_3997,N_2709,N_3004);
nor U3998 (N_3998,N_3133,N_2964);
nand U3999 (N_3999,N_2812,N_3053);
nand U4000 (N_4000,N_3598,N_3892);
or U4001 (N_4001,N_3629,N_3878);
or U4002 (N_4002,N_3224,N_3500);
and U4003 (N_4003,N_3453,N_3783);
or U4004 (N_4004,N_3718,N_3918);
nand U4005 (N_4005,N_3348,N_3543);
or U4006 (N_4006,N_3904,N_3868);
and U4007 (N_4007,N_3472,N_3391);
or U4008 (N_4008,N_3206,N_3404);
xnor U4009 (N_4009,N_3355,N_3753);
nand U4010 (N_4010,N_3401,N_3493);
xnor U4011 (N_4011,N_3634,N_3287);
xnor U4012 (N_4012,N_3388,N_3200);
xor U4013 (N_4013,N_3235,N_3730);
or U4014 (N_4014,N_3569,N_3648);
or U4015 (N_4015,N_3907,N_3911);
nand U4016 (N_4016,N_3956,N_3310);
nand U4017 (N_4017,N_3673,N_3899);
xnor U4018 (N_4018,N_3835,N_3769);
and U4019 (N_4019,N_3877,N_3656);
xor U4020 (N_4020,N_3549,N_3269);
and U4021 (N_4021,N_3865,N_3901);
and U4022 (N_4022,N_3467,N_3245);
nor U4023 (N_4023,N_3278,N_3624);
nor U4024 (N_4024,N_3759,N_3740);
nand U4025 (N_4025,N_3226,N_3346);
nor U4026 (N_4026,N_3443,N_3921);
nand U4027 (N_4027,N_3218,N_3494);
or U4028 (N_4028,N_3462,N_3264);
nor U4029 (N_4029,N_3266,N_3729);
or U4030 (N_4030,N_3488,N_3447);
nand U4031 (N_4031,N_3779,N_3208);
or U4032 (N_4032,N_3382,N_3283);
xor U4033 (N_4033,N_3708,N_3936);
and U4034 (N_4034,N_3327,N_3812);
nand U4035 (N_4035,N_3314,N_3645);
and U4036 (N_4036,N_3498,N_3703);
and U4037 (N_4037,N_3442,N_3216);
and U4038 (N_4038,N_3585,N_3896);
or U4039 (N_4039,N_3428,N_3933);
nand U4040 (N_4040,N_3396,N_3610);
and U4041 (N_4041,N_3600,N_3836);
nor U4042 (N_4042,N_3309,N_3288);
xnor U4043 (N_4043,N_3803,N_3222);
nor U4044 (N_4044,N_3939,N_3885);
xnor U4045 (N_4045,N_3484,N_3840);
nor U4046 (N_4046,N_3211,N_3652);
and U4047 (N_4047,N_3675,N_3659);
xor U4048 (N_4048,N_3870,N_3797);
xnor U4049 (N_4049,N_3565,N_3203);
and U4050 (N_4050,N_3379,N_3728);
nor U4051 (N_4051,N_3525,N_3412);
nand U4052 (N_4052,N_3946,N_3829);
or U4053 (N_4053,N_3586,N_3672);
xnor U4054 (N_4054,N_3906,N_3699);
and U4055 (N_4055,N_3244,N_3455);
and U4056 (N_4056,N_3377,N_3613);
nand U4057 (N_4057,N_3281,N_3786);
and U4058 (N_4058,N_3332,N_3997);
nand U4059 (N_4059,N_3661,N_3541);
or U4060 (N_4060,N_3646,N_3952);
nand U4061 (N_4061,N_3239,N_3805);
or U4062 (N_4062,N_3810,N_3426);
nand U4063 (N_4063,N_3948,N_3509);
or U4064 (N_4064,N_3260,N_3739);
and U4065 (N_4065,N_3968,N_3290);
or U4066 (N_4066,N_3285,N_3750);
and U4067 (N_4067,N_3882,N_3463);
xor U4068 (N_4068,N_3255,N_3220);
xnor U4069 (N_4069,N_3555,N_3347);
xor U4070 (N_4070,N_3817,N_3249);
nor U4071 (N_4071,N_3717,N_3606);
nand U4072 (N_4072,N_3594,N_3791);
and U4073 (N_4073,N_3573,N_3479);
nand U4074 (N_4074,N_3984,N_3205);
nand U4075 (N_4075,N_3261,N_3507);
and U4076 (N_4076,N_3307,N_3670);
or U4077 (N_4077,N_3660,N_3461);
nor U4078 (N_4078,N_3611,N_3638);
and U4079 (N_4079,N_3774,N_3316);
xnor U4080 (N_4080,N_3427,N_3771);
nand U4081 (N_4081,N_3898,N_3697);
nor U4082 (N_4082,N_3851,N_3380);
nor U4083 (N_4083,N_3857,N_3809);
nand U4084 (N_4084,N_3441,N_3210);
xnor U4085 (N_4085,N_3978,N_3213);
xor U4086 (N_4086,N_3983,N_3518);
nor U4087 (N_4087,N_3470,N_3340);
xor U4088 (N_4088,N_3207,N_3691);
and U4089 (N_4089,N_3924,N_3991);
and U4090 (N_4090,N_3971,N_3482);
and U4091 (N_4091,N_3344,N_3458);
nor U4092 (N_4092,N_3400,N_3834);
nand U4093 (N_4093,N_3905,N_3735);
xnor U4094 (N_4094,N_3209,N_3228);
nor U4095 (N_4095,N_3874,N_3254);
xnor U4096 (N_4096,N_3958,N_3623);
nand U4097 (N_4097,N_3696,N_3929);
nand U4098 (N_4098,N_3231,N_3826);
nand U4099 (N_4099,N_3233,N_3736);
xnor U4100 (N_4100,N_3620,N_3987);
or U4101 (N_4101,N_3553,N_3796);
nand U4102 (N_4102,N_3642,N_3303);
and U4103 (N_4103,N_3478,N_3841);
nor U4104 (N_4104,N_3557,N_3671);
nand U4105 (N_4105,N_3602,N_3650);
nor U4106 (N_4106,N_3782,N_3201);
nand U4107 (N_4107,N_3330,N_3754);
nor U4108 (N_4108,N_3279,N_3732);
or U4109 (N_4109,N_3731,N_3867);
nor U4110 (N_4110,N_3527,N_3848);
nand U4111 (N_4111,N_3842,N_3253);
xor U4112 (N_4112,N_3275,N_3505);
and U4113 (N_4113,N_3849,N_3425);
or U4114 (N_4114,N_3497,N_3241);
nor U4115 (N_4115,N_3859,N_3988);
and U4116 (N_4116,N_3698,N_3420);
nor U4117 (N_4117,N_3430,N_3654);
and U4118 (N_4118,N_3574,N_3516);
xnor U4119 (N_4119,N_3561,N_3940);
nand U4120 (N_4120,N_3433,N_3435);
nor U4121 (N_4121,N_3267,N_3726);
nor U4122 (N_4122,N_3350,N_3223);
nor U4123 (N_4123,N_3402,N_3589);
nand U4124 (N_4124,N_3980,N_3993);
and U4125 (N_4125,N_3491,N_3446);
or U4126 (N_4126,N_3888,N_3571);
xor U4127 (N_4127,N_3334,N_3300);
or U4128 (N_4128,N_3421,N_3657);
or U4129 (N_4129,N_3437,N_3333);
nor U4130 (N_4130,N_3236,N_3282);
or U4131 (N_4131,N_3965,N_3234);
xor U4132 (N_4132,N_3432,N_3838);
nor U4133 (N_4133,N_3941,N_3832);
nand U4134 (N_4134,N_3523,N_3374);
nor U4135 (N_4135,N_3506,N_3329);
xnor U4136 (N_4136,N_3568,N_3331);
and U4137 (N_4137,N_3431,N_3250);
nand U4138 (N_4138,N_3318,N_3601);
xor U4139 (N_4139,N_3534,N_3631);
and U4140 (N_4140,N_3407,N_3361);
nor U4141 (N_4141,N_3913,N_3723);
or U4142 (N_4142,N_3853,N_3296);
nand U4143 (N_4143,N_3595,N_3592);
xor U4144 (N_4144,N_3544,N_3342);
or U4145 (N_4145,N_3639,N_3879);
or U4146 (N_4146,N_3452,N_3238);
nor U4147 (N_4147,N_3385,N_3312);
nand U4148 (N_4148,N_3531,N_3398);
nor U4149 (N_4149,N_3864,N_3454);
nand U4150 (N_4150,N_3489,N_3326);
nor U4151 (N_4151,N_3212,N_3890);
xor U4152 (N_4152,N_3225,N_3576);
nor U4153 (N_4153,N_3360,N_3405);
xnor U4154 (N_4154,N_3604,N_3818);
nand U4155 (N_4155,N_3693,N_3217);
xor U4156 (N_4156,N_3994,N_3837);
nand U4157 (N_4157,N_3880,N_3511);
xor U4158 (N_4158,N_3655,N_3503);
nor U4159 (N_4159,N_3674,N_3724);
xnor U4160 (N_4160,N_3747,N_3647);
nor U4161 (N_4161,N_3635,N_3944);
xnor U4162 (N_4162,N_3756,N_3351);
nor U4163 (N_4163,N_3596,N_3785);
nand U4164 (N_4164,N_3846,N_3664);
or U4165 (N_4165,N_3869,N_3532);
xor U4166 (N_4166,N_3324,N_3284);
nand U4167 (N_4167,N_3977,N_3770);
nor U4168 (N_4168,N_3802,N_3304);
nand U4169 (N_4169,N_3475,N_3335);
nand U4170 (N_4170,N_3358,N_3341);
nand U4171 (N_4171,N_3343,N_3298);
nor U4172 (N_4172,N_3788,N_3550);
and U4173 (N_4173,N_3845,N_3910);
nand U4174 (N_4174,N_3422,N_3483);
or U4175 (N_4175,N_3367,N_3737);
or U4176 (N_4176,N_3519,N_3630);
or U4177 (N_4177,N_3701,N_3925);
nand U4178 (N_4178,N_3273,N_3690);
and U4179 (N_4179,N_3781,N_3821);
nand U4180 (N_4180,N_3584,N_3745);
xor U4181 (N_4181,N_3668,N_3395);
and U4182 (N_4182,N_3808,N_3844);
xor U4183 (N_4183,N_3597,N_3727);
xnor U4184 (N_4184,N_3251,N_3860);
nor U4185 (N_4185,N_3376,N_3247);
or U4186 (N_4186,N_3775,N_3345);
nor U4187 (N_4187,N_3955,N_3378);
nor U4188 (N_4188,N_3976,N_3406);
nand U4189 (N_4189,N_3982,N_3593);
or U4190 (N_4190,N_3354,N_3272);
xnor U4191 (N_4191,N_3567,N_3689);
and U4192 (N_4192,N_3651,N_3530);
or U4193 (N_4193,N_3436,N_3587);
nand U4194 (N_4194,N_3363,N_3469);
and U4195 (N_4195,N_3219,N_3581);
xor U4196 (N_4196,N_3789,N_3556);
nand U4197 (N_4197,N_3619,N_3622);
nand U4198 (N_4198,N_3308,N_3700);
and U4199 (N_4199,N_3237,N_3712);
or U4200 (N_4200,N_3986,N_3321);
and U4201 (N_4201,N_3823,N_3477);
nand U4202 (N_4202,N_3492,N_3383);
nor U4203 (N_4203,N_3716,N_3915);
nand U4204 (N_4204,N_3637,N_3258);
and U4205 (N_4205,N_3336,N_3685);
nand U4206 (N_4206,N_3612,N_3445);
xnor U4207 (N_4207,N_3268,N_3418);
and U4208 (N_4208,N_3502,N_3871);
nand U4209 (N_4209,N_3824,N_3909);
and U4210 (N_4210,N_3669,N_3807);
and U4211 (N_4211,N_3424,N_3636);
or U4212 (N_4212,N_3914,N_3713);
and U4213 (N_4213,N_3787,N_3605);
xnor U4214 (N_4214,N_3353,N_3830);
xor U4215 (N_4215,N_3419,N_3369);
nor U4216 (N_4216,N_3487,N_3917);
and U4217 (N_4217,N_3741,N_3852);
and U4218 (N_4218,N_3572,N_3547);
xnor U4219 (N_4219,N_3257,N_3466);
nand U4220 (N_4220,N_3240,N_3277);
and U4221 (N_4221,N_3804,N_3926);
nor U4222 (N_4222,N_3265,N_3459);
or U4223 (N_4223,N_3937,N_3680);
nor U4224 (N_4224,N_3773,N_3763);
nor U4225 (N_4225,N_3533,N_3570);
or U4226 (N_4226,N_3995,N_3545);
xor U4227 (N_4227,N_3384,N_3625);
and U4228 (N_4228,N_3537,N_3999);
nand U4229 (N_4229,N_3352,N_3504);
nor U4230 (N_4230,N_3473,N_3720);
and U4231 (N_4231,N_3934,N_3644);
nand U4232 (N_4232,N_3524,N_3665);
and U4233 (N_4233,N_3370,N_3816);
or U4234 (N_4234,N_3311,N_3632);
nand U4235 (N_4235,N_3748,N_3411);
and U4236 (N_4236,N_3485,N_3764);
or U4237 (N_4237,N_3695,N_3315);
nor U4238 (N_4238,N_3626,N_3954);
and U4239 (N_4239,N_3481,N_3975);
xnor U4240 (N_4240,N_3559,N_3854);
nor U4241 (N_4241,N_3451,N_3746);
nor U4242 (N_4242,N_3694,N_3951);
or U4243 (N_4243,N_3884,N_3616);
and U4244 (N_4244,N_3349,N_3399);
or U4245 (N_4245,N_3998,N_3919);
and U4246 (N_4246,N_3889,N_3563);
nor U4247 (N_4247,N_3963,N_3725);
nor U4248 (N_4248,N_3683,N_3535);
xor U4249 (N_4249,N_3820,N_3762);
xor U4250 (N_4250,N_3520,N_3947);
and U4251 (N_4251,N_3438,N_3649);
xor U4252 (N_4252,N_3444,N_3409);
nor U4253 (N_4253,N_3881,N_3248);
and U4254 (N_4254,N_3738,N_3633);
xnor U4255 (N_4255,N_3923,N_3614);
or U4256 (N_4256,N_3938,N_3902);
nand U4257 (N_4257,N_3752,N_3552);
and U4258 (N_4258,N_3658,N_3702);
nand U4259 (N_4259,N_3591,N_3768);
nand U4260 (N_4260,N_3960,N_3439);
xnor U4261 (N_4261,N_3897,N_3548);
xor U4262 (N_4262,N_3429,N_3371);
nor U4263 (N_4263,N_3621,N_3386);
nand U4264 (N_4264,N_3767,N_3578);
or U4265 (N_4265,N_3560,N_3289);
and U4266 (N_4266,N_3667,N_3204);
and U4267 (N_4267,N_3449,N_3715);
or U4268 (N_4268,N_3684,N_3526);
xnor U4269 (N_4269,N_3707,N_3811);
nor U4270 (N_4270,N_3930,N_3368);
and U4271 (N_4271,N_3387,N_3843);
and U4272 (N_4272,N_3794,N_3761);
and U4273 (N_4273,N_3323,N_3413);
xnor U4274 (N_4274,N_3790,N_3476);
or U4275 (N_4275,N_3822,N_3608);
and U4276 (N_4276,N_3474,N_3903);
xor U4277 (N_4277,N_3232,N_3299);
xor U4278 (N_4278,N_3357,N_3825);
xor U4279 (N_4279,N_3873,N_3677);
xnor U4280 (N_4280,N_3931,N_3972);
and U4281 (N_4281,N_3508,N_3590);
xnor U4282 (N_4282,N_3302,N_3501);
or U4283 (N_4283,N_3434,N_3397);
nor U4284 (N_4284,N_3850,N_3392);
and U4285 (N_4285,N_3862,N_3522);
xnor U4286 (N_4286,N_3891,N_3389);
nand U4287 (N_4287,N_3468,N_3858);
nand U4288 (N_4288,N_3471,N_3256);
nor U4289 (N_4289,N_3408,N_3227);
nor U4290 (N_4290,N_3229,N_3973);
xnor U4291 (N_4291,N_3364,N_3306);
xor U4292 (N_4292,N_3793,N_3262);
or U4293 (N_4293,N_3706,N_3847);
xnor U4294 (N_4294,N_3799,N_3640);
and U4295 (N_4295,N_3856,N_3618);
nand U4296 (N_4296,N_3861,N_3935);
nand U4297 (N_4297,N_3969,N_3765);
xnor U4298 (N_4298,N_3839,N_3800);
and U4299 (N_4299,N_3678,N_3757);
and U4300 (N_4300,N_3221,N_3554);
or U4301 (N_4301,N_3628,N_3989);
and U4302 (N_4302,N_3528,N_3366);
nor U4303 (N_4303,N_3577,N_3362);
or U4304 (N_4304,N_3760,N_3957);
xnor U4305 (N_4305,N_3710,N_3744);
xor U4306 (N_4306,N_3666,N_3813);
nand U4307 (N_4307,N_3751,N_3393);
or U4308 (N_4308,N_3415,N_3719);
or U4309 (N_4309,N_3546,N_3894);
nand U4310 (N_4310,N_3876,N_3863);
nor U4311 (N_4311,N_3961,N_3943);
xnor U4312 (N_4312,N_3778,N_3450);
and U4313 (N_4313,N_3676,N_3339);
or U4314 (N_4314,N_3722,N_3679);
nor U4315 (N_4315,N_3259,N_3833);
xor U4316 (N_4316,N_3920,N_3819);
nand U4317 (N_4317,N_3682,N_3280);
xor U4318 (N_4318,N_3692,N_3681);
xnor U4319 (N_4319,N_3539,N_3579);
or U4320 (N_4320,N_3990,N_3337);
and U4321 (N_4321,N_3580,N_3495);
nand U4322 (N_4322,N_3582,N_3270);
nor U4323 (N_4323,N_3291,N_3743);
or U4324 (N_4324,N_3996,N_3855);
nand U4325 (N_4325,N_3286,N_3514);
nand U4326 (N_4326,N_3798,N_3932);
nor U4327 (N_4327,N_3607,N_3414);
and U4328 (N_4328,N_3643,N_3801);
or U4329 (N_4329,N_3942,N_3513);
nor U4330 (N_4330,N_3962,N_3301);
nand U4331 (N_4331,N_3480,N_3295);
nand U4332 (N_4332,N_3928,N_3417);
or U4333 (N_4333,N_3887,N_3230);
and U4334 (N_4334,N_3714,N_3320);
nand U4335 (N_4335,N_3653,N_3866);
xnor U4336 (N_4336,N_3900,N_3815);
xnor U4337 (N_4337,N_3246,N_3912);
xnor U4338 (N_4338,N_3365,N_3536);
nor U4339 (N_4339,N_3448,N_3294);
nor U4340 (N_4340,N_3922,N_3373);
and U4341 (N_4341,N_3381,N_3734);
xnor U4342 (N_4342,N_3992,N_3515);
nand U4343 (N_4343,N_3202,N_3772);
nor U4344 (N_4344,N_3529,N_3964);
and U4345 (N_4345,N_3416,N_3875);
xor U4346 (N_4346,N_3603,N_3372);
or U4347 (N_4347,N_3540,N_3953);
nand U4348 (N_4348,N_3886,N_3486);
nand U4349 (N_4349,N_3828,N_3403);
xnor U4350 (N_4350,N_3641,N_3686);
or U4351 (N_4351,N_3627,N_3517);
nor U4352 (N_4352,N_3512,N_3872);
or U4353 (N_4353,N_3711,N_3893);
nor U4354 (N_4354,N_3465,N_3945);
nor U4355 (N_4355,N_3338,N_3319);
and U4356 (N_4356,N_3317,N_3687);
or U4357 (N_4357,N_3766,N_3985);
nand U4358 (N_4358,N_3243,N_3276);
or U4359 (N_4359,N_3776,N_3795);
and U4360 (N_4360,N_3709,N_3831);
or U4361 (N_4361,N_3575,N_3908);
nand U4362 (N_4362,N_3981,N_3966);
xnor U4363 (N_4363,N_3558,N_3305);
nor U4364 (N_4364,N_3521,N_3827);
nand U4365 (N_4365,N_3293,N_3499);
and U4366 (N_4366,N_3423,N_3883);
nand U4367 (N_4367,N_3440,N_3792);
or U4368 (N_4368,N_3313,N_3967);
nor U4369 (N_4369,N_3615,N_3274);
nand U4370 (N_4370,N_3704,N_3375);
and U4371 (N_4371,N_3895,N_3457);
nor U4372 (N_4372,N_3970,N_3721);
xor U4373 (N_4373,N_3542,N_3297);
xnor U4374 (N_4374,N_3214,N_3599);
and U4375 (N_4375,N_3325,N_3328);
nand U4376 (N_4376,N_3758,N_3749);
nand U4377 (N_4377,N_3617,N_3410);
and U4378 (N_4378,N_3814,N_3662);
and U4379 (N_4379,N_3464,N_3263);
nor U4380 (N_4380,N_3974,N_3490);
and U4381 (N_4381,N_3755,N_3609);
or U4382 (N_4382,N_3359,N_3949);
and U4383 (N_4383,N_3496,N_3394);
nand U4384 (N_4384,N_3742,N_3927);
nor U4385 (N_4385,N_3784,N_3916);
xnor U4386 (N_4386,N_3733,N_3959);
nor U4387 (N_4387,N_3356,N_3322);
nor U4388 (N_4388,N_3252,N_3583);
xnor U4389 (N_4389,N_3777,N_3460);
or U4390 (N_4390,N_3271,N_3551);
and U4391 (N_4391,N_3215,N_3688);
or U4392 (N_4392,N_3242,N_3705);
nor U4393 (N_4393,N_3562,N_3780);
nand U4394 (N_4394,N_3390,N_3564);
and U4395 (N_4395,N_3806,N_3663);
nand U4396 (N_4396,N_3566,N_3292);
and U4397 (N_4397,N_3979,N_3510);
xor U4398 (N_4398,N_3456,N_3950);
nor U4399 (N_4399,N_3538,N_3588);
nand U4400 (N_4400,N_3723,N_3950);
or U4401 (N_4401,N_3802,N_3544);
xnor U4402 (N_4402,N_3445,N_3239);
or U4403 (N_4403,N_3752,N_3541);
and U4404 (N_4404,N_3215,N_3865);
or U4405 (N_4405,N_3216,N_3555);
xor U4406 (N_4406,N_3811,N_3350);
xor U4407 (N_4407,N_3273,N_3474);
and U4408 (N_4408,N_3366,N_3301);
nor U4409 (N_4409,N_3905,N_3344);
nand U4410 (N_4410,N_3433,N_3731);
and U4411 (N_4411,N_3829,N_3907);
xnor U4412 (N_4412,N_3444,N_3220);
and U4413 (N_4413,N_3637,N_3278);
and U4414 (N_4414,N_3872,N_3472);
xor U4415 (N_4415,N_3379,N_3525);
nand U4416 (N_4416,N_3852,N_3826);
nor U4417 (N_4417,N_3694,N_3308);
nor U4418 (N_4418,N_3714,N_3416);
or U4419 (N_4419,N_3809,N_3468);
xnor U4420 (N_4420,N_3826,N_3956);
and U4421 (N_4421,N_3347,N_3930);
and U4422 (N_4422,N_3651,N_3611);
nor U4423 (N_4423,N_3628,N_3544);
or U4424 (N_4424,N_3571,N_3599);
or U4425 (N_4425,N_3913,N_3272);
nand U4426 (N_4426,N_3998,N_3553);
or U4427 (N_4427,N_3816,N_3237);
and U4428 (N_4428,N_3281,N_3439);
or U4429 (N_4429,N_3418,N_3243);
xnor U4430 (N_4430,N_3721,N_3899);
nor U4431 (N_4431,N_3553,N_3659);
or U4432 (N_4432,N_3213,N_3572);
nor U4433 (N_4433,N_3661,N_3696);
xnor U4434 (N_4434,N_3446,N_3790);
xnor U4435 (N_4435,N_3627,N_3316);
nor U4436 (N_4436,N_3424,N_3900);
nor U4437 (N_4437,N_3884,N_3792);
and U4438 (N_4438,N_3434,N_3926);
and U4439 (N_4439,N_3874,N_3238);
nand U4440 (N_4440,N_3467,N_3435);
and U4441 (N_4441,N_3901,N_3507);
xor U4442 (N_4442,N_3341,N_3784);
nor U4443 (N_4443,N_3804,N_3848);
nor U4444 (N_4444,N_3816,N_3843);
nand U4445 (N_4445,N_3234,N_3222);
xnor U4446 (N_4446,N_3559,N_3978);
nor U4447 (N_4447,N_3600,N_3894);
or U4448 (N_4448,N_3664,N_3271);
nand U4449 (N_4449,N_3820,N_3886);
nand U4450 (N_4450,N_3499,N_3614);
nand U4451 (N_4451,N_3279,N_3385);
xnor U4452 (N_4452,N_3716,N_3438);
xnor U4453 (N_4453,N_3682,N_3790);
nand U4454 (N_4454,N_3513,N_3541);
or U4455 (N_4455,N_3469,N_3707);
xnor U4456 (N_4456,N_3540,N_3798);
or U4457 (N_4457,N_3349,N_3337);
nand U4458 (N_4458,N_3288,N_3582);
xor U4459 (N_4459,N_3402,N_3600);
or U4460 (N_4460,N_3370,N_3788);
or U4461 (N_4461,N_3499,N_3237);
xnor U4462 (N_4462,N_3376,N_3331);
nor U4463 (N_4463,N_3318,N_3787);
xor U4464 (N_4464,N_3267,N_3724);
xnor U4465 (N_4465,N_3622,N_3661);
and U4466 (N_4466,N_3317,N_3757);
and U4467 (N_4467,N_3221,N_3894);
nand U4468 (N_4468,N_3325,N_3575);
or U4469 (N_4469,N_3801,N_3957);
xnor U4470 (N_4470,N_3989,N_3531);
nor U4471 (N_4471,N_3371,N_3670);
xnor U4472 (N_4472,N_3556,N_3902);
nor U4473 (N_4473,N_3767,N_3958);
nor U4474 (N_4474,N_3668,N_3570);
and U4475 (N_4475,N_3497,N_3371);
xnor U4476 (N_4476,N_3262,N_3721);
nand U4477 (N_4477,N_3665,N_3477);
nor U4478 (N_4478,N_3290,N_3512);
and U4479 (N_4479,N_3737,N_3229);
nand U4480 (N_4480,N_3933,N_3330);
and U4481 (N_4481,N_3772,N_3952);
nand U4482 (N_4482,N_3303,N_3217);
xnor U4483 (N_4483,N_3901,N_3270);
nand U4484 (N_4484,N_3650,N_3865);
or U4485 (N_4485,N_3940,N_3440);
nor U4486 (N_4486,N_3442,N_3892);
or U4487 (N_4487,N_3598,N_3380);
and U4488 (N_4488,N_3726,N_3486);
and U4489 (N_4489,N_3645,N_3785);
and U4490 (N_4490,N_3230,N_3724);
nand U4491 (N_4491,N_3711,N_3415);
and U4492 (N_4492,N_3716,N_3211);
and U4493 (N_4493,N_3763,N_3921);
xnor U4494 (N_4494,N_3653,N_3294);
or U4495 (N_4495,N_3206,N_3567);
xor U4496 (N_4496,N_3856,N_3491);
xor U4497 (N_4497,N_3342,N_3454);
or U4498 (N_4498,N_3751,N_3712);
nand U4499 (N_4499,N_3659,N_3373);
and U4500 (N_4500,N_3546,N_3268);
or U4501 (N_4501,N_3344,N_3716);
and U4502 (N_4502,N_3237,N_3369);
nor U4503 (N_4503,N_3757,N_3823);
nand U4504 (N_4504,N_3652,N_3376);
xor U4505 (N_4505,N_3322,N_3401);
or U4506 (N_4506,N_3550,N_3580);
nor U4507 (N_4507,N_3985,N_3630);
and U4508 (N_4508,N_3417,N_3482);
or U4509 (N_4509,N_3353,N_3241);
nor U4510 (N_4510,N_3660,N_3705);
and U4511 (N_4511,N_3603,N_3965);
nor U4512 (N_4512,N_3742,N_3325);
or U4513 (N_4513,N_3784,N_3922);
nand U4514 (N_4514,N_3505,N_3582);
xnor U4515 (N_4515,N_3780,N_3393);
nor U4516 (N_4516,N_3249,N_3881);
xnor U4517 (N_4517,N_3814,N_3569);
or U4518 (N_4518,N_3757,N_3987);
nand U4519 (N_4519,N_3742,N_3836);
and U4520 (N_4520,N_3843,N_3666);
nor U4521 (N_4521,N_3657,N_3368);
nor U4522 (N_4522,N_3653,N_3340);
and U4523 (N_4523,N_3737,N_3974);
xnor U4524 (N_4524,N_3818,N_3380);
nor U4525 (N_4525,N_3855,N_3488);
nor U4526 (N_4526,N_3610,N_3448);
nor U4527 (N_4527,N_3303,N_3379);
and U4528 (N_4528,N_3826,N_3547);
and U4529 (N_4529,N_3602,N_3801);
xnor U4530 (N_4530,N_3489,N_3474);
xnor U4531 (N_4531,N_3759,N_3308);
nand U4532 (N_4532,N_3603,N_3797);
nand U4533 (N_4533,N_3456,N_3260);
and U4534 (N_4534,N_3286,N_3328);
and U4535 (N_4535,N_3842,N_3494);
nor U4536 (N_4536,N_3674,N_3277);
nand U4537 (N_4537,N_3445,N_3522);
xnor U4538 (N_4538,N_3919,N_3403);
nor U4539 (N_4539,N_3352,N_3849);
nor U4540 (N_4540,N_3587,N_3254);
nor U4541 (N_4541,N_3671,N_3955);
xor U4542 (N_4542,N_3314,N_3584);
nor U4543 (N_4543,N_3395,N_3906);
and U4544 (N_4544,N_3698,N_3968);
xor U4545 (N_4545,N_3649,N_3651);
xor U4546 (N_4546,N_3436,N_3367);
or U4547 (N_4547,N_3626,N_3403);
nand U4548 (N_4548,N_3839,N_3548);
or U4549 (N_4549,N_3275,N_3202);
or U4550 (N_4550,N_3276,N_3735);
and U4551 (N_4551,N_3532,N_3494);
nand U4552 (N_4552,N_3203,N_3596);
and U4553 (N_4553,N_3270,N_3422);
and U4554 (N_4554,N_3610,N_3788);
nand U4555 (N_4555,N_3571,N_3757);
nor U4556 (N_4556,N_3353,N_3683);
xnor U4557 (N_4557,N_3574,N_3906);
nor U4558 (N_4558,N_3528,N_3433);
and U4559 (N_4559,N_3350,N_3902);
nand U4560 (N_4560,N_3944,N_3215);
and U4561 (N_4561,N_3255,N_3634);
and U4562 (N_4562,N_3675,N_3448);
xnor U4563 (N_4563,N_3783,N_3218);
nand U4564 (N_4564,N_3774,N_3972);
xnor U4565 (N_4565,N_3394,N_3907);
nor U4566 (N_4566,N_3605,N_3517);
nor U4567 (N_4567,N_3981,N_3399);
xnor U4568 (N_4568,N_3730,N_3370);
or U4569 (N_4569,N_3981,N_3358);
nor U4570 (N_4570,N_3285,N_3232);
or U4571 (N_4571,N_3250,N_3913);
or U4572 (N_4572,N_3435,N_3627);
nand U4573 (N_4573,N_3467,N_3294);
or U4574 (N_4574,N_3581,N_3621);
nor U4575 (N_4575,N_3612,N_3355);
xnor U4576 (N_4576,N_3353,N_3651);
nand U4577 (N_4577,N_3743,N_3689);
or U4578 (N_4578,N_3741,N_3544);
and U4579 (N_4579,N_3884,N_3902);
nor U4580 (N_4580,N_3238,N_3296);
nand U4581 (N_4581,N_3863,N_3540);
or U4582 (N_4582,N_3293,N_3243);
xnor U4583 (N_4583,N_3228,N_3721);
or U4584 (N_4584,N_3944,N_3876);
nor U4585 (N_4585,N_3769,N_3795);
and U4586 (N_4586,N_3956,N_3940);
nor U4587 (N_4587,N_3962,N_3828);
and U4588 (N_4588,N_3498,N_3841);
or U4589 (N_4589,N_3518,N_3697);
or U4590 (N_4590,N_3213,N_3762);
or U4591 (N_4591,N_3256,N_3227);
nand U4592 (N_4592,N_3896,N_3301);
nand U4593 (N_4593,N_3208,N_3333);
or U4594 (N_4594,N_3677,N_3270);
or U4595 (N_4595,N_3787,N_3861);
nand U4596 (N_4596,N_3731,N_3630);
or U4597 (N_4597,N_3653,N_3588);
nor U4598 (N_4598,N_3304,N_3497);
and U4599 (N_4599,N_3537,N_3549);
xnor U4600 (N_4600,N_3630,N_3520);
nand U4601 (N_4601,N_3762,N_3355);
xnor U4602 (N_4602,N_3815,N_3694);
nand U4603 (N_4603,N_3876,N_3593);
or U4604 (N_4604,N_3989,N_3610);
xor U4605 (N_4605,N_3540,N_3895);
nor U4606 (N_4606,N_3990,N_3836);
nand U4607 (N_4607,N_3603,N_3486);
xnor U4608 (N_4608,N_3915,N_3753);
nor U4609 (N_4609,N_3629,N_3513);
nor U4610 (N_4610,N_3746,N_3907);
nor U4611 (N_4611,N_3671,N_3580);
nand U4612 (N_4612,N_3485,N_3688);
nand U4613 (N_4613,N_3424,N_3627);
or U4614 (N_4614,N_3683,N_3367);
xnor U4615 (N_4615,N_3654,N_3807);
xnor U4616 (N_4616,N_3224,N_3576);
nor U4617 (N_4617,N_3699,N_3896);
xor U4618 (N_4618,N_3896,N_3496);
and U4619 (N_4619,N_3472,N_3229);
or U4620 (N_4620,N_3212,N_3878);
xor U4621 (N_4621,N_3613,N_3553);
nand U4622 (N_4622,N_3497,N_3205);
xor U4623 (N_4623,N_3540,N_3968);
or U4624 (N_4624,N_3686,N_3542);
and U4625 (N_4625,N_3435,N_3967);
xor U4626 (N_4626,N_3499,N_3813);
or U4627 (N_4627,N_3847,N_3591);
or U4628 (N_4628,N_3537,N_3894);
nor U4629 (N_4629,N_3927,N_3632);
xor U4630 (N_4630,N_3465,N_3685);
nand U4631 (N_4631,N_3541,N_3780);
nand U4632 (N_4632,N_3512,N_3221);
and U4633 (N_4633,N_3565,N_3592);
or U4634 (N_4634,N_3888,N_3635);
or U4635 (N_4635,N_3366,N_3534);
nand U4636 (N_4636,N_3352,N_3728);
nand U4637 (N_4637,N_3609,N_3713);
xor U4638 (N_4638,N_3737,N_3912);
xor U4639 (N_4639,N_3577,N_3863);
and U4640 (N_4640,N_3947,N_3478);
nand U4641 (N_4641,N_3594,N_3785);
nand U4642 (N_4642,N_3772,N_3573);
and U4643 (N_4643,N_3621,N_3920);
nand U4644 (N_4644,N_3756,N_3759);
nor U4645 (N_4645,N_3651,N_3939);
nor U4646 (N_4646,N_3753,N_3869);
nand U4647 (N_4647,N_3805,N_3474);
and U4648 (N_4648,N_3605,N_3727);
or U4649 (N_4649,N_3828,N_3252);
or U4650 (N_4650,N_3927,N_3714);
and U4651 (N_4651,N_3711,N_3890);
and U4652 (N_4652,N_3307,N_3569);
and U4653 (N_4653,N_3927,N_3738);
nor U4654 (N_4654,N_3982,N_3908);
and U4655 (N_4655,N_3969,N_3665);
xnor U4656 (N_4656,N_3464,N_3302);
nor U4657 (N_4657,N_3893,N_3295);
nand U4658 (N_4658,N_3204,N_3237);
xnor U4659 (N_4659,N_3445,N_3791);
and U4660 (N_4660,N_3424,N_3529);
nor U4661 (N_4661,N_3362,N_3416);
nand U4662 (N_4662,N_3893,N_3989);
xor U4663 (N_4663,N_3236,N_3540);
xnor U4664 (N_4664,N_3395,N_3456);
xor U4665 (N_4665,N_3750,N_3444);
xor U4666 (N_4666,N_3518,N_3595);
xor U4667 (N_4667,N_3435,N_3602);
and U4668 (N_4668,N_3877,N_3864);
nor U4669 (N_4669,N_3732,N_3848);
nand U4670 (N_4670,N_3555,N_3731);
or U4671 (N_4671,N_3400,N_3904);
nand U4672 (N_4672,N_3780,N_3392);
nor U4673 (N_4673,N_3844,N_3717);
nand U4674 (N_4674,N_3782,N_3908);
nand U4675 (N_4675,N_3571,N_3778);
or U4676 (N_4676,N_3959,N_3641);
xnor U4677 (N_4677,N_3241,N_3206);
nor U4678 (N_4678,N_3328,N_3993);
nor U4679 (N_4679,N_3843,N_3565);
and U4680 (N_4680,N_3983,N_3625);
and U4681 (N_4681,N_3955,N_3516);
and U4682 (N_4682,N_3540,N_3707);
nor U4683 (N_4683,N_3616,N_3443);
nor U4684 (N_4684,N_3438,N_3858);
nand U4685 (N_4685,N_3740,N_3948);
nand U4686 (N_4686,N_3680,N_3913);
nand U4687 (N_4687,N_3289,N_3373);
or U4688 (N_4688,N_3291,N_3628);
nor U4689 (N_4689,N_3629,N_3343);
xnor U4690 (N_4690,N_3826,N_3981);
nand U4691 (N_4691,N_3359,N_3478);
nor U4692 (N_4692,N_3240,N_3799);
and U4693 (N_4693,N_3929,N_3269);
xor U4694 (N_4694,N_3258,N_3809);
nand U4695 (N_4695,N_3652,N_3241);
xor U4696 (N_4696,N_3597,N_3736);
nor U4697 (N_4697,N_3285,N_3836);
nor U4698 (N_4698,N_3835,N_3999);
nand U4699 (N_4699,N_3675,N_3900);
and U4700 (N_4700,N_3755,N_3822);
nor U4701 (N_4701,N_3781,N_3696);
and U4702 (N_4702,N_3732,N_3795);
xnor U4703 (N_4703,N_3231,N_3330);
and U4704 (N_4704,N_3692,N_3262);
and U4705 (N_4705,N_3556,N_3623);
xnor U4706 (N_4706,N_3772,N_3700);
xnor U4707 (N_4707,N_3268,N_3344);
and U4708 (N_4708,N_3363,N_3890);
nand U4709 (N_4709,N_3965,N_3787);
nand U4710 (N_4710,N_3961,N_3431);
and U4711 (N_4711,N_3814,N_3970);
and U4712 (N_4712,N_3535,N_3309);
or U4713 (N_4713,N_3260,N_3273);
nor U4714 (N_4714,N_3719,N_3671);
nand U4715 (N_4715,N_3213,N_3731);
or U4716 (N_4716,N_3644,N_3576);
nor U4717 (N_4717,N_3612,N_3805);
nor U4718 (N_4718,N_3320,N_3876);
nand U4719 (N_4719,N_3494,N_3212);
and U4720 (N_4720,N_3402,N_3927);
nand U4721 (N_4721,N_3688,N_3779);
or U4722 (N_4722,N_3731,N_3302);
nand U4723 (N_4723,N_3438,N_3409);
xor U4724 (N_4724,N_3470,N_3514);
or U4725 (N_4725,N_3498,N_3397);
and U4726 (N_4726,N_3434,N_3877);
nand U4727 (N_4727,N_3514,N_3768);
and U4728 (N_4728,N_3245,N_3933);
or U4729 (N_4729,N_3628,N_3766);
or U4730 (N_4730,N_3352,N_3917);
xor U4731 (N_4731,N_3705,N_3425);
nand U4732 (N_4732,N_3676,N_3774);
xnor U4733 (N_4733,N_3668,N_3871);
or U4734 (N_4734,N_3974,N_3237);
or U4735 (N_4735,N_3686,N_3447);
and U4736 (N_4736,N_3436,N_3921);
nor U4737 (N_4737,N_3516,N_3534);
nor U4738 (N_4738,N_3880,N_3731);
nand U4739 (N_4739,N_3469,N_3865);
xnor U4740 (N_4740,N_3932,N_3806);
and U4741 (N_4741,N_3307,N_3896);
xor U4742 (N_4742,N_3314,N_3909);
and U4743 (N_4743,N_3458,N_3956);
or U4744 (N_4744,N_3958,N_3305);
or U4745 (N_4745,N_3725,N_3276);
and U4746 (N_4746,N_3884,N_3448);
or U4747 (N_4747,N_3311,N_3573);
nor U4748 (N_4748,N_3700,N_3967);
or U4749 (N_4749,N_3203,N_3945);
nor U4750 (N_4750,N_3386,N_3660);
and U4751 (N_4751,N_3215,N_3335);
or U4752 (N_4752,N_3497,N_3646);
xor U4753 (N_4753,N_3225,N_3911);
nand U4754 (N_4754,N_3585,N_3562);
nand U4755 (N_4755,N_3752,N_3445);
nor U4756 (N_4756,N_3526,N_3802);
or U4757 (N_4757,N_3238,N_3755);
and U4758 (N_4758,N_3372,N_3321);
or U4759 (N_4759,N_3372,N_3229);
nand U4760 (N_4760,N_3776,N_3665);
and U4761 (N_4761,N_3825,N_3946);
nand U4762 (N_4762,N_3705,N_3789);
xnor U4763 (N_4763,N_3867,N_3970);
and U4764 (N_4764,N_3995,N_3564);
and U4765 (N_4765,N_3685,N_3456);
or U4766 (N_4766,N_3296,N_3900);
nand U4767 (N_4767,N_3990,N_3927);
and U4768 (N_4768,N_3683,N_3524);
and U4769 (N_4769,N_3490,N_3696);
or U4770 (N_4770,N_3730,N_3361);
xor U4771 (N_4771,N_3874,N_3601);
and U4772 (N_4772,N_3354,N_3244);
and U4773 (N_4773,N_3920,N_3933);
nand U4774 (N_4774,N_3209,N_3757);
nand U4775 (N_4775,N_3879,N_3334);
nand U4776 (N_4776,N_3320,N_3763);
or U4777 (N_4777,N_3991,N_3600);
xor U4778 (N_4778,N_3493,N_3251);
and U4779 (N_4779,N_3277,N_3697);
and U4780 (N_4780,N_3839,N_3643);
or U4781 (N_4781,N_3502,N_3717);
xor U4782 (N_4782,N_3862,N_3289);
and U4783 (N_4783,N_3490,N_3869);
nor U4784 (N_4784,N_3880,N_3641);
xor U4785 (N_4785,N_3997,N_3869);
or U4786 (N_4786,N_3506,N_3945);
xor U4787 (N_4787,N_3365,N_3430);
or U4788 (N_4788,N_3957,N_3718);
nand U4789 (N_4789,N_3236,N_3332);
nand U4790 (N_4790,N_3411,N_3807);
xnor U4791 (N_4791,N_3733,N_3813);
nor U4792 (N_4792,N_3845,N_3767);
nor U4793 (N_4793,N_3626,N_3842);
nor U4794 (N_4794,N_3275,N_3576);
and U4795 (N_4795,N_3291,N_3622);
xnor U4796 (N_4796,N_3535,N_3435);
nor U4797 (N_4797,N_3603,N_3985);
xor U4798 (N_4798,N_3915,N_3373);
xnor U4799 (N_4799,N_3495,N_3761);
and U4800 (N_4800,N_4646,N_4288);
nor U4801 (N_4801,N_4115,N_4536);
nand U4802 (N_4802,N_4648,N_4465);
nor U4803 (N_4803,N_4377,N_4329);
nand U4804 (N_4804,N_4152,N_4642);
or U4805 (N_4805,N_4511,N_4728);
xnor U4806 (N_4806,N_4497,N_4272);
nor U4807 (N_4807,N_4373,N_4610);
and U4808 (N_4808,N_4585,N_4296);
nand U4809 (N_4809,N_4142,N_4518);
or U4810 (N_4810,N_4643,N_4565);
nor U4811 (N_4811,N_4561,N_4470);
or U4812 (N_4812,N_4572,N_4651);
nor U4813 (N_4813,N_4127,N_4614);
nand U4814 (N_4814,N_4611,N_4169);
and U4815 (N_4815,N_4394,N_4302);
nand U4816 (N_4816,N_4184,N_4521);
or U4817 (N_4817,N_4589,N_4051);
xor U4818 (N_4818,N_4056,N_4334);
nand U4819 (N_4819,N_4254,N_4710);
nor U4820 (N_4820,N_4206,N_4111);
or U4821 (N_4821,N_4683,N_4258);
nor U4822 (N_4822,N_4598,N_4059);
nand U4823 (N_4823,N_4792,N_4780);
or U4824 (N_4824,N_4649,N_4125);
nand U4825 (N_4825,N_4149,N_4139);
xnor U4826 (N_4826,N_4242,N_4338);
nor U4827 (N_4827,N_4742,N_4011);
nor U4828 (N_4828,N_4312,N_4336);
or U4829 (N_4829,N_4375,N_4692);
xor U4830 (N_4830,N_4550,N_4037);
nand U4831 (N_4831,N_4596,N_4501);
nor U4832 (N_4832,N_4458,N_4775);
nand U4833 (N_4833,N_4279,N_4695);
xnor U4834 (N_4834,N_4349,N_4238);
xor U4835 (N_4835,N_4739,N_4007);
nor U4836 (N_4836,N_4182,N_4694);
and U4837 (N_4837,N_4021,N_4447);
and U4838 (N_4838,N_4240,N_4116);
and U4839 (N_4839,N_4018,N_4028);
xnor U4840 (N_4840,N_4108,N_4453);
xor U4841 (N_4841,N_4367,N_4268);
or U4842 (N_4842,N_4395,N_4460);
nor U4843 (N_4843,N_4569,N_4584);
nand U4844 (N_4844,N_4330,N_4389);
and U4845 (N_4845,N_4563,N_4210);
and U4846 (N_4846,N_4661,N_4492);
nand U4847 (N_4847,N_4793,N_4622);
and U4848 (N_4848,N_4160,N_4174);
xor U4849 (N_4849,N_4426,N_4445);
and U4850 (N_4850,N_4045,N_4117);
or U4851 (N_4851,N_4345,N_4118);
and U4852 (N_4852,N_4163,N_4135);
xnor U4853 (N_4853,N_4653,N_4269);
and U4854 (N_4854,N_4637,N_4402);
nand U4855 (N_4855,N_4164,N_4382);
or U4856 (N_4856,N_4574,N_4079);
and U4857 (N_4857,N_4295,N_4278);
nand U4858 (N_4858,N_4093,N_4043);
xor U4859 (N_4859,N_4244,N_4541);
nor U4860 (N_4860,N_4300,N_4299);
xor U4861 (N_4861,N_4487,N_4428);
and U4862 (N_4862,N_4157,N_4309);
or U4863 (N_4863,N_4446,N_4600);
nor U4864 (N_4864,N_4361,N_4180);
and U4865 (N_4865,N_4176,N_4228);
and U4866 (N_4866,N_4359,N_4229);
or U4867 (N_4867,N_4190,N_4746);
and U4868 (N_4868,N_4619,N_4062);
nand U4869 (N_4869,N_4727,N_4623);
nand U4870 (N_4870,N_4721,N_4378);
xor U4871 (N_4871,N_4151,N_4401);
or U4872 (N_4872,N_4613,N_4686);
nor U4873 (N_4873,N_4509,N_4650);
nor U4874 (N_4874,N_4355,N_4666);
nand U4875 (N_4875,N_4488,N_4433);
xor U4876 (N_4876,N_4621,N_4473);
or U4877 (N_4877,N_4540,N_4348);
nor U4878 (N_4878,N_4413,N_4523);
nand U4879 (N_4879,N_4143,N_4124);
nand U4880 (N_4880,N_4734,N_4101);
nand U4881 (N_4881,N_4570,N_4554);
nor U4882 (N_4882,N_4194,N_4150);
xor U4883 (N_4883,N_4067,N_4567);
nor U4884 (N_4884,N_4073,N_4145);
xnor U4885 (N_4885,N_4726,N_4631);
nand U4886 (N_4886,N_4220,N_4679);
and U4887 (N_4887,N_4015,N_4027);
nand U4888 (N_4888,N_4105,N_4070);
and U4889 (N_4889,N_4205,N_4645);
nand U4890 (N_4890,N_4740,N_4230);
and U4891 (N_4891,N_4404,N_4717);
nor U4892 (N_4892,N_4581,N_4400);
and U4893 (N_4893,N_4071,N_4577);
nor U4894 (N_4894,N_4232,N_4781);
nor U4895 (N_4895,N_4219,N_4779);
and U4896 (N_4896,N_4467,N_4195);
nor U4897 (N_4897,N_4094,N_4575);
or U4898 (N_4898,N_4434,N_4385);
and U4899 (N_4899,N_4544,N_4328);
xor U4900 (N_4900,N_4767,N_4215);
nand U4901 (N_4901,N_4159,N_4669);
nand U4902 (N_4902,N_4436,N_4390);
xor U4903 (N_4903,N_4632,N_4791);
nand U4904 (N_4904,N_4351,N_4306);
or U4905 (N_4905,N_4353,N_4660);
nand U4906 (N_4906,N_4211,N_4256);
xnor U4907 (N_4907,N_4044,N_4667);
or U4908 (N_4908,N_4136,N_4588);
and U4909 (N_4909,N_4038,N_4741);
nand U4910 (N_4910,N_4250,N_4415);
nand U4911 (N_4911,N_4578,N_4462);
nor U4912 (N_4912,N_4644,N_4054);
or U4913 (N_4913,N_4264,N_4366);
and U4914 (N_4914,N_4247,N_4448);
xor U4915 (N_4915,N_4370,N_4451);
or U4916 (N_4916,N_4292,N_4301);
nor U4917 (N_4917,N_4612,N_4416);
and U4918 (N_4918,N_4281,N_4409);
xnor U4919 (N_4919,N_4693,N_4347);
xor U4920 (N_4920,N_4699,N_4773);
and U4921 (N_4921,N_4714,N_4325);
or U4922 (N_4922,N_4641,N_4736);
nor U4923 (N_4923,N_4607,N_4315);
nor U4924 (N_4924,N_4560,N_4091);
nor U4925 (N_4925,N_4333,N_4130);
and U4926 (N_4926,N_4757,N_4481);
or U4927 (N_4927,N_4539,N_4123);
nand U4928 (N_4928,N_4738,N_4128);
and U4929 (N_4929,N_4399,N_4609);
or U4930 (N_4930,N_4750,N_4769);
nor U4931 (N_4931,N_4562,N_4034);
xor U4932 (N_4932,N_4223,N_4617);
nand U4933 (N_4933,N_4058,N_4285);
nand U4934 (N_4934,N_4510,N_4469);
or U4935 (N_4935,N_4237,N_4483);
nand U4936 (N_4936,N_4566,N_4291);
nor U4937 (N_4937,N_4280,N_4690);
nor U4938 (N_4938,N_4543,N_4033);
and U4939 (N_4939,N_4039,N_4731);
xnor U4940 (N_4940,N_4689,N_4046);
xnor U4941 (N_4941,N_4674,N_4049);
and U4942 (N_4942,N_4430,N_4099);
xor U4943 (N_4943,N_4177,N_4010);
and U4944 (N_4944,N_4696,N_4466);
xor U4945 (N_4945,N_4322,N_4534);
xnor U4946 (N_4946,N_4035,N_4311);
xor U4947 (N_4947,N_4319,N_4393);
xor U4948 (N_4948,N_4207,N_4659);
or U4949 (N_4949,N_4104,N_4316);
or U4950 (N_4950,N_4006,N_4016);
nor U4951 (N_4951,N_4005,N_4327);
or U4952 (N_4952,N_4652,N_4564);
nor U4953 (N_4953,N_4042,N_4673);
nand U4954 (N_4954,N_4131,N_4030);
and U4955 (N_4955,N_4654,N_4095);
or U4956 (N_4956,N_4732,N_4245);
and U4957 (N_4957,N_4000,N_4340);
xor U4958 (N_4958,N_4551,N_4025);
nor U4959 (N_4959,N_4014,N_4764);
xor U4960 (N_4960,N_4248,N_4403);
xor U4961 (N_4961,N_4363,N_4197);
or U4962 (N_4962,N_4531,N_4593);
nor U4963 (N_4963,N_4431,N_4022);
xor U4964 (N_4964,N_4723,N_4798);
nand U4965 (N_4965,N_4417,N_4535);
or U4966 (N_4966,N_4002,N_4754);
nand U4967 (N_4967,N_4026,N_4435);
nor U4968 (N_4968,N_4580,N_4471);
nor U4969 (N_4969,N_4208,N_4298);
nand U4970 (N_4970,N_4004,N_4552);
or U4971 (N_4971,N_4100,N_4120);
and U4972 (N_4972,N_4422,N_4065);
or U4973 (N_4973,N_4633,N_4358);
or U4974 (N_4974,N_4066,N_4266);
xnor U4975 (N_4975,N_4707,N_4595);
nand U4976 (N_4976,N_4786,N_4425);
or U4977 (N_4977,N_4321,N_4533);
nand U4978 (N_4978,N_4384,N_4725);
and U4979 (N_4979,N_4715,N_4606);
or U4980 (N_4980,N_4583,N_4107);
nand U4981 (N_4981,N_4098,N_4318);
xnor U4982 (N_4982,N_4172,N_4307);
nor U4983 (N_4983,N_4132,N_4376);
or U4984 (N_4984,N_4133,N_4308);
nand U4985 (N_4985,N_4050,N_4144);
xor U4986 (N_4986,N_4282,N_4362);
nand U4987 (N_4987,N_4201,N_4147);
or U4988 (N_4988,N_4703,N_4087);
or U4989 (N_4989,N_4776,N_4092);
xor U4990 (N_4990,N_4513,N_4218);
or U4991 (N_4991,N_4672,N_4675);
and U4992 (N_4992,N_4148,N_4406);
nor U4993 (N_4993,N_4763,N_4676);
or U4994 (N_4994,N_4008,N_4424);
nand U4995 (N_4995,N_4503,N_4368);
xnor U4996 (N_4996,N_4064,N_4500);
nor U4997 (N_4997,N_4711,N_4608);
xor U4998 (N_4998,N_4331,N_4183);
nand U4999 (N_4999,N_4722,N_4530);
nand U5000 (N_5000,N_4752,N_4724);
xnor U5001 (N_5001,N_4031,N_4122);
nor U5002 (N_5002,N_4520,N_4502);
and U5003 (N_5003,N_4797,N_4785);
xnor U5004 (N_5004,N_4259,N_4001);
and U5005 (N_5005,N_4202,N_4525);
nor U5006 (N_5006,N_4788,N_4350);
nand U5007 (N_5007,N_4705,N_4778);
nand U5008 (N_5008,N_4227,N_4153);
or U5009 (N_5009,N_4656,N_4199);
xnor U5010 (N_5010,N_4636,N_4494);
nor U5011 (N_5011,N_4185,N_4276);
nand U5012 (N_5012,N_4200,N_4074);
or U5013 (N_5013,N_4512,N_4383);
nor U5014 (N_5014,N_4320,N_4297);
xnor U5015 (N_5015,N_4450,N_4304);
and U5016 (N_5016,N_4480,N_4161);
nand U5017 (N_5017,N_4084,N_4138);
and U5018 (N_5018,N_4186,N_4379);
xor U5019 (N_5019,N_4720,N_4078);
and U5020 (N_5020,N_4129,N_4464);
and U5021 (N_5021,N_4293,N_4181);
and U5022 (N_5022,N_4794,N_4233);
nor U5023 (N_5023,N_4526,N_4419);
nor U5024 (N_5024,N_4137,N_4187);
nor U5025 (N_5025,N_4744,N_4708);
xnor U5026 (N_5026,N_4516,N_4020);
or U5027 (N_5027,N_4081,N_4113);
or U5028 (N_5028,N_4505,N_4704);
or U5029 (N_5029,N_4771,N_4438);
and U5030 (N_5030,N_4457,N_4354);
and U5031 (N_5031,N_4796,N_4524);
xnor U5032 (N_5032,N_4277,N_4126);
or U5033 (N_5033,N_4287,N_4678);
xor U5034 (N_5034,N_4003,N_4655);
and U5035 (N_5035,N_4243,N_4640);
nor U5036 (N_5036,N_4134,N_4568);
xor U5037 (N_5037,N_4212,N_4063);
xor U5038 (N_5038,N_4167,N_4663);
nor U5039 (N_5039,N_4203,N_4542);
and U5040 (N_5040,N_4372,N_4077);
and U5041 (N_5041,N_4214,N_4369);
nand U5042 (N_5042,N_4407,N_4141);
xnor U5043 (N_5043,N_4615,N_4691);
or U5044 (N_5044,N_4225,N_4313);
or U5045 (N_5045,N_4371,N_4053);
xor U5046 (N_5046,N_4756,N_4777);
nor U5047 (N_5047,N_4706,N_4772);
nand U5048 (N_5048,N_4226,N_4036);
or U5049 (N_5049,N_4337,N_4270);
nor U5050 (N_5050,N_4665,N_4040);
nor U5051 (N_5051,N_4774,N_4421);
or U5052 (N_5052,N_4317,N_4075);
nor U5053 (N_5053,N_4191,N_4442);
or U5054 (N_5054,N_4255,N_4396);
and U5055 (N_5055,N_4357,N_4398);
xor U5056 (N_5056,N_4166,N_4783);
and U5057 (N_5057,N_4274,N_4271);
nor U5058 (N_5058,N_4743,N_4745);
and U5059 (N_5059,N_4729,N_4484);
and U5060 (N_5060,N_4486,N_4068);
xor U5061 (N_5061,N_4765,N_4506);
and U5062 (N_5062,N_4241,N_4013);
and U5063 (N_5063,N_4346,N_4273);
and U5064 (N_5064,N_4532,N_4427);
and U5065 (N_5065,N_4175,N_4085);
and U5066 (N_5066,N_4170,N_4388);
and U5067 (N_5067,N_4097,N_4119);
or U5068 (N_5068,N_4265,N_4478);
nor U5069 (N_5069,N_4052,N_4253);
nand U5070 (N_5070,N_4455,N_4517);
nand U5071 (N_5071,N_4605,N_4323);
nor U5072 (N_5072,N_4341,N_4490);
nor U5073 (N_5073,N_4702,N_4260);
nand U5074 (N_5074,N_4514,N_4381);
and U5075 (N_5075,N_4294,N_4762);
nor U5076 (N_5076,N_4408,N_4635);
nand U5077 (N_5077,N_4209,N_4537);
nor U5078 (N_5078,N_4173,N_4213);
xnor U5079 (N_5079,N_4198,N_4733);
and U5080 (N_5080,N_4410,N_4735);
nor U5081 (N_5081,N_4491,N_4236);
nand U5082 (N_5082,N_4224,N_4755);
nand U5083 (N_5083,N_4677,N_4597);
nand U5084 (N_5084,N_4590,N_4630);
or U5085 (N_5085,N_4657,N_4364);
nor U5086 (N_5086,N_4670,N_4751);
and U5087 (N_5087,N_4468,N_4461);
xnor U5088 (N_5088,N_4680,N_4069);
xor U5089 (N_5089,N_4456,N_4165);
xor U5090 (N_5090,N_4060,N_4339);
or U5091 (N_5091,N_4499,N_4140);
and U5092 (N_5092,N_4601,N_4048);
and U5093 (N_5093,N_4012,N_4759);
nand U5094 (N_5094,N_4546,N_4420);
xnor U5095 (N_5095,N_4257,N_4668);
xor U5096 (N_5096,N_4289,N_4594);
and U5097 (N_5097,N_4682,N_4009);
nand U5098 (N_5098,N_4647,N_4103);
xnor U5099 (N_5099,N_4096,N_4628);
and U5100 (N_5100,N_4441,N_4082);
nand U5101 (N_5101,N_4770,N_4267);
nand U5102 (N_5102,N_4527,N_4671);
or U5103 (N_5103,N_4571,N_4110);
nand U5104 (N_5104,N_4545,N_4504);
xnor U5105 (N_5105,N_4076,N_4557);
nor U5106 (N_5106,N_4559,N_4171);
xnor U5107 (N_5107,N_4324,N_4629);
nor U5108 (N_5108,N_4032,N_4493);
nor U5109 (N_5109,N_4089,N_4023);
and U5110 (N_5110,N_4658,N_4429);
or U5111 (N_5111,N_4222,N_4789);
nor U5112 (N_5112,N_4365,N_4475);
nand U5113 (N_5113,N_4439,N_4753);
and U5114 (N_5114,N_4476,N_4627);
and U5115 (N_5115,N_4437,N_4681);
or U5116 (N_5116,N_4716,N_4352);
xor U5117 (N_5117,N_4088,N_4263);
or U5118 (N_5118,N_4418,N_4444);
nor U5119 (N_5119,N_4760,N_4179);
or U5120 (N_5120,N_4547,N_4452);
and U5121 (N_5121,N_4360,N_4662);
or U5122 (N_5122,N_4231,N_4414);
and U5123 (N_5123,N_4799,N_4719);
and U5124 (N_5124,N_4698,N_4782);
xnor U5125 (N_5125,N_4625,N_4314);
nand U5126 (N_5126,N_4749,N_4558);
xor U5127 (N_5127,N_4405,N_4221);
and U5128 (N_5128,N_4795,N_4495);
xnor U5129 (N_5129,N_4604,N_4477);
nand U5130 (N_5130,N_4747,N_4090);
xnor U5131 (N_5131,N_4335,N_4162);
nor U5132 (N_5132,N_4474,N_4192);
or U5133 (N_5133,N_4538,N_4283);
nand U5134 (N_5134,N_4624,N_4528);
and U5135 (N_5135,N_4235,N_4239);
nor U5136 (N_5136,N_4432,N_4262);
xnor U5137 (N_5137,N_4529,N_4343);
or U5138 (N_5138,N_4761,N_4154);
and U5139 (N_5139,N_4790,N_4155);
or U5140 (N_5140,N_4303,N_4498);
nand U5141 (N_5141,N_4519,N_4041);
nand U5142 (N_5142,N_4114,N_4784);
or U5143 (N_5143,N_4463,N_4047);
xnor U5144 (N_5144,N_4109,N_4556);
nor U5145 (N_5145,N_4599,N_4638);
nor U5146 (N_5146,N_4305,N_4196);
xor U5147 (N_5147,N_4700,N_4548);
or U5148 (N_5148,N_4508,N_4616);
and U5149 (N_5149,N_4387,N_4688);
or U5150 (N_5150,N_4024,N_4029);
and U5151 (N_5151,N_4086,N_4712);
nor U5152 (N_5152,N_4356,N_4391);
nor U5153 (N_5153,N_4586,N_4168);
or U5154 (N_5154,N_4522,N_4582);
and U5155 (N_5155,N_4121,N_4768);
and U5156 (N_5156,N_4290,N_4057);
or U5157 (N_5157,N_4766,N_4252);
nor U5158 (N_5158,N_4718,N_4576);
nand U5159 (N_5159,N_4454,N_4397);
nor U5160 (N_5160,N_4344,N_4737);
nor U5161 (N_5161,N_4489,N_4251);
nand U5162 (N_5162,N_4423,N_4443);
or U5163 (N_5163,N_4618,N_4412);
and U5164 (N_5164,N_4193,N_4449);
xor U5165 (N_5165,N_4146,N_4411);
nand U5166 (N_5166,N_4579,N_4061);
nand U5167 (N_5167,N_4485,N_4758);
and U5168 (N_5168,N_4234,N_4592);
and U5169 (N_5169,N_4713,N_4684);
nor U5170 (N_5170,N_4479,N_4482);
and U5171 (N_5171,N_4083,N_4701);
nor U5172 (N_5172,N_4286,N_4602);
xor U5173 (N_5173,N_4730,N_4178);
nor U5174 (N_5174,N_4392,N_4188);
or U5175 (N_5175,N_4472,N_4249);
xor U5176 (N_5176,N_4620,N_4634);
and U5177 (N_5177,N_4158,N_4310);
and U5178 (N_5178,N_4626,N_4553);
or U5179 (N_5179,N_4326,N_4591);
nor U5180 (N_5180,N_4102,N_4386);
xor U5181 (N_5181,N_4507,N_4709);
or U5182 (N_5182,N_4017,N_4204);
nand U5183 (N_5183,N_4332,N_4697);
xor U5184 (N_5184,N_4072,N_4106);
and U5185 (N_5185,N_4246,N_4496);
or U5186 (N_5186,N_4555,N_4019);
and U5187 (N_5187,N_4380,N_4189);
nand U5188 (N_5188,N_4587,N_4080);
nor U5189 (N_5189,N_4549,N_4515);
xnor U5190 (N_5190,N_4639,N_4685);
nand U5191 (N_5191,N_4787,N_4440);
nand U5192 (N_5192,N_4112,N_4156);
or U5193 (N_5193,N_4573,N_4748);
and U5194 (N_5194,N_4374,N_4275);
nand U5195 (N_5195,N_4687,N_4342);
xnor U5196 (N_5196,N_4459,N_4216);
nand U5197 (N_5197,N_4055,N_4217);
or U5198 (N_5198,N_4284,N_4664);
and U5199 (N_5199,N_4603,N_4261);
xnor U5200 (N_5200,N_4332,N_4598);
nor U5201 (N_5201,N_4078,N_4035);
nor U5202 (N_5202,N_4379,N_4575);
nand U5203 (N_5203,N_4788,N_4480);
or U5204 (N_5204,N_4769,N_4711);
nand U5205 (N_5205,N_4052,N_4278);
xor U5206 (N_5206,N_4307,N_4672);
and U5207 (N_5207,N_4183,N_4082);
or U5208 (N_5208,N_4255,N_4144);
nor U5209 (N_5209,N_4376,N_4450);
or U5210 (N_5210,N_4106,N_4201);
nor U5211 (N_5211,N_4469,N_4724);
nor U5212 (N_5212,N_4005,N_4656);
nand U5213 (N_5213,N_4364,N_4794);
or U5214 (N_5214,N_4067,N_4723);
nor U5215 (N_5215,N_4000,N_4090);
or U5216 (N_5216,N_4708,N_4693);
nand U5217 (N_5217,N_4473,N_4318);
nor U5218 (N_5218,N_4564,N_4286);
nand U5219 (N_5219,N_4711,N_4201);
nand U5220 (N_5220,N_4610,N_4728);
and U5221 (N_5221,N_4650,N_4536);
or U5222 (N_5222,N_4226,N_4331);
xnor U5223 (N_5223,N_4724,N_4460);
xor U5224 (N_5224,N_4102,N_4791);
xnor U5225 (N_5225,N_4679,N_4103);
xnor U5226 (N_5226,N_4047,N_4468);
nor U5227 (N_5227,N_4248,N_4099);
xnor U5228 (N_5228,N_4695,N_4792);
nand U5229 (N_5229,N_4565,N_4603);
nor U5230 (N_5230,N_4580,N_4767);
xor U5231 (N_5231,N_4215,N_4394);
xor U5232 (N_5232,N_4429,N_4415);
and U5233 (N_5233,N_4460,N_4488);
xor U5234 (N_5234,N_4217,N_4704);
and U5235 (N_5235,N_4685,N_4533);
nand U5236 (N_5236,N_4211,N_4261);
nand U5237 (N_5237,N_4419,N_4700);
or U5238 (N_5238,N_4681,N_4175);
and U5239 (N_5239,N_4291,N_4625);
nor U5240 (N_5240,N_4442,N_4658);
xor U5241 (N_5241,N_4377,N_4650);
xor U5242 (N_5242,N_4267,N_4048);
nand U5243 (N_5243,N_4680,N_4709);
or U5244 (N_5244,N_4798,N_4281);
nor U5245 (N_5245,N_4293,N_4332);
nand U5246 (N_5246,N_4351,N_4688);
and U5247 (N_5247,N_4350,N_4404);
nand U5248 (N_5248,N_4455,N_4262);
and U5249 (N_5249,N_4337,N_4136);
nor U5250 (N_5250,N_4361,N_4654);
nand U5251 (N_5251,N_4389,N_4087);
and U5252 (N_5252,N_4006,N_4707);
nor U5253 (N_5253,N_4040,N_4496);
xor U5254 (N_5254,N_4557,N_4376);
nand U5255 (N_5255,N_4458,N_4466);
and U5256 (N_5256,N_4135,N_4110);
nand U5257 (N_5257,N_4371,N_4544);
nand U5258 (N_5258,N_4304,N_4023);
or U5259 (N_5259,N_4091,N_4470);
xor U5260 (N_5260,N_4044,N_4075);
or U5261 (N_5261,N_4564,N_4083);
nor U5262 (N_5262,N_4700,N_4758);
or U5263 (N_5263,N_4080,N_4611);
or U5264 (N_5264,N_4723,N_4108);
nand U5265 (N_5265,N_4209,N_4608);
or U5266 (N_5266,N_4331,N_4778);
nand U5267 (N_5267,N_4776,N_4072);
nand U5268 (N_5268,N_4630,N_4289);
or U5269 (N_5269,N_4519,N_4058);
nor U5270 (N_5270,N_4650,N_4582);
nor U5271 (N_5271,N_4266,N_4512);
xnor U5272 (N_5272,N_4111,N_4473);
and U5273 (N_5273,N_4205,N_4495);
and U5274 (N_5274,N_4726,N_4022);
nand U5275 (N_5275,N_4400,N_4267);
or U5276 (N_5276,N_4467,N_4785);
nor U5277 (N_5277,N_4504,N_4275);
nor U5278 (N_5278,N_4728,N_4354);
nand U5279 (N_5279,N_4541,N_4779);
xor U5280 (N_5280,N_4046,N_4094);
xnor U5281 (N_5281,N_4544,N_4755);
and U5282 (N_5282,N_4528,N_4582);
nand U5283 (N_5283,N_4068,N_4147);
and U5284 (N_5284,N_4774,N_4794);
xor U5285 (N_5285,N_4037,N_4518);
nand U5286 (N_5286,N_4008,N_4188);
nand U5287 (N_5287,N_4482,N_4669);
nand U5288 (N_5288,N_4742,N_4760);
and U5289 (N_5289,N_4176,N_4106);
xnor U5290 (N_5290,N_4758,N_4013);
or U5291 (N_5291,N_4688,N_4089);
and U5292 (N_5292,N_4788,N_4007);
nor U5293 (N_5293,N_4370,N_4291);
xor U5294 (N_5294,N_4166,N_4484);
nand U5295 (N_5295,N_4357,N_4159);
or U5296 (N_5296,N_4359,N_4535);
and U5297 (N_5297,N_4457,N_4027);
or U5298 (N_5298,N_4057,N_4103);
nor U5299 (N_5299,N_4617,N_4133);
and U5300 (N_5300,N_4154,N_4791);
and U5301 (N_5301,N_4622,N_4625);
nand U5302 (N_5302,N_4335,N_4795);
xor U5303 (N_5303,N_4643,N_4251);
and U5304 (N_5304,N_4344,N_4526);
or U5305 (N_5305,N_4782,N_4634);
xor U5306 (N_5306,N_4613,N_4081);
nor U5307 (N_5307,N_4422,N_4364);
xnor U5308 (N_5308,N_4780,N_4318);
xor U5309 (N_5309,N_4738,N_4602);
nand U5310 (N_5310,N_4508,N_4135);
and U5311 (N_5311,N_4347,N_4083);
nand U5312 (N_5312,N_4459,N_4145);
nor U5313 (N_5313,N_4329,N_4222);
xor U5314 (N_5314,N_4625,N_4177);
nand U5315 (N_5315,N_4401,N_4064);
nand U5316 (N_5316,N_4756,N_4314);
nand U5317 (N_5317,N_4724,N_4761);
nor U5318 (N_5318,N_4667,N_4178);
nor U5319 (N_5319,N_4504,N_4516);
xor U5320 (N_5320,N_4156,N_4741);
nand U5321 (N_5321,N_4763,N_4217);
nor U5322 (N_5322,N_4543,N_4105);
xor U5323 (N_5323,N_4637,N_4677);
nand U5324 (N_5324,N_4431,N_4120);
and U5325 (N_5325,N_4104,N_4583);
nand U5326 (N_5326,N_4519,N_4053);
nand U5327 (N_5327,N_4554,N_4304);
or U5328 (N_5328,N_4776,N_4636);
and U5329 (N_5329,N_4370,N_4436);
nand U5330 (N_5330,N_4209,N_4200);
nand U5331 (N_5331,N_4525,N_4560);
and U5332 (N_5332,N_4788,N_4549);
nand U5333 (N_5333,N_4628,N_4163);
nor U5334 (N_5334,N_4632,N_4783);
xnor U5335 (N_5335,N_4498,N_4511);
nor U5336 (N_5336,N_4617,N_4565);
or U5337 (N_5337,N_4602,N_4206);
nand U5338 (N_5338,N_4455,N_4571);
xor U5339 (N_5339,N_4288,N_4675);
nor U5340 (N_5340,N_4414,N_4648);
nor U5341 (N_5341,N_4399,N_4131);
nor U5342 (N_5342,N_4190,N_4204);
and U5343 (N_5343,N_4366,N_4265);
or U5344 (N_5344,N_4446,N_4419);
nor U5345 (N_5345,N_4129,N_4768);
nor U5346 (N_5346,N_4267,N_4004);
or U5347 (N_5347,N_4680,N_4379);
or U5348 (N_5348,N_4178,N_4722);
and U5349 (N_5349,N_4345,N_4371);
nand U5350 (N_5350,N_4121,N_4368);
nand U5351 (N_5351,N_4769,N_4550);
nand U5352 (N_5352,N_4535,N_4607);
xnor U5353 (N_5353,N_4146,N_4020);
nand U5354 (N_5354,N_4759,N_4020);
nor U5355 (N_5355,N_4571,N_4355);
and U5356 (N_5356,N_4651,N_4154);
xnor U5357 (N_5357,N_4075,N_4002);
or U5358 (N_5358,N_4377,N_4288);
and U5359 (N_5359,N_4467,N_4725);
and U5360 (N_5360,N_4698,N_4116);
xor U5361 (N_5361,N_4154,N_4609);
or U5362 (N_5362,N_4576,N_4617);
nand U5363 (N_5363,N_4260,N_4351);
or U5364 (N_5364,N_4592,N_4679);
xnor U5365 (N_5365,N_4781,N_4398);
nor U5366 (N_5366,N_4520,N_4278);
xor U5367 (N_5367,N_4065,N_4153);
or U5368 (N_5368,N_4006,N_4255);
nand U5369 (N_5369,N_4503,N_4594);
and U5370 (N_5370,N_4115,N_4411);
and U5371 (N_5371,N_4534,N_4254);
nand U5372 (N_5372,N_4628,N_4465);
nand U5373 (N_5373,N_4128,N_4507);
xor U5374 (N_5374,N_4393,N_4352);
xor U5375 (N_5375,N_4000,N_4739);
nand U5376 (N_5376,N_4054,N_4558);
or U5377 (N_5377,N_4551,N_4191);
or U5378 (N_5378,N_4045,N_4602);
nand U5379 (N_5379,N_4156,N_4261);
or U5380 (N_5380,N_4507,N_4063);
and U5381 (N_5381,N_4143,N_4184);
xnor U5382 (N_5382,N_4581,N_4645);
or U5383 (N_5383,N_4125,N_4510);
xnor U5384 (N_5384,N_4714,N_4752);
or U5385 (N_5385,N_4676,N_4546);
nand U5386 (N_5386,N_4173,N_4016);
nor U5387 (N_5387,N_4597,N_4276);
and U5388 (N_5388,N_4221,N_4463);
nor U5389 (N_5389,N_4358,N_4574);
and U5390 (N_5390,N_4540,N_4051);
xnor U5391 (N_5391,N_4221,N_4574);
nand U5392 (N_5392,N_4573,N_4563);
or U5393 (N_5393,N_4784,N_4233);
nand U5394 (N_5394,N_4272,N_4233);
xnor U5395 (N_5395,N_4012,N_4313);
xnor U5396 (N_5396,N_4014,N_4562);
nor U5397 (N_5397,N_4743,N_4554);
xor U5398 (N_5398,N_4315,N_4621);
xnor U5399 (N_5399,N_4549,N_4678);
and U5400 (N_5400,N_4286,N_4147);
nor U5401 (N_5401,N_4599,N_4617);
nor U5402 (N_5402,N_4794,N_4763);
xor U5403 (N_5403,N_4051,N_4774);
xor U5404 (N_5404,N_4257,N_4404);
nor U5405 (N_5405,N_4693,N_4774);
and U5406 (N_5406,N_4504,N_4720);
and U5407 (N_5407,N_4310,N_4116);
nand U5408 (N_5408,N_4419,N_4764);
nand U5409 (N_5409,N_4545,N_4112);
nand U5410 (N_5410,N_4274,N_4512);
and U5411 (N_5411,N_4321,N_4448);
xnor U5412 (N_5412,N_4716,N_4083);
nor U5413 (N_5413,N_4228,N_4654);
nor U5414 (N_5414,N_4704,N_4326);
xor U5415 (N_5415,N_4310,N_4212);
and U5416 (N_5416,N_4043,N_4195);
or U5417 (N_5417,N_4632,N_4406);
and U5418 (N_5418,N_4422,N_4512);
or U5419 (N_5419,N_4527,N_4372);
xnor U5420 (N_5420,N_4680,N_4359);
xor U5421 (N_5421,N_4397,N_4699);
xnor U5422 (N_5422,N_4647,N_4477);
or U5423 (N_5423,N_4301,N_4024);
nor U5424 (N_5424,N_4000,N_4439);
and U5425 (N_5425,N_4510,N_4553);
and U5426 (N_5426,N_4004,N_4152);
nand U5427 (N_5427,N_4712,N_4279);
or U5428 (N_5428,N_4023,N_4796);
xor U5429 (N_5429,N_4137,N_4378);
xnor U5430 (N_5430,N_4668,N_4527);
and U5431 (N_5431,N_4209,N_4091);
xor U5432 (N_5432,N_4696,N_4666);
nor U5433 (N_5433,N_4674,N_4129);
nand U5434 (N_5434,N_4704,N_4498);
nor U5435 (N_5435,N_4796,N_4557);
or U5436 (N_5436,N_4323,N_4198);
xor U5437 (N_5437,N_4482,N_4043);
or U5438 (N_5438,N_4523,N_4190);
or U5439 (N_5439,N_4016,N_4081);
nand U5440 (N_5440,N_4434,N_4376);
and U5441 (N_5441,N_4347,N_4066);
nand U5442 (N_5442,N_4324,N_4796);
or U5443 (N_5443,N_4015,N_4508);
nor U5444 (N_5444,N_4314,N_4650);
nand U5445 (N_5445,N_4321,N_4121);
nand U5446 (N_5446,N_4274,N_4056);
nor U5447 (N_5447,N_4715,N_4558);
nor U5448 (N_5448,N_4558,N_4400);
or U5449 (N_5449,N_4642,N_4485);
nor U5450 (N_5450,N_4532,N_4484);
xor U5451 (N_5451,N_4735,N_4774);
and U5452 (N_5452,N_4738,N_4021);
nand U5453 (N_5453,N_4526,N_4512);
and U5454 (N_5454,N_4026,N_4307);
nor U5455 (N_5455,N_4334,N_4027);
nor U5456 (N_5456,N_4566,N_4671);
nand U5457 (N_5457,N_4254,N_4372);
nand U5458 (N_5458,N_4396,N_4733);
nor U5459 (N_5459,N_4769,N_4055);
nor U5460 (N_5460,N_4534,N_4139);
xor U5461 (N_5461,N_4515,N_4430);
nand U5462 (N_5462,N_4210,N_4637);
or U5463 (N_5463,N_4044,N_4679);
xnor U5464 (N_5464,N_4001,N_4477);
nand U5465 (N_5465,N_4201,N_4287);
and U5466 (N_5466,N_4371,N_4182);
and U5467 (N_5467,N_4589,N_4149);
and U5468 (N_5468,N_4625,N_4677);
or U5469 (N_5469,N_4381,N_4499);
xor U5470 (N_5470,N_4237,N_4356);
nor U5471 (N_5471,N_4485,N_4609);
xor U5472 (N_5472,N_4497,N_4318);
and U5473 (N_5473,N_4552,N_4218);
nand U5474 (N_5474,N_4625,N_4055);
nor U5475 (N_5475,N_4456,N_4283);
and U5476 (N_5476,N_4602,N_4322);
xor U5477 (N_5477,N_4527,N_4382);
or U5478 (N_5478,N_4665,N_4104);
or U5479 (N_5479,N_4011,N_4633);
and U5480 (N_5480,N_4387,N_4326);
nor U5481 (N_5481,N_4270,N_4111);
xnor U5482 (N_5482,N_4320,N_4150);
nand U5483 (N_5483,N_4288,N_4046);
nand U5484 (N_5484,N_4259,N_4516);
xor U5485 (N_5485,N_4286,N_4439);
nor U5486 (N_5486,N_4284,N_4567);
nor U5487 (N_5487,N_4144,N_4550);
nor U5488 (N_5488,N_4139,N_4152);
nor U5489 (N_5489,N_4058,N_4787);
xor U5490 (N_5490,N_4394,N_4768);
xor U5491 (N_5491,N_4342,N_4156);
nor U5492 (N_5492,N_4273,N_4407);
or U5493 (N_5493,N_4206,N_4640);
and U5494 (N_5494,N_4194,N_4784);
nand U5495 (N_5495,N_4183,N_4219);
or U5496 (N_5496,N_4500,N_4283);
nand U5497 (N_5497,N_4167,N_4482);
nand U5498 (N_5498,N_4550,N_4087);
nor U5499 (N_5499,N_4091,N_4612);
or U5500 (N_5500,N_4449,N_4101);
and U5501 (N_5501,N_4123,N_4233);
nor U5502 (N_5502,N_4784,N_4059);
or U5503 (N_5503,N_4485,N_4338);
nor U5504 (N_5504,N_4204,N_4769);
nor U5505 (N_5505,N_4246,N_4459);
nand U5506 (N_5506,N_4098,N_4677);
xor U5507 (N_5507,N_4723,N_4580);
xnor U5508 (N_5508,N_4336,N_4224);
or U5509 (N_5509,N_4642,N_4035);
or U5510 (N_5510,N_4425,N_4414);
nand U5511 (N_5511,N_4625,N_4168);
nand U5512 (N_5512,N_4263,N_4026);
nand U5513 (N_5513,N_4440,N_4415);
nand U5514 (N_5514,N_4253,N_4093);
or U5515 (N_5515,N_4471,N_4339);
xnor U5516 (N_5516,N_4210,N_4078);
nor U5517 (N_5517,N_4532,N_4220);
or U5518 (N_5518,N_4513,N_4348);
nor U5519 (N_5519,N_4268,N_4560);
or U5520 (N_5520,N_4132,N_4495);
nor U5521 (N_5521,N_4722,N_4088);
and U5522 (N_5522,N_4718,N_4257);
and U5523 (N_5523,N_4092,N_4791);
or U5524 (N_5524,N_4722,N_4302);
nand U5525 (N_5525,N_4763,N_4297);
and U5526 (N_5526,N_4681,N_4134);
xor U5527 (N_5527,N_4290,N_4083);
or U5528 (N_5528,N_4295,N_4604);
nor U5529 (N_5529,N_4246,N_4042);
xor U5530 (N_5530,N_4130,N_4719);
nand U5531 (N_5531,N_4081,N_4794);
or U5532 (N_5532,N_4490,N_4684);
or U5533 (N_5533,N_4531,N_4019);
and U5534 (N_5534,N_4602,N_4562);
xor U5535 (N_5535,N_4787,N_4158);
nand U5536 (N_5536,N_4157,N_4642);
nand U5537 (N_5537,N_4122,N_4603);
or U5538 (N_5538,N_4556,N_4285);
nand U5539 (N_5539,N_4614,N_4522);
xor U5540 (N_5540,N_4469,N_4744);
nand U5541 (N_5541,N_4013,N_4023);
nand U5542 (N_5542,N_4776,N_4398);
nand U5543 (N_5543,N_4605,N_4072);
nand U5544 (N_5544,N_4726,N_4707);
and U5545 (N_5545,N_4109,N_4155);
or U5546 (N_5546,N_4464,N_4773);
xor U5547 (N_5547,N_4439,N_4480);
nor U5548 (N_5548,N_4386,N_4588);
nand U5549 (N_5549,N_4578,N_4170);
nand U5550 (N_5550,N_4083,N_4034);
xnor U5551 (N_5551,N_4782,N_4707);
nand U5552 (N_5552,N_4638,N_4187);
nor U5553 (N_5553,N_4690,N_4018);
and U5554 (N_5554,N_4461,N_4588);
xor U5555 (N_5555,N_4441,N_4255);
nand U5556 (N_5556,N_4124,N_4585);
nor U5557 (N_5557,N_4112,N_4221);
xnor U5558 (N_5558,N_4765,N_4288);
xor U5559 (N_5559,N_4107,N_4040);
or U5560 (N_5560,N_4556,N_4172);
nand U5561 (N_5561,N_4681,N_4237);
xor U5562 (N_5562,N_4557,N_4797);
and U5563 (N_5563,N_4251,N_4200);
nor U5564 (N_5564,N_4557,N_4730);
nand U5565 (N_5565,N_4317,N_4221);
and U5566 (N_5566,N_4164,N_4292);
nand U5567 (N_5567,N_4538,N_4442);
or U5568 (N_5568,N_4222,N_4634);
or U5569 (N_5569,N_4646,N_4467);
nand U5570 (N_5570,N_4108,N_4069);
xnor U5571 (N_5571,N_4714,N_4244);
xor U5572 (N_5572,N_4087,N_4405);
nand U5573 (N_5573,N_4260,N_4449);
or U5574 (N_5574,N_4742,N_4426);
and U5575 (N_5575,N_4338,N_4112);
and U5576 (N_5576,N_4127,N_4508);
and U5577 (N_5577,N_4525,N_4426);
and U5578 (N_5578,N_4615,N_4358);
and U5579 (N_5579,N_4103,N_4514);
xnor U5580 (N_5580,N_4412,N_4366);
or U5581 (N_5581,N_4456,N_4640);
nor U5582 (N_5582,N_4631,N_4034);
nor U5583 (N_5583,N_4771,N_4506);
nand U5584 (N_5584,N_4484,N_4404);
xor U5585 (N_5585,N_4452,N_4140);
or U5586 (N_5586,N_4410,N_4613);
and U5587 (N_5587,N_4128,N_4711);
nand U5588 (N_5588,N_4779,N_4409);
and U5589 (N_5589,N_4212,N_4247);
xor U5590 (N_5590,N_4180,N_4112);
xor U5591 (N_5591,N_4622,N_4712);
nor U5592 (N_5592,N_4072,N_4557);
nand U5593 (N_5593,N_4101,N_4140);
xor U5594 (N_5594,N_4279,N_4569);
or U5595 (N_5595,N_4298,N_4511);
or U5596 (N_5596,N_4630,N_4342);
and U5597 (N_5597,N_4771,N_4177);
xor U5598 (N_5598,N_4778,N_4723);
nand U5599 (N_5599,N_4131,N_4073);
nand U5600 (N_5600,N_5446,N_5253);
xor U5601 (N_5601,N_5267,N_4903);
xnor U5602 (N_5602,N_4930,N_4956);
nand U5603 (N_5603,N_4926,N_5552);
or U5604 (N_5604,N_4877,N_5046);
nor U5605 (N_5605,N_4803,N_5090);
or U5606 (N_5606,N_5403,N_5340);
nor U5607 (N_5607,N_5490,N_4876);
and U5608 (N_5608,N_5401,N_5540);
nand U5609 (N_5609,N_5445,N_5058);
or U5610 (N_5610,N_5281,N_5397);
xor U5611 (N_5611,N_5580,N_5183);
and U5612 (N_5612,N_5169,N_5032);
xnor U5613 (N_5613,N_5219,N_5459);
or U5614 (N_5614,N_5440,N_5044);
or U5615 (N_5615,N_5101,N_4970);
or U5616 (N_5616,N_4874,N_5180);
or U5617 (N_5617,N_5417,N_4906);
and U5618 (N_5618,N_4963,N_4986);
nor U5619 (N_5619,N_4967,N_4855);
nor U5620 (N_5620,N_5249,N_5235);
or U5621 (N_5621,N_5404,N_4948);
nor U5622 (N_5622,N_5163,N_5578);
or U5623 (N_5623,N_4849,N_4814);
and U5624 (N_5624,N_5413,N_4987);
xnor U5625 (N_5625,N_5184,N_5213);
nand U5626 (N_5626,N_5188,N_4910);
xnor U5627 (N_5627,N_4887,N_5530);
or U5628 (N_5628,N_4856,N_5501);
and U5629 (N_5629,N_5096,N_5551);
xor U5630 (N_5630,N_5233,N_5458);
and U5631 (N_5631,N_5041,N_5051);
and U5632 (N_5632,N_5433,N_5149);
or U5633 (N_5633,N_4827,N_5504);
and U5634 (N_5634,N_5415,N_5400);
xnor U5635 (N_5635,N_5001,N_4811);
nand U5636 (N_5636,N_5088,N_5048);
and U5637 (N_5637,N_5547,N_5229);
nand U5638 (N_5638,N_5443,N_4944);
or U5639 (N_5639,N_5174,N_5170);
xnor U5640 (N_5640,N_4808,N_4936);
nor U5641 (N_5641,N_5211,N_4823);
xor U5642 (N_5642,N_5338,N_5224);
or U5643 (N_5643,N_4960,N_4833);
nor U5644 (N_5644,N_4990,N_5526);
nor U5645 (N_5645,N_5316,N_4866);
nor U5646 (N_5646,N_5270,N_5296);
and U5647 (N_5647,N_5061,N_5276);
nor U5648 (N_5648,N_5099,N_5008);
nand U5649 (N_5649,N_5015,N_4820);
or U5650 (N_5650,N_5082,N_5065);
nor U5651 (N_5651,N_5587,N_4891);
nor U5652 (N_5652,N_4805,N_5287);
xnor U5653 (N_5653,N_5579,N_5437);
or U5654 (N_5654,N_4882,N_5487);
nand U5655 (N_5655,N_5478,N_4983);
or U5656 (N_5656,N_4994,N_5531);
or U5657 (N_5657,N_5215,N_5042);
nor U5658 (N_5658,N_5411,N_5200);
xnor U5659 (N_5659,N_5012,N_5039);
or U5660 (N_5660,N_5535,N_5595);
nand U5661 (N_5661,N_5473,N_5262);
or U5662 (N_5662,N_5185,N_5310);
and U5663 (N_5663,N_4872,N_5289);
nor U5664 (N_5664,N_5545,N_5223);
xnor U5665 (N_5665,N_5343,N_5141);
xor U5666 (N_5666,N_5391,N_5585);
and U5667 (N_5667,N_4974,N_5366);
xnor U5668 (N_5668,N_5512,N_5286);
xnor U5669 (N_5669,N_5410,N_5346);
xnor U5670 (N_5670,N_5546,N_5221);
xor U5671 (N_5671,N_5383,N_5306);
nor U5672 (N_5672,N_5399,N_4892);
xnor U5673 (N_5673,N_4865,N_5152);
nor U5674 (N_5674,N_5384,N_5029);
and U5675 (N_5675,N_5536,N_4888);
xor U5676 (N_5676,N_4928,N_5105);
nor U5677 (N_5677,N_5034,N_4869);
and U5678 (N_5678,N_4884,N_5124);
nand U5679 (N_5679,N_5006,N_5145);
or U5680 (N_5680,N_4980,N_4992);
nand U5681 (N_5681,N_5130,N_5293);
xnor U5682 (N_5682,N_5351,N_4819);
or U5683 (N_5683,N_4900,N_5059);
or U5684 (N_5684,N_5414,N_4879);
or U5685 (N_5685,N_5158,N_5495);
and U5686 (N_5686,N_4896,N_5576);
nor U5687 (N_5687,N_5325,N_5011);
nor U5688 (N_5688,N_5481,N_5568);
nand U5689 (N_5689,N_5322,N_5005);
nor U5690 (N_5690,N_4800,N_5218);
xnor U5691 (N_5691,N_5412,N_5592);
and U5692 (N_5692,N_5497,N_5376);
or U5693 (N_5693,N_5146,N_4802);
or U5694 (N_5694,N_5225,N_5055);
nor U5695 (N_5695,N_4828,N_5070);
or U5696 (N_5696,N_5004,N_5189);
nand U5697 (N_5697,N_5147,N_5460);
nor U5698 (N_5698,N_5066,N_5181);
and U5699 (N_5699,N_4871,N_4890);
xor U5700 (N_5700,N_5024,N_5398);
and U5701 (N_5701,N_5419,N_4821);
xor U5702 (N_5702,N_5331,N_5596);
or U5703 (N_5703,N_5395,N_5332);
nand U5704 (N_5704,N_4950,N_5407);
and U5705 (N_5705,N_5110,N_5354);
or U5706 (N_5706,N_5186,N_5301);
nor U5707 (N_5707,N_5379,N_5361);
or U5708 (N_5708,N_5447,N_5421);
nand U5709 (N_5709,N_5555,N_5360);
or U5710 (N_5710,N_4964,N_5291);
or U5711 (N_5711,N_5216,N_5484);
or U5712 (N_5712,N_4846,N_5236);
nand U5713 (N_5713,N_5341,N_5556);
or U5714 (N_5714,N_4925,N_4893);
xor U5715 (N_5715,N_4985,N_5052);
nor U5716 (N_5716,N_4895,N_5190);
or U5717 (N_5717,N_5599,N_5247);
xor U5718 (N_5718,N_5021,N_5314);
and U5719 (N_5719,N_5230,N_4920);
and U5720 (N_5720,N_4946,N_4966);
and U5721 (N_5721,N_5295,N_5272);
and U5722 (N_5722,N_5258,N_5309);
or U5723 (N_5723,N_5378,N_5388);
and U5724 (N_5724,N_5476,N_5122);
and U5725 (N_5725,N_4839,N_5373);
nor U5726 (N_5726,N_5570,N_5496);
nor U5727 (N_5727,N_5102,N_5329);
and U5728 (N_5728,N_5468,N_5483);
or U5729 (N_5729,N_5420,N_5246);
nor U5730 (N_5730,N_4894,N_4873);
xor U5731 (N_5731,N_5464,N_5299);
xor U5732 (N_5732,N_5479,N_5566);
and U5733 (N_5733,N_4982,N_5517);
and U5734 (N_5734,N_5462,N_4947);
nand U5735 (N_5735,N_4911,N_5320);
nor U5736 (N_5736,N_5493,N_4813);
and U5737 (N_5737,N_5371,N_5591);
nand U5738 (N_5738,N_5164,N_4861);
and U5739 (N_5739,N_5231,N_5173);
nor U5740 (N_5740,N_5486,N_5358);
xor U5741 (N_5741,N_5520,N_5393);
nand U5742 (N_5742,N_5598,N_5569);
or U5743 (N_5743,N_4853,N_5285);
and U5744 (N_5744,N_5007,N_4968);
nor U5745 (N_5745,N_5503,N_5157);
or U5746 (N_5746,N_5423,N_5313);
nand U5747 (N_5747,N_4868,N_5385);
nor U5748 (N_5748,N_5434,N_5359);
and U5749 (N_5749,N_4996,N_4862);
or U5750 (N_5750,N_5060,N_5129);
nor U5751 (N_5751,N_4914,N_5557);
and U5752 (N_5752,N_5162,N_5513);
or U5753 (N_5753,N_4999,N_5264);
xnor U5754 (N_5754,N_4935,N_5212);
nand U5755 (N_5755,N_5121,N_5037);
nand U5756 (N_5756,N_5192,N_5357);
nand U5757 (N_5757,N_5352,N_5553);
xnor U5758 (N_5758,N_5594,N_4850);
or U5759 (N_5759,N_5138,N_5337);
nand U5760 (N_5760,N_4810,N_5047);
or U5761 (N_5761,N_4918,N_4975);
xor U5762 (N_5762,N_5097,N_5374);
and U5763 (N_5763,N_5127,N_5333);
and U5764 (N_5764,N_4934,N_5210);
or U5765 (N_5765,N_5197,N_5133);
xor U5766 (N_5766,N_4834,N_5155);
or U5767 (N_5767,N_5193,N_5448);
nor U5768 (N_5768,N_5307,N_5382);
or U5769 (N_5769,N_4816,N_5087);
nand U5770 (N_5770,N_5550,N_4817);
xor U5771 (N_5771,N_5475,N_4881);
xnor U5772 (N_5772,N_4848,N_5139);
or U5773 (N_5773,N_5069,N_5115);
or U5774 (N_5774,N_4940,N_5456);
xor U5775 (N_5775,N_5284,N_5261);
nand U5776 (N_5776,N_5593,N_5525);
nand U5777 (N_5777,N_4984,N_5406);
xor U5778 (N_5778,N_4860,N_5117);
and U5779 (N_5779,N_5134,N_5143);
or U5780 (N_5780,N_5118,N_4991);
nand U5781 (N_5781,N_5237,N_4883);
and U5782 (N_5782,N_5040,N_5156);
nand U5783 (N_5783,N_5315,N_5450);
nand U5784 (N_5784,N_5377,N_4922);
nor U5785 (N_5785,N_5418,N_5187);
xor U5786 (N_5786,N_5111,N_5031);
and U5787 (N_5787,N_5241,N_5150);
nor U5788 (N_5788,N_5436,N_5516);
or U5789 (N_5789,N_5319,N_4942);
nor U5790 (N_5790,N_4943,N_5000);
and U5791 (N_5791,N_5502,N_5120);
or U5792 (N_5792,N_5126,N_5489);
xor U5793 (N_5793,N_5084,N_4806);
nor U5794 (N_5794,N_5292,N_5288);
nand U5795 (N_5795,N_5494,N_5523);
xor U5796 (N_5796,N_5349,N_4864);
or U5797 (N_5797,N_4953,N_4863);
xor U5798 (N_5798,N_4945,N_5203);
nand U5799 (N_5799,N_5030,N_4878);
nor U5800 (N_5800,N_4807,N_5144);
xnor U5801 (N_5801,N_5266,N_5112);
and U5802 (N_5802,N_4841,N_5348);
nand U5803 (N_5803,N_5022,N_5471);
and U5804 (N_5804,N_5256,N_5098);
xnor U5805 (N_5805,N_5424,N_5064);
nand U5806 (N_5806,N_4858,N_5511);
and U5807 (N_5807,N_5466,N_5137);
nand U5808 (N_5808,N_4976,N_5375);
and U5809 (N_5809,N_4949,N_5506);
nor U5810 (N_5810,N_5431,N_5049);
nand U5811 (N_5811,N_5567,N_4957);
xnor U5812 (N_5812,N_5364,N_5106);
and U5813 (N_5813,N_4885,N_5027);
xor U5814 (N_5814,N_4978,N_4919);
and U5815 (N_5815,N_4826,N_4916);
nor U5816 (N_5816,N_4835,N_5532);
nor U5817 (N_5817,N_5191,N_5581);
xor U5818 (N_5818,N_5271,N_4837);
nand U5819 (N_5819,N_5571,N_4954);
nor U5820 (N_5820,N_5075,N_5019);
nand U5821 (N_5821,N_5275,N_5202);
nor U5822 (N_5822,N_5076,N_5508);
nand U5823 (N_5823,N_5500,N_5527);
nor U5824 (N_5824,N_4815,N_5470);
nor U5825 (N_5825,N_5543,N_5318);
nor U5826 (N_5826,N_5442,N_5323);
nand U5827 (N_5827,N_5154,N_5043);
nor U5828 (N_5828,N_5148,N_5123);
nand U5829 (N_5829,N_5482,N_5251);
or U5830 (N_5830,N_5263,N_5480);
nand U5831 (N_5831,N_5367,N_5577);
xor U5832 (N_5832,N_4981,N_5025);
nand U5833 (N_5833,N_5350,N_4962);
xor U5834 (N_5834,N_4843,N_5588);
xor U5835 (N_5835,N_5334,N_5204);
or U5836 (N_5836,N_5018,N_5441);
and U5837 (N_5837,N_5104,N_5582);
xor U5838 (N_5838,N_5438,N_5386);
xnor U5839 (N_5839,N_4908,N_5159);
nor U5840 (N_5840,N_5558,N_5160);
xnor U5841 (N_5841,N_5166,N_5227);
and U5842 (N_5842,N_5045,N_5245);
nor U5843 (N_5843,N_5091,N_5273);
and U5844 (N_5844,N_4838,N_5505);
and U5845 (N_5845,N_5387,N_5402);
or U5846 (N_5846,N_5259,N_5542);
and U5847 (N_5847,N_5426,N_5089);
xnor U5848 (N_5848,N_5498,N_4915);
xor U5849 (N_5849,N_4857,N_5073);
and U5850 (N_5850,N_5232,N_4917);
nand U5851 (N_5851,N_5208,N_5297);
and U5852 (N_5852,N_5394,N_4899);
nor U5853 (N_5853,N_5209,N_4804);
nand U5854 (N_5854,N_5549,N_5078);
nor U5855 (N_5855,N_5584,N_5002);
and U5856 (N_5856,N_5269,N_5151);
and U5857 (N_5857,N_5093,N_5336);
nor U5858 (N_5858,N_5108,N_5092);
or U5859 (N_5859,N_5194,N_5422);
and U5860 (N_5860,N_4965,N_5339);
nand U5861 (N_5861,N_5474,N_5226);
nor U5862 (N_5862,N_5353,N_5198);
xnor U5863 (N_5863,N_5100,N_5079);
and U5864 (N_5864,N_5453,N_5279);
xnor U5865 (N_5865,N_5242,N_5063);
nand U5866 (N_5866,N_5303,N_4847);
xor U5867 (N_5867,N_4842,N_5107);
nor U5868 (N_5868,N_5363,N_5589);
nor U5869 (N_5869,N_5205,N_5548);
or U5870 (N_5870,N_5068,N_5435);
and U5871 (N_5871,N_4897,N_5563);
nand U5872 (N_5872,N_5176,N_5268);
nor U5873 (N_5873,N_4845,N_5081);
xor U5874 (N_5874,N_4886,N_5033);
and U5875 (N_5875,N_5326,N_5425);
and U5876 (N_5876,N_5228,N_5294);
and U5877 (N_5877,N_5214,N_4822);
nand U5878 (N_5878,N_5153,N_5035);
xnor U5879 (N_5879,N_5392,N_5522);
or U5880 (N_5880,N_5240,N_5572);
or U5881 (N_5881,N_5175,N_4938);
xnor U5882 (N_5882,N_4927,N_4812);
nand U5883 (N_5883,N_5491,N_5086);
and U5884 (N_5884,N_4840,N_5128);
xnor U5885 (N_5885,N_4952,N_5463);
or U5886 (N_5886,N_5564,N_5539);
xnor U5887 (N_5887,N_5455,N_5510);
xor U5888 (N_5888,N_5537,N_5283);
or U5889 (N_5889,N_4844,N_5072);
nor U5890 (N_5890,N_5389,N_5586);
xnor U5891 (N_5891,N_5300,N_5161);
or U5892 (N_5892,N_5003,N_5023);
nand U5893 (N_5893,N_5590,N_5195);
nand U5894 (N_5894,N_5290,N_5172);
nand U5895 (N_5895,N_5499,N_4832);
or U5896 (N_5896,N_4901,N_5477);
xnor U5897 (N_5897,N_5238,N_5432);
nor U5898 (N_5898,N_5196,N_5461);
nor U5899 (N_5899,N_5524,N_5243);
or U5900 (N_5900,N_4995,N_4997);
xor U5901 (N_5901,N_5125,N_5429);
xnor U5902 (N_5902,N_5171,N_5178);
nor U5903 (N_5903,N_5427,N_4972);
xnor U5904 (N_5904,N_4924,N_5013);
or U5905 (N_5905,N_5344,N_4958);
nand U5906 (N_5906,N_5597,N_5472);
or U5907 (N_5907,N_5328,N_4830);
or U5908 (N_5908,N_5050,N_5492);
nand U5909 (N_5909,N_4955,N_5408);
nor U5910 (N_5910,N_5182,N_5298);
and U5911 (N_5911,N_5368,N_4898);
nand U5912 (N_5912,N_5330,N_5509);
or U5913 (N_5913,N_5206,N_5083);
or U5914 (N_5914,N_5282,N_4979);
xnor U5915 (N_5915,N_5365,N_5380);
nand U5916 (N_5916,N_4932,N_5053);
nor U5917 (N_5917,N_5136,N_5405);
and U5918 (N_5918,N_5485,N_5324);
nand U5919 (N_5919,N_5177,N_5428);
nand U5920 (N_5920,N_5519,N_4977);
nand U5921 (N_5921,N_5062,N_4902);
nor U5922 (N_5922,N_5521,N_5056);
xor U5923 (N_5923,N_5559,N_4824);
and U5924 (N_5924,N_4889,N_5317);
xnor U5925 (N_5925,N_5109,N_4961);
or U5926 (N_5926,N_5057,N_5560);
nor U5927 (N_5927,N_5217,N_5356);
xnor U5928 (N_5928,N_5469,N_5095);
nor U5929 (N_5929,N_4859,N_5507);
or U5930 (N_5930,N_5515,N_5038);
nand U5931 (N_5931,N_4913,N_5074);
and U5932 (N_5932,N_5538,N_4951);
xor U5933 (N_5933,N_5142,N_5451);
or U5934 (N_5934,N_5009,N_5449);
and U5935 (N_5935,N_5321,N_5454);
nand U5936 (N_5936,N_5179,N_5430);
or U5937 (N_5937,N_4831,N_5244);
nor U5938 (N_5938,N_5119,N_5071);
or U5939 (N_5939,N_5248,N_4941);
nand U5940 (N_5940,N_4973,N_5103);
or U5941 (N_5941,N_4875,N_5278);
nor U5942 (N_5942,N_5311,N_5312);
and U5943 (N_5943,N_5201,N_4939);
xnor U5944 (N_5944,N_5080,N_5304);
or U5945 (N_5945,N_5010,N_4912);
nor U5946 (N_5946,N_5544,N_5573);
or U5947 (N_5947,N_4801,N_5014);
nand U5948 (N_5948,N_4851,N_5583);
nand U5949 (N_5949,N_5094,N_5467);
nand U5950 (N_5950,N_5529,N_5575);
nor U5951 (N_5951,N_5132,N_5199);
and U5952 (N_5952,N_4971,N_5554);
xnor U5953 (N_5953,N_5077,N_4989);
or U5954 (N_5954,N_5239,N_5265);
and U5955 (N_5955,N_5280,N_5054);
and U5956 (N_5956,N_5308,N_5207);
nor U5957 (N_5957,N_5355,N_5302);
or U5958 (N_5958,N_5345,N_5565);
nor U5959 (N_5959,N_5257,N_5116);
nand U5960 (N_5960,N_4852,N_4993);
or U5961 (N_5961,N_5342,N_5347);
nor U5962 (N_5962,N_5234,N_4937);
xnor U5963 (N_5963,N_4867,N_5114);
nor U5964 (N_5964,N_5335,N_5518);
nand U5965 (N_5965,N_5465,N_5409);
xnor U5966 (N_5966,N_4923,N_5561);
nor U5967 (N_5967,N_4931,N_5131);
and U5968 (N_5968,N_5372,N_5533);
or U5969 (N_5969,N_4909,N_5305);
nand U5970 (N_5970,N_5416,N_5541);
or U5971 (N_5971,N_5113,N_5255);
nand U5972 (N_5972,N_5140,N_5067);
and U5973 (N_5973,N_5167,N_4929);
or U5974 (N_5974,N_5085,N_5444);
xnor U5975 (N_5975,N_4825,N_5362);
xnor U5976 (N_5976,N_5026,N_5168);
nand U5977 (N_5977,N_5135,N_5222);
xor U5978 (N_5978,N_4988,N_5488);
xor U5979 (N_5979,N_5250,N_5452);
and U5980 (N_5980,N_5017,N_4969);
nor U5981 (N_5981,N_5036,N_5254);
xor U5982 (N_5982,N_5252,N_4921);
or U5983 (N_5983,N_5370,N_5327);
or U5984 (N_5984,N_5020,N_4905);
xor U5985 (N_5985,N_5369,N_4959);
nor U5986 (N_5986,N_4870,N_5562);
nand U5987 (N_5987,N_5574,N_4809);
xnor U5988 (N_5988,N_4854,N_5396);
nand U5989 (N_5989,N_5260,N_5390);
or U5990 (N_5990,N_5274,N_4880);
nand U5991 (N_5991,N_5534,N_5016);
xor U5992 (N_5992,N_4836,N_5165);
xor U5993 (N_5993,N_4998,N_4904);
nand U5994 (N_5994,N_4907,N_5277);
xor U5995 (N_5995,N_5457,N_5220);
and U5996 (N_5996,N_4829,N_5439);
xor U5997 (N_5997,N_5514,N_5381);
nor U5998 (N_5998,N_4818,N_5028);
nor U5999 (N_5999,N_4933,N_5528);
or U6000 (N_6000,N_5407,N_5206);
xor U6001 (N_6001,N_5294,N_5425);
xor U6002 (N_6002,N_5429,N_4962);
or U6003 (N_6003,N_5426,N_5036);
or U6004 (N_6004,N_5069,N_5128);
xor U6005 (N_6005,N_5459,N_5036);
nor U6006 (N_6006,N_5145,N_5200);
and U6007 (N_6007,N_5246,N_5421);
or U6008 (N_6008,N_5312,N_5591);
nor U6009 (N_6009,N_4935,N_4944);
nand U6010 (N_6010,N_5415,N_5132);
or U6011 (N_6011,N_5284,N_5306);
xnor U6012 (N_6012,N_5240,N_5537);
nor U6013 (N_6013,N_5148,N_5227);
xnor U6014 (N_6014,N_5033,N_5248);
xor U6015 (N_6015,N_5287,N_4881);
and U6016 (N_6016,N_5132,N_4884);
and U6017 (N_6017,N_5385,N_4880);
nor U6018 (N_6018,N_5188,N_5550);
nand U6019 (N_6019,N_5001,N_5396);
nor U6020 (N_6020,N_5196,N_4836);
and U6021 (N_6021,N_5010,N_4877);
or U6022 (N_6022,N_5015,N_4801);
nor U6023 (N_6023,N_4993,N_5526);
xnor U6024 (N_6024,N_4845,N_5401);
or U6025 (N_6025,N_5382,N_5179);
xnor U6026 (N_6026,N_5473,N_5571);
or U6027 (N_6027,N_5339,N_5480);
or U6028 (N_6028,N_5394,N_5364);
and U6029 (N_6029,N_5144,N_5157);
and U6030 (N_6030,N_5182,N_5315);
nor U6031 (N_6031,N_5153,N_4836);
nor U6032 (N_6032,N_5117,N_5508);
xnor U6033 (N_6033,N_5036,N_4901);
and U6034 (N_6034,N_5446,N_4859);
nor U6035 (N_6035,N_5102,N_5139);
or U6036 (N_6036,N_5584,N_5519);
and U6037 (N_6037,N_5093,N_5447);
nor U6038 (N_6038,N_5248,N_5041);
or U6039 (N_6039,N_4974,N_5021);
nor U6040 (N_6040,N_5060,N_5546);
xor U6041 (N_6041,N_5096,N_5021);
nor U6042 (N_6042,N_5395,N_5567);
or U6043 (N_6043,N_5107,N_5071);
nand U6044 (N_6044,N_5149,N_4982);
nand U6045 (N_6045,N_5082,N_5450);
nor U6046 (N_6046,N_5086,N_4925);
nand U6047 (N_6047,N_5391,N_5498);
nand U6048 (N_6048,N_4886,N_4877);
nor U6049 (N_6049,N_5130,N_5043);
nand U6050 (N_6050,N_5278,N_4829);
or U6051 (N_6051,N_4820,N_5220);
xnor U6052 (N_6052,N_5185,N_4965);
and U6053 (N_6053,N_5111,N_5036);
nand U6054 (N_6054,N_5158,N_4850);
nor U6055 (N_6055,N_5290,N_5138);
nand U6056 (N_6056,N_4977,N_5221);
xnor U6057 (N_6057,N_5333,N_4813);
or U6058 (N_6058,N_5222,N_5086);
or U6059 (N_6059,N_4800,N_4882);
and U6060 (N_6060,N_5466,N_5245);
xnor U6061 (N_6061,N_5549,N_4932);
nor U6062 (N_6062,N_5289,N_4855);
xor U6063 (N_6063,N_5493,N_5411);
and U6064 (N_6064,N_4977,N_5154);
nand U6065 (N_6065,N_5000,N_5526);
and U6066 (N_6066,N_5064,N_5252);
xnor U6067 (N_6067,N_5223,N_4912);
nand U6068 (N_6068,N_5185,N_5444);
xnor U6069 (N_6069,N_5128,N_5017);
and U6070 (N_6070,N_5186,N_5515);
nor U6071 (N_6071,N_5042,N_4804);
xnor U6072 (N_6072,N_5084,N_5576);
xor U6073 (N_6073,N_5383,N_5589);
nand U6074 (N_6074,N_5384,N_5433);
nand U6075 (N_6075,N_4823,N_5324);
nand U6076 (N_6076,N_5174,N_5126);
nand U6077 (N_6077,N_5455,N_4978);
and U6078 (N_6078,N_5444,N_5340);
and U6079 (N_6079,N_5140,N_5007);
nand U6080 (N_6080,N_5078,N_4972);
nor U6081 (N_6081,N_4908,N_5002);
or U6082 (N_6082,N_4819,N_5047);
xnor U6083 (N_6083,N_4850,N_5502);
and U6084 (N_6084,N_5276,N_4936);
or U6085 (N_6085,N_5416,N_5008);
xnor U6086 (N_6086,N_5117,N_5328);
nand U6087 (N_6087,N_4857,N_5494);
or U6088 (N_6088,N_5456,N_5136);
or U6089 (N_6089,N_5469,N_5224);
or U6090 (N_6090,N_5107,N_5547);
nor U6091 (N_6091,N_4967,N_5338);
nor U6092 (N_6092,N_5511,N_5568);
nand U6093 (N_6093,N_5205,N_5002);
nand U6094 (N_6094,N_5076,N_4916);
or U6095 (N_6095,N_5415,N_5402);
or U6096 (N_6096,N_5135,N_5430);
nand U6097 (N_6097,N_5485,N_5214);
nor U6098 (N_6098,N_5199,N_5045);
and U6099 (N_6099,N_5356,N_4806);
nand U6100 (N_6100,N_4965,N_4890);
and U6101 (N_6101,N_5408,N_5201);
xor U6102 (N_6102,N_5358,N_5373);
and U6103 (N_6103,N_5200,N_5383);
or U6104 (N_6104,N_4958,N_5555);
or U6105 (N_6105,N_5060,N_5554);
or U6106 (N_6106,N_5155,N_4946);
or U6107 (N_6107,N_5215,N_4964);
xnor U6108 (N_6108,N_5075,N_5558);
nand U6109 (N_6109,N_5304,N_5510);
or U6110 (N_6110,N_5074,N_4837);
or U6111 (N_6111,N_5281,N_5163);
xnor U6112 (N_6112,N_5391,N_5342);
xnor U6113 (N_6113,N_4881,N_5053);
nand U6114 (N_6114,N_5253,N_5523);
nand U6115 (N_6115,N_4912,N_5471);
xnor U6116 (N_6116,N_5039,N_5235);
nand U6117 (N_6117,N_5381,N_5018);
nand U6118 (N_6118,N_5053,N_5455);
nand U6119 (N_6119,N_4881,N_5028);
or U6120 (N_6120,N_5078,N_4853);
nand U6121 (N_6121,N_5073,N_5569);
and U6122 (N_6122,N_5336,N_5446);
or U6123 (N_6123,N_5461,N_5568);
nor U6124 (N_6124,N_5098,N_4802);
or U6125 (N_6125,N_4867,N_5260);
nor U6126 (N_6126,N_4876,N_5597);
nand U6127 (N_6127,N_5420,N_4806);
or U6128 (N_6128,N_4942,N_5144);
or U6129 (N_6129,N_4811,N_5433);
nor U6130 (N_6130,N_5502,N_5109);
nand U6131 (N_6131,N_4964,N_5413);
xor U6132 (N_6132,N_5202,N_4955);
and U6133 (N_6133,N_4821,N_5178);
xnor U6134 (N_6134,N_4975,N_5372);
nor U6135 (N_6135,N_4916,N_5403);
nand U6136 (N_6136,N_4914,N_5079);
or U6137 (N_6137,N_4878,N_5445);
nand U6138 (N_6138,N_5309,N_5378);
and U6139 (N_6139,N_5428,N_4852);
or U6140 (N_6140,N_5273,N_5108);
nor U6141 (N_6141,N_5337,N_5128);
xnor U6142 (N_6142,N_5110,N_5220);
and U6143 (N_6143,N_5400,N_4820);
nor U6144 (N_6144,N_5448,N_5372);
or U6145 (N_6145,N_5558,N_5413);
xnor U6146 (N_6146,N_5397,N_5029);
nor U6147 (N_6147,N_5162,N_5457);
or U6148 (N_6148,N_4860,N_4896);
or U6149 (N_6149,N_5140,N_5464);
or U6150 (N_6150,N_5326,N_5226);
nor U6151 (N_6151,N_5116,N_5502);
nor U6152 (N_6152,N_4893,N_5559);
nand U6153 (N_6153,N_5092,N_5220);
xnor U6154 (N_6154,N_5090,N_4897);
xor U6155 (N_6155,N_5403,N_5156);
or U6156 (N_6156,N_5094,N_5163);
and U6157 (N_6157,N_5349,N_5113);
and U6158 (N_6158,N_5175,N_5526);
nor U6159 (N_6159,N_5383,N_5269);
nand U6160 (N_6160,N_5006,N_5427);
or U6161 (N_6161,N_5316,N_4876);
nor U6162 (N_6162,N_5581,N_5042);
and U6163 (N_6163,N_5053,N_5477);
nor U6164 (N_6164,N_4953,N_5436);
and U6165 (N_6165,N_4997,N_5052);
nand U6166 (N_6166,N_5114,N_5502);
and U6167 (N_6167,N_4957,N_5485);
nand U6168 (N_6168,N_5249,N_5209);
or U6169 (N_6169,N_4879,N_5148);
xor U6170 (N_6170,N_5390,N_5113);
or U6171 (N_6171,N_5494,N_4847);
or U6172 (N_6172,N_5440,N_5368);
xor U6173 (N_6173,N_4879,N_5430);
nor U6174 (N_6174,N_5101,N_5338);
and U6175 (N_6175,N_4963,N_5130);
nor U6176 (N_6176,N_5425,N_5557);
xnor U6177 (N_6177,N_5044,N_5551);
nor U6178 (N_6178,N_4851,N_5037);
and U6179 (N_6179,N_5064,N_5036);
nor U6180 (N_6180,N_4851,N_5568);
xor U6181 (N_6181,N_5590,N_5349);
nand U6182 (N_6182,N_4913,N_5369);
nor U6183 (N_6183,N_5219,N_5450);
or U6184 (N_6184,N_5258,N_5549);
nor U6185 (N_6185,N_5442,N_5274);
or U6186 (N_6186,N_5301,N_5077);
or U6187 (N_6187,N_5292,N_5170);
nor U6188 (N_6188,N_5421,N_5040);
xor U6189 (N_6189,N_5588,N_4957);
or U6190 (N_6190,N_5584,N_5489);
xnor U6191 (N_6191,N_5195,N_5533);
nor U6192 (N_6192,N_5153,N_5563);
nand U6193 (N_6193,N_5591,N_5032);
nand U6194 (N_6194,N_5349,N_4872);
nand U6195 (N_6195,N_4934,N_5582);
or U6196 (N_6196,N_4954,N_5172);
nand U6197 (N_6197,N_5239,N_5457);
and U6198 (N_6198,N_5490,N_4980);
or U6199 (N_6199,N_5125,N_4839);
nor U6200 (N_6200,N_4888,N_5126);
xor U6201 (N_6201,N_4860,N_5463);
xor U6202 (N_6202,N_4967,N_4954);
nand U6203 (N_6203,N_5240,N_5588);
and U6204 (N_6204,N_5206,N_4824);
or U6205 (N_6205,N_5280,N_5368);
and U6206 (N_6206,N_4925,N_5593);
nor U6207 (N_6207,N_5411,N_5314);
xor U6208 (N_6208,N_5217,N_5529);
nand U6209 (N_6209,N_5540,N_4945);
nor U6210 (N_6210,N_5122,N_4972);
and U6211 (N_6211,N_5276,N_5581);
and U6212 (N_6212,N_4815,N_5403);
nand U6213 (N_6213,N_5308,N_5574);
nor U6214 (N_6214,N_5080,N_5322);
and U6215 (N_6215,N_4921,N_4867);
nand U6216 (N_6216,N_4840,N_5144);
nor U6217 (N_6217,N_5047,N_5063);
or U6218 (N_6218,N_5564,N_4880);
nor U6219 (N_6219,N_5502,N_4802);
xnor U6220 (N_6220,N_5372,N_5043);
nor U6221 (N_6221,N_5155,N_4951);
or U6222 (N_6222,N_5153,N_5265);
nand U6223 (N_6223,N_5384,N_5274);
nand U6224 (N_6224,N_5580,N_5079);
nand U6225 (N_6225,N_5580,N_5269);
nand U6226 (N_6226,N_5134,N_4867);
and U6227 (N_6227,N_5573,N_5278);
or U6228 (N_6228,N_5482,N_5590);
nand U6229 (N_6229,N_5296,N_5127);
or U6230 (N_6230,N_5229,N_4931);
nor U6231 (N_6231,N_5277,N_5030);
nand U6232 (N_6232,N_4946,N_5208);
or U6233 (N_6233,N_5097,N_5211);
or U6234 (N_6234,N_5126,N_5302);
and U6235 (N_6235,N_4910,N_5360);
nor U6236 (N_6236,N_5250,N_5222);
or U6237 (N_6237,N_5148,N_5088);
nand U6238 (N_6238,N_4922,N_4913);
nand U6239 (N_6239,N_5598,N_4806);
nand U6240 (N_6240,N_5018,N_5456);
nor U6241 (N_6241,N_5229,N_4894);
and U6242 (N_6242,N_4933,N_5476);
xnor U6243 (N_6243,N_5470,N_5018);
xnor U6244 (N_6244,N_4829,N_5355);
nor U6245 (N_6245,N_5378,N_5401);
or U6246 (N_6246,N_5198,N_5555);
nor U6247 (N_6247,N_4944,N_5145);
and U6248 (N_6248,N_5336,N_5260);
or U6249 (N_6249,N_5188,N_5269);
nor U6250 (N_6250,N_4863,N_5406);
or U6251 (N_6251,N_4959,N_5367);
xnor U6252 (N_6252,N_4951,N_4814);
nand U6253 (N_6253,N_5433,N_5484);
or U6254 (N_6254,N_4953,N_5172);
or U6255 (N_6255,N_5260,N_4919);
or U6256 (N_6256,N_5166,N_5538);
nor U6257 (N_6257,N_4965,N_5353);
nand U6258 (N_6258,N_4849,N_4859);
and U6259 (N_6259,N_4955,N_5156);
nor U6260 (N_6260,N_5083,N_5138);
nor U6261 (N_6261,N_5374,N_5030);
or U6262 (N_6262,N_5455,N_5491);
xor U6263 (N_6263,N_5410,N_5375);
xor U6264 (N_6264,N_5087,N_4930);
nor U6265 (N_6265,N_5568,N_5329);
or U6266 (N_6266,N_5418,N_4966);
nor U6267 (N_6267,N_5391,N_4824);
and U6268 (N_6268,N_5003,N_5241);
nor U6269 (N_6269,N_4948,N_5082);
or U6270 (N_6270,N_5576,N_4981);
nand U6271 (N_6271,N_4974,N_5562);
xor U6272 (N_6272,N_5118,N_5443);
nor U6273 (N_6273,N_4884,N_5031);
or U6274 (N_6274,N_5375,N_5381);
and U6275 (N_6275,N_5062,N_5086);
xnor U6276 (N_6276,N_4960,N_4871);
nor U6277 (N_6277,N_5293,N_5491);
nand U6278 (N_6278,N_4883,N_5100);
nor U6279 (N_6279,N_5524,N_5464);
nor U6280 (N_6280,N_5149,N_5466);
and U6281 (N_6281,N_5355,N_5438);
nor U6282 (N_6282,N_5127,N_5213);
xnor U6283 (N_6283,N_5554,N_5151);
nand U6284 (N_6284,N_5303,N_5120);
nor U6285 (N_6285,N_4975,N_5287);
nand U6286 (N_6286,N_5314,N_5383);
and U6287 (N_6287,N_4831,N_5510);
nand U6288 (N_6288,N_5149,N_5455);
nand U6289 (N_6289,N_5158,N_5460);
xor U6290 (N_6290,N_5259,N_5507);
and U6291 (N_6291,N_5232,N_5080);
nor U6292 (N_6292,N_5421,N_5294);
and U6293 (N_6293,N_5436,N_5086);
xor U6294 (N_6294,N_5025,N_5236);
and U6295 (N_6295,N_5535,N_5332);
nand U6296 (N_6296,N_4898,N_5205);
nand U6297 (N_6297,N_5090,N_4831);
nor U6298 (N_6298,N_5397,N_4863);
nor U6299 (N_6299,N_5533,N_4965);
or U6300 (N_6300,N_4927,N_5148);
or U6301 (N_6301,N_5014,N_5534);
nor U6302 (N_6302,N_5564,N_5572);
xor U6303 (N_6303,N_5158,N_5444);
nor U6304 (N_6304,N_5100,N_5493);
and U6305 (N_6305,N_5570,N_5043);
or U6306 (N_6306,N_5561,N_5488);
xor U6307 (N_6307,N_4834,N_5045);
or U6308 (N_6308,N_4912,N_4969);
nand U6309 (N_6309,N_5247,N_5184);
and U6310 (N_6310,N_5322,N_5536);
xnor U6311 (N_6311,N_4959,N_5295);
xor U6312 (N_6312,N_4842,N_5316);
and U6313 (N_6313,N_5254,N_5407);
nand U6314 (N_6314,N_5078,N_5261);
and U6315 (N_6315,N_4991,N_4852);
and U6316 (N_6316,N_5451,N_5119);
nor U6317 (N_6317,N_5119,N_5213);
and U6318 (N_6318,N_5099,N_5115);
xnor U6319 (N_6319,N_5251,N_5529);
nand U6320 (N_6320,N_5422,N_5167);
xor U6321 (N_6321,N_5177,N_5386);
and U6322 (N_6322,N_5007,N_5475);
nand U6323 (N_6323,N_4831,N_5597);
xor U6324 (N_6324,N_5290,N_5276);
nor U6325 (N_6325,N_5161,N_4959);
xnor U6326 (N_6326,N_5238,N_5206);
nor U6327 (N_6327,N_5538,N_5589);
or U6328 (N_6328,N_4811,N_5452);
and U6329 (N_6329,N_5302,N_5277);
xor U6330 (N_6330,N_5149,N_4849);
xor U6331 (N_6331,N_4979,N_5293);
nand U6332 (N_6332,N_4916,N_5284);
xnor U6333 (N_6333,N_4821,N_4906);
nand U6334 (N_6334,N_5157,N_5346);
and U6335 (N_6335,N_4909,N_5388);
xor U6336 (N_6336,N_4900,N_4813);
xnor U6337 (N_6337,N_5368,N_5570);
or U6338 (N_6338,N_5215,N_4864);
nor U6339 (N_6339,N_5447,N_5275);
nor U6340 (N_6340,N_5078,N_4895);
nor U6341 (N_6341,N_5289,N_5191);
and U6342 (N_6342,N_4951,N_5465);
or U6343 (N_6343,N_4834,N_5020);
or U6344 (N_6344,N_5024,N_5349);
nor U6345 (N_6345,N_5445,N_5008);
nand U6346 (N_6346,N_5306,N_5109);
and U6347 (N_6347,N_4931,N_4963);
nor U6348 (N_6348,N_5426,N_5432);
nor U6349 (N_6349,N_5181,N_4866);
nand U6350 (N_6350,N_4892,N_5275);
or U6351 (N_6351,N_5380,N_5150);
nor U6352 (N_6352,N_5021,N_5127);
xnor U6353 (N_6353,N_5074,N_5041);
nand U6354 (N_6354,N_4817,N_5094);
xnor U6355 (N_6355,N_5442,N_5116);
and U6356 (N_6356,N_5171,N_5046);
nand U6357 (N_6357,N_5175,N_5122);
and U6358 (N_6358,N_5221,N_4938);
and U6359 (N_6359,N_5127,N_5532);
nor U6360 (N_6360,N_5187,N_4824);
nand U6361 (N_6361,N_4970,N_5028);
xnor U6362 (N_6362,N_5410,N_4903);
nor U6363 (N_6363,N_5345,N_4800);
nand U6364 (N_6364,N_4883,N_4901);
or U6365 (N_6365,N_5371,N_4871);
nand U6366 (N_6366,N_5015,N_5184);
nand U6367 (N_6367,N_5537,N_5157);
and U6368 (N_6368,N_5305,N_5130);
and U6369 (N_6369,N_4888,N_5423);
or U6370 (N_6370,N_5394,N_5431);
nor U6371 (N_6371,N_5369,N_4935);
or U6372 (N_6372,N_5226,N_5287);
and U6373 (N_6373,N_5483,N_4990);
xor U6374 (N_6374,N_4988,N_5439);
xor U6375 (N_6375,N_4911,N_4952);
xnor U6376 (N_6376,N_4950,N_5293);
or U6377 (N_6377,N_5281,N_4867);
nor U6378 (N_6378,N_4986,N_5164);
xnor U6379 (N_6379,N_5004,N_5049);
or U6380 (N_6380,N_4827,N_5046);
xor U6381 (N_6381,N_5393,N_5016);
or U6382 (N_6382,N_5568,N_5183);
nand U6383 (N_6383,N_5596,N_4973);
or U6384 (N_6384,N_5183,N_4904);
or U6385 (N_6385,N_5508,N_5582);
or U6386 (N_6386,N_5397,N_5524);
nand U6387 (N_6387,N_5454,N_5195);
xnor U6388 (N_6388,N_5510,N_5262);
or U6389 (N_6389,N_5252,N_5016);
nor U6390 (N_6390,N_5185,N_5564);
nor U6391 (N_6391,N_5529,N_5360);
nor U6392 (N_6392,N_4863,N_4919);
or U6393 (N_6393,N_5596,N_5187);
and U6394 (N_6394,N_5299,N_5537);
and U6395 (N_6395,N_5287,N_5386);
and U6396 (N_6396,N_5404,N_4901);
and U6397 (N_6397,N_5278,N_5515);
and U6398 (N_6398,N_4824,N_5398);
and U6399 (N_6399,N_5357,N_5566);
nor U6400 (N_6400,N_5790,N_5879);
nand U6401 (N_6401,N_5789,N_6142);
xnor U6402 (N_6402,N_6134,N_5867);
nor U6403 (N_6403,N_6206,N_6166);
and U6404 (N_6404,N_6129,N_6091);
xor U6405 (N_6405,N_5955,N_5835);
nand U6406 (N_6406,N_6309,N_6095);
nand U6407 (N_6407,N_6094,N_6261);
nand U6408 (N_6408,N_6149,N_5911);
and U6409 (N_6409,N_6375,N_5933);
nor U6410 (N_6410,N_5984,N_5767);
nor U6411 (N_6411,N_6194,N_5753);
or U6412 (N_6412,N_5854,N_5842);
and U6413 (N_6413,N_5997,N_5917);
nand U6414 (N_6414,N_6305,N_5874);
or U6415 (N_6415,N_6364,N_6037);
or U6416 (N_6416,N_6066,N_6060);
or U6417 (N_6417,N_5644,N_6225);
nand U6418 (N_6418,N_5970,N_5729);
nor U6419 (N_6419,N_5870,N_6250);
nor U6420 (N_6420,N_6077,N_6033);
xnor U6421 (N_6421,N_5849,N_5672);
nor U6422 (N_6422,N_6328,N_5732);
and U6423 (N_6423,N_5748,N_6287);
nand U6424 (N_6424,N_6004,N_5900);
nand U6425 (N_6425,N_6351,N_6269);
xor U6426 (N_6426,N_6242,N_6219);
nor U6427 (N_6427,N_6383,N_5827);
xor U6428 (N_6428,N_6034,N_5634);
nor U6429 (N_6429,N_5629,N_6127);
and U6430 (N_6430,N_6200,N_6158);
nand U6431 (N_6431,N_5905,N_5863);
and U6432 (N_6432,N_5718,N_5639);
nor U6433 (N_6433,N_6196,N_6110);
nand U6434 (N_6434,N_6378,N_6182);
and U6435 (N_6435,N_5885,N_6275);
nand U6436 (N_6436,N_6359,N_5922);
xor U6437 (N_6437,N_5944,N_5730);
and U6438 (N_6438,N_6340,N_6205);
or U6439 (N_6439,N_6162,N_6227);
or U6440 (N_6440,N_5657,N_5803);
and U6441 (N_6441,N_6363,N_6080);
nor U6442 (N_6442,N_5875,N_5702);
and U6443 (N_6443,N_6115,N_6185);
or U6444 (N_6444,N_5909,N_5707);
nand U6445 (N_6445,N_6389,N_6356);
nand U6446 (N_6446,N_5681,N_6350);
nor U6447 (N_6447,N_5719,N_6298);
nand U6448 (N_6448,N_5692,N_6308);
nand U6449 (N_6449,N_6174,N_6210);
nand U6450 (N_6450,N_6349,N_6238);
xor U6451 (N_6451,N_5979,N_5674);
and U6452 (N_6452,N_6169,N_6044);
nand U6453 (N_6453,N_5693,N_5815);
nand U6454 (N_6454,N_6140,N_5738);
and U6455 (N_6455,N_5655,N_5756);
and U6456 (N_6456,N_5614,N_6329);
or U6457 (N_6457,N_6092,N_5943);
nand U6458 (N_6458,N_5888,N_5865);
xor U6459 (N_6459,N_5628,N_5667);
nand U6460 (N_6460,N_5936,N_6118);
and U6461 (N_6461,N_5620,N_5699);
or U6462 (N_6462,N_6198,N_5828);
or U6463 (N_6463,N_5770,N_5747);
xnor U6464 (N_6464,N_5619,N_5797);
and U6465 (N_6465,N_6057,N_6161);
nor U6466 (N_6466,N_5777,N_6218);
and U6467 (N_6467,N_6214,N_5621);
nand U6468 (N_6468,N_6156,N_5873);
nor U6469 (N_6469,N_6191,N_6342);
xnor U6470 (N_6470,N_6096,N_5878);
and U6471 (N_6471,N_6252,N_5887);
nor U6472 (N_6472,N_6302,N_6143);
or U6473 (N_6473,N_5882,N_6019);
and U6474 (N_6474,N_5742,N_5973);
and U6475 (N_6475,N_5641,N_6106);
nand U6476 (N_6476,N_5959,N_6000);
or U6477 (N_6477,N_5838,N_5627);
and U6478 (N_6478,N_5662,N_6144);
and U6479 (N_6479,N_6024,N_5966);
and U6480 (N_6480,N_5953,N_6254);
nor U6481 (N_6481,N_6193,N_6015);
and U6482 (N_6482,N_6086,N_6330);
xor U6483 (N_6483,N_5688,N_5774);
or U6484 (N_6484,N_6321,N_5991);
nand U6485 (N_6485,N_5706,N_6368);
xnor U6486 (N_6486,N_6029,N_5683);
nor U6487 (N_6487,N_5811,N_5666);
or U6488 (N_6488,N_6304,N_6325);
xnor U6489 (N_6489,N_6168,N_6257);
and U6490 (N_6490,N_5763,N_5960);
nand U6491 (N_6491,N_5892,N_6105);
or U6492 (N_6492,N_6117,N_5822);
or U6493 (N_6493,N_6043,N_5847);
xor U6494 (N_6494,N_5602,N_5799);
and U6495 (N_6495,N_6195,N_6372);
and U6496 (N_6496,N_5600,N_5801);
nor U6497 (N_6497,N_6361,N_5851);
nor U6498 (N_6498,N_6175,N_6085);
nor U6499 (N_6499,N_6267,N_5798);
nand U6500 (N_6500,N_6343,N_5647);
or U6501 (N_6501,N_5890,N_5989);
or U6502 (N_6502,N_5787,N_6047);
and U6503 (N_6503,N_5834,N_6319);
nor U6504 (N_6504,N_6027,N_5603);
and U6505 (N_6505,N_6002,N_5859);
or U6506 (N_6506,N_6399,N_5745);
or U6507 (N_6507,N_6026,N_6190);
nand U6508 (N_6508,N_5894,N_5986);
nand U6509 (N_6509,N_6387,N_5935);
nor U6510 (N_6510,N_5857,N_6229);
nand U6511 (N_6511,N_5755,N_6307);
xnor U6512 (N_6512,N_6025,N_5987);
nand U6513 (N_6513,N_5845,N_6226);
nor U6514 (N_6514,N_6192,N_5677);
nand U6515 (N_6515,N_6065,N_5848);
nand U6516 (N_6516,N_6005,N_6130);
nand U6517 (N_6517,N_5924,N_5915);
or U6518 (N_6518,N_6099,N_5934);
or U6519 (N_6519,N_5823,N_5819);
or U6520 (N_6520,N_5840,N_5605);
nor U6521 (N_6521,N_6202,N_6279);
nor U6522 (N_6522,N_6067,N_6203);
and U6523 (N_6523,N_5650,N_6068);
nor U6524 (N_6524,N_5992,N_6204);
and U6525 (N_6525,N_5661,N_6069);
or U6526 (N_6526,N_6320,N_6082);
and U6527 (N_6527,N_5609,N_5687);
nor U6528 (N_6528,N_5809,N_5833);
nand U6529 (N_6529,N_5938,N_5623);
and U6530 (N_6530,N_6338,N_5947);
or U6531 (N_6531,N_5750,N_5858);
and U6532 (N_6532,N_6197,N_6014);
xor U6533 (N_6533,N_6377,N_6113);
xnor U6534 (N_6534,N_5717,N_5994);
xor U6535 (N_6535,N_6285,N_5678);
nor U6536 (N_6536,N_5949,N_5923);
nor U6537 (N_6537,N_5784,N_5685);
nand U6538 (N_6538,N_5700,N_6051);
xor U6539 (N_6539,N_6098,N_6295);
and U6540 (N_6540,N_5780,N_6097);
nand U6541 (N_6541,N_6052,N_5733);
nand U6542 (N_6542,N_5788,N_5932);
xor U6543 (N_6543,N_6394,N_5910);
xnor U6544 (N_6544,N_6048,N_6055);
nand U6545 (N_6545,N_5794,N_5637);
nand U6546 (N_6546,N_5734,N_6331);
nand U6547 (N_6547,N_6126,N_6186);
xor U6548 (N_6548,N_5804,N_5843);
nand U6549 (N_6549,N_5715,N_6102);
or U6550 (N_6550,N_6036,N_6222);
nor U6551 (N_6551,N_6132,N_5826);
xnor U6552 (N_6552,N_6266,N_6259);
and U6553 (N_6553,N_5613,N_6012);
nand U6554 (N_6554,N_5829,N_5975);
or U6555 (N_6555,N_6178,N_6180);
or U6556 (N_6556,N_5704,N_5744);
or U6557 (N_6557,N_5972,N_6274);
and U6558 (N_6558,N_6201,N_6396);
or U6559 (N_6559,N_5886,N_5956);
and U6560 (N_6560,N_5864,N_6018);
nor U6561 (N_6561,N_5649,N_6327);
and U6562 (N_6562,N_6016,N_6154);
or U6563 (N_6563,N_5836,N_6299);
nand U6564 (N_6564,N_6059,N_6114);
nor U6565 (N_6565,N_6217,N_6253);
xor U6566 (N_6566,N_6112,N_5682);
nor U6567 (N_6567,N_6141,N_6355);
xor U6568 (N_6568,N_5844,N_5711);
nor U6569 (N_6569,N_6138,N_5645);
nand U6570 (N_6570,N_6173,N_5726);
and U6571 (N_6571,N_6021,N_6151);
or U6572 (N_6572,N_5813,N_5807);
and U6573 (N_6573,N_6075,N_5850);
nor U6574 (N_6574,N_6146,N_6341);
and U6575 (N_6575,N_5725,N_6301);
nor U6576 (N_6576,N_6353,N_6076);
nor U6577 (N_6577,N_6345,N_5679);
xor U6578 (N_6578,N_6334,N_6376);
nand U6579 (N_6579,N_6256,N_5861);
nor U6580 (N_6580,N_6346,N_6392);
and U6581 (N_6581,N_5775,N_6365);
nand U6582 (N_6582,N_6211,N_5806);
nor U6583 (N_6583,N_6040,N_6183);
and U6584 (N_6584,N_5980,N_6172);
xor U6585 (N_6585,N_6153,N_6170);
or U6586 (N_6586,N_6122,N_6271);
xnor U6587 (N_6587,N_6073,N_6234);
nand U6588 (N_6588,N_6381,N_6006);
nand U6589 (N_6589,N_6049,N_6288);
nand U6590 (N_6590,N_5724,N_6103);
or U6591 (N_6591,N_6312,N_6313);
nand U6592 (N_6592,N_6088,N_5893);
nand U6593 (N_6593,N_6171,N_6030);
or U6594 (N_6594,N_5786,N_6282);
and U6595 (N_6595,N_6317,N_5976);
and U6596 (N_6596,N_6101,N_5872);
or U6597 (N_6597,N_5746,N_5721);
xnor U6598 (N_6598,N_5999,N_6137);
nand U6599 (N_6599,N_5884,N_6042);
nand U6600 (N_6600,N_5630,N_6239);
xor U6601 (N_6601,N_6354,N_6022);
nand U6602 (N_6602,N_5772,N_5761);
or U6603 (N_6603,N_5760,N_6270);
nand U6604 (N_6604,N_5927,N_6155);
nor U6605 (N_6605,N_6284,N_5610);
and U6606 (N_6606,N_6293,N_5633);
xor U6607 (N_6607,N_5957,N_6380);
xor U6608 (N_6608,N_6181,N_5652);
nand U6609 (N_6609,N_6243,N_6221);
and U6610 (N_6610,N_6236,N_5824);
nor U6611 (N_6611,N_5616,N_5624);
nand U6612 (N_6612,N_6045,N_6324);
nor U6613 (N_6613,N_5812,N_6072);
or U6614 (N_6614,N_6276,N_6007);
nor U6615 (N_6615,N_5686,N_5963);
xor U6616 (N_6616,N_6344,N_6316);
xnor U6617 (N_6617,N_5995,N_5846);
nand U6618 (N_6618,N_5769,N_5877);
or U6619 (N_6619,N_6120,N_6001);
xor U6620 (N_6620,N_5684,N_6286);
and U6621 (N_6621,N_5902,N_5622);
nor U6622 (N_6622,N_6011,N_5618);
or U6623 (N_6623,N_6337,N_6318);
xnor U6624 (N_6624,N_5825,N_5871);
or U6625 (N_6625,N_5940,N_5920);
and U6626 (N_6626,N_5810,N_6209);
nand U6627 (N_6627,N_5856,N_5795);
xnor U6628 (N_6628,N_6152,N_5898);
nor U6629 (N_6629,N_5907,N_6220);
nor U6630 (N_6630,N_6028,N_5971);
nand U6631 (N_6631,N_5611,N_6207);
and U6632 (N_6632,N_6031,N_5728);
or U6633 (N_6633,N_5658,N_6233);
and U6634 (N_6634,N_5626,N_6306);
and U6635 (N_6635,N_5896,N_6136);
nand U6636 (N_6636,N_6291,N_5705);
or U6637 (N_6637,N_6335,N_6083);
nand U6638 (N_6638,N_5939,N_5654);
or U6639 (N_6639,N_5855,N_6184);
nor U6640 (N_6640,N_5671,N_6164);
and U6641 (N_6641,N_6241,N_6213);
xnor U6642 (N_6642,N_6148,N_6362);
nor U6643 (N_6643,N_5749,N_5759);
and U6644 (N_6644,N_5740,N_6109);
nand U6645 (N_6645,N_6089,N_5736);
and U6646 (N_6646,N_5831,N_5821);
or U6647 (N_6647,N_6260,N_5876);
nand U6648 (N_6648,N_5779,N_6315);
nor U6649 (N_6649,N_5914,N_5636);
nor U6650 (N_6650,N_5737,N_6003);
nand U6651 (N_6651,N_6246,N_5903);
xnor U6652 (N_6652,N_6216,N_5768);
and U6653 (N_6653,N_6056,N_6009);
nor U6654 (N_6654,N_6145,N_6251);
nand U6655 (N_6655,N_6087,N_6093);
xor U6656 (N_6656,N_5974,N_5830);
xor U6657 (N_6657,N_5778,N_5659);
nor U6658 (N_6658,N_5978,N_6133);
nor U6659 (N_6659,N_6123,N_5703);
xor U6660 (N_6660,N_5642,N_6157);
xnor U6661 (N_6661,N_5928,N_6303);
and U6662 (N_6662,N_5670,N_5723);
and U6663 (N_6663,N_6119,N_6074);
xor U6664 (N_6664,N_5814,N_6081);
and U6665 (N_6665,N_6063,N_5739);
nor U6666 (N_6666,N_5766,N_6326);
and U6667 (N_6667,N_5818,N_6053);
nor U6668 (N_6668,N_6071,N_6023);
xor U6669 (N_6669,N_6188,N_5757);
or U6670 (N_6670,N_6248,N_5607);
nand U6671 (N_6671,N_6244,N_6121);
or U6672 (N_6672,N_5841,N_5697);
xnor U6673 (N_6673,N_6189,N_5996);
and U6674 (N_6674,N_5612,N_5709);
nor U6675 (N_6675,N_5817,N_5802);
nand U6676 (N_6676,N_6310,N_5752);
nand U6677 (N_6677,N_6300,N_6061);
nor U6678 (N_6678,N_5908,N_5983);
and U6679 (N_6679,N_5977,N_5839);
xor U6680 (N_6680,N_5990,N_6369);
or U6681 (N_6681,N_5796,N_5668);
xnor U6682 (N_6682,N_5866,N_5837);
xor U6683 (N_6683,N_6078,N_6358);
and U6684 (N_6684,N_6391,N_5656);
and U6685 (N_6685,N_6176,N_6323);
and U6686 (N_6686,N_5773,N_6084);
nand U6687 (N_6687,N_5741,N_5781);
and U6688 (N_6688,N_5853,N_6371);
xnor U6689 (N_6689,N_6263,N_6124);
and U6690 (N_6690,N_5921,N_5988);
or U6691 (N_6691,N_5604,N_6070);
or U6692 (N_6692,N_5716,N_6289);
or U6693 (N_6693,N_5690,N_5950);
or U6694 (N_6694,N_6167,N_5664);
or U6695 (N_6695,N_5793,N_5860);
nand U6696 (N_6696,N_5925,N_5808);
nor U6697 (N_6697,N_5660,N_6100);
and U6698 (N_6698,N_5648,N_6264);
and U6699 (N_6699,N_5676,N_5862);
nor U6700 (N_6700,N_5695,N_5751);
nand U6701 (N_6701,N_6273,N_6224);
nand U6702 (N_6702,N_6357,N_5899);
and U6703 (N_6703,N_6296,N_6322);
and U6704 (N_6704,N_5651,N_5820);
nor U6705 (N_6705,N_6366,N_5930);
nand U6706 (N_6706,N_5880,N_6360);
nand U6707 (N_6707,N_5635,N_5783);
or U6708 (N_6708,N_6008,N_5954);
xnor U6709 (N_6709,N_6339,N_5919);
nor U6710 (N_6710,N_5743,N_6297);
xor U6711 (N_6711,N_5805,N_5881);
nand U6712 (N_6712,N_6032,N_5631);
xnor U6713 (N_6713,N_5640,N_6179);
nor U6714 (N_6714,N_5722,N_6163);
and U6715 (N_6715,N_6290,N_5852);
nand U6716 (N_6716,N_6232,N_6107);
nand U6717 (N_6717,N_5771,N_5969);
nor U6718 (N_6718,N_6013,N_5913);
or U6719 (N_6719,N_5653,N_6332);
or U6720 (N_6720,N_6373,N_6393);
nand U6721 (N_6721,N_6277,N_5929);
xor U6722 (N_6722,N_5776,N_5632);
nor U6723 (N_6723,N_6041,N_5958);
nor U6724 (N_6724,N_5952,N_6054);
nor U6725 (N_6725,N_5764,N_5696);
nand U6726 (N_6726,N_5961,N_5720);
nand U6727 (N_6727,N_6386,N_6079);
nor U6728 (N_6728,N_6294,N_6017);
nand U6729 (N_6729,N_6398,N_5762);
nand U6730 (N_6730,N_6046,N_5918);
or U6731 (N_6731,N_5912,N_6020);
nand U6732 (N_6732,N_6265,N_6379);
nor U6733 (N_6733,N_5646,N_6352);
nand U6734 (N_6734,N_6116,N_5982);
nand U6735 (N_6735,N_6311,N_5617);
nand U6736 (N_6736,N_5889,N_5869);
xnor U6737 (N_6737,N_6397,N_5964);
xor U6738 (N_6738,N_6160,N_5985);
nand U6739 (N_6739,N_6384,N_5663);
xor U6740 (N_6740,N_5937,N_6038);
and U6741 (N_6741,N_5669,N_5800);
xor U6742 (N_6742,N_5608,N_6131);
xor U6743 (N_6743,N_6139,N_6108);
and U6744 (N_6744,N_6268,N_5791);
or U6745 (N_6745,N_6228,N_6231);
and U6746 (N_6746,N_6150,N_6262);
nand U6747 (N_6747,N_5868,N_5816);
nor U6748 (N_6748,N_6235,N_6064);
nand U6749 (N_6749,N_5951,N_6128);
nor U6750 (N_6750,N_6388,N_5965);
xnor U6751 (N_6751,N_6104,N_6336);
and U6752 (N_6752,N_5832,N_6278);
xor U6753 (N_6753,N_6230,N_6208);
and U6754 (N_6754,N_5946,N_5689);
nand U6755 (N_6755,N_5714,N_5948);
nor U6756 (N_6756,N_5731,N_6050);
nand U6757 (N_6757,N_6215,N_6280);
xor U6758 (N_6758,N_6135,N_6283);
nor U6759 (N_6759,N_5916,N_5785);
xnor U6760 (N_6760,N_5665,N_6223);
or U6761 (N_6761,N_5981,N_6247);
or U6762 (N_6762,N_6385,N_5883);
nand U6763 (N_6763,N_5792,N_6010);
nand U6764 (N_6764,N_6111,N_5713);
nand U6765 (N_6765,N_6199,N_5942);
nor U6766 (N_6766,N_5993,N_5615);
or U6767 (N_6767,N_5673,N_5891);
nand U6768 (N_6768,N_6390,N_6090);
and U6769 (N_6769,N_6258,N_5708);
or U6770 (N_6770,N_5962,N_6314);
or U6771 (N_6771,N_5754,N_6177);
nand U6772 (N_6772,N_5901,N_5698);
or U6773 (N_6773,N_5643,N_6367);
xor U6774 (N_6774,N_5727,N_5710);
nand U6775 (N_6775,N_6347,N_5941);
and U6776 (N_6776,N_6272,N_5967);
or U6777 (N_6777,N_5625,N_5895);
xor U6778 (N_6778,N_6348,N_5758);
and U6779 (N_6779,N_6255,N_5712);
nand U6780 (N_6780,N_6187,N_5926);
nor U6781 (N_6781,N_6058,N_6240);
xnor U6782 (N_6782,N_6370,N_6159);
and U6783 (N_6783,N_5765,N_6147);
and U6784 (N_6784,N_5601,N_6245);
nand U6785 (N_6785,N_5638,N_5694);
xor U6786 (N_6786,N_5998,N_6249);
nand U6787 (N_6787,N_6035,N_6125);
or U6788 (N_6788,N_5968,N_6395);
or U6789 (N_6789,N_6333,N_6212);
and U6790 (N_6790,N_6281,N_5906);
or U6791 (N_6791,N_6237,N_5782);
and U6792 (N_6792,N_6039,N_5606);
or U6793 (N_6793,N_5691,N_5897);
nor U6794 (N_6794,N_6062,N_5735);
or U6795 (N_6795,N_5931,N_6374);
or U6796 (N_6796,N_5945,N_5904);
nand U6797 (N_6797,N_6382,N_5680);
nor U6798 (N_6798,N_5675,N_6292);
xor U6799 (N_6799,N_5701,N_6165);
or U6800 (N_6800,N_6214,N_6316);
nor U6801 (N_6801,N_5857,N_6239);
nor U6802 (N_6802,N_5786,N_6092);
and U6803 (N_6803,N_6374,N_6019);
and U6804 (N_6804,N_6157,N_5640);
nor U6805 (N_6805,N_5788,N_6153);
nor U6806 (N_6806,N_6239,N_5749);
xor U6807 (N_6807,N_5785,N_6346);
nor U6808 (N_6808,N_5730,N_5722);
nor U6809 (N_6809,N_6067,N_5985);
nor U6810 (N_6810,N_6316,N_5725);
or U6811 (N_6811,N_5903,N_6114);
and U6812 (N_6812,N_5659,N_5803);
nor U6813 (N_6813,N_6055,N_6306);
nor U6814 (N_6814,N_6185,N_6313);
and U6815 (N_6815,N_6317,N_6328);
nor U6816 (N_6816,N_5714,N_6365);
or U6817 (N_6817,N_5701,N_5806);
nor U6818 (N_6818,N_6200,N_5617);
or U6819 (N_6819,N_5714,N_6163);
and U6820 (N_6820,N_5972,N_5708);
nor U6821 (N_6821,N_5764,N_5761);
nand U6822 (N_6822,N_6395,N_6045);
nor U6823 (N_6823,N_5902,N_6021);
nor U6824 (N_6824,N_5850,N_6002);
nor U6825 (N_6825,N_6129,N_5738);
and U6826 (N_6826,N_5894,N_6303);
xor U6827 (N_6827,N_6391,N_6331);
nor U6828 (N_6828,N_6042,N_5655);
nand U6829 (N_6829,N_6388,N_5835);
and U6830 (N_6830,N_6121,N_6027);
nand U6831 (N_6831,N_6139,N_5996);
nor U6832 (N_6832,N_6276,N_5686);
nand U6833 (N_6833,N_6125,N_6054);
and U6834 (N_6834,N_6265,N_5913);
xnor U6835 (N_6835,N_5626,N_6213);
and U6836 (N_6836,N_6268,N_6261);
xnor U6837 (N_6837,N_6054,N_6000);
and U6838 (N_6838,N_6011,N_5934);
nor U6839 (N_6839,N_6154,N_6162);
and U6840 (N_6840,N_6255,N_6163);
nor U6841 (N_6841,N_5860,N_5835);
and U6842 (N_6842,N_6356,N_6050);
nand U6843 (N_6843,N_6041,N_5961);
xnor U6844 (N_6844,N_6182,N_5642);
or U6845 (N_6845,N_5625,N_5934);
and U6846 (N_6846,N_6315,N_6076);
nor U6847 (N_6847,N_6121,N_5615);
xor U6848 (N_6848,N_5937,N_6080);
or U6849 (N_6849,N_5607,N_5738);
xnor U6850 (N_6850,N_6251,N_6282);
and U6851 (N_6851,N_5887,N_6182);
and U6852 (N_6852,N_5770,N_5852);
xor U6853 (N_6853,N_6198,N_5714);
nor U6854 (N_6854,N_6358,N_6176);
nand U6855 (N_6855,N_5661,N_5637);
nand U6856 (N_6856,N_5813,N_5947);
or U6857 (N_6857,N_5933,N_5873);
xor U6858 (N_6858,N_5790,N_6196);
and U6859 (N_6859,N_6287,N_6358);
nand U6860 (N_6860,N_6186,N_6289);
xor U6861 (N_6861,N_6168,N_6236);
nand U6862 (N_6862,N_5607,N_5736);
and U6863 (N_6863,N_5845,N_6121);
nor U6864 (N_6864,N_6176,N_6353);
nor U6865 (N_6865,N_5873,N_5686);
xor U6866 (N_6866,N_5842,N_6138);
xnor U6867 (N_6867,N_6183,N_6369);
nand U6868 (N_6868,N_6127,N_5785);
or U6869 (N_6869,N_5975,N_5885);
and U6870 (N_6870,N_6005,N_5783);
or U6871 (N_6871,N_6277,N_6261);
nor U6872 (N_6872,N_5662,N_6363);
and U6873 (N_6873,N_6367,N_6317);
xnor U6874 (N_6874,N_5723,N_5870);
nor U6875 (N_6875,N_5772,N_5675);
and U6876 (N_6876,N_6265,N_5988);
or U6877 (N_6877,N_5940,N_6167);
nor U6878 (N_6878,N_5801,N_5776);
xnor U6879 (N_6879,N_5622,N_5830);
nor U6880 (N_6880,N_6311,N_5830);
or U6881 (N_6881,N_5733,N_5902);
xnor U6882 (N_6882,N_6291,N_5972);
xnor U6883 (N_6883,N_6023,N_5835);
xnor U6884 (N_6884,N_5614,N_6209);
or U6885 (N_6885,N_5801,N_5637);
xnor U6886 (N_6886,N_5656,N_5649);
or U6887 (N_6887,N_5819,N_6284);
or U6888 (N_6888,N_5614,N_6061);
xor U6889 (N_6889,N_6086,N_6009);
xor U6890 (N_6890,N_6311,N_6324);
and U6891 (N_6891,N_6056,N_6222);
xnor U6892 (N_6892,N_6324,N_5622);
or U6893 (N_6893,N_6138,N_5824);
xor U6894 (N_6894,N_6056,N_6066);
or U6895 (N_6895,N_5611,N_6340);
and U6896 (N_6896,N_6138,N_5919);
nor U6897 (N_6897,N_6214,N_6174);
nand U6898 (N_6898,N_5864,N_5795);
nor U6899 (N_6899,N_5989,N_6300);
xor U6900 (N_6900,N_5851,N_6258);
xor U6901 (N_6901,N_6248,N_5935);
nor U6902 (N_6902,N_6194,N_6256);
and U6903 (N_6903,N_6107,N_5837);
xnor U6904 (N_6904,N_6299,N_5766);
or U6905 (N_6905,N_5791,N_6224);
and U6906 (N_6906,N_6333,N_6158);
and U6907 (N_6907,N_5848,N_6036);
nand U6908 (N_6908,N_5967,N_6105);
xor U6909 (N_6909,N_6032,N_6370);
or U6910 (N_6910,N_5846,N_6284);
xor U6911 (N_6911,N_6367,N_5624);
xnor U6912 (N_6912,N_5876,N_5974);
or U6913 (N_6913,N_5862,N_6167);
nand U6914 (N_6914,N_6097,N_6316);
nand U6915 (N_6915,N_5655,N_6393);
nand U6916 (N_6916,N_6171,N_5618);
nor U6917 (N_6917,N_5702,N_5880);
and U6918 (N_6918,N_6353,N_5795);
or U6919 (N_6919,N_5969,N_5719);
nand U6920 (N_6920,N_6066,N_6063);
xor U6921 (N_6921,N_5732,N_5883);
and U6922 (N_6922,N_6238,N_6105);
nand U6923 (N_6923,N_6184,N_6268);
nand U6924 (N_6924,N_5819,N_5609);
nand U6925 (N_6925,N_5707,N_5736);
xor U6926 (N_6926,N_6110,N_6208);
xor U6927 (N_6927,N_6293,N_6184);
and U6928 (N_6928,N_6299,N_6357);
and U6929 (N_6929,N_6075,N_6317);
nand U6930 (N_6930,N_6008,N_5904);
xnor U6931 (N_6931,N_5727,N_5834);
or U6932 (N_6932,N_5947,N_5778);
or U6933 (N_6933,N_6368,N_5715);
nor U6934 (N_6934,N_6177,N_6192);
nor U6935 (N_6935,N_6317,N_6103);
xor U6936 (N_6936,N_5731,N_6356);
nor U6937 (N_6937,N_5775,N_5872);
nand U6938 (N_6938,N_5900,N_6373);
or U6939 (N_6939,N_6163,N_5791);
and U6940 (N_6940,N_6320,N_6078);
nand U6941 (N_6941,N_6072,N_5973);
and U6942 (N_6942,N_6393,N_5776);
xnor U6943 (N_6943,N_6166,N_5777);
or U6944 (N_6944,N_6056,N_6341);
xor U6945 (N_6945,N_5631,N_5617);
or U6946 (N_6946,N_6204,N_6049);
and U6947 (N_6947,N_6263,N_6187);
nor U6948 (N_6948,N_5858,N_6230);
nor U6949 (N_6949,N_6035,N_6095);
nor U6950 (N_6950,N_6306,N_6121);
or U6951 (N_6951,N_5864,N_6176);
xnor U6952 (N_6952,N_5859,N_6347);
nand U6953 (N_6953,N_6383,N_6041);
xor U6954 (N_6954,N_6397,N_6003);
nand U6955 (N_6955,N_6023,N_6167);
or U6956 (N_6956,N_6247,N_6126);
or U6957 (N_6957,N_5650,N_5945);
nand U6958 (N_6958,N_5819,N_6380);
nor U6959 (N_6959,N_5974,N_6148);
xor U6960 (N_6960,N_6148,N_5894);
xnor U6961 (N_6961,N_6185,N_5631);
and U6962 (N_6962,N_6159,N_5979);
or U6963 (N_6963,N_6021,N_5613);
or U6964 (N_6964,N_6170,N_5708);
nor U6965 (N_6965,N_6017,N_5987);
and U6966 (N_6966,N_5630,N_6286);
xnor U6967 (N_6967,N_6122,N_6061);
or U6968 (N_6968,N_5671,N_5696);
or U6969 (N_6969,N_6054,N_5654);
nor U6970 (N_6970,N_6151,N_6169);
nand U6971 (N_6971,N_5730,N_6068);
xor U6972 (N_6972,N_5890,N_6001);
or U6973 (N_6973,N_5909,N_5977);
nand U6974 (N_6974,N_5792,N_6170);
xnor U6975 (N_6975,N_5813,N_5698);
nor U6976 (N_6976,N_6115,N_5796);
and U6977 (N_6977,N_6349,N_6034);
nand U6978 (N_6978,N_6266,N_5969);
nor U6979 (N_6979,N_5904,N_5851);
or U6980 (N_6980,N_5821,N_6053);
or U6981 (N_6981,N_6079,N_6223);
nor U6982 (N_6982,N_5709,N_5851);
nor U6983 (N_6983,N_6263,N_5811);
or U6984 (N_6984,N_6065,N_5919);
xor U6985 (N_6985,N_6156,N_6335);
nand U6986 (N_6986,N_5738,N_6200);
or U6987 (N_6987,N_6375,N_6366);
xnor U6988 (N_6988,N_6386,N_5757);
or U6989 (N_6989,N_6290,N_5700);
and U6990 (N_6990,N_6072,N_6112);
nand U6991 (N_6991,N_5644,N_5613);
nor U6992 (N_6992,N_6037,N_6132);
nand U6993 (N_6993,N_6123,N_6040);
xor U6994 (N_6994,N_6026,N_5985);
xnor U6995 (N_6995,N_6323,N_5922);
and U6996 (N_6996,N_5715,N_6114);
or U6997 (N_6997,N_6097,N_6295);
nor U6998 (N_6998,N_5706,N_5886);
nor U6999 (N_6999,N_6181,N_6015);
xnor U7000 (N_7000,N_6022,N_6015);
and U7001 (N_7001,N_5803,N_6054);
or U7002 (N_7002,N_6369,N_6127);
and U7003 (N_7003,N_6017,N_5681);
and U7004 (N_7004,N_6061,N_5702);
or U7005 (N_7005,N_5928,N_5878);
and U7006 (N_7006,N_5657,N_5810);
xnor U7007 (N_7007,N_5961,N_6165);
or U7008 (N_7008,N_6241,N_6287);
nor U7009 (N_7009,N_6245,N_5605);
nor U7010 (N_7010,N_6368,N_6392);
and U7011 (N_7011,N_5637,N_5902);
and U7012 (N_7012,N_5852,N_5855);
nand U7013 (N_7013,N_6310,N_5913);
or U7014 (N_7014,N_6374,N_5731);
nand U7015 (N_7015,N_5966,N_6330);
nand U7016 (N_7016,N_6133,N_5879);
or U7017 (N_7017,N_5782,N_6069);
xor U7018 (N_7018,N_6359,N_6176);
or U7019 (N_7019,N_6350,N_5738);
and U7020 (N_7020,N_5649,N_6050);
nor U7021 (N_7021,N_6150,N_5897);
xor U7022 (N_7022,N_6045,N_6115);
and U7023 (N_7023,N_5895,N_6230);
xnor U7024 (N_7024,N_6175,N_5798);
and U7025 (N_7025,N_5783,N_5819);
and U7026 (N_7026,N_5699,N_5778);
xnor U7027 (N_7027,N_6247,N_6318);
nor U7028 (N_7028,N_6305,N_5853);
nand U7029 (N_7029,N_5642,N_6380);
or U7030 (N_7030,N_5940,N_6014);
and U7031 (N_7031,N_5808,N_6120);
nor U7032 (N_7032,N_5939,N_6236);
xnor U7033 (N_7033,N_5850,N_6276);
or U7034 (N_7034,N_6286,N_6193);
and U7035 (N_7035,N_5980,N_5789);
xnor U7036 (N_7036,N_6031,N_6157);
and U7037 (N_7037,N_5841,N_5801);
or U7038 (N_7038,N_5696,N_6081);
nor U7039 (N_7039,N_6317,N_6206);
or U7040 (N_7040,N_5707,N_5678);
nor U7041 (N_7041,N_6072,N_6373);
and U7042 (N_7042,N_6205,N_5763);
nor U7043 (N_7043,N_6382,N_6398);
nor U7044 (N_7044,N_6333,N_5667);
nor U7045 (N_7045,N_5769,N_6338);
xnor U7046 (N_7046,N_6029,N_6353);
xnor U7047 (N_7047,N_5761,N_5742);
nand U7048 (N_7048,N_6359,N_6053);
xor U7049 (N_7049,N_6303,N_6108);
xor U7050 (N_7050,N_5620,N_6190);
nand U7051 (N_7051,N_5683,N_6298);
xnor U7052 (N_7052,N_5707,N_6159);
nor U7053 (N_7053,N_5910,N_5947);
xnor U7054 (N_7054,N_6304,N_6056);
and U7055 (N_7055,N_6048,N_5881);
or U7056 (N_7056,N_6161,N_5814);
and U7057 (N_7057,N_5843,N_6230);
and U7058 (N_7058,N_6266,N_5989);
nor U7059 (N_7059,N_5840,N_5942);
nand U7060 (N_7060,N_6282,N_6227);
xor U7061 (N_7061,N_5689,N_6312);
or U7062 (N_7062,N_5998,N_5652);
nand U7063 (N_7063,N_5691,N_5724);
nor U7064 (N_7064,N_5981,N_5785);
xor U7065 (N_7065,N_5672,N_5779);
nor U7066 (N_7066,N_5641,N_5857);
nor U7067 (N_7067,N_5730,N_5715);
xor U7068 (N_7068,N_6259,N_6319);
or U7069 (N_7069,N_6085,N_5728);
nand U7070 (N_7070,N_5878,N_6078);
xnor U7071 (N_7071,N_6038,N_5685);
xnor U7072 (N_7072,N_6176,N_6264);
xor U7073 (N_7073,N_6343,N_6129);
or U7074 (N_7074,N_6078,N_5775);
nand U7075 (N_7075,N_5649,N_5739);
nor U7076 (N_7076,N_6257,N_6261);
and U7077 (N_7077,N_6160,N_5818);
nor U7078 (N_7078,N_6234,N_5888);
xor U7079 (N_7079,N_5967,N_6176);
nand U7080 (N_7080,N_5616,N_5878);
or U7081 (N_7081,N_5790,N_6009);
nand U7082 (N_7082,N_6130,N_5800);
nor U7083 (N_7083,N_5709,N_5686);
or U7084 (N_7084,N_5954,N_6027);
xnor U7085 (N_7085,N_6347,N_5669);
nand U7086 (N_7086,N_6194,N_6336);
xnor U7087 (N_7087,N_5641,N_6293);
or U7088 (N_7088,N_6307,N_6231);
and U7089 (N_7089,N_6320,N_5674);
nor U7090 (N_7090,N_5936,N_6093);
nand U7091 (N_7091,N_6103,N_5892);
xnor U7092 (N_7092,N_5918,N_5730);
nand U7093 (N_7093,N_6196,N_5680);
or U7094 (N_7094,N_6304,N_6039);
nor U7095 (N_7095,N_6025,N_5827);
and U7096 (N_7096,N_5924,N_5606);
and U7097 (N_7097,N_5629,N_6285);
nand U7098 (N_7098,N_5808,N_5611);
or U7099 (N_7099,N_6157,N_6385);
xnor U7100 (N_7100,N_5688,N_5679);
and U7101 (N_7101,N_5899,N_6366);
nand U7102 (N_7102,N_6112,N_5928);
nand U7103 (N_7103,N_5619,N_6226);
xnor U7104 (N_7104,N_6391,N_6330);
and U7105 (N_7105,N_6051,N_5718);
nor U7106 (N_7106,N_6028,N_5619);
and U7107 (N_7107,N_5822,N_6192);
nor U7108 (N_7108,N_6177,N_5955);
or U7109 (N_7109,N_6044,N_6062);
nand U7110 (N_7110,N_6121,N_5867);
xnor U7111 (N_7111,N_5890,N_5686);
nor U7112 (N_7112,N_5812,N_5837);
nand U7113 (N_7113,N_6216,N_5647);
xor U7114 (N_7114,N_5661,N_5819);
or U7115 (N_7115,N_6245,N_6164);
and U7116 (N_7116,N_6378,N_5817);
or U7117 (N_7117,N_5659,N_5776);
or U7118 (N_7118,N_5824,N_5654);
nand U7119 (N_7119,N_6358,N_6128);
xor U7120 (N_7120,N_6314,N_5699);
nor U7121 (N_7121,N_6080,N_5728);
nor U7122 (N_7122,N_5790,N_5665);
or U7123 (N_7123,N_6173,N_5800);
xor U7124 (N_7124,N_6179,N_5873);
xnor U7125 (N_7125,N_6264,N_5780);
and U7126 (N_7126,N_6272,N_5822);
xor U7127 (N_7127,N_5943,N_6126);
nor U7128 (N_7128,N_5846,N_6297);
nand U7129 (N_7129,N_6246,N_5623);
xnor U7130 (N_7130,N_5933,N_5717);
nand U7131 (N_7131,N_6286,N_6091);
and U7132 (N_7132,N_6194,N_6352);
xor U7133 (N_7133,N_5858,N_5726);
and U7134 (N_7134,N_6252,N_5641);
and U7135 (N_7135,N_6240,N_6018);
and U7136 (N_7136,N_6053,N_5781);
or U7137 (N_7137,N_5677,N_5878);
nor U7138 (N_7138,N_6312,N_5676);
nor U7139 (N_7139,N_5981,N_5824);
xnor U7140 (N_7140,N_5762,N_6117);
nor U7141 (N_7141,N_5799,N_6049);
xnor U7142 (N_7142,N_6014,N_6124);
or U7143 (N_7143,N_6104,N_6319);
nor U7144 (N_7144,N_6050,N_6034);
nor U7145 (N_7145,N_6164,N_6066);
nand U7146 (N_7146,N_6127,N_6394);
and U7147 (N_7147,N_5889,N_6279);
and U7148 (N_7148,N_6001,N_5758);
nand U7149 (N_7149,N_5642,N_6387);
nand U7150 (N_7150,N_5897,N_6372);
nor U7151 (N_7151,N_6117,N_5698);
and U7152 (N_7152,N_6014,N_5817);
nor U7153 (N_7153,N_6262,N_6230);
and U7154 (N_7154,N_6280,N_5779);
nand U7155 (N_7155,N_6360,N_5643);
xnor U7156 (N_7156,N_5686,N_6271);
or U7157 (N_7157,N_5988,N_6376);
xnor U7158 (N_7158,N_5972,N_6282);
and U7159 (N_7159,N_5818,N_5759);
or U7160 (N_7160,N_5721,N_5635);
nand U7161 (N_7161,N_5822,N_6374);
and U7162 (N_7162,N_5654,N_6358);
xor U7163 (N_7163,N_6315,N_5932);
and U7164 (N_7164,N_6149,N_5733);
nor U7165 (N_7165,N_6220,N_6085);
nor U7166 (N_7166,N_5949,N_5708);
nand U7167 (N_7167,N_5715,N_5816);
and U7168 (N_7168,N_6175,N_5662);
nor U7169 (N_7169,N_5781,N_5827);
and U7170 (N_7170,N_6115,N_6266);
nand U7171 (N_7171,N_6319,N_6039);
or U7172 (N_7172,N_5749,N_5725);
or U7173 (N_7173,N_6226,N_6106);
and U7174 (N_7174,N_5880,N_5718);
nor U7175 (N_7175,N_6169,N_6085);
nand U7176 (N_7176,N_5920,N_5958);
and U7177 (N_7177,N_6270,N_6096);
or U7178 (N_7178,N_5949,N_5630);
xnor U7179 (N_7179,N_6180,N_6207);
nor U7180 (N_7180,N_5846,N_5789);
xnor U7181 (N_7181,N_5710,N_6020);
and U7182 (N_7182,N_5949,N_5835);
and U7183 (N_7183,N_6113,N_6227);
nor U7184 (N_7184,N_5924,N_6310);
and U7185 (N_7185,N_6085,N_6289);
xnor U7186 (N_7186,N_6393,N_6199);
nor U7187 (N_7187,N_5813,N_6082);
nand U7188 (N_7188,N_6208,N_5724);
and U7189 (N_7189,N_5969,N_5925);
xnor U7190 (N_7190,N_6056,N_5734);
nand U7191 (N_7191,N_6363,N_6258);
xor U7192 (N_7192,N_5841,N_5716);
nor U7193 (N_7193,N_6146,N_6322);
nand U7194 (N_7194,N_5713,N_6214);
and U7195 (N_7195,N_6026,N_5866);
and U7196 (N_7196,N_6144,N_6239);
and U7197 (N_7197,N_5999,N_6013);
and U7198 (N_7198,N_6058,N_6303);
or U7199 (N_7199,N_5791,N_6006);
nor U7200 (N_7200,N_6706,N_6496);
or U7201 (N_7201,N_6471,N_6410);
xnor U7202 (N_7202,N_6563,N_6890);
or U7203 (N_7203,N_6949,N_6577);
and U7204 (N_7204,N_6963,N_6925);
xor U7205 (N_7205,N_6919,N_7107);
and U7206 (N_7206,N_7070,N_6809);
xnor U7207 (N_7207,N_6710,N_6435);
xor U7208 (N_7208,N_6585,N_6802);
nor U7209 (N_7209,N_6443,N_7145);
nor U7210 (N_7210,N_7039,N_6836);
and U7211 (N_7211,N_6812,N_6634);
xor U7212 (N_7212,N_6436,N_7061);
and U7213 (N_7213,N_7040,N_6954);
xor U7214 (N_7214,N_6827,N_6484);
or U7215 (N_7215,N_6854,N_7105);
or U7216 (N_7216,N_7155,N_6975);
and U7217 (N_7217,N_7158,N_6842);
and U7218 (N_7218,N_6520,N_7035);
xnor U7219 (N_7219,N_6796,N_6625);
or U7220 (N_7220,N_6527,N_6492);
nand U7221 (N_7221,N_6833,N_7130);
nor U7222 (N_7222,N_6961,N_6654);
or U7223 (N_7223,N_7118,N_6426);
or U7224 (N_7224,N_6645,N_6879);
nand U7225 (N_7225,N_7180,N_6658);
xor U7226 (N_7226,N_6897,N_6934);
nand U7227 (N_7227,N_6576,N_6623);
xor U7228 (N_7228,N_6519,N_6875);
and U7229 (N_7229,N_7012,N_7137);
and U7230 (N_7230,N_6512,N_6733);
or U7231 (N_7231,N_7075,N_6679);
nand U7232 (N_7232,N_7147,N_6662);
and U7233 (N_7233,N_6939,N_7037);
xor U7234 (N_7234,N_6567,N_7098);
xor U7235 (N_7235,N_7101,N_6700);
and U7236 (N_7236,N_6818,N_7124);
nand U7237 (N_7237,N_6545,N_7071);
nand U7238 (N_7238,N_7009,N_7189);
xnor U7239 (N_7239,N_7050,N_6848);
or U7240 (N_7240,N_6839,N_6999);
or U7241 (N_7241,N_6612,N_6859);
nand U7242 (N_7242,N_6799,N_6761);
and U7243 (N_7243,N_7041,N_6540);
nor U7244 (N_7244,N_6464,N_6971);
or U7245 (N_7245,N_6955,N_7125);
nor U7246 (N_7246,N_6950,N_6795);
nor U7247 (N_7247,N_6843,N_7056);
xnor U7248 (N_7248,N_6417,N_6621);
nor U7249 (N_7249,N_6513,N_6852);
nand U7250 (N_7250,N_6559,N_6981);
or U7251 (N_7251,N_7132,N_6862);
nand U7252 (N_7252,N_6425,N_6587);
or U7253 (N_7253,N_7184,N_7191);
xor U7254 (N_7254,N_6936,N_6990);
nand U7255 (N_7255,N_6806,N_6656);
nor U7256 (N_7256,N_7022,N_7024);
nand U7257 (N_7257,N_6607,N_6644);
or U7258 (N_7258,N_6771,N_6446);
nand U7259 (N_7259,N_6459,N_6794);
xnor U7260 (N_7260,N_6499,N_6995);
nor U7261 (N_7261,N_7136,N_6619);
nand U7262 (N_7262,N_6528,N_6603);
or U7263 (N_7263,N_6709,N_7015);
nand U7264 (N_7264,N_6766,N_6616);
or U7265 (N_7265,N_7077,N_7087);
nor U7266 (N_7266,N_6650,N_6977);
xor U7267 (N_7267,N_6819,N_6595);
nor U7268 (N_7268,N_6651,N_6599);
xor U7269 (N_7269,N_6923,N_6835);
or U7270 (N_7270,N_6776,N_6912);
nor U7271 (N_7271,N_6661,N_6867);
and U7272 (N_7272,N_6543,N_6407);
nand U7273 (N_7273,N_6521,N_6667);
nor U7274 (N_7274,N_6896,N_6641);
xnor U7275 (N_7275,N_6537,N_7079);
and U7276 (N_7276,N_6825,N_6404);
or U7277 (N_7277,N_6747,N_6834);
xnor U7278 (N_7278,N_6914,N_6707);
or U7279 (N_7279,N_6631,N_6952);
nor U7280 (N_7280,N_6774,N_6804);
nor U7281 (N_7281,N_6597,N_7083);
and U7282 (N_7282,N_7149,N_6401);
xor U7283 (N_7283,N_6716,N_6686);
nor U7284 (N_7284,N_6866,N_6449);
and U7285 (N_7285,N_6571,N_7074);
or U7286 (N_7286,N_6980,N_6458);
and U7287 (N_7287,N_6855,N_6778);
nor U7288 (N_7288,N_6687,N_6985);
nand U7289 (N_7289,N_7043,N_6578);
nand U7290 (N_7290,N_6719,N_7163);
nand U7291 (N_7291,N_6507,N_6523);
and U7292 (N_7292,N_6666,N_6501);
xor U7293 (N_7293,N_6826,N_6811);
nor U7294 (N_7294,N_6942,N_6857);
nor U7295 (N_7295,N_6472,N_6622);
and U7296 (N_7296,N_6663,N_6538);
xnor U7297 (N_7297,N_6788,N_6676);
nand U7298 (N_7298,N_6624,N_7193);
xor U7299 (N_7299,N_6926,N_6989);
xor U7300 (N_7300,N_6636,N_6902);
or U7301 (N_7301,N_7057,N_6511);
xor U7302 (N_7302,N_6470,N_6891);
nor U7303 (N_7303,N_6960,N_6596);
xor U7304 (N_7304,N_7046,N_7086);
or U7305 (N_7305,N_6730,N_6831);
xor U7306 (N_7306,N_7036,N_7069);
nor U7307 (N_7307,N_6544,N_6898);
nor U7308 (N_7308,N_6629,N_6531);
or U7309 (N_7309,N_6697,N_6944);
or U7310 (N_7310,N_6957,N_6638);
xnor U7311 (N_7311,N_7044,N_6781);
xnor U7312 (N_7312,N_7129,N_7062);
nand U7313 (N_7313,N_7081,N_6972);
or U7314 (N_7314,N_6910,N_7097);
and U7315 (N_7315,N_6782,N_6639);
xnor U7316 (N_7316,N_6966,N_6845);
nand U7317 (N_7317,N_7106,N_6429);
or U7318 (N_7318,N_7188,N_6557);
nor U7319 (N_7319,N_6648,N_7123);
and U7320 (N_7320,N_6979,N_6592);
nor U7321 (N_7321,N_6466,N_7064);
nor U7322 (N_7322,N_6455,N_6889);
xor U7323 (N_7323,N_7045,N_6454);
xnor U7324 (N_7324,N_6750,N_6529);
and U7325 (N_7325,N_6970,N_6605);
nor U7326 (N_7326,N_6533,N_6974);
or U7327 (N_7327,N_6993,N_6718);
or U7328 (N_7328,N_6784,N_7002);
and U7329 (N_7329,N_7038,N_7197);
nand U7330 (N_7330,N_6894,N_6920);
or U7331 (N_7331,N_6851,N_7148);
nor U7332 (N_7332,N_7127,N_6525);
xor U7333 (N_7333,N_6664,N_6868);
and U7334 (N_7334,N_7177,N_6440);
or U7335 (N_7335,N_6828,N_6413);
xnor U7336 (N_7336,N_6673,N_7082);
nor U7337 (N_7337,N_7152,N_6553);
nor U7338 (N_7338,N_7108,N_6640);
or U7339 (N_7339,N_6448,N_6468);
and U7340 (N_7340,N_6793,N_6675);
and U7341 (N_7341,N_6727,N_7187);
xor U7342 (N_7342,N_7140,N_6505);
xor U7343 (N_7343,N_6503,N_6935);
nand U7344 (N_7344,N_7194,N_6692);
and U7345 (N_7345,N_7067,N_6737);
and U7346 (N_7346,N_6518,N_6699);
nor U7347 (N_7347,N_7042,N_6618);
nand U7348 (N_7348,N_6473,N_7060);
nor U7349 (N_7349,N_7139,N_6988);
nand U7350 (N_7350,N_6690,N_6465);
xnor U7351 (N_7351,N_6924,N_7066);
and U7352 (N_7352,N_6941,N_6749);
and U7353 (N_7353,N_7165,N_6556);
xnor U7354 (N_7354,N_6508,N_6476);
or U7355 (N_7355,N_6689,N_7150);
xor U7356 (N_7356,N_6560,N_7091);
nor U7357 (N_7357,N_6504,N_6416);
xor U7358 (N_7358,N_6973,N_6704);
nor U7359 (N_7359,N_7021,N_6905);
nor U7360 (N_7360,N_7167,N_6581);
and U7361 (N_7361,N_6541,N_6715);
and U7362 (N_7362,N_6853,N_6570);
xor U7363 (N_7363,N_6997,N_6758);
nor U7364 (N_7364,N_7099,N_7052);
and U7365 (N_7365,N_6886,N_7153);
xnor U7366 (N_7366,N_6702,N_6703);
nor U7367 (N_7367,N_7113,N_6453);
or U7368 (N_7368,N_6824,N_6983);
nand U7369 (N_7369,N_6450,N_6943);
nand U7370 (N_7370,N_6551,N_6669);
nand U7371 (N_7371,N_6647,N_6877);
xnor U7372 (N_7372,N_6978,N_7031);
xor U7373 (N_7373,N_6633,N_6813);
nand U7374 (N_7374,N_7161,N_7003);
or U7375 (N_7375,N_6442,N_6608);
nor U7376 (N_7376,N_7126,N_6956);
or U7377 (N_7377,N_6695,N_7102);
xor U7378 (N_7378,N_6615,N_6844);
or U7379 (N_7379,N_6887,N_6477);
nand U7380 (N_7380,N_6967,N_6402);
and U7381 (N_7381,N_6756,N_6767);
nor U7382 (N_7382,N_7016,N_6791);
or U7383 (N_7383,N_6933,N_6445);
and U7384 (N_7384,N_7085,N_7076);
xnor U7385 (N_7385,N_6764,N_7058);
and U7386 (N_7386,N_6463,N_6418);
xor U7387 (N_7387,N_6849,N_6451);
xnor U7388 (N_7388,N_6907,N_6420);
nand U7389 (N_7389,N_6938,N_6701);
and U7390 (N_7390,N_6927,N_6899);
xnor U7391 (N_7391,N_6738,N_6610);
nand U7392 (N_7392,N_6515,N_6414);
and U7393 (N_7393,N_6814,N_6509);
xor U7394 (N_7394,N_6591,N_6723);
nand U7395 (N_7395,N_6741,N_6424);
xnor U7396 (N_7396,N_7073,N_6916);
and U7397 (N_7397,N_6482,N_7018);
nand U7398 (N_7398,N_6526,N_6604);
nand U7399 (N_7399,N_6883,N_7100);
nand U7400 (N_7400,N_6474,N_7199);
or U7401 (N_7401,N_7055,N_7092);
and U7402 (N_7402,N_6475,N_6432);
or U7403 (N_7403,N_7179,N_6439);
nor U7404 (N_7404,N_6549,N_6601);
nor U7405 (N_7405,N_6510,N_6860);
nor U7406 (N_7406,N_6447,N_6685);
nor U7407 (N_7407,N_7115,N_7030);
nand U7408 (N_7408,N_6547,N_7088);
nand U7409 (N_7409,N_6816,N_6817);
xor U7410 (N_7410,N_7104,N_6415);
or U7411 (N_7411,N_6837,N_6722);
and U7412 (N_7412,N_7181,N_6561);
nand U7413 (N_7413,N_6840,N_6421);
nor U7414 (N_7414,N_6913,N_6871);
xor U7415 (N_7415,N_6452,N_7017);
xnor U7416 (N_7416,N_7128,N_6400);
xor U7417 (N_7417,N_6542,N_6562);
nor U7418 (N_7418,N_6808,N_6683);
xnor U7419 (N_7419,N_6746,N_6969);
nand U7420 (N_7420,N_6823,N_6682);
nand U7421 (N_7421,N_6580,N_6487);
xor U7422 (N_7422,N_6665,N_6885);
nor U7423 (N_7423,N_6937,N_6951);
and U7424 (N_7424,N_6881,N_7133);
nor U7425 (N_7425,N_7172,N_7144);
and U7426 (N_7426,N_6740,N_7084);
nand U7427 (N_7427,N_6787,N_6670);
nor U7428 (N_7428,N_6932,N_6628);
or U7429 (N_7429,N_6801,N_6589);
nor U7430 (N_7430,N_6752,N_6829);
or U7431 (N_7431,N_6412,N_6655);
nand U7432 (N_7432,N_6732,N_6986);
and U7433 (N_7433,N_7116,N_6620);
xnor U7434 (N_7434,N_6770,N_6637);
nor U7435 (N_7435,N_6783,N_6965);
and U7436 (N_7436,N_6958,N_6456);
nand U7437 (N_7437,N_6968,N_6611);
nor U7438 (N_7438,N_6588,N_6947);
nor U7439 (N_7439,N_7198,N_6478);
or U7440 (N_7440,N_7154,N_6488);
xor U7441 (N_7441,N_6903,N_6461);
nand U7442 (N_7442,N_6590,N_7112);
nor U7443 (N_7443,N_6922,N_6550);
nand U7444 (N_7444,N_7089,N_6653);
and U7445 (N_7445,N_7134,N_6457);
or U7446 (N_7446,N_6946,N_7094);
or U7447 (N_7447,N_6630,N_6792);
or U7448 (N_7448,N_6409,N_7033);
or U7449 (N_7449,N_6945,N_6863);
nor U7450 (N_7450,N_6915,N_6874);
nor U7451 (N_7451,N_7174,N_7051);
nor U7452 (N_7452,N_7119,N_7166);
nand U7453 (N_7453,N_6635,N_7164);
xor U7454 (N_7454,N_7090,N_6713);
or U7455 (N_7455,N_7117,N_6674);
nand U7456 (N_7456,N_6514,N_6873);
nand U7457 (N_7457,N_6688,N_7011);
xor U7458 (N_7458,N_7168,N_6953);
nand U7459 (N_7459,N_7047,N_7131);
nand U7460 (N_7460,N_6726,N_6904);
nand U7461 (N_7461,N_6744,N_6724);
nand U7462 (N_7462,N_6876,N_6493);
xor U7463 (N_7463,N_7159,N_7103);
nor U7464 (N_7464,N_7093,N_6438);
xor U7465 (N_7465,N_6428,N_6671);
nor U7466 (N_7466,N_7151,N_6524);
nand U7467 (N_7467,N_6568,N_6491);
xnor U7468 (N_7468,N_6769,N_6554);
or U7469 (N_7469,N_6754,N_6921);
xor U7470 (N_7470,N_6882,N_7186);
xor U7471 (N_7471,N_6803,N_6495);
nand U7472 (N_7472,N_6575,N_6602);
or U7473 (N_7473,N_7143,N_7049);
or U7474 (N_7474,N_7027,N_6929);
or U7475 (N_7475,N_6757,N_6626);
nand U7476 (N_7476,N_7178,N_6861);
xor U7477 (N_7477,N_6534,N_6992);
or U7478 (N_7478,N_7135,N_6517);
and U7479 (N_7479,N_6516,N_6884);
and U7480 (N_7480,N_6546,N_6486);
nand U7481 (N_7481,N_6659,N_6433);
nand U7482 (N_7482,N_7196,N_6600);
and U7483 (N_7483,N_6780,N_7162);
nor U7484 (N_7484,N_6864,N_6696);
or U7485 (N_7485,N_6810,N_6900);
xnor U7486 (N_7486,N_6931,N_6821);
xnor U7487 (N_7487,N_7122,N_6502);
xnor U7488 (N_7488,N_7006,N_6632);
nor U7489 (N_7489,N_6573,N_6856);
nor U7490 (N_7490,N_6419,N_7138);
nand U7491 (N_7491,N_7000,N_6739);
or U7492 (N_7492,N_6613,N_6427);
xor U7493 (N_7493,N_6660,N_6735);
nor U7494 (N_7494,N_6717,N_6725);
nand U7495 (N_7495,N_6606,N_6480);
and U7496 (N_7496,N_7110,N_6530);
xor U7497 (N_7497,N_6755,N_7023);
and U7498 (N_7498,N_7020,N_6712);
xnor U7499 (N_7499,N_6646,N_7059);
or U7500 (N_7500,N_7029,N_6850);
or U7501 (N_7501,N_6668,N_7072);
and U7502 (N_7502,N_7008,N_6909);
and U7503 (N_7503,N_6652,N_6408);
and U7504 (N_7504,N_6930,N_6672);
nand U7505 (N_7505,N_7007,N_6405);
and U7506 (N_7506,N_6532,N_6569);
and U7507 (N_7507,N_6786,N_7034);
nor U7508 (N_7508,N_7183,N_6558);
or U7509 (N_7509,N_6431,N_6731);
xnor U7510 (N_7510,N_7170,N_6962);
nor U7511 (N_7511,N_7013,N_6830);
nor U7512 (N_7512,N_6564,N_6694);
nor U7513 (N_7513,N_7095,N_6982);
nor U7514 (N_7514,N_7080,N_6422);
nor U7515 (N_7515,N_7190,N_7068);
nand U7516 (N_7516,N_6964,N_7109);
nor U7517 (N_7517,N_7025,N_7063);
and U7518 (N_7518,N_7160,N_7141);
or U7519 (N_7519,N_6406,N_6759);
nand U7520 (N_7520,N_7156,N_7096);
nor U7521 (N_7521,N_6838,N_6467);
and U7522 (N_7522,N_6779,N_6579);
xnor U7523 (N_7523,N_7028,N_6649);
nor U7524 (N_7524,N_6609,N_6996);
nand U7525 (N_7525,N_6991,N_6798);
and U7526 (N_7526,N_6479,N_6797);
or U7527 (N_7527,N_7171,N_6745);
and U7528 (N_7528,N_7053,N_6772);
xnor U7529 (N_7529,N_7157,N_6911);
nand U7530 (N_7530,N_6711,N_7175);
or U7531 (N_7531,N_6762,N_7195);
nor U7532 (N_7532,N_6908,N_7111);
xnor U7533 (N_7533,N_7001,N_6586);
or U7534 (N_7534,N_6643,N_6460);
and U7535 (N_7535,N_6751,N_6872);
xnor U7536 (N_7536,N_6498,N_6893);
xor U7537 (N_7537,N_6497,N_6720);
nand U7538 (N_7538,N_6987,N_7185);
xnor U7539 (N_7539,N_6708,N_6627);
nand U7540 (N_7540,N_6765,N_6869);
xnor U7541 (N_7541,N_6742,N_6469);
nand U7542 (N_7542,N_7054,N_6763);
nor U7543 (N_7543,N_7004,N_6729);
or U7544 (N_7544,N_7121,N_6485);
or U7545 (N_7545,N_6959,N_6789);
nand U7546 (N_7546,N_6820,N_6584);
nor U7547 (N_7547,N_6680,N_6566);
or U7548 (N_7548,N_6918,N_6805);
or U7549 (N_7549,N_6594,N_6878);
nand U7550 (N_7550,N_6940,N_7014);
nor U7551 (N_7551,N_6481,N_6728);
nor U7552 (N_7552,N_6506,N_6858);
and U7553 (N_7553,N_6714,N_6444);
nor U7554 (N_7554,N_6753,N_6483);
and U7555 (N_7555,N_6583,N_6555);
xor U7556 (N_7556,N_6657,N_6736);
nand U7557 (N_7557,N_6494,N_6677);
nand U7558 (N_7558,N_7114,N_6865);
nor U7559 (N_7559,N_7182,N_7010);
nand U7560 (N_7560,N_6847,N_7173);
nor U7561 (N_7561,N_6434,N_7146);
xor U7562 (N_7562,N_6832,N_7078);
nor U7563 (N_7563,N_6822,N_6880);
nand U7564 (N_7564,N_6489,N_6522);
nand U7565 (N_7565,N_7019,N_6536);
nand U7566 (N_7566,N_6705,N_6691);
nand U7567 (N_7567,N_6411,N_6785);
nor U7568 (N_7568,N_6870,N_7192);
nor U7569 (N_7569,N_7169,N_7026);
nand U7570 (N_7570,N_6698,N_6800);
nor U7571 (N_7571,N_6565,N_6775);
or U7572 (N_7572,N_6593,N_6693);
or U7573 (N_7573,N_6790,N_6807);
nor U7574 (N_7574,N_6721,N_6888);
nor U7575 (N_7575,N_6928,N_6948);
xnor U7576 (N_7576,N_6572,N_6642);
or U7577 (N_7577,N_6614,N_6841);
and U7578 (N_7578,N_6917,N_6815);
nand U7579 (N_7579,N_6462,N_6552);
nand U7580 (N_7580,N_6490,N_6773);
or U7581 (N_7581,N_6678,N_6906);
nand U7582 (N_7582,N_6984,N_6895);
nand U7583 (N_7583,N_7032,N_6437);
nand U7584 (N_7584,N_6548,N_6734);
or U7585 (N_7585,N_6998,N_6430);
or U7586 (N_7586,N_6598,N_6743);
nor U7587 (N_7587,N_7176,N_6994);
nor U7588 (N_7588,N_6976,N_6423);
nor U7589 (N_7589,N_6500,N_7005);
or U7590 (N_7590,N_6892,N_6768);
nand U7591 (N_7591,N_7048,N_6582);
and U7592 (N_7592,N_6760,N_6441);
nand U7593 (N_7593,N_6846,N_6684);
nor U7594 (N_7594,N_7065,N_6901);
xor U7595 (N_7595,N_6748,N_6777);
or U7596 (N_7596,N_6403,N_7120);
or U7597 (N_7597,N_6617,N_6535);
nand U7598 (N_7598,N_6539,N_6574);
xnor U7599 (N_7599,N_7142,N_6681);
nand U7600 (N_7600,N_6755,N_6709);
or U7601 (N_7601,N_6517,N_7130);
and U7602 (N_7602,N_6853,N_6899);
nand U7603 (N_7603,N_6800,N_6754);
nor U7604 (N_7604,N_6751,N_7024);
xor U7605 (N_7605,N_6533,N_7048);
nor U7606 (N_7606,N_6418,N_6690);
nor U7607 (N_7607,N_7031,N_6854);
and U7608 (N_7608,N_6473,N_6854);
nor U7609 (N_7609,N_6656,N_7140);
and U7610 (N_7610,N_6745,N_6824);
xor U7611 (N_7611,N_6858,N_6940);
and U7612 (N_7612,N_6869,N_7055);
or U7613 (N_7613,N_6448,N_6835);
nor U7614 (N_7614,N_6502,N_6827);
nor U7615 (N_7615,N_6400,N_7016);
or U7616 (N_7616,N_7075,N_6669);
nor U7617 (N_7617,N_6651,N_7119);
nor U7618 (N_7618,N_7006,N_7062);
nand U7619 (N_7619,N_7120,N_6469);
and U7620 (N_7620,N_6662,N_6552);
xor U7621 (N_7621,N_6693,N_6534);
xor U7622 (N_7622,N_7055,N_7195);
nor U7623 (N_7623,N_6963,N_6499);
xor U7624 (N_7624,N_6688,N_7153);
xnor U7625 (N_7625,N_6811,N_6636);
xnor U7626 (N_7626,N_6936,N_6428);
and U7627 (N_7627,N_6508,N_6566);
nand U7628 (N_7628,N_7139,N_6701);
nor U7629 (N_7629,N_7197,N_6911);
or U7630 (N_7630,N_6837,N_6972);
nor U7631 (N_7631,N_7001,N_7184);
xor U7632 (N_7632,N_6623,N_6540);
xor U7633 (N_7633,N_7199,N_6774);
nor U7634 (N_7634,N_6668,N_6718);
nand U7635 (N_7635,N_6503,N_6874);
and U7636 (N_7636,N_6944,N_6740);
xnor U7637 (N_7637,N_7153,N_6574);
xnor U7638 (N_7638,N_6977,N_6787);
nor U7639 (N_7639,N_6732,N_6782);
nor U7640 (N_7640,N_6944,N_7131);
or U7641 (N_7641,N_6501,N_6911);
nor U7642 (N_7642,N_6904,N_6937);
xnor U7643 (N_7643,N_7041,N_6736);
and U7644 (N_7644,N_7016,N_6676);
nor U7645 (N_7645,N_6588,N_6478);
nand U7646 (N_7646,N_6953,N_7079);
xor U7647 (N_7647,N_6872,N_7049);
nor U7648 (N_7648,N_7049,N_6603);
nand U7649 (N_7649,N_6590,N_7026);
nand U7650 (N_7650,N_7189,N_6867);
xnor U7651 (N_7651,N_6854,N_6971);
or U7652 (N_7652,N_6695,N_6865);
nor U7653 (N_7653,N_6619,N_6584);
and U7654 (N_7654,N_7010,N_7125);
or U7655 (N_7655,N_6597,N_6429);
nand U7656 (N_7656,N_6473,N_7008);
xor U7657 (N_7657,N_7185,N_6958);
nor U7658 (N_7658,N_6879,N_6458);
xor U7659 (N_7659,N_6640,N_6985);
nor U7660 (N_7660,N_6786,N_6427);
nor U7661 (N_7661,N_6415,N_6670);
and U7662 (N_7662,N_7155,N_6706);
nor U7663 (N_7663,N_6833,N_6416);
xor U7664 (N_7664,N_6424,N_6510);
nand U7665 (N_7665,N_7004,N_6847);
and U7666 (N_7666,N_7170,N_6483);
xnor U7667 (N_7667,N_6951,N_6979);
nand U7668 (N_7668,N_6825,N_6997);
nand U7669 (N_7669,N_7007,N_6478);
and U7670 (N_7670,N_7081,N_6651);
nor U7671 (N_7671,N_6800,N_6994);
nor U7672 (N_7672,N_6908,N_6843);
nor U7673 (N_7673,N_6623,N_6962);
nor U7674 (N_7674,N_6899,N_7186);
nor U7675 (N_7675,N_6537,N_7111);
nand U7676 (N_7676,N_7040,N_6797);
nand U7677 (N_7677,N_6413,N_7087);
xnor U7678 (N_7678,N_7007,N_6667);
xor U7679 (N_7679,N_6875,N_6963);
and U7680 (N_7680,N_6748,N_6653);
nor U7681 (N_7681,N_6452,N_7155);
nand U7682 (N_7682,N_6956,N_6467);
and U7683 (N_7683,N_6718,N_6675);
nand U7684 (N_7684,N_6448,N_6784);
nor U7685 (N_7685,N_6853,N_6960);
or U7686 (N_7686,N_6464,N_6985);
xor U7687 (N_7687,N_7069,N_6538);
nor U7688 (N_7688,N_6862,N_6537);
nand U7689 (N_7689,N_7144,N_6935);
xnor U7690 (N_7690,N_6596,N_6669);
nor U7691 (N_7691,N_6869,N_6591);
xor U7692 (N_7692,N_6651,N_6682);
and U7693 (N_7693,N_7185,N_6729);
or U7694 (N_7694,N_6860,N_6708);
nor U7695 (N_7695,N_7164,N_7102);
nor U7696 (N_7696,N_7057,N_6666);
nor U7697 (N_7697,N_6941,N_6540);
or U7698 (N_7698,N_6683,N_6840);
or U7699 (N_7699,N_6907,N_6698);
or U7700 (N_7700,N_7185,N_6800);
xor U7701 (N_7701,N_6978,N_6906);
xnor U7702 (N_7702,N_6907,N_6998);
nor U7703 (N_7703,N_7025,N_6420);
or U7704 (N_7704,N_6667,N_7107);
nand U7705 (N_7705,N_6544,N_6879);
and U7706 (N_7706,N_7161,N_6971);
nand U7707 (N_7707,N_6655,N_6572);
xnor U7708 (N_7708,N_7010,N_6836);
nor U7709 (N_7709,N_6572,N_6640);
or U7710 (N_7710,N_6713,N_6856);
xnor U7711 (N_7711,N_7015,N_6836);
xor U7712 (N_7712,N_7160,N_6841);
nand U7713 (N_7713,N_6885,N_6474);
xor U7714 (N_7714,N_6823,N_6717);
and U7715 (N_7715,N_6529,N_7196);
and U7716 (N_7716,N_6423,N_6417);
or U7717 (N_7717,N_6815,N_7163);
nand U7718 (N_7718,N_6902,N_7127);
or U7719 (N_7719,N_6873,N_7116);
nand U7720 (N_7720,N_7114,N_7162);
xor U7721 (N_7721,N_6682,N_6708);
nor U7722 (N_7722,N_7102,N_6979);
and U7723 (N_7723,N_6815,N_6838);
or U7724 (N_7724,N_6652,N_7029);
xor U7725 (N_7725,N_6973,N_6765);
xnor U7726 (N_7726,N_6801,N_7159);
nor U7727 (N_7727,N_6481,N_6573);
nor U7728 (N_7728,N_6942,N_6555);
xnor U7729 (N_7729,N_7085,N_6790);
nand U7730 (N_7730,N_6756,N_6846);
nor U7731 (N_7731,N_6779,N_6704);
xnor U7732 (N_7732,N_7018,N_6412);
or U7733 (N_7733,N_6416,N_6418);
xor U7734 (N_7734,N_6568,N_7017);
nor U7735 (N_7735,N_6799,N_6470);
xnor U7736 (N_7736,N_6508,N_6855);
nor U7737 (N_7737,N_6577,N_6762);
and U7738 (N_7738,N_6655,N_7001);
xor U7739 (N_7739,N_6744,N_6469);
nor U7740 (N_7740,N_7079,N_6858);
and U7741 (N_7741,N_6967,N_7159);
nor U7742 (N_7742,N_6924,N_7166);
and U7743 (N_7743,N_6499,N_6423);
nor U7744 (N_7744,N_6459,N_6624);
nor U7745 (N_7745,N_6834,N_6944);
xor U7746 (N_7746,N_6527,N_7183);
xnor U7747 (N_7747,N_6777,N_6889);
nor U7748 (N_7748,N_6772,N_6693);
or U7749 (N_7749,N_6656,N_7155);
nand U7750 (N_7750,N_6943,N_6460);
xnor U7751 (N_7751,N_7002,N_6540);
xnor U7752 (N_7752,N_6659,N_6797);
and U7753 (N_7753,N_6402,N_7077);
and U7754 (N_7754,N_7114,N_6400);
xor U7755 (N_7755,N_6417,N_7145);
nand U7756 (N_7756,N_7143,N_6854);
and U7757 (N_7757,N_7116,N_7118);
xor U7758 (N_7758,N_6432,N_7145);
nand U7759 (N_7759,N_6570,N_6591);
nor U7760 (N_7760,N_7148,N_6472);
or U7761 (N_7761,N_6912,N_6961);
or U7762 (N_7762,N_6572,N_6899);
nor U7763 (N_7763,N_7087,N_6975);
nand U7764 (N_7764,N_7033,N_7109);
nand U7765 (N_7765,N_7139,N_7083);
xnor U7766 (N_7766,N_6820,N_6642);
and U7767 (N_7767,N_6902,N_6892);
xnor U7768 (N_7768,N_6927,N_6696);
nand U7769 (N_7769,N_6438,N_7182);
nor U7770 (N_7770,N_6929,N_7158);
or U7771 (N_7771,N_7113,N_7005);
or U7772 (N_7772,N_6548,N_6681);
or U7773 (N_7773,N_7100,N_7130);
and U7774 (N_7774,N_6749,N_6686);
or U7775 (N_7775,N_6528,N_6602);
nand U7776 (N_7776,N_6548,N_6633);
nand U7777 (N_7777,N_7134,N_6607);
xnor U7778 (N_7778,N_6401,N_6580);
or U7779 (N_7779,N_7100,N_6488);
and U7780 (N_7780,N_7071,N_6713);
or U7781 (N_7781,N_6583,N_6445);
xnor U7782 (N_7782,N_6906,N_6654);
nand U7783 (N_7783,N_6683,N_6855);
nand U7784 (N_7784,N_6792,N_7129);
nor U7785 (N_7785,N_7084,N_7040);
and U7786 (N_7786,N_6727,N_6619);
xor U7787 (N_7787,N_7181,N_6744);
nand U7788 (N_7788,N_6644,N_7187);
nor U7789 (N_7789,N_6957,N_6958);
nand U7790 (N_7790,N_6433,N_6924);
nand U7791 (N_7791,N_6824,N_6932);
xnor U7792 (N_7792,N_6968,N_6429);
or U7793 (N_7793,N_7140,N_6600);
or U7794 (N_7794,N_6991,N_6437);
and U7795 (N_7795,N_7072,N_6982);
nor U7796 (N_7796,N_7060,N_7017);
nor U7797 (N_7797,N_7198,N_6543);
nand U7798 (N_7798,N_6969,N_7133);
and U7799 (N_7799,N_7115,N_7164);
xnor U7800 (N_7800,N_7106,N_6541);
or U7801 (N_7801,N_6765,N_7183);
nor U7802 (N_7802,N_6562,N_6696);
nor U7803 (N_7803,N_6649,N_7123);
nand U7804 (N_7804,N_6492,N_6826);
and U7805 (N_7805,N_6850,N_6859);
or U7806 (N_7806,N_6749,N_6890);
or U7807 (N_7807,N_7055,N_7113);
or U7808 (N_7808,N_6847,N_6988);
nor U7809 (N_7809,N_6854,N_6717);
xnor U7810 (N_7810,N_6596,N_7105);
and U7811 (N_7811,N_6438,N_7147);
nand U7812 (N_7812,N_6980,N_6726);
or U7813 (N_7813,N_7145,N_6560);
nand U7814 (N_7814,N_6503,N_7023);
nand U7815 (N_7815,N_6744,N_6818);
and U7816 (N_7816,N_7026,N_7045);
or U7817 (N_7817,N_7176,N_6676);
or U7818 (N_7818,N_6842,N_6969);
nand U7819 (N_7819,N_6908,N_6958);
and U7820 (N_7820,N_6546,N_6981);
nor U7821 (N_7821,N_7036,N_6634);
or U7822 (N_7822,N_6757,N_7036);
xnor U7823 (N_7823,N_6942,N_7169);
nand U7824 (N_7824,N_7124,N_6868);
nand U7825 (N_7825,N_6832,N_6972);
nand U7826 (N_7826,N_6557,N_7135);
and U7827 (N_7827,N_6799,N_6552);
nand U7828 (N_7828,N_6530,N_6673);
nand U7829 (N_7829,N_6891,N_6509);
and U7830 (N_7830,N_6480,N_6783);
xor U7831 (N_7831,N_6698,N_6617);
nand U7832 (N_7832,N_6669,N_7031);
or U7833 (N_7833,N_6635,N_6584);
xor U7834 (N_7834,N_6911,N_6420);
and U7835 (N_7835,N_6761,N_6938);
nor U7836 (N_7836,N_6640,N_6685);
xor U7837 (N_7837,N_7184,N_6509);
or U7838 (N_7838,N_7162,N_6938);
and U7839 (N_7839,N_6749,N_7083);
nand U7840 (N_7840,N_6414,N_6834);
nor U7841 (N_7841,N_7186,N_7164);
or U7842 (N_7842,N_6865,N_7113);
xor U7843 (N_7843,N_6935,N_6739);
nor U7844 (N_7844,N_6715,N_7116);
or U7845 (N_7845,N_7150,N_6937);
xnor U7846 (N_7846,N_7147,N_6568);
or U7847 (N_7847,N_6714,N_6948);
xnor U7848 (N_7848,N_6497,N_7195);
nor U7849 (N_7849,N_7029,N_6695);
nand U7850 (N_7850,N_6810,N_7088);
nand U7851 (N_7851,N_7038,N_7021);
nor U7852 (N_7852,N_6647,N_6987);
nor U7853 (N_7853,N_6899,N_6818);
or U7854 (N_7854,N_6794,N_7118);
nor U7855 (N_7855,N_6984,N_6973);
or U7856 (N_7856,N_6708,N_6418);
or U7857 (N_7857,N_6902,N_6849);
nand U7858 (N_7858,N_7199,N_6758);
nor U7859 (N_7859,N_6619,N_6775);
xnor U7860 (N_7860,N_6431,N_6703);
or U7861 (N_7861,N_6569,N_6653);
nand U7862 (N_7862,N_6851,N_6553);
nand U7863 (N_7863,N_6499,N_7059);
and U7864 (N_7864,N_6878,N_6473);
nand U7865 (N_7865,N_6760,N_6599);
nand U7866 (N_7866,N_7175,N_6491);
or U7867 (N_7867,N_7098,N_6695);
nand U7868 (N_7868,N_6452,N_6638);
and U7869 (N_7869,N_7050,N_6723);
or U7870 (N_7870,N_6524,N_6618);
or U7871 (N_7871,N_6490,N_6650);
xor U7872 (N_7872,N_6506,N_6804);
xnor U7873 (N_7873,N_7120,N_6782);
or U7874 (N_7874,N_6705,N_6893);
and U7875 (N_7875,N_6907,N_7142);
and U7876 (N_7876,N_6557,N_6846);
xor U7877 (N_7877,N_6881,N_6647);
nand U7878 (N_7878,N_6671,N_6755);
nand U7879 (N_7879,N_6736,N_6883);
xnor U7880 (N_7880,N_7105,N_6661);
and U7881 (N_7881,N_7009,N_6545);
nand U7882 (N_7882,N_6878,N_6753);
nand U7883 (N_7883,N_7188,N_6733);
nand U7884 (N_7884,N_6890,N_6434);
xnor U7885 (N_7885,N_6828,N_7150);
xnor U7886 (N_7886,N_6471,N_6603);
xor U7887 (N_7887,N_6644,N_6884);
and U7888 (N_7888,N_6873,N_6875);
or U7889 (N_7889,N_7059,N_6865);
or U7890 (N_7890,N_7100,N_6947);
or U7891 (N_7891,N_7030,N_6484);
and U7892 (N_7892,N_6506,N_6694);
xnor U7893 (N_7893,N_6993,N_6554);
nand U7894 (N_7894,N_6738,N_6787);
nor U7895 (N_7895,N_6598,N_7009);
nand U7896 (N_7896,N_6520,N_6526);
xor U7897 (N_7897,N_7009,N_6622);
nand U7898 (N_7898,N_7021,N_6977);
nor U7899 (N_7899,N_6544,N_7043);
or U7900 (N_7900,N_7075,N_6629);
xor U7901 (N_7901,N_6965,N_6547);
and U7902 (N_7902,N_6673,N_6496);
and U7903 (N_7903,N_7132,N_6406);
xor U7904 (N_7904,N_6485,N_6489);
and U7905 (N_7905,N_6454,N_7031);
nor U7906 (N_7906,N_6756,N_7193);
and U7907 (N_7907,N_6568,N_7084);
nand U7908 (N_7908,N_6700,N_7033);
and U7909 (N_7909,N_7168,N_6623);
nor U7910 (N_7910,N_6496,N_6828);
xor U7911 (N_7911,N_6926,N_7177);
xnor U7912 (N_7912,N_6874,N_6838);
or U7913 (N_7913,N_6619,N_6881);
or U7914 (N_7914,N_6454,N_6570);
nor U7915 (N_7915,N_6474,N_6625);
xor U7916 (N_7916,N_6901,N_7189);
nand U7917 (N_7917,N_6784,N_7019);
nor U7918 (N_7918,N_7102,N_6767);
xnor U7919 (N_7919,N_6481,N_6528);
or U7920 (N_7920,N_6642,N_6802);
or U7921 (N_7921,N_7193,N_7028);
and U7922 (N_7922,N_6734,N_7031);
and U7923 (N_7923,N_6890,N_6773);
and U7924 (N_7924,N_6759,N_6666);
or U7925 (N_7925,N_6847,N_7061);
xor U7926 (N_7926,N_6702,N_7057);
and U7927 (N_7927,N_7021,N_7168);
and U7928 (N_7928,N_6679,N_6667);
or U7929 (N_7929,N_6704,N_6883);
xnor U7930 (N_7930,N_6499,N_6646);
nand U7931 (N_7931,N_6795,N_6788);
nor U7932 (N_7932,N_6840,N_6726);
and U7933 (N_7933,N_7065,N_7177);
xor U7934 (N_7934,N_6770,N_6985);
nor U7935 (N_7935,N_7146,N_6838);
nand U7936 (N_7936,N_7170,N_6923);
nand U7937 (N_7937,N_6764,N_6922);
nand U7938 (N_7938,N_6922,N_6457);
nand U7939 (N_7939,N_7194,N_7141);
xor U7940 (N_7940,N_6650,N_7044);
nor U7941 (N_7941,N_6867,N_6478);
xor U7942 (N_7942,N_6874,N_6516);
xor U7943 (N_7943,N_6633,N_6785);
xor U7944 (N_7944,N_6987,N_6993);
and U7945 (N_7945,N_6903,N_6641);
or U7946 (N_7946,N_6412,N_6924);
nor U7947 (N_7947,N_6993,N_6570);
xnor U7948 (N_7948,N_7165,N_6648);
nand U7949 (N_7949,N_6883,N_6957);
nor U7950 (N_7950,N_6939,N_6660);
nand U7951 (N_7951,N_6689,N_6830);
or U7952 (N_7952,N_6640,N_6983);
and U7953 (N_7953,N_6900,N_6882);
and U7954 (N_7954,N_7048,N_6579);
nand U7955 (N_7955,N_6681,N_6536);
or U7956 (N_7956,N_6760,N_6425);
xnor U7957 (N_7957,N_6711,N_6968);
nand U7958 (N_7958,N_6605,N_6769);
or U7959 (N_7959,N_7046,N_7187);
xnor U7960 (N_7960,N_6642,N_6949);
or U7961 (N_7961,N_6838,N_6506);
and U7962 (N_7962,N_6779,N_6492);
nand U7963 (N_7963,N_7033,N_7089);
nand U7964 (N_7964,N_6441,N_6653);
or U7965 (N_7965,N_6747,N_6917);
or U7966 (N_7966,N_7175,N_6961);
nand U7967 (N_7967,N_7147,N_7188);
nand U7968 (N_7968,N_6627,N_6451);
and U7969 (N_7969,N_6744,N_7081);
xnor U7970 (N_7970,N_7025,N_6917);
xor U7971 (N_7971,N_6566,N_6446);
xnor U7972 (N_7972,N_6749,N_6472);
and U7973 (N_7973,N_6881,N_6780);
nand U7974 (N_7974,N_7110,N_7111);
nand U7975 (N_7975,N_6688,N_6778);
or U7976 (N_7976,N_6405,N_6807);
and U7977 (N_7977,N_6430,N_6572);
nand U7978 (N_7978,N_6661,N_6796);
or U7979 (N_7979,N_7147,N_7068);
nand U7980 (N_7980,N_6430,N_7096);
and U7981 (N_7981,N_6759,N_6638);
nor U7982 (N_7982,N_6754,N_6412);
and U7983 (N_7983,N_6523,N_6755);
xor U7984 (N_7984,N_6476,N_6886);
nand U7985 (N_7985,N_7160,N_7012);
xnor U7986 (N_7986,N_6567,N_6917);
nor U7987 (N_7987,N_7051,N_6926);
nand U7988 (N_7988,N_7100,N_6946);
and U7989 (N_7989,N_7002,N_6682);
nor U7990 (N_7990,N_6801,N_6869);
or U7991 (N_7991,N_6760,N_6606);
xor U7992 (N_7992,N_6858,N_6959);
nand U7993 (N_7993,N_6681,N_7117);
and U7994 (N_7994,N_6632,N_6819);
or U7995 (N_7995,N_7082,N_6958);
xnor U7996 (N_7996,N_7014,N_6835);
nor U7997 (N_7997,N_6408,N_6748);
nand U7998 (N_7998,N_6439,N_6734);
and U7999 (N_7999,N_6692,N_6890);
and U8000 (N_8000,N_7438,N_7964);
xor U8001 (N_8001,N_7821,N_7374);
nor U8002 (N_8002,N_7809,N_7486);
nor U8003 (N_8003,N_7680,N_7969);
and U8004 (N_8004,N_7842,N_7246);
and U8005 (N_8005,N_7824,N_7553);
xor U8006 (N_8006,N_7443,N_7993);
nor U8007 (N_8007,N_7463,N_7274);
nor U8008 (N_8008,N_7696,N_7768);
and U8009 (N_8009,N_7854,N_7554);
xor U8010 (N_8010,N_7217,N_7365);
nand U8011 (N_8011,N_7644,N_7602);
and U8012 (N_8012,N_7725,N_7379);
or U8013 (N_8013,N_7745,N_7356);
nand U8014 (N_8014,N_7886,N_7785);
nor U8015 (N_8015,N_7892,N_7241);
nand U8016 (N_8016,N_7520,N_7867);
and U8017 (N_8017,N_7899,N_7701);
and U8018 (N_8018,N_7669,N_7782);
or U8019 (N_8019,N_7385,N_7593);
or U8020 (N_8020,N_7400,N_7411);
xnor U8021 (N_8021,N_7209,N_7851);
nor U8022 (N_8022,N_7789,N_7618);
xnor U8023 (N_8023,N_7600,N_7539);
and U8024 (N_8024,N_7818,N_7883);
and U8025 (N_8025,N_7447,N_7849);
nand U8026 (N_8026,N_7659,N_7406);
xor U8027 (N_8027,N_7691,N_7902);
and U8028 (N_8028,N_7927,N_7645);
nor U8029 (N_8029,N_7698,N_7757);
nand U8030 (N_8030,N_7586,N_7257);
xor U8031 (N_8031,N_7943,N_7233);
xnor U8032 (N_8032,N_7777,N_7709);
nand U8033 (N_8033,N_7956,N_7778);
xor U8034 (N_8034,N_7873,N_7200);
nor U8035 (N_8035,N_7389,N_7332);
nand U8036 (N_8036,N_7278,N_7773);
nor U8037 (N_8037,N_7948,N_7479);
or U8038 (N_8038,N_7499,N_7605);
xor U8039 (N_8039,N_7682,N_7910);
xor U8040 (N_8040,N_7531,N_7350);
and U8041 (N_8041,N_7419,N_7878);
xnor U8042 (N_8042,N_7940,N_7668);
or U8043 (N_8043,N_7937,N_7476);
and U8044 (N_8044,N_7321,N_7421);
xnor U8045 (N_8045,N_7863,N_7325);
or U8046 (N_8046,N_7399,N_7387);
nor U8047 (N_8047,N_7547,N_7997);
and U8048 (N_8048,N_7306,N_7326);
or U8049 (N_8049,N_7596,N_7633);
and U8050 (N_8050,N_7548,N_7265);
and U8051 (N_8051,N_7764,N_7654);
nor U8052 (N_8052,N_7660,N_7907);
or U8053 (N_8053,N_7527,N_7630);
or U8054 (N_8054,N_7951,N_7347);
or U8055 (N_8055,N_7670,N_7928);
nand U8056 (N_8056,N_7792,N_7378);
nor U8057 (N_8057,N_7995,N_7571);
xnor U8058 (N_8058,N_7311,N_7584);
nor U8059 (N_8059,N_7500,N_7360);
and U8060 (N_8060,N_7846,N_7252);
nand U8061 (N_8061,N_7860,N_7423);
and U8062 (N_8062,N_7800,N_7472);
and U8063 (N_8063,N_7296,N_7231);
nand U8064 (N_8064,N_7601,N_7739);
nand U8065 (N_8065,N_7493,N_7512);
nor U8066 (N_8066,N_7312,N_7895);
xor U8067 (N_8067,N_7555,N_7258);
or U8068 (N_8068,N_7716,N_7461);
xor U8069 (N_8069,N_7578,N_7333);
nand U8070 (N_8070,N_7575,N_7475);
xor U8071 (N_8071,N_7533,N_7297);
xnor U8072 (N_8072,N_7566,N_7408);
nand U8073 (N_8073,N_7637,N_7544);
or U8074 (N_8074,N_7636,N_7576);
nand U8075 (N_8075,N_7383,N_7699);
or U8076 (N_8076,N_7985,N_7609);
or U8077 (N_8077,N_7308,N_7715);
xnor U8078 (N_8078,N_7595,N_7759);
nor U8079 (N_8079,N_7449,N_7666);
xnor U8080 (N_8080,N_7727,N_7433);
nor U8081 (N_8081,N_7524,N_7638);
nor U8082 (N_8082,N_7407,N_7888);
nor U8083 (N_8083,N_7761,N_7319);
or U8084 (N_8084,N_7808,N_7359);
xor U8085 (N_8085,N_7288,N_7460);
or U8086 (N_8086,N_7429,N_7795);
or U8087 (N_8087,N_7410,N_7291);
or U8088 (N_8088,N_7958,N_7445);
and U8089 (N_8089,N_7677,N_7362);
nand U8090 (N_8090,N_7317,N_7405);
nor U8091 (N_8091,N_7482,N_7371);
and U8092 (N_8092,N_7642,N_7884);
or U8093 (N_8093,N_7661,N_7442);
nor U8094 (N_8094,N_7926,N_7237);
nor U8095 (N_8095,N_7511,N_7213);
or U8096 (N_8096,N_7890,N_7690);
xnor U8097 (N_8097,N_7372,N_7386);
nor U8098 (N_8098,N_7626,N_7802);
nand U8099 (N_8099,N_7728,N_7409);
nor U8100 (N_8100,N_7913,N_7313);
nor U8101 (N_8101,N_7718,N_7971);
and U8102 (N_8102,N_7263,N_7205);
nor U8103 (N_8103,N_7283,N_7494);
and U8104 (N_8104,N_7403,N_7394);
nor U8105 (N_8105,N_7304,N_7369);
nand U8106 (N_8106,N_7700,N_7562);
and U8107 (N_8107,N_7435,N_7623);
nand U8108 (N_8108,N_7906,N_7517);
or U8109 (N_8109,N_7489,N_7495);
nand U8110 (N_8110,N_7552,N_7624);
and U8111 (N_8111,N_7814,N_7545);
nand U8112 (N_8112,N_7535,N_7398);
or U8113 (N_8113,N_7478,N_7572);
xnor U8114 (N_8114,N_7504,N_7261);
xor U8115 (N_8115,N_7227,N_7949);
and U8116 (N_8116,N_7650,N_7567);
xnor U8117 (N_8117,N_7829,N_7464);
xnor U8118 (N_8118,N_7996,N_7806);
nand U8119 (N_8119,N_7747,N_7243);
xor U8120 (N_8120,N_7392,N_7542);
or U8121 (N_8121,N_7384,N_7991);
nor U8122 (N_8122,N_7760,N_7798);
and U8123 (N_8123,N_7268,N_7255);
nand U8124 (N_8124,N_7345,N_7856);
nor U8125 (N_8125,N_7961,N_7836);
or U8126 (N_8126,N_7735,N_7973);
and U8127 (N_8127,N_7862,N_7574);
nand U8128 (N_8128,N_7202,N_7339);
nor U8129 (N_8129,N_7525,N_7934);
nand U8130 (N_8130,N_7783,N_7483);
nor U8131 (N_8131,N_7331,N_7414);
or U8132 (N_8132,N_7388,N_7316);
xor U8133 (N_8133,N_7646,N_7242);
and U8134 (N_8134,N_7767,N_7613);
xnor U8135 (N_8135,N_7327,N_7397);
or U8136 (N_8136,N_7712,N_7451);
xor U8137 (N_8137,N_7556,N_7729);
nand U8138 (N_8138,N_7540,N_7929);
nor U8139 (N_8139,N_7695,N_7484);
or U8140 (N_8140,N_7876,N_7868);
and U8141 (N_8141,N_7568,N_7580);
or U8142 (N_8142,N_7828,N_7416);
nand U8143 (N_8143,N_7367,N_7726);
or U8144 (N_8144,N_7216,N_7507);
and U8145 (N_8145,N_7905,N_7582);
nand U8146 (N_8146,N_7830,N_7281);
nor U8147 (N_8147,N_7557,N_7551);
or U8148 (N_8148,N_7422,N_7864);
nor U8149 (N_8149,N_7244,N_7959);
xor U8150 (N_8150,N_7225,N_7226);
or U8151 (N_8151,N_7919,N_7275);
nor U8152 (N_8152,N_7505,N_7960);
xnor U8153 (N_8153,N_7625,N_7276);
and U8154 (N_8154,N_7466,N_7239);
and U8155 (N_8155,N_7742,N_7523);
and U8156 (N_8156,N_7901,N_7965);
nor U8157 (N_8157,N_7678,N_7685);
nand U8158 (N_8158,N_7672,N_7270);
nor U8159 (N_8159,N_7620,N_7285);
xnor U8160 (N_8160,N_7404,N_7541);
or U8161 (N_8161,N_7208,N_7381);
or U8162 (N_8162,N_7390,N_7247);
nand U8163 (N_8163,N_7355,N_7301);
or U8164 (N_8164,N_7318,N_7513);
nand U8165 (N_8165,N_7396,N_7315);
and U8166 (N_8166,N_7870,N_7748);
nand U8167 (N_8167,N_7713,N_7850);
nand U8168 (N_8168,N_7647,N_7269);
nand U8169 (N_8169,N_7791,N_7826);
or U8170 (N_8170,N_7653,N_7945);
or U8171 (N_8171,N_7819,N_7978);
xor U8172 (N_8172,N_7214,N_7245);
and U8173 (N_8173,N_7338,N_7236);
or U8174 (N_8174,N_7402,N_7323);
or U8175 (N_8175,N_7346,N_7815);
or U8176 (N_8176,N_7223,N_7840);
or U8177 (N_8177,N_7248,N_7457);
and U8178 (N_8178,N_7984,N_7454);
or U8179 (N_8179,N_7855,N_7229);
nor U8180 (N_8180,N_7234,N_7675);
nand U8181 (N_8181,N_7879,N_7272);
or U8182 (N_8182,N_7260,N_7847);
nor U8183 (N_8183,N_7564,N_7219);
xnor U8184 (N_8184,N_7731,N_7284);
and U8185 (N_8185,N_7320,N_7694);
nor U8186 (N_8186,N_7758,N_7627);
nand U8187 (N_8187,N_7775,N_7375);
nand U8188 (N_8188,N_7538,N_7914);
or U8189 (N_8189,N_7635,N_7287);
nand U8190 (N_8190,N_7615,N_7634);
and U8191 (N_8191,N_7865,N_7335);
xnor U8192 (N_8192,N_7790,N_7770);
nor U8193 (N_8193,N_7508,N_7866);
nand U8194 (N_8194,N_7684,N_7834);
or U8195 (N_8195,N_7652,N_7490);
xor U8196 (N_8196,N_7841,N_7293);
and U8197 (N_8197,N_7998,N_7262);
or U8198 (N_8198,N_7591,N_7752);
or U8199 (N_8199,N_7444,N_7577);
and U8200 (N_8200,N_7732,N_7762);
nand U8201 (N_8201,N_7616,N_7756);
or U8202 (N_8202,N_7631,N_7215);
xor U8203 (N_8203,N_7825,N_7665);
nor U8204 (N_8204,N_7295,N_7519);
xnor U8205 (N_8205,N_7707,N_7336);
nand U8206 (N_8206,N_7502,N_7933);
and U8207 (N_8207,N_7689,N_7380);
nand U8208 (N_8208,N_7772,N_7755);
xnor U8209 (N_8209,N_7376,N_7474);
nor U8210 (N_8210,N_7710,N_7455);
nand U8211 (N_8211,N_7947,N_7614);
nand U8212 (N_8212,N_7807,N_7763);
and U8213 (N_8213,N_7722,N_7990);
or U8214 (N_8214,N_7207,N_7881);
xor U8215 (N_8215,N_7664,N_7657);
or U8216 (N_8216,N_7393,N_7203);
and U8217 (N_8217,N_7655,N_7714);
or U8218 (N_8218,N_7885,N_7228);
xnor U8219 (N_8219,N_7453,N_7787);
xor U8220 (N_8220,N_7900,N_7897);
nand U8221 (N_8221,N_7342,N_7981);
xor U8222 (N_8222,N_7530,N_7820);
or U8223 (N_8223,N_7779,N_7412);
or U8224 (N_8224,N_7708,N_7277);
nand U8225 (N_8225,N_7737,N_7908);
nor U8226 (N_8226,N_7944,N_7280);
xor U8227 (N_8227,N_7251,N_7741);
or U8228 (N_8228,N_7711,N_7521);
xnor U8229 (N_8229,N_7509,N_7797);
or U8230 (N_8230,N_7324,N_7253);
or U8231 (N_8231,N_7939,N_7462);
nand U8232 (N_8232,N_7750,N_7796);
nor U8233 (N_8233,N_7617,N_7330);
xnor U8234 (N_8234,N_7608,N_7343);
or U8235 (N_8235,N_7230,N_7497);
nor U8236 (N_8236,N_7621,N_7279);
nor U8237 (N_8237,N_7922,N_7843);
nor U8238 (N_8238,N_7977,N_7989);
or U8239 (N_8239,N_7271,N_7559);
xnor U8240 (N_8240,N_7587,N_7799);
or U8241 (N_8241,N_7592,N_7703);
xnor U8242 (N_8242,N_7629,N_7204);
xnor U8243 (N_8243,N_7290,N_7292);
xnor U8244 (N_8244,N_7832,N_7719);
or U8245 (N_8245,N_7999,N_7861);
nor U8246 (N_8246,N_7780,N_7358);
xor U8247 (N_8247,N_7692,N_7667);
nand U8248 (N_8248,N_7982,N_7966);
or U8249 (N_8249,N_7480,N_7496);
and U8250 (N_8250,N_7754,N_7218);
or U8251 (N_8251,N_7781,N_7477);
xor U8252 (N_8252,N_7310,N_7534);
nand U8253 (N_8253,N_7425,N_7848);
nand U8254 (N_8254,N_7979,N_7721);
nand U8255 (N_8255,N_7370,N_7952);
nor U8256 (N_8256,N_7839,N_7329);
and U8257 (N_8257,N_7351,N_7932);
and U8258 (N_8258,N_7769,N_7417);
and U8259 (N_8259,N_7603,N_7904);
or U8260 (N_8260,N_7314,N_7220);
and U8261 (N_8261,N_7882,N_7891);
or U8262 (N_8262,N_7874,N_7286);
or U8263 (N_8263,N_7515,N_7349);
or U8264 (N_8264,N_7481,N_7210);
or U8265 (N_8265,N_7663,N_7923);
or U8266 (N_8266,N_7693,N_7859);
nor U8267 (N_8267,N_7606,N_7467);
xnor U8268 (N_8268,N_7305,N_7309);
xor U8269 (N_8269,N_7784,N_7546);
and U8270 (N_8270,N_7232,N_7528);
and U8271 (N_8271,N_7986,N_7340);
and U8272 (N_8272,N_7373,N_7456);
nand U8273 (N_8273,N_7604,N_7844);
xor U8274 (N_8274,N_7766,N_7887);
nand U8275 (N_8275,N_7734,N_7471);
or U8276 (N_8276,N_7681,N_7341);
xnor U8277 (N_8277,N_7898,N_7793);
or U8278 (N_8278,N_7501,N_7235);
nand U8279 (N_8279,N_7730,N_7240);
and U8280 (N_8280,N_7487,N_7550);
and U8281 (N_8281,N_7720,N_7440);
nor U8282 (N_8282,N_7622,N_7597);
or U8283 (N_8283,N_7869,N_7516);
and U8284 (N_8284,N_7212,N_7853);
or U8285 (N_8285,N_7671,N_7954);
and U8286 (N_8286,N_7628,N_7298);
nand U8287 (N_8287,N_7250,N_7201);
or U8288 (N_8288,N_7931,N_7915);
and U8289 (N_8289,N_7238,N_7683);
or U8290 (N_8290,N_7801,N_7794);
or U8291 (N_8291,N_7871,N_7590);
and U8292 (N_8292,N_7299,N_7938);
nand U8293 (N_8293,N_7746,N_7771);
nor U8294 (N_8294,N_7941,N_7401);
and U8295 (N_8295,N_7619,N_7676);
xnor U8296 (N_8296,N_7987,N_7537);
nor U8297 (N_8297,N_7413,N_7649);
or U8298 (N_8298,N_7302,N_7366);
xnor U8299 (N_8299,N_7450,N_7561);
nor U8300 (N_8300,N_7328,N_7266);
and U8301 (N_8301,N_7415,N_7599);
nor U8302 (N_8302,N_7852,N_7872);
xor U8303 (N_8303,N_7889,N_7289);
or U8304 (N_8304,N_7594,N_7822);
xnor U8305 (N_8305,N_7470,N_7452);
or U8306 (N_8306,N_7382,N_7465);
and U8307 (N_8307,N_7492,N_7988);
nand U8308 (N_8308,N_7503,N_7560);
nand U8309 (N_8309,N_7632,N_7570);
and U8310 (N_8310,N_7588,N_7514);
xnor U8311 (N_8311,N_7857,N_7536);
xor U8312 (N_8312,N_7448,N_7532);
and U8313 (N_8313,N_7804,N_7439);
nand U8314 (N_8314,N_7858,N_7723);
nor U8315 (N_8315,N_7221,N_7776);
and U8316 (N_8316,N_7607,N_7976);
nand U8317 (N_8317,N_7583,N_7563);
or U8318 (N_8318,N_7364,N_7975);
nand U8319 (N_8319,N_7651,N_7894);
and U8320 (N_8320,N_7222,N_7835);
nand U8321 (N_8321,N_7662,N_7935);
nor U8322 (N_8322,N_7686,N_7377);
xnor U8323 (N_8323,N_7968,N_7573);
nand U8324 (N_8324,N_7811,N_7877);
nand U8325 (N_8325,N_7294,N_7459);
and U8326 (N_8326,N_7611,N_7827);
nor U8327 (N_8327,N_7498,N_7909);
nor U8328 (N_8328,N_7980,N_7610);
nand U8329 (N_8329,N_7744,N_7344);
nand U8330 (N_8330,N_7648,N_7925);
and U8331 (N_8331,N_7921,N_7549);
or U8332 (N_8332,N_7434,N_7743);
nand U8333 (N_8333,N_7273,N_7640);
and U8334 (N_8334,N_7918,N_7936);
nor U8335 (N_8335,N_7348,N_7953);
xnor U8336 (N_8336,N_7446,N_7363);
nor U8337 (N_8337,N_7337,N_7983);
and U8338 (N_8338,N_7353,N_7427);
nand U8339 (N_8339,N_7585,N_7749);
and U8340 (N_8340,N_7352,N_7970);
and U8341 (N_8341,N_7643,N_7812);
and U8342 (N_8342,N_7837,N_7424);
or U8343 (N_8343,N_7704,N_7788);
or U8344 (N_8344,N_7673,N_7706);
xnor U8345 (N_8345,N_7522,N_7491);
nand U8346 (N_8346,N_7431,N_7441);
and U8347 (N_8347,N_7803,N_7805);
and U8348 (N_8348,N_7598,N_7823);
nor U8349 (N_8349,N_7724,N_7224);
nor U8350 (N_8350,N_7920,N_7436);
or U8351 (N_8351,N_7432,N_7418);
nand U8352 (N_8352,N_7994,N_7206);
and U8353 (N_8353,N_7967,N_7765);
xnor U8354 (N_8354,N_7430,N_7211);
or U8355 (N_8355,N_7426,N_7705);
nand U8356 (N_8356,N_7354,N_7813);
xor U8357 (N_8357,N_7697,N_7817);
nand U8358 (N_8358,N_7579,N_7946);
xnor U8359 (N_8359,N_7473,N_7656);
and U8360 (N_8360,N_7845,N_7893);
and U8361 (N_8361,N_7972,N_7903);
and U8362 (N_8362,N_7911,N_7838);
nor U8363 (N_8363,N_7485,N_7518);
nor U8364 (N_8364,N_7688,N_7917);
nand U8365 (N_8365,N_7880,N_7740);
xnor U8366 (N_8366,N_7589,N_7254);
and U8367 (N_8367,N_7930,N_7391);
nand U8368 (N_8368,N_7733,N_7974);
nand U8369 (N_8369,N_7992,N_7488);
nor U8370 (N_8370,N_7322,N_7963);
nor U8371 (N_8371,N_7831,N_7957);
xor U8372 (N_8372,N_7916,N_7529);
xnor U8373 (N_8373,N_7526,N_7420);
and U8374 (N_8374,N_7702,N_7612);
and U8375 (N_8375,N_7458,N_7658);
or U8376 (N_8376,N_7674,N_7833);
and U8377 (N_8377,N_7912,N_7942);
and U8378 (N_8378,N_7428,N_7639);
xor U8379 (N_8379,N_7924,N_7565);
nor U8380 (N_8380,N_7259,N_7469);
nand U8381 (N_8381,N_7955,N_7896);
and U8382 (N_8382,N_7581,N_7437);
nand U8383 (N_8383,N_7753,N_7687);
and U8384 (N_8384,N_7543,N_7264);
nand U8385 (N_8385,N_7816,N_7774);
xnor U8386 (N_8386,N_7357,N_7810);
and U8387 (N_8387,N_7300,N_7468);
and U8388 (N_8388,N_7641,N_7875);
or U8389 (N_8389,N_7361,N_7267);
xnor U8390 (N_8390,N_7510,N_7736);
nand U8391 (N_8391,N_7558,N_7395);
nand U8392 (N_8392,N_7738,N_7506);
and U8393 (N_8393,N_7950,N_7256);
or U8394 (N_8394,N_7679,N_7786);
xnor U8395 (N_8395,N_7307,N_7569);
nor U8396 (N_8396,N_7303,N_7962);
nand U8397 (N_8397,N_7368,N_7249);
nand U8398 (N_8398,N_7334,N_7751);
nand U8399 (N_8399,N_7282,N_7717);
or U8400 (N_8400,N_7768,N_7900);
or U8401 (N_8401,N_7266,N_7464);
and U8402 (N_8402,N_7552,N_7942);
nor U8403 (N_8403,N_7843,N_7201);
and U8404 (N_8404,N_7881,N_7728);
nor U8405 (N_8405,N_7560,N_7755);
nand U8406 (N_8406,N_7822,N_7849);
nor U8407 (N_8407,N_7960,N_7961);
or U8408 (N_8408,N_7608,N_7297);
or U8409 (N_8409,N_7840,N_7293);
nor U8410 (N_8410,N_7515,N_7282);
xor U8411 (N_8411,N_7681,N_7560);
nor U8412 (N_8412,N_7733,N_7681);
or U8413 (N_8413,N_7602,N_7392);
nand U8414 (N_8414,N_7667,N_7815);
or U8415 (N_8415,N_7711,N_7565);
nand U8416 (N_8416,N_7961,N_7580);
or U8417 (N_8417,N_7341,N_7769);
nand U8418 (N_8418,N_7957,N_7544);
xnor U8419 (N_8419,N_7382,N_7455);
nand U8420 (N_8420,N_7900,N_7268);
or U8421 (N_8421,N_7968,N_7239);
nor U8422 (N_8422,N_7519,N_7891);
nor U8423 (N_8423,N_7795,N_7239);
xnor U8424 (N_8424,N_7739,N_7317);
or U8425 (N_8425,N_7524,N_7357);
nor U8426 (N_8426,N_7894,N_7468);
or U8427 (N_8427,N_7857,N_7664);
nor U8428 (N_8428,N_7447,N_7264);
and U8429 (N_8429,N_7573,N_7664);
nand U8430 (N_8430,N_7267,N_7649);
nor U8431 (N_8431,N_7618,N_7661);
nand U8432 (N_8432,N_7732,N_7812);
and U8433 (N_8433,N_7456,N_7960);
or U8434 (N_8434,N_7279,N_7431);
xor U8435 (N_8435,N_7540,N_7326);
or U8436 (N_8436,N_7922,N_7406);
nor U8437 (N_8437,N_7809,N_7717);
nor U8438 (N_8438,N_7403,N_7298);
or U8439 (N_8439,N_7975,N_7837);
nand U8440 (N_8440,N_7517,N_7557);
xor U8441 (N_8441,N_7563,N_7714);
and U8442 (N_8442,N_7494,N_7750);
nand U8443 (N_8443,N_7209,N_7917);
nand U8444 (N_8444,N_7750,N_7930);
or U8445 (N_8445,N_7342,N_7632);
xnor U8446 (N_8446,N_7335,N_7745);
and U8447 (N_8447,N_7243,N_7944);
and U8448 (N_8448,N_7246,N_7971);
nor U8449 (N_8449,N_7842,N_7478);
or U8450 (N_8450,N_7984,N_7969);
xor U8451 (N_8451,N_7825,N_7353);
and U8452 (N_8452,N_7943,N_7973);
or U8453 (N_8453,N_7689,N_7710);
or U8454 (N_8454,N_7665,N_7706);
and U8455 (N_8455,N_7411,N_7669);
xor U8456 (N_8456,N_7279,N_7314);
and U8457 (N_8457,N_7922,N_7479);
or U8458 (N_8458,N_7962,N_7505);
xnor U8459 (N_8459,N_7933,N_7677);
xor U8460 (N_8460,N_7343,N_7204);
xor U8461 (N_8461,N_7241,N_7212);
xor U8462 (N_8462,N_7901,N_7779);
nor U8463 (N_8463,N_7461,N_7598);
xor U8464 (N_8464,N_7283,N_7576);
xor U8465 (N_8465,N_7370,N_7434);
nor U8466 (N_8466,N_7435,N_7871);
and U8467 (N_8467,N_7575,N_7520);
xnor U8468 (N_8468,N_7355,N_7584);
and U8469 (N_8469,N_7924,N_7577);
nand U8470 (N_8470,N_7265,N_7671);
xnor U8471 (N_8471,N_7894,N_7717);
and U8472 (N_8472,N_7447,N_7549);
or U8473 (N_8473,N_7206,N_7672);
or U8474 (N_8474,N_7395,N_7408);
and U8475 (N_8475,N_7953,N_7530);
or U8476 (N_8476,N_7331,N_7552);
or U8477 (N_8477,N_7206,N_7631);
xnor U8478 (N_8478,N_7609,N_7910);
nand U8479 (N_8479,N_7589,N_7412);
xor U8480 (N_8480,N_7626,N_7970);
xnor U8481 (N_8481,N_7958,N_7549);
nor U8482 (N_8482,N_7263,N_7522);
and U8483 (N_8483,N_7656,N_7963);
xnor U8484 (N_8484,N_7210,N_7295);
nand U8485 (N_8485,N_7200,N_7924);
xor U8486 (N_8486,N_7318,N_7579);
nand U8487 (N_8487,N_7323,N_7934);
or U8488 (N_8488,N_7418,N_7763);
or U8489 (N_8489,N_7402,N_7557);
nor U8490 (N_8490,N_7952,N_7407);
xnor U8491 (N_8491,N_7309,N_7958);
or U8492 (N_8492,N_7234,N_7756);
nand U8493 (N_8493,N_7824,N_7533);
and U8494 (N_8494,N_7253,N_7709);
or U8495 (N_8495,N_7577,N_7524);
nor U8496 (N_8496,N_7261,N_7412);
nand U8497 (N_8497,N_7385,N_7394);
or U8498 (N_8498,N_7501,N_7917);
or U8499 (N_8499,N_7364,N_7278);
nand U8500 (N_8500,N_7744,N_7845);
and U8501 (N_8501,N_7583,N_7816);
nor U8502 (N_8502,N_7571,N_7514);
or U8503 (N_8503,N_7789,N_7501);
or U8504 (N_8504,N_7878,N_7763);
xor U8505 (N_8505,N_7584,N_7327);
and U8506 (N_8506,N_7987,N_7272);
nand U8507 (N_8507,N_7798,N_7291);
xnor U8508 (N_8508,N_7720,N_7981);
nor U8509 (N_8509,N_7253,N_7827);
and U8510 (N_8510,N_7858,N_7416);
or U8511 (N_8511,N_7266,N_7706);
nor U8512 (N_8512,N_7422,N_7258);
and U8513 (N_8513,N_7445,N_7677);
nand U8514 (N_8514,N_7497,N_7498);
nand U8515 (N_8515,N_7698,N_7819);
or U8516 (N_8516,N_7755,N_7496);
nor U8517 (N_8517,N_7648,N_7261);
or U8518 (N_8518,N_7249,N_7859);
xor U8519 (N_8519,N_7233,N_7792);
nor U8520 (N_8520,N_7752,N_7281);
and U8521 (N_8521,N_7896,N_7436);
or U8522 (N_8522,N_7655,N_7999);
and U8523 (N_8523,N_7819,N_7906);
and U8524 (N_8524,N_7860,N_7991);
or U8525 (N_8525,N_7780,N_7341);
nand U8526 (N_8526,N_7285,N_7765);
and U8527 (N_8527,N_7609,N_7581);
and U8528 (N_8528,N_7443,N_7551);
xnor U8529 (N_8529,N_7791,N_7692);
nor U8530 (N_8530,N_7867,N_7422);
xor U8531 (N_8531,N_7405,N_7331);
xnor U8532 (N_8532,N_7585,N_7559);
nor U8533 (N_8533,N_7448,N_7390);
xor U8534 (N_8534,N_7820,N_7518);
or U8535 (N_8535,N_7337,N_7213);
or U8536 (N_8536,N_7691,N_7475);
and U8537 (N_8537,N_7398,N_7304);
and U8538 (N_8538,N_7648,N_7277);
or U8539 (N_8539,N_7985,N_7322);
nand U8540 (N_8540,N_7707,N_7648);
and U8541 (N_8541,N_7951,N_7262);
xor U8542 (N_8542,N_7979,N_7798);
nor U8543 (N_8543,N_7258,N_7469);
xnor U8544 (N_8544,N_7813,N_7317);
or U8545 (N_8545,N_7623,N_7452);
nor U8546 (N_8546,N_7490,N_7414);
or U8547 (N_8547,N_7516,N_7308);
xor U8548 (N_8548,N_7834,N_7585);
nor U8549 (N_8549,N_7287,N_7465);
nor U8550 (N_8550,N_7330,N_7659);
nand U8551 (N_8551,N_7387,N_7900);
nand U8552 (N_8552,N_7934,N_7724);
or U8553 (N_8553,N_7698,N_7813);
and U8554 (N_8554,N_7223,N_7615);
and U8555 (N_8555,N_7592,N_7253);
nand U8556 (N_8556,N_7556,N_7856);
and U8557 (N_8557,N_7587,N_7844);
nor U8558 (N_8558,N_7760,N_7655);
xnor U8559 (N_8559,N_7785,N_7200);
and U8560 (N_8560,N_7893,N_7831);
nand U8561 (N_8561,N_7247,N_7980);
and U8562 (N_8562,N_7664,N_7419);
nor U8563 (N_8563,N_7215,N_7715);
nor U8564 (N_8564,N_7497,N_7668);
or U8565 (N_8565,N_7262,N_7874);
xnor U8566 (N_8566,N_7850,N_7534);
nor U8567 (N_8567,N_7621,N_7544);
nor U8568 (N_8568,N_7268,N_7254);
or U8569 (N_8569,N_7703,N_7506);
xnor U8570 (N_8570,N_7910,N_7941);
nand U8571 (N_8571,N_7502,N_7838);
nand U8572 (N_8572,N_7708,N_7449);
nor U8573 (N_8573,N_7883,N_7539);
nand U8574 (N_8574,N_7924,N_7632);
nor U8575 (N_8575,N_7881,N_7311);
nor U8576 (N_8576,N_7734,N_7371);
nand U8577 (N_8577,N_7919,N_7203);
nand U8578 (N_8578,N_7608,N_7616);
nor U8579 (N_8579,N_7303,N_7329);
nor U8580 (N_8580,N_7578,N_7227);
nor U8581 (N_8581,N_7911,N_7285);
nand U8582 (N_8582,N_7563,N_7683);
nor U8583 (N_8583,N_7559,N_7789);
and U8584 (N_8584,N_7649,N_7463);
nor U8585 (N_8585,N_7727,N_7529);
nor U8586 (N_8586,N_7298,N_7773);
xnor U8587 (N_8587,N_7414,N_7863);
or U8588 (N_8588,N_7469,N_7204);
or U8589 (N_8589,N_7813,N_7855);
and U8590 (N_8590,N_7796,N_7468);
or U8591 (N_8591,N_7743,N_7796);
and U8592 (N_8592,N_7793,N_7602);
nand U8593 (N_8593,N_7480,N_7787);
nor U8594 (N_8594,N_7456,N_7474);
and U8595 (N_8595,N_7691,N_7606);
nand U8596 (N_8596,N_7941,N_7416);
or U8597 (N_8597,N_7866,N_7987);
nor U8598 (N_8598,N_7771,N_7951);
or U8599 (N_8599,N_7506,N_7342);
and U8600 (N_8600,N_7530,N_7310);
and U8601 (N_8601,N_7395,N_7583);
nor U8602 (N_8602,N_7249,N_7571);
nor U8603 (N_8603,N_7655,N_7464);
xor U8604 (N_8604,N_7502,N_7464);
and U8605 (N_8605,N_7397,N_7369);
nor U8606 (N_8606,N_7627,N_7633);
nand U8607 (N_8607,N_7533,N_7250);
or U8608 (N_8608,N_7291,N_7873);
nor U8609 (N_8609,N_7809,N_7801);
xnor U8610 (N_8610,N_7525,N_7674);
and U8611 (N_8611,N_7383,N_7605);
or U8612 (N_8612,N_7491,N_7802);
nand U8613 (N_8613,N_7760,N_7497);
nor U8614 (N_8614,N_7712,N_7260);
and U8615 (N_8615,N_7437,N_7981);
nand U8616 (N_8616,N_7935,N_7611);
nand U8617 (N_8617,N_7300,N_7268);
nor U8618 (N_8618,N_7979,N_7401);
nor U8619 (N_8619,N_7664,N_7985);
or U8620 (N_8620,N_7634,N_7702);
nand U8621 (N_8621,N_7633,N_7967);
xor U8622 (N_8622,N_7241,N_7767);
and U8623 (N_8623,N_7893,N_7721);
or U8624 (N_8624,N_7665,N_7447);
and U8625 (N_8625,N_7938,N_7356);
nor U8626 (N_8626,N_7356,N_7500);
nor U8627 (N_8627,N_7525,N_7564);
and U8628 (N_8628,N_7215,N_7672);
and U8629 (N_8629,N_7961,N_7342);
and U8630 (N_8630,N_7513,N_7787);
nand U8631 (N_8631,N_7910,N_7524);
nor U8632 (N_8632,N_7429,N_7419);
or U8633 (N_8633,N_7653,N_7673);
xnor U8634 (N_8634,N_7520,N_7864);
nor U8635 (N_8635,N_7614,N_7909);
or U8636 (N_8636,N_7576,N_7683);
or U8637 (N_8637,N_7581,N_7818);
nand U8638 (N_8638,N_7310,N_7818);
xnor U8639 (N_8639,N_7708,N_7736);
xor U8640 (N_8640,N_7817,N_7273);
and U8641 (N_8641,N_7875,N_7999);
nor U8642 (N_8642,N_7301,N_7587);
nor U8643 (N_8643,N_7505,N_7732);
or U8644 (N_8644,N_7765,N_7361);
nand U8645 (N_8645,N_7370,N_7312);
xor U8646 (N_8646,N_7896,N_7910);
and U8647 (N_8647,N_7579,N_7830);
nand U8648 (N_8648,N_7539,N_7698);
xnor U8649 (N_8649,N_7571,N_7793);
or U8650 (N_8650,N_7619,N_7797);
xor U8651 (N_8651,N_7263,N_7567);
nor U8652 (N_8652,N_7700,N_7524);
xor U8653 (N_8653,N_7568,N_7381);
xor U8654 (N_8654,N_7729,N_7350);
xor U8655 (N_8655,N_7520,N_7700);
xor U8656 (N_8656,N_7953,N_7978);
nand U8657 (N_8657,N_7376,N_7414);
xor U8658 (N_8658,N_7884,N_7230);
and U8659 (N_8659,N_7264,N_7528);
and U8660 (N_8660,N_7804,N_7503);
and U8661 (N_8661,N_7318,N_7492);
xnor U8662 (N_8662,N_7746,N_7842);
xor U8663 (N_8663,N_7562,N_7915);
and U8664 (N_8664,N_7669,N_7455);
xnor U8665 (N_8665,N_7621,N_7508);
and U8666 (N_8666,N_7611,N_7757);
or U8667 (N_8667,N_7557,N_7630);
nand U8668 (N_8668,N_7985,N_7536);
and U8669 (N_8669,N_7985,N_7776);
nand U8670 (N_8670,N_7807,N_7556);
nand U8671 (N_8671,N_7690,N_7826);
xor U8672 (N_8672,N_7905,N_7870);
or U8673 (N_8673,N_7803,N_7958);
nor U8674 (N_8674,N_7558,N_7866);
nand U8675 (N_8675,N_7965,N_7871);
nand U8676 (N_8676,N_7763,N_7824);
and U8677 (N_8677,N_7674,N_7611);
or U8678 (N_8678,N_7297,N_7801);
nand U8679 (N_8679,N_7246,N_7575);
xnor U8680 (N_8680,N_7398,N_7205);
and U8681 (N_8681,N_7454,N_7322);
nor U8682 (N_8682,N_7200,N_7884);
nand U8683 (N_8683,N_7220,N_7461);
or U8684 (N_8684,N_7746,N_7465);
xnor U8685 (N_8685,N_7976,N_7604);
nand U8686 (N_8686,N_7569,N_7957);
nor U8687 (N_8687,N_7398,N_7962);
or U8688 (N_8688,N_7611,N_7873);
and U8689 (N_8689,N_7489,N_7678);
and U8690 (N_8690,N_7243,N_7267);
and U8691 (N_8691,N_7984,N_7505);
nor U8692 (N_8692,N_7431,N_7863);
nand U8693 (N_8693,N_7755,N_7375);
xnor U8694 (N_8694,N_7537,N_7505);
or U8695 (N_8695,N_7506,N_7895);
xor U8696 (N_8696,N_7286,N_7207);
nand U8697 (N_8697,N_7581,N_7925);
xnor U8698 (N_8698,N_7551,N_7320);
or U8699 (N_8699,N_7985,N_7205);
or U8700 (N_8700,N_7492,N_7814);
or U8701 (N_8701,N_7825,N_7928);
nor U8702 (N_8702,N_7873,N_7606);
nand U8703 (N_8703,N_7790,N_7391);
xnor U8704 (N_8704,N_7640,N_7537);
or U8705 (N_8705,N_7457,N_7893);
nor U8706 (N_8706,N_7343,N_7282);
xnor U8707 (N_8707,N_7249,N_7323);
xnor U8708 (N_8708,N_7662,N_7623);
nor U8709 (N_8709,N_7734,N_7275);
and U8710 (N_8710,N_7736,N_7899);
xor U8711 (N_8711,N_7727,N_7919);
nand U8712 (N_8712,N_7909,N_7344);
nand U8713 (N_8713,N_7682,N_7697);
nand U8714 (N_8714,N_7505,N_7649);
nand U8715 (N_8715,N_7938,N_7218);
or U8716 (N_8716,N_7736,N_7206);
nor U8717 (N_8717,N_7961,N_7364);
and U8718 (N_8718,N_7501,N_7358);
and U8719 (N_8719,N_7470,N_7233);
xor U8720 (N_8720,N_7341,N_7963);
and U8721 (N_8721,N_7493,N_7421);
nor U8722 (N_8722,N_7314,N_7461);
or U8723 (N_8723,N_7529,N_7482);
or U8724 (N_8724,N_7883,N_7382);
xnor U8725 (N_8725,N_7695,N_7221);
xor U8726 (N_8726,N_7824,N_7777);
nor U8727 (N_8727,N_7864,N_7731);
and U8728 (N_8728,N_7817,N_7688);
or U8729 (N_8729,N_7471,N_7727);
nor U8730 (N_8730,N_7439,N_7251);
nand U8731 (N_8731,N_7922,N_7556);
nand U8732 (N_8732,N_7317,N_7710);
and U8733 (N_8733,N_7444,N_7321);
nand U8734 (N_8734,N_7258,N_7417);
or U8735 (N_8735,N_7795,N_7616);
and U8736 (N_8736,N_7982,N_7926);
or U8737 (N_8737,N_7503,N_7255);
and U8738 (N_8738,N_7404,N_7730);
nand U8739 (N_8739,N_7352,N_7864);
and U8740 (N_8740,N_7666,N_7740);
and U8741 (N_8741,N_7346,N_7412);
and U8742 (N_8742,N_7763,N_7276);
nand U8743 (N_8743,N_7689,N_7789);
nor U8744 (N_8744,N_7782,N_7685);
nand U8745 (N_8745,N_7995,N_7370);
xnor U8746 (N_8746,N_7858,N_7539);
xor U8747 (N_8747,N_7770,N_7679);
nand U8748 (N_8748,N_7830,N_7850);
nor U8749 (N_8749,N_7487,N_7704);
and U8750 (N_8750,N_7951,N_7954);
xnor U8751 (N_8751,N_7592,N_7806);
nand U8752 (N_8752,N_7776,N_7354);
xor U8753 (N_8753,N_7388,N_7321);
or U8754 (N_8754,N_7501,N_7387);
nand U8755 (N_8755,N_7809,N_7864);
nor U8756 (N_8756,N_7300,N_7569);
or U8757 (N_8757,N_7403,N_7455);
or U8758 (N_8758,N_7790,N_7974);
nor U8759 (N_8759,N_7287,N_7399);
and U8760 (N_8760,N_7475,N_7923);
nor U8761 (N_8761,N_7212,N_7673);
nor U8762 (N_8762,N_7422,N_7616);
xnor U8763 (N_8763,N_7659,N_7970);
nor U8764 (N_8764,N_7806,N_7284);
or U8765 (N_8765,N_7813,N_7405);
and U8766 (N_8766,N_7958,N_7267);
nand U8767 (N_8767,N_7553,N_7211);
nor U8768 (N_8768,N_7462,N_7459);
or U8769 (N_8769,N_7713,N_7685);
nor U8770 (N_8770,N_7684,N_7754);
and U8771 (N_8771,N_7681,N_7320);
xor U8772 (N_8772,N_7431,N_7584);
and U8773 (N_8773,N_7572,N_7711);
nor U8774 (N_8774,N_7339,N_7718);
nand U8775 (N_8775,N_7962,N_7611);
xnor U8776 (N_8776,N_7271,N_7675);
nand U8777 (N_8777,N_7459,N_7457);
or U8778 (N_8778,N_7707,N_7578);
or U8779 (N_8779,N_7394,N_7780);
or U8780 (N_8780,N_7390,N_7673);
nand U8781 (N_8781,N_7274,N_7381);
and U8782 (N_8782,N_7994,N_7683);
nor U8783 (N_8783,N_7597,N_7335);
or U8784 (N_8784,N_7664,N_7949);
xor U8785 (N_8785,N_7598,N_7613);
xnor U8786 (N_8786,N_7877,N_7215);
and U8787 (N_8787,N_7293,N_7943);
nor U8788 (N_8788,N_7443,N_7720);
nor U8789 (N_8789,N_7869,N_7802);
and U8790 (N_8790,N_7615,N_7433);
and U8791 (N_8791,N_7909,N_7705);
nand U8792 (N_8792,N_7703,N_7997);
nor U8793 (N_8793,N_7908,N_7834);
or U8794 (N_8794,N_7844,N_7742);
nor U8795 (N_8795,N_7520,N_7317);
or U8796 (N_8796,N_7678,N_7609);
or U8797 (N_8797,N_7683,N_7458);
and U8798 (N_8798,N_7455,N_7787);
nand U8799 (N_8799,N_7589,N_7221);
xor U8800 (N_8800,N_8644,N_8088);
nand U8801 (N_8801,N_8341,N_8419);
nand U8802 (N_8802,N_8460,N_8672);
nand U8803 (N_8803,N_8423,N_8440);
and U8804 (N_8804,N_8037,N_8430);
or U8805 (N_8805,N_8123,N_8707);
and U8806 (N_8806,N_8784,N_8477);
xor U8807 (N_8807,N_8732,N_8578);
xnor U8808 (N_8808,N_8696,N_8275);
and U8809 (N_8809,N_8655,N_8541);
xor U8810 (N_8810,N_8693,N_8555);
nand U8811 (N_8811,N_8794,N_8520);
nor U8812 (N_8812,N_8431,N_8399);
or U8813 (N_8813,N_8038,N_8730);
and U8814 (N_8814,N_8749,N_8428);
nand U8815 (N_8815,N_8156,N_8270);
and U8816 (N_8816,N_8791,N_8225);
and U8817 (N_8817,N_8393,N_8512);
xnor U8818 (N_8818,N_8280,N_8635);
nor U8819 (N_8819,N_8326,N_8146);
xnor U8820 (N_8820,N_8770,N_8669);
nand U8821 (N_8821,N_8528,N_8789);
and U8822 (N_8822,N_8467,N_8473);
nand U8823 (N_8823,N_8623,N_8165);
xnor U8824 (N_8824,N_8614,N_8637);
and U8825 (N_8825,N_8367,N_8666);
nor U8826 (N_8826,N_8765,N_8487);
nor U8827 (N_8827,N_8233,N_8774);
nand U8828 (N_8828,N_8650,N_8778);
nand U8829 (N_8829,N_8617,N_8040);
nor U8830 (N_8830,N_8621,N_8407);
nand U8831 (N_8831,N_8020,N_8539);
nand U8832 (N_8832,N_8099,N_8556);
and U8833 (N_8833,N_8200,N_8249);
and U8834 (N_8834,N_8334,N_8036);
and U8835 (N_8835,N_8530,N_8119);
nand U8836 (N_8836,N_8527,N_8365);
or U8837 (N_8837,N_8247,N_8612);
and U8838 (N_8838,N_8490,N_8754);
xor U8839 (N_8839,N_8733,N_8207);
nor U8840 (N_8840,N_8143,N_8421);
or U8841 (N_8841,N_8299,N_8759);
or U8842 (N_8842,N_8498,N_8435);
and U8843 (N_8843,N_8570,N_8258);
nor U8844 (N_8844,N_8149,N_8436);
and U8845 (N_8845,N_8057,N_8722);
nor U8846 (N_8846,N_8379,N_8357);
nand U8847 (N_8847,N_8736,N_8771);
or U8848 (N_8848,N_8226,N_8668);
xnor U8849 (N_8849,N_8402,N_8297);
xor U8850 (N_8850,N_8700,N_8538);
or U8851 (N_8851,N_8799,N_8508);
and U8852 (N_8852,N_8214,N_8027);
xor U8853 (N_8853,N_8479,N_8288);
nand U8854 (N_8854,N_8241,N_8380);
and U8855 (N_8855,N_8744,N_8132);
nand U8856 (N_8856,N_8093,N_8102);
or U8857 (N_8857,N_8150,N_8375);
nand U8858 (N_8858,N_8590,N_8568);
nand U8859 (N_8859,N_8321,N_8138);
nor U8860 (N_8860,N_8418,N_8389);
nor U8861 (N_8861,N_8386,N_8329);
nand U8862 (N_8862,N_8320,N_8608);
or U8863 (N_8863,N_8281,N_8118);
xor U8864 (N_8864,N_8602,N_8327);
or U8865 (N_8865,N_8176,N_8113);
nand U8866 (N_8866,N_8335,N_8363);
nand U8867 (N_8867,N_8352,N_8634);
xnor U8868 (N_8868,N_8464,N_8006);
or U8869 (N_8869,N_8441,N_8033);
nor U8870 (N_8870,N_8569,N_8661);
xnor U8871 (N_8871,N_8290,N_8208);
xor U8872 (N_8872,N_8412,N_8444);
nand U8873 (N_8873,N_8303,N_8346);
xor U8874 (N_8874,N_8348,N_8619);
xnor U8875 (N_8875,N_8395,N_8652);
nor U8876 (N_8876,N_8111,N_8776);
nand U8877 (N_8877,N_8211,N_8713);
nand U8878 (N_8878,N_8780,N_8000);
or U8879 (N_8879,N_8022,N_8725);
xnor U8880 (N_8880,N_8246,N_8576);
or U8881 (N_8881,N_8332,N_8628);
nor U8882 (N_8882,N_8454,N_8302);
nor U8883 (N_8883,N_8282,N_8345);
xor U8884 (N_8884,N_8007,N_8446);
or U8885 (N_8885,N_8550,N_8064);
nor U8886 (N_8886,N_8310,N_8383);
xor U8887 (N_8887,N_8372,N_8212);
or U8888 (N_8888,N_8307,N_8004);
nor U8889 (N_8889,N_8025,N_8315);
nand U8890 (N_8890,N_8748,N_8228);
or U8891 (N_8891,N_8083,N_8783);
and U8892 (N_8892,N_8674,N_8168);
or U8893 (N_8893,N_8698,N_8545);
or U8894 (N_8894,N_8021,N_8078);
and U8895 (N_8895,N_8710,N_8486);
or U8896 (N_8896,N_8114,N_8642);
and U8897 (N_8897,N_8174,N_8041);
xnor U8898 (N_8898,N_8731,N_8723);
nor U8899 (N_8899,N_8359,N_8283);
and U8900 (N_8900,N_8260,N_8178);
nand U8901 (N_8901,N_8092,N_8567);
and U8902 (N_8902,N_8458,N_8681);
and U8903 (N_8903,N_8468,N_8499);
xor U8904 (N_8904,N_8170,N_8437);
and U8905 (N_8905,N_8256,N_8003);
nor U8906 (N_8906,N_8456,N_8048);
nand U8907 (N_8907,N_8134,N_8662);
nor U8908 (N_8908,N_8414,N_8009);
nand U8909 (N_8909,N_8101,N_8404);
nor U8910 (N_8910,N_8793,N_8318);
nor U8911 (N_8911,N_8719,N_8366);
nand U8912 (N_8912,N_8071,N_8104);
nor U8913 (N_8913,N_8583,N_8442);
or U8914 (N_8914,N_8167,N_8300);
xor U8915 (N_8915,N_8394,N_8298);
xor U8916 (N_8916,N_8589,N_8471);
and U8917 (N_8917,N_8263,N_8139);
nand U8918 (N_8918,N_8096,N_8495);
nand U8919 (N_8919,N_8059,N_8551);
or U8920 (N_8920,N_8796,N_8429);
or U8921 (N_8921,N_8704,N_8355);
xnor U8922 (N_8922,N_8604,N_8218);
and U8923 (N_8923,N_8002,N_8264);
nand U8924 (N_8924,N_8209,N_8203);
nand U8925 (N_8925,N_8342,N_8517);
and U8926 (N_8926,N_8639,N_8144);
or U8927 (N_8927,N_8100,N_8023);
nor U8928 (N_8928,N_8239,N_8052);
xnor U8929 (N_8929,N_8177,N_8080);
nor U8930 (N_8930,N_8554,N_8559);
and U8931 (N_8931,N_8154,N_8409);
xor U8932 (N_8932,N_8109,N_8401);
and U8933 (N_8933,N_8561,N_8463);
nor U8934 (N_8934,N_8592,N_8449);
and U8935 (N_8935,N_8411,N_8254);
nand U8936 (N_8936,N_8746,N_8433);
xnor U8937 (N_8937,N_8739,N_8760);
nand U8938 (N_8938,N_8523,N_8136);
nand U8939 (N_8939,N_8245,N_8074);
and U8940 (N_8940,N_8728,N_8609);
and U8941 (N_8941,N_8358,N_8008);
nand U8942 (N_8942,N_8129,N_8549);
xnor U8943 (N_8943,N_8432,N_8232);
xor U8944 (N_8944,N_8788,N_8610);
nand U8945 (N_8945,N_8012,N_8516);
nor U8946 (N_8946,N_8761,N_8503);
or U8947 (N_8947,N_8277,N_8781);
xor U8948 (N_8948,N_8360,N_8511);
and U8949 (N_8949,N_8595,N_8684);
nand U8950 (N_8950,N_8660,N_8510);
nand U8951 (N_8951,N_8014,N_8271);
nand U8952 (N_8952,N_8124,N_8019);
xor U8953 (N_8953,N_8518,N_8647);
and U8954 (N_8954,N_8242,N_8257);
and U8955 (N_8955,N_8526,N_8373);
xor U8956 (N_8956,N_8658,N_8265);
nor U8957 (N_8957,N_8340,N_8183);
and U8958 (N_8958,N_8724,N_8391);
xor U8959 (N_8959,N_8267,N_8159);
xor U8960 (N_8960,N_8224,N_8304);
and U8961 (N_8961,N_8137,N_8331);
xor U8962 (N_8962,N_8613,N_8667);
nor U8963 (N_8963,N_8148,N_8145);
and U8964 (N_8964,N_8142,N_8173);
nor U8965 (N_8965,N_8544,N_8750);
xor U8966 (N_8966,N_8105,N_8675);
and U8967 (N_8967,N_8687,N_8127);
or U8968 (N_8968,N_8699,N_8362);
or U8969 (N_8969,N_8067,N_8534);
or U8970 (N_8970,N_8398,N_8076);
xor U8971 (N_8971,N_8587,N_8653);
nor U8972 (N_8972,N_8061,N_8546);
or U8973 (N_8973,N_8151,N_8206);
xnor U8974 (N_8974,N_8417,N_8155);
and U8975 (N_8975,N_8566,N_8255);
nor U8976 (N_8976,N_8797,N_8708);
and U8977 (N_8977,N_8356,N_8586);
nor U8978 (N_8978,N_8248,N_8175);
or U8979 (N_8979,N_8636,N_8035);
xnor U8980 (N_8980,N_8659,N_8115);
nand U8981 (N_8981,N_8054,N_8164);
or U8982 (N_8982,N_8447,N_8370);
nor U8983 (N_8983,N_8469,N_8643);
and U8984 (N_8984,N_8611,N_8714);
nand U8985 (N_8985,N_8287,N_8325);
nand U8986 (N_8986,N_8184,N_8677);
nand U8987 (N_8987,N_8032,N_8694);
and U8988 (N_8988,N_8396,N_8481);
xor U8989 (N_8989,N_8213,N_8751);
or U8990 (N_8990,N_8507,N_8483);
nor U8991 (N_8991,N_8237,N_8600);
nor U8992 (N_8992,N_8631,N_8285);
nand U8993 (N_8993,N_8034,N_8042);
nand U8994 (N_8994,N_8573,N_8221);
xnor U8995 (N_8995,N_8191,N_8376);
nand U8996 (N_8996,N_8439,N_8296);
xor U8997 (N_8997,N_8339,N_8266);
xor U8998 (N_8998,N_8438,N_8734);
nor U8999 (N_8999,N_8272,N_8787);
xnor U9000 (N_9000,N_8095,N_8065);
and U9001 (N_9001,N_8089,N_8795);
and U9002 (N_9002,N_8222,N_8056);
or U9003 (N_9003,N_8777,N_8491);
and U9004 (N_9004,N_8727,N_8347);
nor U9005 (N_9005,N_8082,N_8547);
xnor U9006 (N_9006,N_8024,N_8729);
or U9007 (N_9007,N_8311,N_8599);
xnor U9008 (N_9008,N_8755,N_8504);
nand U9009 (N_9009,N_8641,N_8575);
and U9010 (N_9010,N_8215,N_8651);
nor U9011 (N_9011,N_8524,N_8112);
xor U9012 (N_9012,N_8475,N_8273);
nor U9013 (N_9013,N_8645,N_8536);
or U9014 (N_9014,N_8349,N_8501);
xor U9015 (N_9015,N_8030,N_8090);
or U9016 (N_9016,N_8702,N_8664);
and U9017 (N_9017,N_8194,N_8336);
xnor U9018 (N_9018,N_8603,N_8403);
nand U9019 (N_9019,N_8584,N_8601);
and U9020 (N_9020,N_8210,N_8160);
nor U9021 (N_9021,N_8261,N_8676);
nand U9022 (N_9022,N_8616,N_8465);
or U9023 (N_9023,N_8654,N_8606);
nor U9024 (N_9024,N_8351,N_8186);
and U9025 (N_9025,N_8279,N_8262);
nor U9026 (N_9026,N_8535,N_8202);
nand U9027 (N_9027,N_8622,N_8779);
xor U9028 (N_9028,N_8286,N_8505);
nand U9029 (N_9029,N_8588,N_8294);
and U9030 (N_9030,N_8097,N_8010);
nor U9031 (N_9031,N_8615,N_8679);
or U9032 (N_9032,N_8462,N_8029);
nor U9033 (N_9033,N_8250,N_8678);
nand U9034 (N_9034,N_8764,N_8152);
and U9035 (N_9035,N_8532,N_8378);
or U9036 (N_9036,N_8049,N_8790);
nor U9037 (N_9037,N_8068,N_8459);
and U9038 (N_9038,N_8043,N_8408);
nand U9039 (N_9039,N_8742,N_8240);
and U9040 (N_9040,N_8697,N_8244);
or U9041 (N_9041,N_8564,N_8497);
nand U9042 (N_9042,N_8309,N_8709);
xor U9043 (N_9043,N_8513,N_8274);
nand U9044 (N_9044,N_8201,N_8354);
and U9045 (N_9045,N_8632,N_8182);
nor U9046 (N_9046,N_8166,N_8786);
nand U9047 (N_9047,N_8140,N_8514);
and U9048 (N_9048,N_8072,N_8392);
xor U9049 (N_9049,N_8542,N_8768);
and U9050 (N_9050,N_8716,N_8663);
nor U9051 (N_9051,N_8276,N_8682);
and U9052 (N_9052,N_8529,N_8133);
nand U9053 (N_9053,N_8251,N_8470);
xnor U9054 (N_9054,N_8085,N_8457);
nand U9055 (N_9055,N_8594,N_8044);
xnor U9056 (N_9056,N_8434,N_8405);
and U9057 (N_9057,N_8633,N_8116);
nand U9058 (N_9058,N_8344,N_8087);
nor U9059 (N_9059,N_8740,N_8673);
nor U9060 (N_9060,N_8525,N_8792);
xnor U9061 (N_9061,N_8492,N_8451);
nor U9062 (N_9062,N_8098,N_8427);
nand U9063 (N_9063,N_8762,N_8328);
and U9064 (N_9064,N_8130,N_8343);
xnor U9065 (N_9065,N_8553,N_8015);
nand U9066 (N_9066,N_8618,N_8188);
nand U9067 (N_9067,N_8016,N_8579);
xor U9068 (N_9068,N_8316,N_8323);
nand U9069 (N_9069,N_8598,N_8607);
and U9070 (N_9070,N_8195,N_8053);
nand U9071 (N_9071,N_8045,N_8718);
xor U9072 (N_9072,N_8077,N_8235);
nand U9073 (N_9073,N_8543,N_8135);
nand U9074 (N_9074,N_8190,N_8005);
or U9075 (N_9075,N_8521,N_8425);
and U9076 (N_9076,N_8063,N_8747);
xnor U9077 (N_9077,N_8688,N_8752);
nand U9078 (N_9078,N_8073,N_8585);
nand U9079 (N_9079,N_8665,N_8591);
xnor U9080 (N_9080,N_8397,N_8153);
or U9081 (N_9081,N_8001,N_8337);
nand U9082 (N_9082,N_8110,N_8324);
nor U9083 (N_9083,N_8686,N_8670);
nand U9084 (N_9084,N_8086,N_8482);
or U9085 (N_9085,N_8701,N_8291);
xnor U9086 (N_9086,N_8220,N_8253);
and U9087 (N_9087,N_8147,N_8306);
nand U9088 (N_9088,N_8785,N_8798);
nor U9089 (N_9089,N_8268,N_8120);
nor U9090 (N_9090,N_8572,N_8406);
and U9091 (N_9091,N_8531,N_8489);
xor U9092 (N_9092,N_8741,N_8199);
xor U9093 (N_9093,N_8715,N_8013);
nand U9094 (N_9094,N_8453,N_8743);
and U9095 (N_9095,N_8108,N_8314);
nand U9096 (N_9096,N_8782,N_8685);
nand U9097 (N_9097,N_8292,N_8361);
or U9098 (N_9098,N_8562,N_8624);
nor U9099 (N_9099,N_8705,N_8192);
and U9100 (N_9100,N_8767,N_8478);
nand U9101 (N_9101,N_8219,N_8091);
or U9102 (N_9102,N_8626,N_8070);
nand U9103 (N_9103,N_8364,N_8646);
xor U9104 (N_9104,N_8317,N_8476);
nand U9105 (N_9105,N_8560,N_8028);
nand U9106 (N_9106,N_8047,N_8313);
nand U9107 (N_9107,N_8066,N_8766);
or U9108 (N_9108,N_8128,N_8377);
or U9109 (N_9109,N_8197,N_8582);
and U9110 (N_9110,N_8301,N_8548);
nand U9111 (N_9111,N_8695,N_8690);
or U9112 (N_9112,N_8485,N_8390);
xnor U9113 (N_9113,N_8756,N_8079);
nand U9114 (N_9114,N_8494,N_8496);
or U9115 (N_9115,N_8493,N_8216);
nor U9116 (N_9116,N_8333,N_8236);
nand U9117 (N_9117,N_8243,N_8293);
and U9118 (N_9118,N_8671,N_8018);
nand U9119 (N_9119,N_8424,N_8757);
or U9120 (N_9120,N_8500,N_8450);
and U9121 (N_9121,N_8515,N_8062);
or U9122 (N_9122,N_8121,N_8422);
or U9123 (N_9123,N_8745,N_8410);
xor U9124 (N_9124,N_8163,N_8381);
nor U9125 (N_9125,N_8169,N_8400);
and U9126 (N_9126,N_8353,N_8758);
nor U9127 (N_9127,N_8691,N_8577);
or U9128 (N_9128,N_8330,N_8338);
nand U9129 (N_9129,N_8252,N_8103);
xor U9130 (N_9130,N_8571,N_8502);
xor U9131 (N_9131,N_8574,N_8051);
xor U9132 (N_9132,N_8131,N_8519);
nor U9133 (N_9133,N_8125,N_8187);
xor U9134 (N_9134,N_8231,N_8075);
or U9135 (N_9135,N_8107,N_8217);
nor U9136 (N_9136,N_8627,N_8480);
xor U9137 (N_9137,N_8769,N_8117);
or U9138 (N_9138,N_8726,N_8648);
xor U9139 (N_9139,N_8179,N_8558);
and U9140 (N_9140,N_8656,N_8374);
xor U9141 (N_9141,N_8060,N_8735);
nor U9142 (N_9142,N_8162,N_8448);
nor U9143 (N_9143,N_8017,N_8557);
nor U9144 (N_9144,N_8581,N_8420);
nand U9145 (N_9145,N_8039,N_8563);
and U9146 (N_9146,N_8753,N_8689);
nand U9147 (N_9147,N_8593,N_8312);
xnor U9148 (N_9148,N_8703,N_8385);
or U9149 (N_9149,N_8509,N_8657);
and U9150 (N_9150,N_8171,N_8484);
xnor U9151 (N_9151,N_8620,N_8721);
nand U9152 (N_9152,N_8238,N_8308);
nor U9153 (N_9153,N_8289,N_8181);
or U9154 (N_9154,N_8205,N_8680);
xnor U9155 (N_9155,N_8185,N_8106);
and U9156 (N_9156,N_8706,N_8229);
nand U9157 (N_9157,N_8522,N_8552);
nor U9158 (N_9158,N_8537,N_8058);
xnor U9159 (N_9159,N_8426,N_8466);
nand U9160 (N_9160,N_8069,N_8384);
and U9161 (N_9161,N_8773,N_8050);
nand U9162 (N_9162,N_8638,N_8046);
nor U9163 (N_9163,N_8772,N_8382);
nand U9164 (N_9164,N_8461,N_8720);
nor U9165 (N_9165,N_8605,N_8692);
or U9166 (N_9166,N_8269,N_8026);
nand U9167 (N_9167,N_8625,N_8227);
and U9168 (N_9168,N_8738,N_8597);
nand U9169 (N_9169,N_8158,N_8649);
nor U9170 (N_9170,N_8126,N_8540);
nor U9171 (N_9171,N_8506,N_8737);
or U9172 (N_9172,N_8443,N_8368);
and U9173 (N_9173,N_8284,N_8319);
nor U9174 (N_9174,N_8413,N_8416);
xnor U9175 (N_9175,N_8640,N_8278);
xnor U9176 (N_9176,N_8122,N_8630);
and U9177 (N_9177,N_8445,N_8474);
or U9178 (N_9178,N_8305,N_8196);
xnor U9179 (N_9179,N_8415,N_8712);
nor U9180 (N_9180,N_8180,N_8533);
nor U9181 (N_9181,N_8717,N_8596);
nand U9182 (N_9182,N_8230,N_8350);
nor U9183 (N_9183,N_8488,N_8081);
nand U9184 (N_9184,N_8094,N_8369);
nand U9185 (N_9185,N_8161,N_8371);
nor U9186 (N_9186,N_8683,N_8455);
xor U9187 (N_9187,N_8189,N_8204);
or U9188 (N_9188,N_8234,N_8580);
or U9189 (N_9189,N_8322,N_8388);
xnor U9190 (N_9190,N_8031,N_8711);
xnor U9191 (N_9191,N_8295,N_8011);
nand U9192 (N_9192,N_8084,N_8198);
and U9193 (N_9193,N_8193,N_8259);
or U9194 (N_9194,N_8055,N_8387);
nor U9195 (N_9195,N_8775,N_8141);
xnor U9196 (N_9196,N_8565,N_8157);
and U9197 (N_9197,N_8223,N_8763);
nor U9198 (N_9198,N_8472,N_8629);
or U9199 (N_9199,N_8172,N_8452);
xnor U9200 (N_9200,N_8470,N_8526);
nor U9201 (N_9201,N_8001,N_8374);
nor U9202 (N_9202,N_8173,N_8656);
or U9203 (N_9203,N_8047,N_8346);
xor U9204 (N_9204,N_8744,N_8647);
or U9205 (N_9205,N_8392,N_8129);
nor U9206 (N_9206,N_8791,N_8352);
nor U9207 (N_9207,N_8042,N_8590);
and U9208 (N_9208,N_8608,N_8714);
or U9209 (N_9209,N_8790,N_8018);
nand U9210 (N_9210,N_8623,N_8276);
xnor U9211 (N_9211,N_8643,N_8257);
nand U9212 (N_9212,N_8579,N_8504);
nor U9213 (N_9213,N_8052,N_8482);
xnor U9214 (N_9214,N_8352,N_8406);
xor U9215 (N_9215,N_8529,N_8136);
nand U9216 (N_9216,N_8581,N_8055);
xor U9217 (N_9217,N_8575,N_8461);
nand U9218 (N_9218,N_8262,N_8220);
nor U9219 (N_9219,N_8451,N_8493);
and U9220 (N_9220,N_8609,N_8024);
or U9221 (N_9221,N_8302,N_8408);
xnor U9222 (N_9222,N_8554,N_8460);
xor U9223 (N_9223,N_8382,N_8565);
xor U9224 (N_9224,N_8631,N_8328);
xor U9225 (N_9225,N_8423,N_8377);
xnor U9226 (N_9226,N_8212,N_8011);
or U9227 (N_9227,N_8442,N_8197);
nand U9228 (N_9228,N_8368,N_8544);
xor U9229 (N_9229,N_8627,N_8745);
xnor U9230 (N_9230,N_8624,N_8413);
or U9231 (N_9231,N_8758,N_8242);
nor U9232 (N_9232,N_8535,N_8267);
nor U9233 (N_9233,N_8429,N_8601);
nor U9234 (N_9234,N_8292,N_8456);
xnor U9235 (N_9235,N_8670,N_8251);
and U9236 (N_9236,N_8657,N_8489);
xnor U9237 (N_9237,N_8404,N_8218);
nand U9238 (N_9238,N_8133,N_8218);
or U9239 (N_9239,N_8548,N_8653);
nand U9240 (N_9240,N_8633,N_8033);
or U9241 (N_9241,N_8065,N_8013);
xnor U9242 (N_9242,N_8567,N_8101);
xor U9243 (N_9243,N_8472,N_8138);
nand U9244 (N_9244,N_8347,N_8604);
or U9245 (N_9245,N_8265,N_8747);
xnor U9246 (N_9246,N_8610,N_8780);
or U9247 (N_9247,N_8135,N_8226);
nand U9248 (N_9248,N_8719,N_8251);
nand U9249 (N_9249,N_8500,N_8776);
nor U9250 (N_9250,N_8771,N_8266);
nor U9251 (N_9251,N_8349,N_8125);
xnor U9252 (N_9252,N_8226,N_8002);
and U9253 (N_9253,N_8225,N_8179);
xnor U9254 (N_9254,N_8655,N_8089);
xor U9255 (N_9255,N_8568,N_8022);
and U9256 (N_9256,N_8727,N_8601);
or U9257 (N_9257,N_8239,N_8628);
or U9258 (N_9258,N_8409,N_8106);
or U9259 (N_9259,N_8589,N_8301);
nor U9260 (N_9260,N_8769,N_8708);
and U9261 (N_9261,N_8214,N_8174);
nor U9262 (N_9262,N_8701,N_8788);
xor U9263 (N_9263,N_8073,N_8179);
and U9264 (N_9264,N_8708,N_8109);
and U9265 (N_9265,N_8575,N_8171);
and U9266 (N_9266,N_8242,N_8584);
nand U9267 (N_9267,N_8520,N_8323);
nand U9268 (N_9268,N_8679,N_8347);
xnor U9269 (N_9269,N_8599,N_8164);
xnor U9270 (N_9270,N_8547,N_8167);
nor U9271 (N_9271,N_8245,N_8401);
nand U9272 (N_9272,N_8479,N_8651);
nor U9273 (N_9273,N_8036,N_8538);
or U9274 (N_9274,N_8303,N_8386);
or U9275 (N_9275,N_8711,N_8761);
nor U9276 (N_9276,N_8131,N_8403);
or U9277 (N_9277,N_8298,N_8220);
nor U9278 (N_9278,N_8302,N_8154);
and U9279 (N_9279,N_8445,N_8233);
and U9280 (N_9280,N_8231,N_8436);
and U9281 (N_9281,N_8767,N_8548);
and U9282 (N_9282,N_8422,N_8695);
or U9283 (N_9283,N_8679,N_8556);
nor U9284 (N_9284,N_8477,N_8386);
and U9285 (N_9285,N_8540,N_8665);
or U9286 (N_9286,N_8623,N_8028);
and U9287 (N_9287,N_8224,N_8460);
and U9288 (N_9288,N_8530,N_8065);
or U9289 (N_9289,N_8134,N_8280);
and U9290 (N_9290,N_8123,N_8357);
and U9291 (N_9291,N_8745,N_8215);
and U9292 (N_9292,N_8497,N_8364);
nor U9293 (N_9293,N_8393,N_8780);
nand U9294 (N_9294,N_8259,N_8655);
nor U9295 (N_9295,N_8288,N_8033);
and U9296 (N_9296,N_8308,N_8490);
or U9297 (N_9297,N_8207,N_8650);
xnor U9298 (N_9298,N_8772,N_8569);
xnor U9299 (N_9299,N_8451,N_8735);
nor U9300 (N_9300,N_8191,N_8757);
xor U9301 (N_9301,N_8485,N_8309);
nor U9302 (N_9302,N_8320,N_8362);
nand U9303 (N_9303,N_8199,N_8375);
xnor U9304 (N_9304,N_8284,N_8546);
and U9305 (N_9305,N_8088,N_8622);
nand U9306 (N_9306,N_8676,N_8457);
xor U9307 (N_9307,N_8467,N_8030);
xor U9308 (N_9308,N_8162,N_8492);
and U9309 (N_9309,N_8590,N_8745);
xnor U9310 (N_9310,N_8003,N_8283);
nand U9311 (N_9311,N_8630,N_8437);
or U9312 (N_9312,N_8216,N_8787);
or U9313 (N_9313,N_8462,N_8566);
xor U9314 (N_9314,N_8299,N_8055);
nor U9315 (N_9315,N_8425,N_8229);
nor U9316 (N_9316,N_8571,N_8495);
xor U9317 (N_9317,N_8699,N_8353);
or U9318 (N_9318,N_8037,N_8668);
and U9319 (N_9319,N_8380,N_8173);
and U9320 (N_9320,N_8414,N_8547);
xnor U9321 (N_9321,N_8366,N_8198);
nor U9322 (N_9322,N_8198,N_8788);
or U9323 (N_9323,N_8791,N_8249);
nand U9324 (N_9324,N_8528,N_8612);
and U9325 (N_9325,N_8546,N_8066);
and U9326 (N_9326,N_8526,N_8247);
nand U9327 (N_9327,N_8526,N_8591);
xnor U9328 (N_9328,N_8468,N_8730);
or U9329 (N_9329,N_8215,N_8152);
nor U9330 (N_9330,N_8608,N_8586);
nor U9331 (N_9331,N_8671,N_8379);
and U9332 (N_9332,N_8078,N_8288);
nor U9333 (N_9333,N_8579,N_8783);
and U9334 (N_9334,N_8199,N_8183);
xnor U9335 (N_9335,N_8472,N_8499);
or U9336 (N_9336,N_8770,N_8789);
and U9337 (N_9337,N_8795,N_8476);
and U9338 (N_9338,N_8102,N_8514);
nand U9339 (N_9339,N_8563,N_8063);
and U9340 (N_9340,N_8132,N_8124);
or U9341 (N_9341,N_8115,N_8502);
and U9342 (N_9342,N_8513,N_8325);
or U9343 (N_9343,N_8790,N_8765);
and U9344 (N_9344,N_8124,N_8279);
or U9345 (N_9345,N_8437,N_8580);
and U9346 (N_9346,N_8679,N_8140);
xor U9347 (N_9347,N_8662,N_8767);
xor U9348 (N_9348,N_8045,N_8374);
nor U9349 (N_9349,N_8081,N_8733);
xor U9350 (N_9350,N_8437,N_8521);
and U9351 (N_9351,N_8331,N_8368);
or U9352 (N_9352,N_8634,N_8786);
nor U9353 (N_9353,N_8448,N_8016);
xor U9354 (N_9354,N_8376,N_8159);
xnor U9355 (N_9355,N_8484,N_8035);
and U9356 (N_9356,N_8219,N_8680);
nand U9357 (N_9357,N_8605,N_8447);
xor U9358 (N_9358,N_8295,N_8157);
nand U9359 (N_9359,N_8335,N_8218);
nand U9360 (N_9360,N_8773,N_8159);
or U9361 (N_9361,N_8143,N_8171);
xor U9362 (N_9362,N_8572,N_8617);
nor U9363 (N_9363,N_8567,N_8341);
nand U9364 (N_9364,N_8076,N_8053);
nor U9365 (N_9365,N_8391,N_8334);
xnor U9366 (N_9366,N_8290,N_8153);
and U9367 (N_9367,N_8190,N_8289);
and U9368 (N_9368,N_8451,N_8475);
and U9369 (N_9369,N_8313,N_8491);
nor U9370 (N_9370,N_8316,N_8703);
nand U9371 (N_9371,N_8134,N_8349);
xnor U9372 (N_9372,N_8218,N_8772);
nor U9373 (N_9373,N_8256,N_8572);
xor U9374 (N_9374,N_8428,N_8215);
xnor U9375 (N_9375,N_8496,N_8775);
nor U9376 (N_9376,N_8347,N_8711);
xnor U9377 (N_9377,N_8063,N_8542);
and U9378 (N_9378,N_8050,N_8244);
nand U9379 (N_9379,N_8730,N_8144);
xnor U9380 (N_9380,N_8312,N_8441);
xnor U9381 (N_9381,N_8705,N_8227);
or U9382 (N_9382,N_8102,N_8167);
nor U9383 (N_9383,N_8368,N_8261);
nand U9384 (N_9384,N_8208,N_8532);
nand U9385 (N_9385,N_8014,N_8497);
nor U9386 (N_9386,N_8545,N_8446);
or U9387 (N_9387,N_8008,N_8158);
nand U9388 (N_9388,N_8454,N_8122);
xor U9389 (N_9389,N_8294,N_8015);
xnor U9390 (N_9390,N_8570,N_8441);
nor U9391 (N_9391,N_8240,N_8667);
xor U9392 (N_9392,N_8711,N_8597);
and U9393 (N_9393,N_8718,N_8088);
or U9394 (N_9394,N_8152,N_8038);
nor U9395 (N_9395,N_8510,N_8614);
and U9396 (N_9396,N_8120,N_8195);
nand U9397 (N_9397,N_8794,N_8111);
and U9398 (N_9398,N_8166,N_8260);
or U9399 (N_9399,N_8044,N_8487);
xnor U9400 (N_9400,N_8019,N_8666);
and U9401 (N_9401,N_8780,N_8777);
or U9402 (N_9402,N_8577,N_8512);
xor U9403 (N_9403,N_8216,N_8093);
nor U9404 (N_9404,N_8140,N_8610);
and U9405 (N_9405,N_8691,N_8464);
nand U9406 (N_9406,N_8000,N_8579);
nand U9407 (N_9407,N_8039,N_8354);
xnor U9408 (N_9408,N_8032,N_8129);
nand U9409 (N_9409,N_8452,N_8474);
and U9410 (N_9410,N_8505,N_8079);
and U9411 (N_9411,N_8349,N_8540);
and U9412 (N_9412,N_8647,N_8783);
xnor U9413 (N_9413,N_8770,N_8499);
nand U9414 (N_9414,N_8207,N_8164);
nor U9415 (N_9415,N_8287,N_8006);
nand U9416 (N_9416,N_8483,N_8513);
nor U9417 (N_9417,N_8283,N_8560);
xor U9418 (N_9418,N_8203,N_8158);
xnor U9419 (N_9419,N_8402,N_8572);
or U9420 (N_9420,N_8524,N_8788);
nand U9421 (N_9421,N_8495,N_8133);
or U9422 (N_9422,N_8626,N_8102);
xnor U9423 (N_9423,N_8626,N_8298);
nor U9424 (N_9424,N_8493,N_8281);
nor U9425 (N_9425,N_8177,N_8516);
nor U9426 (N_9426,N_8560,N_8548);
xnor U9427 (N_9427,N_8589,N_8162);
nand U9428 (N_9428,N_8414,N_8334);
xnor U9429 (N_9429,N_8424,N_8567);
or U9430 (N_9430,N_8218,N_8346);
nand U9431 (N_9431,N_8724,N_8195);
nor U9432 (N_9432,N_8128,N_8763);
or U9433 (N_9433,N_8693,N_8786);
nor U9434 (N_9434,N_8452,N_8176);
nand U9435 (N_9435,N_8053,N_8495);
nand U9436 (N_9436,N_8023,N_8385);
or U9437 (N_9437,N_8274,N_8237);
xor U9438 (N_9438,N_8295,N_8048);
nand U9439 (N_9439,N_8432,N_8528);
xor U9440 (N_9440,N_8246,N_8076);
nor U9441 (N_9441,N_8455,N_8624);
nor U9442 (N_9442,N_8649,N_8034);
nor U9443 (N_9443,N_8356,N_8711);
nor U9444 (N_9444,N_8082,N_8598);
nor U9445 (N_9445,N_8786,N_8161);
or U9446 (N_9446,N_8363,N_8068);
or U9447 (N_9447,N_8207,N_8589);
nand U9448 (N_9448,N_8511,N_8583);
and U9449 (N_9449,N_8276,N_8034);
nand U9450 (N_9450,N_8399,N_8531);
or U9451 (N_9451,N_8408,N_8369);
nand U9452 (N_9452,N_8342,N_8133);
or U9453 (N_9453,N_8715,N_8001);
and U9454 (N_9454,N_8736,N_8091);
or U9455 (N_9455,N_8028,N_8435);
nor U9456 (N_9456,N_8466,N_8290);
xor U9457 (N_9457,N_8218,N_8186);
nand U9458 (N_9458,N_8610,N_8692);
nand U9459 (N_9459,N_8370,N_8356);
or U9460 (N_9460,N_8399,N_8447);
nand U9461 (N_9461,N_8360,N_8559);
nand U9462 (N_9462,N_8201,N_8457);
and U9463 (N_9463,N_8703,N_8090);
nor U9464 (N_9464,N_8663,N_8475);
and U9465 (N_9465,N_8070,N_8510);
nand U9466 (N_9466,N_8135,N_8501);
nand U9467 (N_9467,N_8539,N_8372);
xnor U9468 (N_9468,N_8461,N_8677);
nor U9469 (N_9469,N_8306,N_8243);
or U9470 (N_9470,N_8353,N_8461);
nor U9471 (N_9471,N_8212,N_8710);
nand U9472 (N_9472,N_8530,N_8458);
nor U9473 (N_9473,N_8133,N_8242);
nand U9474 (N_9474,N_8119,N_8000);
or U9475 (N_9475,N_8604,N_8664);
nor U9476 (N_9476,N_8378,N_8538);
and U9477 (N_9477,N_8550,N_8008);
nor U9478 (N_9478,N_8103,N_8379);
nand U9479 (N_9479,N_8207,N_8360);
nor U9480 (N_9480,N_8414,N_8026);
and U9481 (N_9481,N_8702,N_8714);
xnor U9482 (N_9482,N_8181,N_8270);
nor U9483 (N_9483,N_8781,N_8331);
or U9484 (N_9484,N_8178,N_8771);
xor U9485 (N_9485,N_8027,N_8357);
and U9486 (N_9486,N_8715,N_8231);
and U9487 (N_9487,N_8038,N_8758);
and U9488 (N_9488,N_8712,N_8571);
xnor U9489 (N_9489,N_8242,N_8170);
nand U9490 (N_9490,N_8443,N_8562);
nor U9491 (N_9491,N_8692,N_8511);
nor U9492 (N_9492,N_8568,N_8258);
xor U9493 (N_9493,N_8368,N_8707);
nand U9494 (N_9494,N_8153,N_8377);
nor U9495 (N_9495,N_8273,N_8011);
and U9496 (N_9496,N_8765,N_8783);
nand U9497 (N_9497,N_8510,N_8092);
nand U9498 (N_9498,N_8476,N_8308);
nor U9499 (N_9499,N_8303,N_8770);
xnor U9500 (N_9500,N_8531,N_8449);
xnor U9501 (N_9501,N_8396,N_8232);
nor U9502 (N_9502,N_8710,N_8482);
nand U9503 (N_9503,N_8202,N_8777);
nand U9504 (N_9504,N_8598,N_8100);
nand U9505 (N_9505,N_8496,N_8743);
and U9506 (N_9506,N_8275,N_8553);
or U9507 (N_9507,N_8014,N_8236);
nor U9508 (N_9508,N_8486,N_8106);
and U9509 (N_9509,N_8061,N_8326);
nor U9510 (N_9510,N_8721,N_8338);
xor U9511 (N_9511,N_8201,N_8731);
xnor U9512 (N_9512,N_8787,N_8139);
and U9513 (N_9513,N_8594,N_8677);
nand U9514 (N_9514,N_8455,N_8439);
nand U9515 (N_9515,N_8592,N_8257);
nor U9516 (N_9516,N_8585,N_8394);
and U9517 (N_9517,N_8513,N_8573);
and U9518 (N_9518,N_8622,N_8467);
xor U9519 (N_9519,N_8104,N_8221);
nor U9520 (N_9520,N_8076,N_8485);
or U9521 (N_9521,N_8300,N_8107);
nor U9522 (N_9522,N_8438,N_8162);
nand U9523 (N_9523,N_8539,N_8231);
or U9524 (N_9524,N_8017,N_8467);
nand U9525 (N_9525,N_8439,N_8049);
nand U9526 (N_9526,N_8257,N_8446);
xor U9527 (N_9527,N_8798,N_8561);
and U9528 (N_9528,N_8563,N_8198);
nand U9529 (N_9529,N_8682,N_8481);
and U9530 (N_9530,N_8675,N_8290);
nand U9531 (N_9531,N_8661,N_8130);
and U9532 (N_9532,N_8445,N_8668);
nor U9533 (N_9533,N_8271,N_8151);
or U9534 (N_9534,N_8613,N_8072);
nor U9535 (N_9535,N_8458,N_8529);
xor U9536 (N_9536,N_8068,N_8532);
xor U9537 (N_9537,N_8787,N_8774);
nand U9538 (N_9538,N_8374,N_8437);
xnor U9539 (N_9539,N_8261,N_8341);
nor U9540 (N_9540,N_8786,N_8002);
or U9541 (N_9541,N_8541,N_8586);
or U9542 (N_9542,N_8162,N_8011);
nor U9543 (N_9543,N_8757,N_8241);
xnor U9544 (N_9544,N_8488,N_8024);
xnor U9545 (N_9545,N_8300,N_8331);
or U9546 (N_9546,N_8018,N_8059);
or U9547 (N_9547,N_8339,N_8568);
and U9548 (N_9548,N_8309,N_8620);
or U9549 (N_9549,N_8057,N_8216);
nand U9550 (N_9550,N_8183,N_8027);
xnor U9551 (N_9551,N_8547,N_8348);
or U9552 (N_9552,N_8788,N_8733);
nor U9553 (N_9553,N_8547,N_8717);
or U9554 (N_9554,N_8390,N_8113);
or U9555 (N_9555,N_8287,N_8023);
nor U9556 (N_9556,N_8133,N_8021);
or U9557 (N_9557,N_8566,N_8120);
xnor U9558 (N_9558,N_8549,N_8019);
xnor U9559 (N_9559,N_8372,N_8481);
or U9560 (N_9560,N_8248,N_8592);
and U9561 (N_9561,N_8332,N_8471);
xnor U9562 (N_9562,N_8498,N_8555);
or U9563 (N_9563,N_8564,N_8126);
nand U9564 (N_9564,N_8336,N_8785);
xnor U9565 (N_9565,N_8422,N_8635);
and U9566 (N_9566,N_8322,N_8407);
nor U9567 (N_9567,N_8256,N_8790);
xnor U9568 (N_9568,N_8294,N_8470);
xnor U9569 (N_9569,N_8168,N_8196);
or U9570 (N_9570,N_8258,N_8437);
nand U9571 (N_9571,N_8412,N_8358);
and U9572 (N_9572,N_8287,N_8730);
nand U9573 (N_9573,N_8741,N_8608);
nor U9574 (N_9574,N_8279,N_8068);
nor U9575 (N_9575,N_8740,N_8664);
nor U9576 (N_9576,N_8075,N_8558);
nand U9577 (N_9577,N_8451,N_8306);
or U9578 (N_9578,N_8486,N_8423);
xor U9579 (N_9579,N_8733,N_8625);
or U9580 (N_9580,N_8297,N_8105);
or U9581 (N_9581,N_8309,N_8473);
or U9582 (N_9582,N_8266,N_8315);
xor U9583 (N_9583,N_8214,N_8696);
xor U9584 (N_9584,N_8268,N_8427);
or U9585 (N_9585,N_8669,N_8642);
xnor U9586 (N_9586,N_8516,N_8476);
xor U9587 (N_9587,N_8028,N_8410);
or U9588 (N_9588,N_8048,N_8773);
nor U9589 (N_9589,N_8014,N_8701);
or U9590 (N_9590,N_8181,N_8283);
and U9591 (N_9591,N_8233,N_8217);
nor U9592 (N_9592,N_8340,N_8690);
nor U9593 (N_9593,N_8438,N_8132);
xor U9594 (N_9594,N_8764,N_8401);
and U9595 (N_9595,N_8721,N_8717);
and U9596 (N_9596,N_8607,N_8463);
or U9597 (N_9597,N_8211,N_8351);
or U9598 (N_9598,N_8495,N_8238);
or U9599 (N_9599,N_8152,N_8578);
and U9600 (N_9600,N_9301,N_9373);
or U9601 (N_9601,N_8964,N_9144);
and U9602 (N_9602,N_9315,N_9138);
and U9603 (N_9603,N_9199,N_9309);
and U9604 (N_9604,N_9344,N_8969);
xnor U9605 (N_9605,N_9079,N_9335);
xor U9606 (N_9606,N_9096,N_8972);
and U9607 (N_9607,N_9143,N_8902);
nand U9608 (N_9608,N_9302,N_9493);
or U9609 (N_9609,N_9191,N_8854);
nand U9610 (N_9610,N_8982,N_8816);
or U9611 (N_9611,N_9348,N_8909);
or U9612 (N_9612,N_8956,N_9072);
nand U9613 (N_9613,N_9537,N_8837);
xor U9614 (N_9614,N_8992,N_9027);
nor U9615 (N_9615,N_9416,N_9329);
and U9616 (N_9616,N_9317,N_9179);
and U9617 (N_9617,N_9100,N_9424);
and U9618 (N_9618,N_9193,N_9089);
nor U9619 (N_9619,N_9422,N_8937);
or U9620 (N_9620,N_9585,N_9380);
or U9621 (N_9621,N_8878,N_9375);
and U9622 (N_9622,N_9565,N_9261);
xnor U9623 (N_9623,N_9439,N_9256);
nor U9624 (N_9624,N_9248,N_9002);
nor U9625 (N_9625,N_9466,N_9107);
or U9626 (N_9626,N_9052,N_9112);
nand U9627 (N_9627,N_9201,N_9205);
or U9628 (N_9628,N_8965,N_9550);
xnor U9629 (N_9629,N_9022,N_9579);
nor U9630 (N_9630,N_9246,N_8876);
nor U9631 (N_9631,N_9404,N_9483);
xor U9632 (N_9632,N_9181,N_9127);
and U9633 (N_9633,N_9004,N_8825);
xor U9634 (N_9634,N_9133,N_9043);
nor U9635 (N_9635,N_9073,N_8974);
xnor U9636 (N_9636,N_9507,N_9474);
or U9637 (N_9637,N_8973,N_8840);
nand U9638 (N_9638,N_8946,N_9521);
and U9639 (N_9639,N_9170,N_9533);
xor U9640 (N_9640,N_9365,N_9054);
and U9641 (N_9641,N_9131,N_9172);
and U9642 (N_9642,N_8961,N_8872);
nor U9643 (N_9643,N_9018,N_9345);
or U9644 (N_9644,N_9279,N_9586);
or U9645 (N_9645,N_9599,N_8826);
nand U9646 (N_9646,N_9498,N_9406);
and U9647 (N_9647,N_8813,N_9058);
nor U9648 (N_9648,N_9413,N_9526);
or U9649 (N_9649,N_8870,N_9462);
and U9650 (N_9650,N_9254,N_9552);
and U9651 (N_9651,N_9129,N_8980);
nand U9652 (N_9652,N_9253,N_8806);
or U9653 (N_9653,N_9025,N_9470);
nand U9654 (N_9654,N_8987,N_9051);
nand U9655 (N_9655,N_8811,N_9557);
or U9656 (N_9656,N_8905,N_8831);
and U9657 (N_9657,N_9480,N_8950);
and U9658 (N_9658,N_9473,N_8908);
xnor U9659 (N_9659,N_9346,N_8868);
nor U9660 (N_9660,N_9490,N_9288);
and U9661 (N_9661,N_9192,N_9296);
or U9662 (N_9662,N_8986,N_9593);
nand U9663 (N_9663,N_8845,N_9103);
or U9664 (N_9664,N_9281,N_9056);
and U9665 (N_9665,N_9275,N_8881);
and U9666 (N_9666,N_9241,N_9083);
xnor U9667 (N_9667,N_8993,N_9469);
nor U9668 (N_9668,N_9313,N_9361);
nand U9669 (N_9669,N_8952,N_9321);
or U9670 (N_9670,N_9595,N_8838);
nand U9671 (N_9671,N_9578,N_9150);
nor U9672 (N_9672,N_9488,N_8927);
and U9673 (N_9673,N_9169,N_9023);
nor U9674 (N_9674,N_8829,N_9341);
xor U9675 (N_9675,N_9527,N_9377);
nand U9676 (N_9676,N_8917,N_9146);
nor U9677 (N_9677,N_9088,N_9095);
or U9678 (N_9678,N_9298,N_9177);
nor U9679 (N_9679,N_9401,N_9075);
nand U9680 (N_9680,N_9419,N_9260);
xnor U9681 (N_9681,N_9086,N_9568);
or U9682 (N_9682,N_9525,N_8985);
and U9683 (N_9683,N_9234,N_9399);
nor U9684 (N_9684,N_8896,N_9292);
and U9685 (N_9685,N_9496,N_9572);
and U9686 (N_9686,N_9139,N_9582);
nor U9687 (N_9687,N_9384,N_9325);
and U9688 (N_9688,N_9030,N_9354);
or U9689 (N_9689,N_9378,N_9124);
and U9690 (N_9690,N_9236,N_9487);
nand U9691 (N_9691,N_8884,N_9020);
nor U9692 (N_9692,N_9262,N_9269);
nand U9693 (N_9693,N_8941,N_9338);
nor U9694 (N_9694,N_9414,N_9102);
nand U9695 (N_9695,N_9409,N_9417);
and U9696 (N_9696,N_8955,N_9062);
or U9697 (N_9697,N_9125,N_9528);
nand U9698 (N_9698,N_8802,N_9195);
or U9699 (N_9699,N_8886,N_9464);
and U9700 (N_9700,N_8847,N_9598);
nor U9701 (N_9701,N_9478,N_9232);
and U9702 (N_9702,N_9012,N_8968);
nand U9703 (N_9703,N_8893,N_9295);
nor U9704 (N_9704,N_8991,N_9167);
nor U9705 (N_9705,N_8978,N_9000);
or U9706 (N_9706,N_8879,N_9505);
or U9707 (N_9707,N_9303,N_9364);
and U9708 (N_9708,N_9502,N_9251);
and U9709 (N_9709,N_8910,N_9554);
nand U9710 (N_9710,N_9531,N_8940);
and U9711 (N_9711,N_9575,N_9116);
xor U9712 (N_9712,N_8916,N_9064);
and U9713 (N_9713,N_8859,N_9060);
and U9714 (N_9714,N_9596,N_8810);
xor U9715 (N_9715,N_9265,N_9482);
and U9716 (N_9716,N_8979,N_9541);
and U9717 (N_9717,N_8867,N_8808);
xnor U9718 (N_9718,N_9589,N_8830);
nand U9719 (N_9719,N_9322,N_9036);
or U9720 (N_9720,N_9320,N_9220);
nand U9721 (N_9721,N_9190,N_9080);
nand U9722 (N_9722,N_9558,N_9277);
nor U9723 (N_9723,N_9115,N_8824);
xnor U9724 (N_9724,N_9007,N_9412);
nor U9725 (N_9725,N_8919,N_9436);
xor U9726 (N_9726,N_9046,N_9398);
and U9727 (N_9727,N_8915,N_9461);
and U9728 (N_9728,N_9147,N_8954);
xnor U9729 (N_9729,N_9119,N_9368);
and U9730 (N_9730,N_9421,N_8912);
nand U9731 (N_9731,N_9187,N_8809);
xor U9732 (N_9732,N_8981,N_9524);
xor U9733 (N_9733,N_9418,N_9494);
xnor U9734 (N_9734,N_9045,N_8836);
nand U9735 (N_9735,N_9397,N_9327);
nor U9736 (N_9736,N_8827,N_8938);
nor U9737 (N_9737,N_9238,N_8839);
and U9738 (N_9738,N_9209,N_8821);
nand U9739 (N_9739,N_9071,N_9009);
and U9740 (N_9740,N_9591,N_9135);
and U9741 (N_9741,N_9352,N_9429);
nand U9742 (N_9742,N_9032,N_9435);
xor U9743 (N_9743,N_8874,N_9411);
or U9744 (N_9744,N_9299,N_8846);
or U9745 (N_9745,N_8818,N_9061);
nand U9746 (N_9746,N_9420,N_9123);
nor U9747 (N_9747,N_8835,N_9529);
and U9748 (N_9748,N_9231,N_9158);
nand U9749 (N_9749,N_9316,N_9161);
nand U9750 (N_9750,N_9166,N_9442);
nand U9751 (N_9751,N_9546,N_9471);
and U9752 (N_9752,N_9349,N_9492);
or U9753 (N_9753,N_8988,N_9386);
xor U9754 (N_9754,N_9441,N_9110);
nor U9755 (N_9755,N_9068,N_9185);
and U9756 (N_9756,N_9148,N_9266);
nand U9757 (N_9757,N_8866,N_8819);
and U9758 (N_9758,N_8834,N_9567);
xnor U9759 (N_9759,N_9577,N_8924);
and U9760 (N_9760,N_9395,N_9287);
xor U9761 (N_9761,N_9021,N_9136);
or U9762 (N_9762,N_9211,N_8865);
nand U9763 (N_9763,N_8807,N_9297);
or U9764 (N_9764,N_9446,N_9559);
nand U9765 (N_9765,N_8892,N_9258);
nor U9766 (N_9766,N_9214,N_8820);
nand U9767 (N_9767,N_9433,N_9132);
and U9768 (N_9768,N_9081,N_9314);
nor U9769 (N_9769,N_9164,N_9540);
or U9770 (N_9770,N_9153,N_9370);
xnor U9771 (N_9771,N_8863,N_9070);
xnor U9772 (N_9772,N_9491,N_9434);
and U9773 (N_9773,N_8928,N_9458);
or U9774 (N_9774,N_9006,N_9067);
nand U9775 (N_9775,N_9029,N_9440);
nor U9776 (N_9776,N_9244,N_9035);
nand U9777 (N_9777,N_9113,N_9109);
xor U9778 (N_9778,N_9245,N_9311);
or U9779 (N_9779,N_8853,N_9207);
nor U9780 (N_9780,N_9485,N_9358);
nor U9781 (N_9781,N_9091,N_9233);
or U9782 (N_9782,N_9069,N_9118);
and U9783 (N_9783,N_8990,N_8862);
or U9784 (N_9784,N_9014,N_9049);
nand U9785 (N_9785,N_9504,N_9379);
nor U9786 (N_9786,N_8957,N_8959);
and U9787 (N_9787,N_8967,N_9114);
or U9788 (N_9788,N_9475,N_9188);
xnor U9789 (N_9789,N_9141,N_9182);
xor U9790 (N_9790,N_9210,N_9590);
nand U9791 (N_9791,N_8907,N_9282);
nor U9792 (N_9792,N_9180,N_8843);
xor U9793 (N_9793,N_9212,N_9323);
or U9794 (N_9794,N_8945,N_9084);
nor U9795 (N_9795,N_9184,N_9519);
xnor U9796 (N_9796,N_8857,N_9028);
xor U9797 (N_9797,N_9337,N_9534);
xnor U9798 (N_9798,N_9451,N_9351);
xor U9799 (N_9799,N_9237,N_8963);
and U9800 (N_9800,N_9447,N_8922);
nor U9801 (N_9801,N_8890,N_9425);
or U9802 (N_9802,N_8960,N_9553);
nand U9803 (N_9803,N_9548,N_9495);
or U9804 (N_9804,N_8888,N_8833);
or U9805 (N_9805,N_9396,N_9176);
or U9806 (N_9806,N_9134,N_9512);
nor U9807 (N_9807,N_9369,N_9592);
nand U9808 (N_9808,N_8856,N_9217);
nand U9809 (N_9809,N_9142,N_9250);
xor U9810 (N_9810,N_9339,N_9539);
nor U9811 (N_9811,N_8869,N_9165);
xnor U9812 (N_9812,N_9597,N_9410);
or U9813 (N_9813,N_9273,N_9569);
nor U9814 (N_9814,N_9532,N_8828);
nor U9815 (N_9815,N_9383,N_9518);
nand U9816 (N_9816,N_9571,N_9449);
nor U9817 (N_9817,N_9162,N_9555);
nor U9818 (N_9818,N_9218,N_9448);
or U9819 (N_9819,N_8920,N_9221);
and U9820 (N_9820,N_9503,N_9149);
and U9821 (N_9821,N_9168,N_8977);
nor U9822 (N_9822,N_8842,N_9264);
and U9823 (N_9823,N_9390,N_9357);
nor U9824 (N_9824,N_9216,N_9561);
xnor U9825 (N_9825,N_9223,N_9038);
or U9826 (N_9826,N_9003,N_9255);
xor U9827 (N_9827,N_8944,N_9268);
and U9828 (N_9828,N_9319,N_9055);
or U9829 (N_9829,N_9024,N_8804);
nand U9830 (N_9830,N_9001,N_8903);
and U9831 (N_9831,N_8971,N_9484);
or U9832 (N_9832,N_9120,N_9090);
and U9833 (N_9833,N_8898,N_9310);
and U9834 (N_9834,N_8958,N_9208);
and U9835 (N_9835,N_9031,N_9500);
or U9836 (N_9836,N_9355,N_8932);
nor U9837 (N_9837,N_9479,N_9326);
xor U9838 (N_9838,N_9366,N_9291);
or U9839 (N_9839,N_9359,N_9042);
or U9840 (N_9840,N_9108,N_9126);
nor U9841 (N_9841,N_9034,N_9226);
nor U9842 (N_9842,N_8914,N_9570);
and U9843 (N_9843,N_9497,N_9228);
and U9844 (N_9844,N_8844,N_8894);
and U9845 (N_9845,N_9085,N_9506);
or U9846 (N_9846,N_9230,N_8995);
and U9847 (N_9847,N_8887,N_8994);
xnor U9848 (N_9848,N_9290,N_9382);
or U9849 (N_9849,N_8975,N_9385);
nand U9850 (N_9850,N_9459,N_8947);
xor U9851 (N_9851,N_8976,N_8933);
nor U9852 (N_9852,N_8989,N_9186);
and U9853 (N_9853,N_9427,N_8882);
and U9854 (N_9854,N_8983,N_9300);
and U9855 (N_9855,N_9583,N_8899);
nor U9856 (N_9856,N_9536,N_8895);
nand U9857 (N_9857,N_9098,N_8871);
nand U9858 (N_9858,N_8923,N_8930);
nor U9859 (N_9859,N_9517,N_9306);
nand U9860 (N_9860,N_9015,N_9145);
and U9861 (N_9861,N_9453,N_8925);
and U9862 (N_9862,N_9580,N_9267);
nand U9863 (N_9863,N_9438,N_8805);
xnor U9864 (N_9864,N_9274,N_9039);
or U9865 (N_9865,N_9376,N_9252);
nand U9866 (N_9866,N_9155,N_9477);
nand U9867 (N_9867,N_8970,N_8900);
and U9868 (N_9868,N_9293,N_9171);
xor U9869 (N_9869,N_8997,N_9367);
nor U9870 (N_9870,N_9026,N_8904);
xnor U9871 (N_9871,N_9016,N_9574);
or U9872 (N_9872,N_9175,N_9157);
xor U9873 (N_9873,N_9286,N_9111);
nand U9874 (N_9874,N_8953,N_9432);
nor U9875 (N_9875,N_9128,N_9040);
nand U9876 (N_9876,N_9183,N_9222);
xor U9877 (N_9877,N_9332,N_9545);
nor U9878 (N_9878,N_9063,N_8812);
and U9879 (N_9879,N_9160,N_9202);
nor U9880 (N_9880,N_9400,N_8875);
nor U9881 (N_9881,N_9078,N_8848);
and U9882 (N_9882,N_9005,N_9249);
or U9883 (N_9883,N_9224,N_8901);
nor U9884 (N_9884,N_8935,N_9530);
nor U9885 (N_9885,N_8860,N_9394);
nand U9886 (N_9886,N_9393,N_9543);
xor U9887 (N_9887,N_9408,N_9362);
xor U9888 (N_9888,N_8911,N_9225);
nand U9889 (N_9889,N_9308,N_9305);
and U9890 (N_9890,N_9239,N_9444);
or U9891 (N_9891,N_9342,N_8936);
and U9892 (N_9892,N_9392,N_8889);
and U9893 (N_9893,N_9499,N_9074);
or U9894 (N_9894,N_9047,N_8801);
or U9895 (N_9895,N_8883,N_9510);
xnor U9896 (N_9896,N_9520,N_9227);
or U9897 (N_9897,N_9033,N_8913);
nand U9898 (N_9898,N_9066,N_9137);
nor U9899 (N_9899,N_9472,N_9371);
or U9900 (N_9900,N_9560,N_8817);
nand U9901 (N_9901,N_9304,N_9197);
nor U9902 (N_9902,N_8858,N_9562);
or U9903 (N_9903,N_9189,N_9271);
or U9904 (N_9904,N_9457,N_9247);
nor U9905 (N_9905,N_9280,N_9556);
nand U9906 (N_9906,N_9318,N_9391);
nand U9907 (N_9907,N_9152,N_9263);
nand U9908 (N_9908,N_8873,N_9324);
nor U9909 (N_9909,N_9523,N_9173);
and U9910 (N_9910,N_8885,N_9200);
or U9911 (N_9911,N_9513,N_9334);
nand U9912 (N_9912,N_9415,N_9094);
and U9913 (N_9913,N_8841,N_8861);
and U9914 (N_9914,N_9087,N_9460);
nand U9915 (N_9915,N_9121,N_8951);
or U9916 (N_9916,N_9122,N_9174);
xor U9917 (N_9917,N_9587,N_9041);
nand U9918 (N_9918,N_9456,N_8921);
xor U9919 (N_9919,N_9566,N_9538);
or U9920 (N_9920,N_9011,N_9285);
xor U9921 (N_9921,N_9544,N_9509);
xor U9922 (N_9922,N_8852,N_9381);
or U9923 (N_9923,N_9426,N_8823);
nor U9924 (N_9924,N_9343,N_9229);
or U9925 (N_9925,N_9455,N_9388);
nand U9926 (N_9926,N_9057,N_9476);
xor U9927 (N_9927,N_9563,N_9547);
or U9928 (N_9928,N_9278,N_9203);
nand U9929 (N_9929,N_9240,N_8999);
xor U9930 (N_9930,N_9452,N_9106);
xor U9931 (N_9931,N_9178,N_8891);
and U9932 (N_9932,N_9594,N_8906);
and U9933 (N_9933,N_8855,N_9235);
and U9934 (N_9934,N_9008,N_9551);
nand U9935 (N_9935,N_9289,N_9454);
nor U9936 (N_9936,N_9387,N_9053);
nor U9937 (N_9937,N_9159,N_9204);
and U9938 (N_9938,N_9564,N_9307);
or U9939 (N_9939,N_9501,N_8822);
and U9940 (N_9940,N_9196,N_9328);
nor U9941 (N_9941,N_9336,N_9481);
xnor U9942 (N_9942,N_8814,N_9065);
nor U9943 (N_9943,N_9219,N_9489);
or U9944 (N_9944,N_9353,N_9431);
and U9945 (N_9945,N_9584,N_9140);
and U9946 (N_9946,N_9340,N_9372);
or U9947 (N_9947,N_9092,N_8849);
nand U9948 (N_9948,N_9099,N_9356);
xnor U9949 (N_9949,N_9389,N_9010);
nor U9950 (N_9950,N_8948,N_8966);
nand U9951 (N_9951,N_9194,N_9573);
nor U9952 (N_9952,N_9515,N_8864);
nand U9953 (N_9953,N_8803,N_8943);
nand U9954 (N_9954,N_9312,N_9468);
nand U9955 (N_9955,N_9430,N_9516);
xnor U9956 (N_9956,N_8880,N_8897);
nor U9957 (N_9957,N_8800,N_9059);
nor U9958 (N_9958,N_8998,N_9076);
nor U9959 (N_9959,N_9511,N_9017);
or U9960 (N_9960,N_9486,N_9276);
or U9961 (N_9961,N_9101,N_8877);
or U9962 (N_9962,N_9104,N_8918);
or U9963 (N_9963,N_9363,N_9156);
and U9964 (N_9964,N_8934,N_9549);
and U9965 (N_9965,N_9467,N_9163);
and U9966 (N_9966,N_9463,N_9130);
nor U9967 (N_9967,N_9465,N_9019);
or U9968 (N_9968,N_9403,N_9050);
nor U9969 (N_9969,N_9522,N_8926);
nor U9970 (N_9970,N_9443,N_8832);
nand U9971 (N_9971,N_8962,N_8996);
or U9972 (N_9972,N_9283,N_9350);
and U9973 (N_9973,N_8931,N_9374);
xnor U9974 (N_9974,N_9097,N_8929);
nor U9975 (N_9975,N_9270,N_9259);
xor U9976 (N_9976,N_9082,N_9272);
or U9977 (N_9977,N_9423,N_9206);
xor U9978 (N_9978,N_8942,N_9508);
nor U9979 (N_9979,N_8815,N_9542);
nor U9980 (N_9980,N_9535,N_9151);
and U9981 (N_9981,N_9044,N_9284);
and U9982 (N_9982,N_9581,N_9333);
nor U9983 (N_9983,N_9576,N_8984);
nand U9984 (N_9984,N_8949,N_9360);
nor U9985 (N_9985,N_9037,N_9450);
or U9986 (N_9986,N_9257,N_9198);
or U9987 (N_9987,N_9077,N_9242);
nor U9988 (N_9988,N_9428,N_9407);
or U9989 (N_9989,N_9105,N_9294);
and U9990 (N_9990,N_9093,N_9013);
and U9991 (N_9991,N_9215,N_9154);
xnor U9992 (N_9992,N_9048,N_9437);
xor U9993 (N_9993,N_9405,N_8851);
xnor U9994 (N_9994,N_9330,N_8939);
xnor U9995 (N_9995,N_9514,N_9243);
nand U9996 (N_9996,N_9117,N_8850);
nor U9997 (N_9997,N_9445,N_9213);
nor U9998 (N_9998,N_9331,N_9347);
nor U9999 (N_9999,N_9402,N_9588);
or U10000 (N_10000,N_9341,N_9315);
and U10001 (N_10001,N_9340,N_9507);
or U10002 (N_10002,N_9319,N_8822);
and U10003 (N_10003,N_9048,N_9191);
xor U10004 (N_10004,N_8852,N_9419);
or U10005 (N_10005,N_9578,N_8812);
and U10006 (N_10006,N_9011,N_9096);
nand U10007 (N_10007,N_9557,N_9430);
nor U10008 (N_10008,N_9501,N_9400);
nor U10009 (N_10009,N_9258,N_9138);
and U10010 (N_10010,N_8895,N_9181);
xnor U10011 (N_10011,N_9527,N_8881);
nor U10012 (N_10012,N_9482,N_9211);
nor U10013 (N_10013,N_9184,N_9256);
or U10014 (N_10014,N_9246,N_9437);
nor U10015 (N_10015,N_8894,N_9356);
nor U10016 (N_10016,N_9062,N_9383);
nand U10017 (N_10017,N_8907,N_9402);
and U10018 (N_10018,N_8963,N_9382);
and U10019 (N_10019,N_9023,N_9142);
and U10020 (N_10020,N_9181,N_9154);
or U10021 (N_10021,N_8853,N_9005);
nor U10022 (N_10022,N_9358,N_8917);
nand U10023 (N_10023,N_8896,N_9500);
nor U10024 (N_10024,N_9099,N_9157);
or U10025 (N_10025,N_8891,N_9251);
nor U10026 (N_10026,N_9594,N_9058);
nand U10027 (N_10027,N_9218,N_9214);
and U10028 (N_10028,N_9226,N_9576);
nand U10029 (N_10029,N_8963,N_8837);
nand U10030 (N_10030,N_9047,N_9302);
xnor U10031 (N_10031,N_9249,N_8983);
nor U10032 (N_10032,N_9313,N_8897);
nand U10033 (N_10033,N_9413,N_9142);
xor U10034 (N_10034,N_9343,N_9194);
nand U10035 (N_10035,N_9304,N_8813);
and U10036 (N_10036,N_9035,N_8838);
and U10037 (N_10037,N_9009,N_8848);
nor U10038 (N_10038,N_9527,N_9086);
or U10039 (N_10039,N_9090,N_9009);
nor U10040 (N_10040,N_9300,N_9522);
nand U10041 (N_10041,N_9072,N_8824);
nor U10042 (N_10042,N_8858,N_9397);
or U10043 (N_10043,N_8948,N_9217);
nor U10044 (N_10044,N_9433,N_9009);
nand U10045 (N_10045,N_8808,N_9589);
or U10046 (N_10046,N_9165,N_9095);
nand U10047 (N_10047,N_9481,N_9324);
nand U10048 (N_10048,N_9060,N_9074);
xnor U10049 (N_10049,N_9016,N_9564);
or U10050 (N_10050,N_8835,N_8926);
or U10051 (N_10051,N_9213,N_8940);
or U10052 (N_10052,N_8940,N_9340);
xnor U10053 (N_10053,N_8917,N_9251);
nor U10054 (N_10054,N_9230,N_9507);
or U10055 (N_10055,N_9386,N_8890);
or U10056 (N_10056,N_9556,N_9411);
nor U10057 (N_10057,N_9009,N_9516);
xor U10058 (N_10058,N_9363,N_9437);
xor U10059 (N_10059,N_8940,N_9297);
or U10060 (N_10060,N_9186,N_9001);
nor U10061 (N_10061,N_9301,N_8962);
and U10062 (N_10062,N_9141,N_9034);
nand U10063 (N_10063,N_9381,N_8891);
or U10064 (N_10064,N_9327,N_9513);
or U10065 (N_10065,N_9472,N_9076);
nand U10066 (N_10066,N_8962,N_8826);
nor U10067 (N_10067,N_8803,N_9171);
nand U10068 (N_10068,N_8817,N_9368);
nor U10069 (N_10069,N_9586,N_9440);
nand U10070 (N_10070,N_9001,N_8895);
xor U10071 (N_10071,N_9087,N_9369);
nor U10072 (N_10072,N_9494,N_9043);
and U10073 (N_10073,N_9478,N_9239);
and U10074 (N_10074,N_9361,N_9487);
xor U10075 (N_10075,N_9217,N_9294);
and U10076 (N_10076,N_9134,N_8985);
xnor U10077 (N_10077,N_8835,N_8868);
xor U10078 (N_10078,N_8823,N_9057);
or U10079 (N_10079,N_9305,N_9593);
and U10080 (N_10080,N_8816,N_9279);
xnor U10081 (N_10081,N_8883,N_8956);
nor U10082 (N_10082,N_9362,N_9599);
nand U10083 (N_10083,N_9542,N_9287);
nand U10084 (N_10084,N_8878,N_9477);
or U10085 (N_10085,N_8850,N_9043);
and U10086 (N_10086,N_9330,N_8894);
or U10087 (N_10087,N_9563,N_9465);
or U10088 (N_10088,N_9144,N_9337);
nand U10089 (N_10089,N_8875,N_9126);
xor U10090 (N_10090,N_8909,N_9542);
and U10091 (N_10091,N_9425,N_9329);
nor U10092 (N_10092,N_9131,N_8905);
xor U10093 (N_10093,N_9455,N_8801);
nand U10094 (N_10094,N_9488,N_9084);
or U10095 (N_10095,N_9571,N_8976);
and U10096 (N_10096,N_9280,N_9506);
or U10097 (N_10097,N_9579,N_8801);
or U10098 (N_10098,N_9139,N_8989);
or U10099 (N_10099,N_9513,N_8994);
and U10100 (N_10100,N_9082,N_9449);
nor U10101 (N_10101,N_9509,N_9590);
nand U10102 (N_10102,N_9466,N_9393);
and U10103 (N_10103,N_8844,N_8938);
xnor U10104 (N_10104,N_9423,N_9017);
and U10105 (N_10105,N_8927,N_9296);
nor U10106 (N_10106,N_8849,N_9125);
and U10107 (N_10107,N_9155,N_9309);
nor U10108 (N_10108,N_9378,N_9532);
nand U10109 (N_10109,N_9010,N_9276);
or U10110 (N_10110,N_9492,N_9528);
nand U10111 (N_10111,N_9085,N_9261);
xnor U10112 (N_10112,N_9538,N_9301);
xnor U10113 (N_10113,N_9327,N_8970);
and U10114 (N_10114,N_9242,N_8872);
nor U10115 (N_10115,N_9098,N_8916);
and U10116 (N_10116,N_8917,N_8874);
nor U10117 (N_10117,N_9512,N_9490);
and U10118 (N_10118,N_8909,N_8890);
nor U10119 (N_10119,N_9380,N_9061);
xnor U10120 (N_10120,N_9196,N_8800);
xnor U10121 (N_10121,N_8903,N_8827);
nor U10122 (N_10122,N_9155,N_9436);
nand U10123 (N_10123,N_9385,N_9011);
and U10124 (N_10124,N_9306,N_9348);
or U10125 (N_10125,N_9002,N_9565);
xnor U10126 (N_10126,N_8971,N_8853);
and U10127 (N_10127,N_9360,N_9133);
and U10128 (N_10128,N_9212,N_8831);
nand U10129 (N_10129,N_9229,N_9518);
and U10130 (N_10130,N_9337,N_8996);
xnor U10131 (N_10131,N_9065,N_9459);
nor U10132 (N_10132,N_8921,N_9512);
xor U10133 (N_10133,N_9302,N_9169);
xnor U10134 (N_10134,N_9395,N_9330);
or U10135 (N_10135,N_9159,N_9359);
or U10136 (N_10136,N_9418,N_9187);
nand U10137 (N_10137,N_9014,N_9196);
nor U10138 (N_10138,N_9558,N_9056);
xnor U10139 (N_10139,N_9153,N_9043);
xnor U10140 (N_10140,N_8826,N_9511);
or U10141 (N_10141,N_9593,N_8815);
nor U10142 (N_10142,N_9425,N_9244);
and U10143 (N_10143,N_9060,N_9299);
or U10144 (N_10144,N_9591,N_9006);
nor U10145 (N_10145,N_9052,N_9390);
nand U10146 (N_10146,N_9184,N_9575);
nor U10147 (N_10147,N_9503,N_9178);
xor U10148 (N_10148,N_9431,N_8803);
nor U10149 (N_10149,N_9042,N_9250);
xor U10150 (N_10150,N_8995,N_9448);
nand U10151 (N_10151,N_9059,N_9173);
or U10152 (N_10152,N_9180,N_9291);
nand U10153 (N_10153,N_8921,N_9406);
xnor U10154 (N_10154,N_9375,N_9327);
and U10155 (N_10155,N_8923,N_9245);
or U10156 (N_10156,N_9204,N_9060);
or U10157 (N_10157,N_8820,N_8826);
or U10158 (N_10158,N_8978,N_9156);
xor U10159 (N_10159,N_8914,N_9279);
and U10160 (N_10160,N_9014,N_9326);
nor U10161 (N_10161,N_8840,N_9406);
nor U10162 (N_10162,N_8879,N_9395);
xnor U10163 (N_10163,N_9589,N_8904);
or U10164 (N_10164,N_9311,N_9301);
or U10165 (N_10165,N_9047,N_8814);
nand U10166 (N_10166,N_9422,N_9181);
nand U10167 (N_10167,N_9226,N_9480);
and U10168 (N_10168,N_9035,N_9186);
or U10169 (N_10169,N_9168,N_9417);
xnor U10170 (N_10170,N_8829,N_9340);
nor U10171 (N_10171,N_9386,N_8847);
nand U10172 (N_10172,N_9564,N_9413);
or U10173 (N_10173,N_8807,N_9012);
xnor U10174 (N_10174,N_9175,N_8809);
xor U10175 (N_10175,N_9569,N_9207);
and U10176 (N_10176,N_9313,N_9222);
nand U10177 (N_10177,N_9505,N_9553);
nand U10178 (N_10178,N_9230,N_9223);
xor U10179 (N_10179,N_8908,N_9494);
xor U10180 (N_10180,N_8824,N_9289);
or U10181 (N_10181,N_8881,N_9289);
and U10182 (N_10182,N_9507,N_9082);
or U10183 (N_10183,N_9124,N_9178);
xnor U10184 (N_10184,N_9202,N_8986);
nor U10185 (N_10185,N_9352,N_9426);
or U10186 (N_10186,N_9432,N_9156);
nand U10187 (N_10187,N_9458,N_8936);
or U10188 (N_10188,N_8868,N_8848);
xnor U10189 (N_10189,N_9240,N_9116);
nand U10190 (N_10190,N_8860,N_9580);
nor U10191 (N_10191,N_9236,N_9181);
xor U10192 (N_10192,N_9341,N_9048);
nor U10193 (N_10193,N_8952,N_9259);
or U10194 (N_10194,N_9349,N_9397);
nand U10195 (N_10195,N_8966,N_9445);
and U10196 (N_10196,N_9408,N_9235);
and U10197 (N_10197,N_9242,N_9587);
nor U10198 (N_10198,N_9345,N_8978);
xnor U10199 (N_10199,N_9042,N_9530);
nand U10200 (N_10200,N_9556,N_9525);
or U10201 (N_10201,N_9493,N_9504);
and U10202 (N_10202,N_9487,N_8892);
xnor U10203 (N_10203,N_9422,N_9230);
nand U10204 (N_10204,N_8929,N_8879);
nand U10205 (N_10205,N_8878,N_8895);
or U10206 (N_10206,N_9583,N_8975);
nor U10207 (N_10207,N_9154,N_8825);
nand U10208 (N_10208,N_9086,N_9569);
or U10209 (N_10209,N_9119,N_9172);
or U10210 (N_10210,N_8866,N_8974);
or U10211 (N_10211,N_9393,N_9113);
or U10212 (N_10212,N_9122,N_8827);
nor U10213 (N_10213,N_8960,N_9240);
nor U10214 (N_10214,N_8915,N_9433);
or U10215 (N_10215,N_8904,N_8977);
xor U10216 (N_10216,N_9029,N_9023);
xnor U10217 (N_10217,N_9563,N_9190);
and U10218 (N_10218,N_8981,N_9450);
xor U10219 (N_10219,N_9321,N_9208);
and U10220 (N_10220,N_9056,N_9247);
nor U10221 (N_10221,N_9357,N_8896);
nand U10222 (N_10222,N_9102,N_9376);
and U10223 (N_10223,N_9133,N_9071);
nor U10224 (N_10224,N_8885,N_9285);
nand U10225 (N_10225,N_9446,N_9489);
or U10226 (N_10226,N_8958,N_9126);
nor U10227 (N_10227,N_8858,N_9015);
and U10228 (N_10228,N_8875,N_9045);
and U10229 (N_10229,N_8984,N_9127);
xor U10230 (N_10230,N_8860,N_9040);
or U10231 (N_10231,N_8861,N_9204);
nand U10232 (N_10232,N_9289,N_9511);
nand U10233 (N_10233,N_8878,N_8915);
xnor U10234 (N_10234,N_8988,N_9280);
or U10235 (N_10235,N_9530,N_9006);
xnor U10236 (N_10236,N_9493,N_9390);
nor U10237 (N_10237,N_9352,N_9272);
xnor U10238 (N_10238,N_9203,N_9572);
xnor U10239 (N_10239,N_9176,N_9337);
nand U10240 (N_10240,N_8966,N_9224);
nand U10241 (N_10241,N_9163,N_9365);
xnor U10242 (N_10242,N_9030,N_9361);
and U10243 (N_10243,N_8967,N_9281);
nor U10244 (N_10244,N_9144,N_9240);
nand U10245 (N_10245,N_9256,N_9065);
and U10246 (N_10246,N_9371,N_8875);
and U10247 (N_10247,N_9438,N_9473);
nand U10248 (N_10248,N_9052,N_9457);
nand U10249 (N_10249,N_9185,N_8942);
nand U10250 (N_10250,N_8904,N_9524);
or U10251 (N_10251,N_9326,N_9305);
or U10252 (N_10252,N_9504,N_9553);
nand U10253 (N_10253,N_8927,N_9027);
nand U10254 (N_10254,N_9028,N_9260);
nor U10255 (N_10255,N_9189,N_9555);
or U10256 (N_10256,N_8819,N_9201);
nand U10257 (N_10257,N_8842,N_9504);
xnor U10258 (N_10258,N_9257,N_9247);
or U10259 (N_10259,N_9414,N_9097);
or U10260 (N_10260,N_8971,N_9052);
and U10261 (N_10261,N_9384,N_9449);
nor U10262 (N_10262,N_8870,N_9013);
or U10263 (N_10263,N_9526,N_9230);
nand U10264 (N_10264,N_9069,N_9423);
xor U10265 (N_10265,N_9289,N_9590);
nor U10266 (N_10266,N_9143,N_9514);
nor U10267 (N_10267,N_9471,N_9159);
nand U10268 (N_10268,N_9412,N_8825);
or U10269 (N_10269,N_9419,N_9049);
or U10270 (N_10270,N_8858,N_8847);
xnor U10271 (N_10271,N_9371,N_9384);
nor U10272 (N_10272,N_8947,N_9242);
nand U10273 (N_10273,N_8876,N_9592);
and U10274 (N_10274,N_9447,N_8817);
and U10275 (N_10275,N_8937,N_9420);
or U10276 (N_10276,N_8949,N_9414);
or U10277 (N_10277,N_8815,N_9096);
or U10278 (N_10278,N_9498,N_9201);
or U10279 (N_10279,N_9526,N_8845);
and U10280 (N_10280,N_9326,N_9555);
nand U10281 (N_10281,N_9054,N_9294);
and U10282 (N_10282,N_9519,N_9003);
nand U10283 (N_10283,N_8960,N_9473);
xnor U10284 (N_10284,N_9167,N_8864);
nor U10285 (N_10285,N_8972,N_9080);
xor U10286 (N_10286,N_9216,N_8876);
nor U10287 (N_10287,N_8862,N_9423);
or U10288 (N_10288,N_9336,N_9546);
and U10289 (N_10289,N_8853,N_8842);
xnor U10290 (N_10290,N_9487,N_9246);
or U10291 (N_10291,N_9357,N_9049);
nor U10292 (N_10292,N_9517,N_9274);
nand U10293 (N_10293,N_9551,N_9539);
xor U10294 (N_10294,N_9230,N_9490);
xnor U10295 (N_10295,N_9380,N_8860);
or U10296 (N_10296,N_9452,N_9281);
xor U10297 (N_10297,N_8806,N_9072);
and U10298 (N_10298,N_9094,N_9354);
nor U10299 (N_10299,N_9115,N_9596);
nand U10300 (N_10300,N_9162,N_8850);
nand U10301 (N_10301,N_9589,N_9585);
nand U10302 (N_10302,N_8957,N_8903);
nand U10303 (N_10303,N_8983,N_9392);
and U10304 (N_10304,N_9370,N_9177);
xor U10305 (N_10305,N_9213,N_9438);
and U10306 (N_10306,N_9142,N_9259);
or U10307 (N_10307,N_8963,N_8875);
or U10308 (N_10308,N_8942,N_8911);
and U10309 (N_10309,N_9271,N_9173);
and U10310 (N_10310,N_8998,N_8819);
or U10311 (N_10311,N_9000,N_8933);
nor U10312 (N_10312,N_8846,N_8990);
and U10313 (N_10313,N_9258,N_9000);
nor U10314 (N_10314,N_9316,N_9518);
and U10315 (N_10315,N_9161,N_9074);
or U10316 (N_10316,N_9540,N_9396);
and U10317 (N_10317,N_9455,N_9219);
nor U10318 (N_10318,N_9562,N_9475);
nor U10319 (N_10319,N_9226,N_9121);
nor U10320 (N_10320,N_8803,N_9068);
and U10321 (N_10321,N_9275,N_8842);
nand U10322 (N_10322,N_9332,N_9135);
nand U10323 (N_10323,N_8816,N_9068);
nand U10324 (N_10324,N_8980,N_8852);
and U10325 (N_10325,N_9241,N_9085);
nand U10326 (N_10326,N_9497,N_9051);
or U10327 (N_10327,N_9557,N_9365);
xnor U10328 (N_10328,N_8839,N_8915);
xnor U10329 (N_10329,N_9239,N_9102);
nand U10330 (N_10330,N_9412,N_9335);
nand U10331 (N_10331,N_9416,N_9057);
nand U10332 (N_10332,N_9178,N_8841);
and U10333 (N_10333,N_9067,N_9107);
nor U10334 (N_10334,N_8917,N_9340);
xnor U10335 (N_10335,N_9244,N_9279);
nor U10336 (N_10336,N_9388,N_8849);
nand U10337 (N_10337,N_9514,N_9594);
nor U10338 (N_10338,N_9327,N_9516);
nor U10339 (N_10339,N_8881,N_9033);
nand U10340 (N_10340,N_9383,N_9255);
nand U10341 (N_10341,N_9213,N_8804);
xor U10342 (N_10342,N_9530,N_9154);
xnor U10343 (N_10343,N_9529,N_9017);
and U10344 (N_10344,N_8998,N_9197);
nand U10345 (N_10345,N_9562,N_9462);
nand U10346 (N_10346,N_9161,N_9370);
nand U10347 (N_10347,N_9010,N_8994);
nand U10348 (N_10348,N_9540,N_8815);
xnor U10349 (N_10349,N_8874,N_9010);
and U10350 (N_10350,N_9214,N_8933);
nand U10351 (N_10351,N_9011,N_9121);
xor U10352 (N_10352,N_9184,N_8809);
xor U10353 (N_10353,N_9454,N_9272);
xor U10354 (N_10354,N_8887,N_9426);
nor U10355 (N_10355,N_9130,N_9499);
nand U10356 (N_10356,N_9147,N_8838);
xnor U10357 (N_10357,N_9067,N_8909);
or U10358 (N_10358,N_9056,N_8869);
nor U10359 (N_10359,N_8941,N_8931);
or U10360 (N_10360,N_9321,N_8894);
or U10361 (N_10361,N_9437,N_9294);
and U10362 (N_10362,N_8922,N_9167);
nor U10363 (N_10363,N_9514,N_9270);
xor U10364 (N_10364,N_9406,N_9372);
xnor U10365 (N_10365,N_9284,N_9462);
xor U10366 (N_10366,N_9107,N_9495);
or U10367 (N_10367,N_9404,N_9050);
or U10368 (N_10368,N_9062,N_8809);
xor U10369 (N_10369,N_9463,N_9540);
and U10370 (N_10370,N_9058,N_9387);
or U10371 (N_10371,N_8918,N_9150);
and U10372 (N_10372,N_9084,N_9495);
or U10373 (N_10373,N_9023,N_9416);
nor U10374 (N_10374,N_9478,N_9291);
nor U10375 (N_10375,N_9215,N_9157);
nor U10376 (N_10376,N_9229,N_8940);
and U10377 (N_10377,N_9301,N_8828);
and U10378 (N_10378,N_9162,N_9590);
nor U10379 (N_10379,N_9478,N_9547);
and U10380 (N_10380,N_9019,N_8819);
nand U10381 (N_10381,N_9237,N_8864);
xnor U10382 (N_10382,N_8846,N_9222);
and U10383 (N_10383,N_8909,N_9270);
and U10384 (N_10384,N_9080,N_9157);
or U10385 (N_10385,N_9230,N_9284);
or U10386 (N_10386,N_9096,N_9325);
nand U10387 (N_10387,N_8871,N_9599);
xnor U10388 (N_10388,N_9210,N_9587);
nor U10389 (N_10389,N_9274,N_9012);
nand U10390 (N_10390,N_8815,N_9107);
nand U10391 (N_10391,N_9108,N_9159);
nand U10392 (N_10392,N_8998,N_8876);
nand U10393 (N_10393,N_9348,N_9555);
xnor U10394 (N_10394,N_9451,N_9456);
or U10395 (N_10395,N_9023,N_9470);
nor U10396 (N_10396,N_9303,N_9548);
or U10397 (N_10397,N_8908,N_9045);
and U10398 (N_10398,N_9436,N_8933);
nor U10399 (N_10399,N_9043,N_8908);
nand U10400 (N_10400,N_10079,N_9779);
nand U10401 (N_10401,N_10281,N_10297);
xor U10402 (N_10402,N_9989,N_9631);
and U10403 (N_10403,N_9661,N_10019);
nand U10404 (N_10404,N_9956,N_10090);
xnor U10405 (N_10405,N_9942,N_10046);
or U10406 (N_10406,N_9608,N_9884);
and U10407 (N_10407,N_10132,N_10384);
nand U10408 (N_10408,N_10073,N_9890);
nand U10409 (N_10409,N_10306,N_10372);
nand U10410 (N_10410,N_9792,N_9704);
nor U10411 (N_10411,N_10258,N_9717);
nand U10412 (N_10412,N_9778,N_10088);
or U10413 (N_10413,N_9943,N_9684);
and U10414 (N_10414,N_10111,N_9851);
nor U10415 (N_10415,N_10315,N_9782);
or U10416 (N_10416,N_10373,N_9690);
nand U10417 (N_10417,N_10193,N_10244);
or U10418 (N_10418,N_9655,N_10291);
nand U10419 (N_10419,N_9692,N_9862);
nand U10420 (N_10420,N_10093,N_9856);
nand U10421 (N_10421,N_10380,N_10135);
and U10422 (N_10422,N_9848,N_10217);
nand U10423 (N_10423,N_10230,N_10322);
nand U10424 (N_10424,N_9694,N_10148);
nand U10425 (N_10425,N_9858,N_10238);
nor U10426 (N_10426,N_9986,N_10105);
and U10427 (N_10427,N_10374,N_9997);
xor U10428 (N_10428,N_9893,N_9695);
nand U10429 (N_10429,N_10245,N_9955);
xnor U10430 (N_10430,N_10350,N_9909);
nand U10431 (N_10431,N_9828,N_9727);
or U10432 (N_10432,N_9747,N_10303);
and U10433 (N_10433,N_10299,N_10390);
and U10434 (N_10434,N_10052,N_9861);
xor U10435 (N_10435,N_10136,N_9895);
xor U10436 (N_10436,N_10359,N_9816);
or U10437 (N_10437,N_9677,N_9983);
and U10438 (N_10438,N_9801,N_9847);
xnor U10439 (N_10439,N_10164,N_10080);
or U10440 (N_10440,N_10176,N_10298);
or U10441 (N_10441,N_10273,N_9836);
nor U10442 (N_10442,N_10199,N_9889);
xor U10443 (N_10443,N_9662,N_10386);
nand U10444 (N_10444,N_10369,N_10159);
nor U10445 (N_10445,N_10066,N_10234);
xnor U10446 (N_10446,N_10127,N_9953);
nor U10447 (N_10447,N_10048,N_10331);
nand U10448 (N_10448,N_9671,N_9645);
or U10449 (N_10449,N_9870,N_9991);
or U10450 (N_10450,N_9627,N_9680);
nor U10451 (N_10451,N_9756,N_10030);
or U10452 (N_10452,N_10357,N_10361);
nor U10453 (N_10453,N_10006,N_10107);
xor U10454 (N_10454,N_9927,N_9971);
nand U10455 (N_10455,N_10292,N_10186);
xor U10456 (N_10456,N_10077,N_10279);
nor U10457 (N_10457,N_9970,N_9979);
xor U10458 (N_10458,N_10190,N_9935);
xor U10459 (N_10459,N_9740,N_9961);
xor U10460 (N_10460,N_9881,N_10340);
and U10461 (N_10461,N_10116,N_10059);
nand U10462 (N_10462,N_9984,N_9839);
or U10463 (N_10463,N_9741,N_10023);
nor U10464 (N_10464,N_9910,N_10293);
xnor U10465 (N_10465,N_9886,N_9622);
nand U10466 (N_10466,N_10276,N_10389);
nor U10467 (N_10467,N_9761,N_9749);
nand U10468 (N_10468,N_10069,N_9688);
xnor U10469 (N_10469,N_9771,N_9777);
or U10470 (N_10470,N_9738,N_10326);
nor U10471 (N_10471,N_10287,N_9606);
or U10472 (N_10472,N_10047,N_10086);
nor U10473 (N_10473,N_10057,N_10318);
nor U10474 (N_10474,N_9911,N_9874);
xor U10475 (N_10475,N_10197,N_9745);
or U10476 (N_10476,N_10010,N_10356);
and U10477 (N_10477,N_10064,N_9674);
nor U10478 (N_10478,N_10041,N_10165);
or U10479 (N_10479,N_10145,N_10202);
nand U10480 (N_10480,N_10074,N_10203);
nand U10481 (N_10481,N_9826,N_9638);
and U10482 (N_10482,N_9999,N_10260);
nand U10483 (N_10483,N_9744,N_9652);
xor U10484 (N_10484,N_10108,N_10339);
nor U10485 (N_10485,N_9678,N_10209);
and U10486 (N_10486,N_9748,N_10115);
nand U10487 (N_10487,N_9885,N_9940);
and U10488 (N_10488,N_9743,N_9985);
and U10489 (N_10489,N_9954,N_10128);
nand U10490 (N_10490,N_9876,N_9959);
nand U10491 (N_10491,N_9775,N_10255);
nor U10492 (N_10492,N_9706,N_10087);
xor U10493 (N_10493,N_9992,N_9710);
or U10494 (N_10494,N_9952,N_9683);
nand U10495 (N_10495,N_9835,N_9859);
nand U10496 (N_10496,N_9648,N_9987);
and U10497 (N_10497,N_10268,N_9716);
nor U10498 (N_10498,N_10257,N_9863);
and U10499 (N_10499,N_9797,N_10348);
or U10500 (N_10500,N_10101,N_9900);
nand U10501 (N_10501,N_10321,N_10329);
nor U10502 (N_10502,N_9903,N_9894);
and U10503 (N_10503,N_9994,N_9619);
nor U10504 (N_10504,N_9819,N_9702);
and U10505 (N_10505,N_9791,N_10347);
nand U10506 (N_10506,N_9823,N_10335);
nand U10507 (N_10507,N_9672,N_9875);
or U10508 (N_10508,N_9735,N_9921);
and U10509 (N_10509,N_10252,N_10133);
or U10510 (N_10510,N_9917,N_10017);
nor U10511 (N_10511,N_10024,N_10168);
and U10512 (N_10512,N_10031,N_9718);
and U10513 (N_10513,N_9646,N_10126);
xor U10514 (N_10514,N_9613,N_9629);
nand U10515 (N_10515,N_10214,N_9902);
xnor U10516 (N_10516,N_10366,N_9887);
nor U10517 (N_10517,N_9751,N_9905);
xnor U10518 (N_10518,N_10343,N_10185);
xor U10519 (N_10519,N_9603,N_9669);
and U10520 (N_10520,N_10143,N_9636);
or U10521 (N_10521,N_9867,N_10235);
or U10522 (N_10522,N_9762,N_10063);
nor U10523 (N_10523,N_9809,N_9611);
or U10524 (N_10524,N_9794,N_9604);
nor U10525 (N_10525,N_9705,N_9676);
nor U10526 (N_10526,N_9939,N_10289);
or U10527 (N_10527,N_10387,N_9929);
and U10528 (N_10528,N_10316,N_9981);
nand U10529 (N_10529,N_9708,N_9980);
nand U10530 (N_10530,N_9691,N_9844);
and U10531 (N_10531,N_10313,N_10177);
or U10532 (N_10532,N_10078,N_9947);
and U10533 (N_10533,N_10237,N_10095);
nand U10534 (N_10534,N_10242,N_10137);
nor U10535 (N_10535,N_10324,N_10033);
nor U10536 (N_10536,N_10084,N_9898);
nor U10537 (N_10537,N_9786,N_10210);
xnor U10538 (N_10538,N_9620,N_10042);
and U10539 (N_10539,N_10034,N_10249);
or U10540 (N_10540,N_9776,N_10007);
xor U10541 (N_10541,N_10266,N_10198);
xnor U10542 (N_10542,N_10188,N_9643);
nand U10543 (N_10543,N_9830,N_10302);
or U10544 (N_10544,N_10312,N_9944);
or U10545 (N_10545,N_10354,N_10004);
or U10546 (N_10546,N_10375,N_9736);
nor U10547 (N_10547,N_9896,N_9995);
and U10548 (N_10548,N_10385,N_10008);
nand U10549 (N_10549,N_10001,N_10091);
and U10550 (N_10550,N_9746,N_9649);
nor U10551 (N_10551,N_9937,N_10263);
xnor U10552 (N_10552,N_10157,N_10227);
nor U10553 (N_10553,N_9617,N_9864);
nor U10554 (N_10554,N_10000,N_9628);
nor U10555 (N_10555,N_10345,N_9637);
or U10556 (N_10556,N_9770,N_9855);
nand U10557 (N_10557,N_9803,N_10365);
xor U10558 (N_10558,N_9721,N_9998);
xor U10559 (N_10559,N_10060,N_9854);
nor U10560 (N_10560,N_10204,N_9891);
and U10561 (N_10561,N_9789,N_9882);
nor U10562 (N_10562,N_10261,N_10005);
and U10563 (N_10563,N_9968,N_9988);
or U10564 (N_10564,N_9610,N_10044);
xnor U10565 (N_10565,N_10028,N_10212);
and U10566 (N_10566,N_9838,N_9774);
nand U10567 (N_10567,N_9825,N_9635);
nand U10568 (N_10568,N_10243,N_10098);
xor U10569 (N_10569,N_10355,N_10222);
or U10570 (N_10570,N_9977,N_9820);
or U10571 (N_10571,N_9714,N_9877);
nand U10572 (N_10572,N_10120,N_10224);
or U10573 (N_10573,N_9908,N_10391);
xor U10574 (N_10574,N_10219,N_10265);
or U10575 (N_10575,N_9897,N_10179);
or U10576 (N_10576,N_10392,N_9696);
or U10577 (N_10577,N_10262,N_9679);
and U10578 (N_10578,N_9703,N_9616);
xnor U10579 (N_10579,N_9934,N_10039);
xnor U10580 (N_10580,N_10134,N_10036);
nand U10581 (N_10581,N_10274,N_9842);
nand U10582 (N_10582,N_9852,N_10320);
and U10583 (N_10583,N_9922,N_9760);
nor U10584 (N_10584,N_9883,N_10184);
nand U10585 (N_10585,N_9633,N_10332);
nand U10586 (N_10586,N_10172,N_10141);
xor U10587 (N_10587,N_10067,N_10393);
nand U10588 (N_10588,N_10123,N_10351);
and U10589 (N_10589,N_10162,N_10275);
xor U10590 (N_10590,N_10038,N_9713);
nor U10591 (N_10591,N_10323,N_10360);
or U10592 (N_10592,N_9664,N_10027);
xor U10593 (N_10593,N_9879,N_9682);
nand U10594 (N_10594,N_9798,N_9615);
nor U10595 (N_10595,N_10267,N_10341);
or U10596 (N_10596,N_10352,N_9958);
xor U10597 (N_10597,N_10022,N_10149);
nand U10598 (N_10598,N_9918,N_10140);
nand U10599 (N_10599,N_10112,N_9681);
nor U10600 (N_10600,N_9769,N_9621);
nand U10601 (N_10601,N_10200,N_10294);
and U10602 (N_10602,N_9693,N_10085);
or U10603 (N_10603,N_9966,N_10013);
and U10604 (N_10604,N_10029,N_9753);
nand U10605 (N_10605,N_9719,N_10284);
xor U10606 (N_10606,N_10037,N_9765);
nand U10607 (N_10607,N_10208,N_10388);
xor U10608 (N_10608,N_9609,N_10353);
nand U10609 (N_10609,N_9697,N_9673);
and U10610 (N_10610,N_10364,N_9860);
nand U10611 (N_10611,N_10271,N_9624);
xnor U10612 (N_10612,N_9667,N_10158);
nor U10613 (N_10613,N_10122,N_9892);
or U10614 (N_10614,N_10015,N_9871);
and U10615 (N_10615,N_10307,N_9960);
or U10616 (N_10616,N_9846,N_9853);
nand U10617 (N_10617,N_10110,N_10102);
or U10618 (N_10618,N_10109,N_10121);
nand U10619 (N_10619,N_9783,N_10003);
and U10620 (N_10620,N_10070,N_9764);
and U10621 (N_10621,N_9759,N_9899);
xnor U10622 (N_10622,N_10216,N_10035);
or U10623 (N_10623,N_10377,N_9666);
xnor U10624 (N_10624,N_9730,N_9701);
xor U10625 (N_10625,N_9601,N_10304);
or U10626 (N_10626,N_9907,N_10083);
nand U10627 (N_10627,N_9781,N_9707);
and U10628 (N_10628,N_10282,N_10251);
nand U10629 (N_10629,N_9837,N_9811);
or U10630 (N_10630,N_10213,N_9930);
xnor U10631 (N_10631,N_10223,N_10218);
xnor U10632 (N_10632,N_9685,N_10072);
nand U10633 (N_10633,N_10328,N_10338);
nand U10634 (N_10634,N_10280,N_10269);
xnor U10635 (N_10635,N_9993,N_10192);
nor U10636 (N_10636,N_10175,N_10337);
or U10637 (N_10637,N_10075,N_9967);
and U10638 (N_10638,N_9951,N_9878);
and U10639 (N_10639,N_10272,N_10049);
nand U10640 (N_10640,N_10398,N_10317);
nor U10641 (N_10641,N_9623,N_10183);
or U10642 (N_10642,N_10205,N_9651);
and U10643 (N_10643,N_10082,N_10016);
or U10644 (N_10644,N_9787,N_9654);
xnor U10645 (N_10645,N_9928,N_10114);
nor U10646 (N_10646,N_9700,N_10290);
or U10647 (N_10647,N_9656,N_10233);
and U10648 (N_10648,N_10288,N_9602);
nand U10649 (N_10649,N_9817,N_10300);
and U10650 (N_10650,N_10113,N_9768);
and U10651 (N_10651,N_9709,N_10191);
nand U10652 (N_10652,N_9924,N_10187);
or U10653 (N_10653,N_10173,N_9849);
nand U10654 (N_10654,N_10100,N_10146);
or U10655 (N_10655,N_9919,N_10119);
nand U10656 (N_10656,N_10383,N_10014);
xor U10657 (N_10657,N_10189,N_9640);
nor U10658 (N_10658,N_9824,N_10215);
or U10659 (N_10659,N_10104,N_9634);
nor U10660 (N_10660,N_9686,N_9923);
nand U10661 (N_10661,N_9866,N_9969);
nor U10662 (N_10662,N_9818,N_10254);
or U10663 (N_10663,N_9614,N_10256);
or U10664 (N_10664,N_10081,N_9873);
or U10665 (N_10665,N_10096,N_10248);
xor U10666 (N_10666,N_10076,N_9600);
xnor U10667 (N_10667,N_9796,N_9653);
nor U10668 (N_10668,N_9804,N_9822);
or U10669 (N_10669,N_9632,N_10270);
xnor U10670 (N_10670,N_10117,N_10394);
and U10671 (N_10671,N_9869,N_10139);
nor U10672 (N_10672,N_9806,N_9843);
xor U10673 (N_10673,N_9974,N_10363);
nor U10674 (N_10674,N_9799,N_9945);
nand U10675 (N_10675,N_10068,N_9904);
xor U10676 (N_10676,N_10206,N_9689);
or U10677 (N_10677,N_9880,N_10285);
nand U10678 (N_10678,N_9933,N_10160);
or U10679 (N_10679,N_9964,N_10278);
or U10680 (N_10680,N_9813,N_10319);
nand U10681 (N_10681,N_10232,N_9742);
or U10682 (N_10682,N_9766,N_9990);
and U10683 (N_10683,N_9773,N_10362);
and U10684 (N_10684,N_9687,N_10368);
and U10685 (N_10685,N_10043,N_10050);
or U10686 (N_10686,N_9641,N_9865);
xor U10687 (N_10687,N_9785,N_10178);
and U10688 (N_10688,N_9965,N_10381);
xor U10689 (N_10689,N_10045,N_10296);
nor U10690 (N_10690,N_9829,N_9931);
nor U10691 (N_10691,N_10026,N_9888);
xor U10692 (N_10692,N_10062,N_10283);
and U10693 (N_10693,N_9805,N_10131);
xor U10694 (N_10694,N_10147,N_10138);
xor U10695 (N_10695,N_9914,N_10310);
xor U10696 (N_10696,N_10247,N_9868);
and U10697 (N_10697,N_10056,N_10211);
nand U10698 (N_10698,N_9639,N_10395);
nand U10699 (N_10699,N_10396,N_9800);
or U10700 (N_10700,N_10253,N_10378);
nand U10701 (N_10701,N_10195,N_9936);
and U10702 (N_10702,N_10055,N_9650);
and U10703 (N_10703,N_9767,N_10171);
and U10704 (N_10704,N_9647,N_9938);
or U10705 (N_10705,N_10229,N_10002);
and U10706 (N_10706,N_10161,N_10152);
or U10707 (N_10707,N_10065,N_9946);
nand U10708 (N_10708,N_10012,N_10336);
and U10709 (N_10709,N_9833,N_9975);
and U10710 (N_10710,N_9626,N_9723);
nand U10711 (N_10711,N_9763,N_9807);
and U10712 (N_10712,N_10376,N_9831);
nor U10713 (N_10713,N_10330,N_9726);
nor U10714 (N_10714,N_10325,N_9739);
or U10715 (N_10715,N_10239,N_10106);
nor U10716 (N_10716,N_10311,N_10308);
or U10717 (N_10717,N_9976,N_10166);
or U10718 (N_10718,N_9784,N_10220);
nor U10719 (N_10719,N_9788,N_10301);
and U10720 (N_10720,N_10314,N_9642);
and U10721 (N_10721,N_10124,N_9957);
nand U10722 (N_10722,N_9750,N_9660);
and U10723 (N_10723,N_10379,N_10250);
and U10724 (N_10724,N_10032,N_9630);
nor U10725 (N_10725,N_10151,N_9722);
xnor U10726 (N_10726,N_10144,N_10103);
nor U10727 (N_10727,N_9857,N_10349);
nor U10728 (N_10728,N_9802,N_9978);
nand U10729 (N_10729,N_9644,N_9926);
nor U10730 (N_10730,N_9618,N_10011);
nand U10731 (N_10731,N_10153,N_10201);
or U10732 (N_10732,N_9737,N_10156);
nor U10733 (N_10733,N_9841,N_10231);
nor U10734 (N_10734,N_9732,N_9605);
xnor U10735 (N_10735,N_10053,N_10236);
nor U10736 (N_10736,N_9752,N_9913);
nor U10737 (N_10737,N_9658,N_10094);
nand U10738 (N_10738,N_10382,N_10344);
xnor U10739 (N_10739,N_9872,N_10327);
nand U10740 (N_10740,N_10009,N_10163);
and U10741 (N_10741,N_9810,N_9972);
xnor U10742 (N_10742,N_10358,N_9941);
or U10743 (N_10743,N_10241,N_10018);
nand U10744 (N_10744,N_10342,N_9698);
xor U10745 (N_10745,N_10170,N_9657);
or U10746 (N_10746,N_10089,N_10099);
nand U10747 (N_10747,N_9901,N_9757);
xnor U10748 (N_10748,N_9668,N_10054);
or U10749 (N_10749,N_10021,N_9612);
or U10750 (N_10750,N_10155,N_9920);
and U10751 (N_10751,N_10167,N_9670);
and U10752 (N_10752,N_9720,N_9724);
and U10753 (N_10753,N_10371,N_9915);
nand U10754 (N_10754,N_9731,N_10071);
or U10755 (N_10755,N_10174,N_10295);
xnor U10756 (N_10756,N_10226,N_9906);
nor U10757 (N_10757,N_10154,N_10221);
or U10758 (N_10758,N_9996,N_9827);
or U10759 (N_10759,N_10305,N_9815);
and U10760 (N_10760,N_9754,N_10346);
xor U10761 (N_10761,N_9850,N_9780);
xor U10762 (N_10762,N_10058,N_9982);
nor U10763 (N_10763,N_10181,N_9821);
nand U10764 (N_10764,N_10246,N_9733);
nand U10765 (N_10765,N_9949,N_9728);
xor U10766 (N_10766,N_9665,N_9725);
nand U10767 (N_10767,N_10040,N_9948);
xor U10768 (N_10768,N_9912,N_9758);
xor U10769 (N_10769,N_10334,N_9916);
or U10770 (N_10770,N_9963,N_9711);
or U10771 (N_10771,N_10225,N_10196);
nand U10772 (N_10772,N_10367,N_9675);
and U10773 (N_10773,N_10333,N_9845);
and U10774 (N_10774,N_10020,N_10097);
xnor U10775 (N_10775,N_9793,N_10207);
xor U10776 (N_10776,N_9812,N_9663);
xor U10777 (N_10777,N_10264,N_10240);
xnor U10778 (N_10778,N_9808,N_9832);
nor U10779 (N_10779,N_10025,N_10182);
nor U10780 (N_10780,N_10180,N_10092);
nand U10781 (N_10781,N_9840,N_9715);
or U10782 (N_10782,N_9734,N_9790);
xnor U10783 (N_10783,N_10370,N_10228);
and U10784 (N_10784,N_10150,N_9625);
nor U10785 (N_10785,N_9925,N_10259);
nand U10786 (N_10786,N_10125,N_9712);
nand U10787 (N_10787,N_10130,N_10118);
nor U10788 (N_10788,N_10397,N_9607);
nor U10789 (N_10789,N_9772,N_10194);
and U10790 (N_10790,N_10061,N_9755);
nand U10791 (N_10791,N_10309,N_9659);
nor U10792 (N_10792,N_9932,N_9962);
nand U10793 (N_10793,N_10399,N_10142);
and U10794 (N_10794,N_10051,N_9699);
nand U10795 (N_10795,N_10169,N_10286);
nand U10796 (N_10796,N_9973,N_9950);
xor U10797 (N_10797,N_9814,N_10277);
nor U10798 (N_10798,N_9795,N_9834);
xor U10799 (N_10799,N_9729,N_10129);
nor U10800 (N_10800,N_10340,N_10046);
or U10801 (N_10801,N_10102,N_10241);
nor U10802 (N_10802,N_10011,N_9771);
xor U10803 (N_10803,N_9960,N_10036);
nor U10804 (N_10804,N_10249,N_9711);
nand U10805 (N_10805,N_9905,N_9947);
and U10806 (N_10806,N_9939,N_9931);
xor U10807 (N_10807,N_9629,N_9739);
and U10808 (N_10808,N_10031,N_10278);
and U10809 (N_10809,N_9989,N_10253);
nor U10810 (N_10810,N_9620,N_9957);
nand U10811 (N_10811,N_10319,N_10116);
or U10812 (N_10812,N_10387,N_9659);
and U10813 (N_10813,N_10116,N_10238);
xnor U10814 (N_10814,N_9987,N_9896);
and U10815 (N_10815,N_9882,N_10284);
nor U10816 (N_10816,N_10108,N_10129);
or U10817 (N_10817,N_10119,N_9811);
nand U10818 (N_10818,N_9766,N_9653);
nor U10819 (N_10819,N_10374,N_10014);
nor U10820 (N_10820,N_10064,N_10010);
xor U10821 (N_10821,N_10398,N_10360);
nand U10822 (N_10822,N_10130,N_10387);
nand U10823 (N_10823,N_10040,N_10024);
nand U10824 (N_10824,N_10198,N_9678);
and U10825 (N_10825,N_10246,N_10202);
or U10826 (N_10826,N_10382,N_9878);
nor U10827 (N_10827,N_10356,N_9968);
or U10828 (N_10828,N_9789,N_9693);
nand U10829 (N_10829,N_10018,N_9735);
xor U10830 (N_10830,N_9981,N_9678);
xnor U10831 (N_10831,N_9770,N_9818);
nand U10832 (N_10832,N_9824,N_10016);
nor U10833 (N_10833,N_10187,N_9672);
xnor U10834 (N_10834,N_9913,N_9934);
or U10835 (N_10835,N_10274,N_9846);
nor U10836 (N_10836,N_9738,N_9727);
or U10837 (N_10837,N_9904,N_10294);
or U10838 (N_10838,N_10039,N_9884);
or U10839 (N_10839,N_9632,N_10027);
and U10840 (N_10840,N_9997,N_10269);
nor U10841 (N_10841,N_9798,N_9968);
nand U10842 (N_10842,N_10323,N_10203);
xnor U10843 (N_10843,N_10236,N_9857);
and U10844 (N_10844,N_10288,N_10213);
or U10845 (N_10845,N_9655,N_9998);
xor U10846 (N_10846,N_9639,N_9791);
xnor U10847 (N_10847,N_9930,N_9696);
nor U10848 (N_10848,N_10030,N_10094);
nor U10849 (N_10849,N_10176,N_9608);
nand U10850 (N_10850,N_9930,N_9633);
and U10851 (N_10851,N_10354,N_9656);
nor U10852 (N_10852,N_9807,N_10200);
and U10853 (N_10853,N_10125,N_9995);
xor U10854 (N_10854,N_9605,N_10274);
and U10855 (N_10855,N_9934,N_9811);
xnor U10856 (N_10856,N_9843,N_9629);
xnor U10857 (N_10857,N_10088,N_9723);
nand U10858 (N_10858,N_10344,N_9766);
nand U10859 (N_10859,N_10303,N_10207);
xnor U10860 (N_10860,N_9922,N_9802);
and U10861 (N_10861,N_9878,N_10244);
nand U10862 (N_10862,N_10259,N_10227);
xor U10863 (N_10863,N_9608,N_9819);
nand U10864 (N_10864,N_10069,N_10388);
nor U10865 (N_10865,N_9816,N_10216);
nor U10866 (N_10866,N_9791,N_10174);
and U10867 (N_10867,N_9669,N_10212);
and U10868 (N_10868,N_10060,N_10165);
xnor U10869 (N_10869,N_9928,N_10076);
or U10870 (N_10870,N_9958,N_10001);
nor U10871 (N_10871,N_10218,N_9639);
and U10872 (N_10872,N_10338,N_9833);
nor U10873 (N_10873,N_9995,N_10270);
xor U10874 (N_10874,N_10389,N_10173);
nor U10875 (N_10875,N_9838,N_10011);
and U10876 (N_10876,N_9822,N_10238);
xnor U10877 (N_10877,N_9945,N_10238);
xnor U10878 (N_10878,N_9670,N_10118);
nand U10879 (N_10879,N_9850,N_9621);
nor U10880 (N_10880,N_9792,N_10256);
xnor U10881 (N_10881,N_9768,N_10177);
or U10882 (N_10882,N_10167,N_9747);
nand U10883 (N_10883,N_9926,N_10182);
nor U10884 (N_10884,N_9608,N_9897);
or U10885 (N_10885,N_10188,N_9655);
nor U10886 (N_10886,N_9909,N_9831);
and U10887 (N_10887,N_10337,N_10179);
nor U10888 (N_10888,N_9671,N_10124);
xor U10889 (N_10889,N_10072,N_10199);
and U10890 (N_10890,N_9694,N_9685);
nand U10891 (N_10891,N_9836,N_9668);
and U10892 (N_10892,N_9695,N_10335);
nand U10893 (N_10893,N_10310,N_10147);
xnor U10894 (N_10894,N_10361,N_9958);
or U10895 (N_10895,N_9816,N_10388);
or U10896 (N_10896,N_9795,N_10373);
nor U10897 (N_10897,N_10080,N_10318);
and U10898 (N_10898,N_9657,N_9912);
or U10899 (N_10899,N_10006,N_9917);
nor U10900 (N_10900,N_10170,N_9627);
nor U10901 (N_10901,N_10338,N_9930);
xor U10902 (N_10902,N_10003,N_10179);
or U10903 (N_10903,N_9676,N_10005);
and U10904 (N_10904,N_10331,N_9941);
and U10905 (N_10905,N_10015,N_10238);
nor U10906 (N_10906,N_10396,N_10177);
nor U10907 (N_10907,N_10129,N_9962);
xor U10908 (N_10908,N_9659,N_10073);
nor U10909 (N_10909,N_10296,N_10389);
nand U10910 (N_10910,N_10206,N_9699);
and U10911 (N_10911,N_10330,N_10007);
and U10912 (N_10912,N_10275,N_9616);
nand U10913 (N_10913,N_9883,N_10059);
xnor U10914 (N_10914,N_10149,N_10001);
and U10915 (N_10915,N_9652,N_10203);
xnor U10916 (N_10916,N_10194,N_10385);
nand U10917 (N_10917,N_9845,N_10344);
and U10918 (N_10918,N_9964,N_9894);
or U10919 (N_10919,N_9782,N_9941);
xor U10920 (N_10920,N_10056,N_9641);
and U10921 (N_10921,N_9873,N_9683);
or U10922 (N_10922,N_10294,N_9698);
nand U10923 (N_10923,N_10137,N_10014);
nand U10924 (N_10924,N_10271,N_9997);
and U10925 (N_10925,N_9662,N_10255);
and U10926 (N_10926,N_9954,N_10085);
nor U10927 (N_10927,N_9828,N_9632);
or U10928 (N_10928,N_9625,N_9711);
nor U10929 (N_10929,N_10157,N_9700);
and U10930 (N_10930,N_9718,N_10067);
xnor U10931 (N_10931,N_10316,N_9686);
nand U10932 (N_10932,N_10051,N_10206);
or U10933 (N_10933,N_10197,N_9967);
nand U10934 (N_10934,N_10251,N_9752);
nand U10935 (N_10935,N_9620,N_10146);
nor U10936 (N_10936,N_9833,N_9788);
and U10937 (N_10937,N_10336,N_9759);
nand U10938 (N_10938,N_10079,N_10084);
xor U10939 (N_10939,N_10315,N_9930);
and U10940 (N_10940,N_10341,N_9654);
nor U10941 (N_10941,N_9625,N_9602);
and U10942 (N_10942,N_10145,N_10361);
xnor U10943 (N_10943,N_10219,N_9901);
xor U10944 (N_10944,N_10089,N_10170);
xnor U10945 (N_10945,N_9711,N_9688);
xor U10946 (N_10946,N_9784,N_9797);
nand U10947 (N_10947,N_10393,N_10290);
nand U10948 (N_10948,N_9847,N_10297);
xnor U10949 (N_10949,N_10146,N_10359);
nand U10950 (N_10950,N_10327,N_10352);
xor U10951 (N_10951,N_9757,N_10207);
nor U10952 (N_10952,N_10002,N_9701);
xor U10953 (N_10953,N_9807,N_9700);
or U10954 (N_10954,N_10096,N_10072);
nor U10955 (N_10955,N_10008,N_9855);
xnor U10956 (N_10956,N_10235,N_10001);
and U10957 (N_10957,N_9832,N_10099);
and U10958 (N_10958,N_10056,N_9776);
or U10959 (N_10959,N_9939,N_10362);
nor U10960 (N_10960,N_9873,N_10166);
or U10961 (N_10961,N_9638,N_10025);
and U10962 (N_10962,N_9992,N_10015);
xor U10963 (N_10963,N_9900,N_9820);
xor U10964 (N_10964,N_9757,N_10102);
and U10965 (N_10965,N_9979,N_9849);
xor U10966 (N_10966,N_10148,N_10016);
nor U10967 (N_10967,N_10197,N_10196);
nand U10968 (N_10968,N_10244,N_9899);
or U10969 (N_10969,N_10058,N_10055);
nand U10970 (N_10970,N_9632,N_10139);
and U10971 (N_10971,N_9660,N_10195);
xnor U10972 (N_10972,N_9985,N_9657);
nand U10973 (N_10973,N_10342,N_9807);
and U10974 (N_10974,N_9610,N_10329);
and U10975 (N_10975,N_10099,N_10175);
nand U10976 (N_10976,N_9834,N_10005);
nand U10977 (N_10977,N_10236,N_10060);
or U10978 (N_10978,N_9607,N_9992);
and U10979 (N_10979,N_10070,N_9986);
and U10980 (N_10980,N_10015,N_10299);
and U10981 (N_10981,N_10349,N_10171);
nor U10982 (N_10982,N_9697,N_9810);
nor U10983 (N_10983,N_10377,N_9961);
xor U10984 (N_10984,N_10255,N_10345);
and U10985 (N_10985,N_10171,N_10271);
xor U10986 (N_10986,N_9632,N_9627);
or U10987 (N_10987,N_9964,N_9728);
or U10988 (N_10988,N_9832,N_10228);
or U10989 (N_10989,N_9622,N_10053);
or U10990 (N_10990,N_9696,N_9905);
and U10991 (N_10991,N_9879,N_9948);
or U10992 (N_10992,N_10211,N_10174);
xnor U10993 (N_10993,N_9867,N_10130);
xor U10994 (N_10994,N_9621,N_10087);
nor U10995 (N_10995,N_10380,N_10111);
or U10996 (N_10996,N_10011,N_9786);
and U10997 (N_10997,N_9699,N_9673);
xor U10998 (N_10998,N_9949,N_9754);
xnor U10999 (N_10999,N_9601,N_10061);
nand U11000 (N_11000,N_10190,N_9652);
and U11001 (N_11001,N_9940,N_9699);
or U11002 (N_11002,N_10384,N_9611);
xor U11003 (N_11003,N_10270,N_10075);
nor U11004 (N_11004,N_9727,N_10140);
or U11005 (N_11005,N_10107,N_9907);
xor U11006 (N_11006,N_10121,N_10157);
or U11007 (N_11007,N_9801,N_10350);
and U11008 (N_11008,N_10102,N_10015);
nand U11009 (N_11009,N_10017,N_10363);
nor U11010 (N_11010,N_10057,N_10195);
or U11011 (N_11011,N_10279,N_9645);
xor U11012 (N_11012,N_9617,N_9894);
nand U11013 (N_11013,N_10204,N_10106);
nand U11014 (N_11014,N_10377,N_10039);
or U11015 (N_11015,N_10398,N_10246);
nand U11016 (N_11016,N_9976,N_10390);
nor U11017 (N_11017,N_10231,N_9764);
xor U11018 (N_11018,N_10150,N_10153);
or U11019 (N_11019,N_9941,N_9634);
nand U11020 (N_11020,N_9623,N_10374);
xnor U11021 (N_11021,N_10224,N_10359);
or U11022 (N_11022,N_9805,N_9678);
and U11023 (N_11023,N_10142,N_10274);
and U11024 (N_11024,N_10117,N_10299);
nand U11025 (N_11025,N_10132,N_10011);
or U11026 (N_11026,N_10007,N_9924);
or U11027 (N_11027,N_9923,N_9854);
nor U11028 (N_11028,N_10113,N_9880);
or U11029 (N_11029,N_10251,N_9986);
xnor U11030 (N_11030,N_10210,N_9784);
nor U11031 (N_11031,N_9656,N_10121);
nor U11032 (N_11032,N_10160,N_9788);
and U11033 (N_11033,N_9766,N_9971);
nor U11034 (N_11034,N_10109,N_9945);
nand U11035 (N_11035,N_9897,N_9813);
xor U11036 (N_11036,N_10179,N_9705);
and U11037 (N_11037,N_10310,N_10230);
or U11038 (N_11038,N_9644,N_9847);
nand U11039 (N_11039,N_10245,N_9784);
or U11040 (N_11040,N_10223,N_10107);
xor U11041 (N_11041,N_9804,N_9879);
nand U11042 (N_11042,N_9963,N_10264);
nand U11043 (N_11043,N_10008,N_9614);
nand U11044 (N_11044,N_10345,N_9859);
and U11045 (N_11045,N_9882,N_9652);
nor U11046 (N_11046,N_9893,N_9767);
xor U11047 (N_11047,N_9868,N_10387);
and U11048 (N_11048,N_9878,N_9683);
or U11049 (N_11049,N_10120,N_9826);
and U11050 (N_11050,N_9970,N_10237);
nor U11051 (N_11051,N_9646,N_9657);
xor U11052 (N_11052,N_10188,N_9782);
nand U11053 (N_11053,N_10272,N_9797);
xnor U11054 (N_11054,N_9873,N_9628);
nand U11055 (N_11055,N_9933,N_9736);
nand U11056 (N_11056,N_10285,N_9701);
nand U11057 (N_11057,N_10021,N_10379);
and U11058 (N_11058,N_10234,N_10158);
nand U11059 (N_11059,N_10241,N_9810);
nor U11060 (N_11060,N_9910,N_10291);
nand U11061 (N_11061,N_9984,N_9625);
and U11062 (N_11062,N_9694,N_10341);
and U11063 (N_11063,N_9677,N_10077);
xor U11064 (N_11064,N_10262,N_10346);
nor U11065 (N_11065,N_10294,N_10225);
and U11066 (N_11066,N_9795,N_9925);
nand U11067 (N_11067,N_9729,N_9650);
and U11068 (N_11068,N_10368,N_9789);
nor U11069 (N_11069,N_10357,N_10202);
nor U11070 (N_11070,N_10152,N_10008);
and U11071 (N_11071,N_10227,N_10094);
or U11072 (N_11072,N_10395,N_9714);
nor U11073 (N_11073,N_9881,N_9867);
nor U11074 (N_11074,N_10003,N_9906);
nor U11075 (N_11075,N_9756,N_9747);
and U11076 (N_11076,N_10012,N_9799);
and U11077 (N_11077,N_9904,N_9923);
nand U11078 (N_11078,N_10329,N_9622);
or U11079 (N_11079,N_10110,N_9641);
or U11080 (N_11080,N_10077,N_10311);
nand U11081 (N_11081,N_9910,N_9921);
xor U11082 (N_11082,N_9663,N_9909);
and U11083 (N_11083,N_10093,N_10022);
nand U11084 (N_11084,N_10332,N_10040);
or U11085 (N_11085,N_10155,N_9752);
nand U11086 (N_11086,N_10031,N_9982);
nand U11087 (N_11087,N_9814,N_9727);
and U11088 (N_11088,N_10002,N_10308);
or U11089 (N_11089,N_10107,N_9955);
nand U11090 (N_11090,N_10092,N_9707);
nand U11091 (N_11091,N_10294,N_10378);
nand U11092 (N_11092,N_9934,N_10230);
and U11093 (N_11093,N_10367,N_9647);
xor U11094 (N_11094,N_10114,N_10338);
xor U11095 (N_11095,N_9606,N_10359);
nand U11096 (N_11096,N_10184,N_10116);
nand U11097 (N_11097,N_9775,N_10356);
nor U11098 (N_11098,N_10048,N_10168);
nand U11099 (N_11099,N_9793,N_10063);
or U11100 (N_11100,N_9724,N_10028);
or U11101 (N_11101,N_10145,N_10277);
nand U11102 (N_11102,N_9630,N_9696);
xor U11103 (N_11103,N_9682,N_10279);
or U11104 (N_11104,N_10000,N_9607);
or U11105 (N_11105,N_9613,N_9944);
xnor U11106 (N_11106,N_10341,N_9885);
xor U11107 (N_11107,N_10112,N_10328);
xor U11108 (N_11108,N_9710,N_10016);
nor U11109 (N_11109,N_9634,N_9998);
or U11110 (N_11110,N_10357,N_10350);
and U11111 (N_11111,N_10075,N_10295);
nor U11112 (N_11112,N_10093,N_10351);
nand U11113 (N_11113,N_10129,N_10087);
nor U11114 (N_11114,N_10261,N_10389);
nand U11115 (N_11115,N_10309,N_10205);
or U11116 (N_11116,N_10239,N_10071);
xor U11117 (N_11117,N_9875,N_10291);
nand U11118 (N_11118,N_9771,N_9707);
or U11119 (N_11119,N_10146,N_9888);
nand U11120 (N_11120,N_10207,N_9929);
nand U11121 (N_11121,N_10298,N_9967);
nand U11122 (N_11122,N_9966,N_10271);
nand U11123 (N_11123,N_9975,N_9801);
nor U11124 (N_11124,N_10357,N_10294);
nor U11125 (N_11125,N_10347,N_10396);
nor U11126 (N_11126,N_10223,N_10195);
or U11127 (N_11127,N_10014,N_10070);
nand U11128 (N_11128,N_9817,N_9902);
xor U11129 (N_11129,N_9672,N_9972);
nor U11130 (N_11130,N_9921,N_9736);
or U11131 (N_11131,N_9766,N_9716);
and U11132 (N_11132,N_9610,N_9868);
nand U11133 (N_11133,N_9644,N_9907);
or U11134 (N_11134,N_9787,N_10124);
nor U11135 (N_11135,N_9919,N_9618);
and U11136 (N_11136,N_9702,N_9782);
nor U11137 (N_11137,N_9950,N_9649);
or U11138 (N_11138,N_9864,N_9758);
xnor U11139 (N_11139,N_9843,N_10181);
nand U11140 (N_11140,N_9634,N_9901);
or U11141 (N_11141,N_9738,N_9798);
nand U11142 (N_11142,N_10259,N_9983);
nor U11143 (N_11143,N_9947,N_10316);
nor U11144 (N_11144,N_9650,N_9912);
nor U11145 (N_11145,N_10257,N_9892);
and U11146 (N_11146,N_10033,N_10137);
xnor U11147 (N_11147,N_9841,N_10235);
nand U11148 (N_11148,N_10241,N_10059);
xnor U11149 (N_11149,N_9764,N_10274);
and U11150 (N_11150,N_10388,N_9936);
nand U11151 (N_11151,N_9716,N_9823);
and U11152 (N_11152,N_10065,N_9999);
xnor U11153 (N_11153,N_9801,N_9811);
nand U11154 (N_11154,N_10219,N_9934);
nand U11155 (N_11155,N_9909,N_9933);
xnor U11156 (N_11156,N_10066,N_9712);
nor U11157 (N_11157,N_9648,N_9849);
and U11158 (N_11158,N_9762,N_9970);
nor U11159 (N_11159,N_9946,N_9987);
nor U11160 (N_11160,N_9931,N_9947);
xor U11161 (N_11161,N_9744,N_9644);
and U11162 (N_11162,N_9720,N_9905);
nor U11163 (N_11163,N_10161,N_10207);
xor U11164 (N_11164,N_10202,N_10324);
and U11165 (N_11165,N_9883,N_9743);
nor U11166 (N_11166,N_10129,N_10205);
xor U11167 (N_11167,N_10197,N_9621);
xnor U11168 (N_11168,N_9625,N_10124);
and U11169 (N_11169,N_9907,N_9624);
and U11170 (N_11170,N_10180,N_9684);
nand U11171 (N_11171,N_9723,N_10073);
or U11172 (N_11172,N_9754,N_9911);
xor U11173 (N_11173,N_10148,N_10076);
xnor U11174 (N_11174,N_9987,N_10105);
nand U11175 (N_11175,N_9758,N_10014);
nor U11176 (N_11176,N_9893,N_9806);
xor U11177 (N_11177,N_9848,N_10125);
nand U11178 (N_11178,N_10286,N_9841);
or U11179 (N_11179,N_10213,N_10140);
nor U11180 (N_11180,N_9931,N_10262);
or U11181 (N_11181,N_10020,N_9842);
nand U11182 (N_11182,N_10293,N_9668);
nand U11183 (N_11183,N_9883,N_10356);
and U11184 (N_11184,N_9863,N_9867);
nand U11185 (N_11185,N_10238,N_9738);
and U11186 (N_11186,N_10357,N_10345);
and U11187 (N_11187,N_9639,N_9737);
nor U11188 (N_11188,N_10326,N_10298);
or U11189 (N_11189,N_10348,N_9880);
and U11190 (N_11190,N_9614,N_10273);
or U11191 (N_11191,N_10129,N_9663);
or U11192 (N_11192,N_10066,N_9952);
and U11193 (N_11193,N_10033,N_10252);
nand U11194 (N_11194,N_9704,N_10298);
xnor U11195 (N_11195,N_10319,N_9972);
nand U11196 (N_11196,N_9834,N_10322);
and U11197 (N_11197,N_9634,N_10026);
nor U11198 (N_11198,N_10002,N_9983);
nor U11199 (N_11199,N_9789,N_9624);
nand U11200 (N_11200,N_10684,N_10419);
and U11201 (N_11201,N_11167,N_10928);
nor U11202 (N_11202,N_11130,N_10648);
nand U11203 (N_11203,N_10481,N_10647);
nand U11204 (N_11204,N_10955,N_10806);
and U11205 (N_11205,N_10580,N_10552);
xor U11206 (N_11206,N_10704,N_10697);
nand U11207 (N_11207,N_11067,N_11190);
nor U11208 (N_11208,N_10968,N_11191);
xnor U11209 (N_11209,N_10510,N_10960);
nor U11210 (N_11210,N_10724,N_11162);
and U11211 (N_11211,N_11106,N_11182);
nor U11212 (N_11212,N_11132,N_11107);
or U11213 (N_11213,N_10599,N_10987);
or U11214 (N_11214,N_10855,N_10637);
xor U11215 (N_11215,N_11144,N_10834);
and U11216 (N_11216,N_10755,N_10541);
nor U11217 (N_11217,N_10471,N_10813);
or U11218 (N_11218,N_11126,N_11154);
and U11219 (N_11219,N_10948,N_11021);
or U11220 (N_11220,N_11145,N_10621);
xor U11221 (N_11221,N_10750,N_10915);
nor U11222 (N_11222,N_10420,N_10656);
and U11223 (N_11223,N_10433,N_10469);
or U11224 (N_11224,N_11159,N_11036);
and U11225 (N_11225,N_10448,N_11189);
or U11226 (N_11226,N_11072,N_10989);
or U11227 (N_11227,N_10429,N_10897);
and U11228 (N_11228,N_11031,N_10836);
nand U11229 (N_11229,N_11051,N_10726);
or U11230 (N_11230,N_10464,N_10734);
nor U11231 (N_11231,N_10486,N_10454);
and U11232 (N_11232,N_10493,N_10479);
nor U11233 (N_11233,N_10563,N_10706);
or U11234 (N_11234,N_10498,N_11065);
or U11235 (N_11235,N_10767,N_10931);
or U11236 (N_11236,N_11063,N_10571);
nor U11237 (N_11237,N_10625,N_11155);
and U11238 (N_11238,N_10600,N_10550);
xnor U11239 (N_11239,N_10747,N_10876);
nor U11240 (N_11240,N_10634,N_10413);
nand U11241 (N_11241,N_10640,N_10785);
nor U11242 (N_11242,N_10430,N_11094);
or U11243 (N_11243,N_10722,N_10774);
or U11244 (N_11244,N_10545,N_11011);
or U11245 (N_11245,N_10994,N_11052);
and U11246 (N_11246,N_10439,N_10477);
or U11247 (N_11247,N_10743,N_10515);
xor U11248 (N_11248,N_10654,N_10460);
and U11249 (N_11249,N_10615,N_11168);
xnor U11250 (N_11250,N_10740,N_10679);
nand U11251 (N_11251,N_10718,N_10804);
or U11252 (N_11252,N_10936,N_11108);
or U11253 (N_11253,N_11117,N_10961);
xnor U11254 (N_11254,N_10958,N_10831);
nor U11255 (N_11255,N_10665,N_10551);
nand U11256 (N_11256,N_10472,N_11058);
xnor U11257 (N_11257,N_11102,N_11074);
xor U11258 (N_11258,N_10675,N_10524);
and U11259 (N_11259,N_11071,N_10427);
or U11260 (N_11260,N_11133,N_10459);
nor U11261 (N_11261,N_10555,N_11068);
or U11262 (N_11262,N_10607,N_10887);
and U11263 (N_11263,N_10560,N_10632);
nor U11264 (N_11264,N_11002,N_10520);
or U11265 (N_11265,N_10548,N_10466);
xnor U11266 (N_11266,N_10888,N_10771);
xnor U11267 (N_11267,N_10696,N_11013);
nand U11268 (N_11268,N_11142,N_10966);
or U11269 (N_11269,N_10764,N_10638);
and U11270 (N_11270,N_10890,N_10962);
and U11271 (N_11271,N_11089,N_11043);
nor U11272 (N_11272,N_11038,N_10456);
nand U11273 (N_11273,N_10916,N_11044);
nand U11274 (N_11274,N_10801,N_11005);
xnor U11275 (N_11275,N_10883,N_11033);
and U11276 (N_11276,N_10485,N_11087);
and U11277 (N_11277,N_10416,N_10816);
or U11278 (N_11278,N_10932,N_10609);
xnor U11279 (N_11279,N_10593,N_10532);
nand U11280 (N_11280,N_11134,N_11016);
nor U11281 (N_11281,N_10759,N_10963);
and U11282 (N_11282,N_11128,N_10846);
nand U11283 (N_11283,N_10789,N_10438);
nor U11284 (N_11284,N_10701,N_10408);
or U11285 (N_11285,N_10797,N_10851);
nand U11286 (N_11286,N_10453,N_10494);
nand U11287 (N_11287,N_10959,N_10886);
or U11288 (N_11288,N_10569,N_11118);
or U11289 (N_11289,N_11194,N_10680);
and U11290 (N_11290,N_10972,N_11040);
and U11291 (N_11291,N_10500,N_10901);
and U11292 (N_11292,N_10484,N_11125);
and U11293 (N_11293,N_11129,N_10773);
nor U11294 (N_11294,N_10799,N_10745);
nor U11295 (N_11295,N_10980,N_11039);
nor U11296 (N_11296,N_10604,N_11122);
nor U11297 (N_11297,N_10997,N_10974);
xor U11298 (N_11298,N_10798,N_10415);
or U11299 (N_11299,N_10713,N_10975);
nand U11300 (N_11300,N_10753,N_10933);
or U11301 (N_11301,N_10424,N_10480);
or U11302 (N_11302,N_10768,N_11095);
xor U11303 (N_11303,N_10410,N_11019);
and U11304 (N_11304,N_10613,N_10492);
and U11305 (N_11305,N_10570,N_11111);
and U11306 (N_11306,N_10461,N_10957);
xor U11307 (N_11307,N_10885,N_10881);
xor U11308 (N_11308,N_11081,N_11056);
xnor U11309 (N_11309,N_10482,N_10409);
or U11310 (N_11310,N_10708,N_10852);
or U11311 (N_11311,N_10940,N_10659);
nor U11312 (N_11312,N_10516,N_10926);
nand U11313 (N_11313,N_10751,N_10733);
xor U11314 (N_11314,N_10508,N_10739);
or U11315 (N_11315,N_10451,N_11086);
xor U11316 (N_11316,N_10819,N_10951);
or U11317 (N_11317,N_10611,N_10872);
or U11318 (N_11318,N_11008,N_10712);
and U11319 (N_11319,N_10450,N_10690);
nor U11320 (N_11320,N_10711,N_11001);
xor U11321 (N_11321,N_10910,N_10919);
or U11322 (N_11322,N_10929,N_11096);
and U11323 (N_11323,N_11042,N_10761);
nor U11324 (N_11324,N_10578,N_10629);
or U11325 (N_11325,N_10984,N_10673);
xnor U11326 (N_11326,N_10826,N_10810);
or U11327 (N_11327,N_10729,N_11059);
and U11328 (N_11328,N_11152,N_10996);
xnor U11329 (N_11329,N_11034,N_10805);
or U11330 (N_11330,N_11027,N_10502);
and U11331 (N_11331,N_11198,N_10720);
nor U11332 (N_11332,N_10730,N_10436);
xnor U11333 (N_11333,N_11103,N_11143);
nand U11334 (N_11334,N_10802,N_10535);
nor U11335 (N_11335,N_10573,N_10820);
xnor U11336 (N_11336,N_11025,N_11113);
xnor U11337 (N_11337,N_11199,N_10657);
and U11338 (N_11338,N_10976,N_10788);
nor U11339 (N_11339,N_10681,N_10754);
xor U11340 (N_11340,N_10889,N_10749);
xnor U11341 (N_11341,N_11188,N_10698);
xnor U11342 (N_11342,N_10833,N_10642);
or U11343 (N_11343,N_10655,N_11187);
xnor U11344 (N_11344,N_10589,N_10918);
nor U11345 (N_11345,N_10445,N_10737);
xor U11346 (N_11346,N_10930,N_10981);
xor U11347 (N_11347,N_10663,N_11119);
nor U11348 (N_11348,N_11093,N_11060);
or U11349 (N_11349,N_11186,N_10863);
nor U11350 (N_11350,N_10891,N_10978);
and U11351 (N_11351,N_11146,N_10631);
nand U11352 (N_11352,N_10623,N_10902);
nor U11353 (N_11353,N_11176,N_10909);
or U11354 (N_11354,N_10939,N_10495);
nand U11355 (N_11355,N_10988,N_10867);
or U11356 (N_11356,N_11100,N_10544);
or U11357 (N_11357,N_10871,N_10425);
xor U11358 (N_11358,N_11064,N_11179);
and U11359 (N_11359,N_10870,N_10517);
and U11360 (N_11360,N_10934,N_10501);
or U11361 (N_11361,N_10567,N_10736);
or U11362 (N_11362,N_10503,N_10403);
nand U11363 (N_11363,N_11026,N_10945);
nor U11364 (N_11364,N_11050,N_11147);
xor U11365 (N_11365,N_10908,N_10763);
or U11366 (N_11366,N_11069,N_10840);
xor U11367 (N_11367,N_11170,N_10766);
nand U11368 (N_11368,N_10509,N_10991);
and U11369 (N_11369,N_11032,N_11097);
xor U11370 (N_11370,N_10896,N_10964);
nor U11371 (N_11371,N_10525,N_10884);
nand U11372 (N_11372,N_11127,N_10463);
or U11373 (N_11373,N_10792,N_10686);
nor U11374 (N_11374,N_10434,N_10823);
or U11375 (N_11375,N_10861,N_10473);
xnor U11376 (N_11376,N_10598,N_11045);
xnor U11377 (N_11377,N_10458,N_11017);
and U11378 (N_11378,N_10842,N_11020);
or U11379 (N_11379,N_10973,N_11078);
or U11380 (N_11380,N_10576,N_10967);
and U11381 (N_11381,N_10591,N_10772);
and U11382 (N_11382,N_10719,N_10594);
nor U11383 (N_11383,N_10407,N_11061);
nor U11384 (N_11384,N_10941,N_10705);
nand U11385 (N_11385,N_10995,N_10983);
nand U11386 (N_11386,N_10618,N_10911);
nor U11387 (N_11387,N_11151,N_10619);
xnor U11388 (N_11388,N_11101,N_10979);
nand U11389 (N_11389,N_10418,N_10531);
and U11390 (N_11390,N_10732,N_10894);
and U11391 (N_11391,N_10470,N_10682);
or U11392 (N_11392,N_10946,N_11003);
nor U11393 (N_11393,N_10622,N_11156);
nand U11394 (N_11394,N_10757,N_10595);
nor U11395 (N_11395,N_10566,N_10899);
xor U11396 (N_11396,N_10444,N_10582);
or U11397 (N_11397,N_10794,N_10814);
and U11398 (N_11398,N_10558,N_10937);
and U11399 (N_11399,N_10923,N_10850);
nand U11400 (N_11400,N_10790,N_10547);
nand U11401 (N_11401,N_11135,N_10649);
and U11402 (N_11402,N_10447,N_10822);
or U11403 (N_11403,N_11163,N_10664);
nor U11404 (N_11404,N_10653,N_11158);
xor U11405 (N_11405,N_10956,N_10568);
or U11406 (N_11406,N_10553,N_10412);
nor U11407 (N_11407,N_10462,N_10858);
xnor U11408 (N_11408,N_10400,N_10489);
and U11409 (N_11409,N_10422,N_11076);
nand U11410 (N_11410,N_10542,N_10862);
xor U11411 (N_11411,N_10791,N_10449);
nor U11412 (N_11412,N_10401,N_10818);
nand U11413 (N_11413,N_11009,N_10954);
nand U11414 (N_11414,N_10683,N_11048);
nor U11415 (N_11415,N_10709,N_10920);
and U11416 (N_11416,N_10935,N_10917);
xnor U11417 (N_11417,N_10702,N_10921);
and U11418 (N_11418,N_10841,N_10514);
and U11419 (N_11419,N_10830,N_10778);
or U11420 (N_11420,N_10710,N_10832);
nor U11421 (N_11421,N_11195,N_11148);
nor U11422 (N_11422,N_10942,N_10859);
nand U11423 (N_11423,N_10856,N_10970);
xor U11424 (N_11424,N_10716,N_10695);
and U11425 (N_11425,N_10783,N_10635);
nor U11426 (N_11426,N_10837,N_10985);
nor U11427 (N_11427,N_10630,N_10483);
nand U11428 (N_11428,N_10676,N_10953);
xor U11429 (N_11429,N_10824,N_10441);
or U11430 (N_11430,N_10487,N_10584);
xnor U11431 (N_11431,N_10913,N_11183);
xnor U11432 (N_11432,N_10411,N_11160);
nand U11433 (N_11433,N_10848,N_10868);
or U11434 (N_11434,N_10691,N_10857);
nor U11435 (N_11435,N_10646,N_11084);
nand U11436 (N_11436,N_10924,N_10949);
xor U11437 (N_11437,N_11006,N_10452);
nand U11438 (N_11438,N_10624,N_10900);
nand U11439 (N_11439,N_10717,N_10432);
xnor U11440 (N_11440,N_10556,N_10603);
nor U11441 (N_11441,N_10543,N_10998);
xnor U11442 (N_11442,N_11085,N_11090);
and U11443 (N_11443,N_10561,N_10905);
xor U11444 (N_11444,N_11079,N_10644);
xnor U11445 (N_11445,N_10597,N_10670);
nand U11446 (N_11446,N_10874,N_10575);
or U11447 (N_11447,N_10440,N_11029);
nor U11448 (N_11448,N_10721,N_11178);
nand U11449 (N_11449,N_10678,N_11070);
and U11450 (N_11450,N_10574,N_10835);
nor U11451 (N_11451,N_10950,N_10406);
nand U11452 (N_11452,N_10617,N_11083);
and U11453 (N_11453,N_10402,N_10756);
or U11454 (N_11454,N_10808,N_10744);
nand U11455 (N_11455,N_10610,N_10728);
xor U11456 (N_11456,N_10476,N_10825);
and U11457 (N_11457,N_10478,N_11012);
or U11458 (N_11458,N_11024,N_10999);
or U11459 (N_11459,N_10758,N_11121);
and U11460 (N_11460,N_11014,N_11098);
xnor U11461 (N_11461,N_11192,N_10669);
nand U11462 (N_11462,N_10925,N_11104);
and U11463 (N_11463,N_10893,N_10530);
nor U11464 (N_11464,N_10853,N_10829);
and U11465 (N_11465,N_10431,N_10986);
or U11466 (N_11466,N_10496,N_10943);
nor U11467 (N_11467,N_10777,N_11066);
or U11468 (N_11468,N_10780,N_10849);
xor U11469 (N_11469,N_11047,N_11171);
and U11470 (N_11470,N_11092,N_10760);
or U11471 (N_11471,N_10457,N_10735);
xnor U11472 (N_11472,N_11175,N_11172);
nand U11473 (N_11473,N_10914,N_10793);
nand U11474 (N_11474,N_10800,N_10786);
xor U11475 (N_11475,N_10612,N_11080);
xor U11476 (N_11476,N_10677,N_10748);
or U11477 (N_11477,N_11049,N_10443);
xor U11478 (N_11478,N_11166,N_10421);
xnor U11479 (N_11479,N_10405,N_10992);
or U11480 (N_11480,N_10442,N_10650);
and U11481 (N_11481,N_10882,N_10414);
xor U11482 (N_11482,N_10581,N_10775);
or U11483 (N_11483,N_11053,N_10592);
and U11484 (N_11484,N_11161,N_11054);
nor U11485 (N_11485,N_10742,N_10528);
nor U11486 (N_11486,N_10435,N_10714);
nand U11487 (N_11487,N_11141,N_10626);
nand U11488 (N_11488,N_10437,N_10865);
nor U11489 (N_11489,N_10828,N_11112);
or U11490 (N_11490,N_10877,N_10572);
or U11491 (N_11491,N_10674,N_11075);
or U11492 (N_11492,N_10505,N_10554);
nand U11493 (N_11493,N_10854,N_10769);
nor U11494 (N_11494,N_10661,N_10455);
xor U11495 (N_11495,N_10579,N_10534);
nand U11496 (N_11496,N_10601,N_10596);
xnor U11497 (N_11497,N_10662,N_10467);
xnor U11498 (N_11498,N_11137,N_10549);
nor U11499 (N_11499,N_10869,N_10927);
or U11500 (N_11500,N_10536,N_11149);
xnor U11501 (N_11501,N_10614,N_10860);
nand U11502 (N_11502,N_10965,N_10523);
or U11503 (N_11503,N_10468,N_10526);
and U11504 (N_11504,N_10504,N_10969);
nor U11505 (N_11505,N_10685,N_10539);
or U11506 (N_11506,N_10583,N_10971);
xor U11507 (N_11507,N_10562,N_11140);
nor U11508 (N_11508,N_10587,N_11124);
nor U11509 (N_11509,N_10880,N_10529);
xnor U11510 (N_11510,N_10488,N_11105);
or U11511 (N_11511,N_10694,N_10633);
nand U11512 (N_11512,N_11055,N_11174);
nor U11513 (N_11513,N_10658,N_11109);
nor U11514 (N_11514,N_10559,N_11169);
xor U11515 (N_11515,N_10538,N_10491);
nor U11516 (N_11516,N_11150,N_10922);
and U11517 (N_11517,N_11115,N_10636);
nand U11518 (N_11518,N_10795,N_10616);
nor U11519 (N_11519,N_10511,N_11091);
xor U11520 (N_11520,N_10417,N_10779);
and U11521 (N_11521,N_10847,N_10907);
nand U11522 (N_11522,N_10947,N_10423);
nor U11523 (N_11523,N_10428,N_10518);
xnor U11524 (N_11524,N_10727,N_10404);
nand U11525 (N_11525,N_10590,N_11088);
xor U11526 (N_11526,N_10903,N_10776);
xnor U11527 (N_11527,N_10904,N_10537);
nor U11528 (N_11528,N_10811,N_10898);
and U11529 (N_11529,N_10787,N_11181);
nor U11530 (N_11530,N_10873,N_11018);
and U11531 (N_11531,N_11153,N_11010);
nand U11532 (N_11532,N_10689,N_11138);
and U11533 (N_11533,N_11082,N_10577);
xor U11534 (N_11534,N_10944,N_11157);
or U11535 (N_11535,N_10723,N_11099);
and U11536 (N_11536,N_10620,N_10827);
or U11537 (N_11537,N_10875,N_11062);
and U11538 (N_11538,N_10707,N_10641);
xor U11539 (N_11539,N_10781,N_10977);
or U11540 (N_11540,N_10512,N_11193);
nor U11541 (N_11541,N_10513,N_10725);
and U11542 (N_11542,N_10660,N_10879);
nor U11543 (N_11543,N_11177,N_10938);
xor U11544 (N_11544,N_11184,N_10527);
nor U11545 (N_11545,N_10605,N_10807);
xnor U11546 (N_11546,N_10606,N_10645);
nor U11547 (N_11547,N_10703,N_11022);
xor U11548 (N_11548,N_10843,N_10892);
xor U11549 (N_11549,N_10809,N_10839);
nor U11550 (N_11550,N_10475,N_11023);
nand U11551 (N_11551,N_11173,N_10557);
or U11552 (N_11552,N_10608,N_10465);
and U11553 (N_11553,N_10497,N_11123);
nor U11554 (N_11554,N_10864,N_10895);
xor U11555 (N_11555,N_10752,N_11165);
xor U11556 (N_11556,N_10533,N_11116);
nor U11557 (N_11557,N_10715,N_10446);
and U11558 (N_11558,N_10693,N_11114);
and U11559 (N_11559,N_11004,N_11136);
xor U11560 (N_11560,N_10521,N_11120);
nor U11561 (N_11561,N_10815,N_11007);
xnor U11562 (N_11562,N_10817,N_11041);
xor U11563 (N_11563,N_10845,N_10506);
xnor U11564 (N_11564,N_10652,N_11073);
nand U11565 (N_11565,N_10699,N_10565);
xnor U11566 (N_11566,N_10627,N_10784);
xnor U11567 (N_11567,N_10731,N_10564);
nor U11568 (N_11568,N_10668,N_10585);
or U11569 (N_11569,N_10540,N_10499);
xor U11570 (N_11570,N_10762,N_10796);
and U11571 (N_11571,N_11030,N_10866);
or U11572 (N_11572,N_11131,N_10651);
xor U11573 (N_11573,N_11185,N_11110);
or U11574 (N_11574,N_10993,N_10906);
xor U11575 (N_11575,N_10782,N_10667);
nand U11576 (N_11576,N_10426,N_10803);
nand U11577 (N_11577,N_11000,N_10687);
or U11578 (N_11578,N_11057,N_10844);
nor U11579 (N_11579,N_10639,N_10474);
and U11580 (N_11580,N_10522,N_11077);
nand U11581 (N_11581,N_11015,N_10519);
nor U11582 (N_11582,N_11028,N_10490);
nor U11583 (N_11583,N_10738,N_11046);
xor U11584 (N_11584,N_10990,N_10507);
xor U11585 (N_11585,N_11196,N_10643);
and U11586 (N_11586,N_11164,N_10666);
nand U11587 (N_11587,N_10692,N_11037);
xor U11588 (N_11588,N_10628,N_10700);
xnor U11589 (N_11589,N_10688,N_10838);
nor U11590 (N_11590,N_10821,N_11180);
or U11591 (N_11591,N_11197,N_10671);
and U11592 (N_11592,N_10741,N_10588);
and U11593 (N_11593,N_10546,N_10770);
nor U11594 (N_11594,N_10982,N_11139);
nand U11595 (N_11595,N_10746,N_10765);
or U11596 (N_11596,N_10602,N_10586);
or U11597 (N_11597,N_10672,N_10812);
xor U11598 (N_11598,N_10952,N_10912);
nand U11599 (N_11599,N_10878,N_11035);
nor U11600 (N_11600,N_10458,N_10888);
nand U11601 (N_11601,N_10467,N_11138);
nand U11602 (N_11602,N_11099,N_10626);
nand U11603 (N_11603,N_10567,N_11198);
or U11604 (N_11604,N_11142,N_11077);
or U11605 (N_11605,N_10990,N_10873);
or U11606 (N_11606,N_10649,N_11102);
and U11607 (N_11607,N_11025,N_11075);
or U11608 (N_11608,N_10477,N_11065);
or U11609 (N_11609,N_11081,N_11197);
and U11610 (N_11610,N_10772,N_10984);
or U11611 (N_11611,N_10856,N_11063);
xor U11612 (N_11612,N_11136,N_10713);
nor U11613 (N_11613,N_11012,N_11135);
nand U11614 (N_11614,N_11116,N_10804);
or U11615 (N_11615,N_11021,N_10792);
xor U11616 (N_11616,N_10841,N_10709);
and U11617 (N_11617,N_10835,N_10947);
and U11618 (N_11618,N_10963,N_10443);
and U11619 (N_11619,N_10946,N_10403);
nand U11620 (N_11620,N_10695,N_10517);
xor U11621 (N_11621,N_10677,N_10993);
or U11622 (N_11622,N_10945,N_11033);
nand U11623 (N_11623,N_10975,N_10588);
nor U11624 (N_11624,N_10892,N_10709);
xor U11625 (N_11625,N_10972,N_10533);
or U11626 (N_11626,N_10857,N_10841);
nor U11627 (N_11627,N_10734,N_10638);
or U11628 (N_11628,N_10646,N_11023);
or U11629 (N_11629,N_10851,N_10891);
or U11630 (N_11630,N_10970,N_10783);
or U11631 (N_11631,N_10995,N_10965);
nor U11632 (N_11632,N_10901,N_11184);
or U11633 (N_11633,N_10451,N_11023);
nand U11634 (N_11634,N_11154,N_10516);
or U11635 (N_11635,N_10862,N_10691);
xor U11636 (N_11636,N_10818,N_11181);
xnor U11637 (N_11637,N_11098,N_10838);
or U11638 (N_11638,N_10621,N_11096);
and U11639 (N_11639,N_11054,N_10574);
nand U11640 (N_11640,N_10918,N_11106);
and U11641 (N_11641,N_10883,N_10866);
nand U11642 (N_11642,N_10642,N_10651);
nor U11643 (N_11643,N_10939,N_11108);
nor U11644 (N_11644,N_11181,N_10623);
nor U11645 (N_11645,N_11128,N_10952);
xor U11646 (N_11646,N_11045,N_10768);
or U11647 (N_11647,N_10895,N_11182);
and U11648 (N_11648,N_11060,N_10586);
xnor U11649 (N_11649,N_11068,N_10568);
nor U11650 (N_11650,N_10786,N_10612);
xnor U11651 (N_11651,N_10715,N_10613);
nand U11652 (N_11652,N_11151,N_10713);
or U11653 (N_11653,N_10547,N_11061);
nor U11654 (N_11654,N_10881,N_10763);
nor U11655 (N_11655,N_10912,N_10485);
nand U11656 (N_11656,N_11054,N_11107);
or U11657 (N_11657,N_11188,N_10458);
or U11658 (N_11658,N_11011,N_10782);
nand U11659 (N_11659,N_10786,N_10734);
nor U11660 (N_11660,N_11049,N_10576);
nand U11661 (N_11661,N_10454,N_10855);
nand U11662 (N_11662,N_11156,N_11147);
or U11663 (N_11663,N_10605,N_10899);
nor U11664 (N_11664,N_10785,N_10496);
nor U11665 (N_11665,N_11175,N_10685);
or U11666 (N_11666,N_11031,N_10729);
and U11667 (N_11667,N_10944,N_11087);
nor U11668 (N_11668,N_10433,N_10946);
or U11669 (N_11669,N_10746,N_10414);
nor U11670 (N_11670,N_10709,N_10793);
xor U11671 (N_11671,N_10660,N_11006);
xor U11672 (N_11672,N_10988,N_10623);
xor U11673 (N_11673,N_10839,N_10748);
nand U11674 (N_11674,N_11163,N_10618);
xor U11675 (N_11675,N_10715,N_10454);
and U11676 (N_11676,N_10554,N_10644);
nor U11677 (N_11677,N_11103,N_11108);
and U11678 (N_11678,N_11128,N_10686);
nor U11679 (N_11679,N_11189,N_10458);
nand U11680 (N_11680,N_11029,N_10905);
xnor U11681 (N_11681,N_11093,N_11125);
nor U11682 (N_11682,N_11040,N_11057);
nor U11683 (N_11683,N_11128,N_11108);
and U11684 (N_11684,N_10449,N_10994);
or U11685 (N_11685,N_10699,N_10412);
nand U11686 (N_11686,N_10723,N_10767);
nand U11687 (N_11687,N_10804,N_10514);
nor U11688 (N_11688,N_10418,N_10899);
xor U11689 (N_11689,N_10738,N_10525);
nor U11690 (N_11690,N_11061,N_10769);
nor U11691 (N_11691,N_10727,N_10801);
xor U11692 (N_11692,N_10667,N_10924);
or U11693 (N_11693,N_11064,N_11115);
nor U11694 (N_11694,N_10479,N_11133);
and U11695 (N_11695,N_11115,N_11118);
nand U11696 (N_11696,N_11156,N_11036);
nand U11697 (N_11697,N_10710,N_10484);
or U11698 (N_11698,N_10730,N_10873);
xnor U11699 (N_11699,N_10564,N_11107);
or U11700 (N_11700,N_10815,N_11070);
and U11701 (N_11701,N_11134,N_10483);
or U11702 (N_11702,N_10853,N_10801);
nand U11703 (N_11703,N_10577,N_10925);
nand U11704 (N_11704,N_11167,N_10497);
nor U11705 (N_11705,N_10698,N_10764);
or U11706 (N_11706,N_10999,N_10928);
xor U11707 (N_11707,N_10968,N_10926);
nand U11708 (N_11708,N_11148,N_10621);
nand U11709 (N_11709,N_11123,N_10499);
nand U11710 (N_11710,N_11070,N_10723);
nand U11711 (N_11711,N_10457,N_10711);
xor U11712 (N_11712,N_10631,N_10415);
and U11713 (N_11713,N_10675,N_10593);
xor U11714 (N_11714,N_10705,N_11036);
or U11715 (N_11715,N_10673,N_10486);
nor U11716 (N_11716,N_10853,N_10615);
nand U11717 (N_11717,N_11198,N_10672);
xor U11718 (N_11718,N_10557,N_10674);
nor U11719 (N_11719,N_10817,N_10733);
xor U11720 (N_11720,N_11120,N_10546);
or U11721 (N_11721,N_10436,N_10420);
or U11722 (N_11722,N_10508,N_10459);
and U11723 (N_11723,N_10956,N_10450);
or U11724 (N_11724,N_10928,N_10866);
nand U11725 (N_11725,N_11016,N_10728);
nand U11726 (N_11726,N_11064,N_10622);
nor U11727 (N_11727,N_10923,N_10481);
xor U11728 (N_11728,N_10702,N_11082);
and U11729 (N_11729,N_10551,N_10679);
nand U11730 (N_11730,N_10758,N_10507);
xor U11731 (N_11731,N_10960,N_10442);
nor U11732 (N_11732,N_10856,N_10671);
nand U11733 (N_11733,N_10548,N_10912);
and U11734 (N_11734,N_10403,N_10887);
xnor U11735 (N_11735,N_10909,N_11021);
xor U11736 (N_11736,N_10684,N_10977);
xor U11737 (N_11737,N_10421,N_10903);
nor U11738 (N_11738,N_10914,N_10469);
xor U11739 (N_11739,N_11056,N_10839);
nand U11740 (N_11740,N_11045,N_10584);
nor U11741 (N_11741,N_11164,N_10670);
and U11742 (N_11742,N_10921,N_10644);
xor U11743 (N_11743,N_11101,N_11028);
nor U11744 (N_11744,N_10417,N_10408);
nor U11745 (N_11745,N_10966,N_10711);
xor U11746 (N_11746,N_10534,N_10442);
nand U11747 (N_11747,N_10440,N_10509);
xnor U11748 (N_11748,N_11129,N_10539);
and U11749 (N_11749,N_10732,N_11108);
and U11750 (N_11750,N_11118,N_10582);
nand U11751 (N_11751,N_10607,N_11097);
and U11752 (N_11752,N_10820,N_11146);
nor U11753 (N_11753,N_10847,N_11159);
and U11754 (N_11754,N_10919,N_10543);
or U11755 (N_11755,N_10866,N_10872);
or U11756 (N_11756,N_10767,N_10614);
and U11757 (N_11757,N_10683,N_10425);
or U11758 (N_11758,N_10607,N_10826);
nand U11759 (N_11759,N_10428,N_11182);
xnor U11760 (N_11760,N_10854,N_10439);
or U11761 (N_11761,N_10921,N_11047);
xnor U11762 (N_11762,N_10512,N_10766);
nor U11763 (N_11763,N_11190,N_11056);
xnor U11764 (N_11764,N_10658,N_10686);
or U11765 (N_11765,N_11073,N_10625);
nor U11766 (N_11766,N_10840,N_10589);
nor U11767 (N_11767,N_10943,N_10777);
xnor U11768 (N_11768,N_11139,N_11081);
nand U11769 (N_11769,N_10560,N_10919);
or U11770 (N_11770,N_10665,N_10658);
xnor U11771 (N_11771,N_10553,N_11163);
nand U11772 (N_11772,N_10519,N_10928);
nand U11773 (N_11773,N_10944,N_10635);
and U11774 (N_11774,N_10520,N_10576);
and U11775 (N_11775,N_10770,N_10812);
nand U11776 (N_11776,N_10943,N_10824);
xnor U11777 (N_11777,N_10899,N_10905);
or U11778 (N_11778,N_10451,N_10756);
and U11779 (N_11779,N_10564,N_11101);
and U11780 (N_11780,N_10508,N_10805);
nor U11781 (N_11781,N_10646,N_10905);
or U11782 (N_11782,N_10476,N_11197);
nand U11783 (N_11783,N_10977,N_10839);
xnor U11784 (N_11784,N_10954,N_10612);
nor U11785 (N_11785,N_11115,N_10683);
nand U11786 (N_11786,N_10640,N_10888);
and U11787 (N_11787,N_10925,N_10628);
and U11788 (N_11788,N_10701,N_10455);
nor U11789 (N_11789,N_11056,N_10557);
nand U11790 (N_11790,N_10714,N_11094);
or U11791 (N_11791,N_10789,N_10753);
nor U11792 (N_11792,N_11025,N_10402);
nand U11793 (N_11793,N_11115,N_10424);
nand U11794 (N_11794,N_10894,N_11120);
nor U11795 (N_11795,N_10968,N_11179);
and U11796 (N_11796,N_10790,N_11117);
nand U11797 (N_11797,N_11118,N_10896);
nand U11798 (N_11798,N_11099,N_10503);
nor U11799 (N_11799,N_11123,N_11054);
nor U11800 (N_11800,N_10988,N_10671);
xnor U11801 (N_11801,N_10690,N_10838);
and U11802 (N_11802,N_11098,N_10496);
xor U11803 (N_11803,N_10817,N_10730);
or U11804 (N_11804,N_10950,N_10865);
xnor U11805 (N_11805,N_10994,N_10965);
nor U11806 (N_11806,N_10619,N_11107);
xor U11807 (N_11807,N_11145,N_11147);
and U11808 (N_11808,N_11169,N_10763);
and U11809 (N_11809,N_11162,N_10863);
or U11810 (N_11810,N_11162,N_10459);
nand U11811 (N_11811,N_10494,N_10731);
or U11812 (N_11812,N_10869,N_11092);
and U11813 (N_11813,N_10610,N_10875);
xnor U11814 (N_11814,N_10449,N_10971);
nand U11815 (N_11815,N_10969,N_10748);
or U11816 (N_11816,N_11095,N_10867);
nor U11817 (N_11817,N_10925,N_10953);
or U11818 (N_11818,N_11092,N_10785);
nor U11819 (N_11819,N_11050,N_10427);
nand U11820 (N_11820,N_10573,N_10915);
nor U11821 (N_11821,N_10710,N_10630);
or U11822 (N_11822,N_11065,N_10623);
and U11823 (N_11823,N_10917,N_10636);
and U11824 (N_11824,N_10885,N_10615);
nand U11825 (N_11825,N_11018,N_10884);
or U11826 (N_11826,N_11103,N_10976);
nand U11827 (N_11827,N_11018,N_10838);
xor U11828 (N_11828,N_10971,N_11153);
nor U11829 (N_11829,N_11073,N_11180);
xor U11830 (N_11830,N_10846,N_10718);
xnor U11831 (N_11831,N_10512,N_10514);
and U11832 (N_11832,N_10851,N_10842);
xor U11833 (N_11833,N_10620,N_10665);
and U11834 (N_11834,N_11183,N_10826);
and U11835 (N_11835,N_10793,N_10909);
nand U11836 (N_11836,N_11044,N_10958);
nor U11837 (N_11837,N_10633,N_10648);
and U11838 (N_11838,N_10624,N_10988);
nand U11839 (N_11839,N_10905,N_10725);
and U11840 (N_11840,N_11059,N_11064);
or U11841 (N_11841,N_11181,N_10620);
or U11842 (N_11842,N_11023,N_11107);
nand U11843 (N_11843,N_10532,N_11067);
nand U11844 (N_11844,N_10721,N_10556);
nor U11845 (N_11845,N_10458,N_10932);
and U11846 (N_11846,N_11006,N_11108);
nor U11847 (N_11847,N_10671,N_10523);
nor U11848 (N_11848,N_11113,N_10624);
and U11849 (N_11849,N_10672,N_10476);
xnor U11850 (N_11850,N_11028,N_11155);
xor U11851 (N_11851,N_11169,N_11024);
or U11852 (N_11852,N_10770,N_10847);
xnor U11853 (N_11853,N_10571,N_10634);
nand U11854 (N_11854,N_10410,N_10894);
or U11855 (N_11855,N_10771,N_10870);
or U11856 (N_11856,N_10611,N_10615);
xor U11857 (N_11857,N_11100,N_11102);
and U11858 (N_11858,N_10913,N_10868);
and U11859 (N_11859,N_11092,N_11161);
or U11860 (N_11860,N_10676,N_10760);
nor U11861 (N_11861,N_10987,N_10564);
and U11862 (N_11862,N_10481,N_10926);
nor U11863 (N_11863,N_10502,N_10831);
and U11864 (N_11864,N_10953,N_10576);
nor U11865 (N_11865,N_10520,N_10478);
nor U11866 (N_11866,N_10636,N_10817);
or U11867 (N_11867,N_10613,N_10647);
nor U11868 (N_11868,N_10417,N_11059);
nand U11869 (N_11869,N_10419,N_10970);
or U11870 (N_11870,N_11090,N_11025);
xor U11871 (N_11871,N_10671,N_10882);
nor U11872 (N_11872,N_10516,N_10541);
nand U11873 (N_11873,N_10663,N_10903);
nor U11874 (N_11874,N_10728,N_11053);
or U11875 (N_11875,N_10542,N_11077);
or U11876 (N_11876,N_10561,N_10810);
or U11877 (N_11877,N_11058,N_10937);
and U11878 (N_11878,N_10540,N_11172);
nor U11879 (N_11879,N_10854,N_10597);
or U11880 (N_11880,N_10406,N_11133);
nor U11881 (N_11881,N_10816,N_11152);
or U11882 (N_11882,N_11116,N_10743);
nor U11883 (N_11883,N_10723,N_10772);
or U11884 (N_11884,N_10557,N_11034);
and U11885 (N_11885,N_11167,N_10857);
nand U11886 (N_11886,N_10869,N_10816);
or U11887 (N_11887,N_11041,N_10559);
xnor U11888 (N_11888,N_10943,N_10756);
nand U11889 (N_11889,N_10588,N_11163);
nor U11890 (N_11890,N_10976,N_10690);
and U11891 (N_11891,N_10975,N_10868);
nor U11892 (N_11892,N_10660,N_11099);
or U11893 (N_11893,N_11184,N_11193);
nand U11894 (N_11894,N_11028,N_10955);
or U11895 (N_11895,N_10611,N_10661);
nand U11896 (N_11896,N_10624,N_10511);
nand U11897 (N_11897,N_10920,N_11040);
nor U11898 (N_11898,N_10818,N_10916);
nand U11899 (N_11899,N_10964,N_10447);
xnor U11900 (N_11900,N_11139,N_10910);
xnor U11901 (N_11901,N_10718,N_11191);
xnor U11902 (N_11902,N_10867,N_11026);
xor U11903 (N_11903,N_10931,N_10676);
xor U11904 (N_11904,N_11128,N_11078);
xnor U11905 (N_11905,N_10706,N_11182);
xor U11906 (N_11906,N_10921,N_10410);
nor U11907 (N_11907,N_10603,N_10797);
or U11908 (N_11908,N_10984,N_10702);
or U11909 (N_11909,N_11095,N_11135);
nor U11910 (N_11910,N_10728,N_10758);
nand U11911 (N_11911,N_10410,N_10957);
nand U11912 (N_11912,N_10747,N_10850);
and U11913 (N_11913,N_10936,N_10604);
nor U11914 (N_11914,N_10918,N_11052);
xor U11915 (N_11915,N_10830,N_10627);
and U11916 (N_11916,N_10617,N_10573);
nand U11917 (N_11917,N_10784,N_11011);
nor U11918 (N_11918,N_10856,N_10649);
and U11919 (N_11919,N_11143,N_10589);
and U11920 (N_11920,N_10938,N_10584);
and U11921 (N_11921,N_10989,N_10953);
and U11922 (N_11922,N_11139,N_10639);
nand U11923 (N_11923,N_10926,N_10605);
xor U11924 (N_11924,N_11046,N_10965);
nand U11925 (N_11925,N_10881,N_10966);
and U11926 (N_11926,N_10774,N_11018);
and U11927 (N_11927,N_10448,N_11100);
nor U11928 (N_11928,N_11119,N_10606);
xor U11929 (N_11929,N_11045,N_10954);
nor U11930 (N_11930,N_10505,N_11044);
and U11931 (N_11931,N_10445,N_10479);
nor U11932 (N_11932,N_10746,N_10532);
nand U11933 (N_11933,N_10479,N_10977);
nor U11934 (N_11934,N_10816,N_11181);
nor U11935 (N_11935,N_10589,N_10722);
xor U11936 (N_11936,N_10459,N_10752);
nor U11937 (N_11937,N_10937,N_10687);
xnor U11938 (N_11938,N_11110,N_11078);
nor U11939 (N_11939,N_11012,N_10989);
nor U11940 (N_11940,N_10957,N_10951);
xnor U11941 (N_11941,N_10952,N_10858);
nor U11942 (N_11942,N_10967,N_10453);
and U11943 (N_11943,N_10716,N_11031);
and U11944 (N_11944,N_10668,N_10754);
nand U11945 (N_11945,N_10783,N_11184);
or U11946 (N_11946,N_10655,N_10873);
nand U11947 (N_11947,N_10967,N_11193);
nor U11948 (N_11948,N_11145,N_10831);
and U11949 (N_11949,N_10746,N_10614);
xnor U11950 (N_11950,N_10958,N_10873);
nand U11951 (N_11951,N_10566,N_10723);
and U11952 (N_11952,N_11112,N_11184);
or U11953 (N_11953,N_10467,N_10690);
nand U11954 (N_11954,N_11180,N_11022);
nand U11955 (N_11955,N_10628,N_10514);
nand U11956 (N_11956,N_10845,N_11089);
nand U11957 (N_11957,N_10782,N_10434);
xnor U11958 (N_11958,N_10626,N_10527);
or U11959 (N_11959,N_11039,N_11176);
or U11960 (N_11960,N_10519,N_11082);
or U11961 (N_11961,N_10696,N_11038);
or U11962 (N_11962,N_10911,N_11025);
and U11963 (N_11963,N_10916,N_10875);
and U11964 (N_11964,N_10403,N_11157);
nor U11965 (N_11965,N_10465,N_10872);
or U11966 (N_11966,N_10669,N_10887);
xor U11967 (N_11967,N_10544,N_11073);
and U11968 (N_11968,N_10995,N_10634);
nor U11969 (N_11969,N_10929,N_10922);
and U11970 (N_11970,N_11174,N_10596);
or U11971 (N_11971,N_11180,N_11190);
nor U11972 (N_11972,N_10847,N_10828);
xnor U11973 (N_11973,N_11040,N_10717);
nor U11974 (N_11974,N_10768,N_10832);
or U11975 (N_11975,N_10864,N_10429);
nand U11976 (N_11976,N_11020,N_11109);
xnor U11977 (N_11977,N_11195,N_10403);
nor U11978 (N_11978,N_10601,N_10665);
nand U11979 (N_11979,N_10520,N_10670);
or U11980 (N_11980,N_11087,N_10731);
nand U11981 (N_11981,N_10506,N_10989);
or U11982 (N_11982,N_10821,N_10966);
nand U11983 (N_11983,N_11006,N_10809);
and U11984 (N_11984,N_10825,N_10765);
or U11985 (N_11985,N_10784,N_10538);
nor U11986 (N_11986,N_11166,N_10861);
and U11987 (N_11987,N_10678,N_10507);
or U11988 (N_11988,N_10457,N_10587);
or U11989 (N_11989,N_11060,N_10851);
nand U11990 (N_11990,N_11056,N_10652);
nor U11991 (N_11991,N_10917,N_10942);
nor U11992 (N_11992,N_10995,N_10952);
nor U11993 (N_11993,N_10474,N_10986);
xnor U11994 (N_11994,N_10956,N_10973);
nor U11995 (N_11995,N_11168,N_10657);
nand U11996 (N_11996,N_11008,N_11012);
and U11997 (N_11997,N_10472,N_11041);
nor U11998 (N_11998,N_10966,N_10661);
xor U11999 (N_11999,N_10509,N_10909);
or U12000 (N_12000,N_11852,N_11816);
xnor U12001 (N_12001,N_11427,N_11666);
and U12002 (N_12002,N_11465,N_11429);
or U12003 (N_12003,N_11960,N_11447);
and U12004 (N_12004,N_11711,N_11347);
nor U12005 (N_12005,N_11872,N_11702);
nand U12006 (N_12006,N_11586,N_11863);
xnor U12007 (N_12007,N_11869,N_11395);
and U12008 (N_12008,N_11256,N_11599);
and U12009 (N_12009,N_11824,N_11630);
nor U12010 (N_12010,N_11368,N_11227);
xnor U12011 (N_12011,N_11953,N_11941);
and U12012 (N_12012,N_11309,N_11885);
xnor U12013 (N_12013,N_11353,N_11817);
xnor U12014 (N_12014,N_11637,N_11766);
nor U12015 (N_12015,N_11857,N_11482);
xnor U12016 (N_12016,N_11422,N_11237);
nor U12017 (N_12017,N_11278,N_11562);
nand U12018 (N_12018,N_11529,N_11588);
and U12019 (N_12019,N_11458,N_11999);
and U12020 (N_12020,N_11417,N_11846);
nor U12021 (N_12021,N_11547,N_11635);
and U12022 (N_12022,N_11412,N_11283);
and U12023 (N_12023,N_11831,N_11326);
nor U12024 (N_12024,N_11294,N_11284);
xor U12025 (N_12025,N_11856,N_11500);
and U12026 (N_12026,N_11829,N_11976);
or U12027 (N_12027,N_11553,N_11949);
nor U12028 (N_12028,N_11906,N_11834);
or U12029 (N_12029,N_11259,N_11552);
nor U12030 (N_12030,N_11689,N_11223);
nor U12031 (N_12031,N_11501,N_11997);
and U12032 (N_12032,N_11647,N_11518);
or U12033 (N_12033,N_11579,N_11312);
nand U12034 (N_12034,N_11234,N_11339);
nor U12035 (N_12035,N_11989,N_11905);
and U12036 (N_12036,N_11291,N_11491);
nand U12037 (N_12037,N_11937,N_11304);
nor U12038 (N_12038,N_11514,N_11334);
xor U12039 (N_12039,N_11979,N_11456);
nand U12040 (N_12040,N_11750,N_11715);
nand U12041 (N_12041,N_11254,N_11299);
nor U12042 (N_12042,N_11802,N_11649);
and U12043 (N_12043,N_11519,N_11536);
nand U12044 (N_12044,N_11230,N_11964);
nor U12045 (N_12045,N_11933,N_11463);
or U12046 (N_12046,N_11844,N_11765);
nor U12047 (N_12047,N_11571,N_11365);
and U12048 (N_12048,N_11202,N_11469);
or U12049 (N_12049,N_11685,N_11495);
nor U12050 (N_12050,N_11927,N_11681);
nor U12051 (N_12051,N_11734,N_11433);
nor U12052 (N_12052,N_11951,N_11523);
nor U12053 (N_12053,N_11669,N_11542);
nand U12054 (N_12054,N_11873,N_11452);
nand U12055 (N_12055,N_11483,N_11874);
and U12056 (N_12056,N_11535,N_11930);
or U12057 (N_12057,N_11531,N_11358);
and U12058 (N_12058,N_11288,N_11628);
nand U12059 (N_12059,N_11585,N_11748);
xnor U12060 (N_12060,N_11321,N_11867);
or U12061 (N_12061,N_11503,N_11459);
xnor U12062 (N_12062,N_11485,N_11426);
and U12063 (N_12063,N_11892,N_11674);
nand U12064 (N_12064,N_11292,N_11855);
nor U12065 (N_12065,N_11767,N_11664);
nor U12066 (N_12066,N_11981,N_11779);
nand U12067 (N_12067,N_11958,N_11573);
xnor U12068 (N_12068,N_11592,N_11773);
or U12069 (N_12069,N_11807,N_11225);
nor U12070 (N_12070,N_11467,N_11258);
or U12071 (N_12071,N_11827,N_11330);
xor U12072 (N_12072,N_11760,N_11377);
and U12073 (N_12073,N_11904,N_11663);
and U12074 (N_12074,N_11604,N_11203);
or U12075 (N_12075,N_11286,N_11741);
and U12076 (N_12076,N_11771,N_11735);
xor U12077 (N_12077,N_11565,N_11696);
and U12078 (N_12078,N_11655,N_11612);
nor U12079 (N_12079,N_11934,N_11595);
nand U12080 (N_12080,N_11893,N_11860);
nor U12081 (N_12081,N_11252,N_11774);
or U12082 (N_12082,N_11583,N_11790);
nor U12083 (N_12083,N_11875,N_11320);
and U12084 (N_12084,N_11820,N_11492);
or U12085 (N_12085,N_11877,N_11854);
and U12086 (N_12086,N_11224,N_11477);
and U12087 (N_12087,N_11376,N_11371);
or U12088 (N_12088,N_11293,N_11564);
nand U12089 (N_12089,N_11453,N_11889);
xor U12090 (N_12090,N_11727,N_11880);
or U12091 (N_12091,N_11680,N_11200);
and U12092 (N_12092,N_11399,N_11724);
and U12093 (N_12093,N_11446,N_11902);
xor U12094 (N_12094,N_11327,N_11440);
xor U12095 (N_12095,N_11757,N_11903);
or U12096 (N_12096,N_11563,N_11716);
xnor U12097 (N_12097,N_11928,N_11437);
and U12098 (N_12098,N_11204,N_11273);
nor U12099 (N_12099,N_11918,N_11838);
or U12100 (N_12100,N_11944,N_11788);
xor U12101 (N_12101,N_11546,N_11526);
nand U12102 (N_12102,N_11493,N_11801);
nand U12103 (N_12103,N_11795,N_11848);
nand U12104 (N_12104,N_11859,N_11761);
nand U12105 (N_12105,N_11512,N_11822);
and U12106 (N_12106,N_11797,N_11209);
nand U12107 (N_12107,N_11584,N_11349);
nor U12108 (N_12108,N_11386,N_11700);
or U12109 (N_12109,N_11865,N_11919);
nand U12110 (N_12110,N_11645,N_11550);
nor U12111 (N_12111,N_11528,N_11736);
and U12112 (N_12112,N_11993,N_11271);
or U12113 (N_12113,N_11504,N_11616);
nand U12114 (N_12114,N_11614,N_11609);
nand U12115 (N_12115,N_11778,N_11484);
xor U12116 (N_12116,N_11231,N_11781);
nor U12117 (N_12117,N_11434,N_11322);
or U12118 (N_12118,N_11843,N_11354);
nand U12119 (N_12119,N_11749,N_11594);
and U12120 (N_12120,N_11533,N_11699);
or U12121 (N_12121,N_11888,N_11487);
nand U12122 (N_12122,N_11946,N_11360);
nor U12123 (N_12123,N_11789,N_11551);
and U12124 (N_12124,N_11445,N_11763);
xor U12125 (N_12125,N_11963,N_11602);
nor U12126 (N_12126,N_11346,N_11608);
nand U12127 (N_12127,N_11603,N_11280);
xor U12128 (N_12128,N_11894,N_11662);
and U12129 (N_12129,N_11506,N_11210);
xor U12130 (N_12130,N_11733,N_11443);
xor U12131 (N_12131,N_11744,N_11671);
nor U12132 (N_12132,N_11532,N_11522);
nor U12133 (N_12133,N_11241,N_11460);
nand U12134 (N_12134,N_11842,N_11678);
nor U12135 (N_12135,N_11511,N_11796);
nor U12136 (N_12136,N_11943,N_11675);
nor U12137 (N_12137,N_11298,N_11995);
or U12138 (N_12138,N_11538,N_11653);
and U12139 (N_12139,N_11220,N_11502);
or U12140 (N_12140,N_11208,N_11871);
or U12141 (N_12141,N_11998,N_11690);
or U12142 (N_12142,N_11650,N_11593);
nor U12143 (N_12143,N_11701,N_11677);
xnor U12144 (N_12144,N_11505,N_11264);
nor U12145 (N_12145,N_11479,N_11425);
and U12146 (N_12146,N_11707,N_11922);
and U12147 (N_12147,N_11303,N_11554);
or U12148 (N_12148,N_11540,N_11296);
nor U12149 (N_12149,N_11777,N_11580);
or U12150 (N_12150,N_11686,N_11862);
nand U12151 (N_12151,N_11403,N_11361);
and U12152 (N_12152,N_11290,N_11544);
and U12153 (N_12153,N_11367,N_11896);
and U12154 (N_12154,N_11887,N_11978);
and U12155 (N_12155,N_11739,N_11809);
or U12156 (N_12156,N_11833,N_11950);
nor U12157 (N_12157,N_11435,N_11398);
or U12158 (N_12158,N_11670,N_11516);
and U12159 (N_12159,N_11442,N_11858);
or U12160 (N_12160,N_11601,N_11768);
or U12161 (N_12161,N_11965,N_11570);
or U12162 (N_12162,N_11694,N_11471);
nand U12163 (N_12163,N_11814,N_11745);
and U12164 (N_12164,N_11996,N_11620);
and U12165 (N_12165,N_11936,N_11449);
nor U12166 (N_12166,N_11784,N_11692);
nand U12167 (N_12167,N_11421,N_11404);
and U12168 (N_12168,N_11718,N_11955);
nand U12169 (N_12169,N_11821,N_11306);
nor U12170 (N_12170,N_11819,N_11362);
nand U12171 (N_12171,N_11391,N_11730);
nand U12172 (N_12172,N_11380,N_11883);
or U12173 (N_12173,N_11242,N_11394);
nor U12174 (N_12174,N_11229,N_11626);
or U12175 (N_12175,N_11929,N_11703);
nor U12176 (N_12176,N_11697,N_11818);
or U12177 (N_12177,N_11845,N_11792);
nor U12178 (N_12178,N_11597,N_11295);
nand U12179 (N_12179,N_11269,N_11629);
and U12180 (N_12180,N_11695,N_11832);
nand U12181 (N_12181,N_11268,N_11917);
nor U12182 (N_12182,N_11219,N_11474);
and U12183 (N_12183,N_11967,N_11742);
and U12184 (N_12184,N_11324,N_11769);
nor U12185 (N_12185,N_11984,N_11201);
nand U12186 (N_12186,N_11966,N_11509);
or U12187 (N_12187,N_11355,N_11959);
xnor U12188 (N_12188,N_11450,N_11644);
nor U12189 (N_12189,N_11351,N_11559);
nand U12190 (N_12190,N_11555,N_11436);
xnor U12191 (N_12191,N_11406,N_11706);
xnor U12192 (N_12192,N_11798,N_11232);
or U12193 (N_12193,N_11397,N_11357);
xnor U12194 (N_12194,N_11444,N_11390);
nand U12195 (N_12195,N_11924,N_11221);
xnor U12196 (N_12196,N_11962,N_11841);
xor U12197 (N_12197,N_11667,N_11261);
nor U12198 (N_12198,N_11383,N_11302);
and U12199 (N_12199,N_11378,N_11384);
nor U12200 (N_12200,N_11823,N_11751);
nand U12201 (N_12201,N_11881,N_11957);
nand U12202 (N_12202,N_11607,N_11336);
nor U12203 (N_12203,N_11255,N_11462);
and U12204 (N_12204,N_11238,N_11714);
and U12205 (N_12205,N_11372,N_11250);
or U12206 (N_12206,N_11407,N_11762);
and U12207 (N_12207,N_11517,N_11828);
and U12208 (N_12208,N_11494,N_11420);
or U12209 (N_12209,N_11366,N_11359);
nor U12210 (N_12210,N_11277,N_11772);
nand U12211 (N_12211,N_11646,N_11691);
nor U12212 (N_12212,N_11515,N_11900);
nand U12213 (N_12213,N_11611,N_11414);
nor U12214 (N_12214,N_11396,N_11343);
xnor U12215 (N_12215,N_11676,N_11679);
or U12216 (N_12216,N_11605,N_11415);
nand U12217 (N_12217,N_11931,N_11432);
xor U12218 (N_12218,N_11222,N_11882);
xnor U12219 (N_12219,N_11982,N_11786);
nand U12220 (N_12220,N_11267,N_11791);
or U12221 (N_12221,N_11890,N_11665);
nand U12222 (N_12222,N_11537,N_11246);
xor U12223 (N_12223,N_11805,N_11262);
nand U12224 (N_12224,N_11297,N_11861);
or U12225 (N_12225,N_11693,N_11379);
and U12226 (N_12226,N_11980,N_11738);
nand U12227 (N_12227,N_11634,N_11940);
nand U12228 (N_12228,N_11683,N_11496);
nor U12229 (N_12229,N_11581,N_11338);
nand U12230 (N_12230,N_11932,N_11329);
nor U12231 (N_12231,N_11521,N_11475);
nor U12232 (N_12232,N_11206,N_11840);
or U12233 (N_12233,N_11804,N_11549);
nor U12234 (N_12234,N_11853,N_11454);
and U12235 (N_12235,N_11582,N_11698);
nand U12236 (N_12236,N_11388,N_11729);
nor U12237 (N_12237,N_11720,N_11534);
nand U12238 (N_12238,N_11651,N_11236);
nand U12239 (N_12239,N_11332,N_11249);
nand U12240 (N_12240,N_11560,N_11808);
nand U12241 (N_12241,N_11658,N_11480);
and U12242 (N_12242,N_11335,N_11948);
xor U12243 (N_12243,N_11244,N_11619);
xnor U12244 (N_12244,N_11636,N_11561);
xor U12245 (N_12245,N_11746,N_11279);
or U12246 (N_12246,N_11287,N_11418);
and U12247 (N_12247,N_11615,N_11215);
xnor U12248 (N_12248,N_11891,N_11657);
nor U12249 (N_12249,N_11864,N_11837);
nand U12250 (N_12250,N_11214,N_11305);
or U12251 (N_12251,N_11408,N_11970);
nor U12252 (N_12252,N_11587,N_11316);
nor U12253 (N_12253,N_11405,N_11466);
and U12254 (N_12254,N_11728,N_11393);
nand U12255 (N_12255,N_11525,N_11990);
nand U12256 (N_12256,N_11668,N_11622);
nor U12257 (N_12257,N_11569,N_11775);
nor U12258 (N_12258,N_11382,N_11755);
xor U12259 (N_12259,N_11470,N_11884);
nor U12260 (N_12260,N_11387,N_11627);
and U12261 (N_12261,N_11567,N_11969);
nand U12262 (N_12262,N_11638,N_11704);
xnor U12263 (N_12263,N_11276,N_11617);
or U12264 (N_12264,N_11596,N_11411);
nand U12265 (N_12265,N_11914,N_11935);
nand U12266 (N_12266,N_11926,N_11764);
and U12267 (N_12267,N_11527,N_11815);
xnor U12268 (N_12268,N_11974,N_11218);
nor U12269 (N_12269,N_11961,N_11606);
or U12270 (N_12270,N_11508,N_11987);
nand U12271 (N_12271,N_11524,N_11468);
nand U12272 (N_12272,N_11441,N_11886);
nor U12273 (N_12273,N_11737,N_11373);
and U12274 (N_12274,N_11991,N_11826);
nand U12275 (N_12275,N_11239,N_11289);
and U12276 (N_12276,N_11688,N_11731);
nand U12277 (N_12277,N_11257,N_11954);
nor U12278 (N_12278,N_11956,N_11812);
and U12279 (N_12279,N_11705,N_11374);
nand U12280 (N_12280,N_11793,N_11717);
nor U12281 (N_12281,N_11633,N_11545);
and U12282 (N_12282,N_11660,N_11656);
and U12283 (N_12283,N_11925,N_11451);
xnor U12284 (N_12284,N_11947,N_11975);
nor U12285 (N_12285,N_11624,N_11541);
and U12286 (N_12286,N_11275,N_11212);
nor U12287 (N_12287,N_11901,N_11988);
or U12288 (N_12288,N_11598,N_11274);
or U12289 (N_12289,N_11590,N_11687);
xnor U12290 (N_12290,N_11909,N_11331);
or U12291 (N_12291,N_11270,N_11486);
or U12292 (N_12292,N_11578,N_11879);
nand U12293 (N_12293,N_11785,N_11759);
or U12294 (N_12294,N_11575,N_11621);
xnor U12295 (N_12295,N_11803,N_11345);
nand U12296 (N_12296,N_11248,N_11640);
and U12297 (N_12297,N_11253,N_11472);
and U12298 (N_12298,N_11307,N_11591);
nor U12299 (N_12299,N_11301,N_11643);
xnor U12300 (N_12300,N_11740,N_11401);
and U12301 (N_12301,N_11912,N_11548);
xnor U12302 (N_12302,N_11806,N_11648);
or U12303 (N_12303,N_11473,N_11839);
nor U12304 (N_12304,N_11363,N_11313);
nand U12305 (N_12305,N_11226,N_11310);
xnor U12306 (N_12306,N_11318,N_11850);
and U12307 (N_12307,N_11708,N_11770);
nor U12308 (N_12308,N_11281,N_11455);
nand U12309 (N_12309,N_11642,N_11323);
and U12310 (N_12310,N_11375,N_11977);
or U12311 (N_12311,N_11752,N_11568);
and U12312 (N_12312,N_11625,N_11285);
xnor U12313 (N_12313,N_11726,N_11481);
and U12314 (N_12314,N_11572,N_11866);
nor U12315 (N_12315,N_11240,N_11464);
xnor U12316 (N_12316,N_11488,N_11211);
nor U12317 (N_12317,N_11497,N_11847);
nand U12318 (N_12318,N_11836,N_11251);
nand U12319 (N_12319,N_11920,N_11328);
xor U12320 (N_12320,N_11897,N_11973);
and U12321 (N_12321,N_11849,N_11782);
nor U12322 (N_12322,N_11341,N_11350);
xor U12323 (N_12323,N_11217,N_11992);
or U12324 (N_12324,N_11983,N_11409);
nor U12325 (N_12325,N_11754,N_11876);
nand U12326 (N_12326,N_11513,N_11282);
nand U12327 (N_12327,N_11870,N_11672);
nand U12328 (N_12328,N_11205,N_11907);
nor U12329 (N_12329,N_11364,N_11566);
and U12330 (N_12330,N_11756,N_11659);
and U12331 (N_12331,N_11228,N_11913);
or U12332 (N_12332,N_11424,N_11923);
nand U12333 (N_12333,N_11461,N_11558);
nand U12334 (N_12334,N_11416,N_11207);
and U12335 (N_12335,N_11314,N_11337);
nor U12336 (N_12336,N_11813,N_11402);
and U12337 (N_12337,N_11972,N_11719);
and U12338 (N_12338,N_11722,N_11641);
and U12339 (N_12339,N_11631,N_11448);
nand U12340 (N_12340,N_11392,N_11457);
nand U12341 (N_12341,N_11899,N_11352);
nand U12342 (N_12342,N_11213,N_11723);
nand U12343 (N_12343,N_11787,N_11985);
nand U12344 (N_12344,N_11780,N_11308);
nor U12345 (N_12345,N_11776,N_11945);
and U12346 (N_12346,N_11431,N_11243);
and U12347 (N_12347,N_11325,N_11410);
nor U12348 (N_12348,N_11916,N_11911);
nand U12349 (N_12349,N_11340,N_11939);
nand U12350 (N_12350,N_11247,N_11613);
and U12351 (N_12351,N_11413,N_11272);
nand U12352 (N_12352,N_11618,N_11489);
and U12353 (N_12353,N_11898,N_11216);
nand U12354 (N_12354,N_11725,N_11265);
nand U12355 (N_12355,N_11794,N_11713);
and U12356 (N_12356,N_11673,N_11344);
or U12357 (N_12357,N_11577,N_11556);
and U12358 (N_12358,N_11758,N_11348);
nand U12359 (N_12359,N_11732,N_11311);
or U12360 (N_12360,N_11721,N_11610);
and U12361 (N_12361,N_11539,N_11747);
nor U12362 (N_12362,N_11825,N_11895);
nand U12363 (N_12363,N_11600,N_11799);
or U12364 (N_12364,N_11423,N_11652);
or U12365 (N_12365,N_11300,N_11942);
or U12366 (N_12366,N_11263,N_11968);
or U12367 (N_12367,N_11811,N_11661);
nand U12368 (N_12368,N_11428,N_11589);
nand U12369 (N_12369,N_11419,N_11810);
nand U12370 (N_12370,N_11430,N_11632);
and U12371 (N_12371,N_11233,N_11576);
nor U12372 (N_12372,N_11476,N_11682);
nand U12373 (N_12373,N_11499,N_11342);
or U12374 (N_12374,N_11385,N_11910);
nor U12375 (N_12375,N_11439,N_11938);
nor U12376 (N_12376,N_11319,N_11507);
nor U12377 (N_12377,N_11356,N_11709);
and U12378 (N_12378,N_11878,N_11915);
or U12379 (N_12379,N_11800,N_11952);
and U12380 (N_12380,N_11245,N_11317);
and U12381 (N_12381,N_11753,N_11490);
and U12382 (N_12382,N_11835,N_11830);
or U12383 (N_12383,N_11623,N_11315);
xor U12384 (N_12384,N_11557,N_11266);
nor U12385 (N_12385,N_11986,N_11369);
nand U12386 (N_12386,N_11478,N_11921);
or U12387 (N_12387,N_11389,N_11400);
or U12388 (N_12388,N_11438,N_11260);
or U12389 (N_12389,N_11574,N_11520);
and U12390 (N_12390,N_11851,N_11712);
or U12391 (N_12391,N_11639,N_11333);
nor U12392 (N_12392,N_11684,N_11381);
xnor U12393 (N_12393,N_11994,N_11235);
and U12394 (N_12394,N_11743,N_11498);
xor U12395 (N_12395,N_11543,N_11868);
nor U12396 (N_12396,N_11908,N_11971);
nand U12397 (N_12397,N_11654,N_11783);
or U12398 (N_12398,N_11370,N_11530);
or U12399 (N_12399,N_11510,N_11710);
or U12400 (N_12400,N_11303,N_11202);
or U12401 (N_12401,N_11812,N_11390);
nor U12402 (N_12402,N_11752,N_11837);
and U12403 (N_12403,N_11739,N_11414);
and U12404 (N_12404,N_11520,N_11940);
xnor U12405 (N_12405,N_11212,N_11622);
xnor U12406 (N_12406,N_11278,N_11627);
nand U12407 (N_12407,N_11210,N_11542);
nor U12408 (N_12408,N_11721,N_11293);
xor U12409 (N_12409,N_11687,N_11426);
and U12410 (N_12410,N_11378,N_11272);
or U12411 (N_12411,N_11412,N_11519);
nor U12412 (N_12412,N_11224,N_11872);
nor U12413 (N_12413,N_11446,N_11315);
or U12414 (N_12414,N_11489,N_11544);
nand U12415 (N_12415,N_11545,N_11978);
nor U12416 (N_12416,N_11988,N_11999);
nor U12417 (N_12417,N_11808,N_11674);
nand U12418 (N_12418,N_11276,N_11331);
nor U12419 (N_12419,N_11338,N_11610);
nor U12420 (N_12420,N_11328,N_11417);
xnor U12421 (N_12421,N_11905,N_11250);
or U12422 (N_12422,N_11330,N_11984);
nand U12423 (N_12423,N_11284,N_11807);
or U12424 (N_12424,N_11257,N_11534);
xor U12425 (N_12425,N_11942,N_11894);
xor U12426 (N_12426,N_11800,N_11778);
and U12427 (N_12427,N_11468,N_11668);
xor U12428 (N_12428,N_11742,N_11583);
nand U12429 (N_12429,N_11847,N_11662);
or U12430 (N_12430,N_11620,N_11464);
and U12431 (N_12431,N_11775,N_11856);
nor U12432 (N_12432,N_11529,N_11858);
nor U12433 (N_12433,N_11217,N_11810);
nand U12434 (N_12434,N_11887,N_11850);
nor U12435 (N_12435,N_11892,N_11890);
or U12436 (N_12436,N_11562,N_11779);
nand U12437 (N_12437,N_11286,N_11714);
nand U12438 (N_12438,N_11546,N_11554);
xor U12439 (N_12439,N_11471,N_11375);
or U12440 (N_12440,N_11970,N_11356);
nor U12441 (N_12441,N_11989,N_11834);
nor U12442 (N_12442,N_11531,N_11863);
xor U12443 (N_12443,N_11391,N_11804);
and U12444 (N_12444,N_11788,N_11868);
nor U12445 (N_12445,N_11975,N_11985);
nand U12446 (N_12446,N_11472,N_11770);
nand U12447 (N_12447,N_11735,N_11683);
nor U12448 (N_12448,N_11832,N_11965);
or U12449 (N_12449,N_11748,N_11557);
xnor U12450 (N_12450,N_11562,N_11858);
xor U12451 (N_12451,N_11464,N_11666);
and U12452 (N_12452,N_11911,N_11577);
and U12453 (N_12453,N_11851,N_11580);
xnor U12454 (N_12454,N_11617,N_11512);
and U12455 (N_12455,N_11437,N_11304);
or U12456 (N_12456,N_11353,N_11521);
or U12457 (N_12457,N_11536,N_11570);
xnor U12458 (N_12458,N_11717,N_11281);
and U12459 (N_12459,N_11800,N_11320);
nor U12460 (N_12460,N_11204,N_11478);
and U12461 (N_12461,N_11880,N_11213);
or U12462 (N_12462,N_11232,N_11332);
nor U12463 (N_12463,N_11918,N_11473);
and U12464 (N_12464,N_11682,N_11809);
or U12465 (N_12465,N_11974,N_11396);
xnor U12466 (N_12466,N_11840,N_11637);
xor U12467 (N_12467,N_11342,N_11206);
and U12468 (N_12468,N_11620,N_11357);
or U12469 (N_12469,N_11687,N_11293);
and U12470 (N_12470,N_11543,N_11956);
and U12471 (N_12471,N_11925,N_11358);
and U12472 (N_12472,N_11236,N_11278);
and U12473 (N_12473,N_11617,N_11846);
and U12474 (N_12474,N_11623,N_11609);
and U12475 (N_12475,N_11529,N_11242);
xnor U12476 (N_12476,N_11259,N_11901);
nor U12477 (N_12477,N_11603,N_11529);
nand U12478 (N_12478,N_11308,N_11318);
or U12479 (N_12479,N_11561,N_11445);
and U12480 (N_12480,N_11799,N_11961);
xor U12481 (N_12481,N_11900,N_11930);
or U12482 (N_12482,N_11902,N_11746);
or U12483 (N_12483,N_11420,N_11256);
and U12484 (N_12484,N_11333,N_11311);
xor U12485 (N_12485,N_11460,N_11506);
nand U12486 (N_12486,N_11303,N_11224);
nor U12487 (N_12487,N_11565,N_11236);
xor U12488 (N_12488,N_11345,N_11944);
xor U12489 (N_12489,N_11606,N_11490);
and U12490 (N_12490,N_11657,N_11560);
nand U12491 (N_12491,N_11832,N_11924);
xnor U12492 (N_12492,N_11461,N_11436);
nor U12493 (N_12493,N_11513,N_11339);
or U12494 (N_12494,N_11743,N_11352);
nor U12495 (N_12495,N_11578,N_11260);
nor U12496 (N_12496,N_11794,N_11885);
xor U12497 (N_12497,N_11275,N_11557);
xor U12498 (N_12498,N_11616,N_11227);
nor U12499 (N_12499,N_11730,N_11453);
xnor U12500 (N_12500,N_11911,N_11720);
xnor U12501 (N_12501,N_11932,N_11995);
nand U12502 (N_12502,N_11911,N_11948);
nor U12503 (N_12503,N_11249,N_11231);
or U12504 (N_12504,N_11841,N_11663);
xnor U12505 (N_12505,N_11780,N_11507);
nor U12506 (N_12506,N_11493,N_11466);
and U12507 (N_12507,N_11781,N_11580);
and U12508 (N_12508,N_11592,N_11782);
nand U12509 (N_12509,N_11567,N_11622);
and U12510 (N_12510,N_11454,N_11313);
and U12511 (N_12511,N_11531,N_11359);
or U12512 (N_12512,N_11823,N_11546);
nand U12513 (N_12513,N_11412,N_11373);
nor U12514 (N_12514,N_11794,N_11633);
nand U12515 (N_12515,N_11867,N_11695);
xor U12516 (N_12516,N_11479,N_11821);
or U12517 (N_12517,N_11311,N_11475);
xnor U12518 (N_12518,N_11859,N_11736);
xnor U12519 (N_12519,N_11674,N_11898);
xnor U12520 (N_12520,N_11866,N_11353);
nand U12521 (N_12521,N_11523,N_11324);
and U12522 (N_12522,N_11312,N_11581);
xnor U12523 (N_12523,N_11300,N_11705);
nand U12524 (N_12524,N_11304,N_11486);
nand U12525 (N_12525,N_11700,N_11729);
or U12526 (N_12526,N_11531,N_11993);
nand U12527 (N_12527,N_11552,N_11844);
xnor U12528 (N_12528,N_11466,N_11814);
xnor U12529 (N_12529,N_11572,N_11600);
nand U12530 (N_12530,N_11828,N_11753);
nor U12531 (N_12531,N_11873,N_11788);
nand U12532 (N_12532,N_11321,N_11885);
xor U12533 (N_12533,N_11740,N_11500);
nand U12534 (N_12534,N_11757,N_11876);
xnor U12535 (N_12535,N_11646,N_11989);
or U12536 (N_12536,N_11725,N_11490);
nor U12537 (N_12537,N_11295,N_11871);
xnor U12538 (N_12538,N_11332,N_11798);
and U12539 (N_12539,N_11567,N_11812);
xor U12540 (N_12540,N_11946,N_11426);
or U12541 (N_12541,N_11751,N_11933);
xnor U12542 (N_12542,N_11408,N_11619);
or U12543 (N_12543,N_11886,N_11303);
nor U12544 (N_12544,N_11793,N_11329);
nor U12545 (N_12545,N_11924,N_11567);
or U12546 (N_12546,N_11573,N_11438);
nand U12547 (N_12547,N_11494,N_11328);
or U12548 (N_12548,N_11837,N_11937);
nor U12549 (N_12549,N_11591,N_11514);
nand U12550 (N_12550,N_11202,N_11428);
or U12551 (N_12551,N_11879,N_11413);
nand U12552 (N_12552,N_11589,N_11679);
xor U12553 (N_12553,N_11809,N_11763);
or U12554 (N_12554,N_11245,N_11908);
or U12555 (N_12555,N_11418,N_11377);
and U12556 (N_12556,N_11648,N_11529);
nor U12557 (N_12557,N_11542,N_11788);
nor U12558 (N_12558,N_11219,N_11392);
nor U12559 (N_12559,N_11447,N_11733);
nand U12560 (N_12560,N_11766,N_11878);
or U12561 (N_12561,N_11410,N_11750);
nor U12562 (N_12562,N_11609,N_11767);
or U12563 (N_12563,N_11534,N_11221);
nand U12564 (N_12564,N_11718,N_11686);
and U12565 (N_12565,N_11829,N_11468);
xor U12566 (N_12566,N_11202,N_11955);
nor U12567 (N_12567,N_11714,N_11698);
or U12568 (N_12568,N_11214,N_11997);
nor U12569 (N_12569,N_11962,N_11407);
nor U12570 (N_12570,N_11307,N_11956);
nand U12571 (N_12571,N_11946,N_11270);
nor U12572 (N_12572,N_11380,N_11879);
or U12573 (N_12573,N_11753,N_11384);
nor U12574 (N_12574,N_11299,N_11361);
or U12575 (N_12575,N_11257,N_11336);
nand U12576 (N_12576,N_11498,N_11590);
and U12577 (N_12577,N_11384,N_11497);
nor U12578 (N_12578,N_11662,N_11326);
nor U12579 (N_12579,N_11385,N_11873);
and U12580 (N_12580,N_11275,N_11373);
nand U12581 (N_12581,N_11548,N_11519);
nand U12582 (N_12582,N_11570,N_11382);
nand U12583 (N_12583,N_11357,N_11309);
nand U12584 (N_12584,N_11757,N_11921);
nor U12585 (N_12585,N_11553,N_11401);
xnor U12586 (N_12586,N_11431,N_11937);
nor U12587 (N_12587,N_11223,N_11989);
nor U12588 (N_12588,N_11702,N_11777);
xor U12589 (N_12589,N_11959,N_11552);
nor U12590 (N_12590,N_11686,N_11609);
xor U12591 (N_12591,N_11737,N_11220);
and U12592 (N_12592,N_11438,N_11983);
or U12593 (N_12593,N_11575,N_11395);
and U12594 (N_12594,N_11583,N_11396);
nand U12595 (N_12595,N_11512,N_11670);
or U12596 (N_12596,N_11461,N_11571);
xnor U12597 (N_12597,N_11932,N_11711);
nand U12598 (N_12598,N_11442,N_11664);
and U12599 (N_12599,N_11537,N_11271);
and U12600 (N_12600,N_11248,N_11267);
or U12601 (N_12601,N_11249,N_11838);
nand U12602 (N_12602,N_11265,N_11598);
nand U12603 (N_12603,N_11857,N_11514);
and U12604 (N_12604,N_11929,N_11373);
nor U12605 (N_12605,N_11690,N_11719);
and U12606 (N_12606,N_11680,N_11265);
nand U12607 (N_12607,N_11245,N_11348);
xor U12608 (N_12608,N_11922,N_11666);
nand U12609 (N_12609,N_11371,N_11794);
nand U12610 (N_12610,N_11541,N_11970);
and U12611 (N_12611,N_11278,N_11427);
xor U12612 (N_12612,N_11819,N_11619);
nand U12613 (N_12613,N_11694,N_11937);
or U12614 (N_12614,N_11540,N_11649);
nand U12615 (N_12615,N_11728,N_11915);
nor U12616 (N_12616,N_11544,N_11563);
nand U12617 (N_12617,N_11986,N_11722);
xor U12618 (N_12618,N_11761,N_11319);
nor U12619 (N_12619,N_11542,N_11373);
or U12620 (N_12620,N_11204,N_11897);
and U12621 (N_12621,N_11387,N_11793);
nand U12622 (N_12622,N_11360,N_11400);
and U12623 (N_12623,N_11625,N_11841);
nor U12624 (N_12624,N_11436,N_11590);
and U12625 (N_12625,N_11751,N_11574);
and U12626 (N_12626,N_11925,N_11459);
and U12627 (N_12627,N_11725,N_11776);
or U12628 (N_12628,N_11247,N_11255);
and U12629 (N_12629,N_11243,N_11280);
xnor U12630 (N_12630,N_11857,N_11827);
nand U12631 (N_12631,N_11237,N_11486);
nor U12632 (N_12632,N_11582,N_11232);
and U12633 (N_12633,N_11283,N_11554);
or U12634 (N_12634,N_11757,N_11216);
nand U12635 (N_12635,N_11374,N_11757);
nor U12636 (N_12636,N_11979,N_11732);
nor U12637 (N_12637,N_11919,N_11718);
nor U12638 (N_12638,N_11497,N_11653);
xor U12639 (N_12639,N_11784,N_11625);
or U12640 (N_12640,N_11288,N_11458);
xnor U12641 (N_12641,N_11320,N_11725);
nand U12642 (N_12642,N_11316,N_11266);
or U12643 (N_12643,N_11778,N_11281);
or U12644 (N_12644,N_11517,N_11822);
and U12645 (N_12645,N_11473,N_11516);
and U12646 (N_12646,N_11478,N_11618);
and U12647 (N_12647,N_11877,N_11507);
and U12648 (N_12648,N_11541,N_11661);
nand U12649 (N_12649,N_11358,N_11841);
nand U12650 (N_12650,N_11507,N_11598);
or U12651 (N_12651,N_11224,N_11358);
or U12652 (N_12652,N_11254,N_11336);
xnor U12653 (N_12653,N_11557,N_11903);
or U12654 (N_12654,N_11786,N_11385);
nand U12655 (N_12655,N_11487,N_11629);
xor U12656 (N_12656,N_11645,N_11634);
nand U12657 (N_12657,N_11953,N_11282);
and U12658 (N_12658,N_11612,N_11694);
nand U12659 (N_12659,N_11889,N_11452);
and U12660 (N_12660,N_11951,N_11994);
xnor U12661 (N_12661,N_11799,N_11972);
nand U12662 (N_12662,N_11945,N_11432);
or U12663 (N_12663,N_11628,N_11402);
xor U12664 (N_12664,N_11785,N_11709);
nand U12665 (N_12665,N_11324,N_11315);
nor U12666 (N_12666,N_11979,N_11285);
nand U12667 (N_12667,N_11547,N_11891);
or U12668 (N_12668,N_11769,N_11415);
nand U12669 (N_12669,N_11305,N_11355);
or U12670 (N_12670,N_11509,N_11847);
nor U12671 (N_12671,N_11440,N_11671);
or U12672 (N_12672,N_11576,N_11380);
or U12673 (N_12673,N_11451,N_11225);
or U12674 (N_12674,N_11505,N_11625);
nor U12675 (N_12675,N_11273,N_11481);
or U12676 (N_12676,N_11400,N_11566);
xor U12677 (N_12677,N_11212,N_11835);
nor U12678 (N_12678,N_11670,N_11757);
nand U12679 (N_12679,N_11217,N_11466);
or U12680 (N_12680,N_11881,N_11847);
and U12681 (N_12681,N_11479,N_11961);
xnor U12682 (N_12682,N_11540,N_11428);
and U12683 (N_12683,N_11402,N_11558);
xor U12684 (N_12684,N_11969,N_11655);
nand U12685 (N_12685,N_11636,N_11897);
and U12686 (N_12686,N_11723,N_11796);
and U12687 (N_12687,N_11631,N_11718);
and U12688 (N_12688,N_11214,N_11354);
or U12689 (N_12689,N_11479,N_11701);
xor U12690 (N_12690,N_11606,N_11271);
nand U12691 (N_12691,N_11642,N_11919);
xnor U12692 (N_12692,N_11322,N_11425);
or U12693 (N_12693,N_11953,N_11469);
and U12694 (N_12694,N_11927,N_11263);
or U12695 (N_12695,N_11483,N_11715);
nor U12696 (N_12696,N_11509,N_11332);
and U12697 (N_12697,N_11425,N_11521);
and U12698 (N_12698,N_11422,N_11654);
or U12699 (N_12699,N_11780,N_11325);
or U12700 (N_12700,N_11248,N_11935);
nand U12701 (N_12701,N_11224,N_11689);
or U12702 (N_12702,N_11347,N_11443);
and U12703 (N_12703,N_11570,N_11738);
or U12704 (N_12704,N_11331,N_11608);
and U12705 (N_12705,N_11762,N_11325);
nor U12706 (N_12706,N_11663,N_11287);
nor U12707 (N_12707,N_11277,N_11514);
nor U12708 (N_12708,N_11267,N_11483);
nand U12709 (N_12709,N_11218,N_11914);
nand U12710 (N_12710,N_11855,N_11434);
or U12711 (N_12711,N_11460,N_11827);
nor U12712 (N_12712,N_11765,N_11311);
or U12713 (N_12713,N_11419,N_11940);
and U12714 (N_12714,N_11366,N_11378);
or U12715 (N_12715,N_11221,N_11257);
and U12716 (N_12716,N_11932,N_11997);
nand U12717 (N_12717,N_11888,N_11979);
xor U12718 (N_12718,N_11258,N_11624);
and U12719 (N_12719,N_11791,N_11508);
nand U12720 (N_12720,N_11765,N_11263);
nor U12721 (N_12721,N_11913,N_11712);
nand U12722 (N_12722,N_11923,N_11547);
nand U12723 (N_12723,N_11239,N_11848);
xnor U12724 (N_12724,N_11668,N_11385);
nand U12725 (N_12725,N_11656,N_11922);
or U12726 (N_12726,N_11708,N_11557);
nand U12727 (N_12727,N_11665,N_11740);
xnor U12728 (N_12728,N_11235,N_11307);
and U12729 (N_12729,N_11674,N_11243);
nor U12730 (N_12730,N_11641,N_11930);
or U12731 (N_12731,N_11241,N_11828);
or U12732 (N_12732,N_11592,N_11224);
and U12733 (N_12733,N_11214,N_11548);
and U12734 (N_12734,N_11926,N_11214);
xnor U12735 (N_12735,N_11576,N_11460);
nand U12736 (N_12736,N_11447,N_11422);
xnor U12737 (N_12737,N_11608,N_11854);
xnor U12738 (N_12738,N_11260,N_11616);
or U12739 (N_12739,N_11766,N_11455);
or U12740 (N_12740,N_11559,N_11895);
and U12741 (N_12741,N_11960,N_11910);
or U12742 (N_12742,N_11435,N_11657);
and U12743 (N_12743,N_11340,N_11607);
xor U12744 (N_12744,N_11473,N_11907);
nand U12745 (N_12745,N_11706,N_11685);
and U12746 (N_12746,N_11345,N_11495);
or U12747 (N_12747,N_11449,N_11653);
and U12748 (N_12748,N_11622,N_11852);
or U12749 (N_12749,N_11544,N_11938);
nand U12750 (N_12750,N_11865,N_11861);
or U12751 (N_12751,N_11439,N_11266);
nor U12752 (N_12752,N_11840,N_11377);
or U12753 (N_12753,N_11475,N_11443);
nor U12754 (N_12754,N_11467,N_11649);
or U12755 (N_12755,N_11593,N_11714);
xnor U12756 (N_12756,N_11771,N_11920);
xor U12757 (N_12757,N_11897,N_11895);
and U12758 (N_12758,N_11399,N_11829);
or U12759 (N_12759,N_11288,N_11419);
and U12760 (N_12760,N_11513,N_11874);
and U12761 (N_12761,N_11930,N_11387);
nand U12762 (N_12762,N_11205,N_11747);
or U12763 (N_12763,N_11874,N_11714);
nor U12764 (N_12764,N_11266,N_11897);
xor U12765 (N_12765,N_11557,N_11464);
and U12766 (N_12766,N_11682,N_11547);
or U12767 (N_12767,N_11503,N_11252);
nor U12768 (N_12768,N_11531,N_11922);
and U12769 (N_12769,N_11526,N_11308);
nand U12770 (N_12770,N_11964,N_11821);
nor U12771 (N_12771,N_11704,N_11969);
nor U12772 (N_12772,N_11782,N_11633);
nand U12773 (N_12773,N_11600,N_11809);
xnor U12774 (N_12774,N_11668,N_11615);
and U12775 (N_12775,N_11874,N_11660);
nand U12776 (N_12776,N_11745,N_11467);
xnor U12777 (N_12777,N_11786,N_11486);
nor U12778 (N_12778,N_11362,N_11833);
or U12779 (N_12779,N_11547,N_11702);
and U12780 (N_12780,N_11905,N_11369);
nand U12781 (N_12781,N_11777,N_11708);
xnor U12782 (N_12782,N_11511,N_11638);
and U12783 (N_12783,N_11682,N_11715);
or U12784 (N_12784,N_11265,N_11385);
xor U12785 (N_12785,N_11694,N_11359);
or U12786 (N_12786,N_11482,N_11869);
nand U12787 (N_12787,N_11969,N_11621);
nor U12788 (N_12788,N_11683,N_11476);
xnor U12789 (N_12789,N_11251,N_11435);
xnor U12790 (N_12790,N_11350,N_11922);
and U12791 (N_12791,N_11641,N_11406);
nand U12792 (N_12792,N_11510,N_11866);
xnor U12793 (N_12793,N_11235,N_11747);
or U12794 (N_12794,N_11460,N_11701);
nand U12795 (N_12795,N_11895,N_11367);
or U12796 (N_12796,N_11368,N_11230);
nor U12797 (N_12797,N_11319,N_11490);
and U12798 (N_12798,N_11661,N_11864);
xor U12799 (N_12799,N_11775,N_11655);
or U12800 (N_12800,N_12167,N_12751);
nand U12801 (N_12801,N_12672,N_12064);
nor U12802 (N_12802,N_12021,N_12380);
xnor U12803 (N_12803,N_12409,N_12391);
and U12804 (N_12804,N_12622,N_12442);
nor U12805 (N_12805,N_12209,N_12315);
and U12806 (N_12806,N_12038,N_12191);
and U12807 (N_12807,N_12311,N_12240);
xnor U12808 (N_12808,N_12454,N_12121);
nand U12809 (N_12809,N_12224,N_12572);
nand U12810 (N_12810,N_12732,N_12793);
or U12811 (N_12811,N_12693,N_12140);
or U12812 (N_12812,N_12117,N_12290);
or U12813 (N_12813,N_12686,N_12418);
and U12814 (N_12814,N_12199,N_12758);
xor U12815 (N_12815,N_12004,N_12695);
and U12816 (N_12816,N_12359,N_12300);
and U12817 (N_12817,N_12464,N_12610);
xor U12818 (N_12818,N_12178,N_12669);
xnor U12819 (N_12819,N_12502,N_12343);
nand U12820 (N_12820,N_12061,N_12003);
nor U12821 (N_12821,N_12386,N_12242);
nor U12822 (N_12822,N_12376,N_12094);
nand U12823 (N_12823,N_12198,N_12461);
nand U12824 (N_12824,N_12707,N_12645);
and U12825 (N_12825,N_12155,N_12377);
nand U12826 (N_12826,N_12573,N_12568);
and U12827 (N_12827,N_12763,N_12655);
nand U12828 (N_12828,N_12593,N_12028);
and U12829 (N_12829,N_12467,N_12187);
xnor U12830 (N_12830,N_12206,N_12030);
nand U12831 (N_12831,N_12599,N_12284);
nand U12832 (N_12832,N_12754,N_12741);
nor U12833 (N_12833,N_12726,N_12671);
or U12834 (N_12834,N_12656,N_12071);
nand U12835 (N_12835,N_12319,N_12534);
and U12836 (N_12836,N_12116,N_12542);
xor U12837 (N_12837,N_12344,N_12350);
or U12838 (N_12838,N_12156,N_12349);
xnor U12839 (N_12839,N_12182,N_12595);
nand U12840 (N_12840,N_12031,N_12288);
nor U12841 (N_12841,N_12781,N_12479);
xnor U12842 (N_12842,N_12445,N_12483);
and U12843 (N_12843,N_12468,N_12474);
nor U12844 (N_12844,N_12045,N_12497);
nor U12845 (N_12845,N_12421,N_12279);
xor U12846 (N_12846,N_12135,N_12118);
nor U12847 (N_12847,N_12389,N_12145);
and U12848 (N_12848,N_12422,N_12587);
nor U12849 (N_12849,N_12576,N_12473);
or U12850 (N_12850,N_12225,N_12407);
xor U12851 (N_12851,N_12719,N_12362);
nor U12852 (N_12852,N_12077,N_12446);
or U12853 (N_12853,N_12276,N_12498);
or U12854 (N_12854,N_12103,N_12297);
xnor U12855 (N_12855,N_12333,N_12492);
nor U12856 (N_12856,N_12705,N_12411);
and U12857 (N_12857,N_12125,N_12318);
xor U12858 (N_12858,N_12133,N_12605);
and U12859 (N_12859,N_12752,N_12480);
xor U12860 (N_12860,N_12087,N_12110);
nor U12861 (N_12861,N_12513,N_12641);
xnor U12862 (N_12862,N_12316,N_12678);
nand U12863 (N_12863,N_12403,N_12281);
nand U12864 (N_12864,N_12716,N_12334);
xor U12865 (N_12865,N_12217,N_12257);
nor U12866 (N_12866,N_12553,N_12165);
and U12867 (N_12867,N_12580,N_12337);
nand U12868 (N_12868,N_12010,N_12541);
or U12869 (N_12869,N_12684,N_12197);
nor U12870 (N_12870,N_12037,N_12516);
and U12871 (N_12871,N_12168,N_12345);
xor U12872 (N_12872,N_12356,N_12489);
and U12873 (N_12873,N_12395,N_12501);
nand U12874 (N_12874,N_12272,N_12091);
or U12875 (N_12875,N_12636,N_12425);
and U12876 (N_12876,N_12269,N_12238);
nor U12877 (N_12877,N_12302,N_12792);
nor U12878 (N_12878,N_12736,N_12679);
nor U12879 (N_12879,N_12075,N_12002);
or U12880 (N_12880,N_12093,N_12755);
nor U12881 (N_12881,N_12008,N_12438);
nor U12882 (N_12882,N_12363,N_12079);
and U12883 (N_12883,N_12136,N_12430);
or U12884 (N_12884,N_12029,N_12256);
nor U12885 (N_12885,N_12107,N_12760);
nand U12886 (N_12886,N_12289,N_12729);
nor U12887 (N_12887,N_12383,N_12397);
and U12888 (N_12888,N_12073,N_12556);
xor U12889 (N_12889,N_12128,N_12049);
xnor U12890 (N_12890,N_12585,N_12432);
nor U12891 (N_12891,N_12779,N_12042);
or U12892 (N_12892,N_12699,N_12047);
xnor U12893 (N_12893,N_12723,N_12046);
nor U12894 (N_12894,N_12494,N_12646);
nand U12895 (N_12895,N_12650,N_12561);
or U12896 (N_12896,N_12774,N_12465);
or U12897 (N_12897,N_12661,N_12538);
nand U12898 (N_12898,N_12666,N_12552);
xor U12899 (N_12899,N_12180,N_12353);
and U12900 (N_12900,N_12720,N_12569);
xnor U12901 (N_12901,N_12050,N_12083);
xor U12902 (N_12902,N_12499,N_12357);
nor U12903 (N_12903,N_12546,N_12390);
or U12904 (N_12904,N_12163,N_12727);
xor U12905 (N_12905,N_12371,N_12581);
nor U12906 (N_12906,N_12239,N_12067);
and U12907 (N_12907,N_12006,N_12560);
nand U12908 (N_12908,N_12697,N_12711);
xor U12909 (N_12909,N_12055,N_12575);
nand U12910 (N_12910,N_12651,N_12273);
xnor U12911 (N_12911,N_12172,N_12314);
or U12912 (N_12912,N_12586,N_12439);
and U12913 (N_12913,N_12462,N_12161);
nor U12914 (N_12914,N_12746,N_12564);
nor U12915 (N_12915,N_12119,N_12310);
xor U12916 (N_12916,N_12470,N_12336);
nand U12917 (N_12917,N_12266,N_12623);
nor U12918 (N_12918,N_12547,N_12068);
nand U12919 (N_12919,N_12122,N_12387);
xor U12920 (N_12920,N_12780,N_12227);
or U12921 (N_12921,N_12435,N_12277);
nor U12922 (N_12922,N_12275,N_12372);
and U12923 (N_12923,N_12398,N_12216);
or U12924 (N_12924,N_12451,N_12293);
or U12925 (N_12925,N_12081,N_12120);
or U12926 (N_12926,N_12582,N_12591);
nand U12927 (N_12927,N_12151,N_12642);
or U12928 (N_12928,N_12696,N_12260);
and U12929 (N_12929,N_12771,N_12740);
nor U12930 (N_12930,N_12253,N_12708);
and U12931 (N_12931,N_12097,N_12459);
nand U12932 (N_12932,N_12562,N_12417);
nand U12933 (N_12933,N_12134,N_12698);
nand U12934 (N_12934,N_12322,N_12000);
nand U12935 (N_12935,N_12453,N_12132);
nand U12936 (N_12936,N_12258,N_12660);
nor U12937 (N_12937,N_12434,N_12521);
xor U12938 (N_12938,N_12169,N_12080);
or U12939 (N_12939,N_12309,N_12001);
or U12940 (N_12940,N_12412,N_12348);
nor U12941 (N_12941,N_12193,N_12691);
or U12942 (N_12942,N_12195,N_12179);
nor U12943 (N_12943,N_12761,N_12447);
xnor U12944 (N_12944,N_12009,N_12394);
nor U12945 (N_12945,N_12787,N_12016);
nand U12946 (N_12946,N_12431,N_12059);
or U12947 (N_12947,N_12041,N_12065);
nor U12948 (N_12948,N_12665,N_12221);
nand U12949 (N_12949,N_12485,N_12278);
nor U12950 (N_12950,N_12742,N_12101);
nor U12951 (N_12951,N_12084,N_12505);
nor U12952 (N_12952,N_12054,N_12332);
xor U12953 (N_12953,N_12782,N_12476);
and U12954 (N_12954,N_12381,N_12682);
xor U12955 (N_12955,N_12635,N_12177);
nor U12956 (N_12956,N_12096,N_12413);
nand U12957 (N_12957,N_12706,N_12689);
and U12958 (N_12958,N_12373,N_12737);
nor U12959 (N_12959,N_12340,N_12063);
xnor U12960 (N_12960,N_12647,N_12150);
nand U12961 (N_12961,N_12159,N_12231);
or U12962 (N_12962,N_12228,N_12072);
and U12963 (N_12963,N_12274,N_12173);
or U12964 (N_12964,N_12486,N_12088);
nand U12965 (N_12965,N_12361,N_12767);
nand U12966 (N_12966,N_12060,N_12419);
and U12967 (N_12967,N_12620,N_12488);
xnor U12968 (N_12968,N_12222,N_12306);
nor U12969 (N_12969,N_12251,N_12549);
or U12970 (N_12970,N_12694,N_12082);
or U12971 (N_12971,N_12219,N_12607);
and U12972 (N_12972,N_12496,N_12113);
nor U12973 (N_12973,N_12612,N_12157);
and U12974 (N_12974,N_12189,N_12052);
nand U12975 (N_12975,N_12237,N_12011);
or U12976 (N_12976,N_12681,N_12370);
or U12977 (N_12977,N_12617,N_12713);
xor U12978 (N_12978,N_12778,N_12158);
and U12979 (N_12979,N_12654,N_12589);
and U12980 (N_12980,N_12621,N_12313);
nand U12981 (N_12981,N_12263,N_12368);
nand U12982 (N_12982,N_12772,N_12517);
or U12983 (N_12983,N_12229,N_12023);
nand U12984 (N_12984,N_12035,N_12588);
nand U12985 (N_12985,N_12559,N_12185);
and U12986 (N_12986,N_12700,N_12244);
xnor U12987 (N_12987,N_12724,N_12043);
xnor U12988 (N_12988,N_12111,N_12558);
nor U12989 (N_12989,N_12626,N_12282);
and U12990 (N_12990,N_12215,N_12034);
and U12991 (N_12991,N_12085,N_12175);
nor U12992 (N_12992,N_12500,N_12481);
nand U12993 (N_12993,N_12143,N_12785);
nor U12994 (N_12994,N_12335,N_12731);
and U12995 (N_12995,N_12428,N_12652);
and U12996 (N_12996,N_12640,N_12196);
xnor U12997 (N_12997,N_12563,N_12644);
nand U12998 (N_12998,N_12127,N_12139);
nand U12999 (N_12999,N_12526,N_12099);
nand U13000 (N_13000,N_12149,N_12443);
xor U13001 (N_13001,N_12183,N_12205);
nor U13002 (N_13002,N_12355,N_12347);
or U13003 (N_13003,N_12303,N_12797);
nor U13004 (N_13004,N_12305,N_12466);
or U13005 (N_13005,N_12298,N_12188);
nand U13006 (N_13006,N_12414,N_12643);
nor U13007 (N_13007,N_12058,N_12070);
nand U13008 (N_13008,N_12570,N_12789);
nor U13009 (N_13009,N_12773,N_12078);
xor U13010 (N_13010,N_12507,N_12676);
or U13011 (N_13011,N_12744,N_12769);
xor U13012 (N_13012,N_12100,N_12735);
nand U13013 (N_13013,N_12426,N_12074);
or U13014 (N_13014,N_12602,N_12066);
or U13015 (N_13015,N_12448,N_12252);
and U13016 (N_13016,N_12743,N_12250);
or U13017 (N_13017,N_12039,N_12776);
nand U13018 (N_13018,N_12463,N_12543);
nand U13019 (N_13019,N_12709,N_12608);
xor U13020 (N_13020,N_12606,N_12765);
or U13021 (N_13021,N_12579,N_12365);
xnor U13022 (N_13022,N_12076,N_12628);
xor U13023 (N_13023,N_12262,N_12089);
nor U13024 (N_13024,N_12753,N_12631);
nor U13025 (N_13025,N_12270,N_12604);
or U13026 (N_13026,N_12423,N_12280);
and U13027 (N_13027,N_12317,N_12565);
or U13028 (N_13028,N_12057,N_12324);
nand U13029 (N_13029,N_12086,N_12092);
nor U13030 (N_13030,N_12249,N_12733);
nor U13031 (N_13031,N_12566,N_12663);
nand U13032 (N_13032,N_12677,N_12012);
or U13033 (N_13033,N_12603,N_12528);
nor U13034 (N_13034,N_12590,N_12594);
xnor U13035 (N_13035,N_12685,N_12524);
and U13036 (N_13036,N_12509,N_12638);
or U13037 (N_13037,N_12675,N_12584);
and U13038 (N_13038,N_12471,N_12768);
nor U13039 (N_13039,N_12154,N_12291);
or U13040 (N_13040,N_12162,N_12657);
nor U13041 (N_13041,N_12166,N_12379);
or U13042 (N_13042,N_12477,N_12688);
and U13043 (N_13043,N_12235,N_12775);
xor U13044 (N_13044,N_12374,N_12105);
xnor U13045 (N_13045,N_12420,N_12181);
and U13046 (N_13046,N_12633,N_12255);
nand U13047 (N_13047,N_12044,N_12056);
and U13048 (N_13048,N_12523,N_12106);
xor U13049 (N_13049,N_12331,N_12687);
nand U13050 (N_13050,N_12456,N_12514);
nand U13051 (N_13051,N_12321,N_12346);
xnor U13052 (N_13052,N_12354,N_12721);
xnor U13053 (N_13053,N_12051,N_12416);
or U13054 (N_13054,N_12510,N_12295);
xor U13055 (N_13055,N_12794,N_12616);
and U13056 (N_13056,N_12529,N_12490);
or U13057 (N_13057,N_12658,N_12259);
xnor U13058 (N_13058,N_12415,N_12102);
nor U13059 (N_13059,N_12153,N_12022);
xor U13060 (N_13060,N_12320,N_12777);
or U13061 (N_13061,N_12265,N_12583);
or U13062 (N_13062,N_12203,N_12323);
or U13063 (N_13063,N_12515,N_12680);
or U13064 (N_13064,N_12147,N_12738);
nor U13065 (N_13065,N_12271,N_12450);
or U13066 (N_13066,N_12632,N_12126);
nand U13067 (N_13067,N_12220,N_12551);
and U13068 (N_13068,N_12718,N_12405);
nor U13069 (N_13069,N_12614,N_12301);
nand U13070 (N_13070,N_12670,N_12458);
xnor U13071 (N_13071,N_12567,N_12018);
nand U13072 (N_13072,N_12449,N_12730);
xor U13073 (N_13073,N_12378,N_12327);
xnor U13074 (N_13074,N_12784,N_12596);
nor U13075 (N_13075,N_12637,N_12764);
nand U13076 (N_13076,N_12712,N_12750);
xor U13077 (N_13077,N_12098,N_12062);
and U13078 (N_13078,N_12184,N_12200);
nor U13079 (N_13079,N_12226,N_12460);
nand U13080 (N_13080,N_12659,N_12747);
nor U13081 (N_13081,N_12557,N_12032);
or U13082 (N_13082,N_12299,N_12401);
nand U13083 (N_13083,N_12766,N_12429);
nand U13084 (N_13084,N_12358,N_12330);
nor U13085 (N_13085,N_12452,N_12164);
or U13086 (N_13086,N_12017,N_12007);
xor U13087 (N_13087,N_12053,N_12577);
or U13088 (N_13088,N_12487,N_12475);
and U13089 (N_13089,N_12624,N_12539);
nand U13090 (N_13090,N_12396,N_12540);
nand U13091 (N_13091,N_12749,N_12005);
nor U13092 (N_13092,N_12146,N_12506);
nand U13093 (N_13093,N_12796,N_12325);
xnor U13094 (N_13094,N_12307,N_12283);
xor U13095 (N_13095,N_12095,N_12601);
nand U13096 (N_13096,N_12410,N_12437);
nor U13097 (N_13097,N_12522,N_12385);
xor U13098 (N_13098,N_12790,N_12619);
xor U13099 (N_13099,N_12609,N_12491);
or U13100 (N_13100,N_12234,N_12537);
nand U13101 (N_13101,N_12109,N_12717);
nand U13102 (N_13102,N_12527,N_12545);
xnor U13103 (N_13103,N_12544,N_12673);
xnor U13104 (N_13104,N_12639,N_12662);
or U13105 (N_13105,N_12791,N_12069);
or U13106 (N_13106,N_12114,N_12267);
nand U13107 (N_13107,N_12408,N_12015);
or U13108 (N_13108,N_12495,N_12611);
or U13109 (N_13109,N_12457,N_12788);
xnor U13110 (N_13110,N_12201,N_12090);
nor U13111 (N_13111,N_12615,N_12144);
xor U13112 (N_13112,N_12033,N_12048);
xnor U13113 (N_13113,N_12366,N_12247);
and U13114 (N_13114,N_12027,N_12484);
and U13115 (N_13115,N_12194,N_12482);
xnor U13116 (N_13116,N_12399,N_12285);
nand U13117 (N_13117,N_12124,N_12504);
xnor U13118 (N_13118,N_12600,N_12795);
or U13119 (N_13119,N_12375,N_12756);
nand U13120 (N_13120,N_12233,N_12328);
or U13121 (N_13121,N_12243,N_12798);
xor U13122 (N_13122,N_12341,N_12629);
or U13123 (N_13123,N_12714,N_12384);
and U13124 (N_13124,N_12026,N_12400);
nand U13125 (N_13125,N_12236,N_12261);
or U13126 (N_13126,N_12190,N_12648);
or U13127 (N_13127,N_12036,N_12212);
xor U13128 (N_13128,N_12170,N_12393);
nand U13129 (N_13129,N_12440,N_12748);
nand U13130 (N_13130,N_12555,N_12627);
and U13131 (N_13131,N_12531,N_12208);
nor U13132 (N_13132,N_12352,N_12722);
xor U13133 (N_13133,N_12533,N_12503);
and U13134 (N_13134,N_12786,N_12264);
nand U13135 (N_13135,N_12137,N_12254);
and U13136 (N_13136,N_12578,N_12223);
or U13137 (N_13137,N_12020,N_12342);
nor U13138 (N_13138,N_12339,N_12759);
and U13139 (N_13139,N_12211,N_12186);
or U13140 (N_13140,N_12799,N_12668);
and U13141 (N_13141,N_12367,N_12734);
nor U13142 (N_13142,N_12701,N_12702);
nand U13143 (N_13143,N_12019,N_12388);
nor U13144 (N_13144,N_12634,N_12192);
or U13145 (N_13145,N_12683,N_12427);
and U13146 (N_13146,N_12308,N_12338);
and U13147 (N_13147,N_12597,N_12204);
or U13148 (N_13148,N_12245,N_12214);
or U13149 (N_13149,N_12292,N_12613);
or U13150 (N_13150,N_12441,N_12382);
or U13151 (N_13151,N_12014,N_12739);
or U13152 (N_13152,N_12770,N_12294);
and U13153 (N_13153,N_12530,N_12728);
nand U13154 (N_13154,N_12013,N_12493);
nand U13155 (N_13155,N_12690,N_12574);
nand U13156 (N_13156,N_12433,N_12112);
nor U13157 (N_13157,N_12108,N_12207);
xnor U13158 (N_13158,N_12511,N_12406);
or U13159 (N_13159,N_12703,N_12674);
nor U13160 (N_13160,N_12592,N_12286);
and U13161 (N_13161,N_12248,N_12757);
and U13162 (N_13162,N_12625,N_12618);
nand U13163 (N_13163,N_12329,N_12160);
nor U13164 (N_13164,N_12554,N_12131);
and U13165 (N_13165,N_12304,N_12478);
or U13166 (N_13166,N_12025,N_12123);
nor U13167 (N_13167,N_12202,N_12142);
and U13168 (N_13168,N_12218,N_12246);
nor U13169 (N_13169,N_12762,N_12436);
and U13170 (N_13170,N_12519,N_12518);
nand U13171 (N_13171,N_12402,N_12630);
nor U13172 (N_13172,N_12404,N_12536);
nand U13173 (N_13173,N_12171,N_12312);
or U13174 (N_13174,N_12369,N_12213);
nor U13175 (N_13175,N_12745,N_12525);
and U13176 (N_13176,N_12148,N_12715);
nand U13177 (N_13177,N_12520,N_12653);
nand U13178 (N_13178,N_12455,N_12667);
or U13179 (N_13179,N_12141,N_12364);
and U13180 (N_13180,N_12472,N_12210);
or U13181 (N_13181,N_12692,N_12268);
and U13182 (N_13182,N_12174,N_12444);
nor U13183 (N_13183,N_12598,N_12571);
nor U13184 (N_13184,N_12649,N_12710);
xnor U13185 (N_13185,N_12138,N_12351);
or U13186 (N_13186,N_12783,N_12424);
and U13187 (N_13187,N_12232,N_12152);
xnor U13188 (N_13188,N_12550,N_12241);
nor U13189 (N_13189,N_12725,N_12326);
or U13190 (N_13190,N_12287,N_12296);
and U13191 (N_13191,N_12392,N_12115);
or U13192 (N_13192,N_12230,N_12548);
nand U13193 (N_13193,N_12176,N_12535);
nand U13194 (N_13194,N_12024,N_12532);
nand U13195 (N_13195,N_12130,N_12360);
nand U13196 (N_13196,N_12469,N_12129);
or U13197 (N_13197,N_12704,N_12508);
nor U13198 (N_13198,N_12040,N_12512);
nand U13199 (N_13199,N_12664,N_12104);
xor U13200 (N_13200,N_12113,N_12686);
nand U13201 (N_13201,N_12530,N_12694);
and U13202 (N_13202,N_12616,N_12005);
nor U13203 (N_13203,N_12195,N_12706);
nor U13204 (N_13204,N_12697,N_12700);
nand U13205 (N_13205,N_12323,N_12078);
nor U13206 (N_13206,N_12446,N_12253);
or U13207 (N_13207,N_12389,N_12277);
nand U13208 (N_13208,N_12424,N_12699);
xnor U13209 (N_13209,N_12361,N_12483);
and U13210 (N_13210,N_12372,N_12386);
nor U13211 (N_13211,N_12581,N_12788);
nor U13212 (N_13212,N_12204,N_12642);
or U13213 (N_13213,N_12411,N_12140);
or U13214 (N_13214,N_12096,N_12301);
nand U13215 (N_13215,N_12053,N_12737);
or U13216 (N_13216,N_12315,N_12414);
xor U13217 (N_13217,N_12088,N_12771);
or U13218 (N_13218,N_12198,N_12650);
or U13219 (N_13219,N_12255,N_12253);
and U13220 (N_13220,N_12721,N_12597);
nor U13221 (N_13221,N_12295,N_12266);
or U13222 (N_13222,N_12145,N_12797);
nor U13223 (N_13223,N_12216,N_12266);
or U13224 (N_13224,N_12491,N_12467);
or U13225 (N_13225,N_12038,N_12301);
nand U13226 (N_13226,N_12416,N_12717);
or U13227 (N_13227,N_12736,N_12627);
xor U13228 (N_13228,N_12014,N_12797);
nor U13229 (N_13229,N_12114,N_12149);
xnor U13230 (N_13230,N_12766,N_12555);
xor U13231 (N_13231,N_12078,N_12173);
nor U13232 (N_13232,N_12195,N_12474);
and U13233 (N_13233,N_12608,N_12793);
nand U13234 (N_13234,N_12155,N_12684);
and U13235 (N_13235,N_12217,N_12128);
xor U13236 (N_13236,N_12335,N_12251);
or U13237 (N_13237,N_12213,N_12160);
or U13238 (N_13238,N_12644,N_12193);
and U13239 (N_13239,N_12256,N_12631);
nand U13240 (N_13240,N_12592,N_12477);
nor U13241 (N_13241,N_12521,N_12770);
or U13242 (N_13242,N_12286,N_12314);
or U13243 (N_13243,N_12507,N_12481);
nor U13244 (N_13244,N_12127,N_12284);
nand U13245 (N_13245,N_12765,N_12382);
nor U13246 (N_13246,N_12529,N_12112);
nand U13247 (N_13247,N_12429,N_12606);
and U13248 (N_13248,N_12235,N_12275);
and U13249 (N_13249,N_12097,N_12160);
xor U13250 (N_13250,N_12165,N_12458);
and U13251 (N_13251,N_12185,N_12737);
xor U13252 (N_13252,N_12452,N_12654);
xor U13253 (N_13253,N_12526,N_12367);
or U13254 (N_13254,N_12753,N_12273);
nor U13255 (N_13255,N_12228,N_12617);
nor U13256 (N_13256,N_12320,N_12044);
nor U13257 (N_13257,N_12444,N_12056);
xnor U13258 (N_13258,N_12190,N_12235);
nand U13259 (N_13259,N_12242,N_12660);
xnor U13260 (N_13260,N_12104,N_12548);
nand U13261 (N_13261,N_12662,N_12047);
and U13262 (N_13262,N_12015,N_12265);
nor U13263 (N_13263,N_12053,N_12424);
nand U13264 (N_13264,N_12172,N_12305);
nor U13265 (N_13265,N_12292,N_12757);
nand U13266 (N_13266,N_12485,N_12286);
and U13267 (N_13267,N_12430,N_12015);
xnor U13268 (N_13268,N_12105,N_12575);
nor U13269 (N_13269,N_12737,N_12076);
xor U13270 (N_13270,N_12009,N_12727);
nor U13271 (N_13271,N_12590,N_12306);
and U13272 (N_13272,N_12596,N_12074);
nor U13273 (N_13273,N_12791,N_12763);
nor U13274 (N_13274,N_12045,N_12166);
and U13275 (N_13275,N_12540,N_12157);
nor U13276 (N_13276,N_12354,N_12372);
nor U13277 (N_13277,N_12742,N_12784);
nand U13278 (N_13278,N_12680,N_12306);
or U13279 (N_13279,N_12034,N_12676);
or U13280 (N_13280,N_12517,N_12448);
nand U13281 (N_13281,N_12320,N_12441);
nand U13282 (N_13282,N_12326,N_12749);
xnor U13283 (N_13283,N_12107,N_12218);
nand U13284 (N_13284,N_12737,N_12217);
and U13285 (N_13285,N_12266,N_12102);
and U13286 (N_13286,N_12592,N_12595);
or U13287 (N_13287,N_12407,N_12144);
nor U13288 (N_13288,N_12585,N_12130);
nor U13289 (N_13289,N_12053,N_12052);
or U13290 (N_13290,N_12766,N_12389);
and U13291 (N_13291,N_12397,N_12244);
or U13292 (N_13292,N_12115,N_12142);
nor U13293 (N_13293,N_12377,N_12182);
nand U13294 (N_13294,N_12268,N_12762);
and U13295 (N_13295,N_12235,N_12194);
and U13296 (N_13296,N_12521,N_12758);
xor U13297 (N_13297,N_12737,N_12321);
or U13298 (N_13298,N_12700,N_12192);
and U13299 (N_13299,N_12373,N_12350);
and U13300 (N_13300,N_12038,N_12166);
nor U13301 (N_13301,N_12694,N_12345);
xor U13302 (N_13302,N_12289,N_12659);
nor U13303 (N_13303,N_12217,N_12130);
nor U13304 (N_13304,N_12349,N_12105);
nor U13305 (N_13305,N_12312,N_12685);
and U13306 (N_13306,N_12315,N_12356);
nor U13307 (N_13307,N_12206,N_12627);
and U13308 (N_13308,N_12244,N_12717);
nor U13309 (N_13309,N_12715,N_12378);
nor U13310 (N_13310,N_12156,N_12214);
nand U13311 (N_13311,N_12694,N_12024);
or U13312 (N_13312,N_12104,N_12297);
nand U13313 (N_13313,N_12285,N_12757);
nor U13314 (N_13314,N_12497,N_12554);
and U13315 (N_13315,N_12664,N_12591);
nand U13316 (N_13316,N_12726,N_12054);
or U13317 (N_13317,N_12285,N_12650);
nor U13318 (N_13318,N_12271,N_12444);
or U13319 (N_13319,N_12494,N_12608);
xnor U13320 (N_13320,N_12128,N_12333);
xor U13321 (N_13321,N_12286,N_12419);
or U13322 (N_13322,N_12563,N_12464);
or U13323 (N_13323,N_12793,N_12694);
xor U13324 (N_13324,N_12155,N_12790);
or U13325 (N_13325,N_12437,N_12568);
nand U13326 (N_13326,N_12145,N_12275);
xnor U13327 (N_13327,N_12439,N_12109);
or U13328 (N_13328,N_12713,N_12468);
xor U13329 (N_13329,N_12021,N_12423);
xor U13330 (N_13330,N_12512,N_12264);
nand U13331 (N_13331,N_12747,N_12437);
and U13332 (N_13332,N_12590,N_12516);
and U13333 (N_13333,N_12703,N_12520);
nor U13334 (N_13334,N_12528,N_12111);
and U13335 (N_13335,N_12214,N_12205);
xnor U13336 (N_13336,N_12229,N_12110);
nand U13337 (N_13337,N_12005,N_12029);
xor U13338 (N_13338,N_12183,N_12729);
nor U13339 (N_13339,N_12150,N_12026);
xor U13340 (N_13340,N_12354,N_12256);
nand U13341 (N_13341,N_12567,N_12767);
and U13342 (N_13342,N_12764,N_12575);
nand U13343 (N_13343,N_12137,N_12381);
xor U13344 (N_13344,N_12333,N_12768);
nor U13345 (N_13345,N_12224,N_12009);
and U13346 (N_13346,N_12634,N_12071);
nand U13347 (N_13347,N_12195,N_12019);
and U13348 (N_13348,N_12391,N_12040);
nand U13349 (N_13349,N_12693,N_12601);
xnor U13350 (N_13350,N_12532,N_12262);
nor U13351 (N_13351,N_12639,N_12038);
xnor U13352 (N_13352,N_12672,N_12493);
xor U13353 (N_13353,N_12689,N_12661);
or U13354 (N_13354,N_12447,N_12315);
xor U13355 (N_13355,N_12229,N_12310);
xor U13356 (N_13356,N_12761,N_12082);
nor U13357 (N_13357,N_12564,N_12395);
xor U13358 (N_13358,N_12487,N_12648);
nor U13359 (N_13359,N_12253,N_12672);
nor U13360 (N_13360,N_12646,N_12036);
and U13361 (N_13361,N_12422,N_12309);
xor U13362 (N_13362,N_12418,N_12147);
or U13363 (N_13363,N_12665,N_12039);
and U13364 (N_13364,N_12733,N_12461);
nand U13365 (N_13365,N_12316,N_12177);
nor U13366 (N_13366,N_12023,N_12623);
or U13367 (N_13367,N_12267,N_12363);
or U13368 (N_13368,N_12367,N_12123);
nor U13369 (N_13369,N_12527,N_12290);
and U13370 (N_13370,N_12565,N_12481);
xor U13371 (N_13371,N_12065,N_12383);
nor U13372 (N_13372,N_12392,N_12486);
or U13373 (N_13373,N_12389,N_12069);
or U13374 (N_13374,N_12136,N_12777);
nor U13375 (N_13375,N_12794,N_12630);
or U13376 (N_13376,N_12291,N_12525);
xnor U13377 (N_13377,N_12510,N_12056);
nor U13378 (N_13378,N_12213,N_12139);
and U13379 (N_13379,N_12342,N_12639);
nor U13380 (N_13380,N_12153,N_12019);
nand U13381 (N_13381,N_12283,N_12000);
xnor U13382 (N_13382,N_12213,N_12226);
xor U13383 (N_13383,N_12261,N_12487);
and U13384 (N_13384,N_12580,N_12147);
or U13385 (N_13385,N_12661,N_12026);
or U13386 (N_13386,N_12364,N_12438);
nor U13387 (N_13387,N_12318,N_12612);
or U13388 (N_13388,N_12391,N_12493);
or U13389 (N_13389,N_12715,N_12082);
xnor U13390 (N_13390,N_12566,N_12365);
nand U13391 (N_13391,N_12426,N_12756);
xor U13392 (N_13392,N_12220,N_12638);
xnor U13393 (N_13393,N_12078,N_12633);
xor U13394 (N_13394,N_12150,N_12690);
and U13395 (N_13395,N_12148,N_12079);
and U13396 (N_13396,N_12295,N_12691);
nor U13397 (N_13397,N_12280,N_12729);
nor U13398 (N_13398,N_12047,N_12044);
nor U13399 (N_13399,N_12762,N_12373);
nor U13400 (N_13400,N_12741,N_12329);
nand U13401 (N_13401,N_12423,N_12608);
nor U13402 (N_13402,N_12481,N_12703);
nor U13403 (N_13403,N_12236,N_12045);
nor U13404 (N_13404,N_12586,N_12193);
and U13405 (N_13405,N_12047,N_12032);
and U13406 (N_13406,N_12132,N_12778);
and U13407 (N_13407,N_12381,N_12625);
or U13408 (N_13408,N_12231,N_12574);
xnor U13409 (N_13409,N_12682,N_12121);
or U13410 (N_13410,N_12275,N_12351);
nor U13411 (N_13411,N_12653,N_12192);
and U13412 (N_13412,N_12369,N_12142);
or U13413 (N_13413,N_12361,N_12196);
nand U13414 (N_13414,N_12615,N_12286);
nor U13415 (N_13415,N_12098,N_12743);
or U13416 (N_13416,N_12519,N_12634);
xnor U13417 (N_13417,N_12745,N_12785);
xnor U13418 (N_13418,N_12496,N_12656);
and U13419 (N_13419,N_12229,N_12211);
nand U13420 (N_13420,N_12117,N_12212);
and U13421 (N_13421,N_12127,N_12604);
nand U13422 (N_13422,N_12156,N_12352);
xor U13423 (N_13423,N_12523,N_12799);
nand U13424 (N_13424,N_12748,N_12227);
or U13425 (N_13425,N_12618,N_12426);
nand U13426 (N_13426,N_12571,N_12434);
and U13427 (N_13427,N_12255,N_12424);
or U13428 (N_13428,N_12457,N_12442);
xor U13429 (N_13429,N_12234,N_12566);
xor U13430 (N_13430,N_12195,N_12558);
nor U13431 (N_13431,N_12481,N_12303);
nor U13432 (N_13432,N_12798,N_12356);
nand U13433 (N_13433,N_12021,N_12679);
nor U13434 (N_13434,N_12173,N_12195);
xnor U13435 (N_13435,N_12096,N_12261);
xor U13436 (N_13436,N_12405,N_12654);
or U13437 (N_13437,N_12543,N_12136);
and U13438 (N_13438,N_12399,N_12553);
xnor U13439 (N_13439,N_12285,N_12140);
or U13440 (N_13440,N_12587,N_12163);
nor U13441 (N_13441,N_12135,N_12736);
and U13442 (N_13442,N_12308,N_12647);
nor U13443 (N_13443,N_12483,N_12525);
nand U13444 (N_13444,N_12430,N_12360);
and U13445 (N_13445,N_12508,N_12542);
nor U13446 (N_13446,N_12455,N_12002);
nand U13447 (N_13447,N_12604,N_12765);
or U13448 (N_13448,N_12799,N_12433);
or U13449 (N_13449,N_12388,N_12733);
nand U13450 (N_13450,N_12218,N_12608);
or U13451 (N_13451,N_12200,N_12087);
nand U13452 (N_13452,N_12653,N_12740);
or U13453 (N_13453,N_12430,N_12421);
nor U13454 (N_13454,N_12722,N_12795);
nand U13455 (N_13455,N_12685,N_12310);
or U13456 (N_13456,N_12241,N_12707);
nand U13457 (N_13457,N_12368,N_12179);
xnor U13458 (N_13458,N_12789,N_12004);
nand U13459 (N_13459,N_12766,N_12032);
nor U13460 (N_13460,N_12627,N_12074);
nor U13461 (N_13461,N_12315,N_12070);
and U13462 (N_13462,N_12477,N_12648);
and U13463 (N_13463,N_12590,N_12089);
and U13464 (N_13464,N_12757,N_12483);
xnor U13465 (N_13465,N_12775,N_12267);
nand U13466 (N_13466,N_12703,N_12185);
xnor U13467 (N_13467,N_12633,N_12018);
and U13468 (N_13468,N_12168,N_12423);
or U13469 (N_13469,N_12008,N_12419);
nor U13470 (N_13470,N_12638,N_12737);
and U13471 (N_13471,N_12200,N_12318);
nor U13472 (N_13472,N_12102,N_12141);
nor U13473 (N_13473,N_12674,N_12142);
nor U13474 (N_13474,N_12403,N_12742);
and U13475 (N_13475,N_12749,N_12691);
or U13476 (N_13476,N_12023,N_12248);
xnor U13477 (N_13477,N_12630,N_12736);
xor U13478 (N_13478,N_12254,N_12103);
or U13479 (N_13479,N_12761,N_12371);
and U13480 (N_13480,N_12386,N_12582);
or U13481 (N_13481,N_12229,N_12644);
nor U13482 (N_13482,N_12629,N_12525);
and U13483 (N_13483,N_12772,N_12225);
nor U13484 (N_13484,N_12089,N_12522);
nor U13485 (N_13485,N_12208,N_12445);
nand U13486 (N_13486,N_12721,N_12775);
nand U13487 (N_13487,N_12248,N_12721);
nor U13488 (N_13488,N_12545,N_12662);
xnor U13489 (N_13489,N_12699,N_12364);
nor U13490 (N_13490,N_12445,N_12712);
and U13491 (N_13491,N_12047,N_12245);
nand U13492 (N_13492,N_12762,N_12491);
nand U13493 (N_13493,N_12675,N_12398);
xor U13494 (N_13494,N_12620,N_12411);
or U13495 (N_13495,N_12533,N_12209);
and U13496 (N_13496,N_12483,N_12671);
xor U13497 (N_13497,N_12105,N_12255);
and U13498 (N_13498,N_12750,N_12289);
or U13499 (N_13499,N_12297,N_12371);
nand U13500 (N_13500,N_12319,N_12660);
xnor U13501 (N_13501,N_12430,N_12670);
xor U13502 (N_13502,N_12538,N_12126);
or U13503 (N_13503,N_12133,N_12338);
or U13504 (N_13504,N_12497,N_12047);
nor U13505 (N_13505,N_12153,N_12390);
xor U13506 (N_13506,N_12164,N_12227);
xnor U13507 (N_13507,N_12423,N_12147);
xnor U13508 (N_13508,N_12354,N_12605);
xor U13509 (N_13509,N_12661,N_12336);
xnor U13510 (N_13510,N_12552,N_12056);
xor U13511 (N_13511,N_12363,N_12196);
and U13512 (N_13512,N_12232,N_12671);
or U13513 (N_13513,N_12461,N_12308);
or U13514 (N_13514,N_12570,N_12301);
or U13515 (N_13515,N_12538,N_12339);
and U13516 (N_13516,N_12542,N_12207);
and U13517 (N_13517,N_12176,N_12015);
or U13518 (N_13518,N_12260,N_12693);
nor U13519 (N_13519,N_12490,N_12338);
xnor U13520 (N_13520,N_12205,N_12360);
nor U13521 (N_13521,N_12264,N_12346);
nand U13522 (N_13522,N_12490,N_12564);
xor U13523 (N_13523,N_12772,N_12171);
nor U13524 (N_13524,N_12367,N_12639);
xnor U13525 (N_13525,N_12620,N_12530);
and U13526 (N_13526,N_12410,N_12606);
nand U13527 (N_13527,N_12786,N_12452);
nand U13528 (N_13528,N_12490,N_12547);
or U13529 (N_13529,N_12786,N_12550);
and U13530 (N_13530,N_12345,N_12350);
and U13531 (N_13531,N_12707,N_12490);
nand U13532 (N_13532,N_12586,N_12020);
nand U13533 (N_13533,N_12095,N_12033);
xnor U13534 (N_13534,N_12188,N_12279);
and U13535 (N_13535,N_12548,N_12304);
nand U13536 (N_13536,N_12096,N_12395);
nor U13537 (N_13537,N_12073,N_12395);
or U13538 (N_13538,N_12097,N_12283);
nor U13539 (N_13539,N_12618,N_12725);
or U13540 (N_13540,N_12578,N_12140);
nor U13541 (N_13541,N_12533,N_12177);
nor U13542 (N_13542,N_12053,N_12519);
nand U13543 (N_13543,N_12699,N_12593);
and U13544 (N_13544,N_12436,N_12082);
nand U13545 (N_13545,N_12433,N_12793);
nand U13546 (N_13546,N_12251,N_12455);
xnor U13547 (N_13547,N_12133,N_12714);
or U13548 (N_13548,N_12095,N_12157);
and U13549 (N_13549,N_12097,N_12711);
and U13550 (N_13550,N_12453,N_12022);
nand U13551 (N_13551,N_12785,N_12007);
nand U13552 (N_13552,N_12227,N_12310);
and U13553 (N_13553,N_12571,N_12588);
xor U13554 (N_13554,N_12334,N_12684);
and U13555 (N_13555,N_12247,N_12732);
nor U13556 (N_13556,N_12536,N_12407);
xor U13557 (N_13557,N_12778,N_12731);
xnor U13558 (N_13558,N_12664,N_12773);
nand U13559 (N_13559,N_12052,N_12565);
and U13560 (N_13560,N_12695,N_12011);
xor U13561 (N_13561,N_12571,N_12655);
and U13562 (N_13562,N_12615,N_12350);
xnor U13563 (N_13563,N_12590,N_12725);
and U13564 (N_13564,N_12790,N_12617);
xor U13565 (N_13565,N_12684,N_12729);
and U13566 (N_13566,N_12469,N_12210);
or U13567 (N_13567,N_12489,N_12086);
nand U13568 (N_13568,N_12054,N_12783);
or U13569 (N_13569,N_12760,N_12680);
nand U13570 (N_13570,N_12260,N_12547);
or U13571 (N_13571,N_12754,N_12050);
or U13572 (N_13572,N_12394,N_12574);
and U13573 (N_13573,N_12445,N_12191);
nand U13574 (N_13574,N_12596,N_12039);
nor U13575 (N_13575,N_12478,N_12587);
and U13576 (N_13576,N_12758,N_12156);
and U13577 (N_13577,N_12356,N_12424);
and U13578 (N_13578,N_12637,N_12441);
xor U13579 (N_13579,N_12476,N_12272);
or U13580 (N_13580,N_12170,N_12109);
or U13581 (N_13581,N_12764,N_12309);
nand U13582 (N_13582,N_12642,N_12771);
nor U13583 (N_13583,N_12279,N_12663);
and U13584 (N_13584,N_12504,N_12006);
and U13585 (N_13585,N_12145,N_12556);
nor U13586 (N_13586,N_12534,N_12602);
nor U13587 (N_13587,N_12719,N_12438);
xnor U13588 (N_13588,N_12566,N_12597);
nand U13589 (N_13589,N_12120,N_12389);
or U13590 (N_13590,N_12079,N_12796);
xnor U13591 (N_13591,N_12403,N_12653);
or U13592 (N_13592,N_12090,N_12124);
xnor U13593 (N_13593,N_12635,N_12615);
and U13594 (N_13594,N_12663,N_12518);
nand U13595 (N_13595,N_12488,N_12763);
and U13596 (N_13596,N_12468,N_12113);
xnor U13597 (N_13597,N_12016,N_12326);
nand U13598 (N_13598,N_12027,N_12488);
and U13599 (N_13599,N_12723,N_12215);
xnor U13600 (N_13600,N_13423,N_13305);
nor U13601 (N_13601,N_13297,N_13239);
and U13602 (N_13602,N_13387,N_13151);
xor U13603 (N_13603,N_13446,N_13395);
xnor U13604 (N_13604,N_13296,N_13099);
nor U13605 (N_13605,N_13084,N_12969);
xor U13606 (N_13606,N_13579,N_12868);
and U13607 (N_13607,N_13479,N_13263);
xnor U13608 (N_13608,N_13348,N_13216);
or U13609 (N_13609,N_13254,N_13349);
nor U13610 (N_13610,N_13083,N_13052);
xnor U13611 (N_13611,N_13458,N_13086);
nand U13612 (N_13612,N_12899,N_13065);
xor U13613 (N_13613,N_13313,N_13106);
nand U13614 (N_13614,N_13309,N_13535);
and U13615 (N_13615,N_12984,N_12916);
xnor U13616 (N_13616,N_13453,N_13318);
xor U13617 (N_13617,N_12891,N_12852);
and U13618 (N_13618,N_13521,N_13119);
and U13619 (N_13619,N_13252,N_12802);
and U13620 (N_13620,N_13034,N_12857);
or U13621 (N_13621,N_13271,N_13191);
or U13622 (N_13622,N_12896,N_13493);
or U13623 (N_13623,N_13071,N_13381);
and U13624 (N_13624,N_13392,N_13462);
nor U13625 (N_13625,N_12967,N_13031);
or U13626 (N_13626,N_13418,N_13519);
or U13627 (N_13627,N_12911,N_13574);
nand U13628 (N_13628,N_13227,N_13530);
or U13629 (N_13629,N_13286,N_13072);
xnor U13630 (N_13630,N_13333,N_13238);
xnor U13631 (N_13631,N_13287,N_12838);
xnor U13632 (N_13632,N_13012,N_12813);
xor U13633 (N_13633,N_13487,N_13073);
xor U13634 (N_13634,N_13023,N_13112);
or U13635 (N_13635,N_12867,N_12974);
or U13636 (N_13636,N_13322,N_13139);
or U13637 (N_13637,N_13406,N_12900);
nor U13638 (N_13638,N_13378,N_13143);
or U13639 (N_13639,N_12843,N_13511);
nor U13640 (N_13640,N_13098,N_13324);
xnor U13641 (N_13641,N_12938,N_13100);
and U13642 (N_13642,N_13005,N_12918);
nor U13643 (N_13643,N_13193,N_13020);
xnor U13644 (N_13644,N_13138,N_13498);
or U13645 (N_13645,N_12924,N_12956);
or U13646 (N_13646,N_13189,N_13057);
xnor U13647 (N_13647,N_13430,N_12816);
xnor U13648 (N_13648,N_12839,N_13477);
nor U13649 (N_13649,N_13489,N_13523);
nand U13650 (N_13650,N_13269,N_13327);
nand U13651 (N_13651,N_13343,N_13236);
or U13652 (N_13652,N_13030,N_13561);
nand U13653 (N_13653,N_13356,N_13257);
xor U13654 (N_13654,N_13434,N_13404);
nor U13655 (N_13655,N_13551,N_12921);
or U13656 (N_13656,N_12878,N_13543);
and U13657 (N_13657,N_13441,N_12874);
nor U13658 (N_13658,N_13243,N_13179);
nor U13659 (N_13659,N_13301,N_13024);
nor U13660 (N_13660,N_13347,N_13029);
or U13661 (N_13661,N_13077,N_13525);
xor U13662 (N_13662,N_13063,N_13342);
nand U13663 (N_13663,N_12844,N_12806);
nand U13664 (N_13664,N_13061,N_13330);
nor U13665 (N_13665,N_13450,N_13137);
and U13666 (N_13666,N_13562,N_13145);
nor U13667 (N_13667,N_13515,N_12992);
nand U13668 (N_13668,N_13282,N_12825);
nand U13669 (N_13669,N_13147,N_13377);
or U13670 (N_13670,N_13375,N_13398);
xnor U13671 (N_13671,N_13074,N_13520);
xnor U13672 (N_13672,N_13497,N_12875);
or U13673 (N_13673,N_13428,N_12932);
nand U13674 (N_13674,N_13117,N_13113);
nor U13675 (N_13675,N_12883,N_12829);
and U13676 (N_13676,N_13533,N_13021);
nor U13677 (N_13677,N_13186,N_12827);
or U13678 (N_13678,N_13044,N_13482);
and U13679 (N_13679,N_12846,N_13415);
or U13680 (N_13680,N_13213,N_13274);
or U13681 (N_13681,N_12803,N_13541);
or U13682 (N_13682,N_13228,N_13038);
xor U13683 (N_13683,N_12948,N_13501);
and U13684 (N_13684,N_13226,N_13165);
nor U13685 (N_13685,N_12823,N_13502);
and U13686 (N_13686,N_13068,N_13224);
or U13687 (N_13687,N_13455,N_12837);
and U13688 (N_13688,N_13383,N_13091);
or U13689 (N_13689,N_12975,N_13545);
nand U13690 (N_13690,N_13401,N_13568);
nor U13691 (N_13691,N_13303,N_12941);
xnor U13692 (N_13692,N_12970,N_12851);
xor U13693 (N_13693,N_13316,N_13153);
and U13694 (N_13694,N_12863,N_12981);
xor U13695 (N_13695,N_12929,N_13565);
xnor U13696 (N_13696,N_12993,N_13027);
and U13697 (N_13697,N_13474,N_13460);
or U13698 (N_13698,N_13516,N_13312);
and U13699 (N_13699,N_13352,N_13293);
nand U13700 (N_13700,N_13412,N_13555);
or U13701 (N_13701,N_13473,N_12988);
xnor U13702 (N_13702,N_12814,N_12977);
nand U13703 (N_13703,N_13573,N_13341);
nor U13704 (N_13704,N_13419,N_12930);
nor U13705 (N_13705,N_13242,N_13304);
nand U13706 (N_13706,N_13110,N_12926);
xnor U13707 (N_13707,N_13513,N_13247);
nand U13708 (N_13708,N_13484,N_13537);
xnor U13709 (N_13709,N_12840,N_12935);
nor U13710 (N_13710,N_13060,N_13577);
nand U13711 (N_13711,N_13488,N_13081);
nand U13712 (N_13712,N_12925,N_13408);
or U13713 (N_13713,N_13386,N_13433);
and U13714 (N_13714,N_13184,N_13399);
or U13715 (N_13715,N_13294,N_13298);
and U13716 (N_13716,N_13361,N_13288);
nor U13717 (N_13717,N_12898,N_13559);
or U13718 (N_13718,N_13556,N_13111);
nand U13719 (N_13719,N_13045,N_12858);
xnor U13720 (N_13720,N_13411,N_13366);
and U13721 (N_13721,N_13456,N_13041);
and U13722 (N_13722,N_13178,N_13241);
nand U13723 (N_13723,N_13563,N_13200);
and U13724 (N_13724,N_13037,N_13215);
xnor U13725 (N_13725,N_13177,N_13156);
nor U13726 (N_13726,N_12862,N_13325);
xnor U13727 (N_13727,N_13445,N_13276);
xnor U13728 (N_13728,N_13373,N_13194);
nand U13729 (N_13729,N_13529,N_13431);
and U13730 (N_13730,N_12937,N_13008);
or U13731 (N_13731,N_13010,N_13451);
xor U13732 (N_13732,N_13315,N_13203);
or U13733 (N_13733,N_13549,N_13397);
nand U13734 (N_13734,N_13201,N_13187);
xor U13735 (N_13735,N_13101,N_13050);
nand U13736 (N_13736,N_13550,N_13332);
nor U13737 (N_13737,N_13589,N_13232);
xnor U13738 (N_13738,N_13481,N_13266);
and U13739 (N_13739,N_13598,N_12927);
xnor U13740 (N_13740,N_12964,N_13095);
nor U13741 (N_13741,N_13066,N_13087);
and U13742 (N_13742,N_13019,N_13259);
and U13743 (N_13743,N_13326,N_13166);
nand U13744 (N_13744,N_13486,N_13440);
or U13745 (N_13745,N_12884,N_13311);
nor U13746 (N_13746,N_13018,N_12903);
or U13747 (N_13747,N_13043,N_12809);
nand U13748 (N_13748,N_13130,N_13494);
and U13749 (N_13749,N_13026,N_13094);
xor U13750 (N_13750,N_13234,N_13245);
or U13751 (N_13751,N_13306,N_13290);
nand U13752 (N_13752,N_13314,N_13135);
and U13753 (N_13753,N_13133,N_12800);
and U13754 (N_13754,N_13268,N_13011);
xnor U13755 (N_13755,N_13233,N_12866);
nand U13756 (N_13756,N_13466,N_13105);
or U13757 (N_13757,N_13576,N_13134);
or U13758 (N_13758,N_13062,N_13379);
or U13759 (N_13759,N_12973,N_12949);
nand U13760 (N_13760,N_13438,N_13572);
or U13761 (N_13761,N_12853,N_13207);
and U13762 (N_13762,N_13424,N_13526);
xor U13763 (N_13763,N_13210,N_12987);
and U13764 (N_13764,N_13032,N_13118);
nand U13765 (N_13765,N_13492,N_12872);
or U13766 (N_13766,N_12950,N_13040);
or U13767 (N_13767,N_12805,N_13067);
nor U13768 (N_13768,N_13417,N_12980);
nor U13769 (N_13769,N_13013,N_13116);
and U13770 (N_13770,N_13542,N_12901);
nand U13771 (N_13771,N_12848,N_13307);
nand U13772 (N_13772,N_12879,N_13485);
nand U13773 (N_13773,N_13422,N_13517);
or U13774 (N_13774,N_13250,N_12836);
xnor U13775 (N_13775,N_13039,N_13435);
nor U13776 (N_13776,N_13078,N_13248);
and U13777 (N_13777,N_13362,N_12897);
nor U13778 (N_13778,N_13357,N_12859);
nor U13779 (N_13779,N_12847,N_13329);
and U13780 (N_13780,N_12909,N_12960);
and U13781 (N_13781,N_13321,N_12944);
xnor U13782 (N_13782,N_13114,N_13096);
nand U13783 (N_13783,N_12880,N_13219);
xor U13784 (N_13784,N_13033,N_12807);
or U13785 (N_13785,N_13175,N_13380);
or U13786 (N_13786,N_13291,N_13042);
and U13787 (N_13787,N_13531,N_13069);
and U13788 (N_13788,N_13182,N_13506);
and U13789 (N_13789,N_13109,N_13280);
and U13790 (N_13790,N_13337,N_13323);
nor U13791 (N_13791,N_13173,N_13204);
xnor U13792 (N_13792,N_13258,N_13457);
or U13793 (N_13793,N_12908,N_13534);
nand U13794 (N_13794,N_13465,N_13262);
or U13795 (N_13795,N_13246,N_13500);
or U13796 (N_13796,N_13469,N_13218);
or U13797 (N_13797,N_13496,N_12815);
nor U13798 (N_13798,N_12966,N_13102);
xor U13799 (N_13799,N_13354,N_13394);
nand U13800 (N_13800,N_13188,N_12951);
nand U13801 (N_13801,N_13510,N_13413);
nor U13802 (N_13802,N_13454,N_12865);
and U13803 (N_13803,N_13064,N_13051);
and U13804 (N_13804,N_13581,N_13267);
xor U13805 (N_13805,N_12817,N_12912);
xor U13806 (N_13806,N_13499,N_12877);
and U13807 (N_13807,N_13468,N_13364);
xor U13808 (N_13808,N_12820,N_13382);
or U13809 (N_13809,N_12831,N_13202);
nor U13810 (N_13810,N_12945,N_13085);
and U13811 (N_13811,N_13079,N_12986);
nand U13812 (N_13812,N_12885,N_13132);
and U13813 (N_13813,N_13390,N_13584);
and U13814 (N_13814,N_12835,N_12832);
xor U13815 (N_13815,N_13070,N_13229);
or U13816 (N_13816,N_12920,N_13170);
nor U13817 (N_13817,N_13593,N_13261);
nand U13818 (N_13818,N_13585,N_13426);
and U13819 (N_13819,N_13586,N_13463);
nand U13820 (N_13820,N_13583,N_13222);
or U13821 (N_13821,N_13338,N_13560);
nand U13822 (N_13822,N_13538,N_13237);
nor U13823 (N_13823,N_13336,N_13437);
or U13824 (N_13824,N_13374,N_13319);
and U13825 (N_13825,N_13432,N_13388);
and U13826 (N_13826,N_13518,N_12943);
nor U13827 (N_13827,N_13155,N_12996);
nand U13828 (N_13828,N_13253,N_13183);
nor U13829 (N_13829,N_13104,N_12959);
nor U13830 (N_13830,N_13264,N_13595);
nor U13831 (N_13831,N_13080,N_12954);
nand U13832 (N_13832,N_13436,N_13036);
nand U13833 (N_13833,N_13004,N_13076);
or U13834 (N_13834,N_12997,N_12931);
nand U13835 (N_13835,N_12889,N_13223);
nor U13836 (N_13836,N_13528,N_12990);
nand U13837 (N_13837,N_13197,N_12871);
nand U13838 (N_13838,N_13148,N_13478);
and U13839 (N_13839,N_13212,N_12928);
nand U13840 (N_13840,N_13360,N_13588);
or U13841 (N_13841,N_13553,N_13587);
or U13842 (N_13842,N_13090,N_13429);
or U13843 (N_13843,N_13448,N_13281);
and U13844 (N_13844,N_12904,N_13292);
and U13845 (N_13845,N_13265,N_13552);
and U13846 (N_13846,N_13410,N_13273);
or U13847 (N_13847,N_13308,N_12994);
xor U13848 (N_13848,N_13217,N_12919);
nor U13849 (N_13849,N_13400,N_13136);
nand U13850 (N_13850,N_13578,N_12894);
xor U13851 (N_13851,N_13317,N_13120);
and U13852 (N_13852,N_13495,N_13211);
nor U13853 (N_13853,N_12979,N_13174);
nand U13854 (N_13854,N_13490,N_12860);
nor U13855 (N_13855,N_12955,N_13163);
nand U13856 (N_13856,N_13536,N_13370);
and U13857 (N_13857,N_13467,N_13570);
nand U13858 (N_13858,N_12936,N_13442);
nor U13859 (N_13859,N_12882,N_13447);
or U13860 (N_13860,N_12957,N_13142);
and U13861 (N_13861,N_13564,N_13295);
or U13862 (N_13862,N_12826,N_12830);
nor U13863 (N_13863,N_13372,N_12801);
and U13864 (N_13864,N_13554,N_13405);
nand U13865 (N_13865,N_13597,N_13590);
or U13866 (N_13866,N_13206,N_12849);
nand U13867 (N_13867,N_12982,N_13007);
nor U13868 (N_13868,N_13054,N_12934);
and U13869 (N_13869,N_13524,N_13414);
nand U13870 (N_13870,N_13089,N_13196);
and U13871 (N_13871,N_12983,N_13158);
or U13872 (N_13872,N_13459,N_12808);
nor U13873 (N_13873,N_12834,N_13571);
nor U13874 (N_13874,N_13231,N_13162);
nand U13875 (N_13875,N_13393,N_12952);
nand U13876 (N_13876,N_12804,N_13127);
nand U13877 (N_13877,N_13558,N_13532);
or U13878 (N_13878,N_13198,N_13092);
or U13879 (N_13879,N_12821,N_13452);
nor U13880 (N_13880,N_12850,N_12841);
nand U13881 (N_13881,N_13097,N_13527);
nand U13882 (N_13882,N_12818,N_13582);
xnor U13883 (N_13883,N_13345,N_13472);
or U13884 (N_13884,N_12913,N_13409);
or U13885 (N_13885,N_13439,N_12923);
xnor U13886 (N_13886,N_13146,N_13220);
nor U13887 (N_13887,N_13002,N_13035);
and U13888 (N_13888,N_12971,N_12842);
and U13889 (N_13889,N_12907,N_13346);
nor U13890 (N_13890,N_12999,N_13507);
nor U13891 (N_13891,N_12995,N_12946);
xor U13892 (N_13892,N_13505,N_12856);
and U13893 (N_13893,N_12922,N_12958);
and U13894 (N_13894,N_13351,N_13168);
and U13895 (N_13895,N_12991,N_13504);
or U13896 (N_13896,N_13575,N_12845);
xnor U13897 (N_13897,N_13141,N_12972);
xnor U13898 (N_13898,N_13368,N_13088);
nand U13899 (N_13899,N_13367,N_13185);
xor U13900 (N_13900,N_13512,N_13123);
and U13901 (N_13901,N_13594,N_13334);
nand U13902 (N_13902,N_12906,N_13358);
nor U13903 (N_13903,N_13464,N_13402);
and U13904 (N_13904,N_12833,N_13131);
nand U13905 (N_13905,N_13449,N_13461);
or U13906 (N_13906,N_13283,N_12942);
or U13907 (N_13907,N_13221,N_12976);
nand U13908 (N_13908,N_13279,N_13190);
xnor U13909 (N_13909,N_12978,N_12873);
and U13910 (N_13910,N_12855,N_13149);
xor U13911 (N_13911,N_13284,N_13353);
xor U13912 (N_13912,N_12881,N_12892);
xor U13913 (N_13913,N_13328,N_13129);
xnor U13914 (N_13914,N_13365,N_13277);
or U13915 (N_13915,N_13046,N_13150);
nor U13916 (N_13916,N_13421,N_13093);
and U13917 (N_13917,N_13285,N_13167);
and U13918 (N_13918,N_13058,N_13547);
or U13919 (N_13919,N_13017,N_13376);
or U13920 (N_13920,N_13003,N_13115);
or U13921 (N_13921,N_13300,N_12854);
nand U13922 (N_13922,N_13000,N_13580);
or U13923 (N_13923,N_13483,N_12940);
nor U13924 (N_13924,N_13539,N_12914);
and U13925 (N_13925,N_13566,N_13125);
nand U13926 (N_13926,N_12893,N_12870);
and U13927 (N_13927,N_13339,N_13344);
xnor U13928 (N_13928,N_13121,N_12910);
xor U13929 (N_13929,N_13443,N_12953);
xor U13930 (N_13930,N_13299,N_13205);
and U13931 (N_13931,N_12828,N_13128);
and U13932 (N_13932,N_13209,N_13181);
xnor U13933 (N_13933,N_13235,N_13270);
nand U13934 (N_13934,N_12895,N_13025);
nor U13935 (N_13935,N_12998,N_12861);
nand U13936 (N_13936,N_13122,N_13107);
xnor U13937 (N_13937,N_12890,N_13028);
nand U13938 (N_13938,N_13599,N_13272);
xor U13939 (N_13939,N_12822,N_12947);
and U13940 (N_13940,N_13015,N_13140);
and U13941 (N_13941,N_13289,N_13124);
or U13942 (N_13942,N_13592,N_13260);
and U13943 (N_13943,N_13152,N_13048);
or U13944 (N_13944,N_13335,N_13014);
nor U13945 (N_13945,N_13256,N_13350);
or U13946 (N_13946,N_13161,N_13596);
nor U13947 (N_13947,N_13567,N_13310);
xnor U13948 (N_13948,N_13355,N_13208);
nor U13949 (N_13949,N_13103,N_13391);
or U13950 (N_13950,N_13006,N_13369);
and U13951 (N_13951,N_13544,N_13049);
or U13952 (N_13952,N_13508,N_13363);
and U13953 (N_13953,N_13195,N_12887);
xnor U13954 (N_13954,N_13371,N_13403);
and U13955 (N_13955,N_13396,N_13255);
nand U13956 (N_13956,N_13180,N_13503);
nand U13957 (N_13957,N_12915,N_13055);
and U13958 (N_13958,N_13275,N_12963);
and U13959 (N_13959,N_13384,N_12812);
xor U13960 (N_13960,N_12917,N_13340);
and U13961 (N_13961,N_12864,N_13480);
and U13962 (N_13962,N_13126,N_13164);
and U13963 (N_13963,N_13522,N_12824);
nand U13964 (N_13964,N_13476,N_13230);
nor U13965 (N_13965,N_12989,N_13009);
nor U13966 (N_13966,N_13444,N_13154);
nor U13967 (N_13967,N_13169,N_13548);
xnor U13968 (N_13968,N_12876,N_13159);
and U13969 (N_13969,N_13331,N_13540);
and U13970 (N_13970,N_13047,N_13176);
or U13971 (N_13971,N_13022,N_13251);
nand U13972 (N_13972,N_13416,N_12933);
or U13973 (N_13973,N_13053,N_13016);
or U13974 (N_13974,N_12965,N_13082);
and U13975 (N_13975,N_13199,N_13240);
or U13976 (N_13976,N_13075,N_12819);
or U13977 (N_13977,N_13491,N_13302);
or U13978 (N_13978,N_13144,N_13172);
nor U13979 (N_13979,N_12939,N_12985);
and U13980 (N_13980,N_13425,N_13569);
nand U13981 (N_13981,N_13407,N_12810);
nand U13982 (N_13982,N_13514,N_13249);
xnor U13983 (N_13983,N_13420,N_13557);
xnor U13984 (N_13984,N_13108,N_13427);
and U13985 (N_13985,N_13192,N_13389);
xor U13986 (N_13986,N_13470,N_13225);
or U13987 (N_13987,N_12888,N_12869);
nor U13988 (N_13988,N_13056,N_12962);
and U13989 (N_13989,N_13214,N_13475);
xor U13990 (N_13990,N_13244,N_12902);
nand U13991 (N_13991,N_12968,N_12811);
or U13992 (N_13992,N_13385,N_13509);
or U13993 (N_13993,N_13591,N_13157);
xor U13994 (N_13994,N_13546,N_13059);
or U13995 (N_13995,N_12905,N_13001);
and U13996 (N_13996,N_13471,N_13278);
and U13997 (N_13997,N_13359,N_12886);
xor U13998 (N_13998,N_13171,N_13160);
xnor U13999 (N_13999,N_13320,N_12961);
and U14000 (N_14000,N_13135,N_13031);
xor U14001 (N_14001,N_13126,N_13522);
or U14002 (N_14002,N_13383,N_13500);
and U14003 (N_14003,N_13413,N_13575);
or U14004 (N_14004,N_13494,N_13451);
xor U14005 (N_14005,N_13541,N_13585);
or U14006 (N_14006,N_13271,N_13503);
or U14007 (N_14007,N_13254,N_12982);
xor U14008 (N_14008,N_13175,N_13556);
xnor U14009 (N_14009,N_12969,N_12822);
nor U14010 (N_14010,N_12892,N_13336);
xor U14011 (N_14011,N_13072,N_13148);
and U14012 (N_14012,N_12981,N_12931);
nor U14013 (N_14013,N_13165,N_13534);
nand U14014 (N_14014,N_13009,N_13534);
nand U14015 (N_14015,N_12927,N_13581);
xor U14016 (N_14016,N_13421,N_13581);
or U14017 (N_14017,N_13279,N_13238);
nand U14018 (N_14018,N_13437,N_13216);
nor U14019 (N_14019,N_13110,N_13584);
nand U14020 (N_14020,N_13336,N_12997);
and U14021 (N_14021,N_13107,N_13399);
or U14022 (N_14022,N_13248,N_13043);
xnor U14023 (N_14023,N_13552,N_12976);
and U14024 (N_14024,N_12931,N_12819);
and U14025 (N_14025,N_13452,N_12815);
nor U14026 (N_14026,N_13581,N_13016);
xnor U14027 (N_14027,N_13374,N_12977);
and U14028 (N_14028,N_13545,N_13577);
and U14029 (N_14029,N_12897,N_13482);
and U14030 (N_14030,N_13264,N_13089);
or U14031 (N_14031,N_13500,N_13529);
xor U14032 (N_14032,N_12911,N_13306);
and U14033 (N_14033,N_12861,N_13025);
or U14034 (N_14034,N_13017,N_13239);
nand U14035 (N_14035,N_13011,N_12842);
nand U14036 (N_14036,N_13061,N_13275);
or U14037 (N_14037,N_13090,N_13342);
or U14038 (N_14038,N_13015,N_12836);
nor U14039 (N_14039,N_13000,N_13119);
and U14040 (N_14040,N_13138,N_13211);
or U14041 (N_14041,N_13465,N_12855);
xor U14042 (N_14042,N_13092,N_13266);
xnor U14043 (N_14043,N_13539,N_13548);
xor U14044 (N_14044,N_12941,N_13347);
nand U14045 (N_14045,N_12857,N_13514);
xor U14046 (N_14046,N_13133,N_12991);
xnor U14047 (N_14047,N_12839,N_13138);
or U14048 (N_14048,N_13182,N_13279);
or U14049 (N_14049,N_13168,N_12948);
and U14050 (N_14050,N_13001,N_13577);
or U14051 (N_14051,N_13303,N_13272);
xor U14052 (N_14052,N_13346,N_13296);
nand U14053 (N_14053,N_13489,N_13561);
and U14054 (N_14054,N_13158,N_13444);
nor U14055 (N_14055,N_13215,N_12815);
and U14056 (N_14056,N_13290,N_12995);
or U14057 (N_14057,N_13064,N_13219);
or U14058 (N_14058,N_13508,N_13401);
xnor U14059 (N_14059,N_13372,N_12968);
or U14060 (N_14060,N_13503,N_13070);
xnor U14061 (N_14061,N_13157,N_12964);
nand U14062 (N_14062,N_13334,N_13120);
or U14063 (N_14063,N_13037,N_13506);
nor U14064 (N_14064,N_12993,N_13469);
or U14065 (N_14065,N_13405,N_13457);
nand U14066 (N_14066,N_13308,N_12873);
and U14067 (N_14067,N_13552,N_13123);
and U14068 (N_14068,N_13402,N_13012);
and U14069 (N_14069,N_13564,N_13031);
nand U14070 (N_14070,N_13248,N_12946);
xor U14071 (N_14071,N_13270,N_12821);
and U14072 (N_14072,N_13316,N_12858);
and U14073 (N_14073,N_13189,N_12868);
nand U14074 (N_14074,N_13424,N_13327);
xnor U14075 (N_14075,N_13179,N_13246);
or U14076 (N_14076,N_13353,N_13058);
or U14077 (N_14077,N_12903,N_13270);
and U14078 (N_14078,N_13013,N_13283);
nand U14079 (N_14079,N_13086,N_13412);
xnor U14080 (N_14080,N_13434,N_12874);
or U14081 (N_14081,N_13355,N_13301);
nand U14082 (N_14082,N_13397,N_13149);
nor U14083 (N_14083,N_13115,N_13386);
or U14084 (N_14084,N_13349,N_13356);
and U14085 (N_14085,N_12825,N_12877);
xor U14086 (N_14086,N_13053,N_13279);
nor U14087 (N_14087,N_13025,N_13466);
nand U14088 (N_14088,N_12968,N_12809);
xnor U14089 (N_14089,N_12845,N_13420);
or U14090 (N_14090,N_13152,N_13123);
nand U14091 (N_14091,N_13328,N_13079);
and U14092 (N_14092,N_12813,N_12877);
and U14093 (N_14093,N_13441,N_13174);
nor U14094 (N_14094,N_13157,N_12920);
and U14095 (N_14095,N_13263,N_13058);
nor U14096 (N_14096,N_12996,N_13126);
and U14097 (N_14097,N_13207,N_13285);
nand U14098 (N_14098,N_13034,N_12836);
nand U14099 (N_14099,N_13563,N_13264);
or U14100 (N_14100,N_13264,N_12941);
nor U14101 (N_14101,N_13287,N_13133);
and U14102 (N_14102,N_13456,N_13294);
nor U14103 (N_14103,N_13462,N_13439);
nor U14104 (N_14104,N_12830,N_13547);
nor U14105 (N_14105,N_12946,N_13588);
or U14106 (N_14106,N_13585,N_13275);
xor U14107 (N_14107,N_13164,N_13458);
xnor U14108 (N_14108,N_12874,N_13094);
or U14109 (N_14109,N_13174,N_12872);
nor U14110 (N_14110,N_13561,N_13474);
or U14111 (N_14111,N_12846,N_13536);
nand U14112 (N_14112,N_13140,N_12952);
nor U14113 (N_14113,N_13256,N_12951);
nand U14114 (N_14114,N_13437,N_13569);
and U14115 (N_14115,N_13594,N_13205);
nand U14116 (N_14116,N_13584,N_13337);
and U14117 (N_14117,N_13062,N_13560);
xor U14118 (N_14118,N_13173,N_12898);
or U14119 (N_14119,N_12868,N_13035);
and U14120 (N_14120,N_13492,N_12843);
nand U14121 (N_14121,N_13084,N_13158);
nor U14122 (N_14122,N_12925,N_13539);
nand U14123 (N_14123,N_13037,N_13292);
and U14124 (N_14124,N_13252,N_13528);
nand U14125 (N_14125,N_13364,N_13422);
nor U14126 (N_14126,N_13512,N_12821);
nand U14127 (N_14127,N_13524,N_13146);
nor U14128 (N_14128,N_13424,N_13478);
and U14129 (N_14129,N_13497,N_13010);
or U14130 (N_14130,N_13358,N_13149);
or U14131 (N_14131,N_13108,N_12979);
nand U14132 (N_14132,N_13225,N_13223);
xor U14133 (N_14133,N_13247,N_13123);
nor U14134 (N_14134,N_13012,N_13214);
nand U14135 (N_14135,N_12922,N_12998);
or U14136 (N_14136,N_13356,N_13059);
or U14137 (N_14137,N_13565,N_13466);
or U14138 (N_14138,N_13238,N_13534);
or U14139 (N_14139,N_13075,N_13352);
and U14140 (N_14140,N_12820,N_12913);
nand U14141 (N_14141,N_13306,N_12803);
and U14142 (N_14142,N_12981,N_13221);
nand U14143 (N_14143,N_13090,N_13567);
xor U14144 (N_14144,N_13141,N_12804);
xnor U14145 (N_14145,N_13255,N_13133);
xnor U14146 (N_14146,N_13125,N_13117);
and U14147 (N_14147,N_13516,N_13422);
nor U14148 (N_14148,N_13279,N_13032);
nand U14149 (N_14149,N_13396,N_13063);
nor U14150 (N_14150,N_12990,N_13298);
and U14151 (N_14151,N_13096,N_13184);
nor U14152 (N_14152,N_13593,N_12858);
xor U14153 (N_14153,N_13312,N_13360);
and U14154 (N_14154,N_13143,N_12965);
xnor U14155 (N_14155,N_13097,N_12990);
and U14156 (N_14156,N_12907,N_12882);
xnor U14157 (N_14157,N_12976,N_12994);
nor U14158 (N_14158,N_13455,N_13536);
xnor U14159 (N_14159,N_13199,N_13080);
xor U14160 (N_14160,N_13054,N_13282);
nor U14161 (N_14161,N_13118,N_12849);
or U14162 (N_14162,N_12947,N_13479);
xnor U14163 (N_14163,N_13381,N_13231);
and U14164 (N_14164,N_13391,N_12922);
nand U14165 (N_14165,N_12933,N_13091);
nand U14166 (N_14166,N_13382,N_13502);
nor U14167 (N_14167,N_13501,N_12996);
nand U14168 (N_14168,N_13452,N_13000);
or U14169 (N_14169,N_13345,N_13577);
and U14170 (N_14170,N_12992,N_12871);
nor U14171 (N_14171,N_13050,N_12846);
and U14172 (N_14172,N_13278,N_13503);
xnor U14173 (N_14173,N_12801,N_13591);
and U14174 (N_14174,N_13360,N_13566);
xor U14175 (N_14175,N_13355,N_12955);
nor U14176 (N_14176,N_13049,N_13373);
and U14177 (N_14177,N_13450,N_13422);
nor U14178 (N_14178,N_12811,N_13108);
nand U14179 (N_14179,N_13262,N_12820);
xor U14180 (N_14180,N_12834,N_13001);
nand U14181 (N_14181,N_12979,N_13081);
and U14182 (N_14182,N_13038,N_13315);
nand U14183 (N_14183,N_13291,N_13279);
xor U14184 (N_14184,N_13511,N_13221);
nand U14185 (N_14185,N_13462,N_13175);
nor U14186 (N_14186,N_13043,N_13016);
nor U14187 (N_14187,N_13515,N_13109);
nor U14188 (N_14188,N_13208,N_13028);
nand U14189 (N_14189,N_13053,N_13062);
xor U14190 (N_14190,N_13248,N_13126);
xnor U14191 (N_14191,N_13161,N_13333);
nand U14192 (N_14192,N_13411,N_13302);
and U14193 (N_14193,N_13380,N_13136);
nand U14194 (N_14194,N_13101,N_13246);
xnor U14195 (N_14195,N_12983,N_13208);
and U14196 (N_14196,N_13292,N_13281);
xnor U14197 (N_14197,N_12989,N_13178);
nand U14198 (N_14198,N_13163,N_13521);
xnor U14199 (N_14199,N_13043,N_12882);
xnor U14200 (N_14200,N_13405,N_13559);
and U14201 (N_14201,N_13596,N_13107);
and U14202 (N_14202,N_12890,N_12913);
nor U14203 (N_14203,N_13227,N_13114);
or U14204 (N_14204,N_12930,N_12833);
xor U14205 (N_14205,N_13326,N_13001);
nor U14206 (N_14206,N_12849,N_13359);
xnor U14207 (N_14207,N_13507,N_13062);
or U14208 (N_14208,N_13156,N_13219);
or U14209 (N_14209,N_13487,N_13037);
nand U14210 (N_14210,N_13226,N_13455);
nor U14211 (N_14211,N_13033,N_13371);
nand U14212 (N_14212,N_13535,N_12932);
or U14213 (N_14213,N_13069,N_13596);
or U14214 (N_14214,N_13396,N_13102);
xnor U14215 (N_14215,N_13011,N_13139);
xnor U14216 (N_14216,N_13546,N_13127);
nand U14217 (N_14217,N_12992,N_13087);
xor U14218 (N_14218,N_13057,N_13054);
nor U14219 (N_14219,N_13138,N_13283);
xnor U14220 (N_14220,N_12852,N_13235);
nor U14221 (N_14221,N_13182,N_12815);
xor U14222 (N_14222,N_13527,N_13090);
and U14223 (N_14223,N_12849,N_13271);
and U14224 (N_14224,N_13283,N_13578);
nand U14225 (N_14225,N_13472,N_13129);
xor U14226 (N_14226,N_12869,N_13270);
nand U14227 (N_14227,N_13224,N_13086);
or U14228 (N_14228,N_13418,N_13023);
xor U14229 (N_14229,N_13172,N_13435);
or U14230 (N_14230,N_12971,N_13142);
and U14231 (N_14231,N_13248,N_13468);
nor U14232 (N_14232,N_13282,N_13464);
and U14233 (N_14233,N_13444,N_13209);
nand U14234 (N_14234,N_13231,N_13489);
nand U14235 (N_14235,N_13544,N_12801);
nor U14236 (N_14236,N_13147,N_13301);
and U14237 (N_14237,N_13263,N_13509);
or U14238 (N_14238,N_12813,N_12810);
and U14239 (N_14239,N_13102,N_13115);
nand U14240 (N_14240,N_13533,N_13258);
xnor U14241 (N_14241,N_13176,N_13334);
or U14242 (N_14242,N_13236,N_13232);
or U14243 (N_14243,N_12983,N_13445);
or U14244 (N_14244,N_13202,N_13142);
nor U14245 (N_14245,N_13388,N_13081);
nor U14246 (N_14246,N_13113,N_13342);
and U14247 (N_14247,N_13142,N_13178);
nand U14248 (N_14248,N_13101,N_12898);
xor U14249 (N_14249,N_13175,N_13070);
nor U14250 (N_14250,N_13291,N_12831);
nand U14251 (N_14251,N_13347,N_12953);
nor U14252 (N_14252,N_13454,N_13453);
or U14253 (N_14253,N_13073,N_13165);
xor U14254 (N_14254,N_12975,N_12903);
xnor U14255 (N_14255,N_12866,N_13523);
nand U14256 (N_14256,N_13512,N_12808);
nand U14257 (N_14257,N_12879,N_12936);
nor U14258 (N_14258,N_13183,N_13524);
nor U14259 (N_14259,N_13572,N_13371);
xnor U14260 (N_14260,N_13524,N_13035);
xnor U14261 (N_14261,N_13525,N_12860);
or U14262 (N_14262,N_13574,N_13379);
nor U14263 (N_14263,N_13301,N_13284);
and U14264 (N_14264,N_12864,N_13340);
or U14265 (N_14265,N_13025,N_13432);
nor U14266 (N_14266,N_12922,N_12848);
xnor U14267 (N_14267,N_13467,N_13553);
nand U14268 (N_14268,N_13571,N_12873);
nand U14269 (N_14269,N_13437,N_13503);
and U14270 (N_14270,N_13357,N_13149);
nand U14271 (N_14271,N_12981,N_13546);
nor U14272 (N_14272,N_12869,N_13075);
nand U14273 (N_14273,N_13453,N_13524);
and U14274 (N_14274,N_12801,N_13374);
and U14275 (N_14275,N_12969,N_13332);
nor U14276 (N_14276,N_13355,N_12935);
or U14277 (N_14277,N_13490,N_13041);
xnor U14278 (N_14278,N_13429,N_13227);
or U14279 (N_14279,N_13580,N_13042);
xnor U14280 (N_14280,N_13490,N_12873);
xnor U14281 (N_14281,N_13006,N_13391);
xnor U14282 (N_14282,N_13235,N_13374);
and U14283 (N_14283,N_13492,N_12944);
and U14284 (N_14284,N_13330,N_12863);
xnor U14285 (N_14285,N_13582,N_12954);
xor U14286 (N_14286,N_13352,N_13171);
nand U14287 (N_14287,N_12941,N_13240);
xnor U14288 (N_14288,N_12966,N_13021);
xor U14289 (N_14289,N_12881,N_13045);
nand U14290 (N_14290,N_12925,N_13545);
nor U14291 (N_14291,N_13446,N_13597);
nand U14292 (N_14292,N_12967,N_13229);
or U14293 (N_14293,N_12971,N_12960);
nor U14294 (N_14294,N_13422,N_13074);
nand U14295 (N_14295,N_13411,N_13079);
nor U14296 (N_14296,N_13294,N_13363);
nor U14297 (N_14297,N_13441,N_12868);
and U14298 (N_14298,N_13463,N_13432);
and U14299 (N_14299,N_13080,N_13003);
or U14300 (N_14300,N_13116,N_13034);
xnor U14301 (N_14301,N_13404,N_13345);
nand U14302 (N_14302,N_13402,N_13115);
nand U14303 (N_14303,N_12820,N_13059);
nand U14304 (N_14304,N_12918,N_13037);
or U14305 (N_14305,N_13308,N_13436);
nor U14306 (N_14306,N_13513,N_12940);
xor U14307 (N_14307,N_13196,N_12863);
nand U14308 (N_14308,N_13161,N_12951);
xnor U14309 (N_14309,N_12908,N_13303);
xnor U14310 (N_14310,N_12910,N_13109);
and U14311 (N_14311,N_13579,N_13344);
nand U14312 (N_14312,N_13134,N_12802);
or U14313 (N_14313,N_12824,N_13521);
xnor U14314 (N_14314,N_12941,N_13055);
or U14315 (N_14315,N_13293,N_12833);
or U14316 (N_14316,N_12864,N_13352);
nor U14317 (N_14317,N_13435,N_12833);
and U14318 (N_14318,N_12911,N_13299);
nor U14319 (N_14319,N_13283,N_13186);
nor U14320 (N_14320,N_13553,N_12837);
nor U14321 (N_14321,N_13064,N_13369);
and U14322 (N_14322,N_13002,N_13330);
xor U14323 (N_14323,N_13344,N_13588);
or U14324 (N_14324,N_13543,N_13198);
nor U14325 (N_14325,N_12817,N_13331);
or U14326 (N_14326,N_13555,N_13301);
or U14327 (N_14327,N_13368,N_13053);
and U14328 (N_14328,N_13312,N_13222);
or U14329 (N_14329,N_13355,N_13239);
nand U14330 (N_14330,N_13401,N_13065);
xor U14331 (N_14331,N_13339,N_13079);
and U14332 (N_14332,N_13252,N_13267);
or U14333 (N_14333,N_13415,N_13412);
xor U14334 (N_14334,N_12832,N_13215);
and U14335 (N_14335,N_13015,N_13399);
xnor U14336 (N_14336,N_13299,N_13050);
or U14337 (N_14337,N_12961,N_13002);
nand U14338 (N_14338,N_13358,N_13518);
xor U14339 (N_14339,N_12882,N_12809);
and U14340 (N_14340,N_13182,N_13563);
nand U14341 (N_14341,N_13435,N_12841);
xor U14342 (N_14342,N_13551,N_13364);
nand U14343 (N_14343,N_13352,N_13419);
nor U14344 (N_14344,N_13563,N_12971);
nand U14345 (N_14345,N_13024,N_13362);
nand U14346 (N_14346,N_13519,N_12847);
nor U14347 (N_14347,N_13244,N_13020);
nor U14348 (N_14348,N_13559,N_13401);
nor U14349 (N_14349,N_12942,N_13365);
xnor U14350 (N_14350,N_12897,N_13540);
and U14351 (N_14351,N_12913,N_12824);
and U14352 (N_14352,N_13385,N_13491);
and U14353 (N_14353,N_13408,N_13202);
nor U14354 (N_14354,N_13485,N_13019);
or U14355 (N_14355,N_13259,N_12923);
nand U14356 (N_14356,N_13323,N_12834);
and U14357 (N_14357,N_12921,N_13575);
xnor U14358 (N_14358,N_13304,N_13063);
xnor U14359 (N_14359,N_13203,N_13204);
xnor U14360 (N_14360,N_13150,N_13429);
nand U14361 (N_14361,N_13560,N_13444);
nor U14362 (N_14362,N_13379,N_13565);
or U14363 (N_14363,N_13526,N_13281);
nand U14364 (N_14364,N_12888,N_13191);
and U14365 (N_14365,N_13328,N_12903);
nor U14366 (N_14366,N_13439,N_13449);
nor U14367 (N_14367,N_12956,N_12927);
and U14368 (N_14368,N_13393,N_13458);
or U14369 (N_14369,N_13390,N_13226);
and U14370 (N_14370,N_13475,N_13247);
nor U14371 (N_14371,N_13340,N_13404);
xnor U14372 (N_14372,N_13333,N_12815);
xor U14373 (N_14373,N_13320,N_13153);
xor U14374 (N_14374,N_13181,N_13546);
nor U14375 (N_14375,N_13099,N_13120);
nand U14376 (N_14376,N_13219,N_12964);
nor U14377 (N_14377,N_13222,N_13487);
and U14378 (N_14378,N_13150,N_13139);
nand U14379 (N_14379,N_13050,N_13102);
or U14380 (N_14380,N_13105,N_13333);
xor U14381 (N_14381,N_13321,N_13147);
nand U14382 (N_14382,N_12987,N_13030);
xor U14383 (N_14383,N_13506,N_13268);
or U14384 (N_14384,N_13168,N_12896);
and U14385 (N_14385,N_12893,N_13282);
nand U14386 (N_14386,N_13097,N_13530);
or U14387 (N_14387,N_13543,N_13122);
nand U14388 (N_14388,N_12883,N_13212);
or U14389 (N_14389,N_13532,N_12846);
xnor U14390 (N_14390,N_13252,N_13092);
and U14391 (N_14391,N_12825,N_13359);
and U14392 (N_14392,N_13192,N_13158);
and U14393 (N_14393,N_13471,N_13450);
xnor U14394 (N_14394,N_13054,N_13155);
nand U14395 (N_14395,N_13128,N_13296);
or U14396 (N_14396,N_13361,N_12826);
nor U14397 (N_14397,N_12904,N_13132);
xor U14398 (N_14398,N_12826,N_12997);
and U14399 (N_14399,N_13442,N_13247);
xnor U14400 (N_14400,N_13632,N_14184);
and U14401 (N_14401,N_14203,N_14251);
nor U14402 (N_14402,N_14358,N_14013);
xnor U14403 (N_14403,N_14360,N_14172);
or U14404 (N_14404,N_13937,N_13949);
and U14405 (N_14405,N_14367,N_13887);
or U14406 (N_14406,N_13778,N_13888);
and U14407 (N_14407,N_13751,N_13697);
or U14408 (N_14408,N_14258,N_14081);
xnor U14409 (N_14409,N_14376,N_14120);
and U14410 (N_14410,N_14180,N_13869);
nor U14411 (N_14411,N_14338,N_14016);
nand U14412 (N_14412,N_13621,N_14045);
xor U14413 (N_14413,N_13764,N_13940);
or U14414 (N_14414,N_13886,N_14350);
nand U14415 (N_14415,N_14359,N_13923);
nand U14416 (N_14416,N_14344,N_13950);
nor U14417 (N_14417,N_14038,N_13918);
nor U14418 (N_14418,N_14306,N_13772);
or U14419 (N_14419,N_13720,N_13748);
xor U14420 (N_14420,N_14044,N_13699);
nand U14421 (N_14421,N_14288,N_13788);
nand U14422 (N_14422,N_13798,N_14036);
nand U14423 (N_14423,N_13873,N_13759);
xnor U14424 (N_14424,N_14160,N_14062);
xnor U14425 (N_14425,N_14389,N_13885);
nand U14426 (N_14426,N_13954,N_14060);
nor U14427 (N_14427,N_13831,N_13718);
or U14428 (N_14428,N_14006,N_14148);
or U14429 (N_14429,N_13681,N_13855);
xnor U14430 (N_14430,N_14283,N_13682);
nand U14431 (N_14431,N_13928,N_13799);
or U14432 (N_14432,N_14216,N_14284);
and U14433 (N_14433,N_14051,N_13670);
or U14434 (N_14434,N_13825,N_13704);
or U14435 (N_14435,N_14304,N_13616);
nor U14436 (N_14436,N_13803,N_14014);
xnor U14437 (N_14437,N_13776,N_14147);
xnor U14438 (N_14438,N_14012,N_13837);
nor U14439 (N_14439,N_14249,N_13932);
nand U14440 (N_14440,N_14351,N_13696);
xor U14441 (N_14441,N_13854,N_14110);
or U14442 (N_14442,N_14255,N_14276);
or U14443 (N_14443,N_13775,N_13866);
xnor U14444 (N_14444,N_14121,N_14163);
nor U14445 (N_14445,N_14289,N_13677);
or U14446 (N_14446,N_13844,N_14113);
or U14447 (N_14447,N_13847,N_14280);
nand U14448 (N_14448,N_14159,N_14399);
nor U14449 (N_14449,N_14291,N_13868);
xor U14450 (N_14450,N_14073,N_13604);
nor U14451 (N_14451,N_14167,N_14272);
and U14452 (N_14452,N_13979,N_13691);
or U14453 (N_14453,N_14202,N_13724);
or U14454 (N_14454,N_14083,N_14250);
nor U14455 (N_14455,N_13781,N_14293);
nand U14456 (N_14456,N_14310,N_14264);
and U14457 (N_14457,N_13802,N_14221);
and U14458 (N_14458,N_14381,N_13732);
xnor U14459 (N_14459,N_14231,N_13882);
and U14460 (N_14460,N_14212,N_14312);
nor U14461 (N_14461,N_14108,N_13617);
and U14462 (N_14462,N_13782,N_13832);
or U14463 (N_14463,N_13636,N_14087);
or U14464 (N_14464,N_13629,N_13952);
or U14465 (N_14465,N_14240,N_13678);
xnor U14466 (N_14466,N_14232,N_14230);
nand U14467 (N_14467,N_14179,N_14273);
or U14468 (N_14468,N_13602,N_14089);
and U14469 (N_14469,N_14109,N_14329);
nor U14470 (N_14470,N_13785,N_13653);
xnor U14471 (N_14471,N_14186,N_14315);
nor U14472 (N_14472,N_14377,N_14100);
nor U14473 (N_14473,N_13717,N_13660);
nor U14474 (N_14474,N_14365,N_13620);
nand U14475 (N_14475,N_13809,N_14205);
xor U14476 (N_14476,N_13614,N_14257);
nand U14477 (N_14477,N_14352,N_14271);
xnor U14478 (N_14478,N_14104,N_14088);
or U14479 (N_14479,N_14394,N_13944);
nand U14480 (N_14480,N_14197,N_14170);
and U14481 (N_14481,N_13841,N_14064);
nor U14482 (N_14482,N_14139,N_14114);
nor U14483 (N_14483,N_14238,N_13739);
or U14484 (N_14484,N_14227,N_14301);
nor U14485 (N_14485,N_13730,N_13878);
and U14486 (N_14486,N_13679,N_13771);
nand U14487 (N_14487,N_13813,N_13713);
nor U14488 (N_14488,N_14134,N_13702);
nor U14489 (N_14489,N_14026,N_13667);
or U14490 (N_14490,N_14298,N_13919);
nand U14491 (N_14491,N_13880,N_14164);
xnor U14492 (N_14492,N_13669,N_14369);
nand U14493 (N_14493,N_14286,N_13773);
nand U14494 (N_14494,N_14269,N_13715);
or U14495 (N_14495,N_13624,N_14252);
nor U14496 (N_14496,N_14181,N_14387);
xnor U14497 (N_14497,N_13926,N_13845);
or U14498 (N_14498,N_14009,N_13676);
nand U14499 (N_14499,N_14319,N_14029);
or U14500 (N_14500,N_14101,N_14028);
and U14501 (N_14501,N_13904,N_13701);
and U14502 (N_14502,N_13714,N_13839);
and U14503 (N_14503,N_13729,N_13700);
nand U14504 (N_14504,N_13849,N_14018);
and U14505 (N_14505,N_13884,N_13630);
nand U14506 (N_14506,N_13946,N_14347);
nand U14507 (N_14507,N_14124,N_14311);
xor U14508 (N_14508,N_14074,N_14219);
nand U14509 (N_14509,N_14270,N_13687);
or U14510 (N_14510,N_14204,N_13897);
nor U14511 (N_14511,N_14382,N_13953);
nor U14512 (N_14512,N_13978,N_14070);
and U14513 (N_14513,N_13655,N_14063);
or U14514 (N_14514,N_14162,N_13820);
nand U14515 (N_14515,N_13601,N_13605);
xor U14516 (N_14516,N_13685,N_13942);
nor U14517 (N_14517,N_14225,N_14210);
nand U14518 (N_14518,N_14085,N_13684);
nand U14519 (N_14519,N_14396,N_14265);
nand U14520 (N_14520,N_13625,N_14058);
nand U14521 (N_14521,N_13637,N_14052);
and U14522 (N_14522,N_13780,N_13977);
nor U14523 (N_14523,N_13640,N_13826);
nand U14524 (N_14524,N_13902,N_13892);
xnor U14525 (N_14525,N_14322,N_13976);
nor U14526 (N_14526,N_13628,N_14174);
xor U14527 (N_14527,N_14048,N_13984);
nor U14528 (N_14528,N_13657,N_13786);
xor U14529 (N_14529,N_14041,N_13933);
nand U14530 (N_14530,N_14155,N_13931);
or U14531 (N_14531,N_14379,N_13924);
nand U14532 (N_14532,N_14127,N_14046);
nor U14533 (N_14533,N_14395,N_13816);
nor U14534 (N_14534,N_13666,N_14066);
xnor U14535 (N_14535,N_13883,N_14099);
and U14536 (N_14536,N_14175,N_13683);
xnor U14537 (N_14537,N_14326,N_13703);
nand U14538 (N_14538,N_14132,N_13790);
nand U14539 (N_14539,N_13992,N_14072);
xor U14540 (N_14540,N_13642,N_14043);
or U14541 (N_14541,N_13962,N_14300);
or U14542 (N_14542,N_14002,N_13770);
or U14543 (N_14543,N_13765,N_13983);
nor U14544 (N_14544,N_14130,N_14305);
or U14545 (N_14545,N_14171,N_13688);
nand U14546 (N_14546,N_14214,N_14198);
xnor U14547 (N_14547,N_13804,N_13861);
and U14548 (N_14548,N_13757,N_13603);
nand U14549 (N_14549,N_13671,N_14285);
xnor U14550 (N_14550,N_13903,N_14076);
nor U14551 (N_14551,N_13943,N_14321);
xor U14552 (N_14552,N_13857,N_14390);
or U14553 (N_14553,N_14373,N_14111);
and U14554 (N_14554,N_14268,N_14011);
and U14555 (N_14555,N_13999,N_13608);
nor U14556 (N_14556,N_13905,N_14362);
xor U14557 (N_14557,N_13900,N_13870);
nor U14558 (N_14558,N_14299,N_14176);
and U14559 (N_14559,N_13898,N_14146);
xnor U14560 (N_14560,N_13740,N_13945);
xor U14561 (N_14561,N_13758,N_14151);
and U14562 (N_14562,N_14375,N_14342);
nand U14563 (N_14563,N_14126,N_13853);
and U14564 (N_14564,N_13663,N_13830);
xnor U14565 (N_14565,N_13941,N_13735);
or U14566 (N_14566,N_13967,N_13793);
and U14567 (N_14567,N_14364,N_14090);
or U14568 (N_14568,N_13982,N_14363);
and U14569 (N_14569,N_14226,N_13737);
xnor U14570 (N_14570,N_14316,N_13817);
xnor U14571 (N_14571,N_13745,N_14357);
or U14572 (N_14572,N_14247,N_13647);
and U14573 (N_14573,N_13988,N_13912);
xor U14574 (N_14574,N_13760,N_14086);
and U14575 (N_14575,N_13731,N_14281);
nor U14576 (N_14576,N_13960,N_14190);
nand U14577 (N_14577,N_13618,N_14224);
nand U14578 (N_14578,N_14324,N_13695);
xor U14579 (N_14579,N_13925,N_13733);
and U14580 (N_14580,N_14200,N_13889);
nand U14581 (N_14581,N_14333,N_14339);
nor U14582 (N_14582,N_13801,N_14034);
nand U14583 (N_14583,N_13744,N_14267);
xor U14584 (N_14584,N_14196,N_14125);
and U14585 (N_14585,N_14173,N_14095);
or U14586 (N_14586,N_13774,N_14290);
nand U14587 (N_14587,N_13690,N_13795);
or U14588 (N_14588,N_14079,N_14242);
nor U14589 (N_14589,N_13656,N_13843);
nand U14590 (N_14590,N_14065,N_13808);
and U14591 (N_14591,N_14136,N_13694);
nand U14592 (N_14592,N_13929,N_13654);
nor U14593 (N_14593,N_14361,N_14296);
and U14594 (N_14594,N_13749,N_13922);
and U14595 (N_14595,N_14145,N_14010);
and U14596 (N_14596,N_14131,N_13916);
nand U14597 (N_14597,N_14235,N_14030);
or U14598 (N_14598,N_13914,N_13964);
nand U14599 (N_14599,N_14133,N_13867);
nor U14600 (N_14600,N_14335,N_14185);
xor U14601 (N_14601,N_14135,N_13895);
nand U14602 (N_14602,N_14047,N_14022);
xor U14603 (N_14603,N_14187,N_13651);
nand U14604 (N_14604,N_13846,N_13947);
nand U14605 (N_14605,N_13862,N_13917);
or U14606 (N_14606,N_14385,N_13712);
and U14607 (N_14607,N_13692,N_14209);
nand U14608 (N_14608,N_13996,N_13767);
and U14609 (N_14609,N_14031,N_14115);
and U14610 (N_14610,N_14246,N_14093);
nand U14611 (N_14611,N_13973,N_14349);
xor U14612 (N_14612,N_14384,N_13851);
and U14613 (N_14613,N_14330,N_13990);
and U14614 (N_14614,N_14161,N_14017);
nor U14615 (N_14615,N_13934,N_14309);
and U14616 (N_14616,N_13961,N_13913);
xnor U14617 (N_14617,N_13686,N_14348);
and U14618 (N_14618,N_14150,N_14222);
nand U14619 (N_14619,N_13756,N_14112);
nand U14620 (N_14620,N_13958,N_14393);
or U14621 (N_14621,N_14346,N_13645);
and U14622 (N_14622,N_13705,N_13633);
nor U14623 (N_14623,N_14040,N_14292);
xnor U14624 (N_14624,N_14388,N_14194);
nor U14625 (N_14625,N_13815,N_14071);
nand U14626 (N_14626,N_14295,N_14206);
and U14627 (N_14627,N_13622,N_13672);
nor U14628 (N_14628,N_13865,N_14340);
xnor U14629 (N_14629,N_14102,N_13980);
and U14630 (N_14630,N_14117,N_14039);
nand U14631 (N_14631,N_14241,N_14165);
xnor U14632 (N_14632,N_13649,N_13674);
nand U14633 (N_14633,N_13863,N_14239);
nand U14634 (N_14634,N_14201,N_14067);
and U14635 (N_14635,N_13634,N_13859);
nand U14636 (N_14636,N_13787,N_13899);
or U14637 (N_14637,N_14118,N_13728);
and U14638 (N_14638,N_14157,N_14019);
and U14639 (N_14639,N_13709,N_13959);
nor U14640 (N_14640,N_13626,N_13783);
xor U14641 (N_14641,N_14059,N_14211);
nand U14642 (N_14642,N_14182,N_13747);
or U14643 (N_14643,N_14025,N_13907);
nand U14644 (N_14644,N_14094,N_13639);
xor U14645 (N_14645,N_13811,N_14213);
nor U14646 (N_14646,N_13779,N_13675);
nand U14647 (N_14647,N_14138,N_13723);
nor U14648 (N_14648,N_14003,N_14287);
nor U14649 (N_14649,N_14233,N_13908);
xor U14650 (N_14650,N_14137,N_13750);
or U14651 (N_14651,N_13698,N_14374);
nor U14652 (N_14652,N_13741,N_13890);
nor U14653 (N_14653,N_13842,N_14398);
and U14654 (N_14654,N_14106,N_13819);
or U14655 (N_14655,N_14020,N_14005);
nor U14656 (N_14656,N_14103,N_13643);
xor U14657 (N_14657,N_13935,N_14220);
and U14658 (N_14658,N_14237,N_13963);
nand U14659 (N_14659,N_13727,N_13818);
or U14660 (N_14660,N_14218,N_13743);
nor U14661 (N_14661,N_14229,N_13930);
or U14662 (N_14662,N_14116,N_14234);
xor U14663 (N_14663,N_14320,N_13951);
nor U14664 (N_14664,N_14080,N_13650);
nor U14665 (N_14665,N_14015,N_14154);
nor U14666 (N_14666,N_13600,N_14336);
and U14667 (N_14667,N_13829,N_14050);
or U14668 (N_14668,N_14078,N_13769);
xor U14669 (N_14669,N_14279,N_14207);
nor U14670 (N_14670,N_13989,N_13864);
nor U14671 (N_14671,N_14345,N_13822);
and U14672 (N_14672,N_13644,N_14023);
xnor U14673 (N_14673,N_13874,N_13800);
xor U14674 (N_14674,N_13607,N_13693);
xor U14675 (N_14675,N_14366,N_14192);
nor U14676 (N_14676,N_14332,N_14189);
and U14677 (N_14677,N_14323,N_13920);
nand U14678 (N_14678,N_13613,N_13664);
or U14679 (N_14679,N_13646,N_14024);
xnor U14680 (N_14680,N_13661,N_13658);
or U14681 (N_14681,N_14259,N_13840);
xnor U14682 (N_14682,N_13734,N_13668);
or U14683 (N_14683,N_14098,N_13762);
xor U14684 (N_14684,N_13957,N_14027);
or U14685 (N_14685,N_14123,N_14391);
xnor U14686 (N_14686,N_13777,N_13891);
or U14687 (N_14687,N_13761,N_14193);
or U14688 (N_14688,N_13726,N_14314);
nand U14689 (N_14689,N_13796,N_13936);
or U14690 (N_14690,N_14037,N_13986);
or U14691 (N_14691,N_14278,N_13738);
xnor U14692 (N_14692,N_14282,N_13652);
nand U14693 (N_14693,N_13719,N_13966);
xor U14694 (N_14694,N_14128,N_13673);
xor U14695 (N_14695,N_14008,N_14397);
nor U14696 (N_14696,N_13807,N_13623);
or U14697 (N_14697,N_13710,N_13828);
nor U14698 (N_14698,N_13615,N_14069);
xor U14699 (N_14699,N_14077,N_13665);
nor U14700 (N_14700,N_13766,N_13721);
nor U14701 (N_14701,N_13707,N_14354);
xor U14702 (N_14702,N_13994,N_13806);
or U14703 (N_14703,N_14096,N_14318);
nor U14704 (N_14704,N_13906,N_14107);
or U14705 (N_14705,N_13725,N_14277);
and U14706 (N_14706,N_14275,N_13970);
or U14707 (N_14707,N_13894,N_14371);
nand U14708 (N_14708,N_14302,N_14274);
xor U14709 (N_14709,N_14177,N_13974);
xnor U14710 (N_14710,N_14217,N_14004);
nor U14711 (N_14711,N_14254,N_13814);
nand U14712 (N_14712,N_14325,N_13852);
and U14713 (N_14713,N_13827,N_14152);
and U14714 (N_14714,N_13805,N_13755);
xnor U14715 (N_14715,N_14243,N_13948);
and U14716 (N_14716,N_14208,N_14256);
or U14717 (N_14717,N_13875,N_13631);
nor U14718 (N_14718,N_13662,N_14303);
nor U14719 (N_14719,N_13835,N_14119);
or U14720 (N_14720,N_14055,N_13792);
and U14721 (N_14721,N_13838,N_14084);
xor U14722 (N_14722,N_13969,N_13850);
nand U14723 (N_14723,N_14337,N_13911);
xnor U14724 (N_14724,N_13985,N_13768);
xor U14725 (N_14725,N_13641,N_14053);
nor U14726 (N_14726,N_14156,N_14334);
xnor U14727 (N_14727,N_13810,N_14383);
nor U14728 (N_14728,N_14223,N_13821);
and U14729 (N_14729,N_14178,N_14328);
nor U14730 (N_14730,N_13921,N_14392);
and U14731 (N_14731,N_13711,N_13833);
nor U14732 (N_14732,N_14158,N_13909);
xnor U14733 (N_14733,N_14263,N_13789);
xor U14734 (N_14734,N_14032,N_14042);
nand U14735 (N_14735,N_14353,N_13746);
xor U14736 (N_14736,N_13879,N_13659);
nor U14737 (N_14737,N_14035,N_13635);
or U14738 (N_14738,N_14141,N_14356);
nor U14739 (N_14739,N_13824,N_13716);
xor U14740 (N_14740,N_14140,N_14056);
nand U14741 (N_14741,N_14097,N_14199);
or U14742 (N_14742,N_13901,N_13910);
nor U14743 (N_14743,N_13939,N_13872);
nand U14744 (N_14744,N_14236,N_14091);
xor U14745 (N_14745,N_14122,N_13871);
and U14746 (N_14746,N_14380,N_14183);
nand U14747 (N_14747,N_13971,N_13938);
xnor U14748 (N_14748,N_14215,N_13860);
nand U14749 (N_14749,N_14092,N_14355);
nor U14750 (N_14750,N_14143,N_14168);
and U14751 (N_14751,N_14153,N_14372);
nor U14752 (N_14752,N_13610,N_13752);
or U14753 (N_14753,N_13627,N_14191);
nor U14754 (N_14754,N_14308,N_14068);
or U14755 (N_14755,N_14341,N_13611);
nand U14756 (N_14756,N_14169,N_13784);
or U14757 (N_14757,N_13881,N_14331);
nor U14758 (N_14758,N_13791,N_13956);
nand U14759 (N_14759,N_13742,N_14075);
nor U14760 (N_14760,N_13998,N_13856);
nand U14761 (N_14761,N_13708,N_13995);
nor U14762 (N_14762,N_13965,N_14262);
or U14763 (N_14763,N_13997,N_14378);
nor U14764 (N_14764,N_14007,N_14082);
xor U14765 (N_14765,N_13968,N_13893);
nand U14766 (N_14766,N_14188,N_13612);
or U14767 (N_14767,N_14000,N_13794);
xor U14768 (N_14768,N_14144,N_14244);
nand U14769 (N_14769,N_13993,N_14061);
and U14770 (N_14770,N_13754,N_14033);
xor U14771 (N_14771,N_14343,N_13848);
and U14772 (N_14772,N_13877,N_14386);
and U14773 (N_14773,N_14260,N_13915);
nor U14774 (N_14774,N_14368,N_13858);
and U14775 (N_14775,N_14142,N_13834);
nor U14776 (N_14776,N_14266,N_13812);
and U14777 (N_14777,N_13955,N_13609);
xnor U14778 (N_14778,N_13991,N_14253);
and U14779 (N_14779,N_13972,N_13836);
nand U14780 (N_14780,N_14245,N_13736);
and U14781 (N_14781,N_13981,N_14307);
nand U14782 (N_14782,N_14195,N_13797);
xor U14783 (N_14783,N_14294,N_14054);
and U14784 (N_14784,N_14313,N_14327);
xor U14785 (N_14785,N_14297,N_13722);
nor U14786 (N_14786,N_13927,N_13606);
nor U14787 (N_14787,N_14317,N_14057);
nand U14788 (N_14788,N_13876,N_13975);
or U14789 (N_14789,N_13689,N_14228);
and U14790 (N_14790,N_13763,N_13896);
nand U14791 (N_14791,N_13987,N_14248);
and U14792 (N_14792,N_13619,N_14049);
xor U14793 (N_14793,N_13753,N_13823);
nor U14794 (N_14794,N_14261,N_13680);
nor U14795 (N_14795,N_13638,N_13706);
nor U14796 (N_14796,N_14105,N_14021);
and U14797 (N_14797,N_14129,N_13648);
nand U14798 (N_14798,N_14001,N_14166);
and U14799 (N_14799,N_14149,N_14370);
nor U14800 (N_14800,N_13778,N_14004);
nand U14801 (N_14801,N_14331,N_14311);
nand U14802 (N_14802,N_14291,N_14265);
nor U14803 (N_14803,N_13994,N_13953);
xnor U14804 (N_14804,N_14376,N_13642);
nand U14805 (N_14805,N_13821,N_14135);
nor U14806 (N_14806,N_13957,N_13811);
or U14807 (N_14807,N_13724,N_14121);
and U14808 (N_14808,N_13788,N_13691);
nor U14809 (N_14809,N_14162,N_14064);
nand U14810 (N_14810,N_13618,N_13609);
or U14811 (N_14811,N_14322,N_13969);
nand U14812 (N_14812,N_14212,N_14045);
and U14813 (N_14813,N_13970,N_14311);
nor U14814 (N_14814,N_14141,N_14128);
nand U14815 (N_14815,N_13709,N_14288);
xor U14816 (N_14816,N_14270,N_13693);
or U14817 (N_14817,N_14243,N_13836);
nor U14818 (N_14818,N_14370,N_13634);
nor U14819 (N_14819,N_13706,N_14107);
or U14820 (N_14820,N_13798,N_14270);
xor U14821 (N_14821,N_14002,N_13898);
nand U14822 (N_14822,N_14274,N_13688);
and U14823 (N_14823,N_14357,N_13927);
nand U14824 (N_14824,N_13843,N_13727);
and U14825 (N_14825,N_13693,N_13774);
nor U14826 (N_14826,N_13726,N_14189);
nor U14827 (N_14827,N_14166,N_13799);
nor U14828 (N_14828,N_14050,N_14052);
or U14829 (N_14829,N_13967,N_13748);
nand U14830 (N_14830,N_14055,N_14319);
xnor U14831 (N_14831,N_14220,N_14261);
and U14832 (N_14832,N_13713,N_13984);
xnor U14833 (N_14833,N_14046,N_14362);
nor U14834 (N_14834,N_14302,N_13640);
xnor U14835 (N_14835,N_13859,N_14367);
nand U14836 (N_14836,N_14350,N_14033);
xnor U14837 (N_14837,N_14063,N_13711);
or U14838 (N_14838,N_13777,N_14060);
or U14839 (N_14839,N_14399,N_14364);
and U14840 (N_14840,N_13610,N_14283);
nor U14841 (N_14841,N_13748,N_14047);
nor U14842 (N_14842,N_13609,N_13694);
or U14843 (N_14843,N_14272,N_14307);
or U14844 (N_14844,N_14340,N_13821);
xnor U14845 (N_14845,N_14295,N_13756);
or U14846 (N_14846,N_14267,N_14210);
and U14847 (N_14847,N_14204,N_14286);
or U14848 (N_14848,N_14345,N_14327);
and U14849 (N_14849,N_14150,N_13952);
nand U14850 (N_14850,N_14042,N_14184);
nor U14851 (N_14851,N_13749,N_14236);
and U14852 (N_14852,N_13980,N_13602);
and U14853 (N_14853,N_13715,N_13703);
nand U14854 (N_14854,N_14286,N_13663);
nor U14855 (N_14855,N_14217,N_14285);
xnor U14856 (N_14856,N_14135,N_13658);
and U14857 (N_14857,N_13676,N_13862);
xnor U14858 (N_14858,N_14252,N_14200);
and U14859 (N_14859,N_13868,N_13941);
xor U14860 (N_14860,N_14175,N_14038);
or U14861 (N_14861,N_14068,N_13806);
or U14862 (N_14862,N_14151,N_14019);
and U14863 (N_14863,N_14340,N_14135);
nor U14864 (N_14864,N_14367,N_13820);
and U14865 (N_14865,N_13917,N_13600);
or U14866 (N_14866,N_14378,N_14383);
or U14867 (N_14867,N_13724,N_13607);
and U14868 (N_14868,N_13642,N_13787);
nand U14869 (N_14869,N_13785,N_13611);
xor U14870 (N_14870,N_14387,N_13994);
nand U14871 (N_14871,N_13641,N_13992);
or U14872 (N_14872,N_13978,N_14286);
xnor U14873 (N_14873,N_13669,N_14390);
or U14874 (N_14874,N_14146,N_13839);
and U14875 (N_14875,N_13862,N_13841);
nor U14876 (N_14876,N_13829,N_14201);
or U14877 (N_14877,N_14263,N_14040);
nand U14878 (N_14878,N_14112,N_13733);
nor U14879 (N_14879,N_14272,N_13796);
nand U14880 (N_14880,N_14068,N_13975);
and U14881 (N_14881,N_13654,N_13625);
nand U14882 (N_14882,N_14148,N_14198);
or U14883 (N_14883,N_13679,N_13690);
and U14884 (N_14884,N_14276,N_14244);
or U14885 (N_14885,N_14057,N_13726);
xor U14886 (N_14886,N_13867,N_14055);
xor U14887 (N_14887,N_13700,N_14298);
xor U14888 (N_14888,N_14330,N_14151);
or U14889 (N_14889,N_14332,N_14036);
nor U14890 (N_14890,N_13718,N_13749);
and U14891 (N_14891,N_14246,N_13919);
nor U14892 (N_14892,N_13617,N_13825);
nor U14893 (N_14893,N_13736,N_14181);
xor U14894 (N_14894,N_14103,N_13707);
nand U14895 (N_14895,N_13678,N_13915);
and U14896 (N_14896,N_14222,N_14179);
nor U14897 (N_14897,N_13938,N_14081);
and U14898 (N_14898,N_13839,N_13868);
nor U14899 (N_14899,N_13864,N_13957);
and U14900 (N_14900,N_14148,N_14358);
and U14901 (N_14901,N_14397,N_14091);
or U14902 (N_14902,N_14253,N_13654);
nor U14903 (N_14903,N_13964,N_14246);
and U14904 (N_14904,N_13899,N_14380);
nor U14905 (N_14905,N_14103,N_14183);
nand U14906 (N_14906,N_14317,N_14014);
nand U14907 (N_14907,N_14133,N_13992);
nand U14908 (N_14908,N_14280,N_13745);
nand U14909 (N_14909,N_14196,N_13996);
nor U14910 (N_14910,N_13786,N_14351);
xor U14911 (N_14911,N_14188,N_14093);
nand U14912 (N_14912,N_13954,N_13946);
nor U14913 (N_14913,N_14106,N_14024);
nor U14914 (N_14914,N_13867,N_13999);
xor U14915 (N_14915,N_13662,N_14389);
or U14916 (N_14916,N_14189,N_14373);
or U14917 (N_14917,N_14122,N_13669);
or U14918 (N_14918,N_14119,N_13961);
nor U14919 (N_14919,N_14087,N_13724);
nor U14920 (N_14920,N_13794,N_13894);
nand U14921 (N_14921,N_13600,N_13663);
or U14922 (N_14922,N_13635,N_13903);
or U14923 (N_14923,N_13635,N_13722);
nor U14924 (N_14924,N_13926,N_13848);
and U14925 (N_14925,N_13953,N_14338);
nor U14926 (N_14926,N_14372,N_14361);
nand U14927 (N_14927,N_14373,N_13961);
nor U14928 (N_14928,N_13978,N_14392);
nand U14929 (N_14929,N_14295,N_13664);
or U14930 (N_14930,N_14020,N_13786);
nor U14931 (N_14931,N_14021,N_13998);
and U14932 (N_14932,N_14145,N_13848);
nor U14933 (N_14933,N_14053,N_14045);
and U14934 (N_14934,N_14309,N_13978);
nor U14935 (N_14935,N_14341,N_14245);
nor U14936 (N_14936,N_14031,N_14229);
nand U14937 (N_14937,N_13964,N_14391);
and U14938 (N_14938,N_14377,N_13931);
or U14939 (N_14939,N_13981,N_14037);
nand U14940 (N_14940,N_14249,N_14006);
and U14941 (N_14941,N_13806,N_13714);
or U14942 (N_14942,N_14100,N_14124);
and U14943 (N_14943,N_13792,N_14105);
nor U14944 (N_14944,N_13615,N_14199);
and U14945 (N_14945,N_14221,N_13706);
xor U14946 (N_14946,N_14115,N_14336);
and U14947 (N_14947,N_13933,N_13829);
or U14948 (N_14948,N_13978,N_13834);
nor U14949 (N_14949,N_13634,N_13839);
xnor U14950 (N_14950,N_14364,N_14114);
nor U14951 (N_14951,N_13979,N_13616);
or U14952 (N_14952,N_14046,N_13985);
nand U14953 (N_14953,N_14210,N_14169);
xnor U14954 (N_14954,N_13648,N_14340);
nor U14955 (N_14955,N_13784,N_13995);
and U14956 (N_14956,N_13860,N_13939);
nor U14957 (N_14957,N_13838,N_14104);
and U14958 (N_14958,N_13995,N_14064);
xor U14959 (N_14959,N_13796,N_14299);
or U14960 (N_14960,N_13665,N_14269);
and U14961 (N_14961,N_13786,N_14070);
or U14962 (N_14962,N_13610,N_14059);
or U14963 (N_14963,N_14003,N_14294);
nand U14964 (N_14964,N_13952,N_13721);
xnor U14965 (N_14965,N_13874,N_14367);
and U14966 (N_14966,N_14241,N_13751);
nand U14967 (N_14967,N_14264,N_13675);
and U14968 (N_14968,N_13777,N_14191);
and U14969 (N_14969,N_13881,N_13980);
nand U14970 (N_14970,N_13905,N_13847);
and U14971 (N_14971,N_13889,N_14365);
and U14972 (N_14972,N_14064,N_13714);
nand U14973 (N_14973,N_14082,N_13789);
nor U14974 (N_14974,N_14003,N_14141);
xor U14975 (N_14975,N_13614,N_13708);
xor U14976 (N_14976,N_13795,N_14265);
or U14977 (N_14977,N_14266,N_14340);
nand U14978 (N_14978,N_14336,N_14030);
or U14979 (N_14979,N_14361,N_13727);
nand U14980 (N_14980,N_14209,N_14344);
or U14981 (N_14981,N_14347,N_14317);
or U14982 (N_14982,N_13895,N_13796);
nor U14983 (N_14983,N_13619,N_13799);
nand U14984 (N_14984,N_14155,N_13703);
and U14985 (N_14985,N_14366,N_13856);
and U14986 (N_14986,N_14142,N_14253);
and U14987 (N_14987,N_14137,N_13956);
or U14988 (N_14988,N_14098,N_14152);
xnor U14989 (N_14989,N_13810,N_13877);
nand U14990 (N_14990,N_13891,N_13633);
and U14991 (N_14991,N_14164,N_14397);
nand U14992 (N_14992,N_13713,N_14003);
nor U14993 (N_14993,N_14343,N_14392);
nor U14994 (N_14994,N_13691,N_13892);
nand U14995 (N_14995,N_14138,N_14221);
xnor U14996 (N_14996,N_13620,N_13883);
xnor U14997 (N_14997,N_14208,N_13920);
xor U14998 (N_14998,N_13911,N_14285);
xor U14999 (N_14999,N_14175,N_14173);
xnor U15000 (N_15000,N_13805,N_14150);
and U15001 (N_15001,N_13832,N_13888);
or U15002 (N_15002,N_13733,N_14258);
or U15003 (N_15003,N_14375,N_14089);
nor U15004 (N_15004,N_14229,N_13884);
xor U15005 (N_15005,N_14152,N_13938);
nand U15006 (N_15006,N_13613,N_13716);
or U15007 (N_15007,N_14358,N_14036);
nor U15008 (N_15008,N_13913,N_13621);
nor U15009 (N_15009,N_13755,N_13869);
and U15010 (N_15010,N_13845,N_14349);
and U15011 (N_15011,N_14285,N_13669);
or U15012 (N_15012,N_13974,N_14375);
xnor U15013 (N_15013,N_14013,N_14132);
or U15014 (N_15014,N_13821,N_14034);
nand U15015 (N_15015,N_14365,N_14175);
and U15016 (N_15016,N_13701,N_14037);
and U15017 (N_15017,N_14151,N_14087);
or U15018 (N_15018,N_13859,N_13657);
nand U15019 (N_15019,N_14234,N_13918);
nor U15020 (N_15020,N_13899,N_13668);
and U15021 (N_15021,N_14382,N_14307);
nor U15022 (N_15022,N_14388,N_14208);
nor U15023 (N_15023,N_13680,N_14328);
nand U15024 (N_15024,N_13814,N_13630);
xnor U15025 (N_15025,N_14203,N_13863);
and U15026 (N_15026,N_14168,N_14247);
xnor U15027 (N_15027,N_13621,N_13858);
or U15028 (N_15028,N_13954,N_13747);
and U15029 (N_15029,N_14141,N_14305);
xor U15030 (N_15030,N_14112,N_14134);
or U15031 (N_15031,N_13784,N_14061);
or U15032 (N_15032,N_14051,N_13838);
xnor U15033 (N_15033,N_13892,N_13682);
or U15034 (N_15034,N_14303,N_14064);
and U15035 (N_15035,N_13704,N_13810);
nand U15036 (N_15036,N_14314,N_13657);
xnor U15037 (N_15037,N_14351,N_13896);
or U15038 (N_15038,N_14326,N_13990);
or U15039 (N_15039,N_13945,N_14322);
xnor U15040 (N_15040,N_14330,N_14292);
nor U15041 (N_15041,N_14186,N_14202);
xor U15042 (N_15042,N_13722,N_13622);
nor U15043 (N_15043,N_14108,N_14068);
nor U15044 (N_15044,N_14086,N_13962);
and U15045 (N_15045,N_13964,N_13765);
or U15046 (N_15046,N_13997,N_14255);
xnor U15047 (N_15047,N_13995,N_14059);
and U15048 (N_15048,N_14165,N_14146);
and U15049 (N_15049,N_14234,N_13955);
nor U15050 (N_15050,N_13695,N_13721);
or U15051 (N_15051,N_14008,N_14241);
xnor U15052 (N_15052,N_14021,N_14243);
and U15053 (N_15053,N_14132,N_13647);
or U15054 (N_15054,N_14119,N_14387);
and U15055 (N_15055,N_13703,N_13648);
nand U15056 (N_15056,N_13711,N_14109);
or U15057 (N_15057,N_13744,N_13926);
or U15058 (N_15058,N_13720,N_14176);
and U15059 (N_15059,N_14364,N_14073);
nand U15060 (N_15060,N_14337,N_14383);
and U15061 (N_15061,N_14370,N_14338);
or U15062 (N_15062,N_14085,N_14383);
or U15063 (N_15063,N_13989,N_14306);
and U15064 (N_15064,N_13799,N_14100);
and U15065 (N_15065,N_14317,N_13742);
nor U15066 (N_15066,N_14345,N_13789);
or U15067 (N_15067,N_13943,N_13878);
xnor U15068 (N_15068,N_14296,N_14022);
or U15069 (N_15069,N_13624,N_13790);
nor U15070 (N_15070,N_14084,N_13839);
nor U15071 (N_15071,N_13988,N_14370);
and U15072 (N_15072,N_13699,N_13990);
xor U15073 (N_15073,N_14295,N_14012);
nand U15074 (N_15074,N_13961,N_13895);
and U15075 (N_15075,N_13836,N_13752);
or U15076 (N_15076,N_14109,N_14261);
xor U15077 (N_15077,N_14334,N_14311);
nor U15078 (N_15078,N_13676,N_13729);
nand U15079 (N_15079,N_13977,N_14298);
and U15080 (N_15080,N_13619,N_14333);
nor U15081 (N_15081,N_13668,N_14049);
and U15082 (N_15082,N_14034,N_14306);
or U15083 (N_15083,N_14105,N_14304);
xnor U15084 (N_15084,N_14359,N_13962);
and U15085 (N_15085,N_13845,N_13688);
and U15086 (N_15086,N_13969,N_13676);
and U15087 (N_15087,N_13753,N_14224);
and U15088 (N_15088,N_13877,N_13796);
or U15089 (N_15089,N_14342,N_13682);
xnor U15090 (N_15090,N_14140,N_13605);
nand U15091 (N_15091,N_13717,N_13703);
or U15092 (N_15092,N_13744,N_13954);
nand U15093 (N_15093,N_14127,N_13682);
or U15094 (N_15094,N_13798,N_14395);
nor U15095 (N_15095,N_13981,N_14204);
xnor U15096 (N_15096,N_14064,N_13721);
and U15097 (N_15097,N_14050,N_13707);
xnor U15098 (N_15098,N_13666,N_13722);
nor U15099 (N_15099,N_14243,N_14375);
nand U15100 (N_15100,N_13650,N_14360);
nand U15101 (N_15101,N_13796,N_14292);
nor U15102 (N_15102,N_13624,N_14227);
and U15103 (N_15103,N_13817,N_14299);
xor U15104 (N_15104,N_14366,N_14183);
nor U15105 (N_15105,N_14290,N_13938);
nor U15106 (N_15106,N_14035,N_13671);
xnor U15107 (N_15107,N_13871,N_14132);
or U15108 (N_15108,N_13763,N_14228);
or U15109 (N_15109,N_14151,N_13642);
xor U15110 (N_15110,N_14101,N_14020);
nand U15111 (N_15111,N_14143,N_13686);
xor U15112 (N_15112,N_14010,N_14359);
xor U15113 (N_15113,N_14148,N_13731);
and U15114 (N_15114,N_13904,N_14151);
xnor U15115 (N_15115,N_14313,N_13650);
or U15116 (N_15116,N_13667,N_13753);
nor U15117 (N_15117,N_14325,N_13968);
nor U15118 (N_15118,N_14071,N_14149);
nor U15119 (N_15119,N_14349,N_13618);
xnor U15120 (N_15120,N_13673,N_14113);
and U15121 (N_15121,N_14131,N_14089);
xnor U15122 (N_15122,N_13671,N_14130);
nand U15123 (N_15123,N_13896,N_14261);
nor U15124 (N_15124,N_13875,N_14214);
and U15125 (N_15125,N_14177,N_14302);
or U15126 (N_15126,N_14127,N_13705);
and U15127 (N_15127,N_14222,N_14242);
or U15128 (N_15128,N_13976,N_13974);
xor U15129 (N_15129,N_13766,N_13808);
and U15130 (N_15130,N_13669,N_14373);
nand U15131 (N_15131,N_14209,N_13739);
nor U15132 (N_15132,N_13927,N_14244);
and U15133 (N_15133,N_14117,N_13757);
nor U15134 (N_15134,N_13917,N_14041);
or U15135 (N_15135,N_14069,N_13817);
xor U15136 (N_15136,N_14161,N_13750);
xnor U15137 (N_15137,N_14306,N_14105);
xnor U15138 (N_15138,N_13835,N_13886);
and U15139 (N_15139,N_14378,N_14123);
xnor U15140 (N_15140,N_13958,N_14026);
and U15141 (N_15141,N_14018,N_13935);
or U15142 (N_15142,N_13762,N_13993);
nor U15143 (N_15143,N_13717,N_13985);
or U15144 (N_15144,N_13755,N_14362);
or U15145 (N_15145,N_13961,N_13661);
xor U15146 (N_15146,N_14277,N_13849);
or U15147 (N_15147,N_14034,N_13616);
or U15148 (N_15148,N_13852,N_14133);
nand U15149 (N_15149,N_14167,N_13762);
or U15150 (N_15150,N_13639,N_14305);
and U15151 (N_15151,N_13933,N_13951);
or U15152 (N_15152,N_14224,N_13602);
nand U15153 (N_15153,N_14037,N_14159);
nor U15154 (N_15154,N_14048,N_13818);
xnor U15155 (N_15155,N_13701,N_13824);
nor U15156 (N_15156,N_14207,N_13821);
nor U15157 (N_15157,N_14233,N_14356);
or U15158 (N_15158,N_14260,N_14161);
or U15159 (N_15159,N_14173,N_13808);
nor U15160 (N_15160,N_14178,N_13676);
nor U15161 (N_15161,N_14150,N_14004);
nand U15162 (N_15162,N_14388,N_14186);
and U15163 (N_15163,N_13875,N_14280);
nor U15164 (N_15164,N_13795,N_13668);
or U15165 (N_15165,N_14182,N_14349);
and U15166 (N_15166,N_13938,N_14063);
xnor U15167 (N_15167,N_14302,N_13698);
nor U15168 (N_15168,N_14049,N_13691);
xnor U15169 (N_15169,N_13732,N_14013);
and U15170 (N_15170,N_14244,N_14324);
nor U15171 (N_15171,N_13669,N_13771);
nand U15172 (N_15172,N_13928,N_13961);
xor U15173 (N_15173,N_13985,N_14145);
and U15174 (N_15174,N_13920,N_13864);
nor U15175 (N_15175,N_13842,N_14228);
and U15176 (N_15176,N_13735,N_14078);
xnor U15177 (N_15177,N_13701,N_13833);
nor U15178 (N_15178,N_13961,N_13946);
nor U15179 (N_15179,N_14308,N_14037);
nor U15180 (N_15180,N_14180,N_14070);
and U15181 (N_15181,N_13773,N_13607);
nor U15182 (N_15182,N_14201,N_14372);
nand U15183 (N_15183,N_14299,N_14027);
nand U15184 (N_15184,N_13973,N_13608);
or U15185 (N_15185,N_14247,N_14375);
nor U15186 (N_15186,N_14155,N_14391);
nor U15187 (N_15187,N_14144,N_13626);
or U15188 (N_15188,N_14364,N_14212);
nand U15189 (N_15189,N_13700,N_13687);
nand U15190 (N_15190,N_13712,N_13972);
and U15191 (N_15191,N_14383,N_13710);
or U15192 (N_15192,N_13684,N_13991);
xnor U15193 (N_15193,N_13944,N_13993);
nand U15194 (N_15194,N_14009,N_14053);
and U15195 (N_15195,N_14363,N_14294);
nor U15196 (N_15196,N_14033,N_13794);
or U15197 (N_15197,N_13685,N_13956);
xnor U15198 (N_15198,N_14279,N_13835);
or U15199 (N_15199,N_13766,N_14214);
nor U15200 (N_15200,N_14816,N_15049);
xnor U15201 (N_15201,N_14541,N_14763);
nand U15202 (N_15202,N_14943,N_14612);
nand U15203 (N_15203,N_14966,N_15160);
nand U15204 (N_15204,N_14674,N_15040);
or U15205 (N_15205,N_14592,N_15041);
and U15206 (N_15206,N_14620,N_14506);
or U15207 (N_15207,N_14748,N_14964);
xor U15208 (N_15208,N_14536,N_14431);
nand U15209 (N_15209,N_15078,N_14540);
or U15210 (N_15210,N_14512,N_15023);
xor U15211 (N_15211,N_14433,N_14835);
nor U15212 (N_15212,N_15019,N_15178);
or U15213 (N_15213,N_14971,N_15053);
and U15214 (N_15214,N_14455,N_14430);
and U15215 (N_15215,N_14581,N_14962);
nand U15216 (N_15216,N_15082,N_14852);
and U15217 (N_15217,N_14693,N_15180);
xnor U15218 (N_15218,N_14917,N_14619);
xor U15219 (N_15219,N_14798,N_14869);
and U15220 (N_15220,N_15163,N_15139);
nor U15221 (N_15221,N_14965,N_15034);
or U15222 (N_15222,N_14696,N_15105);
nand U15223 (N_15223,N_14569,N_14783);
nand U15224 (N_15224,N_15001,N_15072);
and U15225 (N_15225,N_14854,N_14484);
or U15226 (N_15226,N_14858,N_15156);
and U15227 (N_15227,N_14597,N_15027);
or U15228 (N_15228,N_15002,N_14605);
and U15229 (N_15229,N_14575,N_14675);
nand U15230 (N_15230,N_14772,N_14863);
xor U15231 (N_15231,N_14522,N_14519);
or U15232 (N_15232,N_14654,N_14504);
nand U15233 (N_15233,N_15007,N_14641);
nor U15234 (N_15234,N_14649,N_14400);
and U15235 (N_15235,N_14749,N_14880);
nor U15236 (N_15236,N_14588,N_14846);
nand U15237 (N_15237,N_14981,N_14628);
or U15238 (N_15238,N_14711,N_15145);
nor U15239 (N_15239,N_15080,N_14870);
nor U15240 (N_15240,N_14771,N_14834);
and U15241 (N_15241,N_15020,N_14655);
or U15242 (N_15242,N_14785,N_15127);
xnor U15243 (N_15243,N_14664,N_14411);
and U15244 (N_15244,N_14514,N_14872);
and U15245 (N_15245,N_15032,N_15021);
nor U15246 (N_15246,N_14570,N_14937);
nor U15247 (N_15247,N_14809,N_15169);
nand U15248 (N_15248,N_14996,N_14599);
and U15249 (N_15249,N_14474,N_14551);
or U15250 (N_15250,N_14545,N_15195);
and U15251 (N_15251,N_14889,N_14409);
or U15252 (N_15252,N_15097,N_14583);
nor U15253 (N_15253,N_14482,N_14756);
nand U15254 (N_15254,N_14670,N_14652);
xnor U15255 (N_15255,N_14796,N_14960);
nand U15256 (N_15256,N_14938,N_14918);
or U15257 (N_15257,N_14446,N_14955);
nand U15258 (N_15258,N_14893,N_14841);
nand U15259 (N_15259,N_14924,N_14751);
nor U15260 (N_15260,N_14804,N_14891);
or U15261 (N_15261,N_14406,N_14611);
nand U15262 (N_15262,N_14580,N_14546);
or U15263 (N_15263,N_15181,N_14959);
xor U15264 (N_15264,N_14704,N_14420);
or U15265 (N_15265,N_14454,N_14689);
xnor U15266 (N_15266,N_14470,N_14805);
and U15267 (N_15267,N_14615,N_14463);
or U15268 (N_15268,N_14525,N_14571);
nor U15269 (N_15269,N_15029,N_15164);
xnor U15270 (N_15270,N_14833,N_15043);
nor U15271 (N_15271,N_14505,N_14839);
nor U15272 (N_15272,N_14444,N_14699);
nand U15273 (N_15273,N_14625,N_14626);
nor U15274 (N_15274,N_14990,N_15150);
nand U15275 (N_15275,N_14587,N_15179);
or U15276 (N_15276,N_14537,N_14538);
xor U15277 (N_15277,N_14478,N_15106);
or U15278 (N_15278,N_14912,N_15135);
and U15279 (N_15279,N_14521,N_14553);
nand U15280 (N_15280,N_14679,N_14946);
xor U15281 (N_15281,N_14866,N_15119);
nand U15282 (N_15282,N_15187,N_14415);
nor U15283 (N_15283,N_14426,N_15152);
nor U15284 (N_15284,N_14424,N_14413);
or U15285 (N_15285,N_14567,N_14493);
nand U15286 (N_15286,N_14983,N_15052);
and U15287 (N_15287,N_14724,N_14606);
nor U15288 (N_15288,N_14826,N_14973);
nor U15289 (N_15289,N_15120,N_14665);
and U15290 (N_15290,N_14890,N_15044);
nor U15291 (N_15291,N_14837,N_14766);
nor U15292 (N_15292,N_14781,N_14705);
or U15293 (N_15293,N_14726,N_14523);
xnor U15294 (N_15294,N_14779,N_14487);
xnor U15295 (N_15295,N_14584,N_15109);
and U15296 (N_15296,N_14448,N_14673);
and U15297 (N_15297,N_15062,N_14987);
nor U15298 (N_15298,N_14671,N_15175);
or U15299 (N_15299,N_14860,N_15189);
nor U15300 (N_15300,N_14476,N_14800);
xor U15301 (N_15301,N_14878,N_14643);
nand U15302 (N_15302,N_14862,N_14857);
nand U15303 (N_15303,N_15108,N_15048);
or U15304 (N_15304,N_15026,N_14657);
nor U15305 (N_15305,N_14988,N_14819);
nand U15306 (N_15306,N_14640,N_14492);
xnor U15307 (N_15307,N_14886,N_14591);
nor U15308 (N_15308,N_15129,N_14718);
nand U15309 (N_15309,N_14761,N_14667);
nand U15310 (N_15310,N_15148,N_14466);
or U15311 (N_15311,N_14830,N_14593);
or U15312 (N_15312,N_14725,N_14443);
or U15313 (N_15313,N_15154,N_15077);
xnor U15314 (N_15314,N_14635,N_15098);
or U15315 (N_15315,N_14995,N_15193);
xor U15316 (N_15316,N_14520,N_14922);
or U15317 (N_15317,N_14694,N_14452);
nand U15318 (N_15318,N_14982,N_14622);
and U15319 (N_15319,N_14797,N_14709);
nor U15320 (N_15320,N_14661,N_14842);
xor U15321 (N_15321,N_14740,N_15143);
xor U15322 (N_15322,N_14980,N_14552);
nor U15323 (N_15323,N_15166,N_14867);
nand U15324 (N_15324,N_14914,N_14483);
xor U15325 (N_15325,N_15137,N_15070);
xor U15326 (N_15326,N_14945,N_14490);
nor U15327 (N_15327,N_14876,N_15167);
nand U15328 (N_15328,N_14548,N_14408);
nor U15329 (N_15329,N_14712,N_14594);
xor U15330 (N_15330,N_14480,N_14404);
nor U15331 (N_15331,N_14610,N_14840);
nand U15332 (N_15332,N_15064,N_14488);
or U15333 (N_15333,N_15037,N_14682);
and U15334 (N_15334,N_14813,N_14698);
or U15335 (N_15335,N_14510,N_15117);
nor U15336 (N_15336,N_14423,N_15196);
nand U15337 (N_15337,N_15018,N_14873);
nand U15338 (N_15338,N_14678,N_14899);
nor U15339 (N_15339,N_14562,N_14818);
and U15340 (N_15340,N_14629,N_14847);
or U15341 (N_15341,N_14631,N_14774);
or U15342 (N_15342,N_14735,N_14907);
nor U15343 (N_15343,N_14624,N_15199);
nor U15344 (N_15344,N_14767,N_14757);
and U15345 (N_15345,N_15121,N_15184);
and U15346 (N_15346,N_14515,N_14422);
and U15347 (N_15347,N_15146,N_14403);
nand U15348 (N_15348,N_14472,N_14456);
nand U15349 (N_15349,N_14992,N_14642);
or U15350 (N_15350,N_15118,N_14926);
nor U15351 (N_15351,N_14638,N_14730);
xnor U15352 (N_15352,N_14741,N_14934);
xor U15353 (N_15353,N_14770,N_15000);
and U15354 (N_15354,N_14604,N_15115);
xor U15355 (N_15355,N_15107,N_14526);
nor U15356 (N_15356,N_14658,N_14687);
nand U15357 (N_15357,N_14586,N_14829);
and U15358 (N_15358,N_15005,N_14572);
nor U15359 (N_15359,N_14941,N_15074);
or U15360 (N_15360,N_14904,N_15094);
xor U15361 (N_15361,N_14820,N_14888);
or U15362 (N_15362,N_14453,N_15095);
nor U15363 (N_15363,N_15004,N_15177);
nor U15364 (N_15364,N_15036,N_14887);
and U15365 (N_15365,N_14963,N_15051);
and U15366 (N_15366,N_14630,N_14823);
nor U15367 (N_15367,N_14634,N_14877);
nor U15368 (N_15368,N_14511,N_14432);
nand U15369 (N_15369,N_14951,N_14760);
and U15370 (N_15370,N_15073,N_14776);
xnor U15371 (N_15371,N_14777,N_15066);
nand U15372 (N_15372,N_14738,N_14977);
xor U15373 (N_15373,N_14864,N_14745);
nand U15374 (N_15374,N_14848,N_14688);
nand U15375 (N_15375,N_15054,N_15176);
xnor U15376 (N_15376,N_14831,N_14817);
or U15377 (N_15377,N_15087,N_14722);
or U15378 (N_15378,N_15188,N_14539);
nor U15379 (N_15379,N_14464,N_14849);
or U15380 (N_15380,N_14533,N_15083);
xor U15381 (N_15381,N_14916,N_15192);
xnor U15382 (N_15382,N_14669,N_15183);
or U15383 (N_15383,N_14542,N_14425);
xor U15384 (N_15384,N_14556,N_14547);
nand U15385 (N_15385,N_14677,N_15168);
or U15386 (N_15386,N_14659,N_15136);
nand U15387 (N_15387,N_14952,N_15045);
and U15388 (N_15388,N_14434,N_14884);
and U15389 (N_15389,N_14746,N_14923);
nand U15390 (N_15390,N_15068,N_14903);
or U15391 (N_15391,N_14499,N_14949);
xor U15392 (N_15392,N_14419,N_14529);
nor U15393 (N_15393,N_14498,N_14407);
or U15394 (N_15394,N_15050,N_15033);
nor U15395 (N_15395,N_15092,N_14868);
or U15396 (N_15396,N_14421,N_15096);
nor U15397 (N_15397,N_15017,N_14913);
and U15398 (N_15398,N_14879,N_15038);
xnor U15399 (N_15399,N_15059,N_14824);
nand U15400 (N_15400,N_14577,N_14944);
nor U15401 (N_15401,N_14574,N_15161);
and U15402 (N_15402,N_15102,N_14660);
or U15403 (N_15403,N_14460,N_15142);
nand U15404 (N_15404,N_14734,N_14729);
xnor U15405 (N_15405,N_14639,N_14700);
xor U15406 (N_15406,N_15147,N_14998);
nor U15407 (N_15407,N_15065,N_15099);
nand U15408 (N_15408,N_14897,N_14750);
xnor U15409 (N_15409,N_14695,N_14645);
nand U15410 (N_15410,N_15112,N_15123);
or U15411 (N_15411,N_14778,N_14601);
xor U15412 (N_15412,N_14573,N_14845);
nor U15413 (N_15413,N_14691,N_14978);
and U15414 (N_15414,N_14794,N_14475);
or U15415 (N_15415,N_14439,N_14672);
nand U15416 (N_15416,N_14811,N_15130);
or U15417 (N_15417,N_14881,N_14975);
nor U15418 (N_15418,N_14765,N_14617);
and U15419 (N_15419,N_15028,N_14494);
and U15420 (N_15420,N_14663,N_15170);
and U15421 (N_15421,N_15194,N_15159);
or U15422 (N_15422,N_14892,N_14559);
nor U15423 (N_15423,N_14939,N_14662);
or U15424 (N_15424,N_14527,N_14441);
xor U15425 (N_15425,N_14458,N_14558);
xnor U15426 (N_15426,N_14752,N_15006);
and U15427 (N_15427,N_15174,N_14933);
nand U15428 (N_15428,N_14530,N_15090);
xnor U15429 (N_15429,N_14827,N_14736);
or U15430 (N_15430,N_14560,N_15113);
xnor U15431 (N_15431,N_14467,N_15014);
nor U15432 (N_15432,N_14717,N_14788);
nor U15433 (N_15433,N_14782,N_14927);
nand U15434 (N_15434,N_15197,N_15063);
nand U15435 (N_15435,N_15009,N_14618);
nor U15436 (N_15436,N_14865,N_14633);
or U15437 (N_15437,N_14993,N_14485);
and U15438 (N_15438,N_14859,N_15010);
and U15439 (N_15439,N_14600,N_14609);
or U15440 (N_15440,N_14703,N_14557);
nor U15441 (N_15441,N_14684,N_14497);
or U15442 (N_15442,N_14759,N_14753);
nand U15443 (N_15443,N_15151,N_14896);
xnor U15444 (N_15444,N_14871,N_15056);
nand U15445 (N_15445,N_14555,N_14412);
nand U15446 (N_15446,N_14970,N_14532);
nand U15447 (N_15447,N_14808,N_14825);
xnor U15448 (N_15448,N_15190,N_14416);
xnor U15449 (N_15449,N_14936,N_15016);
and U15450 (N_15450,N_14795,N_15081);
xor U15451 (N_15451,N_14435,N_14731);
xnor U15452 (N_15452,N_14803,N_14895);
nand U15453 (N_15453,N_14815,N_14994);
xor U15454 (N_15454,N_14517,N_14481);
and U15455 (N_15455,N_14784,N_14989);
and U15456 (N_15456,N_14564,N_14690);
xor U15457 (N_15457,N_14961,N_14681);
xor U15458 (N_15458,N_14405,N_14534);
or U15459 (N_15459,N_14554,N_14744);
nand U15460 (N_15460,N_14898,N_14549);
nor U15461 (N_15461,N_14999,N_15132);
and U15462 (N_15462,N_14683,N_14780);
and U15463 (N_15463,N_15058,N_14787);
nor U15464 (N_15464,N_14758,N_14501);
xnor U15465 (N_15465,N_14828,N_15182);
or U15466 (N_15466,N_15055,N_14449);
or U15467 (N_15467,N_14940,N_14883);
and U15468 (N_15468,N_14733,N_14650);
nor U15469 (N_15469,N_14968,N_14942);
or U15470 (N_15470,N_14802,N_15111);
nand U15471 (N_15471,N_14468,N_14616);
xor U15472 (N_15472,N_14921,N_14747);
and U15473 (N_15473,N_14838,N_14929);
nor U15474 (N_15474,N_14732,N_14462);
nand U15475 (N_15475,N_15046,N_14894);
and U15476 (N_15476,N_14810,N_14656);
or U15477 (N_15477,N_14953,N_15125);
nor U15478 (N_15478,N_14856,N_14590);
xor U15479 (N_15479,N_14428,N_15061);
nand U15480 (N_15480,N_15124,N_14653);
xor U15481 (N_15481,N_14632,N_14598);
nor U15482 (N_15482,N_14762,N_14874);
or U15483 (N_15483,N_14806,N_14603);
or U15484 (N_15484,N_15071,N_15134);
and U15485 (N_15485,N_14507,N_14489);
nand U15486 (N_15486,N_14822,N_14902);
nand U15487 (N_15487,N_15079,N_14595);
nand U15488 (N_15488,N_14773,N_15128);
nand U15489 (N_15489,N_14930,N_14972);
xor U15490 (N_15490,N_14928,N_14568);
nor U15491 (N_15491,N_14710,N_15089);
nor U15492 (N_15492,N_14754,N_14666);
and U15493 (N_15493,N_14651,N_14985);
or U15494 (N_15494,N_14925,N_14582);
xnor U15495 (N_15495,N_15126,N_14801);
nor U15496 (N_15496,N_14438,N_14607);
and U15497 (N_15497,N_14566,N_15057);
nor U15498 (N_15498,N_14967,N_14769);
xnor U15499 (N_15499,N_14613,N_14440);
xor U15500 (N_15500,N_15012,N_14701);
nand U15501 (N_15501,N_14550,N_15022);
and U15502 (N_15502,N_14637,N_14812);
nor U15503 (N_15503,N_14958,N_14799);
nor U15504 (N_15504,N_14791,N_14821);
nor U15505 (N_15505,N_14543,N_14720);
nand U15506 (N_15506,N_15131,N_15008);
nor U15507 (N_15507,N_14727,N_14589);
nor U15508 (N_15508,N_14451,N_15086);
or U15509 (N_15509,N_14561,N_14565);
nand U15510 (N_15510,N_14851,N_15093);
or U15511 (N_15511,N_14450,N_15060);
nand U15512 (N_15512,N_15069,N_14855);
or U15513 (N_15513,N_15138,N_14714);
and U15514 (N_15514,N_15173,N_14457);
nand U15515 (N_15515,N_14513,N_14844);
nand U15516 (N_15516,N_14427,N_15133);
nand U15517 (N_15517,N_14447,N_15171);
nor U15518 (N_15518,N_14986,N_14882);
and U15519 (N_15519,N_15084,N_14644);
xnor U15520 (N_15520,N_14459,N_15155);
or U15521 (N_15521,N_14909,N_14491);
or U15522 (N_15522,N_14728,N_14739);
xor U15523 (N_15523,N_15110,N_14585);
or U15524 (N_15524,N_15101,N_14685);
and U15525 (N_15525,N_14706,N_14518);
or U15526 (N_15526,N_15165,N_14436);
and U15527 (N_15527,N_14713,N_15162);
nor U15528 (N_15528,N_14954,N_14647);
or U15529 (N_15529,N_14920,N_14715);
nor U15530 (N_15530,N_14680,N_14935);
nand U15531 (N_15531,N_14905,N_15085);
nand U15532 (N_15532,N_14742,N_15157);
nor U15533 (N_15533,N_14578,N_15141);
nand U15534 (N_15534,N_14947,N_14401);
nand U15535 (N_15535,N_15191,N_14814);
and U15536 (N_15536,N_14509,N_14418);
and U15537 (N_15537,N_14836,N_14768);
or U15538 (N_15538,N_14911,N_14906);
and U15539 (N_15539,N_14417,N_15042);
nor U15540 (N_15540,N_15088,N_14477);
nand U15541 (N_15541,N_14429,N_14861);
or U15542 (N_15542,N_14979,N_14402);
and U15543 (N_15543,N_14479,N_15103);
nor U15544 (N_15544,N_14764,N_14465);
nand U15545 (N_15545,N_14576,N_14496);
nor U15546 (N_15546,N_14535,N_14516);
nand U15547 (N_15547,N_15076,N_14948);
and U15548 (N_15548,N_15114,N_14807);
nand U15549 (N_15549,N_14931,N_14414);
nand U15550 (N_15550,N_14686,N_15011);
or U15551 (N_15551,N_14708,N_14502);
or U15552 (N_15552,N_15144,N_15047);
xor U15553 (N_15553,N_15104,N_14910);
and U15554 (N_15554,N_14528,N_14792);
xnor U15555 (N_15555,N_14900,N_14721);
and U15556 (N_15556,N_14793,N_15031);
nand U15557 (N_15557,N_14697,N_15067);
xor U15558 (N_15558,N_14716,N_15015);
and U15559 (N_15559,N_14885,N_14843);
nor U15560 (N_15560,N_14563,N_14850);
and U15561 (N_15561,N_14410,N_15039);
and U15562 (N_15562,N_14719,N_14950);
xnor U15563 (N_15563,N_14832,N_14997);
or U15564 (N_15564,N_14853,N_15100);
nand U15565 (N_15565,N_14908,N_14743);
xnor U15566 (N_15566,N_14627,N_14636);
or U15567 (N_15567,N_14707,N_15153);
or U15568 (N_15568,N_14442,N_15186);
nor U15569 (N_15569,N_15122,N_14919);
xor U15570 (N_15570,N_14969,N_14676);
nor U15571 (N_15571,N_14957,N_14445);
nor U15572 (N_15572,N_14579,N_14991);
or U15573 (N_15573,N_14471,N_14495);
nor U15574 (N_15574,N_14976,N_14469);
xnor U15575 (N_15575,N_15149,N_15158);
or U15576 (N_15576,N_14614,N_15035);
nand U15577 (N_15577,N_15172,N_14602);
nor U15578 (N_15578,N_15003,N_14596);
and U15579 (N_15579,N_15116,N_15030);
nor U15580 (N_15580,N_14692,N_14503);
nor U15581 (N_15581,N_14646,N_15024);
or U15582 (N_15582,N_15185,N_14723);
and U15583 (N_15583,N_14915,N_14544);
and U15584 (N_15584,N_14755,N_15198);
or U15585 (N_15585,N_14500,N_14524);
and U15586 (N_15586,N_14473,N_14775);
xor U15587 (N_15587,N_14668,N_15091);
xor U15588 (N_15588,N_15075,N_14437);
xor U15589 (N_15589,N_15025,N_14786);
nor U15590 (N_15590,N_14621,N_14956);
nor U15591 (N_15591,N_14901,N_14702);
nand U15592 (N_15592,N_14984,N_14932);
nand U15593 (N_15593,N_14508,N_14648);
or U15594 (N_15594,N_14486,N_15013);
xnor U15595 (N_15595,N_14974,N_14737);
nand U15596 (N_15596,N_14461,N_14790);
or U15597 (N_15597,N_14608,N_14875);
nand U15598 (N_15598,N_14531,N_14623);
and U15599 (N_15599,N_15140,N_14789);
nand U15600 (N_15600,N_14881,N_14589);
xnor U15601 (N_15601,N_14599,N_14977);
nor U15602 (N_15602,N_14944,N_14515);
nand U15603 (N_15603,N_15198,N_14856);
or U15604 (N_15604,N_14782,N_14957);
nor U15605 (N_15605,N_14952,N_15115);
nor U15606 (N_15606,N_15019,N_15173);
or U15607 (N_15607,N_14822,N_15145);
and U15608 (N_15608,N_14617,N_14796);
and U15609 (N_15609,N_15068,N_14500);
or U15610 (N_15610,N_14959,N_15030);
nor U15611 (N_15611,N_15126,N_14624);
nand U15612 (N_15612,N_14859,N_14469);
nand U15613 (N_15613,N_14595,N_15053);
xor U15614 (N_15614,N_14636,N_15121);
nand U15615 (N_15615,N_14634,N_14970);
or U15616 (N_15616,N_14799,N_14730);
nand U15617 (N_15617,N_14756,N_14882);
or U15618 (N_15618,N_15124,N_14596);
or U15619 (N_15619,N_15157,N_14573);
xor U15620 (N_15620,N_15160,N_14548);
nand U15621 (N_15621,N_15067,N_14984);
or U15622 (N_15622,N_15164,N_14927);
nand U15623 (N_15623,N_15150,N_14782);
nor U15624 (N_15624,N_14630,N_14442);
nor U15625 (N_15625,N_14742,N_15160);
nand U15626 (N_15626,N_14954,N_15110);
and U15627 (N_15627,N_14987,N_14848);
nor U15628 (N_15628,N_15001,N_15148);
nor U15629 (N_15629,N_14708,N_15164);
nand U15630 (N_15630,N_14663,N_15066);
and U15631 (N_15631,N_14509,N_15079);
nand U15632 (N_15632,N_14842,N_14617);
xor U15633 (N_15633,N_15171,N_14584);
and U15634 (N_15634,N_14536,N_15103);
nand U15635 (N_15635,N_15132,N_14408);
nand U15636 (N_15636,N_14899,N_15039);
xor U15637 (N_15637,N_14747,N_14408);
or U15638 (N_15638,N_15086,N_15055);
xor U15639 (N_15639,N_15001,N_15175);
xnor U15640 (N_15640,N_15071,N_14817);
xnor U15641 (N_15641,N_14986,N_14592);
or U15642 (N_15642,N_14693,N_15193);
nor U15643 (N_15643,N_14660,N_14944);
or U15644 (N_15644,N_15146,N_14638);
or U15645 (N_15645,N_14792,N_14403);
nor U15646 (N_15646,N_15074,N_14593);
nand U15647 (N_15647,N_14722,N_14979);
nor U15648 (N_15648,N_14747,N_14564);
xor U15649 (N_15649,N_15170,N_14632);
and U15650 (N_15650,N_14600,N_14719);
and U15651 (N_15651,N_14916,N_14628);
nand U15652 (N_15652,N_15122,N_14657);
nor U15653 (N_15653,N_14805,N_15167);
nor U15654 (N_15654,N_14619,N_14402);
or U15655 (N_15655,N_15075,N_14681);
nand U15656 (N_15656,N_14686,N_14975);
or U15657 (N_15657,N_15182,N_15070);
and U15658 (N_15658,N_15181,N_14634);
nand U15659 (N_15659,N_14463,N_14569);
or U15660 (N_15660,N_14985,N_14425);
or U15661 (N_15661,N_14984,N_15016);
or U15662 (N_15662,N_14878,N_14813);
xor U15663 (N_15663,N_14512,N_15097);
and U15664 (N_15664,N_14602,N_14935);
nor U15665 (N_15665,N_14418,N_15075);
xor U15666 (N_15666,N_15198,N_14458);
nand U15667 (N_15667,N_14888,N_15115);
or U15668 (N_15668,N_15127,N_14405);
or U15669 (N_15669,N_14604,N_14811);
nor U15670 (N_15670,N_14798,N_14654);
xnor U15671 (N_15671,N_15171,N_14466);
nor U15672 (N_15672,N_14607,N_15149);
nor U15673 (N_15673,N_14992,N_14562);
xor U15674 (N_15674,N_14893,N_14674);
nor U15675 (N_15675,N_14969,N_14839);
and U15676 (N_15676,N_14870,N_14752);
and U15677 (N_15677,N_14896,N_15022);
nand U15678 (N_15678,N_14853,N_14532);
and U15679 (N_15679,N_14811,N_14801);
xor U15680 (N_15680,N_14990,N_14600);
or U15681 (N_15681,N_14852,N_15146);
or U15682 (N_15682,N_14499,N_14488);
or U15683 (N_15683,N_14906,N_14942);
xnor U15684 (N_15684,N_14983,N_15043);
nor U15685 (N_15685,N_14709,N_14690);
and U15686 (N_15686,N_14414,N_14585);
xor U15687 (N_15687,N_14588,N_14447);
or U15688 (N_15688,N_15154,N_14426);
and U15689 (N_15689,N_14857,N_14777);
nor U15690 (N_15690,N_14506,N_14644);
nand U15691 (N_15691,N_14681,N_15041);
nor U15692 (N_15692,N_14501,N_15098);
or U15693 (N_15693,N_14955,N_15070);
nand U15694 (N_15694,N_14658,N_15179);
xor U15695 (N_15695,N_14602,N_14731);
or U15696 (N_15696,N_14499,N_14648);
nor U15697 (N_15697,N_14868,N_15027);
or U15698 (N_15698,N_14581,N_15056);
or U15699 (N_15699,N_15127,N_14730);
or U15700 (N_15700,N_15138,N_14543);
and U15701 (N_15701,N_14766,N_14486);
nor U15702 (N_15702,N_14789,N_14609);
and U15703 (N_15703,N_14587,N_14415);
nor U15704 (N_15704,N_15088,N_15037);
xnor U15705 (N_15705,N_14537,N_14660);
nand U15706 (N_15706,N_14874,N_14991);
nor U15707 (N_15707,N_15038,N_15147);
and U15708 (N_15708,N_14872,N_14775);
xnor U15709 (N_15709,N_14800,N_14428);
nor U15710 (N_15710,N_14915,N_14530);
and U15711 (N_15711,N_15097,N_14588);
nor U15712 (N_15712,N_14488,N_14884);
or U15713 (N_15713,N_14778,N_14554);
nor U15714 (N_15714,N_14980,N_14953);
or U15715 (N_15715,N_15131,N_15083);
xnor U15716 (N_15716,N_14419,N_14832);
xor U15717 (N_15717,N_14925,N_14723);
or U15718 (N_15718,N_14417,N_15040);
nand U15719 (N_15719,N_14622,N_14454);
nor U15720 (N_15720,N_14696,N_14645);
nand U15721 (N_15721,N_14607,N_15091);
and U15722 (N_15722,N_14700,N_14485);
nand U15723 (N_15723,N_15180,N_15061);
nor U15724 (N_15724,N_15173,N_14819);
or U15725 (N_15725,N_14697,N_14864);
or U15726 (N_15726,N_14581,N_14738);
xor U15727 (N_15727,N_14575,N_14674);
xnor U15728 (N_15728,N_15126,N_14941);
nor U15729 (N_15729,N_14533,N_14936);
xnor U15730 (N_15730,N_14731,N_14441);
nor U15731 (N_15731,N_14882,N_14557);
and U15732 (N_15732,N_14821,N_15146);
nand U15733 (N_15733,N_14493,N_15118);
nor U15734 (N_15734,N_14795,N_14758);
nor U15735 (N_15735,N_14983,N_14687);
nand U15736 (N_15736,N_14925,N_15169);
nand U15737 (N_15737,N_14692,N_14741);
nor U15738 (N_15738,N_14770,N_14900);
and U15739 (N_15739,N_15151,N_14560);
nand U15740 (N_15740,N_14636,N_15188);
xor U15741 (N_15741,N_14679,N_14400);
xnor U15742 (N_15742,N_14894,N_14651);
and U15743 (N_15743,N_15085,N_14584);
nand U15744 (N_15744,N_14900,N_14500);
nor U15745 (N_15745,N_14943,N_14768);
nor U15746 (N_15746,N_15135,N_14461);
or U15747 (N_15747,N_15050,N_15167);
xnor U15748 (N_15748,N_14527,N_14670);
or U15749 (N_15749,N_14732,N_14632);
and U15750 (N_15750,N_14889,N_14588);
xnor U15751 (N_15751,N_14535,N_14853);
xnor U15752 (N_15752,N_15039,N_14740);
and U15753 (N_15753,N_14994,N_14584);
nor U15754 (N_15754,N_14553,N_14492);
or U15755 (N_15755,N_15032,N_14993);
and U15756 (N_15756,N_14814,N_14735);
and U15757 (N_15757,N_14801,N_14621);
and U15758 (N_15758,N_14857,N_15045);
nand U15759 (N_15759,N_15040,N_14615);
and U15760 (N_15760,N_14418,N_15155);
or U15761 (N_15761,N_15056,N_14892);
and U15762 (N_15762,N_14638,N_14698);
and U15763 (N_15763,N_15161,N_14657);
and U15764 (N_15764,N_14527,N_14768);
or U15765 (N_15765,N_14711,N_15033);
and U15766 (N_15766,N_14731,N_14744);
nand U15767 (N_15767,N_14992,N_14546);
xor U15768 (N_15768,N_14425,N_14867);
xnor U15769 (N_15769,N_14985,N_15119);
nand U15770 (N_15770,N_15139,N_14432);
or U15771 (N_15771,N_14743,N_14524);
or U15772 (N_15772,N_14775,N_14981);
xnor U15773 (N_15773,N_14560,N_14451);
and U15774 (N_15774,N_14910,N_15084);
nor U15775 (N_15775,N_14897,N_14414);
nand U15776 (N_15776,N_14758,N_14431);
nand U15777 (N_15777,N_15025,N_15006);
xor U15778 (N_15778,N_15177,N_14949);
and U15779 (N_15779,N_14878,N_14518);
nor U15780 (N_15780,N_14432,N_15137);
nor U15781 (N_15781,N_14669,N_15002);
nand U15782 (N_15782,N_15047,N_15198);
xor U15783 (N_15783,N_14479,N_15026);
nand U15784 (N_15784,N_14865,N_14468);
xnor U15785 (N_15785,N_14471,N_14547);
xor U15786 (N_15786,N_14686,N_14897);
or U15787 (N_15787,N_14541,N_14608);
and U15788 (N_15788,N_15193,N_14952);
or U15789 (N_15789,N_14943,N_15050);
nand U15790 (N_15790,N_14563,N_15165);
xnor U15791 (N_15791,N_15080,N_14688);
or U15792 (N_15792,N_15138,N_14896);
or U15793 (N_15793,N_15109,N_15062);
xor U15794 (N_15794,N_14955,N_15062);
nand U15795 (N_15795,N_14987,N_15109);
nand U15796 (N_15796,N_15168,N_14445);
xor U15797 (N_15797,N_14411,N_14726);
and U15798 (N_15798,N_15100,N_15080);
and U15799 (N_15799,N_14464,N_15011);
nor U15800 (N_15800,N_14792,N_15197);
and U15801 (N_15801,N_14640,N_14893);
xor U15802 (N_15802,N_14804,N_15018);
and U15803 (N_15803,N_15046,N_15062);
nor U15804 (N_15804,N_14943,N_14464);
or U15805 (N_15805,N_14906,N_14407);
xnor U15806 (N_15806,N_15026,N_15088);
nor U15807 (N_15807,N_14757,N_14457);
xor U15808 (N_15808,N_15094,N_14834);
and U15809 (N_15809,N_14622,N_15040);
nor U15810 (N_15810,N_14819,N_14462);
or U15811 (N_15811,N_14880,N_14863);
nor U15812 (N_15812,N_14584,N_14847);
or U15813 (N_15813,N_15174,N_14549);
and U15814 (N_15814,N_15009,N_14513);
xnor U15815 (N_15815,N_14702,N_14645);
and U15816 (N_15816,N_14421,N_14832);
xnor U15817 (N_15817,N_15182,N_14414);
nor U15818 (N_15818,N_14547,N_15083);
nand U15819 (N_15819,N_15079,N_14987);
or U15820 (N_15820,N_14860,N_14581);
nor U15821 (N_15821,N_15047,N_14774);
nand U15822 (N_15822,N_14538,N_14999);
nand U15823 (N_15823,N_14774,N_14921);
and U15824 (N_15824,N_14848,N_14617);
nor U15825 (N_15825,N_14882,N_15173);
nor U15826 (N_15826,N_15071,N_14910);
xor U15827 (N_15827,N_15166,N_14994);
nor U15828 (N_15828,N_14463,N_14794);
nand U15829 (N_15829,N_14600,N_14439);
xnor U15830 (N_15830,N_14768,N_14954);
nand U15831 (N_15831,N_14435,N_15113);
xnor U15832 (N_15832,N_14699,N_15099);
and U15833 (N_15833,N_15009,N_14815);
and U15834 (N_15834,N_14444,N_14489);
or U15835 (N_15835,N_14747,N_15007);
and U15836 (N_15836,N_14400,N_14707);
or U15837 (N_15837,N_14911,N_14876);
nand U15838 (N_15838,N_14538,N_14643);
xor U15839 (N_15839,N_14759,N_14405);
xnor U15840 (N_15840,N_14619,N_14827);
and U15841 (N_15841,N_14957,N_15087);
or U15842 (N_15842,N_14464,N_14896);
xor U15843 (N_15843,N_14640,N_15105);
and U15844 (N_15844,N_14604,N_14593);
xor U15845 (N_15845,N_14982,N_14545);
nor U15846 (N_15846,N_15076,N_14960);
nor U15847 (N_15847,N_15177,N_14656);
or U15848 (N_15848,N_15066,N_14651);
xor U15849 (N_15849,N_14972,N_14781);
xor U15850 (N_15850,N_14618,N_14660);
nand U15851 (N_15851,N_14659,N_14612);
nor U15852 (N_15852,N_15001,N_14701);
xnor U15853 (N_15853,N_15015,N_15066);
nand U15854 (N_15854,N_14933,N_15038);
or U15855 (N_15855,N_15093,N_15002);
or U15856 (N_15856,N_14488,N_14828);
or U15857 (N_15857,N_14524,N_14860);
nand U15858 (N_15858,N_15059,N_14566);
nand U15859 (N_15859,N_14594,N_14471);
or U15860 (N_15860,N_14858,N_14704);
xnor U15861 (N_15861,N_14882,N_15124);
or U15862 (N_15862,N_14944,N_15120);
xor U15863 (N_15863,N_14497,N_14660);
nor U15864 (N_15864,N_15117,N_14475);
xor U15865 (N_15865,N_14804,N_14814);
and U15866 (N_15866,N_14881,N_15055);
and U15867 (N_15867,N_14684,N_14895);
xnor U15868 (N_15868,N_14541,N_14472);
xor U15869 (N_15869,N_14967,N_14828);
and U15870 (N_15870,N_14820,N_14679);
and U15871 (N_15871,N_14502,N_14649);
and U15872 (N_15872,N_14430,N_15079);
or U15873 (N_15873,N_14849,N_14971);
xnor U15874 (N_15874,N_14949,N_14859);
nor U15875 (N_15875,N_14533,N_15147);
and U15876 (N_15876,N_15116,N_15166);
and U15877 (N_15877,N_14777,N_15012);
or U15878 (N_15878,N_15109,N_14944);
or U15879 (N_15879,N_14438,N_14749);
nor U15880 (N_15880,N_14437,N_14415);
xnor U15881 (N_15881,N_14796,N_14531);
or U15882 (N_15882,N_14966,N_14778);
or U15883 (N_15883,N_14706,N_14468);
nand U15884 (N_15884,N_15020,N_14813);
nand U15885 (N_15885,N_15173,N_14993);
nand U15886 (N_15886,N_14971,N_14942);
or U15887 (N_15887,N_14935,N_15145);
and U15888 (N_15888,N_14953,N_14626);
nand U15889 (N_15889,N_14828,N_15051);
or U15890 (N_15890,N_14619,N_14921);
nor U15891 (N_15891,N_14849,N_14559);
nand U15892 (N_15892,N_14402,N_14512);
nor U15893 (N_15893,N_14457,N_14946);
xnor U15894 (N_15894,N_15066,N_14502);
and U15895 (N_15895,N_14703,N_14725);
or U15896 (N_15896,N_14441,N_14734);
nor U15897 (N_15897,N_14656,N_15145);
xnor U15898 (N_15898,N_14412,N_14613);
nor U15899 (N_15899,N_14869,N_14799);
nand U15900 (N_15900,N_14753,N_15022);
nor U15901 (N_15901,N_14497,N_14631);
or U15902 (N_15902,N_14944,N_14752);
or U15903 (N_15903,N_14700,N_15143);
nor U15904 (N_15904,N_14780,N_14971);
and U15905 (N_15905,N_14811,N_14715);
nor U15906 (N_15906,N_14620,N_14538);
or U15907 (N_15907,N_14680,N_14470);
xnor U15908 (N_15908,N_14415,N_14833);
nor U15909 (N_15909,N_15037,N_14901);
xnor U15910 (N_15910,N_14562,N_14482);
nor U15911 (N_15911,N_14567,N_14621);
xnor U15912 (N_15912,N_14487,N_14489);
or U15913 (N_15913,N_14960,N_14706);
xnor U15914 (N_15914,N_14770,N_14736);
nand U15915 (N_15915,N_14721,N_15170);
nand U15916 (N_15916,N_15077,N_15106);
xnor U15917 (N_15917,N_15071,N_15113);
and U15918 (N_15918,N_15113,N_15100);
nand U15919 (N_15919,N_14797,N_14681);
and U15920 (N_15920,N_14753,N_14516);
or U15921 (N_15921,N_14593,N_14938);
or U15922 (N_15922,N_14681,N_14429);
and U15923 (N_15923,N_15071,N_14731);
nand U15924 (N_15924,N_14823,N_14594);
nand U15925 (N_15925,N_14441,N_14647);
nor U15926 (N_15926,N_14824,N_14940);
nor U15927 (N_15927,N_14537,N_14745);
nand U15928 (N_15928,N_15162,N_15112);
and U15929 (N_15929,N_14553,N_14846);
and U15930 (N_15930,N_14914,N_15113);
nor U15931 (N_15931,N_14466,N_14631);
nor U15932 (N_15932,N_14530,N_15131);
or U15933 (N_15933,N_15128,N_14531);
nand U15934 (N_15934,N_15144,N_14794);
nand U15935 (N_15935,N_15023,N_14818);
xnor U15936 (N_15936,N_14878,N_14777);
or U15937 (N_15937,N_14573,N_14653);
xor U15938 (N_15938,N_14731,N_14900);
or U15939 (N_15939,N_14878,N_14914);
nand U15940 (N_15940,N_14896,N_14411);
and U15941 (N_15941,N_14768,N_14504);
and U15942 (N_15942,N_14879,N_14420);
nand U15943 (N_15943,N_15030,N_14888);
nand U15944 (N_15944,N_15016,N_14587);
nor U15945 (N_15945,N_14856,N_14983);
and U15946 (N_15946,N_14705,N_14754);
nor U15947 (N_15947,N_15186,N_14676);
nor U15948 (N_15948,N_14725,N_14980);
xnor U15949 (N_15949,N_14750,N_14833);
nand U15950 (N_15950,N_15031,N_14441);
and U15951 (N_15951,N_14415,N_14701);
nand U15952 (N_15952,N_15027,N_14618);
nand U15953 (N_15953,N_14941,N_14529);
nand U15954 (N_15954,N_14578,N_15097);
or U15955 (N_15955,N_14803,N_14528);
nor U15956 (N_15956,N_14684,N_14787);
nor U15957 (N_15957,N_14792,N_15172);
or U15958 (N_15958,N_14513,N_14667);
xnor U15959 (N_15959,N_15024,N_14994);
nor U15960 (N_15960,N_15124,N_15000);
and U15961 (N_15961,N_15174,N_14794);
and U15962 (N_15962,N_15146,N_14739);
and U15963 (N_15963,N_14801,N_14443);
and U15964 (N_15964,N_15110,N_14777);
nand U15965 (N_15965,N_14898,N_14592);
nand U15966 (N_15966,N_14541,N_14598);
and U15967 (N_15967,N_14954,N_14519);
nor U15968 (N_15968,N_15065,N_14753);
nand U15969 (N_15969,N_14968,N_14615);
and U15970 (N_15970,N_14812,N_14814);
or U15971 (N_15971,N_15139,N_14642);
nor U15972 (N_15972,N_14772,N_14878);
xnor U15973 (N_15973,N_14538,N_15199);
or U15974 (N_15974,N_14681,N_15003);
nor U15975 (N_15975,N_14407,N_14951);
or U15976 (N_15976,N_14775,N_14577);
xor U15977 (N_15977,N_15122,N_14429);
and U15978 (N_15978,N_14801,N_14960);
nand U15979 (N_15979,N_15020,N_14667);
nand U15980 (N_15980,N_14618,N_14836);
and U15981 (N_15981,N_15138,N_14510);
nor U15982 (N_15982,N_15176,N_14749);
nor U15983 (N_15983,N_14673,N_14574);
or U15984 (N_15984,N_14401,N_15143);
xnor U15985 (N_15985,N_15055,N_14801);
nor U15986 (N_15986,N_14552,N_14881);
nand U15987 (N_15987,N_14415,N_15115);
or U15988 (N_15988,N_14896,N_14895);
xnor U15989 (N_15989,N_14735,N_14823);
xnor U15990 (N_15990,N_14930,N_14556);
or U15991 (N_15991,N_14425,N_14969);
nor U15992 (N_15992,N_14781,N_14645);
nand U15993 (N_15993,N_14500,N_15032);
or U15994 (N_15994,N_14544,N_14594);
nand U15995 (N_15995,N_15077,N_14794);
and U15996 (N_15996,N_14855,N_15015);
or U15997 (N_15997,N_14507,N_15065);
xor U15998 (N_15998,N_14887,N_14585);
and U15999 (N_15999,N_14460,N_14587);
or U16000 (N_16000,N_15740,N_15295);
nor U16001 (N_16001,N_15439,N_15917);
or U16002 (N_16002,N_15586,N_15314);
nor U16003 (N_16003,N_15367,N_15371);
nor U16004 (N_16004,N_15827,N_15872);
or U16005 (N_16005,N_15700,N_15507);
xor U16006 (N_16006,N_15289,N_15547);
nand U16007 (N_16007,N_15823,N_15897);
nand U16008 (N_16008,N_15681,N_15683);
nand U16009 (N_16009,N_15541,N_15247);
nor U16010 (N_16010,N_15529,N_15277);
and U16011 (N_16011,N_15401,N_15616);
nor U16012 (N_16012,N_15527,N_15476);
and U16013 (N_16013,N_15426,N_15319);
nor U16014 (N_16014,N_15971,N_15810);
nor U16015 (N_16015,N_15299,N_15479);
and U16016 (N_16016,N_15505,N_15378);
nand U16017 (N_16017,N_15233,N_15407);
xor U16018 (N_16018,N_15656,N_15264);
xnor U16019 (N_16019,N_15565,N_15432);
or U16020 (N_16020,N_15443,N_15931);
and U16021 (N_16021,N_15337,N_15634);
nor U16022 (N_16022,N_15631,N_15761);
and U16023 (N_16023,N_15321,N_15224);
xor U16024 (N_16024,N_15765,N_15974);
or U16025 (N_16025,N_15579,N_15771);
xor U16026 (N_16026,N_15569,N_15228);
nand U16027 (N_16027,N_15686,N_15613);
or U16028 (N_16028,N_15454,N_15366);
or U16029 (N_16029,N_15817,N_15511);
and U16030 (N_16030,N_15294,N_15252);
or U16031 (N_16031,N_15259,N_15865);
nand U16032 (N_16032,N_15288,N_15987);
xor U16033 (N_16033,N_15802,N_15861);
xnor U16034 (N_16034,N_15862,N_15855);
and U16035 (N_16035,N_15414,N_15302);
nand U16036 (N_16036,N_15404,N_15261);
xor U16037 (N_16037,N_15729,N_15420);
and U16038 (N_16038,N_15941,N_15398);
xor U16039 (N_16039,N_15455,N_15839);
and U16040 (N_16040,N_15465,N_15643);
or U16041 (N_16041,N_15637,N_15497);
and U16042 (N_16042,N_15622,N_15304);
or U16043 (N_16043,N_15782,N_15756);
nor U16044 (N_16044,N_15399,N_15967);
xnor U16045 (N_16045,N_15478,N_15836);
nand U16046 (N_16046,N_15453,N_15223);
and U16047 (N_16047,N_15516,N_15303);
nor U16048 (N_16048,N_15991,N_15544);
or U16049 (N_16049,N_15738,N_15308);
xnor U16050 (N_16050,N_15667,N_15781);
xor U16051 (N_16051,N_15945,N_15847);
and U16052 (N_16052,N_15888,N_15920);
nor U16053 (N_16053,N_15447,N_15301);
nand U16054 (N_16054,N_15969,N_15253);
nand U16055 (N_16055,N_15203,N_15627);
xor U16056 (N_16056,N_15682,N_15200);
xnor U16057 (N_16057,N_15947,N_15809);
and U16058 (N_16058,N_15720,N_15585);
nor U16059 (N_16059,N_15481,N_15821);
nor U16060 (N_16060,N_15560,N_15226);
nand U16061 (N_16061,N_15676,N_15361);
and U16062 (N_16062,N_15789,N_15279);
and U16063 (N_16063,N_15572,N_15512);
xor U16064 (N_16064,N_15796,N_15340);
and U16065 (N_16065,N_15548,N_15628);
and U16066 (N_16066,N_15430,N_15928);
nor U16067 (N_16067,N_15229,N_15495);
xor U16068 (N_16068,N_15978,N_15212);
or U16069 (N_16069,N_15778,N_15813);
and U16070 (N_16070,N_15415,N_15514);
xor U16071 (N_16071,N_15678,N_15513);
nor U16072 (N_16072,N_15262,N_15687);
nor U16073 (N_16073,N_15446,N_15214);
and U16074 (N_16074,N_15577,N_15602);
nand U16075 (N_16075,N_15853,N_15835);
and U16076 (N_16076,N_15213,N_15359);
nand U16077 (N_16077,N_15843,N_15311);
and U16078 (N_16078,N_15721,N_15743);
or U16079 (N_16079,N_15763,N_15640);
nand U16080 (N_16080,N_15912,N_15309);
nand U16081 (N_16081,N_15911,N_15671);
nor U16082 (N_16082,N_15292,N_15868);
and U16083 (N_16083,N_15717,N_15388);
nor U16084 (N_16084,N_15764,N_15986);
nor U16085 (N_16085,N_15240,N_15286);
and U16086 (N_16086,N_15387,N_15799);
xnor U16087 (N_16087,N_15329,N_15392);
xnor U16088 (N_16088,N_15298,N_15276);
or U16089 (N_16089,N_15549,N_15451);
nor U16090 (N_16090,N_15612,N_15775);
and U16091 (N_16091,N_15290,N_15840);
nand U16092 (N_16092,N_15900,N_15377);
or U16093 (N_16093,N_15403,N_15747);
xor U16094 (N_16094,N_15578,N_15996);
nand U16095 (N_16095,N_15711,N_15610);
xnor U16096 (N_16096,N_15207,N_15982);
and U16097 (N_16097,N_15472,N_15882);
nand U16098 (N_16098,N_15825,N_15730);
nand U16099 (N_16099,N_15217,N_15929);
nor U16100 (N_16100,N_15425,N_15693);
nand U16101 (N_16101,N_15658,N_15633);
nand U16102 (N_16102,N_15956,N_15755);
xor U16103 (N_16103,N_15770,N_15583);
or U16104 (N_16104,N_15669,N_15632);
nor U16105 (N_16105,N_15339,N_15558);
nor U16106 (N_16106,N_15468,N_15871);
xor U16107 (N_16107,N_15875,N_15604);
nor U16108 (N_16108,N_15551,N_15600);
xor U16109 (N_16109,N_15249,N_15508);
nand U16110 (N_16110,N_15357,N_15341);
nor U16111 (N_16111,N_15829,N_15312);
nor U16112 (N_16112,N_15691,N_15227);
nand U16113 (N_16113,N_15411,N_15570);
xor U16114 (N_16114,N_15533,N_15927);
nor U16115 (N_16115,N_15464,N_15494);
nor U16116 (N_16116,N_15694,N_15762);
or U16117 (N_16117,N_15940,N_15325);
and U16118 (N_16118,N_15305,N_15489);
nand U16119 (N_16119,N_15296,N_15383);
nand U16120 (N_16120,N_15313,N_15488);
nor U16121 (N_16121,N_15716,N_15904);
and U16122 (N_16122,N_15588,N_15343);
xnor U16123 (N_16123,N_15891,N_15381);
or U16124 (N_16124,N_15206,N_15449);
xnor U16125 (N_16125,N_15543,N_15473);
nand U16126 (N_16126,N_15814,N_15930);
nor U16127 (N_16127,N_15863,N_15760);
nor U16128 (N_16128,N_15662,N_15958);
and U16129 (N_16129,N_15221,N_15858);
nand U16130 (N_16130,N_15587,N_15611);
xnor U16131 (N_16131,N_15287,N_15722);
and U16132 (N_16132,N_15718,N_15393);
or U16133 (N_16133,N_15310,N_15910);
nor U16134 (N_16134,N_15406,N_15674);
and U16135 (N_16135,N_15624,N_15396);
nor U16136 (N_16136,N_15499,N_15575);
nand U16137 (N_16137,N_15703,N_15670);
and U16138 (N_16138,N_15737,N_15650);
and U16139 (N_16139,N_15477,N_15556);
nor U16140 (N_16140,N_15554,N_15370);
nor U16141 (N_16141,N_15250,N_15386);
xnor U16142 (N_16142,N_15772,N_15204);
or U16143 (N_16143,N_15757,N_15784);
nor U16144 (N_16144,N_15293,N_15444);
xor U16145 (N_16145,N_15709,N_15780);
xnor U16146 (N_16146,N_15423,N_15812);
and U16147 (N_16147,N_15939,N_15807);
or U16148 (N_16148,N_15883,N_15635);
nor U16149 (N_16149,N_15485,N_15258);
nand U16150 (N_16150,N_15663,N_15648);
nand U16151 (N_16151,N_15651,N_15768);
xor U16152 (N_16152,N_15461,N_15922);
and U16153 (N_16153,N_15838,N_15921);
nand U16154 (N_16154,N_15324,N_15723);
and U16155 (N_16155,N_15269,N_15675);
or U16156 (N_16156,N_15714,N_15470);
and U16157 (N_16157,N_15475,N_15915);
nor U16158 (N_16158,N_15205,N_15382);
nand U16159 (N_16159,N_15774,N_15952);
nand U16160 (N_16160,N_15484,N_15445);
and U16161 (N_16161,N_15608,N_15278);
xor U16162 (N_16162,N_15758,N_15496);
nor U16163 (N_16163,N_15988,N_15788);
nand U16164 (N_16164,N_15246,N_15878);
nand U16165 (N_16165,N_15316,N_15210);
xnor U16166 (N_16166,N_15422,N_15356);
or U16167 (N_16167,N_15615,N_15492);
and U16168 (N_16168,N_15498,N_15211);
nand U16169 (N_16169,N_15800,N_15659);
xor U16170 (N_16170,N_15641,N_15236);
and U16171 (N_16171,N_15673,N_15998);
nor U16172 (N_16172,N_15563,N_15255);
xnor U16173 (N_16173,N_15239,N_15742);
nand U16174 (N_16174,N_15360,N_15850);
xor U16175 (N_16175,N_15344,N_15805);
nand U16176 (N_16176,N_15852,N_15333);
nor U16177 (N_16177,N_15429,N_15448);
and U16178 (N_16178,N_15493,N_15786);
and U16179 (N_16179,N_15741,N_15243);
xnor U16180 (N_16180,N_15935,N_15993);
and U16181 (N_16181,N_15471,N_15906);
and U16182 (N_16182,N_15801,N_15520);
or U16183 (N_16183,N_15968,N_15892);
or U16184 (N_16184,N_15907,N_15725);
and U16185 (N_16185,N_15459,N_15526);
nand U16186 (N_16186,N_15491,N_15502);
xnor U16187 (N_16187,N_15657,N_15525);
xor U16188 (N_16188,N_15363,N_15831);
nand U16189 (N_16189,N_15483,N_15405);
nand U16190 (N_16190,N_15724,N_15894);
nor U16191 (N_16191,N_15625,N_15594);
nand U16192 (N_16192,N_15896,N_15933);
and U16193 (N_16193,N_15617,N_15601);
xnor U16194 (N_16194,N_15826,N_15431);
or U16195 (N_16195,N_15697,N_15591);
xor U16196 (N_16196,N_15260,N_15326);
nor U16197 (N_16197,N_15804,N_15949);
or U16198 (N_16198,N_15649,N_15954);
and U16199 (N_16199,N_15924,N_15402);
nor U16200 (N_16200,N_15873,N_15905);
or U16201 (N_16201,N_15241,N_15561);
or U16202 (N_16202,N_15413,N_15271);
nor U16203 (N_16203,N_15270,N_15620);
xor U16204 (N_16204,N_15965,N_15486);
xnor U16205 (N_16205,N_15469,N_15467);
xnor U16206 (N_16206,N_15267,N_15833);
nor U16207 (N_16207,N_15919,N_15522);
and U16208 (N_16208,N_15946,N_15582);
and U16209 (N_16209,N_15581,N_15934);
or U16210 (N_16210,N_15379,N_15997);
or U16211 (N_16211,N_15745,N_15218);
nor U16212 (N_16212,N_15936,N_15977);
xor U16213 (N_16213,N_15955,N_15734);
or U16214 (N_16214,N_15614,N_15254);
nor U16215 (N_16215,N_15884,N_15690);
xor U16216 (N_16216,N_15530,N_15566);
and U16217 (N_16217,N_15792,N_15731);
xnor U16218 (N_16218,N_15966,N_15441);
or U16219 (N_16219,N_15886,N_15391);
or U16220 (N_16220,N_15732,N_15607);
and U16221 (N_16221,N_15474,N_15668);
nand U16222 (N_16222,N_15281,N_15679);
and U16223 (N_16223,N_15440,N_15854);
nor U16224 (N_16224,N_15960,N_15421);
xnor U16225 (N_16225,N_15848,N_15948);
xnor U16226 (N_16226,N_15452,N_15598);
nor U16227 (N_16227,N_15653,N_15918);
xnor U16228 (N_16228,N_15794,N_15623);
nor U16229 (N_16229,N_15348,N_15553);
nand U16230 (N_16230,N_15975,N_15538);
nand U16231 (N_16231,N_15819,N_15932);
nor U16232 (N_16232,N_15701,N_15593);
nand U16233 (N_16233,N_15973,N_15606);
and U16234 (N_16234,N_15595,N_15428);
nor U16235 (N_16235,N_15707,N_15201);
nor U16236 (N_16236,N_15592,N_15751);
and U16237 (N_16237,N_15487,N_15688);
nor U16238 (N_16238,N_15803,N_15291);
xor U16239 (N_16239,N_15950,N_15903);
or U16240 (N_16240,N_15434,N_15866);
or U16241 (N_16241,N_15272,N_15646);
or U16242 (N_16242,N_15597,N_15713);
or U16243 (N_16243,N_15546,N_15376);
nand U16244 (N_16244,N_15735,N_15989);
nor U16245 (N_16245,N_15590,N_15841);
nor U16246 (N_16246,N_15859,N_15899);
and U16247 (N_16247,N_15545,N_15317);
xor U16248 (N_16248,N_15282,N_15876);
nand U16249 (N_16249,N_15754,N_15573);
xnor U16250 (N_16250,N_15914,N_15696);
or U16251 (N_16251,N_15437,N_15540);
nand U16252 (N_16252,N_15380,N_15564);
xor U16253 (N_16253,N_15216,N_15457);
or U16254 (N_16254,N_15273,N_15834);
xnor U16255 (N_16255,N_15231,N_15300);
nand U16256 (N_16256,N_15787,N_15209);
and U16257 (N_16257,N_15571,N_15698);
and U16258 (N_16258,N_15542,N_15373);
xnor U16259 (N_16259,N_15685,N_15857);
or U16260 (N_16260,N_15394,N_15793);
and U16261 (N_16261,N_15418,N_15744);
xnor U16262 (N_16262,N_15684,N_15318);
and U16263 (N_16263,N_15889,N_15902);
or U16264 (N_16264,N_15925,N_15500);
or U16265 (N_16265,N_15568,N_15664);
or U16266 (N_16266,N_15528,N_15389);
nor U16267 (N_16267,N_15524,N_15335);
nor U16268 (N_16268,N_15712,N_15222);
nor U16269 (N_16269,N_15776,N_15753);
xor U16270 (N_16270,N_15885,N_15962);
xnor U16271 (N_16271,N_15395,N_15364);
or U16272 (N_16272,N_15702,N_15790);
xnor U16273 (N_16273,N_15436,N_15680);
nand U16274 (N_16274,N_15596,N_15976);
nor U16275 (N_16275,N_15957,N_15938);
xnor U16276 (N_16276,N_15944,N_15661);
or U16277 (N_16277,N_15943,N_15518);
nor U16278 (N_16278,N_15342,N_15980);
or U16279 (N_16279,N_15959,N_15797);
and U16280 (N_16280,N_15963,N_15257);
xnor U16281 (N_16281,N_15639,N_15515);
nor U16282 (N_16282,N_15323,N_15759);
or U16283 (N_16283,N_15567,N_15749);
xor U16284 (N_16284,N_15618,N_15879);
or U16285 (N_16285,N_15926,N_15652);
xor U16286 (N_16286,N_15777,N_15412);
nand U16287 (N_16287,N_15985,N_15739);
xnor U16288 (N_16288,N_15202,N_15748);
nand U16289 (N_16289,N_15242,N_15877);
nor U16290 (N_16290,N_15315,N_15630);
xor U16291 (N_16291,N_15346,N_15999);
nor U16292 (N_16292,N_15860,N_15844);
and U16293 (N_16293,N_15867,N_15887);
or U16294 (N_16294,N_15603,N_15208);
nand U16295 (N_16295,N_15283,N_15609);
nor U16296 (N_16296,N_15248,N_15880);
and U16297 (N_16297,N_15951,N_15898);
xor U16298 (N_16298,N_15390,N_15372);
and U16299 (N_16299,N_15766,N_15345);
nor U16300 (N_16300,N_15235,N_15320);
nand U16301 (N_16301,N_15913,N_15795);
nand U16302 (N_16302,N_15708,N_15332);
nand U16303 (N_16303,N_15846,N_15334);
xnor U16304 (N_16304,N_15647,N_15791);
or U16305 (N_16305,N_15306,N_15909);
and U16306 (N_16306,N_15280,N_15984);
nand U16307 (N_16307,N_15728,N_15397);
nor U16308 (N_16308,N_15644,N_15773);
or U16309 (N_16309,N_15665,N_15419);
and U16310 (N_16310,N_15689,N_15580);
and U16311 (N_16311,N_15256,N_15816);
or U16312 (N_16312,N_15562,N_15438);
nand U16313 (N_16313,N_15336,N_15501);
xor U16314 (N_16314,N_15504,N_15535);
nand U16315 (N_16315,N_15266,N_15715);
nand U16316 (N_16316,N_15752,N_15830);
or U16317 (N_16317,N_15869,N_15619);
nand U16318 (N_16318,N_15655,N_15284);
nor U16319 (N_16319,N_15785,N_15350);
or U16320 (N_16320,N_15808,N_15979);
nand U16321 (N_16321,N_15274,N_15510);
xnor U16322 (N_16322,N_15881,N_15400);
and U16323 (N_16323,N_15574,N_15517);
nor U16324 (N_16324,N_15523,N_15820);
xor U16325 (N_16325,N_15727,N_15845);
xnor U16326 (N_16326,N_15338,N_15557);
nand U16327 (N_16327,N_15972,N_15358);
xor U16328 (N_16328,N_15408,N_15417);
nand U16329 (N_16329,N_15937,N_15942);
nand U16330 (N_16330,N_15285,N_15244);
xnor U16331 (N_16331,N_15828,N_15769);
or U16332 (N_16332,N_15695,N_15990);
or U16333 (N_16333,N_15626,N_15456);
or U16334 (N_16334,N_15874,N_15482);
nand U16335 (N_16335,N_15265,N_15552);
xnor U16336 (N_16336,N_15352,N_15832);
nand U16337 (N_16337,N_15442,N_15666);
or U16338 (N_16338,N_15532,N_15427);
nor U16339 (N_16339,N_15531,N_15923);
nor U16340 (N_16340,N_15462,N_15331);
xor U16341 (N_16341,N_15964,N_15353);
nor U16342 (N_16342,N_15837,N_15490);
xor U16343 (N_16343,N_15995,N_15327);
nand U16344 (N_16344,N_15726,N_15706);
xnor U16345 (N_16345,N_15463,N_15234);
nor U16346 (N_16346,N_15719,N_15705);
nand U16347 (N_16347,N_15798,N_15375);
nor U16348 (N_16348,N_15736,N_15297);
xor U16349 (N_16349,N_15642,N_15374);
and U16350 (N_16350,N_15355,N_15433);
or U16351 (N_16351,N_15220,N_15779);
nor U16352 (N_16352,N_15672,N_15576);
or U16353 (N_16353,N_15783,N_15699);
nand U16354 (N_16354,N_15811,N_15368);
nand U16355 (N_16355,N_15645,N_15232);
nand U16356 (N_16356,N_15654,N_15215);
nand U16357 (N_16357,N_15384,N_15307);
or U16358 (N_16358,N_15901,N_15605);
and U16359 (N_16359,N_15385,N_15815);
xnor U16360 (N_16360,N_15851,N_15822);
nor U16361 (N_16361,N_15509,N_15354);
nor U16362 (N_16362,N_15322,N_15369);
or U16363 (N_16363,N_15347,N_15503);
xnor U16364 (N_16364,N_15584,N_15870);
nor U16365 (N_16365,N_15856,N_15424);
xnor U16366 (N_16366,N_15225,N_15245);
nand U16367 (N_16367,N_15994,N_15351);
and U16368 (N_16368,N_15519,N_15636);
and U16369 (N_16369,N_15466,N_15767);
and U16370 (N_16370,N_15746,N_15733);
nand U16371 (N_16371,N_15537,N_15983);
nand U16372 (N_16372,N_15961,N_15330);
and U16373 (N_16373,N_15704,N_15849);
xnor U16374 (N_16374,N_15895,N_15458);
or U16375 (N_16375,N_15710,N_15409);
nand U16376 (N_16376,N_15806,N_15435);
nand U16377 (N_16377,N_15893,N_15692);
nor U16378 (N_16378,N_15521,N_15237);
or U16379 (N_16379,N_15621,N_15629);
and U16380 (N_16380,N_15263,N_15506);
or U16381 (N_16381,N_15589,N_15890);
nand U16382 (N_16382,N_15599,N_15328);
nor U16383 (N_16383,N_15908,N_15916);
xor U16384 (N_16384,N_15362,N_15238);
and U16385 (N_16385,N_15555,N_15219);
nor U16386 (N_16386,N_15638,N_15460);
or U16387 (N_16387,N_15410,N_15550);
nor U16388 (N_16388,N_15534,N_15268);
and U16389 (N_16389,N_15349,N_15660);
and U16390 (N_16390,N_15677,N_15536);
xnor U16391 (N_16391,N_15450,N_15230);
and U16392 (N_16392,N_15539,N_15275);
nor U16393 (N_16393,N_15953,N_15559);
nor U16394 (N_16394,N_15416,N_15750);
xnor U16395 (N_16395,N_15824,N_15480);
nor U16396 (N_16396,N_15992,N_15981);
or U16397 (N_16397,N_15365,N_15970);
nand U16398 (N_16398,N_15842,N_15251);
xnor U16399 (N_16399,N_15864,N_15818);
nor U16400 (N_16400,N_15882,N_15505);
nor U16401 (N_16401,N_15722,N_15689);
and U16402 (N_16402,N_15349,N_15235);
xnor U16403 (N_16403,N_15553,N_15576);
and U16404 (N_16404,N_15636,N_15620);
nor U16405 (N_16405,N_15756,N_15967);
nand U16406 (N_16406,N_15289,N_15887);
nor U16407 (N_16407,N_15772,N_15691);
xor U16408 (N_16408,N_15498,N_15601);
nor U16409 (N_16409,N_15386,N_15749);
xor U16410 (N_16410,N_15294,N_15875);
and U16411 (N_16411,N_15903,N_15985);
or U16412 (N_16412,N_15728,N_15920);
nor U16413 (N_16413,N_15286,N_15799);
and U16414 (N_16414,N_15978,N_15730);
or U16415 (N_16415,N_15224,N_15632);
or U16416 (N_16416,N_15582,N_15927);
and U16417 (N_16417,N_15207,N_15735);
and U16418 (N_16418,N_15609,N_15678);
nand U16419 (N_16419,N_15602,N_15943);
nor U16420 (N_16420,N_15579,N_15770);
nor U16421 (N_16421,N_15325,N_15212);
nand U16422 (N_16422,N_15212,N_15301);
xnor U16423 (N_16423,N_15475,N_15957);
or U16424 (N_16424,N_15512,N_15573);
or U16425 (N_16425,N_15784,N_15311);
and U16426 (N_16426,N_15633,N_15954);
nand U16427 (N_16427,N_15732,N_15545);
and U16428 (N_16428,N_15204,N_15903);
or U16429 (N_16429,N_15923,N_15520);
and U16430 (N_16430,N_15207,N_15261);
or U16431 (N_16431,N_15352,N_15598);
nor U16432 (N_16432,N_15873,N_15511);
xnor U16433 (N_16433,N_15797,N_15936);
nor U16434 (N_16434,N_15269,N_15802);
nor U16435 (N_16435,N_15257,N_15423);
or U16436 (N_16436,N_15712,N_15846);
nor U16437 (N_16437,N_15918,N_15830);
and U16438 (N_16438,N_15463,N_15935);
nor U16439 (N_16439,N_15202,N_15719);
or U16440 (N_16440,N_15541,N_15225);
nor U16441 (N_16441,N_15235,N_15631);
and U16442 (N_16442,N_15470,N_15395);
and U16443 (N_16443,N_15335,N_15868);
nor U16444 (N_16444,N_15572,N_15660);
or U16445 (N_16445,N_15828,N_15551);
or U16446 (N_16446,N_15977,N_15358);
xnor U16447 (N_16447,N_15631,N_15644);
nand U16448 (N_16448,N_15956,N_15446);
xnor U16449 (N_16449,N_15849,N_15260);
or U16450 (N_16450,N_15734,N_15910);
xor U16451 (N_16451,N_15552,N_15499);
or U16452 (N_16452,N_15263,N_15708);
nor U16453 (N_16453,N_15608,N_15999);
and U16454 (N_16454,N_15674,N_15672);
xor U16455 (N_16455,N_15686,N_15552);
nand U16456 (N_16456,N_15537,N_15416);
and U16457 (N_16457,N_15289,N_15794);
xor U16458 (N_16458,N_15336,N_15938);
xnor U16459 (N_16459,N_15545,N_15743);
and U16460 (N_16460,N_15959,N_15790);
or U16461 (N_16461,N_15273,N_15651);
or U16462 (N_16462,N_15408,N_15456);
or U16463 (N_16463,N_15260,N_15690);
xor U16464 (N_16464,N_15925,N_15304);
and U16465 (N_16465,N_15904,N_15228);
and U16466 (N_16466,N_15921,N_15749);
and U16467 (N_16467,N_15254,N_15703);
xor U16468 (N_16468,N_15389,N_15721);
and U16469 (N_16469,N_15921,N_15618);
or U16470 (N_16470,N_15979,N_15997);
and U16471 (N_16471,N_15793,N_15932);
or U16472 (N_16472,N_15934,N_15669);
and U16473 (N_16473,N_15801,N_15540);
nor U16474 (N_16474,N_15228,N_15521);
nor U16475 (N_16475,N_15744,N_15474);
nor U16476 (N_16476,N_15241,N_15502);
xnor U16477 (N_16477,N_15816,N_15312);
nor U16478 (N_16478,N_15239,N_15518);
xor U16479 (N_16479,N_15473,N_15781);
or U16480 (N_16480,N_15979,N_15915);
nor U16481 (N_16481,N_15933,N_15213);
or U16482 (N_16482,N_15412,N_15813);
nor U16483 (N_16483,N_15869,N_15639);
xor U16484 (N_16484,N_15907,N_15713);
or U16485 (N_16485,N_15203,N_15338);
and U16486 (N_16486,N_15418,N_15381);
xor U16487 (N_16487,N_15944,N_15841);
and U16488 (N_16488,N_15466,N_15851);
or U16489 (N_16489,N_15824,N_15489);
nand U16490 (N_16490,N_15994,N_15711);
and U16491 (N_16491,N_15742,N_15482);
xnor U16492 (N_16492,N_15235,N_15501);
xor U16493 (N_16493,N_15816,N_15500);
and U16494 (N_16494,N_15421,N_15536);
nor U16495 (N_16495,N_15275,N_15689);
nand U16496 (N_16496,N_15716,N_15241);
nand U16497 (N_16497,N_15533,N_15996);
nand U16498 (N_16498,N_15261,N_15369);
or U16499 (N_16499,N_15469,N_15221);
or U16500 (N_16500,N_15441,N_15730);
and U16501 (N_16501,N_15949,N_15875);
xor U16502 (N_16502,N_15586,N_15234);
nand U16503 (N_16503,N_15932,N_15341);
nand U16504 (N_16504,N_15976,N_15939);
xor U16505 (N_16505,N_15533,N_15974);
nor U16506 (N_16506,N_15905,N_15876);
and U16507 (N_16507,N_15236,N_15581);
xor U16508 (N_16508,N_15505,N_15974);
or U16509 (N_16509,N_15279,N_15771);
and U16510 (N_16510,N_15806,N_15622);
nand U16511 (N_16511,N_15723,N_15845);
nand U16512 (N_16512,N_15214,N_15375);
nor U16513 (N_16513,N_15816,N_15309);
xor U16514 (N_16514,N_15831,N_15372);
nor U16515 (N_16515,N_15227,N_15928);
nand U16516 (N_16516,N_15236,N_15632);
nor U16517 (N_16517,N_15429,N_15227);
xor U16518 (N_16518,N_15959,N_15698);
nand U16519 (N_16519,N_15689,N_15300);
and U16520 (N_16520,N_15301,N_15795);
nand U16521 (N_16521,N_15787,N_15952);
xnor U16522 (N_16522,N_15261,N_15968);
or U16523 (N_16523,N_15419,N_15399);
nor U16524 (N_16524,N_15907,N_15985);
nor U16525 (N_16525,N_15588,N_15341);
or U16526 (N_16526,N_15469,N_15889);
nor U16527 (N_16527,N_15588,N_15843);
nand U16528 (N_16528,N_15399,N_15346);
nand U16529 (N_16529,N_15797,N_15916);
xnor U16530 (N_16530,N_15825,N_15398);
nor U16531 (N_16531,N_15568,N_15484);
nor U16532 (N_16532,N_15479,N_15657);
nor U16533 (N_16533,N_15697,N_15640);
nor U16534 (N_16534,N_15886,N_15704);
nor U16535 (N_16535,N_15205,N_15840);
or U16536 (N_16536,N_15562,N_15886);
nor U16537 (N_16537,N_15635,N_15830);
nor U16538 (N_16538,N_15592,N_15397);
nand U16539 (N_16539,N_15490,N_15582);
nand U16540 (N_16540,N_15674,N_15845);
xor U16541 (N_16541,N_15831,N_15694);
nor U16542 (N_16542,N_15985,N_15423);
or U16543 (N_16543,N_15424,N_15611);
xor U16544 (N_16544,N_15622,N_15311);
nand U16545 (N_16545,N_15980,N_15996);
and U16546 (N_16546,N_15972,N_15908);
and U16547 (N_16547,N_15224,N_15577);
nor U16548 (N_16548,N_15430,N_15710);
xnor U16549 (N_16549,N_15876,N_15683);
nor U16550 (N_16550,N_15403,N_15445);
or U16551 (N_16551,N_15768,N_15555);
and U16552 (N_16552,N_15213,N_15253);
and U16553 (N_16553,N_15700,N_15610);
xnor U16554 (N_16554,N_15766,N_15665);
nor U16555 (N_16555,N_15501,N_15376);
and U16556 (N_16556,N_15915,N_15388);
nor U16557 (N_16557,N_15340,N_15290);
or U16558 (N_16558,N_15479,N_15871);
xor U16559 (N_16559,N_15552,N_15526);
nand U16560 (N_16560,N_15806,N_15562);
nand U16561 (N_16561,N_15613,N_15216);
and U16562 (N_16562,N_15458,N_15424);
nor U16563 (N_16563,N_15977,N_15389);
xor U16564 (N_16564,N_15373,N_15407);
nor U16565 (N_16565,N_15315,N_15312);
and U16566 (N_16566,N_15503,N_15560);
or U16567 (N_16567,N_15450,N_15908);
or U16568 (N_16568,N_15624,N_15774);
nand U16569 (N_16569,N_15461,N_15743);
and U16570 (N_16570,N_15440,N_15293);
nand U16571 (N_16571,N_15574,N_15855);
nand U16572 (N_16572,N_15724,N_15315);
nand U16573 (N_16573,N_15466,N_15806);
and U16574 (N_16574,N_15851,N_15875);
or U16575 (N_16575,N_15546,N_15848);
and U16576 (N_16576,N_15824,N_15347);
nor U16577 (N_16577,N_15676,N_15496);
and U16578 (N_16578,N_15567,N_15626);
xor U16579 (N_16579,N_15287,N_15792);
nand U16580 (N_16580,N_15924,N_15986);
nor U16581 (N_16581,N_15472,N_15850);
and U16582 (N_16582,N_15526,N_15227);
xor U16583 (N_16583,N_15631,N_15604);
xor U16584 (N_16584,N_15471,N_15542);
and U16585 (N_16585,N_15270,N_15504);
nor U16586 (N_16586,N_15860,N_15312);
nand U16587 (N_16587,N_15607,N_15525);
nor U16588 (N_16588,N_15440,N_15384);
xnor U16589 (N_16589,N_15513,N_15577);
and U16590 (N_16590,N_15418,N_15380);
and U16591 (N_16591,N_15436,N_15785);
or U16592 (N_16592,N_15608,N_15293);
or U16593 (N_16593,N_15245,N_15506);
and U16594 (N_16594,N_15507,N_15325);
nand U16595 (N_16595,N_15492,N_15440);
xor U16596 (N_16596,N_15499,N_15771);
nand U16597 (N_16597,N_15940,N_15729);
nor U16598 (N_16598,N_15662,N_15473);
nor U16599 (N_16599,N_15815,N_15630);
and U16600 (N_16600,N_15628,N_15403);
and U16601 (N_16601,N_15393,N_15661);
and U16602 (N_16602,N_15365,N_15428);
nor U16603 (N_16603,N_15521,N_15547);
nor U16604 (N_16604,N_15668,N_15706);
and U16605 (N_16605,N_15251,N_15788);
nand U16606 (N_16606,N_15928,N_15209);
nand U16607 (N_16607,N_15420,N_15605);
or U16608 (N_16608,N_15254,N_15389);
or U16609 (N_16609,N_15465,N_15601);
xnor U16610 (N_16610,N_15559,N_15239);
nor U16611 (N_16611,N_15421,N_15663);
nor U16612 (N_16612,N_15824,N_15658);
and U16613 (N_16613,N_15772,N_15859);
nor U16614 (N_16614,N_15231,N_15381);
nor U16615 (N_16615,N_15982,N_15837);
xor U16616 (N_16616,N_15670,N_15416);
nand U16617 (N_16617,N_15756,N_15519);
xnor U16618 (N_16618,N_15375,N_15819);
or U16619 (N_16619,N_15856,N_15821);
and U16620 (N_16620,N_15323,N_15200);
nor U16621 (N_16621,N_15508,N_15281);
or U16622 (N_16622,N_15747,N_15987);
and U16623 (N_16623,N_15287,N_15979);
or U16624 (N_16624,N_15471,N_15457);
nor U16625 (N_16625,N_15230,N_15354);
nand U16626 (N_16626,N_15752,N_15698);
nand U16627 (N_16627,N_15253,N_15285);
nand U16628 (N_16628,N_15916,N_15904);
or U16629 (N_16629,N_15267,N_15485);
nand U16630 (N_16630,N_15921,N_15330);
nand U16631 (N_16631,N_15471,N_15258);
or U16632 (N_16632,N_15638,N_15988);
nor U16633 (N_16633,N_15280,N_15832);
or U16634 (N_16634,N_15310,N_15671);
nor U16635 (N_16635,N_15360,N_15538);
xor U16636 (N_16636,N_15538,N_15301);
xor U16637 (N_16637,N_15649,N_15884);
and U16638 (N_16638,N_15247,N_15812);
nand U16639 (N_16639,N_15755,N_15694);
nand U16640 (N_16640,N_15949,N_15297);
or U16641 (N_16641,N_15999,N_15741);
xor U16642 (N_16642,N_15968,N_15970);
and U16643 (N_16643,N_15300,N_15662);
or U16644 (N_16644,N_15772,N_15275);
nor U16645 (N_16645,N_15613,N_15510);
nor U16646 (N_16646,N_15821,N_15959);
and U16647 (N_16647,N_15344,N_15306);
nand U16648 (N_16648,N_15344,N_15291);
and U16649 (N_16649,N_15397,N_15210);
nand U16650 (N_16650,N_15484,N_15449);
or U16651 (N_16651,N_15771,N_15597);
or U16652 (N_16652,N_15955,N_15309);
xnor U16653 (N_16653,N_15889,N_15525);
or U16654 (N_16654,N_15453,N_15891);
nor U16655 (N_16655,N_15600,N_15431);
and U16656 (N_16656,N_15881,N_15762);
and U16657 (N_16657,N_15699,N_15629);
or U16658 (N_16658,N_15336,N_15596);
and U16659 (N_16659,N_15824,N_15401);
nand U16660 (N_16660,N_15522,N_15390);
or U16661 (N_16661,N_15295,N_15480);
nand U16662 (N_16662,N_15250,N_15744);
xor U16663 (N_16663,N_15477,N_15620);
nand U16664 (N_16664,N_15808,N_15215);
nand U16665 (N_16665,N_15213,N_15555);
nand U16666 (N_16666,N_15936,N_15892);
xnor U16667 (N_16667,N_15589,N_15372);
nor U16668 (N_16668,N_15581,N_15653);
xor U16669 (N_16669,N_15656,N_15715);
and U16670 (N_16670,N_15267,N_15777);
nand U16671 (N_16671,N_15735,N_15463);
nor U16672 (N_16672,N_15965,N_15534);
and U16673 (N_16673,N_15931,N_15968);
or U16674 (N_16674,N_15660,N_15890);
or U16675 (N_16675,N_15215,N_15964);
or U16676 (N_16676,N_15913,N_15779);
nor U16677 (N_16677,N_15311,N_15582);
nor U16678 (N_16678,N_15371,N_15999);
and U16679 (N_16679,N_15837,N_15647);
nand U16680 (N_16680,N_15996,N_15308);
nand U16681 (N_16681,N_15393,N_15727);
nand U16682 (N_16682,N_15450,N_15213);
and U16683 (N_16683,N_15974,N_15714);
xnor U16684 (N_16684,N_15779,N_15674);
nor U16685 (N_16685,N_15354,N_15373);
or U16686 (N_16686,N_15695,N_15408);
nor U16687 (N_16687,N_15540,N_15845);
and U16688 (N_16688,N_15760,N_15518);
xnor U16689 (N_16689,N_15253,N_15241);
and U16690 (N_16690,N_15436,N_15221);
or U16691 (N_16691,N_15284,N_15650);
nand U16692 (N_16692,N_15261,N_15925);
or U16693 (N_16693,N_15788,N_15465);
or U16694 (N_16694,N_15839,N_15351);
xnor U16695 (N_16695,N_15815,N_15846);
nand U16696 (N_16696,N_15852,N_15372);
xor U16697 (N_16697,N_15837,N_15751);
and U16698 (N_16698,N_15624,N_15806);
xnor U16699 (N_16699,N_15689,N_15243);
or U16700 (N_16700,N_15691,N_15706);
nor U16701 (N_16701,N_15322,N_15760);
and U16702 (N_16702,N_15969,N_15298);
nor U16703 (N_16703,N_15229,N_15803);
or U16704 (N_16704,N_15658,N_15248);
xor U16705 (N_16705,N_15353,N_15203);
nor U16706 (N_16706,N_15281,N_15479);
nand U16707 (N_16707,N_15718,N_15363);
nor U16708 (N_16708,N_15891,N_15516);
xor U16709 (N_16709,N_15619,N_15382);
nand U16710 (N_16710,N_15659,N_15832);
xnor U16711 (N_16711,N_15678,N_15819);
nor U16712 (N_16712,N_15973,N_15388);
or U16713 (N_16713,N_15330,N_15285);
or U16714 (N_16714,N_15437,N_15293);
xnor U16715 (N_16715,N_15309,N_15267);
nand U16716 (N_16716,N_15804,N_15399);
nor U16717 (N_16717,N_15330,N_15429);
and U16718 (N_16718,N_15388,N_15724);
and U16719 (N_16719,N_15990,N_15599);
nor U16720 (N_16720,N_15320,N_15291);
nor U16721 (N_16721,N_15593,N_15245);
and U16722 (N_16722,N_15558,N_15439);
or U16723 (N_16723,N_15839,N_15478);
or U16724 (N_16724,N_15367,N_15733);
nor U16725 (N_16725,N_15838,N_15868);
or U16726 (N_16726,N_15396,N_15942);
nand U16727 (N_16727,N_15689,N_15652);
xor U16728 (N_16728,N_15447,N_15722);
and U16729 (N_16729,N_15792,N_15605);
nor U16730 (N_16730,N_15477,N_15615);
or U16731 (N_16731,N_15735,N_15538);
nor U16732 (N_16732,N_15256,N_15690);
xnor U16733 (N_16733,N_15499,N_15700);
xor U16734 (N_16734,N_15983,N_15567);
nor U16735 (N_16735,N_15532,N_15320);
nand U16736 (N_16736,N_15743,N_15488);
xnor U16737 (N_16737,N_15248,N_15871);
nand U16738 (N_16738,N_15560,N_15665);
xor U16739 (N_16739,N_15324,N_15678);
nor U16740 (N_16740,N_15683,N_15504);
nand U16741 (N_16741,N_15429,N_15773);
xor U16742 (N_16742,N_15614,N_15462);
and U16743 (N_16743,N_15229,N_15892);
xor U16744 (N_16744,N_15587,N_15879);
xnor U16745 (N_16745,N_15305,N_15554);
and U16746 (N_16746,N_15519,N_15898);
or U16747 (N_16747,N_15215,N_15935);
nor U16748 (N_16748,N_15643,N_15789);
and U16749 (N_16749,N_15932,N_15233);
nor U16750 (N_16750,N_15557,N_15813);
or U16751 (N_16751,N_15537,N_15294);
nor U16752 (N_16752,N_15684,N_15244);
xor U16753 (N_16753,N_15483,N_15225);
nand U16754 (N_16754,N_15685,N_15318);
nand U16755 (N_16755,N_15943,N_15412);
xor U16756 (N_16756,N_15347,N_15925);
nor U16757 (N_16757,N_15353,N_15454);
or U16758 (N_16758,N_15250,N_15963);
xnor U16759 (N_16759,N_15786,N_15294);
xor U16760 (N_16760,N_15769,N_15495);
nor U16761 (N_16761,N_15870,N_15288);
xnor U16762 (N_16762,N_15759,N_15388);
and U16763 (N_16763,N_15620,N_15319);
xnor U16764 (N_16764,N_15226,N_15392);
and U16765 (N_16765,N_15513,N_15874);
nand U16766 (N_16766,N_15570,N_15644);
nand U16767 (N_16767,N_15305,N_15767);
xor U16768 (N_16768,N_15446,N_15812);
and U16769 (N_16769,N_15462,N_15562);
and U16770 (N_16770,N_15767,N_15990);
nand U16771 (N_16771,N_15979,N_15849);
nor U16772 (N_16772,N_15860,N_15490);
nor U16773 (N_16773,N_15237,N_15605);
nor U16774 (N_16774,N_15774,N_15453);
or U16775 (N_16775,N_15856,N_15598);
nand U16776 (N_16776,N_15598,N_15783);
and U16777 (N_16777,N_15920,N_15878);
nand U16778 (N_16778,N_15493,N_15440);
nand U16779 (N_16779,N_15376,N_15493);
or U16780 (N_16780,N_15471,N_15566);
nor U16781 (N_16781,N_15502,N_15222);
nand U16782 (N_16782,N_15328,N_15534);
nor U16783 (N_16783,N_15898,N_15931);
or U16784 (N_16784,N_15579,N_15262);
nand U16785 (N_16785,N_15467,N_15456);
and U16786 (N_16786,N_15393,N_15256);
nand U16787 (N_16787,N_15733,N_15376);
xor U16788 (N_16788,N_15830,N_15275);
nor U16789 (N_16789,N_15831,N_15225);
nor U16790 (N_16790,N_15224,N_15431);
xor U16791 (N_16791,N_15549,N_15544);
or U16792 (N_16792,N_15554,N_15435);
xor U16793 (N_16793,N_15991,N_15845);
nor U16794 (N_16794,N_15538,N_15237);
nand U16795 (N_16795,N_15746,N_15443);
xor U16796 (N_16796,N_15683,N_15662);
or U16797 (N_16797,N_15212,N_15535);
and U16798 (N_16798,N_15366,N_15545);
xnor U16799 (N_16799,N_15448,N_15246);
nor U16800 (N_16800,N_16311,N_16762);
and U16801 (N_16801,N_16003,N_16739);
and U16802 (N_16802,N_16655,N_16179);
or U16803 (N_16803,N_16705,N_16691);
and U16804 (N_16804,N_16635,N_16005);
nand U16805 (N_16805,N_16356,N_16068);
xor U16806 (N_16806,N_16214,N_16359);
nor U16807 (N_16807,N_16141,N_16536);
and U16808 (N_16808,N_16095,N_16243);
or U16809 (N_16809,N_16551,N_16425);
and U16810 (N_16810,N_16046,N_16594);
or U16811 (N_16811,N_16184,N_16372);
nand U16812 (N_16812,N_16326,N_16454);
and U16813 (N_16813,N_16578,N_16297);
nor U16814 (N_16814,N_16440,N_16393);
or U16815 (N_16815,N_16302,N_16123);
nor U16816 (N_16816,N_16421,N_16265);
xnor U16817 (N_16817,N_16228,N_16798);
xnor U16818 (N_16818,N_16499,N_16301);
or U16819 (N_16819,N_16287,N_16185);
or U16820 (N_16820,N_16182,N_16759);
nor U16821 (N_16821,N_16677,N_16639);
xor U16822 (N_16822,N_16164,N_16782);
xnor U16823 (N_16823,N_16176,N_16659);
or U16824 (N_16824,N_16339,N_16065);
and U16825 (N_16825,N_16223,N_16405);
and U16826 (N_16826,N_16073,N_16155);
nand U16827 (N_16827,N_16006,N_16553);
nor U16828 (N_16828,N_16786,N_16709);
nor U16829 (N_16829,N_16037,N_16715);
or U16830 (N_16830,N_16617,N_16266);
xnor U16831 (N_16831,N_16253,N_16545);
nor U16832 (N_16832,N_16523,N_16396);
or U16833 (N_16833,N_16320,N_16699);
nand U16834 (N_16834,N_16186,N_16105);
nor U16835 (N_16835,N_16042,N_16055);
nand U16836 (N_16836,N_16284,N_16086);
nor U16837 (N_16837,N_16035,N_16247);
or U16838 (N_16838,N_16377,N_16525);
nand U16839 (N_16839,N_16118,N_16582);
nor U16840 (N_16840,N_16331,N_16272);
or U16841 (N_16841,N_16726,N_16215);
nor U16842 (N_16842,N_16570,N_16081);
xnor U16843 (N_16843,N_16328,N_16038);
or U16844 (N_16844,N_16506,N_16697);
nor U16845 (N_16845,N_16780,N_16651);
and U16846 (N_16846,N_16197,N_16262);
xor U16847 (N_16847,N_16261,N_16070);
and U16848 (N_16848,N_16758,N_16434);
xor U16849 (N_16849,N_16638,N_16391);
xnor U16850 (N_16850,N_16547,N_16381);
and U16851 (N_16851,N_16206,N_16059);
and U16852 (N_16852,N_16541,N_16149);
nand U16853 (N_16853,N_16652,N_16431);
or U16854 (N_16854,N_16244,N_16143);
nand U16855 (N_16855,N_16486,N_16604);
nor U16856 (N_16856,N_16676,N_16300);
and U16857 (N_16857,N_16057,N_16443);
and U16858 (N_16858,N_16294,N_16531);
nand U16859 (N_16859,N_16233,N_16724);
xnor U16860 (N_16860,N_16587,N_16279);
or U16861 (N_16861,N_16309,N_16508);
or U16862 (N_16862,N_16537,N_16448);
or U16863 (N_16863,N_16074,N_16213);
nand U16864 (N_16864,N_16111,N_16009);
and U16865 (N_16865,N_16256,N_16770);
nand U16866 (N_16866,N_16410,N_16636);
xnor U16867 (N_16867,N_16601,N_16245);
nor U16868 (N_16868,N_16568,N_16121);
and U16869 (N_16869,N_16529,N_16449);
or U16870 (N_16870,N_16656,N_16286);
or U16871 (N_16871,N_16765,N_16152);
nor U16872 (N_16872,N_16592,N_16004);
nand U16873 (N_16873,N_16110,N_16408);
nand U16874 (N_16874,N_16564,N_16530);
or U16875 (N_16875,N_16771,N_16079);
or U16876 (N_16876,N_16706,N_16390);
xnor U16877 (N_16877,N_16583,N_16389);
xnor U16878 (N_16878,N_16535,N_16360);
xor U16879 (N_16879,N_16465,N_16658);
or U16880 (N_16880,N_16435,N_16475);
nor U16881 (N_16881,N_16711,N_16554);
and U16882 (N_16882,N_16159,N_16542);
nand U16883 (N_16883,N_16384,N_16719);
nand U16884 (N_16884,N_16336,N_16533);
nand U16885 (N_16885,N_16364,N_16411);
xnor U16886 (N_16886,N_16313,N_16741);
nand U16887 (N_16887,N_16703,N_16281);
or U16888 (N_16888,N_16794,N_16716);
nand U16889 (N_16889,N_16365,N_16014);
and U16890 (N_16890,N_16464,N_16295);
and U16891 (N_16891,N_16382,N_16283);
nor U16892 (N_16892,N_16474,N_16264);
nor U16893 (N_16893,N_16188,N_16156);
nor U16894 (N_16894,N_16748,N_16373);
nand U16895 (N_16895,N_16512,N_16463);
and U16896 (N_16896,N_16028,N_16543);
or U16897 (N_16897,N_16608,N_16494);
nand U16898 (N_16898,N_16595,N_16227);
nor U16899 (N_16899,N_16787,N_16567);
and U16900 (N_16900,N_16493,N_16045);
nor U16901 (N_16901,N_16769,N_16694);
or U16902 (N_16902,N_16462,N_16238);
or U16903 (N_16903,N_16113,N_16199);
or U16904 (N_16904,N_16556,N_16240);
nor U16905 (N_16905,N_16062,N_16620);
xnor U16906 (N_16906,N_16161,N_16084);
and U16907 (N_16907,N_16735,N_16180);
nor U16908 (N_16908,N_16423,N_16456);
nand U16909 (N_16909,N_16054,N_16166);
nor U16910 (N_16910,N_16076,N_16598);
nor U16911 (N_16911,N_16733,N_16352);
and U16912 (N_16912,N_16222,N_16650);
and U16913 (N_16913,N_16109,N_16510);
xor U16914 (N_16914,N_16581,N_16366);
nor U16915 (N_16915,N_16312,N_16322);
nand U16916 (N_16916,N_16039,N_16544);
or U16917 (N_16917,N_16246,N_16497);
or U16918 (N_16918,N_16133,N_16024);
nor U16919 (N_16919,N_16496,N_16790);
and U16920 (N_16920,N_16696,N_16450);
or U16921 (N_16921,N_16093,N_16753);
and U16922 (N_16922,N_16387,N_16668);
nor U16923 (N_16923,N_16048,N_16096);
and U16924 (N_16924,N_16259,N_16460);
and U16925 (N_16925,N_16789,N_16168);
xnor U16926 (N_16926,N_16483,N_16693);
nor U16927 (N_16927,N_16707,N_16254);
nand U16928 (N_16928,N_16585,N_16056);
xnor U16929 (N_16929,N_16630,N_16632);
nand U16930 (N_16930,N_16341,N_16071);
or U16931 (N_16931,N_16346,N_16607);
nor U16932 (N_16932,N_16734,N_16532);
and U16933 (N_16933,N_16327,N_16783);
nand U16934 (N_16934,N_16157,N_16436);
nor U16935 (N_16935,N_16799,N_16094);
nand U16936 (N_16936,N_16670,N_16458);
nor U16937 (N_16937,N_16461,N_16701);
nand U16938 (N_16938,N_16522,N_16001);
and U16939 (N_16939,N_16649,N_16729);
or U16940 (N_16940,N_16692,N_16513);
nand U16941 (N_16941,N_16559,N_16280);
xnor U16942 (N_16942,N_16424,N_16178);
nor U16943 (N_16943,N_16731,N_16413);
or U16944 (N_16944,N_16170,N_16429);
nand U16945 (N_16945,N_16761,N_16713);
or U16946 (N_16946,N_16267,N_16679);
or U16947 (N_16947,N_16641,N_16018);
and U16948 (N_16948,N_16616,N_16172);
or U16949 (N_16949,N_16654,N_16471);
xor U16950 (N_16950,N_16369,N_16747);
nand U16951 (N_16951,N_16126,N_16211);
xnor U16952 (N_16952,N_16760,N_16402);
and U16953 (N_16953,N_16140,N_16127);
nor U16954 (N_16954,N_16666,N_16250);
and U16955 (N_16955,N_16566,N_16574);
or U16956 (N_16956,N_16524,N_16011);
nor U16957 (N_16957,N_16194,N_16628);
or U16958 (N_16958,N_16702,N_16200);
or U16959 (N_16959,N_16354,N_16257);
and U16960 (N_16960,N_16502,N_16316);
nand U16961 (N_16961,N_16190,N_16437);
nor U16962 (N_16962,N_16150,N_16438);
nand U16963 (N_16963,N_16067,N_16249);
xnor U16964 (N_16964,N_16509,N_16664);
xor U16965 (N_16965,N_16577,N_16239);
and U16966 (N_16966,N_16792,N_16293);
xor U16967 (N_16967,N_16130,N_16400);
nand U16968 (N_16968,N_16146,N_16773);
and U16969 (N_16969,N_16367,N_16100);
or U16970 (N_16970,N_16596,N_16204);
and U16971 (N_16971,N_16744,N_16277);
xor U16972 (N_16972,N_16646,N_16622);
nand U16973 (N_16973,N_16796,N_16298);
and U16974 (N_16974,N_16597,N_16021);
xor U16975 (N_16975,N_16064,N_16092);
xor U16976 (N_16976,N_16669,N_16348);
nand U16977 (N_16977,N_16428,N_16492);
nand U16978 (N_16978,N_16611,N_16218);
xnor U16979 (N_16979,N_16455,N_16198);
xnor U16980 (N_16980,N_16439,N_16593);
and U16981 (N_16981,N_16271,N_16767);
or U16982 (N_16982,N_16538,N_16351);
nor U16983 (N_16983,N_16645,N_16358);
or U16984 (N_16984,N_16777,N_16274);
nand U16985 (N_16985,N_16202,N_16647);
xnor U16986 (N_16986,N_16217,N_16040);
nand U16987 (N_16987,N_16128,N_16329);
or U16988 (N_16988,N_16340,N_16108);
or U16989 (N_16989,N_16047,N_16728);
and U16990 (N_16990,N_16337,N_16131);
xnor U16991 (N_16991,N_16539,N_16334);
xor U16992 (N_16992,N_16154,N_16169);
or U16993 (N_16993,N_16116,N_16484);
nor U16994 (N_16994,N_16629,N_16007);
nand U16995 (N_16995,N_16763,N_16485);
and U16996 (N_16996,N_16285,N_16335);
and U16997 (N_16997,N_16303,N_16732);
and U16998 (N_16998,N_16482,N_16229);
xnor U16999 (N_16999,N_16717,N_16690);
xnor U17000 (N_17000,N_16212,N_16778);
xor U17001 (N_17001,N_16114,N_16447);
and U17002 (N_17002,N_16451,N_16209);
or U17003 (N_17003,N_16386,N_16572);
nand U17004 (N_17004,N_16010,N_16569);
xor U17005 (N_17005,N_16314,N_16026);
xnor U17006 (N_17006,N_16764,N_16324);
or U17007 (N_17007,N_16241,N_16072);
nand U17008 (N_17008,N_16557,N_16580);
nor U17009 (N_17009,N_16627,N_16291);
and U17010 (N_17010,N_16338,N_16614);
or U17011 (N_17011,N_16260,N_16368);
nand U17012 (N_17012,N_16480,N_16251);
nand U17013 (N_17013,N_16151,N_16555);
or U17014 (N_17014,N_16099,N_16442);
and U17015 (N_17015,N_16528,N_16644);
xor U17016 (N_17016,N_16016,N_16220);
nand U17017 (N_17017,N_16549,N_16115);
nor U17018 (N_17018,N_16124,N_16195);
and U17019 (N_17019,N_16637,N_16603);
or U17020 (N_17020,N_16663,N_16061);
xor U17021 (N_17021,N_16002,N_16561);
xor U17022 (N_17022,N_16323,N_16681);
xor U17023 (N_17023,N_16210,N_16175);
and U17024 (N_17024,N_16602,N_16012);
nor U17025 (N_17025,N_16278,N_16615);
xnor U17026 (N_17026,N_16104,N_16671);
or U17027 (N_17027,N_16640,N_16708);
nor U17028 (N_17028,N_16224,N_16098);
and U17029 (N_17029,N_16634,N_16044);
and U17030 (N_17030,N_16565,N_16144);
or U17031 (N_17031,N_16342,N_16208);
xnor U17032 (N_17032,N_16344,N_16695);
nor U17033 (N_17033,N_16631,N_16772);
nand U17034 (N_17034,N_16147,N_16507);
xnor U17035 (N_17035,N_16562,N_16097);
nand U17036 (N_17036,N_16683,N_16017);
nand U17037 (N_17037,N_16307,N_16625);
nor U17038 (N_17038,N_16605,N_16091);
and U17039 (N_17039,N_16743,N_16416);
nor U17040 (N_17040,N_16505,N_16310);
xnor U17041 (N_17041,N_16174,N_16165);
xnor U17042 (N_17042,N_16576,N_16672);
xnor U17043 (N_17043,N_16397,N_16720);
and U17044 (N_17044,N_16621,N_16432);
nand U17045 (N_17045,N_16299,N_16504);
nor U17046 (N_17046,N_16457,N_16183);
or U17047 (N_17047,N_16090,N_16000);
nor U17048 (N_17048,N_16306,N_16153);
or U17049 (N_17049,N_16361,N_16022);
xor U17050 (N_17050,N_16469,N_16350);
nand U17051 (N_17051,N_16452,N_16112);
nand U17052 (N_17052,N_16371,N_16343);
and U17053 (N_17053,N_16558,N_16579);
and U17054 (N_17054,N_16653,N_16201);
xor U17055 (N_17055,N_16318,N_16242);
and U17056 (N_17056,N_16521,N_16275);
xor U17057 (N_17057,N_16129,N_16103);
and U17058 (N_17058,N_16078,N_16205);
and U17059 (N_17059,N_16586,N_16685);
and U17060 (N_17060,N_16252,N_16473);
and U17061 (N_17061,N_16445,N_16173);
or U17062 (N_17062,N_16714,N_16606);
and U17063 (N_17063,N_16526,N_16467);
nor U17064 (N_17064,N_16591,N_16025);
nor U17065 (N_17065,N_16036,N_16219);
xnor U17066 (N_17066,N_16441,N_16347);
nor U17067 (N_17067,N_16476,N_16148);
xnor U17068 (N_17068,N_16137,N_16643);
nand U17069 (N_17069,N_16730,N_16612);
xnor U17070 (N_17070,N_16418,N_16687);
nand U17071 (N_17071,N_16119,N_16563);
nor U17072 (N_17072,N_16237,N_16053);
and U17073 (N_17073,N_16321,N_16230);
xnor U17074 (N_17074,N_16013,N_16468);
or U17075 (N_17075,N_16134,N_16378);
nor U17076 (N_17076,N_16050,N_16120);
and U17077 (N_17077,N_16742,N_16791);
xor U17078 (N_17078,N_16495,N_16375);
or U17079 (N_17079,N_16718,N_16355);
xor U17080 (N_17080,N_16756,N_16041);
nand U17081 (N_17081,N_16752,N_16374);
nor U17082 (N_17082,N_16019,N_16427);
xor U17083 (N_17083,N_16160,N_16162);
or U17084 (N_17084,N_16399,N_16258);
or U17085 (N_17085,N_16409,N_16737);
or U17086 (N_17086,N_16498,N_16226);
or U17087 (N_17087,N_16033,N_16776);
nor U17088 (N_17088,N_16043,N_16269);
and U17089 (N_17089,N_16534,N_16422);
and U17090 (N_17090,N_16785,N_16135);
nor U17091 (N_17091,N_16122,N_16308);
and U17092 (N_17092,N_16305,N_16385);
and U17093 (N_17093,N_16546,N_16420);
xor U17094 (N_17094,N_16029,N_16296);
or U17095 (N_17095,N_16414,N_16618);
and U17096 (N_17096,N_16478,N_16191);
nor U17097 (N_17097,N_16665,N_16500);
or U17098 (N_17098,N_16139,N_16477);
nor U17099 (N_17099,N_16797,N_16087);
or U17100 (N_17100,N_16345,N_16270);
nand U17101 (N_17101,N_16330,N_16779);
or U17102 (N_17102,N_16725,N_16633);
nand U17103 (N_17103,N_16030,N_16203);
or U17104 (N_17104,N_16698,N_16721);
nand U17105 (N_17105,N_16590,N_16489);
and U17106 (N_17106,N_16610,N_16793);
xor U17107 (N_17107,N_16487,N_16584);
or U17108 (N_17108,N_16282,N_16704);
nand U17109 (N_17109,N_16349,N_16187);
xor U17110 (N_17110,N_16395,N_16207);
nand U17111 (N_17111,N_16503,N_16406);
or U17112 (N_17112,N_16540,N_16795);
nand U17113 (N_17113,N_16077,N_16231);
xor U17114 (N_17114,N_16234,N_16740);
nor U17115 (N_17115,N_16255,N_16479);
xnor U17116 (N_17116,N_16117,N_16063);
or U17117 (N_17117,N_16723,N_16774);
and U17118 (N_17118,N_16216,N_16700);
nor U17119 (N_17119,N_16514,N_16276);
nor U17120 (N_17120,N_16660,N_16749);
nor U17121 (N_17121,N_16020,N_16289);
or U17122 (N_17122,N_16268,N_16727);
nor U17123 (N_17123,N_16027,N_16686);
and U17124 (N_17124,N_16662,N_16520);
and U17125 (N_17125,N_16383,N_16192);
or U17126 (N_17126,N_16689,N_16550);
xnor U17127 (N_17127,N_16088,N_16755);
nand U17128 (N_17128,N_16225,N_16023);
and U17129 (N_17129,N_16158,N_16781);
and U17130 (N_17130,N_16142,N_16221);
nand U17131 (N_17131,N_16106,N_16031);
or U17132 (N_17132,N_16325,N_16710);
and U17133 (N_17133,N_16235,N_16332);
nand U17134 (N_17134,N_16459,N_16052);
nor U17135 (N_17135,N_16273,N_16642);
nand U17136 (N_17136,N_16015,N_16069);
or U17137 (N_17137,N_16398,N_16125);
nor U17138 (N_17138,N_16136,N_16599);
and U17139 (N_17139,N_16472,N_16470);
nand U17140 (N_17140,N_16722,N_16145);
nand U17141 (N_17141,N_16080,N_16560);
or U17142 (N_17142,N_16589,N_16518);
or U17143 (N_17143,N_16600,N_16075);
nand U17144 (N_17144,N_16626,N_16315);
nand U17145 (N_17145,N_16661,N_16193);
xnor U17146 (N_17146,N_16304,N_16682);
or U17147 (N_17147,N_16688,N_16138);
or U17148 (N_17148,N_16673,N_16353);
xor U17149 (N_17149,N_16446,N_16588);
and U17150 (N_17150,N_16788,N_16177);
xnor U17151 (N_17151,N_16667,N_16571);
or U17152 (N_17152,N_16674,N_16394);
nand U17153 (N_17153,N_16426,N_16049);
nor U17154 (N_17154,N_16527,N_16388);
and U17155 (N_17155,N_16575,N_16548);
nand U17156 (N_17156,N_16712,N_16236);
nand U17157 (N_17157,N_16552,N_16609);
or U17158 (N_17158,N_16619,N_16613);
or U17159 (N_17159,N_16370,N_16511);
and U17160 (N_17160,N_16519,N_16417);
or U17161 (N_17161,N_16404,N_16380);
xor U17162 (N_17162,N_16032,N_16263);
xnor U17163 (N_17163,N_16624,N_16768);
xnor U17164 (N_17164,N_16684,N_16766);
nand U17165 (N_17165,N_16680,N_16444);
xor U17166 (N_17166,N_16648,N_16196);
or U17167 (N_17167,N_16317,N_16034);
and U17168 (N_17168,N_16060,N_16491);
xnor U17169 (N_17169,N_16623,N_16171);
nor U17170 (N_17170,N_16466,N_16738);
nor U17171 (N_17171,N_16501,N_16517);
and U17172 (N_17172,N_16403,N_16132);
or U17173 (N_17173,N_16379,N_16101);
nor U17174 (N_17174,N_16751,N_16784);
nor U17175 (N_17175,N_16736,N_16319);
nor U17176 (N_17176,N_16357,N_16163);
and U17177 (N_17177,N_16678,N_16376);
xor U17178 (N_17178,N_16083,N_16189);
xor U17179 (N_17179,N_16290,N_16051);
nor U17180 (N_17180,N_16515,N_16453);
and U17181 (N_17181,N_16775,N_16490);
nand U17182 (N_17182,N_16082,N_16066);
nand U17183 (N_17183,N_16362,N_16573);
xor U17184 (N_17184,N_16745,N_16433);
nor U17185 (N_17185,N_16754,N_16657);
and U17186 (N_17186,N_16419,N_16333);
xor U17187 (N_17187,N_16488,N_16415);
xor U17188 (N_17188,N_16008,N_16430);
nor U17189 (N_17189,N_16167,N_16746);
xor U17190 (N_17190,N_16058,N_16412);
and U17191 (N_17191,N_16675,N_16392);
nor U17192 (N_17192,N_16750,N_16102);
or U17193 (N_17193,N_16232,N_16292);
nand U17194 (N_17194,N_16757,N_16288);
nor U17195 (N_17195,N_16363,N_16516);
and U17196 (N_17196,N_16085,N_16407);
and U17197 (N_17197,N_16107,N_16481);
nor U17198 (N_17198,N_16401,N_16248);
xor U17199 (N_17199,N_16089,N_16181);
xnor U17200 (N_17200,N_16692,N_16741);
or U17201 (N_17201,N_16400,N_16157);
nand U17202 (N_17202,N_16497,N_16762);
nand U17203 (N_17203,N_16701,N_16531);
nor U17204 (N_17204,N_16385,N_16628);
and U17205 (N_17205,N_16345,N_16032);
xnor U17206 (N_17206,N_16427,N_16784);
and U17207 (N_17207,N_16257,N_16170);
xnor U17208 (N_17208,N_16033,N_16605);
nand U17209 (N_17209,N_16485,N_16059);
and U17210 (N_17210,N_16340,N_16429);
nor U17211 (N_17211,N_16236,N_16616);
nor U17212 (N_17212,N_16520,N_16424);
and U17213 (N_17213,N_16053,N_16548);
and U17214 (N_17214,N_16301,N_16138);
nor U17215 (N_17215,N_16129,N_16556);
xnor U17216 (N_17216,N_16584,N_16036);
nor U17217 (N_17217,N_16009,N_16547);
and U17218 (N_17218,N_16314,N_16757);
or U17219 (N_17219,N_16211,N_16604);
nor U17220 (N_17220,N_16101,N_16755);
nor U17221 (N_17221,N_16018,N_16746);
or U17222 (N_17222,N_16462,N_16129);
and U17223 (N_17223,N_16460,N_16589);
and U17224 (N_17224,N_16622,N_16398);
or U17225 (N_17225,N_16604,N_16197);
nor U17226 (N_17226,N_16204,N_16488);
nor U17227 (N_17227,N_16750,N_16354);
and U17228 (N_17228,N_16690,N_16133);
xor U17229 (N_17229,N_16366,N_16671);
xnor U17230 (N_17230,N_16773,N_16077);
or U17231 (N_17231,N_16422,N_16614);
nand U17232 (N_17232,N_16414,N_16334);
nor U17233 (N_17233,N_16054,N_16488);
xor U17234 (N_17234,N_16584,N_16352);
or U17235 (N_17235,N_16301,N_16324);
xor U17236 (N_17236,N_16544,N_16376);
and U17237 (N_17237,N_16360,N_16626);
xor U17238 (N_17238,N_16109,N_16555);
or U17239 (N_17239,N_16531,N_16642);
or U17240 (N_17240,N_16178,N_16185);
xor U17241 (N_17241,N_16533,N_16664);
and U17242 (N_17242,N_16244,N_16523);
xor U17243 (N_17243,N_16374,N_16047);
and U17244 (N_17244,N_16081,N_16509);
nor U17245 (N_17245,N_16780,N_16014);
and U17246 (N_17246,N_16185,N_16656);
nor U17247 (N_17247,N_16177,N_16275);
nor U17248 (N_17248,N_16108,N_16281);
and U17249 (N_17249,N_16399,N_16702);
nor U17250 (N_17250,N_16101,N_16266);
and U17251 (N_17251,N_16205,N_16717);
nand U17252 (N_17252,N_16498,N_16617);
and U17253 (N_17253,N_16045,N_16116);
nor U17254 (N_17254,N_16645,N_16655);
and U17255 (N_17255,N_16784,N_16152);
and U17256 (N_17256,N_16336,N_16029);
xor U17257 (N_17257,N_16106,N_16085);
or U17258 (N_17258,N_16236,N_16762);
and U17259 (N_17259,N_16119,N_16438);
or U17260 (N_17260,N_16580,N_16667);
nor U17261 (N_17261,N_16562,N_16471);
nor U17262 (N_17262,N_16156,N_16711);
xnor U17263 (N_17263,N_16401,N_16151);
and U17264 (N_17264,N_16307,N_16784);
nand U17265 (N_17265,N_16606,N_16021);
xor U17266 (N_17266,N_16485,N_16325);
xor U17267 (N_17267,N_16373,N_16309);
xnor U17268 (N_17268,N_16349,N_16109);
or U17269 (N_17269,N_16151,N_16769);
nand U17270 (N_17270,N_16397,N_16206);
nor U17271 (N_17271,N_16218,N_16397);
xor U17272 (N_17272,N_16271,N_16352);
nand U17273 (N_17273,N_16537,N_16391);
nor U17274 (N_17274,N_16787,N_16284);
nor U17275 (N_17275,N_16335,N_16405);
and U17276 (N_17276,N_16214,N_16445);
xnor U17277 (N_17277,N_16544,N_16017);
nor U17278 (N_17278,N_16102,N_16515);
nand U17279 (N_17279,N_16083,N_16261);
and U17280 (N_17280,N_16020,N_16285);
xnor U17281 (N_17281,N_16578,N_16171);
xnor U17282 (N_17282,N_16365,N_16160);
xor U17283 (N_17283,N_16639,N_16598);
nand U17284 (N_17284,N_16689,N_16667);
xor U17285 (N_17285,N_16397,N_16280);
and U17286 (N_17286,N_16498,N_16710);
nand U17287 (N_17287,N_16152,N_16557);
or U17288 (N_17288,N_16070,N_16740);
nor U17289 (N_17289,N_16481,N_16505);
nand U17290 (N_17290,N_16073,N_16444);
and U17291 (N_17291,N_16354,N_16744);
xnor U17292 (N_17292,N_16025,N_16176);
or U17293 (N_17293,N_16628,N_16783);
xnor U17294 (N_17294,N_16661,N_16555);
and U17295 (N_17295,N_16042,N_16129);
nand U17296 (N_17296,N_16702,N_16715);
or U17297 (N_17297,N_16135,N_16271);
or U17298 (N_17298,N_16600,N_16029);
nor U17299 (N_17299,N_16283,N_16410);
nor U17300 (N_17300,N_16643,N_16618);
or U17301 (N_17301,N_16407,N_16764);
xor U17302 (N_17302,N_16211,N_16174);
and U17303 (N_17303,N_16148,N_16043);
nor U17304 (N_17304,N_16648,N_16556);
or U17305 (N_17305,N_16733,N_16604);
and U17306 (N_17306,N_16575,N_16428);
and U17307 (N_17307,N_16681,N_16594);
nand U17308 (N_17308,N_16671,N_16045);
xor U17309 (N_17309,N_16621,N_16280);
and U17310 (N_17310,N_16270,N_16604);
xor U17311 (N_17311,N_16681,N_16488);
nand U17312 (N_17312,N_16389,N_16446);
or U17313 (N_17313,N_16342,N_16222);
xor U17314 (N_17314,N_16504,N_16326);
nor U17315 (N_17315,N_16307,N_16694);
xnor U17316 (N_17316,N_16019,N_16548);
and U17317 (N_17317,N_16401,N_16049);
or U17318 (N_17318,N_16203,N_16388);
xnor U17319 (N_17319,N_16148,N_16212);
or U17320 (N_17320,N_16676,N_16727);
or U17321 (N_17321,N_16117,N_16551);
nand U17322 (N_17322,N_16050,N_16204);
and U17323 (N_17323,N_16177,N_16280);
and U17324 (N_17324,N_16688,N_16611);
nand U17325 (N_17325,N_16695,N_16518);
and U17326 (N_17326,N_16604,N_16665);
nor U17327 (N_17327,N_16689,N_16799);
nor U17328 (N_17328,N_16187,N_16164);
xor U17329 (N_17329,N_16037,N_16591);
nand U17330 (N_17330,N_16752,N_16128);
nor U17331 (N_17331,N_16307,N_16334);
or U17332 (N_17332,N_16625,N_16478);
nand U17333 (N_17333,N_16672,N_16385);
or U17334 (N_17334,N_16039,N_16175);
or U17335 (N_17335,N_16411,N_16193);
nand U17336 (N_17336,N_16672,N_16087);
nor U17337 (N_17337,N_16210,N_16406);
xor U17338 (N_17338,N_16650,N_16678);
or U17339 (N_17339,N_16510,N_16514);
and U17340 (N_17340,N_16232,N_16100);
nor U17341 (N_17341,N_16571,N_16340);
nand U17342 (N_17342,N_16738,N_16303);
nand U17343 (N_17343,N_16233,N_16430);
nand U17344 (N_17344,N_16432,N_16017);
and U17345 (N_17345,N_16140,N_16004);
xor U17346 (N_17346,N_16582,N_16029);
nor U17347 (N_17347,N_16201,N_16620);
nand U17348 (N_17348,N_16321,N_16430);
nand U17349 (N_17349,N_16453,N_16701);
xnor U17350 (N_17350,N_16041,N_16765);
nor U17351 (N_17351,N_16316,N_16681);
nor U17352 (N_17352,N_16000,N_16283);
xnor U17353 (N_17353,N_16398,N_16700);
or U17354 (N_17354,N_16038,N_16342);
or U17355 (N_17355,N_16251,N_16051);
xnor U17356 (N_17356,N_16416,N_16432);
or U17357 (N_17357,N_16712,N_16761);
nand U17358 (N_17358,N_16694,N_16780);
nand U17359 (N_17359,N_16226,N_16780);
nor U17360 (N_17360,N_16759,N_16553);
nand U17361 (N_17361,N_16756,N_16108);
and U17362 (N_17362,N_16291,N_16350);
nor U17363 (N_17363,N_16129,N_16039);
or U17364 (N_17364,N_16489,N_16647);
nor U17365 (N_17365,N_16789,N_16776);
and U17366 (N_17366,N_16275,N_16683);
and U17367 (N_17367,N_16103,N_16691);
nor U17368 (N_17368,N_16307,N_16646);
nand U17369 (N_17369,N_16167,N_16491);
and U17370 (N_17370,N_16470,N_16293);
or U17371 (N_17371,N_16344,N_16379);
xor U17372 (N_17372,N_16008,N_16023);
nor U17373 (N_17373,N_16085,N_16504);
nand U17374 (N_17374,N_16132,N_16668);
xnor U17375 (N_17375,N_16684,N_16120);
xor U17376 (N_17376,N_16430,N_16220);
or U17377 (N_17377,N_16209,N_16059);
or U17378 (N_17378,N_16205,N_16778);
nor U17379 (N_17379,N_16622,N_16012);
or U17380 (N_17380,N_16604,N_16660);
nor U17381 (N_17381,N_16575,N_16707);
nand U17382 (N_17382,N_16112,N_16246);
xnor U17383 (N_17383,N_16488,N_16203);
xnor U17384 (N_17384,N_16538,N_16161);
xnor U17385 (N_17385,N_16360,N_16703);
and U17386 (N_17386,N_16263,N_16571);
or U17387 (N_17387,N_16582,N_16578);
xnor U17388 (N_17388,N_16723,N_16494);
nand U17389 (N_17389,N_16573,N_16279);
nor U17390 (N_17390,N_16018,N_16137);
xnor U17391 (N_17391,N_16286,N_16348);
xnor U17392 (N_17392,N_16266,N_16222);
or U17393 (N_17393,N_16518,N_16593);
nor U17394 (N_17394,N_16182,N_16350);
xnor U17395 (N_17395,N_16703,N_16211);
nand U17396 (N_17396,N_16757,N_16712);
xor U17397 (N_17397,N_16650,N_16721);
nand U17398 (N_17398,N_16309,N_16778);
nand U17399 (N_17399,N_16299,N_16750);
xor U17400 (N_17400,N_16410,N_16572);
or U17401 (N_17401,N_16254,N_16301);
nand U17402 (N_17402,N_16502,N_16338);
and U17403 (N_17403,N_16393,N_16047);
nand U17404 (N_17404,N_16420,N_16555);
or U17405 (N_17405,N_16403,N_16108);
nor U17406 (N_17406,N_16305,N_16417);
nor U17407 (N_17407,N_16577,N_16711);
or U17408 (N_17408,N_16223,N_16463);
nor U17409 (N_17409,N_16700,N_16459);
xnor U17410 (N_17410,N_16601,N_16702);
nor U17411 (N_17411,N_16320,N_16072);
xor U17412 (N_17412,N_16278,N_16028);
xor U17413 (N_17413,N_16644,N_16432);
nand U17414 (N_17414,N_16018,N_16748);
or U17415 (N_17415,N_16438,N_16726);
nor U17416 (N_17416,N_16343,N_16040);
and U17417 (N_17417,N_16754,N_16213);
nor U17418 (N_17418,N_16711,N_16455);
xnor U17419 (N_17419,N_16115,N_16745);
or U17420 (N_17420,N_16214,N_16494);
nand U17421 (N_17421,N_16608,N_16057);
or U17422 (N_17422,N_16756,N_16070);
xnor U17423 (N_17423,N_16091,N_16248);
xor U17424 (N_17424,N_16757,N_16787);
xor U17425 (N_17425,N_16791,N_16710);
xnor U17426 (N_17426,N_16109,N_16475);
and U17427 (N_17427,N_16520,N_16099);
nor U17428 (N_17428,N_16173,N_16179);
nor U17429 (N_17429,N_16411,N_16229);
nor U17430 (N_17430,N_16427,N_16219);
nand U17431 (N_17431,N_16460,N_16177);
and U17432 (N_17432,N_16019,N_16476);
or U17433 (N_17433,N_16468,N_16491);
or U17434 (N_17434,N_16038,N_16691);
or U17435 (N_17435,N_16006,N_16013);
nor U17436 (N_17436,N_16500,N_16144);
or U17437 (N_17437,N_16486,N_16427);
xor U17438 (N_17438,N_16104,N_16341);
nor U17439 (N_17439,N_16355,N_16444);
xor U17440 (N_17440,N_16354,N_16234);
or U17441 (N_17441,N_16267,N_16414);
xor U17442 (N_17442,N_16446,N_16441);
nand U17443 (N_17443,N_16784,N_16396);
xor U17444 (N_17444,N_16649,N_16460);
or U17445 (N_17445,N_16027,N_16205);
nor U17446 (N_17446,N_16208,N_16191);
nor U17447 (N_17447,N_16148,N_16182);
nor U17448 (N_17448,N_16524,N_16127);
nor U17449 (N_17449,N_16040,N_16728);
or U17450 (N_17450,N_16140,N_16597);
xnor U17451 (N_17451,N_16250,N_16396);
nor U17452 (N_17452,N_16047,N_16681);
nand U17453 (N_17453,N_16047,N_16532);
nand U17454 (N_17454,N_16749,N_16310);
xnor U17455 (N_17455,N_16742,N_16431);
nor U17456 (N_17456,N_16399,N_16072);
xnor U17457 (N_17457,N_16714,N_16204);
nor U17458 (N_17458,N_16245,N_16199);
xor U17459 (N_17459,N_16673,N_16235);
nor U17460 (N_17460,N_16562,N_16022);
nand U17461 (N_17461,N_16423,N_16602);
nand U17462 (N_17462,N_16497,N_16695);
and U17463 (N_17463,N_16728,N_16637);
nor U17464 (N_17464,N_16311,N_16683);
nand U17465 (N_17465,N_16099,N_16588);
xnor U17466 (N_17466,N_16389,N_16077);
xnor U17467 (N_17467,N_16742,N_16376);
and U17468 (N_17468,N_16299,N_16011);
nand U17469 (N_17469,N_16648,N_16531);
nor U17470 (N_17470,N_16200,N_16607);
nand U17471 (N_17471,N_16280,N_16333);
or U17472 (N_17472,N_16781,N_16767);
or U17473 (N_17473,N_16172,N_16184);
nor U17474 (N_17474,N_16453,N_16652);
nand U17475 (N_17475,N_16181,N_16039);
or U17476 (N_17476,N_16106,N_16016);
nor U17477 (N_17477,N_16426,N_16153);
or U17478 (N_17478,N_16547,N_16280);
xnor U17479 (N_17479,N_16282,N_16532);
xnor U17480 (N_17480,N_16396,N_16720);
xor U17481 (N_17481,N_16637,N_16161);
xor U17482 (N_17482,N_16119,N_16332);
xnor U17483 (N_17483,N_16424,N_16157);
or U17484 (N_17484,N_16187,N_16308);
nor U17485 (N_17485,N_16767,N_16358);
xor U17486 (N_17486,N_16249,N_16240);
xnor U17487 (N_17487,N_16434,N_16331);
and U17488 (N_17488,N_16394,N_16768);
or U17489 (N_17489,N_16020,N_16258);
nor U17490 (N_17490,N_16378,N_16483);
or U17491 (N_17491,N_16704,N_16397);
nand U17492 (N_17492,N_16758,N_16645);
xor U17493 (N_17493,N_16652,N_16251);
xnor U17494 (N_17494,N_16743,N_16770);
and U17495 (N_17495,N_16110,N_16782);
nand U17496 (N_17496,N_16647,N_16665);
and U17497 (N_17497,N_16426,N_16524);
xnor U17498 (N_17498,N_16420,N_16139);
xnor U17499 (N_17499,N_16435,N_16404);
nor U17500 (N_17500,N_16397,N_16392);
nor U17501 (N_17501,N_16246,N_16634);
and U17502 (N_17502,N_16433,N_16524);
xor U17503 (N_17503,N_16243,N_16386);
xnor U17504 (N_17504,N_16403,N_16541);
and U17505 (N_17505,N_16646,N_16342);
xnor U17506 (N_17506,N_16679,N_16698);
xor U17507 (N_17507,N_16618,N_16334);
and U17508 (N_17508,N_16400,N_16055);
nand U17509 (N_17509,N_16241,N_16600);
xor U17510 (N_17510,N_16060,N_16332);
and U17511 (N_17511,N_16270,N_16376);
and U17512 (N_17512,N_16471,N_16304);
nor U17513 (N_17513,N_16195,N_16201);
nor U17514 (N_17514,N_16662,N_16340);
nor U17515 (N_17515,N_16701,N_16728);
xor U17516 (N_17516,N_16396,N_16786);
and U17517 (N_17517,N_16521,N_16173);
nor U17518 (N_17518,N_16702,N_16240);
nand U17519 (N_17519,N_16594,N_16158);
nand U17520 (N_17520,N_16442,N_16702);
and U17521 (N_17521,N_16381,N_16451);
nand U17522 (N_17522,N_16047,N_16675);
and U17523 (N_17523,N_16755,N_16131);
or U17524 (N_17524,N_16446,N_16275);
nor U17525 (N_17525,N_16261,N_16026);
xor U17526 (N_17526,N_16515,N_16606);
nor U17527 (N_17527,N_16036,N_16459);
nor U17528 (N_17528,N_16671,N_16728);
xor U17529 (N_17529,N_16238,N_16426);
nor U17530 (N_17530,N_16515,N_16342);
or U17531 (N_17531,N_16352,N_16010);
or U17532 (N_17532,N_16141,N_16003);
or U17533 (N_17533,N_16617,N_16113);
and U17534 (N_17534,N_16207,N_16549);
xnor U17535 (N_17535,N_16599,N_16543);
and U17536 (N_17536,N_16544,N_16560);
xnor U17537 (N_17537,N_16792,N_16067);
or U17538 (N_17538,N_16513,N_16413);
nand U17539 (N_17539,N_16511,N_16556);
and U17540 (N_17540,N_16445,N_16653);
nand U17541 (N_17541,N_16770,N_16479);
or U17542 (N_17542,N_16524,N_16272);
nor U17543 (N_17543,N_16366,N_16750);
and U17544 (N_17544,N_16423,N_16685);
and U17545 (N_17545,N_16360,N_16304);
nand U17546 (N_17546,N_16519,N_16437);
or U17547 (N_17547,N_16061,N_16126);
nor U17548 (N_17548,N_16065,N_16722);
nand U17549 (N_17549,N_16109,N_16219);
nand U17550 (N_17550,N_16589,N_16763);
or U17551 (N_17551,N_16167,N_16156);
and U17552 (N_17552,N_16013,N_16231);
or U17553 (N_17553,N_16059,N_16365);
or U17554 (N_17554,N_16091,N_16011);
xor U17555 (N_17555,N_16355,N_16507);
and U17556 (N_17556,N_16309,N_16500);
or U17557 (N_17557,N_16575,N_16576);
nor U17558 (N_17558,N_16525,N_16291);
nor U17559 (N_17559,N_16614,N_16533);
nand U17560 (N_17560,N_16020,N_16759);
and U17561 (N_17561,N_16317,N_16798);
nor U17562 (N_17562,N_16407,N_16403);
or U17563 (N_17563,N_16270,N_16321);
nor U17564 (N_17564,N_16137,N_16165);
xnor U17565 (N_17565,N_16356,N_16685);
nor U17566 (N_17566,N_16601,N_16621);
or U17567 (N_17567,N_16587,N_16048);
nand U17568 (N_17568,N_16144,N_16334);
nor U17569 (N_17569,N_16580,N_16300);
or U17570 (N_17570,N_16175,N_16196);
nor U17571 (N_17571,N_16635,N_16072);
nand U17572 (N_17572,N_16710,N_16453);
nand U17573 (N_17573,N_16181,N_16288);
nand U17574 (N_17574,N_16295,N_16451);
xnor U17575 (N_17575,N_16673,N_16687);
and U17576 (N_17576,N_16355,N_16002);
nor U17577 (N_17577,N_16232,N_16278);
or U17578 (N_17578,N_16180,N_16218);
nor U17579 (N_17579,N_16141,N_16066);
and U17580 (N_17580,N_16261,N_16598);
nand U17581 (N_17581,N_16504,N_16205);
nand U17582 (N_17582,N_16120,N_16754);
nor U17583 (N_17583,N_16359,N_16710);
nor U17584 (N_17584,N_16614,N_16643);
xor U17585 (N_17585,N_16359,N_16797);
and U17586 (N_17586,N_16688,N_16490);
and U17587 (N_17587,N_16536,N_16787);
or U17588 (N_17588,N_16575,N_16107);
and U17589 (N_17589,N_16397,N_16697);
nor U17590 (N_17590,N_16740,N_16299);
nand U17591 (N_17591,N_16321,N_16701);
or U17592 (N_17592,N_16478,N_16495);
xor U17593 (N_17593,N_16353,N_16607);
and U17594 (N_17594,N_16594,N_16012);
nor U17595 (N_17595,N_16771,N_16340);
and U17596 (N_17596,N_16552,N_16689);
nand U17597 (N_17597,N_16174,N_16036);
nand U17598 (N_17598,N_16214,N_16071);
xnor U17599 (N_17599,N_16347,N_16019);
nor U17600 (N_17600,N_17119,N_17194);
nand U17601 (N_17601,N_17259,N_17570);
or U17602 (N_17602,N_17041,N_17391);
nor U17603 (N_17603,N_17014,N_16982);
nand U17604 (N_17604,N_17139,N_17242);
nor U17605 (N_17605,N_17438,N_17267);
or U17606 (N_17606,N_16936,N_16870);
xor U17607 (N_17607,N_16903,N_17284);
and U17608 (N_17608,N_17311,N_17271);
nor U17609 (N_17609,N_17038,N_17401);
or U17610 (N_17610,N_17136,N_17204);
or U17611 (N_17611,N_17441,N_17214);
and U17612 (N_17612,N_17247,N_16845);
and U17613 (N_17613,N_16897,N_17431);
xor U17614 (N_17614,N_17081,N_17013);
nor U17615 (N_17615,N_17053,N_16875);
and U17616 (N_17616,N_17416,N_17168);
nand U17617 (N_17617,N_16872,N_16850);
nand U17618 (N_17618,N_16843,N_17043);
nand U17619 (N_17619,N_17412,N_17051);
nand U17620 (N_17620,N_17140,N_17518);
or U17621 (N_17621,N_17274,N_16917);
xnor U17622 (N_17622,N_16827,N_17358);
and U17623 (N_17623,N_17147,N_17521);
and U17624 (N_17624,N_16995,N_17221);
nor U17625 (N_17625,N_17086,N_17200);
and U17626 (N_17626,N_17548,N_17135);
nor U17627 (N_17627,N_17579,N_17451);
xor U17628 (N_17628,N_16853,N_17343);
nor U17629 (N_17629,N_17179,N_17505);
xnor U17630 (N_17630,N_16987,N_17459);
and U17631 (N_17631,N_17103,N_17535);
xor U17632 (N_17632,N_17035,N_17496);
nor U17633 (N_17633,N_17527,N_16841);
or U17634 (N_17634,N_17529,N_17489);
and U17635 (N_17635,N_17449,N_17209);
nor U17636 (N_17636,N_17185,N_17159);
nand U17637 (N_17637,N_17359,N_17062);
and U17638 (N_17638,N_17127,N_16898);
or U17639 (N_17639,N_17260,N_17215);
nand U17640 (N_17640,N_16918,N_17387);
and U17641 (N_17641,N_17249,N_17004);
nand U17642 (N_17642,N_17161,N_16964);
xor U17643 (N_17643,N_16913,N_17021);
xor U17644 (N_17644,N_17300,N_17094);
xnor U17645 (N_17645,N_17526,N_17181);
nand U17646 (N_17646,N_17176,N_16900);
nor U17647 (N_17647,N_16858,N_17379);
nand U17648 (N_17648,N_16905,N_17054);
nor U17649 (N_17649,N_17167,N_17129);
or U17650 (N_17650,N_17314,N_17039);
xnor U17651 (N_17651,N_17533,N_17323);
nor U17652 (N_17652,N_17225,N_17205);
nor U17653 (N_17653,N_17195,N_17301);
or U17654 (N_17654,N_17375,N_17130);
or U17655 (N_17655,N_17506,N_17228);
nand U17656 (N_17656,N_17405,N_17131);
or U17657 (N_17657,N_17487,N_17397);
xnor U17658 (N_17658,N_16868,N_17490);
nor U17659 (N_17659,N_17120,N_17297);
nand U17660 (N_17660,N_16819,N_16941);
or U17661 (N_17661,N_17427,N_17188);
xnor U17662 (N_17662,N_17085,N_17462);
and U17663 (N_17663,N_16974,N_17166);
nand U17664 (N_17664,N_17403,N_17395);
and U17665 (N_17665,N_17097,N_16828);
nand U17666 (N_17666,N_17572,N_17281);
nor U17667 (N_17667,N_17530,N_17546);
nand U17668 (N_17668,N_17163,N_16834);
xor U17669 (N_17669,N_16867,N_17025);
nand U17670 (N_17670,N_17101,N_17138);
xor U17671 (N_17671,N_16957,N_17160);
and U17672 (N_17672,N_17588,N_17315);
or U17673 (N_17673,N_17580,N_16908);
nand U17674 (N_17674,N_16857,N_16915);
and U17675 (N_17675,N_17199,N_16817);
or U17676 (N_17676,N_16979,N_17132);
nor U17677 (N_17677,N_16876,N_17146);
and U17678 (N_17678,N_16919,N_17393);
nor U17679 (N_17679,N_17059,N_17589);
xor U17680 (N_17680,N_17440,N_17360);
nand U17681 (N_17681,N_17118,N_17364);
nor U17682 (N_17682,N_16971,N_17348);
nand U17683 (N_17683,N_17476,N_17007);
or U17684 (N_17684,N_17064,N_17443);
xnor U17685 (N_17685,N_17394,N_17374);
nor U17686 (N_17686,N_17574,N_16986);
and U17687 (N_17687,N_17210,N_17563);
nand U17688 (N_17688,N_17015,N_16985);
xor U17689 (N_17689,N_16928,N_16849);
xnor U17690 (N_17690,N_16840,N_16992);
nand U17691 (N_17691,N_17218,N_17034);
and U17692 (N_17692,N_17223,N_16864);
nand U17693 (N_17693,N_16891,N_17327);
or U17694 (N_17694,N_17231,N_17112);
nor U17695 (N_17695,N_16955,N_17378);
and U17696 (N_17696,N_17447,N_16862);
or U17697 (N_17697,N_17282,N_17488);
xnor U17698 (N_17698,N_17352,N_17208);
xor U17699 (N_17699,N_17545,N_17596);
nor U17700 (N_17700,N_16976,N_17292);
xor U17701 (N_17701,N_17268,N_17415);
or U17702 (N_17702,N_17321,N_17102);
nand U17703 (N_17703,N_17067,N_17507);
nor U17704 (N_17704,N_17141,N_17425);
and U17705 (N_17705,N_17058,N_17398);
nand U17706 (N_17706,N_16809,N_16895);
xnor U17707 (N_17707,N_17368,N_17150);
and U17708 (N_17708,N_17457,N_17464);
xor U17709 (N_17709,N_16885,N_17114);
and U17710 (N_17710,N_17169,N_17227);
or U17711 (N_17711,N_17399,N_17229);
and U17712 (N_17712,N_17234,N_17313);
nand U17713 (N_17713,N_17116,N_16931);
xor U17714 (N_17714,N_16958,N_17155);
xor U17715 (N_17715,N_17543,N_17304);
or U17716 (N_17716,N_17528,N_16859);
and U17717 (N_17717,N_17508,N_16844);
nand U17718 (N_17718,N_16927,N_17414);
and U17719 (N_17719,N_17582,N_17402);
and U17720 (N_17720,N_17445,N_16938);
and U17721 (N_17721,N_16925,N_16988);
xnor U17722 (N_17722,N_17010,N_17177);
xor U17723 (N_17723,N_16977,N_17063);
or U17724 (N_17724,N_17492,N_16980);
or U17725 (N_17725,N_17512,N_17349);
or U17726 (N_17726,N_17089,N_17419);
nand U17727 (N_17727,N_17331,N_17409);
nand U17728 (N_17728,N_17157,N_16965);
xnor U17729 (N_17729,N_17463,N_16932);
xnor U17730 (N_17730,N_16978,N_17481);
and U17731 (N_17731,N_17511,N_16883);
xor U17732 (N_17732,N_16871,N_17060);
or U17733 (N_17733,N_17143,N_16944);
nand U17734 (N_17734,N_16926,N_17174);
nor U17735 (N_17735,N_17285,N_16815);
or U17736 (N_17736,N_17270,N_17306);
xor U17737 (N_17737,N_17326,N_17318);
nor U17738 (N_17738,N_17406,N_16914);
xor U17739 (N_17739,N_17133,N_17265);
or U17740 (N_17740,N_17503,N_17217);
or U17741 (N_17741,N_17226,N_17201);
nor U17742 (N_17742,N_17407,N_17491);
nand U17743 (N_17743,N_16981,N_17211);
and U17744 (N_17744,N_17494,N_17549);
and U17745 (N_17745,N_17531,N_17045);
nand U17746 (N_17746,N_17590,N_17392);
nand U17747 (N_17747,N_17122,N_17052);
nand U17748 (N_17748,N_17110,N_17008);
or U17749 (N_17749,N_17540,N_17244);
xnor U17750 (N_17750,N_16808,N_17187);
and U17751 (N_17751,N_16820,N_16879);
nor U17752 (N_17752,N_16998,N_17500);
nor U17753 (N_17753,N_16959,N_17026);
or U17754 (N_17754,N_17149,N_17278);
and U17755 (N_17755,N_17197,N_17093);
xor U17756 (N_17756,N_17121,N_17556);
or U17757 (N_17757,N_17469,N_16996);
nor U17758 (N_17758,N_17245,N_17109);
xor U17759 (N_17759,N_17329,N_17212);
and U17760 (N_17760,N_17079,N_17597);
nand U17761 (N_17761,N_17532,N_17519);
nand U17762 (N_17762,N_17198,N_17269);
or U17763 (N_17763,N_17554,N_16935);
xnor U17764 (N_17764,N_17578,N_17389);
nor U17765 (N_17765,N_17277,N_17577);
xor U17766 (N_17766,N_17429,N_17333);
nand U17767 (N_17767,N_16923,N_17032);
xor U17768 (N_17768,N_17203,N_17287);
nand U17769 (N_17769,N_17020,N_17312);
xnor U17770 (N_17770,N_17046,N_17219);
nor U17771 (N_17771,N_17466,N_17009);
nor U17772 (N_17772,N_17296,N_17371);
nand U17773 (N_17773,N_17351,N_17040);
nor U17774 (N_17774,N_17216,N_17107);
nand U17775 (N_17775,N_17257,N_16835);
xor U17776 (N_17776,N_17309,N_16912);
nand U17777 (N_17777,N_17473,N_17123);
or U17778 (N_17778,N_17550,N_17184);
xor U17779 (N_17779,N_17584,N_17384);
nand U17780 (N_17780,N_17551,N_17165);
nand U17781 (N_17781,N_16813,N_17152);
xnor U17782 (N_17782,N_16829,N_16837);
xor U17783 (N_17783,N_17456,N_16910);
or U17784 (N_17784,N_17383,N_17207);
xnor U17785 (N_17785,N_17583,N_16937);
nand U17786 (N_17786,N_17319,N_17250);
xor U17787 (N_17787,N_16806,N_17299);
and U17788 (N_17788,N_17290,N_17088);
xnor U17789 (N_17789,N_17576,N_17486);
nor U17790 (N_17790,N_17144,N_17559);
xnor U17791 (N_17791,N_16948,N_16969);
or U17792 (N_17792,N_17106,N_17361);
nor U17793 (N_17793,N_17365,N_17388);
nand U17794 (N_17794,N_16866,N_17479);
or U17795 (N_17795,N_17396,N_17417);
xnor U17796 (N_17796,N_17595,N_17353);
nor U17797 (N_17797,N_17275,N_16812);
xnor U17798 (N_17798,N_17332,N_16984);
xnor U17799 (N_17799,N_16855,N_17220);
and U17800 (N_17800,N_16884,N_17206);
xnor U17801 (N_17801,N_16833,N_17186);
nor U17802 (N_17802,N_17233,N_17073);
nor U17803 (N_17803,N_17240,N_17087);
nand U17804 (N_17804,N_17156,N_17248);
xor U17805 (N_17805,N_16892,N_17555);
and U17806 (N_17806,N_17042,N_17453);
nor U17807 (N_17807,N_16826,N_17593);
nor U17808 (N_17808,N_16824,N_17202);
xnor U17809 (N_17809,N_16886,N_17279);
xnor U17810 (N_17810,N_17134,N_17376);
nand U17811 (N_17811,N_17498,N_17420);
nor U17812 (N_17812,N_16814,N_16911);
and U17813 (N_17813,N_16823,N_16821);
xnor U17814 (N_17814,N_16807,N_17002);
and U17815 (N_17815,N_17591,N_16887);
nand U17816 (N_17816,N_16888,N_16818);
and U17817 (N_17817,N_16805,N_16877);
nor U17818 (N_17818,N_17557,N_17439);
nand U17819 (N_17819,N_17061,N_17434);
nor U17820 (N_17820,N_17515,N_17224);
nor U17821 (N_17821,N_17362,N_16963);
and U17822 (N_17822,N_17404,N_17162);
nand U17823 (N_17823,N_17478,N_17472);
nor U17824 (N_17824,N_17422,N_17355);
nor U17825 (N_17825,N_17057,N_16881);
or U17826 (N_17826,N_17280,N_16943);
xnor U17827 (N_17827,N_17264,N_17153);
or U17828 (N_17828,N_17504,N_17117);
and U17829 (N_17829,N_17066,N_17037);
nand U17830 (N_17830,N_17370,N_17330);
nand U17831 (N_17831,N_17552,N_17308);
xor U17832 (N_17832,N_17340,N_17000);
xor U17833 (N_17833,N_17075,N_17237);
and U17834 (N_17834,N_17065,N_17298);
and U17835 (N_17835,N_16906,N_17056);
and U17836 (N_17836,N_17544,N_17029);
and U17837 (N_17837,N_17446,N_17090);
nand U17838 (N_17838,N_16902,N_16990);
xor U17839 (N_17839,N_16847,N_17435);
xor U17840 (N_17840,N_17542,N_17585);
xnor U17841 (N_17841,N_17105,N_17251);
and U17842 (N_17842,N_17172,N_17158);
xnor U17843 (N_17843,N_16842,N_17336);
xor U17844 (N_17844,N_17372,N_17154);
nand U17845 (N_17845,N_17562,N_16945);
and U17846 (N_17846,N_17344,N_17024);
nor U17847 (N_17847,N_17108,N_17256);
nand U17848 (N_17848,N_17474,N_17400);
nand U17849 (N_17849,N_17071,N_17510);
or U17850 (N_17850,N_16860,N_17350);
xnor U17851 (N_17851,N_17164,N_16921);
nand U17852 (N_17852,N_16839,N_17125);
or U17853 (N_17853,N_17522,N_17363);
nor U17854 (N_17854,N_17003,N_16942);
and U17855 (N_17855,N_16999,N_16801);
or U17856 (N_17856,N_16893,N_17423);
and U17857 (N_17857,N_17536,N_17534);
nor U17858 (N_17858,N_17483,N_17178);
nand U17859 (N_17859,N_17011,N_17347);
nor U17860 (N_17860,N_16802,N_17322);
xor U17861 (N_17861,N_17484,N_17289);
nand U17862 (N_17862,N_17261,N_17072);
nand U17863 (N_17863,N_17254,N_16836);
xor U17864 (N_17864,N_17524,N_16803);
or U17865 (N_17865,N_17373,N_17031);
nand U17866 (N_17866,N_17230,N_17568);
xnor U17867 (N_17867,N_17316,N_16916);
xor U17868 (N_17868,N_17433,N_17569);
or U17869 (N_17869,N_16909,N_16904);
nand U17870 (N_17870,N_16997,N_17243);
and U17871 (N_17871,N_17276,N_17050);
nor U17872 (N_17872,N_17044,N_17477);
nand U17873 (N_17873,N_17341,N_17183);
or U17874 (N_17874,N_17509,N_17263);
xor U17875 (N_17875,N_17236,N_17345);
xor U17876 (N_17876,N_17272,N_16934);
xor U17877 (N_17877,N_17030,N_16811);
and U17878 (N_17878,N_17180,N_17291);
nand U17879 (N_17879,N_16848,N_17092);
xnor U17880 (N_17880,N_17115,N_17470);
or U17881 (N_17881,N_16989,N_17074);
or U17882 (N_17882,N_17070,N_17541);
nor U17883 (N_17883,N_16838,N_17099);
nor U17884 (N_17884,N_17142,N_16920);
or U17885 (N_17885,N_17452,N_17475);
nand U17886 (N_17886,N_17517,N_17196);
nand U17887 (N_17887,N_17380,N_17418);
and U17888 (N_17888,N_17095,N_17599);
xor U17889 (N_17889,N_17241,N_17111);
or U17890 (N_17890,N_17561,N_16865);
nand U17891 (N_17891,N_17096,N_17255);
and U17892 (N_17892,N_17502,N_17048);
and U17893 (N_17893,N_17036,N_16951);
or U17894 (N_17894,N_17454,N_16940);
xor U17895 (N_17895,N_17148,N_17421);
and U17896 (N_17896,N_17573,N_17377);
xnor U17897 (N_17897,N_17078,N_17525);
and U17898 (N_17898,N_16991,N_17246);
nor U17899 (N_17899,N_17124,N_16922);
or U17900 (N_17900,N_16939,N_16949);
xor U17901 (N_17901,N_17190,N_17354);
xnor U17902 (N_17902,N_16832,N_16831);
nor U17903 (N_17903,N_17235,N_16930);
and U17904 (N_17904,N_17357,N_17342);
nor U17905 (N_17905,N_17273,N_17335);
or U17906 (N_17906,N_17390,N_16851);
or U17907 (N_17907,N_16962,N_17077);
nand U17908 (N_17908,N_16946,N_17033);
or U17909 (N_17909,N_16933,N_17126);
nor U17910 (N_17910,N_17189,N_16816);
nand U17911 (N_17911,N_17049,N_17191);
and U17912 (N_17912,N_17047,N_16970);
and U17913 (N_17913,N_16972,N_17173);
nand U17914 (N_17914,N_17458,N_17558);
or U17915 (N_17915,N_16961,N_16901);
nor U17916 (N_17916,N_16852,N_17450);
nand U17917 (N_17917,N_16975,N_17151);
xnor U17918 (N_17918,N_17460,N_17485);
xnor U17919 (N_17919,N_16956,N_17262);
xor U17920 (N_17920,N_16810,N_17320);
nand U17921 (N_17921,N_17100,N_17437);
nand U17922 (N_17922,N_16924,N_17175);
or U17923 (N_17923,N_17482,N_17560);
xnor U17924 (N_17924,N_17346,N_16889);
xnor U17925 (N_17925,N_17027,N_17369);
nor U17926 (N_17926,N_16869,N_17324);
nor U17927 (N_17927,N_17567,N_17068);
nor U17928 (N_17928,N_17411,N_16822);
xnor U17929 (N_17929,N_16854,N_16846);
or U17930 (N_17930,N_17468,N_17022);
or U17931 (N_17931,N_16960,N_17182);
nand U17932 (N_17932,N_17436,N_17213);
and U17933 (N_17933,N_17293,N_17428);
or U17934 (N_17934,N_17076,N_17080);
or U17935 (N_17935,N_16973,N_17019);
or U17936 (N_17936,N_17028,N_17325);
and U17937 (N_17937,N_17113,N_17317);
xor U17938 (N_17938,N_17455,N_16861);
xor U17939 (N_17939,N_16825,N_17193);
and U17940 (N_17940,N_17565,N_17288);
xnor U17941 (N_17941,N_17082,N_17537);
xor U17942 (N_17942,N_17337,N_17386);
xor U17943 (N_17943,N_17307,N_16863);
and U17944 (N_17944,N_17410,N_16950);
nor U17945 (N_17945,N_17283,N_17367);
or U17946 (N_17946,N_16907,N_16953);
or U17947 (N_17947,N_16899,N_17083);
nand U17948 (N_17948,N_16804,N_17012);
and U17949 (N_17949,N_17513,N_17286);
and U17950 (N_17950,N_16952,N_17017);
and U17951 (N_17951,N_17594,N_17586);
or U17952 (N_17952,N_17432,N_17023);
nand U17953 (N_17953,N_17538,N_17069);
or U17954 (N_17954,N_17497,N_17480);
and U17955 (N_17955,N_17571,N_17547);
xnor U17956 (N_17956,N_17426,N_17305);
and U17957 (N_17957,N_16994,N_17575);
nor U17958 (N_17958,N_17252,N_17430);
and U17959 (N_17959,N_17493,N_17592);
xnor U17960 (N_17960,N_17145,N_16966);
and U17961 (N_17961,N_16954,N_17382);
and U17962 (N_17962,N_16880,N_16967);
nand U17963 (N_17963,N_17016,N_17310);
nand U17964 (N_17964,N_17465,N_17444);
nand U17965 (N_17965,N_17232,N_17385);
nand U17966 (N_17966,N_17338,N_16800);
and U17967 (N_17967,N_17055,N_17408);
xor U17968 (N_17968,N_16968,N_17448);
xor U17969 (N_17969,N_17566,N_17137);
xor U17970 (N_17970,N_17495,N_17598);
nand U17971 (N_17971,N_17514,N_17239);
or U17972 (N_17972,N_17222,N_16890);
and U17973 (N_17973,N_17520,N_17170);
nand U17974 (N_17974,N_16894,N_16830);
xnor U17975 (N_17975,N_17471,N_17413);
xnor U17976 (N_17976,N_17238,N_16873);
or U17977 (N_17977,N_17516,N_16947);
and U17978 (N_17978,N_16874,N_17302);
or U17979 (N_17979,N_17295,N_17461);
nor U17980 (N_17980,N_16993,N_17258);
and U17981 (N_17981,N_17104,N_17266);
nor U17982 (N_17982,N_16882,N_17334);
or U17983 (N_17983,N_17366,N_17581);
or U17984 (N_17984,N_17128,N_17539);
and U17985 (N_17985,N_17381,N_17467);
or U17986 (N_17986,N_17018,N_17328);
or U17987 (N_17987,N_17005,N_17192);
xnor U17988 (N_17988,N_17171,N_17001);
and U17989 (N_17989,N_17523,N_17253);
xor U17990 (N_17990,N_17006,N_16878);
or U17991 (N_17991,N_17587,N_17424);
xor U17992 (N_17992,N_16983,N_17084);
nor U17993 (N_17993,N_17091,N_17356);
nor U17994 (N_17994,N_17294,N_17501);
or U17995 (N_17995,N_17303,N_17499);
and U17996 (N_17996,N_17098,N_17564);
and U17997 (N_17997,N_16929,N_16856);
and U17998 (N_17998,N_16896,N_17553);
xnor U17999 (N_17999,N_17442,N_17339);
nor U18000 (N_18000,N_16927,N_17067);
and U18001 (N_18001,N_17459,N_17511);
nand U18002 (N_18002,N_17041,N_16974);
or U18003 (N_18003,N_17491,N_17218);
nand U18004 (N_18004,N_16889,N_17220);
nor U18005 (N_18005,N_16913,N_17409);
or U18006 (N_18006,N_17402,N_16928);
nor U18007 (N_18007,N_16898,N_16864);
nor U18008 (N_18008,N_16976,N_17359);
nand U18009 (N_18009,N_16965,N_17152);
nor U18010 (N_18010,N_17566,N_17354);
nand U18011 (N_18011,N_17363,N_17146);
and U18012 (N_18012,N_17574,N_17534);
xor U18013 (N_18013,N_17565,N_16949);
nor U18014 (N_18014,N_16919,N_16854);
nor U18015 (N_18015,N_16813,N_17058);
and U18016 (N_18016,N_17090,N_17301);
nand U18017 (N_18017,N_17399,N_17214);
and U18018 (N_18018,N_16887,N_17434);
and U18019 (N_18019,N_16802,N_16872);
nor U18020 (N_18020,N_17202,N_17151);
nor U18021 (N_18021,N_16992,N_17041);
nand U18022 (N_18022,N_17291,N_17293);
and U18023 (N_18023,N_16813,N_17259);
xnor U18024 (N_18024,N_17103,N_17116);
and U18025 (N_18025,N_17033,N_17183);
nor U18026 (N_18026,N_16808,N_17554);
nand U18027 (N_18027,N_17534,N_17374);
or U18028 (N_18028,N_16808,N_17435);
or U18029 (N_18029,N_17402,N_16836);
or U18030 (N_18030,N_17005,N_17177);
or U18031 (N_18031,N_17459,N_17160);
nor U18032 (N_18032,N_17586,N_17508);
or U18033 (N_18033,N_17268,N_16986);
and U18034 (N_18034,N_17201,N_17325);
nor U18035 (N_18035,N_17315,N_17553);
nor U18036 (N_18036,N_16891,N_16884);
or U18037 (N_18037,N_16900,N_17350);
or U18038 (N_18038,N_17440,N_17363);
or U18039 (N_18039,N_17507,N_17465);
xor U18040 (N_18040,N_16964,N_17400);
nand U18041 (N_18041,N_16854,N_16916);
nor U18042 (N_18042,N_17537,N_17376);
and U18043 (N_18043,N_17285,N_16824);
and U18044 (N_18044,N_16816,N_17542);
xor U18045 (N_18045,N_17455,N_17384);
or U18046 (N_18046,N_17587,N_17332);
or U18047 (N_18047,N_17018,N_17407);
nand U18048 (N_18048,N_17560,N_17105);
or U18049 (N_18049,N_17401,N_16961);
and U18050 (N_18050,N_16896,N_17317);
nor U18051 (N_18051,N_17548,N_17043);
and U18052 (N_18052,N_17176,N_16823);
nor U18053 (N_18053,N_17481,N_17469);
nor U18054 (N_18054,N_17438,N_17192);
or U18055 (N_18055,N_17408,N_17003);
xnor U18056 (N_18056,N_16915,N_17500);
and U18057 (N_18057,N_17218,N_17502);
or U18058 (N_18058,N_17466,N_17546);
and U18059 (N_18059,N_17087,N_17284);
xor U18060 (N_18060,N_16921,N_17441);
and U18061 (N_18061,N_17114,N_17115);
nor U18062 (N_18062,N_16863,N_16939);
or U18063 (N_18063,N_17031,N_17035);
xor U18064 (N_18064,N_17179,N_17159);
or U18065 (N_18065,N_17001,N_16812);
and U18066 (N_18066,N_17431,N_16888);
and U18067 (N_18067,N_17171,N_17166);
xor U18068 (N_18068,N_16809,N_16998);
or U18069 (N_18069,N_17537,N_16928);
nand U18070 (N_18070,N_17225,N_16822);
and U18071 (N_18071,N_17157,N_17178);
nand U18072 (N_18072,N_17410,N_17379);
nor U18073 (N_18073,N_16887,N_17503);
and U18074 (N_18074,N_17383,N_17558);
nor U18075 (N_18075,N_16978,N_17285);
nor U18076 (N_18076,N_17169,N_16883);
xnor U18077 (N_18077,N_17112,N_17435);
xor U18078 (N_18078,N_17030,N_16825);
xor U18079 (N_18079,N_17377,N_17499);
or U18080 (N_18080,N_17206,N_16990);
nand U18081 (N_18081,N_16970,N_17501);
nor U18082 (N_18082,N_16862,N_17150);
and U18083 (N_18083,N_16824,N_16876);
and U18084 (N_18084,N_16868,N_17580);
xnor U18085 (N_18085,N_17363,N_16887);
xnor U18086 (N_18086,N_16985,N_16822);
xnor U18087 (N_18087,N_17200,N_17248);
and U18088 (N_18088,N_17578,N_17019);
or U18089 (N_18089,N_17094,N_16876);
xor U18090 (N_18090,N_17134,N_17240);
and U18091 (N_18091,N_17014,N_17253);
and U18092 (N_18092,N_17076,N_17010);
xor U18093 (N_18093,N_17380,N_17007);
xor U18094 (N_18094,N_17282,N_17110);
nor U18095 (N_18095,N_17199,N_16851);
and U18096 (N_18096,N_17504,N_16953);
and U18097 (N_18097,N_16832,N_17154);
nand U18098 (N_18098,N_17317,N_17535);
xor U18099 (N_18099,N_17010,N_17272);
nand U18100 (N_18100,N_17061,N_16967);
nor U18101 (N_18101,N_17148,N_17446);
or U18102 (N_18102,N_16872,N_17554);
or U18103 (N_18103,N_17432,N_17325);
xnor U18104 (N_18104,N_16852,N_17133);
and U18105 (N_18105,N_17342,N_16983);
nor U18106 (N_18106,N_17276,N_17379);
nor U18107 (N_18107,N_16902,N_17438);
or U18108 (N_18108,N_17282,N_17257);
xnor U18109 (N_18109,N_16815,N_17365);
xor U18110 (N_18110,N_17418,N_17422);
nor U18111 (N_18111,N_17249,N_17339);
or U18112 (N_18112,N_17194,N_17180);
or U18113 (N_18113,N_17223,N_17147);
or U18114 (N_18114,N_17006,N_17487);
nor U18115 (N_18115,N_17322,N_17062);
and U18116 (N_18116,N_17193,N_17217);
nand U18117 (N_18117,N_17049,N_17111);
or U18118 (N_18118,N_17024,N_17426);
and U18119 (N_18119,N_16938,N_17476);
or U18120 (N_18120,N_17497,N_17077);
and U18121 (N_18121,N_17571,N_17470);
nor U18122 (N_18122,N_17368,N_16820);
and U18123 (N_18123,N_17033,N_17053);
xnor U18124 (N_18124,N_16911,N_17290);
or U18125 (N_18125,N_17476,N_16994);
and U18126 (N_18126,N_17140,N_17312);
nor U18127 (N_18127,N_17272,N_17556);
nand U18128 (N_18128,N_17324,N_17088);
or U18129 (N_18129,N_17382,N_17158);
nor U18130 (N_18130,N_17408,N_17398);
and U18131 (N_18131,N_17188,N_17345);
nor U18132 (N_18132,N_17083,N_17018);
or U18133 (N_18133,N_17425,N_16830);
or U18134 (N_18134,N_17553,N_16928);
nor U18135 (N_18135,N_16887,N_17123);
xor U18136 (N_18136,N_17567,N_17011);
or U18137 (N_18137,N_16815,N_17141);
nand U18138 (N_18138,N_17068,N_17492);
nor U18139 (N_18139,N_17479,N_17137);
nor U18140 (N_18140,N_17137,N_17238);
nor U18141 (N_18141,N_17225,N_16971);
nor U18142 (N_18142,N_16827,N_17586);
xnor U18143 (N_18143,N_16933,N_16890);
xor U18144 (N_18144,N_17277,N_16927);
nand U18145 (N_18145,N_16963,N_16833);
or U18146 (N_18146,N_17003,N_17095);
or U18147 (N_18147,N_17284,N_17521);
or U18148 (N_18148,N_17476,N_16806);
nor U18149 (N_18149,N_16819,N_17206);
nor U18150 (N_18150,N_17480,N_17416);
and U18151 (N_18151,N_17531,N_17501);
nor U18152 (N_18152,N_17205,N_16870);
and U18153 (N_18153,N_16907,N_17177);
nor U18154 (N_18154,N_16873,N_17500);
or U18155 (N_18155,N_17088,N_16802);
nand U18156 (N_18156,N_17151,N_17156);
nor U18157 (N_18157,N_17413,N_17554);
nand U18158 (N_18158,N_17557,N_16854);
nor U18159 (N_18159,N_17050,N_17016);
or U18160 (N_18160,N_17420,N_17574);
and U18161 (N_18161,N_17285,N_17507);
nand U18162 (N_18162,N_17494,N_17129);
nor U18163 (N_18163,N_17233,N_17410);
nand U18164 (N_18164,N_17101,N_16825);
xor U18165 (N_18165,N_16814,N_16891);
nor U18166 (N_18166,N_17567,N_16873);
or U18167 (N_18167,N_17403,N_17516);
xor U18168 (N_18168,N_16991,N_17085);
xnor U18169 (N_18169,N_16919,N_17083);
xor U18170 (N_18170,N_17280,N_17286);
or U18171 (N_18171,N_17281,N_16905);
or U18172 (N_18172,N_17523,N_17474);
xor U18173 (N_18173,N_17425,N_17348);
xor U18174 (N_18174,N_17212,N_17375);
xnor U18175 (N_18175,N_17592,N_16876);
nand U18176 (N_18176,N_17390,N_17545);
or U18177 (N_18177,N_17178,N_17523);
or U18178 (N_18178,N_17502,N_17109);
xor U18179 (N_18179,N_17527,N_17426);
nor U18180 (N_18180,N_17527,N_16991);
or U18181 (N_18181,N_17318,N_16997);
xnor U18182 (N_18182,N_16830,N_17350);
and U18183 (N_18183,N_17110,N_17362);
nor U18184 (N_18184,N_16834,N_16968);
xnor U18185 (N_18185,N_16943,N_17216);
nand U18186 (N_18186,N_17148,N_17174);
nand U18187 (N_18187,N_17047,N_17347);
xor U18188 (N_18188,N_17236,N_16898);
nand U18189 (N_18189,N_16870,N_17221);
xor U18190 (N_18190,N_17064,N_17012);
xnor U18191 (N_18191,N_17512,N_17283);
nand U18192 (N_18192,N_17567,N_17379);
and U18193 (N_18193,N_17123,N_17597);
or U18194 (N_18194,N_17086,N_17434);
nor U18195 (N_18195,N_17133,N_17547);
nor U18196 (N_18196,N_17031,N_17063);
or U18197 (N_18197,N_16880,N_17487);
and U18198 (N_18198,N_16947,N_17067);
nand U18199 (N_18199,N_17298,N_17127);
nor U18200 (N_18200,N_16841,N_17483);
xor U18201 (N_18201,N_16877,N_17023);
nor U18202 (N_18202,N_17086,N_17391);
or U18203 (N_18203,N_17072,N_17111);
or U18204 (N_18204,N_17210,N_17300);
nor U18205 (N_18205,N_17270,N_17490);
xor U18206 (N_18206,N_16860,N_16832);
nor U18207 (N_18207,N_16879,N_16868);
xor U18208 (N_18208,N_17318,N_17040);
nand U18209 (N_18209,N_17311,N_17368);
and U18210 (N_18210,N_17194,N_16899);
and U18211 (N_18211,N_17347,N_17512);
nand U18212 (N_18212,N_17059,N_17262);
nand U18213 (N_18213,N_16991,N_16864);
nand U18214 (N_18214,N_16840,N_16945);
and U18215 (N_18215,N_17362,N_17022);
or U18216 (N_18216,N_17051,N_16947);
nand U18217 (N_18217,N_17018,N_17073);
nor U18218 (N_18218,N_17201,N_16901);
or U18219 (N_18219,N_17294,N_17371);
and U18220 (N_18220,N_17055,N_17373);
or U18221 (N_18221,N_16820,N_16897);
or U18222 (N_18222,N_17116,N_17347);
nand U18223 (N_18223,N_16815,N_17429);
nand U18224 (N_18224,N_16989,N_17102);
and U18225 (N_18225,N_17061,N_16804);
xor U18226 (N_18226,N_17184,N_17025);
nor U18227 (N_18227,N_17300,N_17322);
xnor U18228 (N_18228,N_17329,N_16987);
nor U18229 (N_18229,N_17001,N_17530);
xor U18230 (N_18230,N_16950,N_17530);
xor U18231 (N_18231,N_17502,N_17471);
nor U18232 (N_18232,N_17436,N_17187);
xor U18233 (N_18233,N_17516,N_17511);
xor U18234 (N_18234,N_17502,N_16821);
nand U18235 (N_18235,N_17190,N_17441);
or U18236 (N_18236,N_17408,N_17139);
or U18237 (N_18237,N_17438,N_16979);
nand U18238 (N_18238,N_17126,N_16807);
or U18239 (N_18239,N_17577,N_17505);
or U18240 (N_18240,N_16855,N_17222);
or U18241 (N_18241,N_17260,N_17321);
xor U18242 (N_18242,N_17542,N_17236);
xor U18243 (N_18243,N_17491,N_16894);
or U18244 (N_18244,N_17583,N_17444);
nor U18245 (N_18245,N_16930,N_17211);
and U18246 (N_18246,N_16906,N_16838);
nand U18247 (N_18247,N_17255,N_16981);
xnor U18248 (N_18248,N_16911,N_16939);
or U18249 (N_18249,N_16815,N_17363);
nor U18250 (N_18250,N_16989,N_17123);
nor U18251 (N_18251,N_17314,N_17225);
xor U18252 (N_18252,N_17004,N_17022);
and U18253 (N_18253,N_16838,N_16823);
xnor U18254 (N_18254,N_16991,N_17516);
nor U18255 (N_18255,N_16884,N_17143);
or U18256 (N_18256,N_17507,N_16851);
xnor U18257 (N_18257,N_17514,N_17432);
or U18258 (N_18258,N_17281,N_17148);
xnor U18259 (N_18259,N_17354,N_17552);
nor U18260 (N_18260,N_17258,N_17205);
nand U18261 (N_18261,N_17201,N_17131);
or U18262 (N_18262,N_17322,N_17041);
nor U18263 (N_18263,N_17395,N_17483);
and U18264 (N_18264,N_17443,N_16859);
nor U18265 (N_18265,N_17216,N_16952);
and U18266 (N_18266,N_17222,N_17477);
and U18267 (N_18267,N_17137,N_16862);
nand U18268 (N_18268,N_16876,N_17599);
nand U18269 (N_18269,N_17007,N_17342);
or U18270 (N_18270,N_17174,N_17034);
xor U18271 (N_18271,N_17494,N_16935);
nand U18272 (N_18272,N_17123,N_17362);
nor U18273 (N_18273,N_17375,N_17023);
nand U18274 (N_18274,N_17457,N_17468);
xor U18275 (N_18275,N_17224,N_17413);
nand U18276 (N_18276,N_16918,N_17464);
nor U18277 (N_18277,N_16920,N_17491);
or U18278 (N_18278,N_17100,N_17248);
nand U18279 (N_18279,N_17158,N_17501);
and U18280 (N_18280,N_16879,N_17231);
and U18281 (N_18281,N_16821,N_16925);
xor U18282 (N_18282,N_17572,N_17534);
and U18283 (N_18283,N_17089,N_16953);
or U18284 (N_18284,N_17521,N_16840);
and U18285 (N_18285,N_17265,N_17077);
nor U18286 (N_18286,N_17232,N_17557);
or U18287 (N_18287,N_16952,N_16950);
nand U18288 (N_18288,N_17041,N_17162);
and U18289 (N_18289,N_17508,N_17243);
or U18290 (N_18290,N_17529,N_17226);
nor U18291 (N_18291,N_16866,N_17451);
nor U18292 (N_18292,N_16873,N_17032);
nand U18293 (N_18293,N_17306,N_17141);
and U18294 (N_18294,N_17084,N_17143);
nor U18295 (N_18295,N_17382,N_17413);
nor U18296 (N_18296,N_17010,N_17275);
and U18297 (N_18297,N_17130,N_16822);
or U18298 (N_18298,N_17546,N_16804);
and U18299 (N_18299,N_16990,N_17389);
nor U18300 (N_18300,N_17183,N_17411);
or U18301 (N_18301,N_16885,N_17226);
or U18302 (N_18302,N_17116,N_17214);
nor U18303 (N_18303,N_16861,N_17085);
or U18304 (N_18304,N_17596,N_17176);
nand U18305 (N_18305,N_17146,N_17543);
and U18306 (N_18306,N_16874,N_17311);
or U18307 (N_18307,N_16920,N_17592);
nor U18308 (N_18308,N_16888,N_17592);
nand U18309 (N_18309,N_17054,N_16976);
xor U18310 (N_18310,N_17469,N_17279);
nand U18311 (N_18311,N_17556,N_17140);
xor U18312 (N_18312,N_17455,N_17340);
xor U18313 (N_18313,N_17547,N_17535);
or U18314 (N_18314,N_17029,N_16858);
or U18315 (N_18315,N_17225,N_17598);
xnor U18316 (N_18316,N_16843,N_17007);
xnor U18317 (N_18317,N_16920,N_16838);
or U18318 (N_18318,N_16921,N_17197);
nor U18319 (N_18319,N_16885,N_17289);
xnor U18320 (N_18320,N_16804,N_17337);
xnor U18321 (N_18321,N_17177,N_16946);
nand U18322 (N_18322,N_16866,N_16959);
and U18323 (N_18323,N_16881,N_17071);
nand U18324 (N_18324,N_17370,N_17328);
or U18325 (N_18325,N_17443,N_17571);
and U18326 (N_18326,N_17335,N_16808);
nor U18327 (N_18327,N_16815,N_16820);
nor U18328 (N_18328,N_17164,N_17590);
or U18329 (N_18329,N_17291,N_17285);
xnor U18330 (N_18330,N_17393,N_16975);
or U18331 (N_18331,N_16948,N_17259);
xor U18332 (N_18332,N_17137,N_17144);
nand U18333 (N_18333,N_17515,N_16840);
and U18334 (N_18334,N_17082,N_17251);
xnor U18335 (N_18335,N_17244,N_17113);
nor U18336 (N_18336,N_17060,N_16883);
or U18337 (N_18337,N_17283,N_17195);
or U18338 (N_18338,N_16986,N_16922);
xnor U18339 (N_18339,N_17040,N_17070);
nor U18340 (N_18340,N_17267,N_16878);
nand U18341 (N_18341,N_16953,N_17394);
or U18342 (N_18342,N_17120,N_16894);
or U18343 (N_18343,N_17446,N_17180);
xor U18344 (N_18344,N_16824,N_17312);
nand U18345 (N_18345,N_17489,N_17591);
or U18346 (N_18346,N_17522,N_17454);
nor U18347 (N_18347,N_17187,N_17475);
nand U18348 (N_18348,N_17198,N_17417);
nand U18349 (N_18349,N_16914,N_17426);
or U18350 (N_18350,N_17526,N_17059);
nand U18351 (N_18351,N_17515,N_17344);
or U18352 (N_18352,N_16921,N_17373);
xnor U18353 (N_18353,N_17243,N_16986);
nor U18354 (N_18354,N_17327,N_17322);
and U18355 (N_18355,N_17139,N_17238);
nor U18356 (N_18356,N_16980,N_17407);
xor U18357 (N_18357,N_17234,N_16977);
or U18358 (N_18358,N_17446,N_17033);
nand U18359 (N_18359,N_17304,N_16957);
and U18360 (N_18360,N_17004,N_17379);
and U18361 (N_18361,N_17349,N_17421);
nand U18362 (N_18362,N_17156,N_17128);
xor U18363 (N_18363,N_17529,N_17203);
nor U18364 (N_18364,N_17325,N_17130);
or U18365 (N_18365,N_16996,N_17020);
nand U18366 (N_18366,N_16915,N_16919);
or U18367 (N_18367,N_17242,N_17384);
nand U18368 (N_18368,N_17333,N_17035);
nand U18369 (N_18369,N_17471,N_17409);
xor U18370 (N_18370,N_17128,N_17129);
or U18371 (N_18371,N_17304,N_17368);
and U18372 (N_18372,N_17153,N_17562);
nand U18373 (N_18373,N_16903,N_17120);
nor U18374 (N_18374,N_17337,N_17164);
and U18375 (N_18375,N_17230,N_17417);
nor U18376 (N_18376,N_17109,N_16929);
and U18377 (N_18377,N_17101,N_17190);
nand U18378 (N_18378,N_17081,N_17011);
and U18379 (N_18379,N_17263,N_17312);
or U18380 (N_18380,N_16871,N_17362);
nand U18381 (N_18381,N_17142,N_17505);
or U18382 (N_18382,N_17539,N_16911);
xnor U18383 (N_18383,N_16940,N_17212);
and U18384 (N_18384,N_17174,N_17099);
and U18385 (N_18385,N_17100,N_17475);
nand U18386 (N_18386,N_16800,N_17083);
nand U18387 (N_18387,N_16815,N_16839);
and U18388 (N_18388,N_17168,N_17285);
nand U18389 (N_18389,N_16813,N_17480);
nand U18390 (N_18390,N_16961,N_17462);
nand U18391 (N_18391,N_17595,N_17492);
nand U18392 (N_18392,N_17511,N_17382);
nor U18393 (N_18393,N_16891,N_17374);
and U18394 (N_18394,N_16997,N_17095);
or U18395 (N_18395,N_17536,N_16934);
or U18396 (N_18396,N_16843,N_16913);
nor U18397 (N_18397,N_16906,N_16972);
nand U18398 (N_18398,N_17216,N_17099);
nand U18399 (N_18399,N_17281,N_17444);
xnor U18400 (N_18400,N_17622,N_18103);
nand U18401 (N_18401,N_17811,N_18200);
xor U18402 (N_18402,N_18273,N_17675);
xnor U18403 (N_18403,N_18272,N_18388);
and U18404 (N_18404,N_17655,N_17804);
or U18405 (N_18405,N_17891,N_17719);
and U18406 (N_18406,N_18338,N_17813);
nor U18407 (N_18407,N_18279,N_17861);
and U18408 (N_18408,N_18005,N_17775);
and U18409 (N_18409,N_18006,N_18092);
nor U18410 (N_18410,N_17643,N_18227);
nor U18411 (N_18411,N_17820,N_18126);
or U18412 (N_18412,N_18398,N_18260);
nand U18413 (N_18413,N_17706,N_18361);
and U18414 (N_18414,N_18231,N_18037);
and U18415 (N_18415,N_18331,N_18186);
or U18416 (N_18416,N_17832,N_18038);
and U18417 (N_18417,N_18147,N_17904);
and U18418 (N_18418,N_17845,N_17866);
nand U18419 (N_18419,N_18163,N_18206);
or U18420 (N_18420,N_17920,N_18019);
or U18421 (N_18421,N_17701,N_17708);
or U18422 (N_18422,N_18230,N_18057);
and U18423 (N_18423,N_17789,N_18300);
nand U18424 (N_18424,N_18214,N_17790);
nand U18425 (N_18425,N_18141,N_17843);
nand U18426 (N_18426,N_18150,N_18267);
and U18427 (N_18427,N_18078,N_18143);
xnor U18428 (N_18428,N_18266,N_18316);
xnor U18429 (N_18429,N_18118,N_18034);
nor U18430 (N_18430,N_18033,N_18086);
nor U18431 (N_18431,N_17688,N_18226);
nor U18432 (N_18432,N_17852,N_18304);
and U18433 (N_18433,N_18275,N_17890);
or U18434 (N_18434,N_18327,N_17628);
nand U18435 (N_18435,N_18156,N_18363);
nor U18436 (N_18436,N_18383,N_18208);
and U18437 (N_18437,N_18323,N_18154);
nand U18438 (N_18438,N_18310,N_17968);
xor U18439 (N_18439,N_17608,N_17858);
and U18440 (N_18440,N_17896,N_17970);
xor U18441 (N_18441,N_17826,N_17644);
and U18442 (N_18442,N_17750,N_17963);
nor U18443 (N_18443,N_17773,N_17652);
and U18444 (N_18444,N_17912,N_18129);
or U18445 (N_18445,N_17934,N_17621);
nand U18446 (N_18446,N_17677,N_17959);
or U18447 (N_18447,N_17840,N_17925);
or U18448 (N_18448,N_17630,N_17803);
or U18449 (N_18449,N_17690,N_17808);
or U18450 (N_18450,N_17636,N_17783);
or U18451 (N_18451,N_17863,N_17637);
and U18452 (N_18452,N_18198,N_18274);
nor U18453 (N_18453,N_18047,N_18018);
and U18454 (N_18454,N_18091,N_17795);
nor U18455 (N_18455,N_17744,N_18318);
nor U18456 (N_18456,N_17850,N_17984);
and U18457 (N_18457,N_17967,N_18305);
nand U18458 (N_18458,N_18209,N_17642);
and U18459 (N_18459,N_18023,N_18097);
nand U18460 (N_18460,N_17767,N_17945);
or U18461 (N_18461,N_17830,N_18211);
xnor U18462 (N_18462,N_17936,N_17838);
nor U18463 (N_18463,N_18251,N_17791);
xnor U18464 (N_18464,N_17741,N_18121);
or U18465 (N_18465,N_18142,N_17699);
xor U18466 (N_18466,N_17757,N_17609);
nand U18467 (N_18467,N_18170,N_17978);
nand U18468 (N_18468,N_18290,N_17825);
and U18469 (N_18469,N_17647,N_18098);
nor U18470 (N_18470,N_18139,N_18375);
xnor U18471 (N_18471,N_17869,N_18149);
nand U18472 (N_18472,N_18377,N_17835);
nand U18473 (N_18473,N_17908,N_18196);
xor U18474 (N_18474,N_17943,N_18113);
and U18475 (N_18475,N_18213,N_17619);
xnor U18476 (N_18476,N_17821,N_18342);
nor U18477 (N_18477,N_17785,N_17625);
and U18478 (N_18478,N_18204,N_18177);
nor U18479 (N_18479,N_17672,N_17842);
or U18480 (N_18480,N_17906,N_18244);
nand U18481 (N_18481,N_18080,N_17695);
xnor U18482 (N_18482,N_17694,N_18120);
or U18483 (N_18483,N_18359,N_18364);
nand U18484 (N_18484,N_18241,N_17932);
and U18485 (N_18485,N_18069,N_18136);
or U18486 (N_18486,N_17926,N_17919);
and U18487 (N_18487,N_18058,N_17903);
or U18488 (N_18488,N_18062,N_17664);
xor U18489 (N_18489,N_17898,N_17818);
xor U18490 (N_18490,N_18010,N_18345);
nor U18491 (N_18491,N_18084,N_17880);
or U18492 (N_18492,N_17895,N_17996);
or U18493 (N_18493,N_17864,N_18216);
or U18494 (N_18494,N_17654,N_18271);
and U18495 (N_18495,N_18334,N_18035);
and U18496 (N_18496,N_18075,N_18157);
nor U18497 (N_18497,N_18050,N_17833);
nand U18498 (N_18498,N_17693,N_17679);
xor U18499 (N_18499,N_18276,N_18042);
nand U18500 (N_18500,N_18232,N_18228);
and U18501 (N_18501,N_18022,N_17823);
or U18502 (N_18502,N_17889,N_17915);
and U18503 (N_18503,N_17776,N_17940);
nor U18504 (N_18504,N_17979,N_17728);
nor U18505 (N_18505,N_18144,N_18253);
nand U18506 (N_18506,N_18393,N_17718);
nand U18507 (N_18507,N_17616,N_18222);
xor U18508 (N_18508,N_18045,N_17933);
nor U18509 (N_18509,N_17986,N_17614);
and U18510 (N_18510,N_18234,N_18224);
xor U18511 (N_18511,N_18320,N_17962);
nand U18512 (N_18512,N_17966,N_17607);
or U18513 (N_18513,N_18162,N_17914);
nand U18514 (N_18514,N_17907,N_18295);
nand U18515 (N_18515,N_18053,N_18242);
or U18516 (N_18516,N_17662,N_17960);
xnor U18517 (N_18517,N_18344,N_18087);
xor U18518 (N_18518,N_18376,N_18263);
or U18519 (N_18519,N_18090,N_18014);
xnor U18520 (N_18520,N_17853,N_18281);
or U18521 (N_18521,N_17604,N_17646);
and U18522 (N_18522,N_18193,N_18130);
xor U18523 (N_18523,N_18061,N_17954);
and U18524 (N_18524,N_18296,N_18108);
nor U18525 (N_18525,N_18060,N_18082);
nor U18526 (N_18526,N_18270,N_17924);
or U18527 (N_18527,N_17849,N_18337);
and U18528 (N_18528,N_18184,N_17602);
xor U18529 (N_18529,N_17922,N_17894);
or U18530 (N_18530,N_18329,N_17689);
nor U18531 (N_18531,N_17711,N_18360);
nand U18532 (N_18532,N_18212,N_17848);
or U18533 (N_18533,N_17999,N_18347);
or U18534 (N_18534,N_18390,N_18127);
xnor U18535 (N_18535,N_17913,N_17686);
or U18536 (N_18536,N_18221,N_18358);
and U18537 (N_18537,N_17753,N_17713);
nor U18538 (N_18538,N_18250,N_17725);
or U18539 (N_18539,N_18194,N_18031);
and U18540 (N_18540,N_17806,N_18104);
or U18541 (N_18541,N_17897,N_17610);
nand U18542 (N_18542,N_17641,N_17947);
xor U18543 (N_18543,N_17730,N_18125);
xnor U18544 (N_18544,N_17839,N_17824);
nor U18545 (N_18545,N_17887,N_18063);
xor U18546 (N_18546,N_17834,N_18399);
xnor U18547 (N_18547,N_17851,N_17819);
nor U18548 (N_18548,N_17831,N_17696);
nor U18549 (N_18549,N_18306,N_17605);
nor U18550 (N_18550,N_18009,N_18265);
or U18551 (N_18551,N_17615,N_18387);
or U18552 (N_18552,N_18085,N_17946);
nor U18553 (N_18553,N_17691,N_17617);
or U18554 (N_18554,N_17632,N_18164);
and U18555 (N_18555,N_17687,N_18352);
xor U18556 (N_18556,N_18044,N_18261);
and U18557 (N_18557,N_17739,N_17964);
and U18558 (N_18558,N_18133,N_17857);
and U18559 (N_18559,N_17668,N_18026);
nand U18560 (N_18560,N_18099,N_17660);
and U18561 (N_18561,N_18225,N_18235);
and U18562 (N_18562,N_18178,N_17988);
nor U18563 (N_18563,N_18003,N_18040);
xor U18564 (N_18564,N_18151,N_18373);
xor U18565 (N_18565,N_17611,N_17633);
xnor U18566 (N_18566,N_18207,N_18166);
and U18567 (N_18567,N_18081,N_17653);
nand U18568 (N_18568,N_17724,N_17770);
nor U18569 (N_18569,N_18029,N_17648);
xnor U18570 (N_18570,N_17714,N_17969);
or U18571 (N_18571,N_17624,N_18039);
and U18572 (N_18572,N_17768,N_17758);
nand U18573 (N_18573,N_18285,N_18094);
and U18574 (N_18574,N_18109,N_18255);
xor U18575 (N_18575,N_18122,N_18074);
nor U18576 (N_18576,N_17909,N_18105);
nand U18577 (N_18577,N_18002,N_17705);
or U18578 (N_18578,N_18089,N_18328);
nor U18579 (N_18579,N_18169,N_18137);
or U18580 (N_18580,N_18343,N_17879);
or U18581 (N_18581,N_17805,N_18189);
nand U18582 (N_18582,N_18257,N_18210);
and U18583 (N_18583,N_17751,N_18321);
nand U18584 (N_18584,N_18293,N_17651);
xor U18585 (N_18585,N_17981,N_17900);
nand U18586 (N_18586,N_17910,N_18000);
xnor U18587 (N_18587,N_18248,N_18135);
xor U18588 (N_18588,N_17674,N_17921);
xnor U18589 (N_18589,N_18048,N_17888);
and U18590 (N_18590,N_18394,N_17854);
nor U18591 (N_18591,N_18220,N_18299);
nor U18592 (N_18592,N_18041,N_18036);
nand U18593 (N_18593,N_17881,N_17883);
nor U18594 (N_18594,N_17747,N_17721);
nor U18595 (N_18595,N_18068,N_17980);
and U18596 (N_18596,N_17623,N_17923);
and U18597 (N_18597,N_18123,N_18382);
nand U18598 (N_18598,N_17973,N_18254);
or U18599 (N_18599,N_18256,N_17697);
and U18600 (N_18600,N_17829,N_18268);
and U18601 (N_18601,N_17704,N_18397);
nand U18602 (N_18602,N_17797,N_17671);
and U18603 (N_18603,N_18183,N_18155);
nand U18604 (N_18604,N_18140,N_17722);
xor U18605 (N_18605,N_17712,N_18366);
nand U18606 (N_18606,N_17807,N_18187);
nor U18607 (N_18607,N_17860,N_17743);
xor U18608 (N_18608,N_17752,N_17737);
and U18609 (N_18609,N_18322,N_17634);
nand U18610 (N_18610,N_17663,N_18012);
nor U18611 (N_18611,N_18369,N_18365);
nand U18612 (N_18612,N_17837,N_18379);
xnor U18613 (N_18613,N_17656,N_18395);
nand U18614 (N_18614,N_18088,N_18341);
or U18615 (N_18615,N_17682,N_18385);
nor U18616 (N_18616,N_18071,N_18203);
nor U18617 (N_18617,N_17603,N_17916);
and U18618 (N_18618,N_18046,N_18020);
nand U18619 (N_18619,N_17709,N_18017);
xor U18620 (N_18620,N_17990,N_17794);
or U18621 (N_18621,N_17918,N_18115);
nor U18622 (N_18622,N_17681,N_18171);
nand U18623 (N_18623,N_18013,N_18028);
nand U18624 (N_18624,N_17998,N_17972);
nor U18625 (N_18625,N_17836,N_18236);
and U18626 (N_18626,N_17991,N_17745);
xor U18627 (N_18627,N_18051,N_18378);
nand U18628 (N_18628,N_18215,N_17673);
nor U18629 (N_18629,N_18350,N_18243);
xor U18630 (N_18630,N_18015,N_17600);
xor U18631 (N_18631,N_18032,N_18278);
or U18632 (N_18632,N_17720,N_17670);
nand U18633 (N_18633,N_18030,N_18070);
and U18634 (N_18634,N_18252,N_17828);
xnor U18635 (N_18635,N_17792,N_18055);
nor U18636 (N_18636,N_17928,N_18396);
nand U18637 (N_18637,N_17886,N_18064);
and U18638 (N_18638,N_18016,N_17601);
or U18639 (N_18639,N_17731,N_18258);
and U18640 (N_18640,N_18066,N_17765);
nand U18641 (N_18641,N_17976,N_18330);
or U18642 (N_18642,N_17736,N_17983);
nor U18643 (N_18643,N_18286,N_17878);
nand U18644 (N_18644,N_18324,N_17938);
nor U18645 (N_18645,N_18181,N_17958);
and U18646 (N_18646,N_17771,N_18145);
nor U18647 (N_18647,N_17875,N_18153);
xnor U18648 (N_18648,N_18240,N_18165);
nand U18649 (N_18649,N_17977,N_18160);
nor U18650 (N_18650,N_17606,N_18110);
nor U18651 (N_18651,N_17942,N_17865);
and U18652 (N_18652,N_17800,N_18175);
and U18653 (N_18653,N_18291,N_17627);
or U18654 (N_18654,N_18001,N_17992);
nand U18655 (N_18655,N_17814,N_18340);
or U18656 (N_18656,N_17661,N_17874);
or U18657 (N_18657,N_17764,N_18168);
and U18658 (N_18658,N_18095,N_17723);
or U18659 (N_18659,N_17944,N_17618);
and U18660 (N_18660,N_18174,N_17989);
and U18661 (N_18661,N_17755,N_17987);
nand U18662 (N_18662,N_17707,N_17801);
nand U18663 (N_18663,N_17905,N_18182);
or U18664 (N_18664,N_17782,N_17762);
xor U18665 (N_18665,N_17774,N_18100);
xnor U18666 (N_18666,N_18303,N_18294);
nand U18667 (N_18667,N_18202,N_18043);
xor U18668 (N_18668,N_18339,N_18134);
xor U18669 (N_18669,N_18239,N_18192);
nand U18670 (N_18670,N_18146,N_17793);
xnor U18671 (N_18671,N_17727,N_17650);
or U18672 (N_18672,N_18333,N_17871);
nand U18673 (N_18673,N_17855,N_17939);
and U18674 (N_18674,N_17778,N_18357);
xor U18675 (N_18675,N_17683,N_18079);
nor U18676 (N_18676,N_18392,N_18238);
and U18677 (N_18677,N_18119,N_17885);
nor U18678 (N_18678,N_18167,N_18355);
or U18679 (N_18679,N_18004,N_17759);
or U18680 (N_18680,N_17657,N_17815);
or U18681 (N_18681,N_18332,N_18314);
and U18682 (N_18682,N_17997,N_18280);
nor U18683 (N_18683,N_17716,N_17957);
and U18684 (N_18684,N_17780,N_18096);
or U18685 (N_18685,N_18301,N_17692);
xor U18686 (N_18686,N_18114,N_18191);
nor U18687 (N_18687,N_17738,N_18384);
nor U18688 (N_18688,N_18386,N_18247);
and U18689 (N_18689,N_18176,N_17766);
nand U18690 (N_18690,N_17733,N_18059);
or U18691 (N_18691,N_17965,N_17678);
nor U18692 (N_18692,N_17809,N_18391);
nand U18693 (N_18693,N_18353,N_17669);
nand U18694 (N_18694,N_17798,N_17639);
or U18695 (N_18695,N_18372,N_18269);
nor U18696 (N_18696,N_18025,N_18117);
or U18697 (N_18697,N_17994,N_17884);
nor U18698 (N_18698,N_17784,N_17729);
nor U18699 (N_18699,N_17666,N_17847);
and U18700 (N_18700,N_17985,N_17930);
xor U18701 (N_18701,N_17876,N_18217);
xnor U18702 (N_18702,N_17956,N_17941);
and U18703 (N_18703,N_18011,N_17867);
or U18704 (N_18704,N_18312,N_17640);
nor U18705 (N_18705,N_17703,N_17953);
and U18706 (N_18706,N_18297,N_18309);
nor U18707 (N_18707,N_17777,N_18195);
nand U18708 (N_18708,N_17612,N_17658);
nor U18709 (N_18709,N_17971,N_18072);
and U18710 (N_18710,N_18124,N_17862);
and U18711 (N_18711,N_18262,N_17872);
nand U18712 (N_18712,N_18259,N_17927);
or U18713 (N_18713,N_18335,N_18315);
nand U18714 (N_18714,N_18152,N_17685);
nand U18715 (N_18715,N_17974,N_17779);
or U18716 (N_18716,N_18148,N_17629);
nor U18717 (N_18717,N_18199,N_17748);
and U18718 (N_18718,N_17715,N_17754);
nand U18719 (N_18719,N_17902,N_18128);
nor U18720 (N_18720,N_17951,N_17877);
and U18721 (N_18721,N_18067,N_17620);
nand U18722 (N_18722,N_17710,N_17742);
or U18723 (N_18723,N_17717,N_17899);
or U18724 (N_18724,N_17868,N_18246);
xor U18725 (N_18725,N_18205,N_17995);
or U18726 (N_18726,N_17955,N_18284);
or U18727 (N_18727,N_17901,N_18336);
and U18728 (N_18728,N_17626,N_18093);
nand U18729 (N_18729,N_17882,N_18367);
nand U18730 (N_18730,N_17817,N_18302);
or U18731 (N_18731,N_18027,N_17781);
and U18732 (N_18732,N_17665,N_18283);
nor U18733 (N_18733,N_18083,N_17812);
and U18734 (N_18734,N_17975,N_17735);
nor U18735 (N_18735,N_18188,N_18106);
and U18736 (N_18736,N_17756,N_18348);
and U18737 (N_18737,N_18102,N_18159);
xor U18738 (N_18738,N_18368,N_17631);
nand U18739 (N_18739,N_18116,N_18112);
nor U18740 (N_18740,N_17952,N_17740);
nand U18741 (N_18741,N_18264,N_17786);
and U18742 (N_18742,N_18054,N_17892);
nor U18743 (N_18743,N_17816,N_17917);
nand U18744 (N_18744,N_18158,N_17749);
xor U18745 (N_18745,N_18138,N_18024);
xor U18746 (N_18746,N_17841,N_18287);
nor U18747 (N_18747,N_17799,N_18052);
nor U18748 (N_18748,N_18288,N_18298);
or U18749 (N_18749,N_18326,N_18179);
or U18750 (N_18750,N_17870,N_17859);
nand U18751 (N_18751,N_18349,N_17961);
xor U18752 (N_18752,N_17763,N_17949);
or U18753 (N_18753,N_17873,N_17613);
and U18754 (N_18754,N_17935,N_18308);
or U18755 (N_18755,N_18131,N_17893);
xor U18756 (N_18756,N_17700,N_18197);
or U18757 (N_18757,N_18201,N_18313);
and U18758 (N_18758,N_18374,N_17680);
nand U18759 (N_18759,N_18076,N_18056);
or U18760 (N_18760,N_18077,N_17822);
nor U18761 (N_18761,N_17810,N_18049);
or U18762 (N_18762,N_18073,N_17796);
or U18763 (N_18763,N_18111,N_18107);
xnor U18764 (N_18764,N_17788,N_17787);
xor U18765 (N_18765,N_17659,N_18325);
nand U18766 (N_18766,N_18277,N_17846);
nor U18767 (N_18767,N_18233,N_17772);
nor U18768 (N_18768,N_17635,N_17726);
nor U18769 (N_18769,N_18008,N_17929);
nor U18770 (N_18770,N_17649,N_18173);
or U18771 (N_18771,N_17734,N_18218);
or U18772 (N_18772,N_17950,N_17761);
nor U18773 (N_18773,N_18180,N_18223);
or U18774 (N_18774,N_18237,N_18356);
and U18775 (N_18775,N_18351,N_18245);
nor U18776 (N_18776,N_18007,N_17684);
nand U18777 (N_18777,N_18172,N_18289);
or U18778 (N_18778,N_18380,N_18370);
and U18779 (N_18779,N_17769,N_18371);
nand U18780 (N_18780,N_18101,N_17844);
or U18781 (N_18781,N_17667,N_18185);
xnor U18782 (N_18782,N_18161,N_18317);
nor U18783 (N_18783,N_17993,N_17676);
and U18784 (N_18784,N_17760,N_17931);
nor U18785 (N_18785,N_18354,N_18307);
nor U18786 (N_18786,N_17911,N_18389);
or U18787 (N_18787,N_17732,N_18362);
nor U18788 (N_18788,N_17702,N_18021);
nor U18789 (N_18789,N_17982,N_18065);
xnor U18790 (N_18790,N_18219,N_17948);
and U18791 (N_18791,N_17698,N_17827);
nor U18792 (N_18792,N_18311,N_18190);
or U18793 (N_18793,N_18229,N_17645);
and U18794 (N_18794,N_18132,N_17856);
nor U18795 (N_18795,N_18249,N_18282);
xnor U18796 (N_18796,N_17802,N_17937);
or U18797 (N_18797,N_17746,N_18319);
nor U18798 (N_18798,N_17638,N_18346);
nand U18799 (N_18799,N_18381,N_18292);
xor U18800 (N_18800,N_18183,N_17875);
xnor U18801 (N_18801,N_18201,N_18059);
nand U18802 (N_18802,N_17989,N_18280);
nand U18803 (N_18803,N_18109,N_17939);
and U18804 (N_18804,N_17961,N_18260);
xor U18805 (N_18805,N_17888,N_18129);
nor U18806 (N_18806,N_17667,N_18194);
or U18807 (N_18807,N_17648,N_17944);
and U18808 (N_18808,N_18337,N_18145);
nor U18809 (N_18809,N_18363,N_17638);
and U18810 (N_18810,N_18202,N_18187);
xnor U18811 (N_18811,N_17767,N_18206);
or U18812 (N_18812,N_18157,N_17665);
xnor U18813 (N_18813,N_17709,N_18128);
or U18814 (N_18814,N_17698,N_18085);
and U18815 (N_18815,N_17896,N_18308);
or U18816 (N_18816,N_18303,N_18394);
nor U18817 (N_18817,N_17820,N_17924);
xnor U18818 (N_18818,N_17730,N_17704);
nor U18819 (N_18819,N_17860,N_18149);
and U18820 (N_18820,N_18394,N_18338);
xor U18821 (N_18821,N_18030,N_18239);
xor U18822 (N_18822,N_17636,N_18042);
or U18823 (N_18823,N_18126,N_17651);
xnor U18824 (N_18824,N_17930,N_17854);
xor U18825 (N_18825,N_18009,N_18032);
or U18826 (N_18826,N_17878,N_17762);
nand U18827 (N_18827,N_18180,N_17720);
nor U18828 (N_18828,N_18360,N_17922);
xnor U18829 (N_18829,N_17739,N_18324);
or U18830 (N_18830,N_17827,N_18260);
xor U18831 (N_18831,N_17866,N_17994);
nor U18832 (N_18832,N_18154,N_18168);
and U18833 (N_18833,N_18371,N_17963);
xor U18834 (N_18834,N_18132,N_18217);
nand U18835 (N_18835,N_17681,N_18274);
nand U18836 (N_18836,N_17867,N_18333);
and U18837 (N_18837,N_18002,N_17880);
nor U18838 (N_18838,N_18221,N_18391);
nand U18839 (N_18839,N_18308,N_18298);
xor U18840 (N_18840,N_17744,N_18302);
nor U18841 (N_18841,N_17801,N_18382);
nor U18842 (N_18842,N_17992,N_17809);
nor U18843 (N_18843,N_18238,N_18035);
nor U18844 (N_18844,N_18003,N_18280);
and U18845 (N_18845,N_18393,N_18011);
nand U18846 (N_18846,N_17676,N_18002);
xor U18847 (N_18847,N_18218,N_17874);
nand U18848 (N_18848,N_18168,N_18369);
and U18849 (N_18849,N_18057,N_17680);
nand U18850 (N_18850,N_17891,N_18105);
xnor U18851 (N_18851,N_17883,N_17773);
xor U18852 (N_18852,N_18368,N_17951);
nor U18853 (N_18853,N_18313,N_17825);
xnor U18854 (N_18854,N_17892,N_18341);
and U18855 (N_18855,N_17644,N_18222);
nand U18856 (N_18856,N_18296,N_18116);
or U18857 (N_18857,N_18179,N_17745);
and U18858 (N_18858,N_18119,N_17718);
or U18859 (N_18859,N_17633,N_18287);
xnor U18860 (N_18860,N_17725,N_18214);
and U18861 (N_18861,N_18336,N_18125);
xnor U18862 (N_18862,N_18054,N_17632);
xnor U18863 (N_18863,N_17970,N_18207);
or U18864 (N_18864,N_18321,N_17630);
and U18865 (N_18865,N_18302,N_17632);
nand U18866 (N_18866,N_18026,N_18257);
xor U18867 (N_18867,N_18040,N_18010);
nor U18868 (N_18868,N_17978,N_18029);
xnor U18869 (N_18869,N_17630,N_17657);
xor U18870 (N_18870,N_18293,N_18385);
nand U18871 (N_18871,N_18392,N_18004);
xor U18872 (N_18872,N_17632,N_17850);
xor U18873 (N_18873,N_17719,N_18195);
nand U18874 (N_18874,N_17971,N_17769);
nor U18875 (N_18875,N_18170,N_17856);
nand U18876 (N_18876,N_17602,N_17896);
or U18877 (N_18877,N_18212,N_18374);
and U18878 (N_18878,N_18149,N_18257);
and U18879 (N_18879,N_17987,N_18391);
xor U18880 (N_18880,N_17988,N_18166);
nand U18881 (N_18881,N_17984,N_18110);
and U18882 (N_18882,N_18274,N_17608);
nand U18883 (N_18883,N_18309,N_17870);
nor U18884 (N_18884,N_18103,N_18345);
nor U18885 (N_18885,N_18232,N_17844);
nor U18886 (N_18886,N_18049,N_17626);
nand U18887 (N_18887,N_18250,N_18272);
and U18888 (N_18888,N_18206,N_18040);
nand U18889 (N_18889,N_17890,N_18370);
or U18890 (N_18890,N_17905,N_18175);
and U18891 (N_18891,N_18059,N_18109);
xor U18892 (N_18892,N_18332,N_18354);
nor U18893 (N_18893,N_17844,N_17971);
xor U18894 (N_18894,N_18217,N_18098);
nand U18895 (N_18895,N_18255,N_18058);
nand U18896 (N_18896,N_18220,N_18180);
and U18897 (N_18897,N_18157,N_18116);
and U18898 (N_18898,N_17641,N_18170);
and U18899 (N_18899,N_17683,N_17931);
nor U18900 (N_18900,N_17987,N_17727);
and U18901 (N_18901,N_17750,N_18063);
and U18902 (N_18902,N_18082,N_17653);
xor U18903 (N_18903,N_17849,N_17738);
and U18904 (N_18904,N_18122,N_17847);
xnor U18905 (N_18905,N_17970,N_18058);
nor U18906 (N_18906,N_18390,N_18218);
xor U18907 (N_18907,N_18326,N_18095);
and U18908 (N_18908,N_17745,N_18399);
or U18909 (N_18909,N_17883,N_18355);
nand U18910 (N_18910,N_18384,N_17646);
xor U18911 (N_18911,N_18299,N_18003);
xnor U18912 (N_18912,N_18179,N_17716);
or U18913 (N_18913,N_17732,N_18319);
and U18914 (N_18914,N_18260,N_18155);
or U18915 (N_18915,N_18148,N_18389);
and U18916 (N_18916,N_17726,N_17622);
xor U18917 (N_18917,N_17732,N_18286);
nor U18918 (N_18918,N_17920,N_18328);
xor U18919 (N_18919,N_18001,N_18022);
nor U18920 (N_18920,N_17774,N_18115);
xnor U18921 (N_18921,N_17659,N_17773);
nor U18922 (N_18922,N_18238,N_18285);
xnor U18923 (N_18923,N_17624,N_18231);
and U18924 (N_18924,N_18312,N_18030);
xnor U18925 (N_18925,N_18061,N_18382);
nand U18926 (N_18926,N_18250,N_17819);
nor U18927 (N_18927,N_17909,N_17957);
and U18928 (N_18928,N_18292,N_18127);
xnor U18929 (N_18929,N_17857,N_18250);
xnor U18930 (N_18930,N_18298,N_18329);
nor U18931 (N_18931,N_17609,N_17779);
and U18932 (N_18932,N_18340,N_17654);
nor U18933 (N_18933,N_18060,N_17789);
and U18934 (N_18934,N_17878,N_17930);
nor U18935 (N_18935,N_18136,N_17694);
nor U18936 (N_18936,N_18252,N_18166);
nand U18937 (N_18937,N_17671,N_17668);
and U18938 (N_18938,N_18007,N_18160);
nand U18939 (N_18939,N_17632,N_18269);
nor U18940 (N_18940,N_18052,N_17646);
nor U18941 (N_18941,N_17698,N_18013);
nor U18942 (N_18942,N_17911,N_17895);
xor U18943 (N_18943,N_17743,N_17899);
and U18944 (N_18944,N_18154,N_17669);
and U18945 (N_18945,N_17921,N_18257);
or U18946 (N_18946,N_18149,N_17830);
or U18947 (N_18947,N_17966,N_17817);
and U18948 (N_18948,N_17815,N_17704);
nor U18949 (N_18949,N_17622,N_17813);
or U18950 (N_18950,N_17753,N_18149);
xnor U18951 (N_18951,N_18244,N_17853);
xnor U18952 (N_18952,N_18312,N_17719);
xnor U18953 (N_18953,N_18357,N_17646);
nand U18954 (N_18954,N_17878,N_18287);
nand U18955 (N_18955,N_18034,N_18102);
nand U18956 (N_18956,N_17974,N_18168);
xor U18957 (N_18957,N_18121,N_17876);
nand U18958 (N_18958,N_18154,N_18144);
and U18959 (N_18959,N_17811,N_17884);
or U18960 (N_18960,N_17690,N_18085);
or U18961 (N_18961,N_17721,N_17806);
xnor U18962 (N_18962,N_17803,N_17944);
nand U18963 (N_18963,N_17707,N_17771);
and U18964 (N_18964,N_17791,N_18049);
or U18965 (N_18965,N_17907,N_17609);
nor U18966 (N_18966,N_17871,N_17761);
nand U18967 (N_18967,N_17757,N_18053);
and U18968 (N_18968,N_17772,N_18318);
and U18969 (N_18969,N_18288,N_18178);
or U18970 (N_18970,N_18202,N_18065);
xor U18971 (N_18971,N_17810,N_17730);
or U18972 (N_18972,N_18258,N_17812);
nand U18973 (N_18973,N_18296,N_18249);
xnor U18974 (N_18974,N_17605,N_17651);
nand U18975 (N_18975,N_18134,N_17773);
or U18976 (N_18976,N_18364,N_17707);
or U18977 (N_18977,N_18006,N_18014);
nor U18978 (N_18978,N_17767,N_18050);
and U18979 (N_18979,N_18301,N_17783);
nand U18980 (N_18980,N_17907,N_17644);
xor U18981 (N_18981,N_18275,N_17661);
xnor U18982 (N_18982,N_17953,N_18123);
or U18983 (N_18983,N_17942,N_17985);
nand U18984 (N_18984,N_18352,N_18213);
nand U18985 (N_18985,N_18088,N_18171);
or U18986 (N_18986,N_17795,N_18328);
nand U18987 (N_18987,N_18361,N_17798);
xnor U18988 (N_18988,N_18106,N_18187);
or U18989 (N_18989,N_17978,N_17841);
and U18990 (N_18990,N_18252,N_18093);
nand U18991 (N_18991,N_17768,N_18343);
or U18992 (N_18992,N_18078,N_17680);
nand U18993 (N_18993,N_18045,N_18211);
nor U18994 (N_18994,N_18215,N_18237);
or U18995 (N_18995,N_17730,N_18058);
and U18996 (N_18996,N_18361,N_18300);
and U18997 (N_18997,N_17771,N_18069);
xor U18998 (N_18998,N_18018,N_18150);
and U18999 (N_18999,N_17843,N_17959);
or U19000 (N_19000,N_17924,N_17830);
and U19001 (N_19001,N_17907,N_18135);
xnor U19002 (N_19002,N_17944,N_17968);
nor U19003 (N_19003,N_18243,N_18378);
or U19004 (N_19004,N_18344,N_17974);
nor U19005 (N_19005,N_18229,N_17989);
and U19006 (N_19006,N_17750,N_18108);
and U19007 (N_19007,N_17852,N_17754);
nand U19008 (N_19008,N_17848,N_18101);
xor U19009 (N_19009,N_17948,N_17674);
xor U19010 (N_19010,N_18355,N_18034);
and U19011 (N_19011,N_18261,N_18026);
or U19012 (N_19012,N_18246,N_18248);
nand U19013 (N_19013,N_18369,N_17683);
and U19014 (N_19014,N_17923,N_17819);
or U19015 (N_19015,N_18100,N_18033);
or U19016 (N_19016,N_18130,N_17605);
and U19017 (N_19017,N_18145,N_18013);
or U19018 (N_19018,N_18294,N_18197);
nor U19019 (N_19019,N_18254,N_18069);
and U19020 (N_19020,N_17663,N_17944);
nor U19021 (N_19021,N_18151,N_18394);
or U19022 (N_19022,N_18017,N_17895);
nor U19023 (N_19023,N_17641,N_18265);
nand U19024 (N_19024,N_18298,N_18035);
nand U19025 (N_19025,N_17971,N_17642);
nand U19026 (N_19026,N_18228,N_17986);
nand U19027 (N_19027,N_17929,N_18292);
xor U19028 (N_19028,N_18020,N_17860);
xor U19029 (N_19029,N_18142,N_17624);
and U19030 (N_19030,N_17687,N_17716);
xnor U19031 (N_19031,N_18027,N_18062);
and U19032 (N_19032,N_17953,N_17706);
nor U19033 (N_19033,N_18050,N_18041);
nor U19034 (N_19034,N_17652,N_18213);
xnor U19035 (N_19035,N_18099,N_17614);
or U19036 (N_19036,N_17956,N_18227);
nand U19037 (N_19037,N_17942,N_17646);
nand U19038 (N_19038,N_17753,N_18003);
or U19039 (N_19039,N_18250,N_18301);
nor U19040 (N_19040,N_18358,N_18171);
and U19041 (N_19041,N_18099,N_17936);
nor U19042 (N_19042,N_18164,N_17637);
and U19043 (N_19043,N_18180,N_18222);
nand U19044 (N_19044,N_18089,N_18347);
nand U19045 (N_19045,N_17759,N_17939);
xor U19046 (N_19046,N_17800,N_17775);
nor U19047 (N_19047,N_17698,N_17768);
xor U19048 (N_19048,N_18155,N_18023);
nor U19049 (N_19049,N_18253,N_18266);
and U19050 (N_19050,N_18128,N_18327);
xor U19051 (N_19051,N_18011,N_18178);
nor U19052 (N_19052,N_18239,N_18236);
or U19053 (N_19053,N_17762,N_17605);
or U19054 (N_19054,N_18069,N_17926);
nand U19055 (N_19055,N_17924,N_17655);
nand U19056 (N_19056,N_18360,N_18048);
and U19057 (N_19057,N_18101,N_17924);
and U19058 (N_19058,N_17808,N_17761);
nand U19059 (N_19059,N_17610,N_17878);
nor U19060 (N_19060,N_17870,N_17906);
and U19061 (N_19061,N_18380,N_17879);
and U19062 (N_19062,N_18241,N_18233);
xnor U19063 (N_19063,N_17864,N_18351);
and U19064 (N_19064,N_18340,N_17697);
nand U19065 (N_19065,N_18243,N_17833);
xor U19066 (N_19066,N_18181,N_17908);
nand U19067 (N_19067,N_18109,N_18240);
or U19068 (N_19068,N_18174,N_18087);
nor U19069 (N_19069,N_18310,N_18359);
or U19070 (N_19070,N_17663,N_17648);
xor U19071 (N_19071,N_17681,N_18013);
nor U19072 (N_19072,N_18078,N_17919);
nand U19073 (N_19073,N_18061,N_18321);
nand U19074 (N_19074,N_17988,N_18151);
nor U19075 (N_19075,N_18224,N_18212);
and U19076 (N_19076,N_18045,N_18162);
and U19077 (N_19077,N_17866,N_17905);
nand U19078 (N_19078,N_18340,N_17801);
nand U19079 (N_19079,N_17607,N_18146);
nand U19080 (N_19080,N_17645,N_18336);
nor U19081 (N_19081,N_18350,N_17718);
xnor U19082 (N_19082,N_17914,N_18116);
and U19083 (N_19083,N_18151,N_18025);
nor U19084 (N_19084,N_18178,N_18089);
xnor U19085 (N_19085,N_18176,N_17925);
or U19086 (N_19086,N_17614,N_18219);
and U19087 (N_19087,N_17913,N_18128);
and U19088 (N_19088,N_18306,N_18144);
xor U19089 (N_19089,N_17880,N_17788);
or U19090 (N_19090,N_17955,N_18386);
nor U19091 (N_19091,N_17861,N_17968);
xor U19092 (N_19092,N_17893,N_18377);
nand U19093 (N_19093,N_18243,N_18369);
and U19094 (N_19094,N_18107,N_17669);
or U19095 (N_19095,N_17827,N_18058);
nand U19096 (N_19096,N_17940,N_17801);
and U19097 (N_19097,N_17817,N_17666);
nand U19098 (N_19098,N_18162,N_18032);
nor U19099 (N_19099,N_17926,N_18161);
and U19100 (N_19100,N_17702,N_18154);
xor U19101 (N_19101,N_18368,N_17814);
nor U19102 (N_19102,N_18008,N_17760);
or U19103 (N_19103,N_18110,N_18022);
or U19104 (N_19104,N_18344,N_17676);
nand U19105 (N_19105,N_17714,N_17773);
xor U19106 (N_19106,N_18082,N_18076);
or U19107 (N_19107,N_17746,N_18321);
and U19108 (N_19108,N_17843,N_18127);
xnor U19109 (N_19109,N_17932,N_17718);
and U19110 (N_19110,N_17855,N_18173);
nand U19111 (N_19111,N_18046,N_18004);
xor U19112 (N_19112,N_18117,N_18174);
or U19113 (N_19113,N_17961,N_17674);
or U19114 (N_19114,N_18121,N_18034);
or U19115 (N_19115,N_18131,N_17635);
xor U19116 (N_19116,N_17828,N_18122);
nor U19117 (N_19117,N_18299,N_17609);
and U19118 (N_19118,N_17648,N_18328);
nand U19119 (N_19119,N_17768,N_17800);
nand U19120 (N_19120,N_18044,N_18281);
nor U19121 (N_19121,N_18359,N_18058);
or U19122 (N_19122,N_17999,N_18337);
xor U19123 (N_19123,N_18167,N_17747);
nor U19124 (N_19124,N_17607,N_17671);
xor U19125 (N_19125,N_17703,N_18131);
or U19126 (N_19126,N_17730,N_18316);
and U19127 (N_19127,N_17756,N_17946);
xor U19128 (N_19128,N_17884,N_18188);
nor U19129 (N_19129,N_18395,N_18224);
and U19130 (N_19130,N_18355,N_17857);
or U19131 (N_19131,N_18270,N_18304);
nand U19132 (N_19132,N_18135,N_17796);
xor U19133 (N_19133,N_17865,N_18032);
nand U19134 (N_19134,N_17965,N_18146);
and U19135 (N_19135,N_18098,N_17742);
nand U19136 (N_19136,N_17780,N_18181);
nor U19137 (N_19137,N_18386,N_18342);
nand U19138 (N_19138,N_18069,N_18050);
nand U19139 (N_19139,N_17943,N_18366);
nand U19140 (N_19140,N_18268,N_17722);
nor U19141 (N_19141,N_18121,N_18096);
nand U19142 (N_19142,N_17908,N_17901);
and U19143 (N_19143,N_18331,N_17647);
and U19144 (N_19144,N_18361,N_17857);
xnor U19145 (N_19145,N_18279,N_18068);
or U19146 (N_19146,N_17713,N_17879);
xnor U19147 (N_19147,N_18320,N_17902);
xnor U19148 (N_19148,N_17707,N_18105);
and U19149 (N_19149,N_18156,N_18166);
xnor U19150 (N_19150,N_18398,N_18396);
nor U19151 (N_19151,N_17947,N_18227);
xor U19152 (N_19152,N_17702,N_17606);
and U19153 (N_19153,N_17604,N_18345);
xnor U19154 (N_19154,N_18009,N_17932);
nand U19155 (N_19155,N_17920,N_17623);
nor U19156 (N_19156,N_17817,N_18216);
nor U19157 (N_19157,N_18339,N_18072);
nor U19158 (N_19158,N_17789,N_18035);
nor U19159 (N_19159,N_18000,N_17915);
nand U19160 (N_19160,N_18263,N_17887);
and U19161 (N_19161,N_18295,N_18327);
nand U19162 (N_19162,N_18262,N_17679);
nor U19163 (N_19163,N_18048,N_17719);
xnor U19164 (N_19164,N_17679,N_17660);
and U19165 (N_19165,N_17761,N_17898);
xor U19166 (N_19166,N_18058,N_18247);
nand U19167 (N_19167,N_18208,N_17666);
or U19168 (N_19168,N_17991,N_17751);
xor U19169 (N_19169,N_18146,N_18236);
nor U19170 (N_19170,N_18022,N_18289);
or U19171 (N_19171,N_18351,N_18371);
nand U19172 (N_19172,N_18379,N_18386);
and U19173 (N_19173,N_18055,N_18338);
nand U19174 (N_19174,N_17980,N_17847);
nor U19175 (N_19175,N_17703,N_17712);
or U19176 (N_19176,N_17736,N_18132);
and U19177 (N_19177,N_17833,N_17789);
xnor U19178 (N_19178,N_18042,N_17661);
and U19179 (N_19179,N_17850,N_17727);
xor U19180 (N_19180,N_17628,N_18108);
or U19181 (N_19181,N_17697,N_17783);
nand U19182 (N_19182,N_18346,N_17643);
and U19183 (N_19183,N_18291,N_17955);
xnor U19184 (N_19184,N_18083,N_18088);
or U19185 (N_19185,N_18275,N_18033);
or U19186 (N_19186,N_17927,N_17747);
xor U19187 (N_19187,N_17925,N_18222);
xor U19188 (N_19188,N_18115,N_18307);
nor U19189 (N_19189,N_18235,N_17696);
nor U19190 (N_19190,N_17762,N_18180);
and U19191 (N_19191,N_17753,N_17849);
and U19192 (N_19192,N_18366,N_18340);
nor U19193 (N_19193,N_18207,N_18148);
or U19194 (N_19194,N_18093,N_17876);
nor U19195 (N_19195,N_18176,N_18034);
nor U19196 (N_19196,N_17635,N_17620);
or U19197 (N_19197,N_17983,N_17908);
nor U19198 (N_19198,N_18330,N_18048);
nor U19199 (N_19199,N_17712,N_18056);
nor U19200 (N_19200,N_19071,N_18831);
and U19201 (N_19201,N_18614,N_18669);
xnor U19202 (N_19202,N_18646,N_18571);
nor U19203 (N_19203,N_18937,N_19193);
or U19204 (N_19204,N_19163,N_18625);
or U19205 (N_19205,N_18678,N_19044);
nand U19206 (N_19206,N_18972,N_19050);
nand U19207 (N_19207,N_18554,N_18406);
and U19208 (N_19208,N_18570,N_18733);
or U19209 (N_19209,N_18963,N_18946);
xor U19210 (N_19210,N_19142,N_18843);
xnor U19211 (N_19211,N_19096,N_18433);
xor U19212 (N_19212,N_18504,N_19082);
nor U19213 (N_19213,N_18720,N_19107);
nor U19214 (N_19214,N_18470,N_18877);
or U19215 (N_19215,N_18777,N_19057);
or U19216 (N_19216,N_19131,N_18754);
and U19217 (N_19217,N_18649,N_19150);
or U19218 (N_19218,N_19144,N_18677);
nand U19219 (N_19219,N_18408,N_18612);
and U19220 (N_19220,N_18999,N_18621);
xor U19221 (N_19221,N_18435,N_18833);
nor U19222 (N_19222,N_18482,N_19058);
nor U19223 (N_19223,N_18726,N_18993);
nor U19224 (N_19224,N_18839,N_19175);
nand U19225 (N_19225,N_19184,N_19046);
or U19226 (N_19226,N_19034,N_18719);
and U19227 (N_19227,N_18431,N_18523);
or U19228 (N_19228,N_18893,N_18468);
nor U19229 (N_19229,N_18815,N_18905);
nor U19230 (N_19230,N_18842,N_18801);
or U19231 (N_19231,N_18871,N_18919);
nand U19232 (N_19232,N_19080,N_18863);
xor U19233 (N_19233,N_18542,N_19077);
or U19234 (N_19234,N_19174,N_19076);
and U19235 (N_19235,N_18721,N_18480);
nor U19236 (N_19236,N_18631,N_18786);
nor U19237 (N_19237,N_18981,N_18787);
or U19238 (N_19238,N_18692,N_18425);
or U19239 (N_19239,N_19191,N_18608);
or U19240 (N_19240,N_18686,N_18716);
xnor U19241 (N_19241,N_18577,N_18434);
nand U19242 (N_19242,N_18913,N_18615);
or U19243 (N_19243,N_18998,N_18463);
or U19244 (N_19244,N_18421,N_18970);
xnor U19245 (N_19245,N_18727,N_18783);
nand U19246 (N_19246,N_18918,N_18962);
or U19247 (N_19247,N_18763,N_18923);
nor U19248 (N_19248,N_18453,N_18792);
nor U19249 (N_19249,N_18524,N_18960);
or U19250 (N_19250,N_18740,N_19164);
nand U19251 (N_19251,N_18735,N_18888);
nor U19252 (N_19252,N_18860,N_18651);
and U19253 (N_19253,N_18867,N_18706);
nor U19254 (N_19254,N_18976,N_18618);
and U19255 (N_19255,N_18628,N_18613);
nand U19256 (N_19256,N_19014,N_18813);
nor U19257 (N_19257,N_18771,N_18619);
xnor U19258 (N_19258,N_19117,N_18683);
nor U19259 (N_19259,N_19104,N_19139);
and U19260 (N_19260,N_19137,N_18507);
or U19261 (N_19261,N_19012,N_18745);
nand U19262 (N_19262,N_18822,N_18797);
and U19263 (N_19263,N_19176,N_18642);
and U19264 (N_19264,N_18640,N_18698);
and U19265 (N_19265,N_18465,N_18685);
xnor U19266 (N_19266,N_19134,N_18714);
xnor U19267 (N_19267,N_18861,N_18729);
and U19268 (N_19268,N_18611,N_18670);
and U19269 (N_19269,N_18997,N_19157);
and U19270 (N_19270,N_18694,N_18782);
or U19271 (N_19271,N_18932,N_18812);
nor U19272 (N_19272,N_18410,N_18420);
and U19273 (N_19273,N_18730,N_19079);
xor U19274 (N_19274,N_18574,N_19083);
or U19275 (N_19275,N_18531,N_18665);
nand U19276 (N_19276,N_18658,N_18989);
and U19277 (N_19277,N_19023,N_18519);
and U19278 (N_19278,N_18681,N_18475);
or U19279 (N_19279,N_19149,N_19189);
or U19280 (N_19280,N_18580,N_19042);
xnor U19281 (N_19281,N_19030,N_18950);
xor U19282 (N_19282,N_19049,N_18679);
or U19283 (N_19283,N_18695,N_19089);
or U19284 (N_19284,N_19006,N_19052);
nand U19285 (N_19285,N_19119,N_19148);
nor U19286 (N_19286,N_19047,N_19099);
and U19287 (N_19287,N_18874,N_18832);
and U19288 (N_19288,N_18451,N_18557);
xor U19289 (N_19289,N_19078,N_18945);
nand U19290 (N_19290,N_18961,N_18447);
nand U19291 (N_19291,N_18939,N_18449);
nor U19292 (N_19292,N_18757,N_19158);
nand U19293 (N_19293,N_18973,N_19008);
and U19294 (N_19294,N_19130,N_19048);
and U19295 (N_19295,N_18700,N_18402);
xnor U19296 (N_19296,N_19198,N_18922);
xnor U19297 (N_19297,N_18485,N_18458);
xnor U19298 (N_19298,N_18423,N_18568);
xnor U19299 (N_19299,N_18750,N_18987);
xor U19300 (N_19300,N_18974,N_18811);
or U19301 (N_19301,N_19147,N_19098);
nand U19302 (N_19302,N_18545,N_18594);
and U19303 (N_19303,N_19040,N_18793);
xor U19304 (N_19304,N_19170,N_19112);
nand U19305 (N_19305,N_18701,N_19151);
and U19306 (N_19306,N_18428,N_18712);
and U19307 (N_19307,N_18713,N_18637);
or U19308 (N_19308,N_18567,N_18912);
xor U19309 (N_19309,N_18598,N_18857);
xnor U19310 (N_19310,N_18865,N_19154);
xnor U19311 (N_19311,N_18804,N_19140);
nand U19312 (N_19312,N_18559,N_18856);
and U19313 (N_19313,N_18538,N_18840);
nor U19314 (N_19314,N_19001,N_19016);
nand U19315 (N_19315,N_18710,N_18718);
xnor U19316 (N_19316,N_18702,N_18828);
or U19317 (N_19317,N_18588,N_18623);
nor U19318 (N_19318,N_19166,N_18941);
nor U19319 (N_19319,N_18823,N_19103);
or U19320 (N_19320,N_18606,N_18781);
nor U19321 (N_19321,N_19004,N_18816);
nor U19322 (N_19322,N_18599,N_18500);
and U19323 (N_19323,N_18483,N_19133);
xor U19324 (N_19324,N_18991,N_18491);
or U19325 (N_19325,N_18800,N_18841);
nor U19326 (N_19326,N_19114,N_18597);
nor U19327 (N_19327,N_18590,N_19186);
and U19328 (N_19328,N_18532,N_18432);
or U19329 (N_19329,N_18990,N_18654);
or U19330 (N_19330,N_18605,N_18897);
xnor U19331 (N_19331,N_18424,N_18688);
and U19332 (N_19332,N_19067,N_18810);
nand U19333 (N_19333,N_18521,N_18766);
nor U19334 (N_19334,N_18659,N_18759);
nand U19335 (N_19335,N_18928,N_18456);
or U19336 (N_19336,N_18547,N_19092);
and U19337 (N_19337,N_19177,N_18907);
nor U19338 (N_19338,N_18663,N_18587);
or U19339 (N_19339,N_18596,N_18838);
nor U19340 (N_19340,N_18761,N_18544);
nand U19341 (N_19341,N_18953,N_19038);
nor U19342 (N_19342,N_18904,N_18788);
nand U19343 (N_19343,N_18758,N_18650);
and U19344 (N_19344,N_18769,N_18940);
and U19345 (N_19345,N_19053,N_18555);
or U19346 (N_19346,N_18589,N_18887);
and U19347 (N_19347,N_19041,N_18473);
or U19348 (N_19348,N_18942,N_18563);
or U19349 (N_19349,N_19173,N_18952);
xor U19350 (N_19350,N_19102,N_18508);
nand U19351 (N_19351,N_18803,N_18772);
nor U19352 (N_19352,N_19036,N_19064);
or U19353 (N_19353,N_18964,N_19109);
nand U19354 (N_19354,N_19002,N_19187);
or U19355 (N_19355,N_18668,N_18417);
nand U19356 (N_19356,N_19074,N_18556);
nand U19357 (N_19357,N_18653,N_19097);
nand U19358 (N_19358,N_19156,N_18603);
xnor U19359 (N_19359,N_18418,N_19039);
and U19360 (N_19360,N_18566,N_18767);
or U19361 (N_19361,N_18807,N_18558);
xnor U19362 (N_19362,N_18440,N_18472);
or U19363 (N_19363,N_18495,N_18722);
nand U19364 (N_19364,N_18884,N_19160);
and U19365 (N_19365,N_18511,N_18864);
or U19366 (N_19366,N_18427,N_18490);
nand U19367 (N_19367,N_18443,N_18609);
xnor U19368 (N_19368,N_18725,N_18572);
xor U19369 (N_19369,N_18927,N_19009);
xnor U19370 (N_19370,N_19194,N_19121);
nand U19371 (N_19371,N_18466,N_19162);
and U19372 (N_19372,N_19141,N_18705);
nand U19373 (N_19373,N_18734,N_19172);
nand U19374 (N_19374,N_19059,N_18461);
nor U19375 (N_19375,N_18513,N_19105);
and U19376 (N_19376,N_18551,N_18667);
xor U19377 (N_19377,N_18641,N_18747);
nand U19378 (N_19378,N_18853,N_18858);
and U19379 (N_19379,N_19022,N_18586);
and U19380 (N_19380,N_18775,N_18814);
and U19381 (N_19381,N_18849,N_18824);
xnor U19382 (N_19382,N_19007,N_19120);
xor U19383 (N_19383,N_18908,N_19183);
nor U19384 (N_19384,N_18749,N_19110);
xnor U19385 (N_19385,N_19084,N_19086);
or U19386 (N_19386,N_18711,N_19122);
nand U19387 (N_19387,N_18446,N_18582);
or U19388 (N_19388,N_18562,N_18818);
nand U19389 (N_19389,N_18452,N_18617);
nand U19390 (N_19390,N_18806,N_18739);
nor U19391 (N_19391,N_18537,N_18929);
nor U19392 (N_19392,N_18966,N_19192);
xnor U19393 (N_19393,N_18916,N_18971);
nand U19394 (N_19394,N_18984,N_18549);
nand U19395 (N_19395,N_19095,N_18643);
or U19396 (N_19396,N_18415,N_18676);
nor U19397 (N_19397,N_19123,N_18690);
and U19398 (N_19398,N_18957,N_19199);
nand U19399 (N_19399,N_18835,N_18880);
nand U19400 (N_19400,N_18645,N_18959);
xnor U19401 (N_19401,N_19061,N_19015);
xnor U19402 (N_19402,N_18836,N_19181);
and U19403 (N_19403,N_18910,N_18883);
xor U19404 (N_19404,N_19182,N_18890);
nand U19405 (N_19405,N_18579,N_18419);
xor U19406 (N_19406,N_19088,N_19113);
xor U19407 (N_19407,N_18644,N_19135);
or U19408 (N_19408,N_18746,N_19178);
or U19409 (N_19409,N_18664,N_18911);
or U19410 (N_19410,N_18737,N_19037);
xnor U19411 (N_19411,N_19019,N_18829);
nor U19412 (N_19412,N_18809,N_18442);
xor U19413 (N_19413,N_19024,N_18752);
nand U19414 (N_19414,N_18827,N_18762);
or U19415 (N_19415,N_18462,N_18866);
and U19416 (N_19416,N_18936,N_18576);
xnor U19417 (N_19417,N_19020,N_18622);
xor U19418 (N_19418,N_18825,N_18675);
xnor U19419 (N_19419,N_18489,N_19115);
xnor U19420 (N_19420,N_18657,N_18467);
nor U19421 (N_19421,N_18915,N_19146);
and U19422 (N_19422,N_18411,N_18983);
nor U19423 (N_19423,N_18607,N_18779);
nand U19424 (N_19424,N_18691,N_18630);
and U19425 (N_19425,N_18847,N_18909);
nand U19426 (N_19426,N_18968,N_19118);
and U19427 (N_19427,N_18751,N_18851);
or U19428 (N_19428,N_18429,N_18503);
or U19429 (N_19429,N_19111,N_18448);
or U19430 (N_19430,N_18527,N_18776);
nor U19431 (N_19431,N_18768,N_18821);
or U19432 (N_19432,N_18765,N_18412);
or U19433 (N_19433,N_18436,N_18943);
and U19434 (N_19434,N_18454,N_18844);
and U19435 (N_19435,N_18684,N_18656);
and U19436 (N_19436,N_18707,N_18510);
xnor U19437 (N_19437,N_18926,N_18879);
and U19438 (N_19438,N_18553,N_18638);
nand U19439 (N_19439,N_19073,N_18891);
nor U19440 (N_19440,N_18591,N_19070);
nor U19441 (N_19441,N_18647,N_18982);
nand U19442 (N_19442,N_18994,N_18774);
or U19443 (N_19443,N_18539,N_19090);
xnor U19444 (N_19444,N_18868,N_18755);
xor U19445 (N_19445,N_18534,N_18409);
or U19446 (N_19446,N_19027,N_19188);
and U19447 (N_19447,N_18808,N_18403);
nand U19448 (N_19448,N_18703,N_18732);
or U19449 (N_19449,N_18789,N_18543);
xnor U19450 (N_19450,N_18660,N_19197);
or U19451 (N_19451,N_18487,N_18593);
nand U19452 (N_19452,N_18826,N_18512);
nor U19453 (N_19453,N_19017,N_19190);
and U19454 (N_19454,N_18837,N_18934);
or U19455 (N_19455,N_18846,N_18636);
and U19456 (N_19456,N_18575,N_18502);
and U19457 (N_19457,N_18986,N_18944);
xor U19458 (N_19458,N_19063,N_18977);
or U19459 (N_19459,N_18484,N_18834);
and U19460 (N_19460,N_19108,N_18995);
or U19461 (N_19461,N_18785,N_19005);
nor U19462 (N_19462,N_19101,N_19155);
nand U19463 (N_19463,N_18949,N_18492);
and U19464 (N_19464,N_18881,N_18457);
nor U19465 (N_19465,N_19126,N_19087);
and U19466 (N_19466,N_19195,N_18933);
xor U19467 (N_19467,N_19180,N_19179);
xor U19468 (N_19468,N_18439,N_18687);
xor U19469 (N_19469,N_19185,N_18756);
or U19470 (N_19470,N_18854,N_18980);
xor U19471 (N_19471,N_18460,N_19075);
nand U19472 (N_19472,N_19129,N_18478);
or U19473 (N_19473,N_18850,N_18535);
nand U19474 (N_19474,N_18680,N_18748);
and U19475 (N_19475,N_19029,N_18723);
xnor U19476 (N_19476,N_18796,N_18516);
xnor U19477 (N_19477,N_18820,N_18526);
nand U19478 (N_19478,N_18624,N_18903);
nand U19479 (N_19479,N_18954,N_18741);
nand U19480 (N_19480,N_18724,N_18947);
nand U19481 (N_19481,N_18548,N_18652);
xor U19482 (N_19482,N_19032,N_18405);
nand U19483 (N_19483,N_18655,N_18930);
xnor U19484 (N_19484,N_18525,N_18648);
and U19485 (N_19485,N_18560,N_18967);
nand U19486 (N_19486,N_18662,N_18931);
nor U19487 (N_19487,N_19116,N_18848);
xnor U19488 (N_19488,N_18498,N_19062);
nand U19489 (N_19489,N_18896,N_18780);
or U19490 (N_19490,N_19021,N_19026);
or U19491 (N_19491,N_18546,N_18885);
nand U19492 (N_19492,N_18764,N_18744);
and U19493 (N_19493,N_19011,N_19168);
and U19494 (N_19494,N_18802,N_18505);
xnor U19495 (N_19495,N_19165,N_18401);
nor U19496 (N_19496,N_18743,N_18682);
nor U19497 (N_19497,N_18499,N_18573);
and U19498 (N_19498,N_18906,N_18875);
and U19499 (N_19499,N_19106,N_18501);
xnor U19500 (N_19500,N_18552,N_18870);
xor U19501 (N_19501,N_18948,N_18770);
and U19502 (N_19502,N_19143,N_18469);
or U19503 (N_19503,N_19065,N_18529);
and U19504 (N_19504,N_19124,N_18697);
and U19505 (N_19505,N_18450,N_18496);
xor U19506 (N_19506,N_18958,N_19068);
nor U19507 (N_19507,N_18672,N_19169);
xor U19508 (N_19508,N_19069,N_19152);
or U19509 (N_19509,N_18773,N_18528);
nor U19510 (N_19510,N_18900,N_18699);
and U19511 (N_19511,N_18935,N_18855);
nand U19512 (N_19512,N_18520,N_18635);
or U19513 (N_19513,N_18515,N_19145);
xnor U19514 (N_19514,N_19028,N_18753);
nor U19515 (N_19515,N_18708,N_18717);
or U19516 (N_19516,N_19025,N_18541);
and U19517 (N_19517,N_18583,N_18476);
xnor U19518 (N_19518,N_19100,N_18561);
xor U19519 (N_19519,N_18494,N_18882);
xor U19520 (N_19520,N_18898,N_19132);
nor U19521 (N_19521,N_19013,N_18889);
nand U19522 (N_19522,N_19010,N_19161);
xor U19523 (N_19523,N_18444,N_18859);
and U19524 (N_19524,N_18601,N_19043);
and U19525 (N_19525,N_18627,N_18920);
nand U19526 (N_19526,N_19138,N_18862);
and U19527 (N_19527,N_18400,N_18517);
xnor U19528 (N_19528,N_18661,N_18459);
or U19529 (N_19529,N_19056,N_19093);
nand U19530 (N_19530,N_19060,N_19125);
or U19531 (N_19531,N_18988,N_18956);
and U19532 (N_19532,N_18709,N_18610);
and U19533 (N_19533,N_18778,N_18925);
or U19534 (N_19534,N_18924,N_18969);
xor U19535 (N_19535,N_18592,N_18715);
and U19536 (N_19536,N_19159,N_18486);
and U19537 (N_19537,N_19003,N_18581);
nor U19538 (N_19538,N_18634,N_18902);
nand U19539 (N_19539,N_18620,N_18892);
or U19540 (N_19540,N_18493,N_18530);
nor U19541 (N_19541,N_18985,N_18616);
or U19542 (N_19542,N_18869,N_18951);
nand U19543 (N_19543,N_19035,N_19196);
and U19544 (N_19544,N_18979,N_18938);
or U19545 (N_19545,N_19000,N_18407);
and U19546 (N_19546,N_18584,N_18790);
nand U19547 (N_19547,N_19167,N_18673);
nor U19548 (N_19548,N_18522,N_18564);
or U19549 (N_19549,N_18671,N_19136);
nand U19550 (N_19550,N_18817,N_18488);
xor U19551 (N_19551,N_18878,N_18872);
nor U19552 (N_19552,N_18550,N_18533);
nor U19553 (N_19553,N_18805,N_18438);
nor U19554 (N_19554,N_18819,N_18481);
xnor U19555 (N_19555,N_18799,N_18514);
or U19556 (N_19556,N_18600,N_19018);
and U19557 (N_19557,N_18917,N_18629);
xnor U19558 (N_19558,N_18895,N_18886);
xor U19559 (N_19559,N_18921,N_18540);
xor U19560 (N_19560,N_19094,N_19128);
or U19561 (N_19561,N_18633,N_18791);
or U19562 (N_19562,N_18742,N_18914);
xnor U19563 (N_19563,N_18728,N_18639);
xor U19564 (N_19564,N_19171,N_18738);
nor U19565 (N_19565,N_18992,N_18666);
xor U19566 (N_19566,N_19153,N_18894);
xor U19567 (N_19567,N_18901,N_18876);
nor U19568 (N_19568,N_18445,N_18852);
nand U19569 (N_19569,N_18696,N_18477);
xor U19570 (N_19570,N_19066,N_18565);
xor U19571 (N_19571,N_18497,N_18602);
xor U19572 (N_19572,N_18674,N_19045);
and U19573 (N_19573,N_18474,N_18585);
and U19574 (N_19574,N_18471,N_18955);
or U19575 (N_19575,N_19085,N_18595);
nor U19576 (N_19576,N_18578,N_18509);
nand U19577 (N_19577,N_18437,N_19033);
nand U19578 (N_19578,N_19051,N_18996);
xnor U19579 (N_19579,N_18798,N_18414);
or U19580 (N_19580,N_18416,N_19031);
and U19581 (N_19581,N_18704,N_19127);
nand U19582 (N_19582,N_18845,N_18760);
nand U19583 (N_19583,N_18975,N_18626);
or U19584 (N_19584,N_18413,N_18422);
xnor U19585 (N_19585,N_18536,N_18873);
or U19586 (N_19586,N_19054,N_18899);
nor U19587 (N_19587,N_18830,N_18430);
or U19588 (N_19588,N_18604,N_18689);
nor U19589 (N_19589,N_18795,N_19081);
nor U19590 (N_19590,N_18464,N_19072);
nor U19591 (N_19591,N_18404,N_18784);
nor U19592 (N_19592,N_18736,N_18506);
nor U19593 (N_19593,N_19091,N_18693);
xor U19594 (N_19594,N_18479,N_18632);
xnor U19595 (N_19595,N_18455,N_18569);
or U19596 (N_19596,N_18965,N_19055);
or U19597 (N_19597,N_18731,N_18978);
and U19598 (N_19598,N_18426,N_18518);
xnor U19599 (N_19599,N_18794,N_18441);
xnor U19600 (N_19600,N_18925,N_18443);
xor U19601 (N_19601,N_18479,N_18443);
xor U19602 (N_19602,N_18411,N_18537);
nand U19603 (N_19603,N_18648,N_18778);
nand U19604 (N_19604,N_18868,N_18635);
nor U19605 (N_19605,N_19093,N_18744);
or U19606 (N_19606,N_18547,N_18679);
and U19607 (N_19607,N_18804,N_18656);
nand U19608 (N_19608,N_18801,N_19056);
xnor U19609 (N_19609,N_19050,N_18756);
and U19610 (N_19610,N_18886,N_19049);
xor U19611 (N_19611,N_18480,N_18668);
xor U19612 (N_19612,N_18492,N_18674);
and U19613 (N_19613,N_18652,N_18808);
nor U19614 (N_19614,N_19194,N_18480);
xnor U19615 (N_19615,N_18442,N_19124);
nand U19616 (N_19616,N_18859,N_18991);
nor U19617 (N_19617,N_18572,N_18464);
and U19618 (N_19618,N_19049,N_18419);
nor U19619 (N_19619,N_18738,N_19137);
nor U19620 (N_19620,N_18934,N_18813);
and U19621 (N_19621,N_18471,N_19173);
nand U19622 (N_19622,N_19002,N_18822);
or U19623 (N_19623,N_19077,N_18890);
xnor U19624 (N_19624,N_18965,N_18898);
nand U19625 (N_19625,N_18651,N_18580);
nand U19626 (N_19626,N_18932,N_19047);
nor U19627 (N_19627,N_18446,N_18713);
xnor U19628 (N_19628,N_18918,N_18488);
nand U19629 (N_19629,N_18983,N_18639);
nor U19630 (N_19630,N_18873,N_18529);
nor U19631 (N_19631,N_18823,N_18950);
or U19632 (N_19632,N_18790,N_18999);
and U19633 (N_19633,N_19054,N_18942);
and U19634 (N_19634,N_18630,N_19022);
nor U19635 (N_19635,N_18501,N_18543);
nor U19636 (N_19636,N_18873,N_18544);
xnor U19637 (N_19637,N_18613,N_18744);
or U19638 (N_19638,N_18974,N_18857);
or U19639 (N_19639,N_18906,N_18636);
nor U19640 (N_19640,N_18844,N_18413);
or U19641 (N_19641,N_19054,N_19021);
xnor U19642 (N_19642,N_18653,N_19193);
nor U19643 (N_19643,N_18896,N_18654);
and U19644 (N_19644,N_18771,N_18898);
and U19645 (N_19645,N_18994,N_18548);
nor U19646 (N_19646,N_18963,N_18837);
and U19647 (N_19647,N_18567,N_19143);
xnor U19648 (N_19648,N_18461,N_18658);
or U19649 (N_19649,N_19036,N_18440);
nor U19650 (N_19650,N_18954,N_19097);
and U19651 (N_19651,N_19172,N_18856);
and U19652 (N_19652,N_18620,N_18664);
xnor U19653 (N_19653,N_18974,N_18703);
and U19654 (N_19654,N_18886,N_19063);
nor U19655 (N_19655,N_18581,N_18981);
xnor U19656 (N_19656,N_18518,N_19073);
xor U19657 (N_19657,N_19017,N_18657);
nand U19658 (N_19658,N_18610,N_18718);
and U19659 (N_19659,N_18764,N_18579);
and U19660 (N_19660,N_19132,N_18697);
xor U19661 (N_19661,N_18629,N_18701);
nor U19662 (N_19662,N_18713,N_18943);
xor U19663 (N_19663,N_18520,N_18782);
nor U19664 (N_19664,N_18816,N_18710);
and U19665 (N_19665,N_19012,N_18558);
and U19666 (N_19666,N_19114,N_18745);
nor U19667 (N_19667,N_19048,N_18734);
nand U19668 (N_19668,N_18997,N_18569);
xor U19669 (N_19669,N_18643,N_19011);
and U19670 (N_19670,N_19021,N_18554);
nor U19671 (N_19671,N_18914,N_19039);
nand U19672 (N_19672,N_18570,N_18944);
nor U19673 (N_19673,N_18834,N_18534);
nor U19674 (N_19674,N_18660,N_18917);
nand U19675 (N_19675,N_19044,N_18762);
and U19676 (N_19676,N_19097,N_19092);
nor U19677 (N_19677,N_18967,N_19102);
nand U19678 (N_19678,N_18913,N_18499);
xor U19679 (N_19679,N_18867,N_18618);
nor U19680 (N_19680,N_18657,N_18480);
nand U19681 (N_19681,N_19148,N_18777);
nor U19682 (N_19682,N_18499,N_18636);
nor U19683 (N_19683,N_19091,N_18523);
nand U19684 (N_19684,N_18861,N_18827);
nor U19685 (N_19685,N_18782,N_18810);
or U19686 (N_19686,N_18677,N_18666);
and U19687 (N_19687,N_18556,N_18728);
nor U19688 (N_19688,N_19025,N_18903);
or U19689 (N_19689,N_19043,N_18913);
and U19690 (N_19690,N_18571,N_19183);
nand U19691 (N_19691,N_18993,N_18825);
xor U19692 (N_19692,N_18700,N_18965);
nand U19693 (N_19693,N_18581,N_18421);
xnor U19694 (N_19694,N_19183,N_18912);
xnor U19695 (N_19695,N_18730,N_19036);
nand U19696 (N_19696,N_19161,N_18713);
xor U19697 (N_19697,N_18959,N_18668);
or U19698 (N_19698,N_19190,N_19035);
nor U19699 (N_19699,N_18911,N_18794);
and U19700 (N_19700,N_19153,N_18658);
nor U19701 (N_19701,N_18620,N_19136);
nand U19702 (N_19702,N_19027,N_18763);
nand U19703 (N_19703,N_18954,N_18565);
xnor U19704 (N_19704,N_18551,N_18600);
xor U19705 (N_19705,N_18794,N_18816);
nor U19706 (N_19706,N_18990,N_19127);
and U19707 (N_19707,N_19058,N_18764);
nor U19708 (N_19708,N_18966,N_18642);
nand U19709 (N_19709,N_18983,N_19191);
or U19710 (N_19710,N_18405,N_18878);
or U19711 (N_19711,N_18637,N_18543);
or U19712 (N_19712,N_18789,N_19001);
and U19713 (N_19713,N_19095,N_18619);
nand U19714 (N_19714,N_18812,N_19128);
nor U19715 (N_19715,N_18832,N_19026);
or U19716 (N_19716,N_18685,N_19038);
nor U19717 (N_19717,N_18758,N_18827);
or U19718 (N_19718,N_18489,N_18772);
and U19719 (N_19719,N_18564,N_18480);
nand U19720 (N_19720,N_18403,N_19181);
nand U19721 (N_19721,N_18730,N_18508);
nand U19722 (N_19722,N_18660,N_19175);
nand U19723 (N_19723,N_18804,N_19016);
nor U19724 (N_19724,N_18944,N_18661);
or U19725 (N_19725,N_19038,N_18493);
and U19726 (N_19726,N_18547,N_18662);
or U19727 (N_19727,N_18695,N_19165);
and U19728 (N_19728,N_19041,N_18992);
xnor U19729 (N_19729,N_18898,N_18810);
or U19730 (N_19730,N_18816,N_19177);
and U19731 (N_19731,N_18637,N_18706);
and U19732 (N_19732,N_18774,N_18825);
and U19733 (N_19733,N_19013,N_19068);
and U19734 (N_19734,N_18666,N_19001);
nor U19735 (N_19735,N_19003,N_19060);
and U19736 (N_19736,N_18429,N_18466);
or U19737 (N_19737,N_18477,N_18687);
and U19738 (N_19738,N_18459,N_19198);
xor U19739 (N_19739,N_18994,N_18519);
nor U19740 (N_19740,N_18594,N_18818);
nor U19741 (N_19741,N_18584,N_18835);
and U19742 (N_19742,N_19034,N_18710);
nor U19743 (N_19743,N_19080,N_18877);
xnor U19744 (N_19744,N_18825,N_18838);
nor U19745 (N_19745,N_18437,N_18609);
or U19746 (N_19746,N_18896,N_18746);
nand U19747 (N_19747,N_18499,N_19029);
nor U19748 (N_19748,N_18922,N_18616);
or U19749 (N_19749,N_18777,N_18955);
or U19750 (N_19750,N_19083,N_19169);
nand U19751 (N_19751,N_18404,N_18457);
xor U19752 (N_19752,N_18853,N_19081);
or U19753 (N_19753,N_19125,N_19170);
nand U19754 (N_19754,N_18659,N_19118);
nand U19755 (N_19755,N_19067,N_19198);
nor U19756 (N_19756,N_18937,N_18891);
nor U19757 (N_19757,N_18667,N_18758);
nand U19758 (N_19758,N_18951,N_18486);
xnor U19759 (N_19759,N_18733,N_18871);
nor U19760 (N_19760,N_18462,N_19056);
nor U19761 (N_19761,N_18676,N_18892);
nor U19762 (N_19762,N_18829,N_18426);
and U19763 (N_19763,N_18494,N_18499);
and U19764 (N_19764,N_18608,N_18740);
and U19765 (N_19765,N_18802,N_18568);
nor U19766 (N_19766,N_18809,N_19191);
xor U19767 (N_19767,N_18408,N_18963);
xnor U19768 (N_19768,N_18944,N_18995);
xnor U19769 (N_19769,N_18456,N_18771);
and U19770 (N_19770,N_18934,N_19027);
nand U19771 (N_19771,N_18778,N_18639);
nand U19772 (N_19772,N_18972,N_18722);
nand U19773 (N_19773,N_18868,N_18882);
or U19774 (N_19774,N_18840,N_18770);
xnor U19775 (N_19775,N_18505,N_19048);
nor U19776 (N_19776,N_19129,N_18759);
nand U19777 (N_19777,N_19028,N_18828);
or U19778 (N_19778,N_18749,N_18413);
or U19779 (N_19779,N_18868,N_18580);
nand U19780 (N_19780,N_19149,N_18591);
nand U19781 (N_19781,N_18500,N_18474);
or U19782 (N_19782,N_18898,N_18623);
xor U19783 (N_19783,N_18486,N_18536);
or U19784 (N_19784,N_18838,N_18433);
and U19785 (N_19785,N_18703,N_19124);
or U19786 (N_19786,N_18604,N_18415);
xnor U19787 (N_19787,N_18926,N_18451);
and U19788 (N_19788,N_18560,N_19181);
nand U19789 (N_19789,N_18818,N_18418);
xnor U19790 (N_19790,N_18660,N_18432);
nand U19791 (N_19791,N_19146,N_18595);
and U19792 (N_19792,N_18427,N_18861);
or U19793 (N_19793,N_18642,N_19009);
and U19794 (N_19794,N_18808,N_18749);
xor U19795 (N_19795,N_18475,N_18608);
nand U19796 (N_19796,N_18425,N_18568);
or U19797 (N_19797,N_18745,N_19172);
or U19798 (N_19798,N_18917,N_18934);
nor U19799 (N_19799,N_18765,N_19020);
nor U19800 (N_19800,N_18421,N_18545);
or U19801 (N_19801,N_18989,N_19133);
nand U19802 (N_19802,N_18607,N_19060);
or U19803 (N_19803,N_18898,N_18401);
nand U19804 (N_19804,N_18942,N_18856);
xnor U19805 (N_19805,N_18425,N_18989);
nor U19806 (N_19806,N_18835,N_18712);
xor U19807 (N_19807,N_19117,N_18618);
or U19808 (N_19808,N_19038,N_18733);
or U19809 (N_19809,N_18685,N_19011);
nor U19810 (N_19810,N_18786,N_18480);
nand U19811 (N_19811,N_18502,N_18485);
or U19812 (N_19812,N_18742,N_18505);
nor U19813 (N_19813,N_18455,N_18666);
nor U19814 (N_19814,N_18693,N_18465);
nor U19815 (N_19815,N_19133,N_18996);
or U19816 (N_19816,N_18660,N_18579);
nor U19817 (N_19817,N_19030,N_18543);
and U19818 (N_19818,N_18630,N_18485);
or U19819 (N_19819,N_19141,N_18429);
xor U19820 (N_19820,N_19170,N_19102);
or U19821 (N_19821,N_18448,N_18761);
nand U19822 (N_19822,N_18822,N_18940);
nor U19823 (N_19823,N_18933,N_18686);
xor U19824 (N_19824,N_18986,N_18941);
and U19825 (N_19825,N_19067,N_18821);
and U19826 (N_19826,N_19115,N_18583);
or U19827 (N_19827,N_18647,N_18764);
nor U19828 (N_19828,N_18455,N_18935);
nand U19829 (N_19829,N_18889,N_18636);
xnor U19830 (N_19830,N_18685,N_18609);
nor U19831 (N_19831,N_19002,N_18465);
or U19832 (N_19832,N_18642,N_18883);
nor U19833 (N_19833,N_18641,N_18997);
xnor U19834 (N_19834,N_19167,N_18521);
xnor U19835 (N_19835,N_18909,N_18903);
xor U19836 (N_19836,N_18605,N_18888);
or U19837 (N_19837,N_18800,N_18464);
or U19838 (N_19838,N_18735,N_18764);
and U19839 (N_19839,N_19099,N_19113);
xor U19840 (N_19840,N_18774,N_19125);
or U19841 (N_19841,N_18833,N_18795);
or U19842 (N_19842,N_18658,N_19198);
and U19843 (N_19843,N_18847,N_18546);
or U19844 (N_19844,N_18679,N_18856);
and U19845 (N_19845,N_18930,N_18937);
xor U19846 (N_19846,N_18804,N_18404);
nor U19847 (N_19847,N_18612,N_18980);
xor U19848 (N_19848,N_18717,N_18452);
nor U19849 (N_19849,N_19137,N_19128);
xor U19850 (N_19850,N_18848,N_18543);
nor U19851 (N_19851,N_18638,N_18897);
and U19852 (N_19852,N_18614,N_18496);
nor U19853 (N_19853,N_18897,N_18698);
xnor U19854 (N_19854,N_18541,N_18849);
nand U19855 (N_19855,N_18862,N_19018);
nand U19856 (N_19856,N_18442,N_18648);
xor U19857 (N_19857,N_19174,N_19195);
or U19858 (N_19858,N_18876,N_18999);
xnor U19859 (N_19859,N_18619,N_18513);
or U19860 (N_19860,N_18517,N_18975);
nand U19861 (N_19861,N_18716,N_18857);
xnor U19862 (N_19862,N_18761,N_18554);
xnor U19863 (N_19863,N_18894,N_18755);
xor U19864 (N_19864,N_19198,N_18417);
xor U19865 (N_19865,N_18439,N_18599);
xnor U19866 (N_19866,N_19175,N_18913);
or U19867 (N_19867,N_18543,N_19057);
and U19868 (N_19868,N_19180,N_19018);
nand U19869 (N_19869,N_18827,N_18578);
and U19870 (N_19870,N_18804,N_18650);
or U19871 (N_19871,N_18542,N_18859);
nor U19872 (N_19872,N_18741,N_18680);
nor U19873 (N_19873,N_18747,N_18975);
and U19874 (N_19874,N_18509,N_18582);
or U19875 (N_19875,N_18425,N_18751);
nand U19876 (N_19876,N_18532,N_19126);
nand U19877 (N_19877,N_18483,N_19067);
nand U19878 (N_19878,N_19013,N_18650);
or U19879 (N_19879,N_19128,N_18482);
nor U19880 (N_19880,N_18442,N_18786);
nand U19881 (N_19881,N_18586,N_18771);
or U19882 (N_19882,N_18634,N_18709);
or U19883 (N_19883,N_18981,N_18756);
nand U19884 (N_19884,N_18543,N_19166);
nand U19885 (N_19885,N_18623,N_18755);
xor U19886 (N_19886,N_18403,N_18828);
xnor U19887 (N_19887,N_19136,N_18634);
and U19888 (N_19888,N_18924,N_18777);
nor U19889 (N_19889,N_18472,N_18795);
xor U19890 (N_19890,N_18983,N_18833);
and U19891 (N_19891,N_18511,N_18891);
or U19892 (N_19892,N_18854,N_18760);
xor U19893 (N_19893,N_18590,N_19096);
nand U19894 (N_19894,N_19126,N_19028);
nor U19895 (N_19895,N_18999,N_18867);
and U19896 (N_19896,N_19146,N_19076);
nor U19897 (N_19897,N_18806,N_18519);
nor U19898 (N_19898,N_18941,N_19088);
or U19899 (N_19899,N_19062,N_18586);
nand U19900 (N_19900,N_18911,N_18489);
nor U19901 (N_19901,N_18464,N_18477);
nand U19902 (N_19902,N_18407,N_18974);
nor U19903 (N_19903,N_18833,N_18586);
xor U19904 (N_19904,N_18720,N_18540);
xor U19905 (N_19905,N_18865,N_18596);
xor U19906 (N_19906,N_18549,N_18799);
xnor U19907 (N_19907,N_18646,N_18985);
or U19908 (N_19908,N_18842,N_18829);
nand U19909 (N_19909,N_19134,N_18629);
and U19910 (N_19910,N_18580,N_18644);
or U19911 (N_19911,N_18543,N_19020);
nand U19912 (N_19912,N_18432,N_18656);
and U19913 (N_19913,N_19030,N_19044);
or U19914 (N_19914,N_19111,N_18755);
or U19915 (N_19915,N_18844,N_18407);
nor U19916 (N_19916,N_18848,N_19005);
nor U19917 (N_19917,N_18526,N_18704);
xnor U19918 (N_19918,N_18580,N_19113);
xor U19919 (N_19919,N_19130,N_18770);
nor U19920 (N_19920,N_18973,N_18934);
nor U19921 (N_19921,N_19109,N_18866);
or U19922 (N_19922,N_19118,N_18444);
or U19923 (N_19923,N_19101,N_18610);
nor U19924 (N_19924,N_18715,N_18531);
xor U19925 (N_19925,N_18897,N_18460);
or U19926 (N_19926,N_18437,N_18584);
nand U19927 (N_19927,N_19175,N_18470);
and U19928 (N_19928,N_19093,N_18643);
nor U19929 (N_19929,N_19041,N_18844);
nor U19930 (N_19930,N_18910,N_18804);
or U19931 (N_19931,N_18681,N_18543);
or U19932 (N_19932,N_19152,N_18657);
xnor U19933 (N_19933,N_18932,N_18749);
xnor U19934 (N_19934,N_18439,N_18572);
nor U19935 (N_19935,N_18952,N_18439);
nand U19936 (N_19936,N_19063,N_19168);
or U19937 (N_19937,N_18502,N_18835);
nor U19938 (N_19938,N_18690,N_18724);
xnor U19939 (N_19939,N_19181,N_19091);
xnor U19940 (N_19940,N_18894,N_19137);
nor U19941 (N_19941,N_18992,N_18754);
or U19942 (N_19942,N_19080,N_18405);
or U19943 (N_19943,N_18484,N_18416);
nor U19944 (N_19944,N_19102,N_18633);
nand U19945 (N_19945,N_18720,N_19193);
xor U19946 (N_19946,N_18464,N_18472);
and U19947 (N_19947,N_18907,N_18700);
nor U19948 (N_19948,N_19192,N_18654);
nor U19949 (N_19949,N_18744,N_18806);
xnor U19950 (N_19950,N_18764,N_18640);
and U19951 (N_19951,N_18416,N_18401);
or U19952 (N_19952,N_18436,N_19050);
nor U19953 (N_19953,N_19135,N_19156);
or U19954 (N_19954,N_19168,N_18457);
nor U19955 (N_19955,N_18942,N_18716);
xor U19956 (N_19956,N_18485,N_18760);
and U19957 (N_19957,N_18921,N_18691);
nor U19958 (N_19958,N_19088,N_18541);
or U19959 (N_19959,N_18913,N_18432);
and U19960 (N_19960,N_18592,N_18922);
or U19961 (N_19961,N_18494,N_18657);
nand U19962 (N_19962,N_19075,N_18682);
nand U19963 (N_19963,N_19058,N_18956);
nor U19964 (N_19964,N_18636,N_19051);
and U19965 (N_19965,N_18569,N_18915);
or U19966 (N_19966,N_18621,N_19162);
xnor U19967 (N_19967,N_18957,N_19197);
xnor U19968 (N_19968,N_19031,N_19101);
or U19969 (N_19969,N_18560,N_18786);
and U19970 (N_19970,N_18658,N_18577);
nor U19971 (N_19971,N_18524,N_19145);
and U19972 (N_19972,N_19016,N_18892);
nand U19973 (N_19973,N_18579,N_18453);
or U19974 (N_19974,N_18733,N_19060);
and U19975 (N_19975,N_19024,N_18856);
xor U19976 (N_19976,N_18511,N_18403);
nand U19977 (N_19977,N_19007,N_19000);
xor U19978 (N_19978,N_18464,N_19119);
xor U19979 (N_19979,N_18662,N_18558);
xnor U19980 (N_19980,N_18567,N_19094);
nand U19981 (N_19981,N_19186,N_19010);
and U19982 (N_19982,N_18769,N_18727);
and U19983 (N_19983,N_18846,N_18825);
and U19984 (N_19984,N_18635,N_18874);
and U19985 (N_19985,N_19165,N_19112);
nand U19986 (N_19986,N_18579,N_18998);
and U19987 (N_19987,N_18638,N_18755);
nand U19988 (N_19988,N_18808,N_18494);
or U19989 (N_19989,N_18509,N_18801);
nor U19990 (N_19990,N_18604,N_18735);
xor U19991 (N_19991,N_19170,N_19156);
and U19992 (N_19992,N_19067,N_18816);
and U19993 (N_19993,N_18732,N_18750);
or U19994 (N_19994,N_19050,N_18720);
nor U19995 (N_19995,N_18612,N_18723);
xnor U19996 (N_19996,N_18655,N_18627);
nand U19997 (N_19997,N_18645,N_18712);
xor U19998 (N_19998,N_18424,N_18748);
xor U19999 (N_19999,N_18742,N_19009);
nand UO_0 (O_0,N_19221,N_19672);
nor UO_1 (O_1,N_19649,N_19244);
and UO_2 (O_2,N_19571,N_19266);
nor UO_3 (O_3,N_19281,N_19291);
nand UO_4 (O_4,N_19771,N_19772);
or UO_5 (O_5,N_19653,N_19636);
or UO_6 (O_6,N_19233,N_19634);
nand UO_7 (O_7,N_19512,N_19617);
nor UO_8 (O_8,N_19396,N_19990);
nor UO_9 (O_9,N_19340,N_19353);
and UO_10 (O_10,N_19367,N_19782);
nand UO_11 (O_11,N_19766,N_19527);
nor UO_12 (O_12,N_19288,N_19324);
nand UO_13 (O_13,N_19648,N_19395);
nand UO_14 (O_14,N_19681,N_19478);
nor UO_15 (O_15,N_19502,N_19282);
xor UO_16 (O_16,N_19295,N_19469);
or UO_17 (O_17,N_19872,N_19615);
xnor UO_18 (O_18,N_19332,N_19850);
nor UO_19 (O_19,N_19948,N_19346);
and UO_20 (O_20,N_19548,N_19287);
and UO_21 (O_21,N_19616,N_19399);
or UO_22 (O_22,N_19865,N_19740);
and UO_23 (O_23,N_19977,N_19613);
xor UO_24 (O_24,N_19858,N_19581);
or UO_25 (O_25,N_19246,N_19430);
or UO_26 (O_26,N_19961,N_19981);
nand UO_27 (O_27,N_19700,N_19733);
or UO_28 (O_28,N_19480,N_19349);
nor UO_29 (O_29,N_19515,N_19953);
nor UO_30 (O_30,N_19524,N_19589);
or UO_31 (O_31,N_19878,N_19748);
or UO_32 (O_32,N_19808,N_19241);
nor UO_33 (O_33,N_19578,N_19505);
and UO_34 (O_34,N_19668,N_19759);
nand UO_35 (O_35,N_19744,N_19510);
xnor UO_36 (O_36,N_19939,N_19780);
or UO_37 (O_37,N_19454,N_19452);
or UO_38 (O_38,N_19864,N_19484);
nor UO_39 (O_39,N_19795,N_19910);
nand UO_40 (O_40,N_19262,N_19600);
nor UO_41 (O_41,N_19911,N_19936);
xor UO_42 (O_42,N_19713,N_19761);
nand UO_43 (O_43,N_19409,N_19568);
or UO_44 (O_44,N_19722,N_19929);
nand UO_45 (O_45,N_19473,N_19921);
xnor UO_46 (O_46,N_19493,N_19586);
xnor UO_47 (O_47,N_19680,N_19875);
nand UO_48 (O_48,N_19200,N_19488);
xor UO_49 (O_49,N_19645,N_19236);
or UO_50 (O_50,N_19552,N_19729);
or UO_51 (O_51,N_19408,N_19857);
nor UO_52 (O_52,N_19205,N_19542);
and UO_53 (O_53,N_19490,N_19877);
and UO_54 (O_54,N_19216,N_19279);
nor UO_55 (O_55,N_19224,N_19982);
nand UO_56 (O_56,N_19496,N_19323);
or UO_57 (O_57,N_19777,N_19688);
or UO_58 (O_58,N_19783,N_19882);
nand UO_59 (O_59,N_19687,N_19978);
nor UO_60 (O_60,N_19704,N_19614);
xnor UO_61 (O_61,N_19249,N_19776);
nor UO_62 (O_62,N_19667,N_19794);
xor UO_63 (O_63,N_19329,N_19689);
or UO_64 (O_64,N_19273,N_19392);
xnor UO_65 (O_65,N_19334,N_19504);
nor UO_66 (O_66,N_19758,N_19537);
and UO_67 (O_67,N_19724,N_19988);
or UO_68 (O_68,N_19419,N_19971);
nand UO_69 (O_69,N_19208,N_19458);
nand UO_70 (O_70,N_19253,N_19647);
nand UO_71 (O_71,N_19705,N_19923);
and UO_72 (O_72,N_19604,N_19342);
nand UO_73 (O_73,N_19931,N_19847);
xnor UO_74 (O_74,N_19973,N_19576);
or UO_75 (O_75,N_19312,N_19540);
nor UO_76 (O_76,N_19341,N_19550);
nand UO_77 (O_77,N_19546,N_19439);
nand UO_78 (O_78,N_19440,N_19453);
or UO_79 (O_79,N_19934,N_19558);
nor UO_80 (O_80,N_19394,N_19514);
nand UO_81 (O_81,N_19815,N_19886);
nand UO_82 (O_82,N_19644,N_19446);
nand UO_83 (O_83,N_19629,N_19796);
or UO_84 (O_84,N_19711,N_19400);
nor UO_85 (O_85,N_19624,N_19894);
or UO_86 (O_86,N_19709,N_19922);
nor UO_87 (O_87,N_19278,N_19431);
or UO_88 (O_88,N_19949,N_19827);
or UO_89 (O_89,N_19856,N_19582);
and UO_90 (O_90,N_19449,N_19966);
and UO_91 (O_91,N_19547,N_19300);
nor UO_92 (O_92,N_19914,N_19924);
or UO_93 (O_93,N_19250,N_19747);
nor UO_94 (O_94,N_19998,N_19657);
xor UO_95 (O_95,N_19401,N_19466);
or UO_96 (O_96,N_19954,N_19967);
nand UO_97 (O_97,N_19870,N_19225);
or UO_98 (O_98,N_19608,N_19209);
nor UO_99 (O_99,N_19927,N_19359);
xor UO_100 (O_100,N_19851,N_19674);
or UO_101 (O_101,N_19293,N_19306);
nand UO_102 (O_102,N_19481,N_19526);
nor UO_103 (O_103,N_19819,N_19317);
nand UO_104 (O_104,N_19360,N_19587);
xor UO_105 (O_105,N_19298,N_19880);
nand UO_106 (O_106,N_19785,N_19338);
xor UO_107 (O_107,N_19650,N_19790);
and UO_108 (O_108,N_19386,N_19612);
xnor UO_109 (O_109,N_19585,N_19773);
xor UO_110 (O_110,N_19946,N_19450);
xor UO_111 (O_111,N_19213,N_19402);
nor UO_112 (O_112,N_19665,N_19311);
or UO_113 (O_113,N_19844,N_19739);
xor UO_114 (O_114,N_19677,N_19623);
xor UO_115 (O_115,N_19701,N_19331);
xnor UO_116 (O_116,N_19326,N_19214);
and UO_117 (O_117,N_19730,N_19276);
or UO_118 (O_118,N_19974,N_19411);
and UO_119 (O_119,N_19919,N_19862);
xor UO_120 (O_120,N_19507,N_19917);
nor UO_121 (O_121,N_19980,N_19218);
nand UO_122 (O_122,N_19390,N_19398);
and UO_123 (O_123,N_19217,N_19373);
and UO_124 (O_124,N_19365,N_19849);
or UO_125 (O_125,N_19363,N_19479);
nor UO_126 (O_126,N_19621,N_19573);
or UO_127 (O_127,N_19348,N_19580);
nor UO_128 (O_128,N_19779,N_19935);
xor UO_129 (O_129,N_19654,N_19951);
nand UO_130 (O_130,N_19885,N_19516);
or UO_131 (O_131,N_19268,N_19405);
nand UO_132 (O_132,N_19567,N_19410);
or UO_133 (O_133,N_19545,N_19968);
and UO_134 (O_134,N_19610,N_19260);
xor UO_135 (O_135,N_19393,N_19406);
xnor UO_136 (O_136,N_19222,N_19603);
nor UO_137 (O_137,N_19442,N_19728);
and UO_138 (O_138,N_19383,N_19397);
nor UO_139 (O_139,N_19664,N_19381);
or UO_140 (O_140,N_19435,N_19319);
nor UO_141 (O_141,N_19223,N_19305);
nor UO_142 (O_142,N_19292,N_19918);
nand UO_143 (O_143,N_19330,N_19628);
and UO_144 (O_144,N_19774,N_19322);
xor UO_145 (O_145,N_19309,N_19908);
and UO_146 (O_146,N_19271,N_19434);
xor UO_147 (O_147,N_19474,N_19267);
nor UO_148 (O_148,N_19750,N_19735);
nand UO_149 (O_149,N_19963,N_19690);
nor UO_150 (O_150,N_19579,N_19420);
and UO_151 (O_151,N_19764,N_19391);
xor UO_152 (O_152,N_19798,N_19854);
nand UO_153 (O_153,N_19685,N_19660);
or UO_154 (O_154,N_19993,N_19652);
nand UO_155 (O_155,N_19595,N_19706);
xnor UO_156 (O_156,N_19712,N_19809);
xor UO_157 (O_157,N_19703,N_19226);
xor UO_158 (O_158,N_19684,N_19638);
nor UO_159 (O_159,N_19601,N_19767);
nand UO_160 (O_160,N_19942,N_19415);
nor UO_161 (O_161,N_19412,N_19955);
nand UO_162 (O_162,N_19792,N_19895);
or UO_163 (O_163,N_19832,N_19531);
or UO_164 (O_164,N_19591,N_19741);
or UO_165 (O_165,N_19307,N_19344);
or UO_166 (O_166,N_19762,N_19763);
nor UO_167 (O_167,N_19959,N_19830);
nor UO_168 (O_168,N_19743,N_19602);
or UO_169 (O_169,N_19482,N_19592);
or UO_170 (O_170,N_19495,N_19793);
nor UO_171 (O_171,N_19725,N_19727);
nor UO_172 (O_172,N_19925,N_19888);
or UO_173 (O_173,N_19708,N_19694);
xor UO_174 (O_174,N_19584,N_19569);
and UO_175 (O_175,N_19828,N_19433);
nor UO_176 (O_176,N_19755,N_19574);
nor UO_177 (O_177,N_19285,N_19497);
or UO_178 (O_178,N_19651,N_19263);
nand UO_179 (O_179,N_19786,N_19228);
nor UO_180 (O_180,N_19239,N_19544);
xor UO_181 (O_181,N_19572,N_19372);
nor UO_182 (O_182,N_19588,N_19598);
and UO_183 (O_183,N_19320,N_19656);
nand UO_184 (O_184,N_19721,N_19521);
xor UO_185 (O_185,N_19775,N_19891);
nor UO_186 (O_186,N_19807,N_19436);
or UO_187 (O_187,N_19388,N_19277);
xnor UO_188 (O_188,N_19655,N_19646);
nand UO_189 (O_189,N_19818,N_19867);
nand UO_190 (O_190,N_19884,N_19461);
xor UO_191 (O_191,N_19347,N_19803);
or UO_192 (O_192,N_19525,N_19445);
nand UO_193 (O_193,N_19302,N_19352);
nor UO_194 (O_194,N_19455,N_19898);
or UO_195 (O_195,N_19965,N_19290);
or UO_196 (O_196,N_19975,N_19806);
or UO_197 (O_197,N_19868,N_19843);
or UO_198 (O_198,N_19475,N_19389);
and UO_199 (O_199,N_19358,N_19999);
and UO_200 (O_200,N_19938,N_19642);
nor UO_201 (O_201,N_19506,N_19991);
or UO_202 (O_202,N_19429,N_19356);
or UO_203 (O_203,N_19248,N_19633);
or UO_204 (O_204,N_19594,N_19303);
nor UO_205 (O_205,N_19465,N_19781);
xor UO_206 (O_206,N_19355,N_19698);
nor UO_207 (O_207,N_19424,N_19380);
xor UO_208 (O_208,N_19622,N_19368);
nand UO_209 (O_209,N_19731,N_19964);
nand UO_210 (O_210,N_19259,N_19297);
or UO_211 (O_211,N_19416,N_19557);
and UO_212 (O_212,N_19866,N_19242);
nor UO_213 (O_213,N_19823,N_19538);
nor UO_214 (O_214,N_19247,N_19952);
or UO_215 (O_215,N_19881,N_19962);
or UO_216 (O_216,N_19810,N_19944);
and UO_217 (O_217,N_19212,N_19518);
xnor UO_218 (O_218,N_19575,N_19836);
or UO_219 (O_219,N_19619,N_19471);
xor UO_220 (O_220,N_19979,N_19464);
and UO_221 (O_221,N_19470,N_19631);
xor UO_222 (O_222,N_19673,N_19535);
nor UO_223 (O_223,N_19447,N_19905);
and UO_224 (O_224,N_19640,N_19369);
nand UO_225 (O_225,N_19520,N_19438);
or UO_226 (O_226,N_19985,N_19983);
or UO_227 (O_227,N_19984,N_19387);
xor UO_228 (O_228,N_19756,N_19996);
nor UO_229 (O_229,N_19742,N_19726);
nand UO_230 (O_230,N_19462,N_19749);
and UO_231 (O_231,N_19563,N_19534);
and UO_232 (O_232,N_19220,N_19354);
nand UO_233 (O_233,N_19425,N_19230);
or UO_234 (O_234,N_19351,N_19876);
and UO_235 (O_235,N_19824,N_19900);
xnor UO_236 (O_236,N_19530,N_19485);
nand UO_237 (O_237,N_19907,N_19328);
nor UO_238 (O_238,N_19835,N_19294);
nor UO_239 (O_239,N_19570,N_19893);
nor UO_240 (O_240,N_19760,N_19801);
and UO_241 (O_241,N_19219,N_19675);
and UO_242 (O_242,N_19997,N_19252);
and UO_243 (O_243,N_19564,N_19627);
or UO_244 (O_244,N_19753,N_19659);
or UO_245 (O_245,N_19956,N_19522);
or UO_246 (O_246,N_19852,N_19283);
nand UO_247 (O_247,N_19280,N_19467);
nor UO_248 (O_248,N_19626,N_19989);
and UO_249 (O_249,N_19498,N_19599);
and UO_250 (O_250,N_19313,N_19611);
xor UO_251 (O_251,N_19784,N_19337);
and UO_252 (O_252,N_19800,N_19970);
xor UO_253 (O_253,N_19765,N_19679);
nand UO_254 (O_254,N_19805,N_19707);
nand UO_255 (O_255,N_19816,N_19609);
or UO_256 (O_256,N_19734,N_19845);
or UO_257 (O_257,N_19301,N_19906);
nor UO_258 (O_258,N_19376,N_19732);
nor UO_259 (O_259,N_19915,N_19529);
or UO_260 (O_260,N_19833,N_19235);
xor UO_261 (O_261,N_19357,N_19940);
and UO_262 (O_262,N_19897,N_19903);
and UO_263 (O_263,N_19274,N_19270);
nand UO_264 (O_264,N_19620,N_19444);
nor UO_265 (O_265,N_19986,N_19362);
and UO_266 (O_266,N_19308,N_19503);
nor UO_267 (O_267,N_19590,N_19427);
and UO_268 (O_268,N_19932,N_19902);
and UO_269 (O_269,N_19375,N_19831);
or UO_270 (O_270,N_19896,N_19232);
and UO_271 (O_271,N_19366,N_19555);
or UO_272 (O_272,N_19799,N_19343);
or UO_273 (O_273,N_19720,N_19286);
and UO_274 (O_274,N_19451,N_19820);
nand UO_275 (O_275,N_19206,N_19203);
or UO_276 (O_276,N_19683,N_19577);
and UO_277 (O_277,N_19215,N_19487);
nand UO_278 (O_278,N_19251,N_19950);
and UO_279 (O_279,N_19201,N_19240);
xor UO_280 (O_280,N_19797,N_19682);
nor UO_281 (O_281,N_19335,N_19869);
and UO_282 (O_282,N_19607,N_19933);
xor UO_283 (O_283,N_19606,N_19842);
or UO_284 (O_284,N_19264,N_19987);
nor UO_285 (O_285,N_19318,N_19551);
xor UO_286 (O_286,N_19871,N_19539);
nand UO_287 (O_287,N_19432,N_19746);
or UO_288 (O_288,N_19691,N_19909);
xnor UO_289 (O_289,N_19255,N_19912);
and UO_290 (O_290,N_19846,N_19508);
and UO_291 (O_291,N_19715,N_19738);
nor UO_292 (O_292,N_19536,N_19463);
nor UO_293 (O_293,N_19477,N_19234);
nor UO_294 (O_294,N_19710,N_19460);
and UO_295 (O_295,N_19597,N_19926);
nor UO_296 (O_296,N_19549,N_19404);
nor UO_297 (O_297,N_19593,N_19204);
nand UO_298 (O_298,N_19812,N_19714);
or UO_299 (O_299,N_19519,N_19699);
or UO_300 (O_300,N_19834,N_19413);
and UO_301 (O_301,N_19254,N_19943);
or UO_302 (O_302,N_19829,N_19605);
or UO_303 (O_303,N_19556,N_19718);
nor UO_304 (O_304,N_19837,N_19848);
nor UO_305 (O_305,N_19422,N_19299);
nor UO_306 (O_306,N_19513,N_19855);
xor UO_307 (O_307,N_19364,N_19379);
nor UO_308 (O_308,N_19913,N_19227);
and UO_309 (O_309,N_19976,N_19757);
and UO_310 (O_310,N_19889,N_19237);
nand UO_311 (O_311,N_19258,N_19533);
xor UO_312 (O_312,N_19768,N_19314);
xnor UO_313 (O_313,N_19517,N_19202);
or UO_314 (O_314,N_19272,N_19890);
or UO_315 (O_315,N_19441,N_19560);
xnor UO_316 (O_316,N_19696,N_19669);
nand UO_317 (O_317,N_19899,N_19541);
xnor UO_318 (O_318,N_19418,N_19261);
nand UO_319 (O_319,N_19840,N_19378);
and UO_320 (O_320,N_19243,N_19632);
or UO_321 (O_321,N_19407,N_19284);
or UO_322 (O_322,N_19327,N_19414);
or UO_323 (O_323,N_19663,N_19625);
or UO_324 (O_324,N_19472,N_19554);
or UO_325 (O_325,N_19423,N_19385);
nor UO_326 (O_326,N_19822,N_19641);
xnor UO_327 (O_327,N_19316,N_19859);
and UO_328 (O_328,N_19321,N_19995);
xnor UO_329 (O_329,N_19863,N_19937);
xnor UO_330 (O_330,N_19930,N_19630);
and UO_331 (O_331,N_19804,N_19561);
nor UO_332 (O_332,N_19789,N_19377);
and UO_333 (O_333,N_19371,N_19325);
or UO_334 (O_334,N_19861,N_19838);
xnor UO_335 (O_335,N_19211,N_19821);
xnor UO_336 (O_336,N_19787,N_19511);
or UO_337 (O_337,N_19817,N_19639);
or UO_338 (O_338,N_19304,N_19994);
and UO_339 (O_339,N_19339,N_19662);
xor UO_340 (O_340,N_19879,N_19716);
nor UO_341 (O_341,N_19658,N_19565);
and UO_342 (O_342,N_19826,N_19443);
nor UO_343 (O_343,N_19374,N_19769);
nor UO_344 (O_344,N_19702,N_19637);
and UO_345 (O_345,N_19770,N_19670);
nand UO_346 (O_346,N_19509,N_19296);
nand UO_347 (O_347,N_19916,N_19210);
nand UO_348 (O_348,N_19839,N_19618);
nor UO_349 (O_349,N_19958,N_19841);
xor UO_350 (O_350,N_19231,N_19813);
or UO_351 (O_351,N_19972,N_19345);
and UO_352 (O_352,N_19494,N_19736);
nor UO_353 (O_353,N_19754,N_19491);
and UO_354 (O_354,N_19468,N_19957);
or UO_355 (O_355,N_19635,N_19583);
nand UO_356 (O_356,N_19437,N_19543);
nor UO_357 (O_357,N_19499,N_19256);
and UO_358 (O_358,N_19501,N_19860);
or UO_359 (O_359,N_19853,N_19887);
nor UO_360 (O_360,N_19814,N_19370);
xnor UO_361 (O_361,N_19457,N_19737);
or UO_362 (O_362,N_19350,N_19532);
and UO_363 (O_363,N_19486,N_19476);
nand UO_364 (O_364,N_19566,N_19553);
or UO_365 (O_365,N_19941,N_19920);
nor UO_366 (O_366,N_19945,N_19333);
nand UO_367 (O_367,N_19719,N_19265);
xnor UO_368 (O_368,N_19483,N_19238);
xor UO_369 (O_369,N_19969,N_19874);
nor UO_370 (O_370,N_19992,N_19417);
xnor UO_371 (O_371,N_19426,N_19289);
or UO_372 (O_372,N_19752,N_19928);
nor UO_373 (O_373,N_19257,N_19275);
nand UO_374 (O_374,N_19717,N_19661);
or UO_375 (O_375,N_19528,N_19315);
nand UO_376 (O_376,N_19456,N_19448);
xnor UO_377 (O_377,N_19676,N_19382);
or UO_378 (O_378,N_19791,N_19904);
nand UO_379 (O_379,N_19245,N_19751);
or UO_380 (O_380,N_19811,N_19459);
and UO_381 (O_381,N_19269,N_19802);
nor UO_382 (O_382,N_19596,N_19489);
xor UO_383 (O_383,N_19562,N_19421);
nand UO_384 (O_384,N_19873,N_19695);
and UO_385 (O_385,N_19947,N_19310);
xor UO_386 (O_386,N_19825,N_19336);
nor UO_387 (O_387,N_19403,N_19692);
xnor UO_388 (O_388,N_19523,N_19745);
and UO_389 (O_389,N_19671,N_19883);
nand UO_390 (O_390,N_19428,N_19723);
and UO_391 (O_391,N_19229,N_19778);
nand UO_392 (O_392,N_19892,N_19697);
or UO_393 (O_393,N_19686,N_19643);
nand UO_394 (O_394,N_19361,N_19500);
and UO_395 (O_395,N_19666,N_19788);
nor UO_396 (O_396,N_19901,N_19960);
or UO_397 (O_397,N_19559,N_19384);
and UO_398 (O_398,N_19492,N_19678);
or UO_399 (O_399,N_19693,N_19207);
nand UO_400 (O_400,N_19859,N_19488);
or UO_401 (O_401,N_19386,N_19492);
xor UO_402 (O_402,N_19352,N_19558);
nor UO_403 (O_403,N_19440,N_19213);
nand UO_404 (O_404,N_19719,N_19294);
nand UO_405 (O_405,N_19551,N_19874);
xnor UO_406 (O_406,N_19627,N_19601);
xnor UO_407 (O_407,N_19396,N_19959);
and UO_408 (O_408,N_19986,N_19281);
nand UO_409 (O_409,N_19982,N_19803);
and UO_410 (O_410,N_19537,N_19885);
xor UO_411 (O_411,N_19635,N_19940);
or UO_412 (O_412,N_19466,N_19764);
nor UO_413 (O_413,N_19314,N_19380);
or UO_414 (O_414,N_19373,N_19580);
or UO_415 (O_415,N_19436,N_19594);
nand UO_416 (O_416,N_19988,N_19759);
or UO_417 (O_417,N_19558,N_19826);
nand UO_418 (O_418,N_19400,N_19490);
nand UO_419 (O_419,N_19672,N_19663);
and UO_420 (O_420,N_19743,N_19772);
xor UO_421 (O_421,N_19935,N_19887);
nor UO_422 (O_422,N_19811,N_19881);
nor UO_423 (O_423,N_19783,N_19513);
nor UO_424 (O_424,N_19892,N_19703);
nand UO_425 (O_425,N_19528,N_19878);
nor UO_426 (O_426,N_19792,N_19460);
nand UO_427 (O_427,N_19374,N_19694);
or UO_428 (O_428,N_19536,N_19894);
nor UO_429 (O_429,N_19951,N_19947);
xor UO_430 (O_430,N_19678,N_19742);
xor UO_431 (O_431,N_19466,N_19235);
and UO_432 (O_432,N_19774,N_19896);
and UO_433 (O_433,N_19427,N_19613);
nor UO_434 (O_434,N_19965,N_19448);
nand UO_435 (O_435,N_19796,N_19404);
or UO_436 (O_436,N_19694,N_19654);
nor UO_437 (O_437,N_19750,N_19209);
nand UO_438 (O_438,N_19721,N_19288);
nand UO_439 (O_439,N_19524,N_19683);
xor UO_440 (O_440,N_19295,N_19390);
or UO_441 (O_441,N_19419,N_19519);
and UO_442 (O_442,N_19690,N_19781);
or UO_443 (O_443,N_19558,N_19674);
xor UO_444 (O_444,N_19433,N_19410);
nand UO_445 (O_445,N_19448,N_19917);
nand UO_446 (O_446,N_19689,N_19269);
or UO_447 (O_447,N_19261,N_19796);
nor UO_448 (O_448,N_19626,N_19900);
nor UO_449 (O_449,N_19219,N_19207);
xor UO_450 (O_450,N_19535,N_19244);
xor UO_451 (O_451,N_19614,N_19266);
xor UO_452 (O_452,N_19898,N_19625);
or UO_453 (O_453,N_19904,N_19928);
or UO_454 (O_454,N_19304,N_19914);
xor UO_455 (O_455,N_19748,N_19367);
xnor UO_456 (O_456,N_19315,N_19737);
or UO_457 (O_457,N_19627,N_19617);
and UO_458 (O_458,N_19482,N_19652);
nand UO_459 (O_459,N_19463,N_19224);
nor UO_460 (O_460,N_19614,N_19243);
or UO_461 (O_461,N_19492,N_19318);
or UO_462 (O_462,N_19749,N_19751);
nor UO_463 (O_463,N_19519,N_19755);
nor UO_464 (O_464,N_19239,N_19832);
or UO_465 (O_465,N_19720,N_19994);
nand UO_466 (O_466,N_19913,N_19868);
nor UO_467 (O_467,N_19736,N_19983);
and UO_468 (O_468,N_19840,N_19652);
nand UO_469 (O_469,N_19349,N_19706);
nand UO_470 (O_470,N_19473,N_19521);
and UO_471 (O_471,N_19252,N_19717);
xnor UO_472 (O_472,N_19896,N_19664);
xnor UO_473 (O_473,N_19395,N_19708);
xnor UO_474 (O_474,N_19583,N_19981);
nand UO_475 (O_475,N_19504,N_19993);
nand UO_476 (O_476,N_19257,N_19321);
or UO_477 (O_477,N_19507,N_19301);
xnor UO_478 (O_478,N_19248,N_19450);
xnor UO_479 (O_479,N_19568,N_19540);
or UO_480 (O_480,N_19677,N_19716);
xor UO_481 (O_481,N_19227,N_19918);
xnor UO_482 (O_482,N_19847,N_19745);
nor UO_483 (O_483,N_19320,N_19227);
xor UO_484 (O_484,N_19955,N_19622);
nor UO_485 (O_485,N_19406,N_19712);
or UO_486 (O_486,N_19587,N_19775);
xor UO_487 (O_487,N_19220,N_19977);
and UO_488 (O_488,N_19807,N_19549);
xor UO_489 (O_489,N_19428,N_19631);
nand UO_490 (O_490,N_19414,N_19343);
xor UO_491 (O_491,N_19412,N_19882);
nand UO_492 (O_492,N_19281,N_19515);
or UO_493 (O_493,N_19270,N_19682);
and UO_494 (O_494,N_19627,N_19415);
nor UO_495 (O_495,N_19880,N_19939);
and UO_496 (O_496,N_19808,N_19800);
or UO_497 (O_497,N_19447,N_19552);
nor UO_498 (O_498,N_19410,N_19587);
nor UO_499 (O_499,N_19498,N_19586);
and UO_500 (O_500,N_19235,N_19444);
nor UO_501 (O_501,N_19718,N_19512);
nand UO_502 (O_502,N_19541,N_19581);
nand UO_503 (O_503,N_19460,N_19248);
or UO_504 (O_504,N_19918,N_19606);
and UO_505 (O_505,N_19590,N_19845);
xor UO_506 (O_506,N_19651,N_19774);
xnor UO_507 (O_507,N_19852,N_19786);
xor UO_508 (O_508,N_19623,N_19995);
and UO_509 (O_509,N_19229,N_19434);
nor UO_510 (O_510,N_19242,N_19699);
nor UO_511 (O_511,N_19702,N_19577);
and UO_512 (O_512,N_19988,N_19781);
xnor UO_513 (O_513,N_19275,N_19351);
and UO_514 (O_514,N_19934,N_19940);
nand UO_515 (O_515,N_19355,N_19984);
xnor UO_516 (O_516,N_19325,N_19277);
nand UO_517 (O_517,N_19542,N_19680);
and UO_518 (O_518,N_19472,N_19325);
xor UO_519 (O_519,N_19304,N_19666);
and UO_520 (O_520,N_19720,N_19285);
or UO_521 (O_521,N_19860,N_19801);
nand UO_522 (O_522,N_19579,N_19641);
nand UO_523 (O_523,N_19564,N_19253);
nand UO_524 (O_524,N_19215,N_19619);
xor UO_525 (O_525,N_19485,N_19520);
xnor UO_526 (O_526,N_19223,N_19997);
or UO_527 (O_527,N_19334,N_19947);
nand UO_528 (O_528,N_19671,N_19896);
nand UO_529 (O_529,N_19605,N_19487);
nor UO_530 (O_530,N_19781,N_19889);
xor UO_531 (O_531,N_19903,N_19404);
and UO_532 (O_532,N_19458,N_19941);
nor UO_533 (O_533,N_19812,N_19790);
xor UO_534 (O_534,N_19775,N_19481);
and UO_535 (O_535,N_19718,N_19623);
nor UO_536 (O_536,N_19442,N_19426);
xor UO_537 (O_537,N_19819,N_19563);
and UO_538 (O_538,N_19489,N_19969);
nand UO_539 (O_539,N_19705,N_19800);
or UO_540 (O_540,N_19321,N_19202);
nand UO_541 (O_541,N_19512,N_19582);
or UO_542 (O_542,N_19979,N_19592);
and UO_543 (O_543,N_19974,N_19533);
xnor UO_544 (O_544,N_19205,N_19211);
nand UO_545 (O_545,N_19539,N_19441);
nor UO_546 (O_546,N_19270,N_19368);
nand UO_547 (O_547,N_19703,N_19474);
nand UO_548 (O_548,N_19200,N_19226);
nand UO_549 (O_549,N_19204,N_19832);
and UO_550 (O_550,N_19458,N_19806);
and UO_551 (O_551,N_19636,N_19948);
xor UO_552 (O_552,N_19232,N_19964);
or UO_553 (O_553,N_19584,N_19765);
or UO_554 (O_554,N_19819,N_19222);
or UO_555 (O_555,N_19773,N_19894);
nor UO_556 (O_556,N_19269,N_19241);
or UO_557 (O_557,N_19792,N_19396);
nor UO_558 (O_558,N_19837,N_19960);
and UO_559 (O_559,N_19670,N_19881);
or UO_560 (O_560,N_19500,N_19593);
nor UO_561 (O_561,N_19979,N_19653);
or UO_562 (O_562,N_19400,N_19432);
nand UO_563 (O_563,N_19457,N_19892);
nor UO_564 (O_564,N_19272,N_19222);
and UO_565 (O_565,N_19601,N_19228);
xnor UO_566 (O_566,N_19327,N_19835);
xnor UO_567 (O_567,N_19756,N_19855);
xor UO_568 (O_568,N_19307,N_19582);
or UO_569 (O_569,N_19231,N_19287);
nor UO_570 (O_570,N_19858,N_19407);
nand UO_571 (O_571,N_19520,N_19266);
nor UO_572 (O_572,N_19785,N_19910);
and UO_573 (O_573,N_19540,N_19871);
xnor UO_574 (O_574,N_19394,N_19309);
and UO_575 (O_575,N_19948,N_19828);
nand UO_576 (O_576,N_19623,N_19717);
xnor UO_577 (O_577,N_19388,N_19786);
xnor UO_578 (O_578,N_19271,N_19218);
xor UO_579 (O_579,N_19877,N_19864);
xor UO_580 (O_580,N_19783,N_19385);
or UO_581 (O_581,N_19855,N_19356);
nand UO_582 (O_582,N_19762,N_19269);
xor UO_583 (O_583,N_19590,N_19739);
and UO_584 (O_584,N_19902,N_19502);
and UO_585 (O_585,N_19631,N_19863);
nand UO_586 (O_586,N_19389,N_19503);
nand UO_587 (O_587,N_19914,N_19349);
nand UO_588 (O_588,N_19887,N_19985);
nor UO_589 (O_589,N_19738,N_19912);
xnor UO_590 (O_590,N_19408,N_19924);
and UO_591 (O_591,N_19947,N_19770);
or UO_592 (O_592,N_19848,N_19428);
and UO_593 (O_593,N_19726,N_19263);
and UO_594 (O_594,N_19850,N_19290);
xnor UO_595 (O_595,N_19364,N_19744);
nor UO_596 (O_596,N_19565,N_19238);
nand UO_597 (O_597,N_19423,N_19518);
xnor UO_598 (O_598,N_19977,N_19810);
and UO_599 (O_599,N_19245,N_19417);
or UO_600 (O_600,N_19436,N_19264);
or UO_601 (O_601,N_19338,N_19428);
or UO_602 (O_602,N_19533,N_19850);
and UO_603 (O_603,N_19819,N_19877);
and UO_604 (O_604,N_19223,N_19739);
xor UO_605 (O_605,N_19972,N_19463);
or UO_606 (O_606,N_19754,N_19402);
xor UO_607 (O_607,N_19772,N_19605);
or UO_608 (O_608,N_19409,N_19509);
nand UO_609 (O_609,N_19679,N_19618);
and UO_610 (O_610,N_19431,N_19561);
xnor UO_611 (O_611,N_19561,N_19613);
nor UO_612 (O_612,N_19469,N_19488);
or UO_613 (O_613,N_19355,N_19962);
nand UO_614 (O_614,N_19373,N_19974);
nor UO_615 (O_615,N_19826,N_19970);
nand UO_616 (O_616,N_19880,N_19786);
or UO_617 (O_617,N_19944,N_19619);
or UO_618 (O_618,N_19694,N_19338);
nor UO_619 (O_619,N_19861,N_19386);
xnor UO_620 (O_620,N_19542,N_19501);
or UO_621 (O_621,N_19684,N_19464);
nor UO_622 (O_622,N_19797,N_19425);
xor UO_623 (O_623,N_19870,N_19650);
nand UO_624 (O_624,N_19435,N_19921);
or UO_625 (O_625,N_19917,N_19646);
and UO_626 (O_626,N_19610,N_19300);
xor UO_627 (O_627,N_19841,N_19456);
nor UO_628 (O_628,N_19586,N_19796);
nor UO_629 (O_629,N_19969,N_19369);
or UO_630 (O_630,N_19460,N_19750);
or UO_631 (O_631,N_19501,N_19275);
xor UO_632 (O_632,N_19662,N_19649);
nand UO_633 (O_633,N_19735,N_19334);
or UO_634 (O_634,N_19835,N_19288);
or UO_635 (O_635,N_19668,N_19985);
nand UO_636 (O_636,N_19203,N_19719);
nor UO_637 (O_637,N_19718,N_19815);
nand UO_638 (O_638,N_19689,N_19944);
nand UO_639 (O_639,N_19996,N_19269);
or UO_640 (O_640,N_19654,N_19473);
nor UO_641 (O_641,N_19990,N_19832);
and UO_642 (O_642,N_19771,N_19752);
and UO_643 (O_643,N_19939,N_19973);
nand UO_644 (O_644,N_19816,N_19826);
nand UO_645 (O_645,N_19648,N_19830);
and UO_646 (O_646,N_19305,N_19685);
nor UO_647 (O_647,N_19595,N_19270);
xor UO_648 (O_648,N_19700,N_19819);
xnor UO_649 (O_649,N_19883,N_19503);
xor UO_650 (O_650,N_19485,N_19588);
or UO_651 (O_651,N_19516,N_19348);
xor UO_652 (O_652,N_19635,N_19381);
or UO_653 (O_653,N_19887,N_19581);
nor UO_654 (O_654,N_19876,N_19832);
xor UO_655 (O_655,N_19348,N_19382);
and UO_656 (O_656,N_19297,N_19542);
xor UO_657 (O_657,N_19207,N_19932);
nand UO_658 (O_658,N_19908,N_19556);
and UO_659 (O_659,N_19482,N_19885);
nor UO_660 (O_660,N_19680,N_19425);
nor UO_661 (O_661,N_19249,N_19697);
nor UO_662 (O_662,N_19878,N_19240);
nand UO_663 (O_663,N_19876,N_19999);
nor UO_664 (O_664,N_19261,N_19723);
and UO_665 (O_665,N_19634,N_19783);
or UO_666 (O_666,N_19296,N_19580);
xnor UO_667 (O_667,N_19794,N_19872);
or UO_668 (O_668,N_19690,N_19733);
or UO_669 (O_669,N_19835,N_19586);
or UO_670 (O_670,N_19858,N_19483);
and UO_671 (O_671,N_19463,N_19487);
xor UO_672 (O_672,N_19284,N_19794);
and UO_673 (O_673,N_19551,N_19581);
and UO_674 (O_674,N_19691,N_19865);
nand UO_675 (O_675,N_19727,N_19232);
xnor UO_676 (O_676,N_19881,N_19901);
nand UO_677 (O_677,N_19773,N_19223);
or UO_678 (O_678,N_19710,N_19897);
and UO_679 (O_679,N_19569,N_19316);
nor UO_680 (O_680,N_19817,N_19569);
or UO_681 (O_681,N_19356,N_19472);
nand UO_682 (O_682,N_19593,N_19214);
or UO_683 (O_683,N_19536,N_19235);
and UO_684 (O_684,N_19785,N_19473);
nand UO_685 (O_685,N_19897,N_19511);
and UO_686 (O_686,N_19889,N_19566);
nor UO_687 (O_687,N_19773,N_19438);
and UO_688 (O_688,N_19692,N_19539);
nor UO_689 (O_689,N_19411,N_19719);
xnor UO_690 (O_690,N_19550,N_19206);
nor UO_691 (O_691,N_19382,N_19422);
nand UO_692 (O_692,N_19758,N_19568);
and UO_693 (O_693,N_19591,N_19607);
xor UO_694 (O_694,N_19627,N_19581);
and UO_695 (O_695,N_19761,N_19235);
nor UO_696 (O_696,N_19616,N_19613);
and UO_697 (O_697,N_19716,N_19570);
nor UO_698 (O_698,N_19519,N_19816);
or UO_699 (O_699,N_19319,N_19814);
nor UO_700 (O_700,N_19623,N_19284);
nand UO_701 (O_701,N_19500,N_19386);
nand UO_702 (O_702,N_19994,N_19490);
xnor UO_703 (O_703,N_19994,N_19468);
nand UO_704 (O_704,N_19801,N_19824);
nor UO_705 (O_705,N_19232,N_19917);
or UO_706 (O_706,N_19425,N_19258);
xor UO_707 (O_707,N_19423,N_19865);
and UO_708 (O_708,N_19670,N_19837);
and UO_709 (O_709,N_19547,N_19745);
nand UO_710 (O_710,N_19344,N_19707);
nor UO_711 (O_711,N_19231,N_19357);
xnor UO_712 (O_712,N_19522,N_19703);
xor UO_713 (O_713,N_19310,N_19241);
or UO_714 (O_714,N_19815,N_19406);
and UO_715 (O_715,N_19627,N_19329);
and UO_716 (O_716,N_19747,N_19897);
nand UO_717 (O_717,N_19765,N_19266);
and UO_718 (O_718,N_19406,N_19739);
and UO_719 (O_719,N_19471,N_19212);
nor UO_720 (O_720,N_19975,N_19997);
nor UO_721 (O_721,N_19318,N_19961);
or UO_722 (O_722,N_19981,N_19283);
and UO_723 (O_723,N_19289,N_19781);
nand UO_724 (O_724,N_19701,N_19301);
or UO_725 (O_725,N_19829,N_19863);
nor UO_726 (O_726,N_19482,N_19462);
nor UO_727 (O_727,N_19394,N_19850);
and UO_728 (O_728,N_19418,N_19491);
nand UO_729 (O_729,N_19581,N_19246);
xor UO_730 (O_730,N_19360,N_19698);
nor UO_731 (O_731,N_19228,N_19482);
nor UO_732 (O_732,N_19778,N_19419);
nor UO_733 (O_733,N_19877,N_19712);
nand UO_734 (O_734,N_19664,N_19938);
nor UO_735 (O_735,N_19206,N_19308);
and UO_736 (O_736,N_19529,N_19221);
and UO_737 (O_737,N_19871,N_19466);
or UO_738 (O_738,N_19326,N_19638);
or UO_739 (O_739,N_19812,N_19481);
nand UO_740 (O_740,N_19770,N_19832);
and UO_741 (O_741,N_19475,N_19228);
nand UO_742 (O_742,N_19824,N_19285);
nand UO_743 (O_743,N_19701,N_19326);
or UO_744 (O_744,N_19500,N_19923);
xor UO_745 (O_745,N_19680,N_19616);
nor UO_746 (O_746,N_19691,N_19632);
or UO_747 (O_747,N_19635,N_19444);
xor UO_748 (O_748,N_19796,N_19797);
or UO_749 (O_749,N_19228,N_19783);
xnor UO_750 (O_750,N_19739,N_19330);
or UO_751 (O_751,N_19303,N_19804);
nor UO_752 (O_752,N_19796,N_19277);
nor UO_753 (O_753,N_19311,N_19485);
or UO_754 (O_754,N_19272,N_19297);
nor UO_755 (O_755,N_19408,N_19232);
xor UO_756 (O_756,N_19512,N_19876);
nor UO_757 (O_757,N_19597,N_19375);
and UO_758 (O_758,N_19900,N_19489);
or UO_759 (O_759,N_19840,N_19309);
or UO_760 (O_760,N_19598,N_19904);
nor UO_761 (O_761,N_19494,N_19757);
or UO_762 (O_762,N_19810,N_19583);
or UO_763 (O_763,N_19772,N_19367);
or UO_764 (O_764,N_19733,N_19880);
nand UO_765 (O_765,N_19314,N_19238);
or UO_766 (O_766,N_19631,N_19223);
xnor UO_767 (O_767,N_19922,N_19334);
nor UO_768 (O_768,N_19325,N_19443);
xnor UO_769 (O_769,N_19352,N_19627);
and UO_770 (O_770,N_19357,N_19385);
nor UO_771 (O_771,N_19406,N_19448);
nand UO_772 (O_772,N_19695,N_19448);
xnor UO_773 (O_773,N_19458,N_19804);
nand UO_774 (O_774,N_19686,N_19265);
xnor UO_775 (O_775,N_19691,N_19785);
nor UO_776 (O_776,N_19935,N_19726);
or UO_777 (O_777,N_19355,N_19868);
nor UO_778 (O_778,N_19342,N_19526);
nor UO_779 (O_779,N_19350,N_19375);
or UO_780 (O_780,N_19500,N_19665);
or UO_781 (O_781,N_19584,N_19239);
and UO_782 (O_782,N_19656,N_19678);
and UO_783 (O_783,N_19709,N_19905);
and UO_784 (O_784,N_19420,N_19747);
xor UO_785 (O_785,N_19848,N_19515);
or UO_786 (O_786,N_19316,N_19561);
nand UO_787 (O_787,N_19943,N_19344);
or UO_788 (O_788,N_19854,N_19229);
xor UO_789 (O_789,N_19289,N_19972);
nor UO_790 (O_790,N_19569,N_19583);
xor UO_791 (O_791,N_19984,N_19415);
or UO_792 (O_792,N_19747,N_19264);
and UO_793 (O_793,N_19507,N_19901);
or UO_794 (O_794,N_19906,N_19607);
xor UO_795 (O_795,N_19254,N_19262);
or UO_796 (O_796,N_19833,N_19700);
nand UO_797 (O_797,N_19737,N_19355);
or UO_798 (O_798,N_19378,N_19516);
or UO_799 (O_799,N_19786,N_19343);
xnor UO_800 (O_800,N_19496,N_19379);
and UO_801 (O_801,N_19358,N_19407);
or UO_802 (O_802,N_19517,N_19639);
nand UO_803 (O_803,N_19390,N_19919);
xor UO_804 (O_804,N_19715,N_19459);
or UO_805 (O_805,N_19704,N_19601);
nand UO_806 (O_806,N_19990,N_19398);
and UO_807 (O_807,N_19734,N_19249);
xnor UO_808 (O_808,N_19209,N_19916);
or UO_809 (O_809,N_19993,N_19390);
or UO_810 (O_810,N_19300,N_19601);
nor UO_811 (O_811,N_19902,N_19415);
or UO_812 (O_812,N_19283,N_19655);
and UO_813 (O_813,N_19975,N_19537);
nand UO_814 (O_814,N_19498,N_19994);
xnor UO_815 (O_815,N_19440,N_19847);
xor UO_816 (O_816,N_19512,N_19511);
and UO_817 (O_817,N_19902,N_19242);
or UO_818 (O_818,N_19814,N_19965);
nand UO_819 (O_819,N_19989,N_19710);
nor UO_820 (O_820,N_19634,N_19512);
or UO_821 (O_821,N_19259,N_19477);
and UO_822 (O_822,N_19431,N_19285);
and UO_823 (O_823,N_19405,N_19813);
xor UO_824 (O_824,N_19992,N_19738);
xnor UO_825 (O_825,N_19822,N_19626);
or UO_826 (O_826,N_19597,N_19747);
nor UO_827 (O_827,N_19278,N_19783);
nand UO_828 (O_828,N_19523,N_19640);
nor UO_829 (O_829,N_19637,N_19235);
or UO_830 (O_830,N_19629,N_19856);
xnor UO_831 (O_831,N_19776,N_19762);
nor UO_832 (O_832,N_19595,N_19266);
nor UO_833 (O_833,N_19521,N_19629);
or UO_834 (O_834,N_19544,N_19985);
nor UO_835 (O_835,N_19275,N_19356);
and UO_836 (O_836,N_19398,N_19819);
or UO_837 (O_837,N_19770,N_19760);
nor UO_838 (O_838,N_19796,N_19643);
or UO_839 (O_839,N_19327,N_19237);
and UO_840 (O_840,N_19749,N_19287);
and UO_841 (O_841,N_19865,N_19411);
or UO_842 (O_842,N_19443,N_19535);
xnor UO_843 (O_843,N_19796,N_19672);
xor UO_844 (O_844,N_19255,N_19244);
nand UO_845 (O_845,N_19608,N_19693);
nand UO_846 (O_846,N_19802,N_19975);
or UO_847 (O_847,N_19879,N_19224);
nor UO_848 (O_848,N_19773,N_19504);
nor UO_849 (O_849,N_19908,N_19628);
nand UO_850 (O_850,N_19241,N_19513);
and UO_851 (O_851,N_19753,N_19671);
or UO_852 (O_852,N_19243,N_19755);
nor UO_853 (O_853,N_19818,N_19986);
or UO_854 (O_854,N_19745,N_19913);
or UO_855 (O_855,N_19761,N_19221);
nor UO_856 (O_856,N_19254,N_19911);
or UO_857 (O_857,N_19487,N_19236);
and UO_858 (O_858,N_19286,N_19233);
and UO_859 (O_859,N_19969,N_19548);
nand UO_860 (O_860,N_19708,N_19583);
and UO_861 (O_861,N_19489,N_19337);
or UO_862 (O_862,N_19404,N_19721);
or UO_863 (O_863,N_19728,N_19922);
nand UO_864 (O_864,N_19500,N_19280);
or UO_865 (O_865,N_19837,N_19869);
or UO_866 (O_866,N_19562,N_19725);
nor UO_867 (O_867,N_19963,N_19544);
nand UO_868 (O_868,N_19698,N_19458);
and UO_869 (O_869,N_19844,N_19532);
nand UO_870 (O_870,N_19705,N_19974);
and UO_871 (O_871,N_19421,N_19962);
and UO_872 (O_872,N_19257,N_19424);
xnor UO_873 (O_873,N_19635,N_19996);
nor UO_874 (O_874,N_19447,N_19500);
nand UO_875 (O_875,N_19253,N_19952);
nor UO_876 (O_876,N_19733,N_19210);
xnor UO_877 (O_877,N_19329,N_19217);
and UO_878 (O_878,N_19333,N_19909);
and UO_879 (O_879,N_19547,N_19699);
nor UO_880 (O_880,N_19316,N_19770);
nor UO_881 (O_881,N_19272,N_19325);
nand UO_882 (O_882,N_19243,N_19380);
nor UO_883 (O_883,N_19328,N_19890);
nand UO_884 (O_884,N_19834,N_19708);
and UO_885 (O_885,N_19563,N_19223);
nor UO_886 (O_886,N_19381,N_19538);
xor UO_887 (O_887,N_19209,N_19930);
and UO_888 (O_888,N_19412,N_19935);
xor UO_889 (O_889,N_19905,N_19379);
and UO_890 (O_890,N_19832,N_19394);
nor UO_891 (O_891,N_19797,N_19946);
nor UO_892 (O_892,N_19809,N_19570);
nor UO_893 (O_893,N_19925,N_19424);
nand UO_894 (O_894,N_19385,N_19770);
nor UO_895 (O_895,N_19708,N_19681);
nand UO_896 (O_896,N_19917,N_19898);
or UO_897 (O_897,N_19980,N_19716);
nor UO_898 (O_898,N_19694,N_19491);
and UO_899 (O_899,N_19470,N_19887);
nand UO_900 (O_900,N_19460,N_19917);
xnor UO_901 (O_901,N_19704,N_19616);
xor UO_902 (O_902,N_19219,N_19477);
or UO_903 (O_903,N_19755,N_19479);
or UO_904 (O_904,N_19885,N_19612);
nand UO_905 (O_905,N_19514,N_19329);
or UO_906 (O_906,N_19806,N_19375);
nor UO_907 (O_907,N_19777,N_19202);
nor UO_908 (O_908,N_19943,N_19788);
and UO_909 (O_909,N_19616,N_19274);
nor UO_910 (O_910,N_19506,N_19629);
or UO_911 (O_911,N_19801,N_19435);
nor UO_912 (O_912,N_19622,N_19389);
nor UO_913 (O_913,N_19780,N_19935);
nor UO_914 (O_914,N_19842,N_19266);
or UO_915 (O_915,N_19811,N_19968);
nand UO_916 (O_916,N_19256,N_19253);
and UO_917 (O_917,N_19846,N_19400);
nor UO_918 (O_918,N_19924,N_19858);
and UO_919 (O_919,N_19648,N_19569);
and UO_920 (O_920,N_19604,N_19379);
nand UO_921 (O_921,N_19379,N_19329);
nor UO_922 (O_922,N_19705,N_19437);
nand UO_923 (O_923,N_19959,N_19319);
or UO_924 (O_924,N_19653,N_19708);
xnor UO_925 (O_925,N_19465,N_19446);
and UO_926 (O_926,N_19589,N_19740);
nand UO_927 (O_927,N_19930,N_19434);
or UO_928 (O_928,N_19943,N_19368);
nand UO_929 (O_929,N_19776,N_19828);
nor UO_930 (O_930,N_19273,N_19533);
nand UO_931 (O_931,N_19897,N_19693);
nor UO_932 (O_932,N_19681,N_19395);
or UO_933 (O_933,N_19940,N_19481);
or UO_934 (O_934,N_19788,N_19926);
or UO_935 (O_935,N_19679,N_19282);
and UO_936 (O_936,N_19348,N_19637);
nand UO_937 (O_937,N_19341,N_19316);
nor UO_938 (O_938,N_19408,N_19722);
nand UO_939 (O_939,N_19645,N_19842);
and UO_940 (O_940,N_19271,N_19467);
and UO_941 (O_941,N_19331,N_19382);
or UO_942 (O_942,N_19539,N_19979);
nor UO_943 (O_943,N_19839,N_19840);
xor UO_944 (O_944,N_19700,N_19310);
xor UO_945 (O_945,N_19613,N_19865);
nand UO_946 (O_946,N_19448,N_19831);
xnor UO_947 (O_947,N_19484,N_19863);
or UO_948 (O_948,N_19350,N_19464);
xnor UO_949 (O_949,N_19669,N_19494);
nor UO_950 (O_950,N_19422,N_19917);
nand UO_951 (O_951,N_19756,N_19439);
or UO_952 (O_952,N_19522,N_19736);
or UO_953 (O_953,N_19796,N_19379);
or UO_954 (O_954,N_19954,N_19355);
or UO_955 (O_955,N_19437,N_19571);
nand UO_956 (O_956,N_19945,N_19997);
and UO_957 (O_957,N_19326,N_19954);
xnor UO_958 (O_958,N_19957,N_19515);
nand UO_959 (O_959,N_19487,N_19286);
or UO_960 (O_960,N_19741,N_19488);
xnor UO_961 (O_961,N_19340,N_19351);
xor UO_962 (O_962,N_19462,N_19467);
nand UO_963 (O_963,N_19434,N_19473);
xnor UO_964 (O_964,N_19611,N_19240);
xor UO_965 (O_965,N_19309,N_19980);
nand UO_966 (O_966,N_19660,N_19266);
xnor UO_967 (O_967,N_19463,N_19836);
or UO_968 (O_968,N_19669,N_19702);
or UO_969 (O_969,N_19890,N_19568);
xor UO_970 (O_970,N_19360,N_19439);
and UO_971 (O_971,N_19742,N_19754);
or UO_972 (O_972,N_19598,N_19783);
xnor UO_973 (O_973,N_19663,N_19814);
or UO_974 (O_974,N_19584,N_19767);
xnor UO_975 (O_975,N_19521,N_19915);
nor UO_976 (O_976,N_19855,N_19984);
nor UO_977 (O_977,N_19759,N_19816);
nor UO_978 (O_978,N_19455,N_19250);
and UO_979 (O_979,N_19467,N_19269);
or UO_980 (O_980,N_19611,N_19524);
nand UO_981 (O_981,N_19443,N_19237);
nor UO_982 (O_982,N_19785,N_19284);
nand UO_983 (O_983,N_19752,N_19273);
xor UO_984 (O_984,N_19351,N_19941);
or UO_985 (O_985,N_19209,N_19612);
and UO_986 (O_986,N_19983,N_19937);
nand UO_987 (O_987,N_19830,N_19979);
nor UO_988 (O_988,N_19486,N_19862);
and UO_989 (O_989,N_19886,N_19895);
nor UO_990 (O_990,N_19320,N_19941);
or UO_991 (O_991,N_19785,N_19432);
and UO_992 (O_992,N_19253,N_19608);
and UO_993 (O_993,N_19686,N_19696);
or UO_994 (O_994,N_19680,N_19395);
or UO_995 (O_995,N_19320,N_19259);
xnor UO_996 (O_996,N_19579,N_19824);
nand UO_997 (O_997,N_19793,N_19868);
and UO_998 (O_998,N_19971,N_19252);
or UO_999 (O_999,N_19495,N_19973);
and UO_1000 (O_1000,N_19466,N_19916);
and UO_1001 (O_1001,N_19944,N_19435);
nor UO_1002 (O_1002,N_19245,N_19623);
nand UO_1003 (O_1003,N_19930,N_19589);
and UO_1004 (O_1004,N_19534,N_19370);
nor UO_1005 (O_1005,N_19980,N_19303);
xnor UO_1006 (O_1006,N_19525,N_19665);
or UO_1007 (O_1007,N_19914,N_19411);
and UO_1008 (O_1008,N_19659,N_19310);
and UO_1009 (O_1009,N_19246,N_19281);
xnor UO_1010 (O_1010,N_19302,N_19563);
nand UO_1011 (O_1011,N_19931,N_19671);
nor UO_1012 (O_1012,N_19996,N_19966);
and UO_1013 (O_1013,N_19813,N_19284);
nand UO_1014 (O_1014,N_19448,N_19374);
or UO_1015 (O_1015,N_19904,N_19885);
or UO_1016 (O_1016,N_19852,N_19967);
xor UO_1017 (O_1017,N_19274,N_19843);
xnor UO_1018 (O_1018,N_19803,N_19775);
nor UO_1019 (O_1019,N_19468,N_19975);
nor UO_1020 (O_1020,N_19873,N_19644);
or UO_1021 (O_1021,N_19479,N_19785);
nor UO_1022 (O_1022,N_19902,N_19565);
xor UO_1023 (O_1023,N_19661,N_19894);
nor UO_1024 (O_1024,N_19773,N_19343);
or UO_1025 (O_1025,N_19723,N_19227);
nand UO_1026 (O_1026,N_19673,N_19993);
xor UO_1027 (O_1027,N_19490,N_19281);
nor UO_1028 (O_1028,N_19767,N_19659);
or UO_1029 (O_1029,N_19934,N_19486);
nand UO_1030 (O_1030,N_19711,N_19949);
nor UO_1031 (O_1031,N_19568,N_19259);
or UO_1032 (O_1032,N_19319,N_19701);
nor UO_1033 (O_1033,N_19384,N_19377);
nor UO_1034 (O_1034,N_19950,N_19583);
nand UO_1035 (O_1035,N_19696,N_19576);
nand UO_1036 (O_1036,N_19921,N_19693);
nand UO_1037 (O_1037,N_19265,N_19647);
xnor UO_1038 (O_1038,N_19529,N_19767);
nand UO_1039 (O_1039,N_19317,N_19327);
nor UO_1040 (O_1040,N_19574,N_19478);
and UO_1041 (O_1041,N_19498,N_19553);
or UO_1042 (O_1042,N_19540,N_19979);
or UO_1043 (O_1043,N_19640,N_19379);
and UO_1044 (O_1044,N_19752,N_19532);
nor UO_1045 (O_1045,N_19716,N_19278);
or UO_1046 (O_1046,N_19656,N_19341);
xnor UO_1047 (O_1047,N_19284,N_19348);
nand UO_1048 (O_1048,N_19905,N_19443);
and UO_1049 (O_1049,N_19864,N_19359);
nor UO_1050 (O_1050,N_19392,N_19408);
xnor UO_1051 (O_1051,N_19594,N_19248);
or UO_1052 (O_1052,N_19403,N_19245);
and UO_1053 (O_1053,N_19533,N_19971);
nor UO_1054 (O_1054,N_19645,N_19843);
or UO_1055 (O_1055,N_19298,N_19685);
and UO_1056 (O_1056,N_19387,N_19430);
and UO_1057 (O_1057,N_19304,N_19363);
or UO_1058 (O_1058,N_19613,N_19546);
xor UO_1059 (O_1059,N_19697,N_19534);
and UO_1060 (O_1060,N_19746,N_19988);
nand UO_1061 (O_1061,N_19370,N_19242);
and UO_1062 (O_1062,N_19506,N_19741);
xnor UO_1063 (O_1063,N_19746,N_19415);
xnor UO_1064 (O_1064,N_19738,N_19317);
and UO_1065 (O_1065,N_19674,N_19972);
or UO_1066 (O_1066,N_19326,N_19916);
or UO_1067 (O_1067,N_19328,N_19338);
nor UO_1068 (O_1068,N_19586,N_19823);
nand UO_1069 (O_1069,N_19646,N_19665);
or UO_1070 (O_1070,N_19968,N_19594);
xor UO_1071 (O_1071,N_19660,N_19875);
xnor UO_1072 (O_1072,N_19300,N_19703);
xnor UO_1073 (O_1073,N_19367,N_19373);
and UO_1074 (O_1074,N_19588,N_19214);
nand UO_1075 (O_1075,N_19839,N_19718);
nand UO_1076 (O_1076,N_19436,N_19542);
or UO_1077 (O_1077,N_19797,N_19754);
or UO_1078 (O_1078,N_19497,N_19209);
xnor UO_1079 (O_1079,N_19242,N_19860);
and UO_1080 (O_1080,N_19826,N_19488);
nand UO_1081 (O_1081,N_19957,N_19345);
xnor UO_1082 (O_1082,N_19534,N_19404);
and UO_1083 (O_1083,N_19515,N_19815);
or UO_1084 (O_1084,N_19480,N_19488);
nand UO_1085 (O_1085,N_19517,N_19802);
or UO_1086 (O_1086,N_19645,N_19568);
xor UO_1087 (O_1087,N_19973,N_19999);
and UO_1088 (O_1088,N_19548,N_19350);
nor UO_1089 (O_1089,N_19873,N_19512);
and UO_1090 (O_1090,N_19637,N_19816);
nor UO_1091 (O_1091,N_19923,N_19662);
nor UO_1092 (O_1092,N_19277,N_19496);
nand UO_1093 (O_1093,N_19390,N_19222);
or UO_1094 (O_1094,N_19380,N_19736);
xnor UO_1095 (O_1095,N_19428,N_19386);
or UO_1096 (O_1096,N_19820,N_19477);
and UO_1097 (O_1097,N_19239,N_19675);
nand UO_1098 (O_1098,N_19269,N_19891);
nor UO_1099 (O_1099,N_19269,N_19667);
or UO_1100 (O_1100,N_19606,N_19240);
or UO_1101 (O_1101,N_19834,N_19553);
and UO_1102 (O_1102,N_19748,N_19406);
and UO_1103 (O_1103,N_19384,N_19798);
and UO_1104 (O_1104,N_19867,N_19395);
xor UO_1105 (O_1105,N_19396,N_19980);
xor UO_1106 (O_1106,N_19982,N_19887);
xnor UO_1107 (O_1107,N_19896,N_19347);
nand UO_1108 (O_1108,N_19456,N_19773);
nand UO_1109 (O_1109,N_19207,N_19781);
and UO_1110 (O_1110,N_19482,N_19790);
nor UO_1111 (O_1111,N_19350,N_19962);
xor UO_1112 (O_1112,N_19803,N_19271);
xor UO_1113 (O_1113,N_19255,N_19258);
nor UO_1114 (O_1114,N_19942,N_19986);
nor UO_1115 (O_1115,N_19391,N_19606);
or UO_1116 (O_1116,N_19894,N_19657);
nor UO_1117 (O_1117,N_19370,N_19720);
and UO_1118 (O_1118,N_19747,N_19815);
xnor UO_1119 (O_1119,N_19679,N_19366);
and UO_1120 (O_1120,N_19200,N_19558);
nor UO_1121 (O_1121,N_19398,N_19939);
nand UO_1122 (O_1122,N_19278,N_19370);
nand UO_1123 (O_1123,N_19906,N_19699);
nor UO_1124 (O_1124,N_19413,N_19387);
and UO_1125 (O_1125,N_19988,N_19310);
xor UO_1126 (O_1126,N_19500,N_19822);
and UO_1127 (O_1127,N_19316,N_19844);
nor UO_1128 (O_1128,N_19559,N_19564);
and UO_1129 (O_1129,N_19685,N_19567);
xor UO_1130 (O_1130,N_19865,N_19875);
nor UO_1131 (O_1131,N_19424,N_19394);
nand UO_1132 (O_1132,N_19675,N_19727);
nor UO_1133 (O_1133,N_19871,N_19429);
nor UO_1134 (O_1134,N_19464,N_19358);
or UO_1135 (O_1135,N_19705,N_19827);
or UO_1136 (O_1136,N_19457,N_19410);
nand UO_1137 (O_1137,N_19716,N_19411);
xor UO_1138 (O_1138,N_19227,N_19779);
nand UO_1139 (O_1139,N_19659,N_19209);
xor UO_1140 (O_1140,N_19472,N_19985);
or UO_1141 (O_1141,N_19314,N_19970);
or UO_1142 (O_1142,N_19249,N_19925);
nor UO_1143 (O_1143,N_19661,N_19915);
xnor UO_1144 (O_1144,N_19683,N_19294);
and UO_1145 (O_1145,N_19986,N_19278);
and UO_1146 (O_1146,N_19539,N_19424);
xor UO_1147 (O_1147,N_19513,N_19603);
nor UO_1148 (O_1148,N_19250,N_19482);
nor UO_1149 (O_1149,N_19270,N_19451);
nor UO_1150 (O_1150,N_19477,N_19391);
xnor UO_1151 (O_1151,N_19625,N_19879);
xor UO_1152 (O_1152,N_19342,N_19710);
nor UO_1153 (O_1153,N_19554,N_19507);
xnor UO_1154 (O_1154,N_19601,N_19483);
nor UO_1155 (O_1155,N_19987,N_19865);
xor UO_1156 (O_1156,N_19970,N_19992);
or UO_1157 (O_1157,N_19971,N_19841);
or UO_1158 (O_1158,N_19865,N_19370);
or UO_1159 (O_1159,N_19597,N_19552);
and UO_1160 (O_1160,N_19822,N_19480);
or UO_1161 (O_1161,N_19635,N_19946);
nor UO_1162 (O_1162,N_19779,N_19899);
and UO_1163 (O_1163,N_19603,N_19759);
and UO_1164 (O_1164,N_19862,N_19238);
nor UO_1165 (O_1165,N_19877,N_19790);
nor UO_1166 (O_1166,N_19337,N_19594);
nor UO_1167 (O_1167,N_19813,N_19678);
or UO_1168 (O_1168,N_19438,N_19678);
or UO_1169 (O_1169,N_19662,N_19392);
or UO_1170 (O_1170,N_19430,N_19291);
nand UO_1171 (O_1171,N_19754,N_19355);
nand UO_1172 (O_1172,N_19923,N_19628);
nor UO_1173 (O_1173,N_19736,N_19356);
nand UO_1174 (O_1174,N_19595,N_19558);
nor UO_1175 (O_1175,N_19708,N_19275);
nand UO_1176 (O_1176,N_19788,N_19866);
xor UO_1177 (O_1177,N_19967,N_19460);
or UO_1178 (O_1178,N_19608,N_19746);
nand UO_1179 (O_1179,N_19459,N_19446);
xor UO_1180 (O_1180,N_19896,N_19403);
xor UO_1181 (O_1181,N_19474,N_19471);
nand UO_1182 (O_1182,N_19429,N_19519);
xor UO_1183 (O_1183,N_19571,N_19559);
or UO_1184 (O_1184,N_19817,N_19998);
xor UO_1185 (O_1185,N_19463,N_19963);
xor UO_1186 (O_1186,N_19763,N_19244);
or UO_1187 (O_1187,N_19447,N_19282);
nor UO_1188 (O_1188,N_19505,N_19334);
nor UO_1189 (O_1189,N_19905,N_19635);
nor UO_1190 (O_1190,N_19515,N_19320);
nor UO_1191 (O_1191,N_19241,N_19837);
and UO_1192 (O_1192,N_19506,N_19348);
nor UO_1193 (O_1193,N_19778,N_19635);
nand UO_1194 (O_1194,N_19569,N_19220);
nand UO_1195 (O_1195,N_19808,N_19752);
xnor UO_1196 (O_1196,N_19309,N_19353);
and UO_1197 (O_1197,N_19913,N_19628);
or UO_1198 (O_1198,N_19663,N_19329);
nor UO_1199 (O_1199,N_19539,N_19490);
nand UO_1200 (O_1200,N_19305,N_19423);
xnor UO_1201 (O_1201,N_19854,N_19358);
or UO_1202 (O_1202,N_19722,N_19427);
xnor UO_1203 (O_1203,N_19691,N_19419);
or UO_1204 (O_1204,N_19982,N_19267);
xor UO_1205 (O_1205,N_19960,N_19780);
nand UO_1206 (O_1206,N_19574,N_19225);
or UO_1207 (O_1207,N_19988,N_19286);
nand UO_1208 (O_1208,N_19581,N_19890);
xnor UO_1209 (O_1209,N_19612,N_19985);
nor UO_1210 (O_1210,N_19786,N_19812);
and UO_1211 (O_1211,N_19991,N_19474);
nor UO_1212 (O_1212,N_19621,N_19958);
nor UO_1213 (O_1213,N_19358,N_19452);
or UO_1214 (O_1214,N_19651,N_19431);
nand UO_1215 (O_1215,N_19428,N_19213);
xnor UO_1216 (O_1216,N_19221,N_19359);
nor UO_1217 (O_1217,N_19666,N_19755);
nor UO_1218 (O_1218,N_19538,N_19262);
nand UO_1219 (O_1219,N_19632,N_19321);
nor UO_1220 (O_1220,N_19209,N_19261);
or UO_1221 (O_1221,N_19399,N_19322);
nor UO_1222 (O_1222,N_19384,N_19300);
or UO_1223 (O_1223,N_19585,N_19893);
nand UO_1224 (O_1224,N_19396,N_19327);
nor UO_1225 (O_1225,N_19273,N_19907);
nor UO_1226 (O_1226,N_19589,N_19756);
xnor UO_1227 (O_1227,N_19248,N_19324);
and UO_1228 (O_1228,N_19997,N_19244);
or UO_1229 (O_1229,N_19650,N_19402);
nand UO_1230 (O_1230,N_19292,N_19206);
nand UO_1231 (O_1231,N_19385,N_19230);
nor UO_1232 (O_1232,N_19602,N_19488);
nor UO_1233 (O_1233,N_19514,N_19340);
and UO_1234 (O_1234,N_19219,N_19409);
nor UO_1235 (O_1235,N_19822,N_19631);
nor UO_1236 (O_1236,N_19716,N_19632);
nand UO_1237 (O_1237,N_19678,N_19411);
or UO_1238 (O_1238,N_19204,N_19429);
xnor UO_1239 (O_1239,N_19398,N_19700);
nor UO_1240 (O_1240,N_19571,N_19325);
and UO_1241 (O_1241,N_19459,N_19283);
and UO_1242 (O_1242,N_19754,N_19421);
nand UO_1243 (O_1243,N_19383,N_19969);
and UO_1244 (O_1244,N_19660,N_19256);
nor UO_1245 (O_1245,N_19592,N_19524);
and UO_1246 (O_1246,N_19869,N_19918);
nor UO_1247 (O_1247,N_19625,N_19322);
xor UO_1248 (O_1248,N_19785,N_19402);
nand UO_1249 (O_1249,N_19816,N_19652);
or UO_1250 (O_1250,N_19946,N_19683);
or UO_1251 (O_1251,N_19696,N_19617);
nor UO_1252 (O_1252,N_19272,N_19289);
xor UO_1253 (O_1253,N_19814,N_19309);
xnor UO_1254 (O_1254,N_19884,N_19992);
or UO_1255 (O_1255,N_19864,N_19896);
and UO_1256 (O_1256,N_19615,N_19689);
nand UO_1257 (O_1257,N_19739,N_19667);
or UO_1258 (O_1258,N_19234,N_19403);
nand UO_1259 (O_1259,N_19222,N_19755);
or UO_1260 (O_1260,N_19912,N_19496);
or UO_1261 (O_1261,N_19880,N_19925);
or UO_1262 (O_1262,N_19375,N_19381);
or UO_1263 (O_1263,N_19230,N_19898);
nor UO_1264 (O_1264,N_19600,N_19546);
nand UO_1265 (O_1265,N_19657,N_19206);
nor UO_1266 (O_1266,N_19249,N_19686);
nor UO_1267 (O_1267,N_19489,N_19948);
and UO_1268 (O_1268,N_19251,N_19507);
nor UO_1269 (O_1269,N_19624,N_19738);
nand UO_1270 (O_1270,N_19562,N_19333);
or UO_1271 (O_1271,N_19719,N_19473);
and UO_1272 (O_1272,N_19939,N_19497);
xor UO_1273 (O_1273,N_19827,N_19332);
nand UO_1274 (O_1274,N_19956,N_19491);
and UO_1275 (O_1275,N_19401,N_19678);
nor UO_1276 (O_1276,N_19500,N_19320);
nand UO_1277 (O_1277,N_19279,N_19900);
xnor UO_1278 (O_1278,N_19581,N_19499);
nand UO_1279 (O_1279,N_19827,N_19321);
or UO_1280 (O_1280,N_19680,N_19261);
and UO_1281 (O_1281,N_19644,N_19865);
and UO_1282 (O_1282,N_19577,N_19312);
and UO_1283 (O_1283,N_19288,N_19397);
nor UO_1284 (O_1284,N_19786,N_19289);
and UO_1285 (O_1285,N_19661,N_19920);
nor UO_1286 (O_1286,N_19768,N_19354);
and UO_1287 (O_1287,N_19783,N_19737);
and UO_1288 (O_1288,N_19503,N_19660);
or UO_1289 (O_1289,N_19634,N_19621);
xnor UO_1290 (O_1290,N_19850,N_19748);
nor UO_1291 (O_1291,N_19897,N_19209);
nor UO_1292 (O_1292,N_19463,N_19597);
nor UO_1293 (O_1293,N_19203,N_19250);
or UO_1294 (O_1294,N_19452,N_19602);
or UO_1295 (O_1295,N_19944,N_19444);
nor UO_1296 (O_1296,N_19914,N_19702);
or UO_1297 (O_1297,N_19253,N_19661);
nand UO_1298 (O_1298,N_19333,N_19764);
nand UO_1299 (O_1299,N_19516,N_19451);
or UO_1300 (O_1300,N_19906,N_19677);
nand UO_1301 (O_1301,N_19720,N_19362);
and UO_1302 (O_1302,N_19873,N_19563);
xor UO_1303 (O_1303,N_19519,N_19974);
and UO_1304 (O_1304,N_19450,N_19241);
and UO_1305 (O_1305,N_19289,N_19573);
and UO_1306 (O_1306,N_19239,N_19472);
nor UO_1307 (O_1307,N_19206,N_19866);
or UO_1308 (O_1308,N_19625,N_19536);
xor UO_1309 (O_1309,N_19893,N_19239);
or UO_1310 (O_1310,N_19906,N_19739);
nand UO_1311 (O_1311,N_19270,N_19366);
xor UO_1312 (O_1312,N_19315,N_19461);
or UO_1313 (O_1313,N_19247,N_19580);
xor UO_1314 (O_1314,N_19547,N_19219);
and UO_1315 (O_1315,N_19681,N_19397);
and UO_1316 (O_1316,N_19978,N_19804);
xnor UO_1317 (O_1317,N_19937,N_19408);
or UO_1318 (O_1318,N_19717,N_19248);
nor UO_1319 (O_1319,N_19249,N_19421);
and UO_1320 (O_1320,N_19686,N_19253);
xor UO_1321 (O_1321,N_19424,N_19728);
and UO_1322 (O_1322,N_19551,N_19577);
nand UO_1323 (O_1323,N_19492,N_19722);
or UO_1324 (O_1324,N_19466,N_19858);
xnor UO_1325 (O_1325,N_19699,N_19538);
and UO_1326 (O_1326,N_19939,N_19539);
xnor UO_1327 (O_1327,N_19444,N_19287);
or UO_1328 (O_1328,N_19214,N_19918);
and UO_1329 (O_1329,N_19933,N_19773);
xor UO_1330 (O_1330,N_19675,N_19939);
or UO_1331 (O_1331,N_19483,N_19500);
nor UO_1332 (O_1332,N_19278,N_19740);
nor UO_1333 (O_1333,N_19509,N_19354);
xnor UO_1334 (O_1334,N_19264,N_19518);
nor UO_1335 (O_1335,N_19445,N_19764);
nor UO_1336 (O_1336,N_19585,N_19517);
nand UO_1337 (O_1337,N_19769,N_19972);
or UO_1338 (O_1338,N_19495,N_19913);
or UO_1339 (O_1339,N_19817,N_19215);
nor UO_1340 (O_1340,N_19303,N_19708);
xnor UO_1341 (O_1341,N_19762,N_19493);
or UO_1342 (O_1342,N_19733,N_19272);
nand UO_1343 (O_1343,N_19962,N_19974);
xor UO_1344 (O_1344,N_19369,N_19690);
and UO_1345 (O_1345,N_19235,N_19478);
xnor UO_1346 (O_1346,N_19556,N_19248);
and UO_1347 (O_1347,N_19573,N_19221);
nor UO_1348 (O_1348,N_19950,N_19851);
and UO_1349 (O_1349,N_19764,N_19227);
nand UO_1350 (O_1350,N_19516,N_19906);
or UO_1351 (O_1351,N_19571,N_19231);
xnor UO_1352 (O_1352,N_19670,N_19955);
nor UO_1353 (O_1353,N_19230,N_19384);
or UO_1354 (O_1354,N_19856,N_19348);
xor UO_1355 (O_1355,N_19343,N_19715);
and UO_1356 (O_1356,N_19925,N_19826);
or UO_1357 (O_1357,N_19917,N_19317);
xor UO_1358 (O_1358,N_19717,N_19381);
or UO_1359 (O_1359,N_19592,N_19414);
or UO_1360 (O_1360,N_19266,N_19324);
xnor UO_1361 (O_1361,N_19264,N_19539);
nand UO_1362 (O_1362,N_19851,N_19594);
xor UO_1363 (O_1363,N_19306,N_19229);
nor UO_1364 (O_1364,N_19370,N_19206);
or UO_1365 (O_1365,N_19992,N_19391);
nand UO_1366 (O_1366,N_19773,N_19693);
nor UO_1367 (O_1367,N_19260,N_19270);
xnor UO_1368 (O_1368,N_19863,N_19792);
nand UO_1369 (O_1369,N_19419,N_19420);
and UO_1370 (O_1370,N_19921,N_19223);
or UO_1371 (O_1371,N_19437,N_19271);
nand UO_1372 (O_1372,N_19758,N_19866);
and UO_1373 (O_1373,N_19232,N_19524);
nor UO_1374 (O_1374,N_19999,N_19315);
nand UO_1375 (O_1375,N_19420,N_19650);
nand UO_1376 (O_1376,N_19707,N_19892);
nand UO_1377 (O_1377,N_19999,N_19432);
nand UO_1378 (O_1378,N_19636,N_19891);
or UO_1379 (O_1379,N_19248,N_19864);
and UO_1380 (O_1380,N_19961,N_19244);
nor UO_1381 (O_1381,N_19240,N_19631);
and UO_1382 (O_1382,N_19974,N_19919);
and UO_1383 (O_1383,N_19425,N_19585);
xor UO_1384 (O_1384,N_19708,N_19959);
xor UO_1385 (O_1385,N_19997,N_19389);
nor UO_1386 (O_1386,N_19627,N_19865);
nor UO_1387 (O_1387,N_19345,N_19390);
nand UO_1388 (O_1388,N_19996,N_19865);
or UO_1389 (O_1389,N_19520,N_19843);
or UO_1390 (O_1390,N_19581,N_19655);
and UO_1391 (O_1391,N_19626,N_19486);
xnor UO_1392 (O_1392,N_19400,N_19517);
nand UO_1393 (O_1393,N_19978,N_19524);
and UO_1394 (O_1394,N_19736,N_19899);
or UO_1395 (O_1395,N_19943,N_19453);
nand UO_1396 (O_1396,N_19302,N_19834);
nand UO_1397 (O_1397,N_19951,N_19852);
nand UO_1398 (O_1398,N_19585,N_19486);
and UO_1399 (O_1399,N_19943,N_19524);
xor UO_1400 (O_1400,N_19856,N_19882);
nand UO_1401 (O_1401,N_19571,N_19679);
and UO_1402 (O_1402,N_19267,N_19415);
nor UO_1403 (O_1403,N_19966,N_19921);
and UO_1404 (O_1404,N_19319,N_19914);
xor UO_1405 (O_1405,N_19303,N_19946);
nand UO_1406 (O_1406,N_19880,N_19260);
nand UO_1407 (O_1407,N_19771,N_19382);
nand UO_1408 (O_1408,N_19567,N_19565);
nor UO_1409 (O_1409,N_19841,N_19995);
or UO_1410 (O_1410,N_19603,N_19870);
nor UO_1411 (O_1411,N_19279,N_19253);
nand UO_1412 (O_1412,N_19515,N_19723);
nor UO_1413 (O_1413,N_19696,N_19317);
or UO_1414 (O_1414,N_19515,N_19849);
and UO_1415 (O_1415,N_19526,N_19865);
nor UO_1416 (O_1416,N_19751,N_19440);
or UO_1417 (O_1417,N_19915,N_19528);
or UO_1418 (O_1418,N_19810,N_19361);
xnor UO_1419 (O_1419,N_19841,N_19242);
and UO_1420 (O_1420,N_19211,N_19594);
nor UO_1421 (O_1421,N_19219,N_19930);
and UO_1422 (O_1422,N_19821,N_19803);
nand UO_1423 (O_1423,N_19565,N_19758);
or UO_1424 (O_1424,N_19781,N_19261);
nor UO_1425 (O_1425,N_19317,N_19277);
nor UO_1426 (O_1426,N_19273,N_19784);
or UO_1427 (O_1427,N_19546,N_19881);
xnor UO_1428 (O_1428,N_19884,N_19983);
nand UO_1429 (O_1429,N_19758,N_19201);
nand UO_1430 (O_1430,N_19889,N_19382);
nand UO_1431 (O_1431,N_19306,N_19986);
xor UO_1432 (O_1432,N_19302,N_19851);
nand UO_1433 (O_1433,N_19489,N_19665);
nor UO_1434 (O_1434,N_19425,N_19798);
and UO_1435 (O_1435,N_19766,N_19823);
nand UO_1436 (O_1436,N_19296,N_19688);
nor UO_1437 (O_1437,N_19275,N_19703);
and UO_1438 (O_1438,N_19755,N_19487);
nor UO_1439 (O_1439,N_19753,N_19660);
or UO_1440 (O_1440,N_19910,N_19432);
or UO_1441 (O_1441,N_19256,N_19291);
nor UO_1442 (O_1442,N_19462,N_19776);
or UO_1443 (O_1443,N_19363,N_19206);
and UO_1444 (O_1444,N_19335,N_19451);
or UO_1445 (O_1445,N_19291,N_19601);
nand UO_1446 (O_1446,N_19891,N_19525);
nand UO_1447 (O_1447,N_19655,N_19373);
nand UO_1448 (O_1448,N_19552,N_19452);
nand UO_1449 (O_1449,N_19512,N_19212);
xor UO_1450 (O_1450,N_19262,N_19665);
xor UO_1451 (O_1451,N_19835,N_19482);
or UO_1452 (O_1452,N_19762,N_19856);
and UO_1453 (O_1453,N_19583,N_19926);
nor UO_1454 (O_1454,N_19209,N_19392);
and UO_1455 (O_1455,N_19717,N_19695);
and UO_1456 (O_1456,N_19865,N_19943);
nand UO_1457 (O_1457,N_19212,N_19729);
xor UO_1458 (O_1458,N_19804,N_19721);
and UO_1459 (O_1459,N_19651,N_19313);
nor UO_1460 (O_1460,N_19835,N_19508);
xnor UO_1461 (O_1461,N_19575,N_19743);
nand UO_1462 (O_1462,N_19752,N_19236);
nor UO_1463 (O_1463,N_19765,N_19665);
or UO_1464 (O_1464,N_19815,N_19674);
nand UO_1465 (O_1465,N_19383,N_19454);
or UO_1466 (O_1466,N_19901,N_19536);
and UO_1467 (O_1467,N_19370,N_19225);
nor UO_1468 (O_1468,N_19931,N_19219);
and UO_1469 (O_1469,N_19431,N_19930);
xnor UO_1470 (O_1470,N_19607,N_19973);
nand UO_1471 (O_1471,N_19929,N_19363);
and UO_1472 (O_1472,N_19589,N_19985);
and UO_1473 (O_1473,N_19454,N_19203);
nor UO_1474 (O_1474,N_19343,N_19814);
or UO_1475 (O_1475,N_19891,N_19537);
nand UO_1476 (O_1476,N_19958,N_19358);
and UO_1477 (O_1477,N_19416,N_19865);
nand UO_1478 (O_1478,N_19819,N_19739);
nor UO_1479 (O_1479,N_19801,N_19838);
and UO_1480 (O_1480,N_19398,N_19843);
nor UO_1481 (O_1481,N_19611,N_19667);
xnor UO_1482 (O_1482,N_19657,N_19638);
xor UO_1483 (O_1483,N_19636,N_19974);
and UO_1484 (O_1484,N_19563,N_19583);
or UO_1485 (O_1485,N_19382,N_19732);
xor UO_1486 (O_1486,N_19293,N_19871);
or UO_1487 (O_1487,N_19533,N_19269);
and UO_1488 (O_1488,N_19931,N_19745);
and UO_1489 (O_1489,N_19462,N_19353);
xor UO_1490 (O_1490,N_19494,N_19946);
and UO_1491 (O_1491,N_19693,N_19611);
and UO_1492 (O_1492,N_19328,N_19621);
nand UO_1493 (O_1493,N_19306,N_19907);
nand UO_1494 (O_1494,N_19568,N_19658);
or UO_1495 (O_1495,N_19252,N_19422);
xnor UO_1496 (O_1496,N_19416,N_19513);
xor UO_1497 (O_1497,N_19674,N_19734);
or UO_1498 (O_1498,N_19580,N_19539);
nand UO_1499 (O_1499,N_19873,N_19391);
nor UO_1500 (O_1500,N_19296,N_19954);
nor UO_1501 (O_1501,N_19998,N_19953);
or UO_1502 (O_1502,N_19830,N_19738);
or UO_1503 (O_1503,N_19873,N_19387);
xnor UO_1504 (O_1504,N_19228,N_19932);
xnor UO_1505 (O_1505,N_19270,N_19383);
xnor UO_1506 (O_1506,N_19492,N_19756);
and UO_1507 (O_1507,N_19813,N_19908);
and UO_1508 (O_1508,N_19951,N_19232);
nand UO_1509 (O_1509,N_19316,N_19807);
and UO_1510 (O_1510,N_19283,N_19597);
nand UO_1511 (O_1511,N_19888,N_19996);
nand UO_1512 (O_1512,N_19856,N_19211);
and UO_1513 (O_1513,N_19978,N_19647);
xor UO_1514 (O_1514,N_19635,N_19201);
and UO_1515 (O_1515,N_19872,N_19368);
and UO_1516 (O_1516,N_19685,N_19429);
nand UO_1517 (O_1517,N_19284,N_19891);
nand UO_1518 (O_1518,N_19631,N_19661);
and UO_1519 (O_1519,N_19921,N_19503);
nor UO_1520 (O_1520,N_19305,N_19388);
and UO_1521 (O_1521,N_19375,N_19456);
or UO_1522 (O_1522,N_19522,N_19292);
and UO_1523 (O_1523,N_19921,N_19522);
and UO_1524 (O_1524,N_19213,N_19877);
nand UO_1525 (O_1525,N_19499,N_19976);
or UO_1526 (O_1526,N_19382,N_19807);
nand UO_1527 (O_1527,N_19816,N_19390);
and UO_1528 (O_1528,N_19727,N_19389);
nor UO_1529 (O_1529,N_19894,N_19384);
or UO_1530 (O_1530,N_19473,N_19917);
nand UO_1531 (O_1531,N_19844,N_19552);
and UO_1532 (O_1532,N_19353,N_19948);
nand UO_1533 (O_1533,N_19924,N_19459);
and UO_1534 (O_1534,N_19645,N_19467);
and UO_1535 (O_1535,N_19957,N_19592);
xnor UO_1536 (O_1536,N_19929,N_19800);
nand UO_1537 (O_1537,N_19277,N_19673);
xor UO_1538 (O_1538,N_19869,N_19765);
nor UO_1539 (O_1539,N_19915,N_19841);
nand UO_1540 (O_1540,N_19973,N_19987);
and UO_1541 (O_1541,N_19867,N_19326);
nor UO_1542 (O_1542,N_19677,N_19731);
xnor UO_1543 (O_1543,N_19296,N_19313);
and UO_1544 (O_1544,N_19393,N_19390);
nor UO_1545 (O_1545,N_19571,N_19383);
and UO_1546 (O_1546,N_19256,N_19556);
or UO_1547 (O_1547,N_19336,N_19228);
xor UO_1548 (O_1548,N_19219,N_19965);
nand UO_1549 (O_1549,N_19394,N_19659);
or UO_1550 (O_1550,N_19767,N_19614);
xnor UO_1551 (O_1551,N_19270,N_19314);
or UO_1552 (O_1552,N_19295,N_19795);
xnor UO_1553 (O_1553,N_19903,N_19417);
and UO_1554 (O_1554,N_19778,N_19754);
and UO_1555 (O_1555,N_19439,N_19690);
nor UO_1556 (O_1556,N_19571,N_19211);
nor UO_1557 (O_1557,N_19790,N_19913);
nand UO_1558 (O_1558,N_19790,N_19448);
nand UO_1559 (O_1559,N_19327,N_19243);
nor UO_1560 (O_1560,N_19268,N_19519);
nand UO_1561 (O_1561,N_19884,N_19576);
or UO_1562 (O_1562,N_19503,N_19952);
or UO_1563 (O_1563,N_19834,N_19610);
nand UO_1564 (O_1564,N_19604,N_19704);
or UO_1565 (O_1565,N_19691,N_19335);
or UO_1566 (O_1566,N_19303,N_19951);
or UO_1567 (O_1567,N_19256,N_19860);
nand UO_1568 (O_1568,N_19398,N_19337);
and UO_1569 (O_1569,N_19632,N_19603);
nor UO_1570 (O_1570,N_19435,N_19764);
and UO_1571 (O_1571,N_19203,N_19932);
xor UO_1572 (O_1572,N_19668,N_19615);
nand UO_1573 (O_1573,N_19886,N_19972);
xor UO_1574 (O_1574,N_19716,N_19797);
nor UO_1575 (O_1575,N_19405,N_19702);
nand UO_1576 (O_1576,N_19287,N_19204);
nor UO_1577 (O_1577,N_19645,N_19671);
nand UO_1578 (O_1578,N_19699,N_19214);
and UO_1579 (O_1579,N_19651,N_19673);
xnor UO_1580 (O_1580,N_19830,N_19472);
or UO_1581 (O_1581,N_19593,N_19715);
nand UO_1582 (O_1582,N_19454,N_19669);
nor UO_1583 (O_1583,N_19240,N_19817);
nor UO_1584 (O_1584,N_19609,N_19261);
nor UO_1585 (O_1585,N_19305,N_19254);
xnor UO_1586 (O_1586,N_19612,N_19480);
nand UO_1587 (O_1587,N_19693,N_19673);
and UO_1588 (O_1588,N_19590,N_19818);
or UO_1589 (O_1589,N_19612,N_19389);
nand UO_1590 (O_1590,N_19598,N_19400);
and UO_1591 (O_1591,N_19445,N_19549);
nor UO_1592 (O_1592,N_19200,N_19817);
xnor UO_1593 (O_1593,N_19417,N_19386);
nor UO_1594 (O_1594,N_19832,N_19444);
xor UO_1595 (O_1595,N_19951,N_19677);
nand UO_1596 (O_1596,N_19892,N_19511);
nand UO_1597 (O_1597,N_19403,N_19364);
nor UO_1598 (O_1598,N_19865,N_19238);
xor UO_1599 (O_1599,N_19855,N_19537);
and UO_1600 (O_1600,N_19270,N_19824);
or UO_1601 (O_1601,N_19891,N_19456);
xnor UO_1602 (O_1602,N_19596,N_19299);
nand UO_1603 (O_1603,N_19402,N_19260);
or UO_1604 (O_1604,N_19956,N_19550);
nor UO_1605 (O_1605,N_19290,N_19599);
nor UO_1606 (O_1606,N_19328,N_19658);
xor UO_1607 (O_1607,N_19603,N_19763);
and UO_1608 (O_1608,N_19434,N_19298);
and UO_1609 (O_1609,N_19972,N_19774);
nand UO_1610 (O_1610,N_19841,N_19781);
and UO_1611 (O_1611,N_19493,N_19744);
or UO_1612 (O_1612,N_19871,N_19956);
nor UO_1613 (O_1613,N_19260,N_19225);
xnor UO_1614 (O_1614,N_19245,N_19583);
nor UO_1615 (O_1615,N_19865,N_19744);
and UO_1616 (O_1616,N_19454,N_19625);
xor UO_1617 (O_1617,N_19484,N_19781);
nor UO_1618 (O_1618,N_19851,N_19366);
xnor UO_1619 (O_1619,N_19208,N_19457);
nor UO_1620 (O_1620,N_19631,N_19541);
nand UO_1621 (O_1621,N_19867,N_19476);
nor UO_1622 (O_1622,N_19903,N_19377);
or UO_1623 (O_1623,N_19290,N_19868);
nor UO_1624 (O_1624,N_19859,N_19687);
xnor UO_1625 (O_1625,N_19999,N_19219);
xor UO_1626 (O_1626,N_19327,N_19811);
nand UO_1627 (O_1627,N_19740,N_19961);
nand UO_1628 (O_1628,N_19932,N_19806);
or UO_1629 (O_1629,N_19605,N_19706);
and UO_1630 (O_1630,N_19597,N_19412);
and UO_1631 (O_1631,N_19241,N_19601);
and UO_1632 (O_1632,N_19404,N_19306);
xor UO_1633 (O_1633,N_19757,N_19873);
nand UO_1634 (O_1634,N_19469,N_19462);
nand UO_1635 (O_1635,N_19682,N_19249);
or UO_1636 (O_1636,N_19865,N_19844);
nand UO_1637 (O_1637,N_19373,N_19677);
nor UO_1638 (O_1638,N_19415,N_19638);
and UO_1639 (O_1639,N_19375,N_19351);
nand UO_1640 (O_1640,N_19697,N_19916);
xnor UO_1641 (O_1641,N_19786,N_19662);
and UO_1642 (O_1642,N_19526,N_19810);
nand UO_1643 (O_1643,N_19802,N_19784);
xnor UO_1644 (O_1644,N_19608,N_19496);
xor UO_1645 (O_1645,N_19900,N_19518);
nand UO_1646 (O_1646,N_19365,N_19503);
and UO_1647 (O_1647,N_19251,N_19324);
nor UO_1648 (O_1648,N_19894,N_19352);
nand UO_1649 (O_1649,N_19922,N_19755);
nor UO_1650 (O_1650,N_19462,N_19395);
nor UO_1651 (O_1651,N_19668,N_19399);
xnor UO_1652 (O_1652,N_19276,N_19686);
xor UO_1653 (O_1653,N_19549,N_19336);
xor UO_1654 (O_1654,N_19778,N_19974);
nor UO_1655 (O_1655,N_19717,N_19260);
nor UO_1656 (O_1656,N_19644,N_19789);
and UO_1657 (O_1657,N_19600,N_19370);
nor UO_1658 (O_1658,N_19678,N_19581);
and UO_1659 (O_1659,N_19889,N_19979);
xor UO_1660 (O_1660,N_19316,N_19901);
and UO_1661 (O_1661,N_19797,N_19782);
and UO_1662 (O_1662,N_19725,N_19307);
or UO_1663 (O_1663,N_19659,N_19815);
nor UO_1664 (O_1664,N_19679,N_19783);
xor UO_1665 (O_1665,N_19248,N_19245);
xor UO_1666 (O_1666,N_19861,N_19321);
nor UO_1667 (O_1667,N_19423,N_19616);
and UO_1668 (O_1668,N_19834,N_19561);
or UO_1669 (O_1669,N_19628,N_19985);
nor UO_1670 (O_1670,N_19275,N_19302);
and UO_1671 (O_1671,N_19965,N_19421);
nand UO_1672 (O_1672,N_19593,N_19444);
and UO_1673 (O_1673,N_19966,N_19251);
and UO_1674 (O_1674,N_19204,N_19325);
xnor UO_1675 (O_1675,N_19566,N_19949);
and UO_1676 (O_1676,N_19636,N_19829);
xnor UO_1677 (O_1677,N_19421,N_19518);
nor UO_1678 (O_1678,N_19947,N_19225);
nand UO_1679 (O_1679,N_19214,N_19434);
and UO_1680 (O_1680,N_19700,N_19551);
or UO_1681 (O_1681,N_19468,N_19383);
and UO_1682 (O_1682,N_19578,N_19898);
xnor UO_1683 (O_1683,N_19866,N_19753);
and UO_1684 (O_1684,N_19661,N_19227);
and UO_1685 (O_1685,N_19423,N_19387);
or UO_1686 (O_1686,N_19927,N_19781);
xor UO_1687 (O_1687,N_19242,N_19230);
nand UO_1688 (O_1688,N_19855,N_19530);
nor UO_1689 (O_1689,N_19239,N_19329);
xnor UO_1690 (O_1690,N_19864,N_19697);
or UO_1691 (O_1691,N_19887,N_19368);
nand UO_1692 (O_1692,N_19655,N_19907);
nand UO_1693 (O_1693,N_19899,N_19493);
nor UO_1694 (O_1694,N_19675,N_19509);
and UO_1695 (O_1695,N_19894,N_19214);
nand UO_1696 (O_1696,N_19736,N_19841);
nand UO_1697 (O_1697,N_19527,N_19278);
and UO_1698 (O_1698,N_19673,N_19859);
and UO_1699 (O_1699,N_19343,N_19775);
nand UO_1700 (O_1700,N_19765,N_19434);
nor UO_1701 (O_1701,N_19835,N_19405);
and UO_1702 (O_1702,N_19408,N_19238);
nand UO_1703 (O_1703,N_19615,N_19435);
nand UO_1704 (O_1704,N_19692,N_19383);
nand UO_1705 (O_1705,N_19249,N_19381);
and UO_1706 (O_1706,N_19726,N_19824);
or UO_1707 (O_1707,N_19708,N_19787);
or UO_1708 (O_1708,N_19486,N_19958);
xor UO_1709 (O_1709,N_19439,N_19919);
and UO_1710 (O_1710,N_19815,N_19699);
nand UO_1711 (O_1711,N_19659,N_19844);
and UO_1712 (O_1712,N_19302,N_19617);
xor UO_1713 (O_1713,N_19285,N_19367);
xor UO_1714 (O_1714,N_19417,N_19814);
nand UO_1715 (O_1715,N_19791,N_19327);
nand UO_1716 (O_1716,N_19905,N_19577);
nor UO_1717 (O_1717,N_19422,N_19639);
nand UO_1718 (O_1718,N_19942,N_19789);
or UO_1719 (O_1719,N_19469,N_19349);
nand UO_1720 (O_1720,N_19424,N_19601);
xor UO_1721 (O_1721,N_19596,N_19576);
nand UO_1722 (O_1722,N_19921,N_19772);
or UO_1723 (O_1723,N_19533,N_19275);
nor UO_1724 (O_1724,N_19303,N_19754);
nor UO_1725 (O_1725,N_19359,N_19539);
or UO_1726 (O_1726,N_19649,N_19955);
nand UO_1727 (O_1727,N_19564,N_19787);
nor UO_1728 (O_1728,N_19362,N_19344);
nand UO_1729 (O_1729,N_19436,N_19211);
nor UO_1730 (O_1730,N_19213,N_19846);
nand UO_1731 (O_1731,N_19391,N_19788);
nand UO_1732 (O_1732,N_19395,N_19306);
nand UO_1733 (O_1733,N_19378,N_19422);
xnor UO_1734 (O_1734,N_19581,N_19697);
nand UO_1735 (O_1735,N_19409,N_19624);
nand UO_1736 (O_1736,N_19293,N_19593);
and UO_1737 (O_1737,N_19926,N_19222);
nand UO_1738 (O_1738,N_19565,N_19635);
nor UO_1739 (O_1739,N_19838,N_19667);
and UO_1740 (O_1740,N_19272,N_19242);
or UO_1741 (O_1741,N_19920,N_19841);
nor UO_1742 (O_1742,N_19629,N_19473);
or UO_1743 (O_1743,N_19533,N_19445);
xor UO_1744 (O_1744,N_19522,N_19814);
and UO_1745 (O_1745,N_19431,N_19523);
xor UO_1746 (O_1746,N_19248,N_19520);
nor UO_1747 (O_1747,N_19851,N_19330);
nand UO_1748 (O_1748,N_19946,N_19429);
or UO_1749 (O_1749,N_19517,N_19825);
nor UO_1750 (O_1750,N_19207,N_19507);
or UO_1751 (O_1751,N_19692,N_19543);
nor UO_1752 (O_1752,N_19678,N_19469);
and UO_1753 (O_1753,N_19726,N_19285);
or UO_1754 (O_1754,N_19631,N_19936);
or UO_1755 (O_1755,N_19508,N_19541);
nor UO_1756 (O_1756,N_19617,N_19724);
nand UO_1757 (O_1757,N_19651,N_19694);
xor UO_1758 (O_1758,N_19528,N_19554);
nand UO_1759 (O_1759,N_19801,N_19533);
nor UO_1760 (O_1760,N_19360,N_19918);
nor UO_1761 (O_1761,N_19661,N_19697);
nor UO_1762 (O_1762,N_19671,N_19506);
nor UO_1763 (O_1763,N_19500,N_19451);
nand UO_1764 (O_1764,N_19218,N_19504);
or UO_1765 (O_1765,N_19362,N_19566);
xnor UO_1766 (O_1766,N_19873,N_19204);
nand UO_1767 (O_1767,N_19398,N_19230);
or UO_1768 (O_1768,N_19765,N_19752);
and UO_1769 (O_1769,N_19489,N_19896);
or UO_1770 (O_1770,N_19487,N_19970);
xnor UO_1771 (O_1771,N_19752,N_19256);
or UO_1772 (O_1772,N_19334,N_19652);
nor UO_1773 (O_1773,N_19239,N_19390);
and UO_1774 (O_1774,N_19702,N_19260);
and UO_1775 (O_1775,N_19261,N_19448);
and UO_1776 (O_1776,N_19793,N_19701);
nand UO_1777 (O_1777,N_19942,N_19903);
or UO_1778 (O_1778,N_19879,N_19610);
nand UO_1779 (O_1779,N_19548,N_19748);
nor UO_1780 (O_1780,N_19330,N_19283);
nand UO_1781 (O_1781,N_19213,N_19656);
and UO_1782 (O_1782,N_19967,N_19208);
and UO_1783 (O_1783,N_19751,N_19401);
nand UO_1784 (O_1784,N_19670,N_19531);
xnor UO_1785 (O_1785,N_19211,N_19599);
and UO_1786 (O_1786,N_19380,N_19688);
nor UO_1787 (O_1787,N_19544,N_19662);
nand UO_1788 (O_1788,N_19829,N_19626);
nor UO_1789 (O_1789,N_19702,N_19748);
and UO_1790 (O_1790,N_19352,N_19614);
nand UO_1791 (O_1791,N_19740,N_19938);
or UO_1792 (O_1792,N_19765,N_19551);
nand UO_1793 (O_1793,N_19959,N_19669);
nand UO_1794 (O_1794,N_19802,N_19400);
or UO_1795 (O_1795,N_19941,N_19563);
nand UO_1796 (O_1796,N_19539,N_19839);
nor UO_1797 (O_1797,N_19722,N_19362);
nand UO_1798 (O_1798,N_19759,N_19809);
nand UO_1799 (O_1799,N_19708,N_19943);
nor UO_1800 (O_1800,N_19246,N_19950);
xnor UO_1801 (O_1801,N_19629,N_19824);
nor UO_1802 (O_1802,N_19685,N_19322);
or UO_1803 (O_1803,N_19617,N_19590);
or UO_1804 (O_1804,N_19723,N_19488);
and UO_1805 (O_1805,N_19343,N_19949);
or UO_1806 (O_1806,N_19291,N_19905);
nand UO_1807 (O_1807,N_19435,N_19385);
xor UO_1808 (O_1808,N_19585,N_19756);
nor UO_1809 (O_1809,N_19871,N_19929);
nor UO_1810 (O_1810,N_19436,N_19233);
and UO_1811 (O_1811,N_19866,N_19254);
or UO_1812 (O_1812,N_19773,N_19750);
and UO_1813 (O_1813,N_19893,N_19648);
nor UO_1814 (O_1814,N_19369,N_19552);
nor UO_1815 (O_1815,N_19824,N_19686);
nand UO_1816 (O_1816,N_19942,N_19929);
nor UO_1817 (O_1817,N_19770,N_19219);
or UO_1818 (O_1818,N_19629,N_19655);
nor UO_1819 (O_1819,N_19297,N_19433);
nor UO_1820 (O_1820,N_19778,N_19641);
nor UO_1821 (O_1821,N_19982,N_19330);
xor UO_1822 (O_1822,N_19831,N_19786);
nor UO_1823 (O_1823,N_19497,N_19826);
or UO_1824 (O_1824,N_19504,N_19368);
nor UO_1825 (O_1825,N_19694,N_19262);
and UO_1826 (O_1826,N_19538,N_19368);
nand UO_1827 (O_1827,N_19734,N_19634);
or UO_1828 (O_1828,N_19271,N_19913);
and UO_1829 (O_1829,N_19693,N_19754);
and UO_1830 (O_1830,N_19840,N_19956);
xor UO_1831 (O_1831,N_19505,N_19374);
nor UO_1832 (O_1832,N_19350,N_19328);
and UO_1833 (O_1833,N_19674,N_19328);
nor UO_1834 (O_1834,N_19466,N_19607);
and UO_1835 (O_1835,N_19610,N_19492);
nand UO_1836 (O_1836,N_19879,N_19455);
xor UO_1837 (O_1837,N_19568,N_19322);
or UO_1838 (O_1838,N_19312,N_19422);
nor UO_1839 (O_1839,N_19465,N_19686);
or UO_1840 (O_1840,N_19860,N_19806);
nand UO_1841 (O_1841,N_19674,N_19277);
nand UO_1842 (O_1842,N_19909,N_19953);
xor UO_1843 (O_1843,N_19606,N_19455);
or UO_1844 (O_1844,N_19204,N_19736);
and UO_1845 (O_1845,N_19912,N_19968);
and UO_1846 (O_1846,N_19269,N_19271);
or UO_1847 (O_1847,N_19974,N_19774);
or UO_1848 (O_1848,N_19740,N_19378);
nand UO_1849 (O_1849,N_19426,N_19394);
nor UO_1850 (O_1850,N_19441,N_19535);
and UO_1851 (O_1851,N_19764,N_19868);
and UO_1852 (O_1852,N_19296,N_19441);
xnor UO_1853 (O_1853,N_19672,N_19337);
and UO_1854 (O_1854,N_19243,N_19955);
and UO_1855 (O_1855,N_19942,N_19383);
and UO_1856 (O_1856,N_19234,N_19470);
and UO_1857 (O_1857,N_19997,N_19336);
nand UO_1858 (O_1858,N_19986,N_19397);
nor UO_1859 (O_1859,N_19564,N_19531);
or UO_1860 (O_1860,N_19385,N_19867);
xnor UO_1861 (O_1861,N_19995,N_19486);
or UO_1862 (O_1862,N_19306,N_19515);
and UO_1863 (O_1863,N_19532,N_19253);
nand UO_1864 (O_1864,N_19267,N_19256);
xor UO_1865 (O_1865,N_19932,N_19534);
nand UO_1866 (O_1866,N_19644,N_19341);
xor UO_1867 (O_1867,N_19819,N_19435);
or UO_1868 (O_1868,N_19229,N_19668);
xnor UO_1869 (O_1869,N_19949,N_19412);
and UO_1870 (O_1870,N_19825,N_19275);
nor UO_1871 (O_1871,N_19960,N_19988);
nor UO_1872 (O_1872,N_19226,N_19531);
xnor UO_1873 (O_1873,N_19212,N_19500);
nor UO_1874 (O_1874,N_19580,N_19758);
nand UO_1875 (O_1875,N_19643,N_19970);
nand UO_1876 (O_1876,N_19542,N_19522);
nand UO_1877 (O_1877,N_19921,N_19989);
and UO_1878 (O_1878,N_19584,N_19320);
xnor UO_1879 (O_1879,N_19344,N_19898);
and UO_1880 (O_1880,N_19309,N_19959);
and UO_1881 (O_1881,N_19571,N_19358);
nor UO_1882 (O_1882,N_19400,N_19309);
nor UO_1883 (O_1883,N_19891,N_19450);
xor UO_1884 (O_1884,N_19889,N_19429);
and UO_1885 (O_1885,N_19486,N_19697);
xor UO_1886 (O_1886,N_19885,N_19778);
or UO_1887 (O_1887,N_19362,N_19296);
nor UO_1888 (O_1888,N_19595,N_19260);
or UO_1889 (O_1889,N_19719,N_19638);
nor UO_1890 (O_1890,N_19827,N_19295);
and UO_1891 (O_1891,N_19548,N_19783);
and UO_1892 (O_1892,N_19211,N_19407);
nor UO_1893 (O_1893,N_19748,N_19610);
nor UO_1894 (O_1894,N_19306,N_19960);
or UO_1895 (O_1895,N_19451,N_19546);
and UO_1896 (O_1896,N_19281,N_19305);
nor UO_1897 (O_1897,N_19620,N_19976);
nand UO_1898 (O_1898,N_19543,N_19888);
or UO_1899 (O_1899,N_19206,N_19717);
nor UO_1900 (O_1900,N_19940,N_19994);
and UO_1901 (O_1901,N_19434,N_19771);
xnor UO_1902 (O_1902,N_19994,N_19861);
nor UO_1903 (O_1903,N_19343,N_19292);
nor UO_1904 (O_1904,N_19925,N_19849);
xnor UO_1905 (O_1905,N_19454,N_19476);
xor UO_1906 (O_1906,N_19451,N_19288);
nor UO_1907 (O_1907,N_19831,N_19209);
or UO_1908 (O_1908,N_19954,N_19736);
nor UO_1909 (O_1909,N_19929,N_19951);
or UO_1910 (O_1910,N_19967,N_19287);
and UO_1911 (O_1911,N_19233,N_19235);
or UO_1912 (O_1912,N_19399,N_19296);
and UO_1913 (O_1913,N_19682,N_19394);
nand UO_1914 (O_1914,N_19984,N_19254);
or UO_1915 (O_1915,N_19361,N_19325);
and UO_1916 (O_1916,N_19253,N_19478);
and UO_1917 (O_1917,N_19693,N_19217);
or UO_1918 (O_1918,N_19544,N_19676);
and UO_1919 (O_1919,N_19859,N_19637);
and UO_1920 (O_1920,N_19458,N_19751);
and UO_1921 (O_1921,N_19392,N_19232);
and UO_1922 (O_1922,N_19407,N_19260);
xnor UO_1923 (O_1923,N_19966,N_19879);
nand UO_1924 (O_1924,N_19278,N_19835);
and UO_1925 (O_1925,N_19577,N_19888);
nor UO_1926 (O_1926,N_19399,N_19423);
nor UO_1927 (O_1927,N_19737,N_19664);
and UO_1928 (O_1928,N_19343,N_19812);
or UO_1929 (O_1929,N_19858,N_19477);
nand UO_1930 (O_1930,N_19404,N_19991);
nand UO_1931 (O_1931,N_19736,N_19986);
nor UO_1932 (O_1932,N_19201,N_19940);
nand UO_1933 (O_1933,N_19201,N_19472);
nand UO_1934 (O_1934,N_19407,N_19543);
and UO_1935 (O_1935,N_19693,N_19523);
nand UO_1936 (O_1936,N_19231,N_19920);
or UO_1937 (O_1937,N_19613,N_19578);
or UO_1938 (O_1938,N_19271,N_19922);
xnor UO_1939 (O_1939,N_19657,N_19954);
nand UO_1940 (O_1940,N_19391,N_19374);
xor UO_1941 (O_1941,N_19502,N_19946);
and UO_1942 (O_1942,N_19644,N_19287);
nor UO_1943 (O_1943,N_19219,N_19911);
and UO_1944 (O_1944,N_19409,N_19783);
or UO_1945 (O_1945,N_19272,N_19564);
xor UO_1946 (O_1946,N_19373,N_19962);
xor UO_1947 (O_1947,N_19437,N_19379);
nor UO_1948 (O_1948,N_19568,N_19557);
nor UO_1949 (O_1949,N_19235,N_19967);
and UO_1950 (O_1950,N_19825,N_19452);
nand UO_1951 (O_1951,N_19774,N_19500);
and UO_1952 (O_1952,N_19310,N_19372);
or UO_1953 (O_1953,N_19999,N_19896);
or UO_1954 (O_1954,N_19853,N_19869);
or UO_1955 (O_1955,N_19442,N_19819);
and UO_1956 (O_1956,N_19565,N_19403);
and UO_1957 (O_1957,N_19477,N_19936);
xnor UO_1958 (O_1958,N_19574,N_19541);
nand UO_1959 (O_1959,N_19766,N_19812);
or UO_1960 (O_1960,N_19909,N_19236);
nand UO_1961 (O_1961,N_19833,N_19663);
and UO_1962 (O_1962,N_19418,N_19755);
or UO_1963 (O_1963,N_19921,N_19742);
nand UO_1964 (O_1964,N_19768,N_19454);
nor UO_1965 (O_1965,N_19340,N_19521);
nand UO_1966 (O_1966,N_19967,N_19652);
or UO_1967 (O_1967,N_19343,N_19457);
nor UO_1968 (O_1968,N_19363,N_19580);
nor UO_1969 (O_1969,N_19972,N_19986);
or UO_1970 (O_1970,N_19899,N_19555);
nand UO_1971 (O_1971,N_19697,N_19566);
xnor UO_1972 (O_1972,N_19271,N_19215);
or UO_1973 (O_1973,N_19543,N_19490);
and UO_1974 (O_1974,N_19926,N_19501);
xnor UO_1975 (O_1975,N_19848,N_19792);
nand UO_1976 (O_1976,N_19815,N_19257);
and UO_1977 (O_1977,N_19637,N_19516);
or UO_1978 (O_1978,N_19347,N_19478);
or UO_1979 (O_1979,N_19587,N_19590);
or UO_1980 (O_1980,N_19234,N_19229);
or UO_1981 (O_1981,N_19599,N_19363);
nor UO_1982 (O_1982,N_19814,N_19941);
and UO_1983 (O_1983,N_19837,N_19868);
and UO_1984 (O_1984,N_19869,N_19385);
and UO_1985 (O_1985,N_19385,N_19626);
and UO_1986 (O_1986,N_19699,N_19324);
nor UO_1987 (O_1987,N_19436,N_19270);
or UO_1988 (O_1988,N_19586,N_19437);
and UO_1989 (O_1989,N_19996,N_19969);
nand UO_1990 (O_1990,N_19949,N_19368);
nand UO_1991 (O_1991,N_19247,N_19559);
or UO_1992 (O_1992,N_19972,N_19979);
nand UO_1993 (O_1993,N_19906,N_19889);
and UO_1994 (O_1994,N_19752,N_19341);
and UO_1995 (O_1995,N_19574,N_19321);
xor UO_1996 (O_1996,N_19323,N_19701);
nand UO_1997 (O_1997,N_19877,N_19588);
xnor UO_1998 (O_1998,N_19250,N_19308);
xnor UO_1999 (O_1999,N_19807,N_19523);
or UO_2000 (O_2000,N_19553,N_19231);
nor UO_2001 (O_2001,N_19798,N_19781);
and UO_2002 (O_2002,N_19963,N_19739);
nand UO_2003 (O_2003,N_19368,N_19584);
nor UO_2004 (O_2004,N_19984,N_19844);
nor UO_2005 (O_2005,N_19790,N_19335);
nand UO_2006 (O_2006,N_19496,N_19488);
nand UO_2007 (O_2007,N_19698,N_19219);
xor UO_2008 (O_2008,N_19270,N_19513);
xor UO_2009 (O_2009,N_19473,N_19916);
nand UO_2010 (O_2010,N_19851,N_19220);
nor UO_2011 (O_2011,N_19389,N_19694);
or UO_2012 (O_2012,N_19259,N_19413);
nor UO_2013 (O_2013,N_19670,N_19282);
or UO_2014 (O_2014,N_19786,N_19546);
nor UO_2015 (O_2015,N_19238,N_19479);
or UO_2016 (O_2016,N_19200,N_19493);
nand UO_2017 (O_2017,N_19355,N_19619);
and UO_2018 (O_2018,N_19870,N_19478);
xnor UO_2019 (O_2019,N_19354,N_19531);
nor UO_2020 (O_2020,N_19513,N_19651);
and UO_2021 (O_2021,N_19474,N_19934);
or UO_2022 (O_2022,N_19605,N_19904);
xor UO_2023 (O_2023,N_19904,N_19536);
xor UO_2024 (O_2024,N_19206,N_19672);
or UO_2025 (O_2025,N_19651,N_19557);
and UO_2026 (O_2026,N_19813,N_19816);
xor UO_2027 (O_2027,N_19948,N_19960);
nor UO_2028 (O_2028,N_19576,N_19639);
nor UO_2029 (O_2029,N_19875,N_19392);
or UO_2030 (O_2030,N_19723,N_19829);
or UO_2031 (O_2031,N_19414,N_19542);
nor UO_2032 (O_2032,N_19514,N_19411);
nand UO_2033 (O_2033,N_19698,N_19700);
xnor UO_2034 (O_2034,N_19361,N_19235);
nand UO_2035 (O_2035,N_19893,N_19656);
nand UO_2036 (O_2036,N_19202,N_19379);
nor UO_2037 (O_2037,N_19935,N_19211);
nor UO_2038 (O_2038,N_19759,N_19233);
nand UO_2039 (O_2039,N_19542,N_19479);
and UO_2040 (O_2040,N_19475,N_19357);
or UO_2041 (O_2041,N_19396,N_19885);
or UO_2042 (O_2042,N_19894,N_19590);
or UO_2043 (O_2043,N_19759,N_19425);
and UO_2044 (O_2044,N_19830,N_19631);
xor UO_2045 (O_2045,N_19332,N_19786);
nand UO_2046 (O_2046,N_19795,N_19393);
xor UO_2047 (O_2047,N_19812,N_19507);
nor UO_2048 (O_2048,N_19462,N_19870);
nand UO_2049 (O_2049,N_19755,N_19890);
and UO_2050 (O_2050,N_19400,N_19643);
nand UO_2051 (O_2051,N_19978,N_19610);
xor UO_2052 (O_2052,N_19320,N_19434);
xnor UO_2053 (O_2053,N_19603,N_19547);
nand UO_2054 (O_2054,N_19922,N_19851);
nand UO_2055 (O_2055,N_19445,N_19565);
nor UO_2056 (O_2056,N_19731,N_19389);
and UO_2057 (O_2057,N_19417,N_19891);
and UO_2058 (O_2058,N_19384,N_19854);
xor UO_2059 (O_2059,N_19793,N_19783);
and UO_2060 (O_2060,N_19843,N_19260);
nor UO_2061 (O_2061,N_19768,N_19203);
nor UO_2062 (O_2062,N_19922,N_19905);
nand UO_2063 (O_2063,N_19954,N_19889);
or UO_2064 (O_2064,N_19455,N_19578);
or UO_2065 (O_2065,N_19382,N_19568);
nand UO_2066 (O_2066,N_19942,N_19268);
nor UO_2067 (O_2067,N_19987,N_19822);
xnor UO_2068 (O_2068,N_19305,N_19911);
or UO_2069 (O_2069,N_19536,N_19643);
or UO_2070 (O_2070,N_19524,N_19537);
nor UO_2071 (O_2071,N_19705,N_19726);
or UO_2072 (O_2072,N_19436,N_19928);
nand UO_2073 (O_2073,N_19295,N_19495);
xnor UO_2074 (O_2074,N_19969,N_19970);
nand UO_2075 (O_2075,N_19416,N_19880);
nor UO_2076 (O_2076,N_19635,N_19640);
nand UO_2077 (O_2077,N_19599,N_19350);
and UO_2078 (O_2078,N_19390,N_19773);
and UO_2079 (O_2079,N_19232,N_19368);
and UO_2080 (O_2080,N_19946,N_19779);
nand UO_2081 (O_2081,N_19817,N_19386);
or UO_2082 (O_2082,N_19992,N_19509);
and UO_2083 (O_2083,N_19848,N_19637);
nand UO_2084 (O_2084,N_19308,N_19624);
nor UO_2085 (O_2085,N_19707,N_19237);
xnor UO_2086 (O_2086,N_19578,N_19902);
or UO_2087 (O_2087,N_19637,N_19965);
nand UO_2088 (O_2088,N_19444,N_19484);
nand UO_2089 (O_2089,N_19872,N_19750);
and UO_2090 (O_2090,N_19949,N_19835);
nand UO_2091 (O_2091,N_19615,N_19570);
nor UO_2092 (O_2092,N_19511,N_19433);
and UO_2093 (O_2093,N_19351,N_19667);
nand UO_2094 (O_2094,N_19784,N_19510);
nor UO_2095 (O_2095,N_19567,N_19493);
nor UO_2096 (O_2096,N_19896,N_19248);
or UO_2097 (O_2097,N_19236,N_19841);
nand UO_2098 (O_2098,N_19597,N_19984);
and UO_2099 (O_2099,N_19690,N_19425);
xor UO_2100 (O_2100,N_19670,N_19307);
xnor UO_2101 (O_2101,N_19888,N_19355);
xnor UO_2102 (O_2102,N_19812,N_19236);
or UO_2103 (O_2103,N_19679,N_19435);
nor UO_2104 (O_2104,N_19311,N_19905);
nor UO_2105 (O_2105,N_19437,N_19734);
and UO_2106 (O_2106,N_19573,N_19624);
nor UO_2107 (O_2107,N_19678,N_19661);
or UO_2108 (O_2108,N_19828,N_19453);
nand UO_2109 (O_2109,N_19338,N_19209);
or UO_2110 (O_2110,N_19619,N_19999);
xnor UO_2111 (O_2111,N_19663,N_19846);
nand UO_2112 (O_2112,N_19765,N_19974);
nor UO_2113 (O_2113,N_19777,N_19373);
nor UO_2114 (O_2114,N_19915,N_19976);
nand UO_2115 (O_2115,N_19902,N_19256);
or UO_2116 (O_2116,N_19832,N_19234);
nand UO_2117 (O_2117,N_19232,N_19622);
nor UO_2118 (O_2118,N_19718,N_19697);
nand UO_2119 (O_2119,N_19696,N_19903);
or UO_2120 (O_2120,N_19349,N_19313);
nand UO_2121 (O_2121,N_19980,N_19249);
xnor UO_2122 (O_2122,N_19989,N_19617);
xor UO_2123 (O_2123,N_19483,N_19738);
nand UO_2124 (O_2124,N_19432,N_19692);
and UO_2125 (O_2125,N_19421,N_19790);
xor UO_2126 (O_2126,N_19579,N_19680);
nor UO_2127 (O_2127,N_19767,N_19789);
nand UO_2128 (O_2128,N_19376,N_19596);
and UO_2129 (O_2129,N_19733,N_19216);
nor UO_2130 (O_2130,N_19513,N_19355);
nor UO_2131 (O_2131,N_19568,N_19492);
or UO_2132 (O_2132,N_19434,N_19516);
and UO_2133 (O_2133,N_19876,N_19937);
or UO_2134 (O_2134,N_19875,N_19238);
nand UO_2135 (O_2135,N_19367,N_19778);
nor UO_2136 (O_2136,N_19553,N_19997);
nor UO_2137 (O_2137,N_19793,N_19850);
and UO_2138 (O_2138,N_19255,N_19715);
and UO_2139 (O_2139,N_19859,N_19380);
nand UO_2140 (O_2140,N_19960,N_19576);
or UO_2141 (O_2141,N_19841,N_19685);
nor UO_2142 (O_2142,N_19382,N_19796);
nor UO_2143 (O_2143,N_19365,N_19839);
and UO_2144 (O_2144,N_19573,N_19354);
nand UO_2145 (O_2145,N_19358,N_19496);
or UO_2146 (O_2146,N_19996,N_19413);
nor UO_2147 (O_2147,N_19286,N_19315);
or UO_2148 (O_2148,N_19354,N_19975);
nor UO_2149 (O_2149,N_19543,N_19855);
nor UO_2150 (O_2150,N_19636,N_19758);
nand UO_2151 (O_2151,N_19368,N_19290);
and UO_2152 (O_2152,N_19701,N_19688);
nand UO_2153 (O_2153,N_19387,N_19930);
nor UO_2154 (O_2154,N_19418,N_19496);
nand UO_2155 (O_2155,N_19717,N_19962);
nor UO_2156 (O_2156,N_19594,N_19442);
xor UO_2157 (O_2157,N_19206,N_19827);
nand UO_2158 (O_2158,N_19320,N_19280);
nor UO_2159 (O_2159,N_19765,N_19543);
and UO_2160 (O_2160,N_19617,N_19747);
or UO_2161 (O_2161,N_19858,N_19281);
and UO_2162 (O_2162,N_19424,N_19243);
and UO_2163 (O_2163,N_19827,N_19924);
nand UO_2164 (O_2164,N_19874,N_19350);
nand UO_2165 (O_2165,N_19775,N_19761);
nand UO_2166 (O_2166,N_19934,N_19535);
or UO_2167 (O_2167,N_19916,N_19533);
or UO_2168 (O_2168,N_19366,N_19815);
and UO_2169 (O_2169,N_19873,N_19589);
or UO_2170 (O_2170,N_19376,N_19915);
nor UO_2171 (O_2171,N_19263,N_19554);
xnor UO_2172 (O_2172,N_19912,N_19260);
or UO_2173 (O_2173,N_19704,N_19443);
or UO_2174 (O_2174,N_19685,N_19358);
nand UO_2175 (O_2175,N_19687,N_19894);
nand UO_2176 (O_2176,N_19692,N_19332);
or UO_2177 (O_2177,N_19567,N_19629);
xor UO_2178 (O_2178,N_19350,N_19850);
nand UO_2179 (O_2179,N_19578,N_19751);
and UO_2180 (O_2180,N_19270,N_19505);
nor UO_2181 (O_2181,N_19918,N_19922);
nor UO_2182 (O_2182,N_19443,N_19207);
or UO_2183 (O_2183,N_19297,N_19346);
nand UO_2184 (O_2184,N_19895,N_19493);
or UO_2185 (O_2185,N_19574,N_19766);
and UO_2186 (O_2186,N_19713,N_19626);
and UO_2187 (O_2187,N_19404,N_19498);
or UO_2188 (O_2188,N_19280,N_19222);
and UO_2189 (O_2189,N_19646,N_19362);
or UO_2190 (O_2190,N_19785,N_19696);
xnor UO_2191 (O_2191,N_19271,N_19379);
xnor UO_2192 (O_2192,N_19930,N_19458);
or UO_2193 (O_2193,N_19366,N_19989);
nand UO_2194 (O_2194,N_19601,N_19368);
or UO_2195 (O_2195,N_19320,N_19769);
and UO_2196 (O_2196,N_19482,N_19967);
nor UO_2197 (O_2197,N_19685,N_19792);
nand UO_2198 (O_2198,N_19316,N_19318);
and UO_2199 (O_2199,N_19478,N_19887);
nand UO_2200 (O_2200,N_19622,N_19747);
xnor UO_2201 (O_2201,N_19918,N_19763);
xnor UO_2202 (O_2202,N_19711,N_19784);
xor UO_2203 (O_2203,N_19965,N_19928);
nand UO_2204 (O_2204,N_19407,N_19799);
and UO_2205 (O_2205,N_19956,N_19357);
and UO_2206 (O_2206,N_19546,N_19756);
xnor UO_2207 (O_2207,N_19486,N_19280);
or UO_2208 (O_2208,N_19290,N_19706);
and UO_2209 (O_2209,N_19636,N_19814);
or UO_2210 (O_2210,N_19622,N_19888);
xor UO_2211 (O_2211,N_19294,N_19969);
and UO_2212 (O_2212,N_19641,N_19460);
and UO_2213 (O_2213,N_19989,N_19346);
xnor UO_2214 (O_2214,N_19925,N_19654);
nor UO_2215 (O_2215,N_19749,N_19280);
and UO_2216 (O_2216,N_19396,N_19526);
nor UO_2217 (O_2217,N_19591,N_19484);
and UO_2218 (O_2218,N_19614,N_19527);
nor UO_2219 (O_2219,N_19260,N_19405);
xor UO_2220 (O_2220,N_19445,N_19722);
nor UO_2221 (O_2221,N_19733,N_19441);
or UO_2222 (O_2222,N_19894,N_19923);
or UO_2223 (O_2223,N_19891,N_19898);
nor UO_2224 (O_2224,N_19443,N_19787);
nand UO_2225 (O_2225,N_19879,N_19249);
nand UO_2226 (O_2226,N_19537,N_19864);
or UO_2227 (O_2227,N_19812,N_19216);
and UO_2228 (O_2228,N_19978,N_19862);
xor UO_2229 (O_2229,N_19673,N_19843);
nor UO_2230 (O_2230,N_19677,N_19958);
nor UO_2231 (O_2231,N_19567,N_19825);
xnor UO_2232 (O_2232,N_19916,N_19781);
or UO_2233 (O_2233,N_19620,N_19599);
nand UO_2234 (O_2234,N_19267,N_19299);
and UO_2235 (O_2235,N_19237,N_19683);
nand UO_2236 (O_2236,N_19962,N_19635);
xnor UO_2237 (O_2237,N_19919,N_19339);
xnor UO_2238 (O_2238,N_19516,N_19616);
and UO_2239 (O_2239,N_19848,N_19627);
or UO_2240 (O_2240,N_19408,N_19852);
nand UO_2241 (O_2241,N_19364,N_19867);
and UO_2242 (O_2242,N_19875,N_19485);
nand UO_2243 (O_2243,N_19579,N_19347);
or UO_2244 (O_2244,N_19904,N_19347);
xnor UO_2245 (O_2245,N_19750,N_19886);
and UO_2246 (O_2246,N_19938,N_19360);
and UO_2247 (O_2247,N_19349,N_19678);
and UO_2248 (O_2248,N_19986,N_19417);
nor UO_2249 (O_2249,N_19911,N_19489);
or UO_2250 (O_2250,N_19482,N_19932);
nor UO_2251 (O_2251,N_19709,N_19747);
and UO_2252 (O_2252,N_19425,N_19263);
xnor UO_2253 (O_2253,N_19783,N_19998);
xnor UO_2254 (O_2254,N_19703,N_19279);
and UO_2255 (O_2255,N_19542,N_19465);
xnor UO_2256 (O_2256,N_19567,N_19201);
or UO_2257 (O_2257,N_19778,N_19356);
xor UO_2258 (O_2258,N_19570,N_19210);
nand UO_2259 (O_2259,N_19312,N_19319);
and UO_2260 (O_2260,N_19756,N_19820);
xnor UO_2261 (O_2261,N_19978,N_19619);
or UO_2262 (O_2262,N_19269,N_19551);
nor UO_2263 (O_2263,N_19927,N_19778);
or UO_2264 (O_2264,N_19720,N_19566);
nand UO_2265 (O_2265,N_19910,N_19820);
and UO_2266 (O_2266,N_19846,N_19608);
and UO_2267 (O_2267,N_19440,N_19249);
and UO_2268 (O_2268,N_19230,N_19399);
nand UO_2269 (O_2269,N_19283,N_19958);
or UO_2270 (O_2270,N_19782,N_19635);
nor UO_2271 (O_2271,N_19737,N_19725);
and UO_2272 (O_2272,N_19692,N_19828);
and UO_2273 (O_2273,N_19964,N_19215);
xor UO_2274 (O_2274,N_19502,N_19953);
or UO_2275 (O_2275,N_19668,N_19994);
or UO_2276 (O_2276,N_19217,N_19739);
xor UO_2277 (O_2277,N_19558,N_19522);
and UO_2278 (O_2278,N_19780,N_19236);
and UO_2279 (O_2279,N_19564,N_19854);
nand UO_2280 (O_2280,N_19317,N_19800);
nor UO_2281 (O_2281,N_19843,N_19278);
nand UO_2282 (O_2282,N_19588,N_19825);
nor UO_2283 (O_2283,N_19284,N_19249);
or UO_2284 (O_2284,N_19255,N_19292);
and UO_2285 (O_2285,N_19300,N_19543);
and UO_2286 (O_2286,N_19371,N_19896);
xnor UO_2287 (O_2287,N_19467,N_19424);
and UO_2288 (O_2288,N_19895,N_19451);
or UO_2289 (O_2289,N_19959,N_19982);
nor UO_2290 (O_2290,N_19451,N_19465);
nand UO_2291 (O_2291,N_19216,N_19811);
xnor UO_2292 (O_2292,N_19365,N_19686);
nand UO_2293 (O_2293,N_19472,N_19924);
xnor UO_2294 (O_2294,N_19731,N_19884);
or UO_2295 (O_2295,N_19806,N_19884);
nor UO_2296 (O_2296,N_19376,N_19231);
and UO_2297 (O_2297,N_19664,N_19648);
xor UO_2298 (O_2298,N_19484,N_19470);
xor UO_2299 (O_2299,N_19570,N_19445);
nand UO_2300 (O_2300,N_19507,N_19363);
and UO_2301 (O_2301,N_19342,N_19747);
nand UO_2302 (O_2302,N_19902,N_19962);
nand UO_2303 (O_2303,N_19363,N_19473);
nor UO_2304 (O_2304,N_19362,N_19996);
nand UO_2305 (O_2305,N_19294,N_19286);
nand UO_2306 (O_2306,N_19600,N_19904);
and UO_2307 (O_2307,N_19922,N_19553);
nor UO_2308 (O_2308,N_19929,N_19433);
and UO_2309 (O_2309,N_19669,N_19931);
and UO_2310 (O_2310,N_19321,N_19808);
nor UO_2311 (O_2311,N_19960,N_19231);
and UO_2312 (O_2312,N_19951,N_19410);
xor UO_2313 (O_2313,N_19390,N_19687);
xor UO_2314 (O_2314,N_19582,N_19683);
or UO_2315 (O_2315,N_19250,N_19907);
nand UO_2316 (O_2316,N_19929,N_19644);
or UO_2317 (O_2317,N_19633,N_19699);
and UO_2318 (O_2318,N_19896,N_19678);
and UO_2319 (O_2319,N_19774,N_19404);
nor UO_2320 (O_2320,N_19898,N_19506);
nand UO_2321 (O_2321,N_19324,N_19900);
and UO_2322 (O_2322,N_19823,N_19309);
and UO_2323 (O_2323,N_19680,N_19664);
or UO_2324 (O_2324,N_19666,N_19953);
nor UO_2325 (O_2325,N_19575,N_19637);
xor UO_2326 (O_2326,N_19480,N_19580);
and UO_2327 (O_2327,N_19309,N_19366);
nand UO_2328 (O_2328,N_19762,N_19398);
nor UO_2329 (O_2329,N_19713,N_19931);
xnor UO_2330 (O_2330,N_19927,N_19415);
and UO_2331 (O_2331,N_19572,N_19860);
nand UO_2332 (O_2332,N_19756,N_19381);
nor UO_2333 (O_2333,N_19855,N_19371);
or UO_2334 (O_2334,N_19292,N_19859);
nand UO_2335 (O_2335,N_19596,N_19247);
nand UO_2336 (O_2336,N_19809,N_19632);
nand UO_2337 (O_2337,N_19311,N_19865);
xnor UO_2338 (O_2338,N_19626,N_19803);
or UO_2339 (O_2339,N_19582,N_19591);
nor UO_2340 (O_2340,N_19478,N_19458);
or UO_2341 (O_2341,N_19297,N_19416);
xor UO_2342 (O_2342,N_19760,N_19930);
and UO_2343 (O_2343,N_19636,N_19629);
xnor UO_2344 (O_2344,N_19922,N_19604);
or UO_2345 (O_2345,N_19925,N_19676);
xor UO_2346 (O_2346,N_19484,N_19255);
or UO_2347 (O_2347,N_19576,N_19231);
or UO_2348 (O_2348,N_19965,N_19663);
or UO_2349 (O_2349,N_19764,N_19887);
nand UO_2350 (O_2350,N_19806,N_19428);
nand UO_2351 (O_2351,N_19527,N_19509);
xor UO_2352 (O_2352,N_19284,N_19553);
xor UO_2353 (O_2353,N_19505,N_19876);
or UO_2354 (O_2354,N_19908,N_19321);
nand UO_2355 (O_2355,N_19734,N_19320);
nand UO_2356 (O_2356,N_19486,N_19852);
xnor UO_2357 (O_2357,N_19319,N_19682);
nand UO_2358 (O_2358,N_19792,N_19787);
or UO_2359 (O_2359,N_19257,N_19741);
nand UO_2360 (O_2360,N_19910,N_19583);
xor UO_2361 (O_2361,N_19604,N_19321);
or UO_2362 (O_2362,N_19408,N_19653);
or UO_2363 (O_2363,N_19582,N_19522);
nor UO_2364 (O_2364,N_19841,N_19310);
nand UO_2365 (O_2365,N_19354,N_19991);
nand UO_2366 (O_2366,N_19711,N_19861);
nor UO_2367 (O_2367,N_19954,N_19795);
nand UO_2368 (O_2368,N_19864,N_19684);
and UO_2369 (O_2369,N_19769,N_19816);
or UO_2370 (O_2370,N_19992,N_19914);
or UO_2371 (O_2371,N_19517,N_19707);
or UO_2372 (O_2372,N_19270,N_19870);
xor UO_2373 (O_2373,N_19254,N_19478);
nor UO_2374 (O_2374,N_19837,N_19582);
and UO_2375 (O_2375,N_19497,N_19925);
nor UO_2376 (O_2376,N_19527,N_19705);
xnor UO_2377 (O_2377,N_19486,N_19989);
xnor UO_2378 (O_2378,N_19640,N_19880);
xor UO_2379 (O_2379,N_19416,N_19663);
or UO_2380 (O_2380,N_19822,N_19216);
nor UO_2381 (O_2381,N_19914,N_19734);
and UO_2382 (O_2382,N_19401,N_19463);
and UO_2383 (O_2383,N_19896,N_19808);
nor UO_2384 (O_2384,N_19323,N_19599);
nor UO_2385 (O_2385,N_19319,N_19433);
nand UO_2386 (O_2386,N_19630,N_19343);
and UO_2387 (O_2387,N_19508,N_19290);
xor UO_2388 (O_2388,N_19237,N_19593);
and UO_2389 (O_2389,N_19860,N_19372);
and UO_2390 (O_2390,N_19234,N_19741);
nor UO_2391 (O_2391,N_19338,N_19202);
xor UO_2392 (O_2392,N_19265,N_19595);
xor UO_2393 (O_2393,N_19805,N_19285);
xnor UO_2394 (O_2394,N_19630,N_19564);
nand UO_2395 (O_2395,N_19404,N_19458);
nor UO_2396 (O_2396,N_19727,N_19334);
or UO_2397 (O_2397,N_19565,N_19329);
and UO_2398 (O_2398,N_19541,N_19407);
xor UO_2399 (O_2399,N_19599,N_19258);
nor UO_2400 (O_2400,N_19579,N_19385);
nand UO_2401 (O_2401,N_19431,N_19846);
nand UO_2402 (O_2402,N_19588,N_19600);
or UO_2403 (O_2403,N_19219,N_19289);
nand UO_2404 (O_2404,N_19237,N_19919);
or UO_2405 (O_2405,N_19872,N_19348);
nor UO_2406 (O_2406,N_19813,N_19880);
or UO_2407 (O_2407,N_19717,N_19451);
and UO_2408 (O_2408,N_19973,N_19608);
nand UO_2409 (O_2409,N_19306,N_19905);
nand UO_2410 (O_2410,N_19356,N_19654);
nand UO_2411 (O_2411,N_19223,N_19560);
nor UO_2412 (O_2412,N_19692,N_19443);
and UO_2413 (O_2413,N_19373,N_19966);
or UO_2414 (O_2414,N_19232,N_19846);
xnor UO_2415 (O_2415,N_19773,N_19498);
and UO_2416 (O_2416,N_19295,N_19984);
or UO_2417 (O_2417,N_19660,N_19956);
or UO_2418 (O_2418,N_19964,N_19448);
nand UO_2419 (O_2419,N_19455,N_19314);
or UO_2420 (O_2420,N_19427,N_19435);
nand UO_2421 (O_2421,N_19775,N_19627);
xor UO_2422 (O_2422,N_19237,N_19800);
xnor UO_2423 (O_2423,N_19861,N_19991);
nor UO_2424 (O_2424,N_19871,N_19762);
or UO_2425 (O_2425,N_19317,N_19602);
nor UO_2426 (O_2426,N_19213,N_19608);
and UO_2427 (O_2427,N_19888,N_19508);
or UO_2428 (O_2428,N_19852,N_19525);
nor UO_2429 (O_2429,N_19413,N_19311);
nor UO_2430 (O_2430,N_19571,N_19285);
and UO_2431 (O_2431,N_19332,N_19378);
or UO_2432 (O_2432,N_19778,N_19786);
nor UO_2433 (O_2433,N_19894,N_19448);
and UO_2434 (O_2434,N_19441,N_19370);
and UO_2435 (O_2435,N_19932,N_19843);
nor UO_2436 (O_2436,N_19295,N_19556);
xnor UO_2437 (O_2437,N_19249,N_19215);
or UO_2438 (O_2438,N_19274,N_19784);
or UO_2439 (O_2439,N_19502,N_19790);
nor UO_2440 (O_2440,N_19550,N_19976);
and UO_2441 (O_2441,N_19295,N_19882);
and UO_2442 (O_2442,N_19384,N_19568);
xor UO_2443 (O_2443,N_19321,N_19879);
nor UO_2444 (O_2444,N_19450,N_19696);
nor UO_2445 (O_2445,N_19466,N_19217);
xnor UO_2446 (O_2446,N_19441,N_19945);
and UO_2447 (O_2447,N_19909,N_19210);
nor UO_2448 (O_2448,N_19467,N_19286);
or UO_2449 (O_2449,N_19461,N_19534);
nand UO_2450 (O_2450,N_19610,N_19305);
xor UO_2451 (O_2451,N_19511,N_19582);
or UO_2452 (O_2452,N_19712,N_19602);
or UO_2453 (O_2453,N_19542,N_19947);
and UO_2454 (O_2454,N_19425,N_19422);
xor UO_2455 (O_2455,N_19661,N_19600);
nor UO_2456 (O_2456,N_19206,N_19502);
and UO_2457 (O_2457,N_19928,N_19797);
or UO_2458 (O_2458,N_19614,N_19512);
or UO_2459 (O_2459,N_19747,N_19630);
nor UO_2460 (O_2460,N_19992,N_19652);
or UO_2461 (O_2461,N_19203,N_19532);
nor UO_2462 (O_2462,N_19820,N_19927);
nand UO_2463 (O_2463,N_19911,N_19740);
and UO_2464 (O_2464,N_19638,N_19308);
xnor UO_2465 (O_2465,N_19848,N_19395);
or UO_2466 (O_2466,N_19684,N_19812);
nand UO_2467 (O_2467,N_19205,N_19729);
or UO_2468 (O_2468,N_19648,N_19283);
or UO_2469 (O_2469,N_19619,N_19870);
and UO_2470 (O_2470,N_19556,N_19529);
nand UO_2471 (O_2471,N_19209,N_19868);
or UO_2472 (O_2472,N_19460,N_19203);
nand UO_2473 (O_2473,N_19771,N_19304);
and UO_2474 (O_2474,N_19318,N_19273);
and UO_2475 (O_2475,N_19799,N_19968);
nand UO_2476 (O_2476,N_19830,N_19526);
xor UO_2477 (O_2477,N_19673,N_19523);
or UO_2478 (O_2478,N_19227,N_19900);
xor UO_2479 (O_2479,N_19373,N_19265);
or UO_2480 (O_2480,N_19876,N_19902);
and UO_2481 (O_2481,N_19907,N_19386);
nor UO_2482 (O_2482,N_19204,N_19474);
nand UO_2483 (O_2483,N_19516,N_19999);
nor UO_2484 (O_2484,N_19277,N_19965);
xor UO_2485 (O_2485,N_19443,N_19432);
xnor UO_2486 (O_2486,N_19339,N_19283);
and UO_2487 (O_2487,N_19646,N_19404);
or UO_2488 (O_2488,N_19295,N_19885);
and UO_2489 (O_2489,N_19714,N_19428);
nand UO_2490 (O_2490,N_19834,N_19470);
xor UO_2491 (O_2491,N_19877,N_19230);
and UO_2492 (O_2492,N_19773,N_19643);
xnor UO_2493 (O_2493,N_19778,N_19263);
xor UO_2494 (O_2494,N_19965,N_19285);
xor UO_2495 (O_2495,N_19882,N_19891);
and UO_2496 (O_2496,N_19334,N_19829);
xnor UO_2497 (O_2497,N_19751,N_19776);
and UO_2498 (O_2498,N_19905,N_19451);
xnor UO_2499 (O_2499,N_19249,N_19219);
endmodule