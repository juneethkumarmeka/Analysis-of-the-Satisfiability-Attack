module basic_1000_10000_1500_5_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_924,In_359);
nor U1 (N_1,In_831,In_634);
and U2 (N_2,In_483,In_139);
nand U3 (N_3,In_234,In_524);
and U4 (N_4,In_218,In_130);
or U5 (N_5,In_616,In_847);
nor U6 (N_6,In_909,In_923);
and U7 (N_7,In_872,In_513);
nor U8 (N_8,In_955,In_785);
nor U9 (N_9,In_538,In_195);
and U10 (N_10,In_669,In_410);
and U11 (N_11,In_986,In_638);
and U12 (N_12,In_445,In_942);
nor U13 (N_13,In_784,In_788);
or U14 (N_14,In_470,In_147);
and U15 (N_15,In_748,In_352);
nor U16 (N_16,In_309,In_862);
nor U17 (N_17,In_506,In_225);
nor U18 (N_18,In_542,In_750);
nor U19 (N_19,In_881,In_260);
nand U20 (N_20,In_546,In_489);
or U21 (N_21,In_471,In_912);
nor U22 (N_22,In_995,In_796);
and U23 (N_23,In_484,In_899);
nand U24 (N_24,In_30,In_49);
or U25 (N_25,In_477,In_536);
nor U26 (N_26,In_464,In_647);
or U27 (N_27,In_209,In_822);
nand U28 (N_28,In_937,In_168);
nor U29 (N_29,In_810,In_361);
nand U30 (N_30,In_947,In_722);
nor U31 (N_31,In_89,In_579);
or U32 (N_32,In_167,In_12);
or U33 (N_33,In_408,In_594);
nand U34 (N_34,In_610,In_375);
nand U35 (N_35,In_52,In_901);
or U36 (N_36,In_206,In_282);
nand U37 (N_37,In_196,In_576);
nand U38 (N_38,In_572,In_349);
nor U39 (N_39,In_879,In_162);
nor U40 (N_40,In_5,In_441);
xnor U41 (N_41,In_957,In_312);
nor U42 (N_42,In_90,In_820);
and U43 (N_43,In_278,In_857);
nor U44 (N_44,In_421,In_717);
nand U45 (N_45,In_617,In_79);
nor U46 (N_46,In_466,In_902);
nand U47 (N_47,In_172,In_863);
nand U48 (N_48,In_759,In_326);
xnor U49 (N_49,In_559,In_545);
and U50 (N_50,In_732,In_36);
nor U51 (N_51,In_733,In_224);
nand U52 (N_52,In_516,In_931);
or U53 (N_53,In_528,In_161);
or U54 (N_54,In_587,In_562);
or U55 (N_55,In_198,In_230);
nor U56 (N_56,In_662,In_391);
or U57 (N_57,In_603,In_56);
nand U58 (N_58,In_121,In_637);
nand U59 (N_59,In_906,In_91);
nand U60 (N_60,In_343,In_183);
nor U61 (N_61,In_884,In_86);
or U62 (N_62,In_381,In_83);
nand U63 (N_63,In_591,In_756);
nor U64 (N_64,In_643,In_80);
or U65 (N_65,In_140,In_734);
and U66 (N_66,In_127,In_987);
and U67 (N_67,In_978,In_549);
nor U68 (N_68,In_488,In_100);
and U69 (N_69,In_163,In_865);
or U70 (N_70,In_60,In_395);
xor U71 (N_71,In_124,In_934);
or U72 (N_72,In_404,In_727);
and U73 (N_73,In_745,In_74);
or U74 (N_74,In_888,In_51);
or U75 (N_75,In_936,In_688);
and U76 (N_76,In_181,In_629);
or U77 (N_77,In_926,In_573);
and U78 (N_78,In_741,In_263);
nor U79 (N_79,In_233,In_128);
and U80 (N_80,In_624,In_744);
or U81 (N_81,In_994,In_311);
nand U82 (N_82,In_406,In_840);
or U83 (N_83,In_21,In_141);
and U84 (N_84,In_649,In_363);
nor U85 (N_85,In_323,In_682);
and U86 (N_86,In_595,In_868);
nor U87 (N_87,In_523,In_302);
nor U88 (N_88,In_802,In_313);
nand U89 (N_89,In_367,In_422);
or U90 (N_90,In_296,In_859);
and U91 (N_91,In_943,In_724);
nand U92 (N_92,In_848,In_336);
and U93 (N_93,In_419,In_818);
nor U94 (N_94,In_277,In_671);
and U95 (N_95,In_844,In_775);
or U96 (N_96,In_673,In_885);
and U97 (N_97,In_574,In_625);
or U98 (N_98,In_84,In_384);
and U99 (N_99,In_284,In_275);
and U100 (N_100,In_14,In_837);
nand U101 (N_101,In_37,In_917);
or U102 (N_102,In_255,In_203);
nand U103 (N_103,In_935,In_606);
nand U104 (N_104,In_258,In_628);
or U105 (N_105,In_158,In_246);
or U106 (N_106,In_96,In_499);
or U107 (N_107,In_244,In_808);
nand U108 (N_108,In_265,In_658);
nand U109 (N_109,In_675,In_256);
and U110 (N_110,In_425,In_269);
nand U111 (N_111,In_589,In_915);
and U112 (N_112,In_622,In_813);
nand U113 (N_113,In_544,In_993);
and U114 (N_114,In_723,In_799);
nand U115 (N_115,In_778,In_151);
nand U116 (N_116,In_975,In_201);
nor U117 (N_117,In_239,In_650);
nand U118 (N_118,In_880,In_997);
and U119 (N_119,In_715,In_611);
and U120 (N_120,In_790,In_67);
or U121 (N_121,In_385,In_135);
or U122 (N_122,In_394,In_533);
nand U123 (N_123,In_792,In_458);
nor U124 (N_124,In_580,In_832);
and U125 (N_125,In_783,In_432);
or U126 (N_126,In_905,In_436);
nand U127 (N_127,In_919,In_362);
nand U128 (N_128,In_821,In_678);
nor U129 (N_129,In_150,In_129);
and U130 (N_130,In_491,In_984);
nand U131 (N_131,In_571,In_786);
or U132 (N_132,In_73,In_189);
nor U133 (N_133,In_358,In_961);
xnor U134 (N_134,In_596,In_766);
nand U135 (N_135,In_493,In_426);
or U136 (N_136,In_485,In_892);
xnor U137 (N_137,In_19,In_386);
nor U138 (N_138,In_213,In_366);
nor U139 (N_139,In_329,In_204);
nand U140 (N_140,In_566,In_428);
nor U141 (N_141,In_304,In_660);
xnor U142 (N_142,In_605,In_478);
nand U143 (N_143,In_219,In_351);
or U144 (N_144,In_577,In_765);
and U145 (N_145,In_920,In_459);
and U146 (N_146,In_679,In_243);
nand U147 (N_147,In_854,In_316);
nor U148 (N_148,In_388,In_583);
or U149 (N_149,In_858,In_298);
or U150 (N_150,In_989,In_187);
nand U151 (N_151,In_701,In_803);
nor U152 (N_152,In_922,In_122);
and U153 (N_153,In_132,In_950);
nor U154 (N_154,In_521,In_856);
or U155 (N_155,In_969,In_293);
and U156 (N_156,In_45,In_43);
nor U157 (N_157,In_382,In_8);
or U158 (N_158,In_928,In_55);
nor U159 (N_159,In_486,In_289);
or U160 (N_160,In_903,In_104);
nand U161 (N_161,In_393,In_816);
and U162 (N_162,In_805,In_76);
nand U163 (N_163,In_268,In_970);
nand U164 (N_164,In_280,In_146);
nor U165 (N_165,In_208,In_563);
and U166 (N_166,In_520,In_780);
or U167 (N_167,In_592,In_214);
xnor U168 (N_168,In_779,In_554);
nand U169 (N_169,In_306,In_613);
and U170 (N_170,In_27,In_415);
nor U171 (N_171,In_692,In_702);
and U172 (N_172,In_346,In_24);
or U173 (N_173,In_15,In_640);
and U174 (N_174,In_855,In_743);
nand U175 (N_175,In_473,In_921);
or U176 (N_176,In_898,In_954);
and U177 (N_177,In_253,In_142);
nand U178 (N_178,In_504,In_370);
or U179 (N_179,In_320,In_494);
and U180 (N_180,In_996,In_264);
or U181 (N_181,In_811,In_69);
nand U182 (N_182,In_31,In_409);
nor U183 (N_183,In_283,In_70);
or U184 (N_184,In_703,In_690);
nor U185 (N_185,In_497,In_353);
and U186 (N_186,In_238,In_951);
nor U187 (N_187,In_891,In_145);
and U188 (N_188,In_449,In_740);
nor U189 (N_189,In_718,In_755);
or U190 (N_190,In_13,In_553);
or U191 (N_191,In_693,In_895);
or U192 (N_192,In_77,In_64);
or U193 (N_193,In_149,In_273);
or U194 (N_194,In_392,In_365);
nand U195 (N_195,In_861,In_990);
nor U196 (N_196,In_34,In_719);
nor U197 (N_197,In_65,In_871);
and U198 (N_198,In_830,In_492);
or U199 (N_199,In_590,In_368);
and U200 (N_200,In_672,In_886);
and U201 (N_201,In_467,In_503);
nand U202 (N_202,In_231,In_804);
and U203 (N_203,In_800,In_176);
or U204 (N_204,In_998,In_869);
or U205 (N_205,In_976,In_41);
or U206 (N_206,In_179,In_911);
nand U207 (N_207,In_946,In_893);
or U208 (N_208,In_442,In_767);
nand U209 (N_209,In_860,In_737);
or U210 (N_210,In_338,In_570);
or U211 (N_211,In_102,In_824);
nand U212 (N_212,In_397,In_763);
nand U213 (N_213,In_413,In_794);
nand U214 (N_214,In_633,In_7);
or U215 (N_215,In_889,In_332);
and U216 (N_216,In_833,In_61);
and U217 (N_217,In_465,In_838);
nor U218 (N_218,In_959,In_532);
and U219 (N_219,In_823,In_707);
nand U220 (N_220,In_424,In_72);
and U221 (N_221,In_548,In_58);
and U222 (N_222,In_330,In_314);
nor U223 (N_223,In_380,In_531);
xnor U224 (N_224,In_918,In_757);
nand U225 (N_225,In_152,In_248);
nand U226 (N_226,In_845,In_94);
nand U227 (N_227,In_771,In_328);
nor U228 (N_228,In_112,In_908);
or U229 (N_229,In_348,In_581);
or U230 (N_230,In_654,In_774);
nor U231 (N_231,In_736,In_819);
nor U232 (N_232,In_347,In_155);
nand U233 (N_233,In_95,In_192);
and U234 (N_234,In_262,In_315);
nor U235 (N_235,In_828,In_188);
nor U236 (N_236,In_968,In_117);
nor U237 (N_237,In_237,In_983);
or U238 (N_238,In_725,In_753);
or U239 (N_239,In_655,In_641);
and U240 (N_240,In_694,In_227);
and U241 (N_241,In_245,In_512);
nor U242 (N_242,In_726,In_480);
nor U243 (N_243,In_383,In_877);
and U244 (N_244,In_403,In_105);
and U245 (N_245,In_476,In_882);
and U246 (N_246,In_297,In_223);
or U247 (N_247,In_564,In_463);
nand U248 (N_248,In_184,In_460);
or U249 (N_249,In_212,In_522);
nand U250 (N_250,In_502,In_171);
and U251 (N_251,In_791,In_390);
nand U252 (N_252,In_541,In_364);
xnor U253 (N_253,In_527,In_705);
nand U254 (N_254,In_608,In_319);
or U255 (N_255,In_875,In_683);
nand U256 (N_256,In_826,In_604);
or U257 (N_257,In_666,In_334);
nand U258 (N_258,In_992,In_839);
and U259 (N_259,In_138,In_980);
nand U260 (N_260,In_170,In_399);
nand U261 (N_261,In_713,In_389);
and U262 (N_262,In_157,In_310);
nor U263 (N_263,In_53,In_691);
nand U264 (N_264,In_420,In_300);
nor U265 (N_265,In_668,In_501);
nor U266 (N_266,In_433,In_874);
and U267 (N_267,In_963,In_475);
nor U268 (N_268,In_526,In_118);
or U269 (N_269,In_23,In_99);
or U270 (N_270,In_461,In_39);
nand U271 (N_271,In_933,In_232);
xor U272 (N_272,In_677,In_207);
or U273 (N_273,In_295,In_164);
or U274 (N_274,In_735,In_93);
and U275 (N_275,In_229,In_444);
nand U276 (N_276,In_761,In_896);
or U277 (N_277,In_772,In_795);
nor U278 (N_278,In_134,In_517);
and U279 (N_279,In_123,In_156);
nand U280 (N_280,In_582,In_48);
nand U281 (N_281,In_585,In_639);
and U282 (N_282,In_2,In_887);
or U283 (N_283,In_175,In_469);
and U284 (N_284,In_327,In_852);
nand U285 (N_285,In_561,In_894);
or U286 (N_286,In_619,In_355);
and U287 (N_287,In_977,In_9);
nand U288 (N_288,In_716,In_401);
or U289 (N_289,In_240,In_510);
and U290 (N_290,In_414,In_940);
or U291 (N_291,In_846,In_398);
nand U292 (N_292,In_948,In_435);
or U293 (N_293,In_40,In_850);
nand U294 (N_294,In_674,In_210);
and U295 (N_295,In_169,In_279);
or U296 (N_296,In_738,In_866);
and U297 (N_297,In_308,In_720);
and U298 (N_298,In_952,In_601);
or U299 (N_299,In_801,In_222);
nand U300 (N_300,In_182,In_930);
nand U301 (N_301,In_789,In_63);
or U302 (N_302,In_956,In_988);
nor U303 (N_303,In_843,In_339);
nor U304 (N_304,In_614,In_372);
and U305 (N_305,In_285,In_114);
nor U306 (N_306,In_126,In_377);
nand U307 (N_307,In_939,In_318);
nand U308 (N_308,In_71,In_103);
and U309 (N_309,In_842,In_305);
nor U310 (N_310,In_773,In_965);
and U311 (N_311,In_38,In_999);
and U312 (N_312,In_173,In_119);
nand U313 (N_313,In_496,In_670);
nor U314 (N_314,In_960,In_864);
nand U315 (N_315,In_281,In_81);
or U316 (N_316,In_534,In_371);
and U317 (N_317,In_651,In_468);
or U318 (N_318,In_787,In_217);
nor U319 (N_319,In_402,In_498);
or U320 (N_320,In_247,In_46);
and U321 (N_321,In_817,In_809);
nor U322 (N_322,In_276,In_452);
or U323 (N_323,In_695,In_430);
xnor U324 (N_324,In_749,In_700);
nor U325 (N_325,In_697,In_665);
or U326 (N_326,In_760,In_199);
and U327 (N_327,In_797,In_221);
or U328 (N_328,In_472,In_913);
xor U329 (N_329,In_714,In_360);
nand U330 (N_330,In_907,In_254);
xnor U331 (N_331,In_423,In_450);
nor U332 (N_332,In_979,In_730);
nand U333 (N_333,In_378,In_18);
or U334 (N_334,In_621,In_890);
and U335 (N_335,In_626,In_661);
or U336 (N_336,In_337,In_518);
or U337 (N_337,In_405,In_22);
or U338 (N_338,In_66,In_897);
nor U339 (N_339,In_333,In_274);
nand U340 (N_340,In_689,In_547);
nor U341 (N_341,In_341,In_825);
xor U342 (N_342,In_652,In_479);
or U343 (N_343,In_57,In_967);
nand U344 (N_344,In_434,In_437);
or U345 (N_345,In_953,In_962);
and U346 (N_346,In_565,In_560);
and U347 (N_347,In_200,In_567);
and U348 (N_348,In_431,In_418);
or U349 (N_349,In_288,In_412);
or U350 (N_350,In_659,In_656);
and U351 (N_351,In_762,In_374);
nor U352 (N_352,In_829,In_299);
nor U353 (N_353,In_120,In_680);
and U354 (N_354,In_453,In_505);
nand U355 (N_355,In_107,In_687);
nor U356 (N_356,In_653,In_340);
and U357 (N_357,In_974,In_109);
xnor U358 (N_358,In_964,In_446);
and U359 (N_359,In_710,In_938);
nor U360 (N_360,In_742,In_75);
nand U361 (N_361,In_32,In_174);
nand U362 (N_362,In_500,In_747);
and U363 (N_363,In_270,In_344);
nand U364 (N_364,In_849,In_853);
or U365 (N_365,In_443,In_33);
and U366 (N_366,In_242,In_317);
nand U367 (N_367,In_286,In_111);
or U368 (N_368,In_685,In_618);
nor U369 (N_369,In_981,In_746);
or U370 (N_370,In_927,In_870);
nor U371 (N_371,In_396,In_525);
and U372 (N_372,In_664,In_113);
and U373 (N_373,In_115,In_646);
nor U374 (N_374,In_407,In_602);
or U375 (N_375,In_751,In_447);
and U376 (N_376,In_944,In_807);
nand U377 (N_377,In_711,In_97);
nor U378 (N_378,In_54,In_728);
or U379 (N_379,In_148,In_376);
or U380 (N_380,In_982,In_454);
or U381 (N_381,In_159,In_914);
nor U382 (N_382,In_627,In_294);
nor U383 (N_383,In_178,In_110);
and U384 (N_384,In_416,In_708);
nand U385 (N_385,In_190,In_236);
and U386 (N_386,In_136,In_68);
nor U387 (N_387,In_211,In_438);
nand U388 (N_388,In_681,In_515);
and U389 (N_389,In_607,In_648);
nor U390 (N_390,In_593,In_644);
and U391 (N_391,In_228,In_557);
or U392 (N_392,In_949,In_44);
xnor U393 (N_393,In_645,In_116);
nand U394 (N_394,In_448,In_770);
and U395 (N_395,In_731,In_568);
and U396 (N_396,In_17,In_815);
nor U397 (N_397,In_0,In_867);
nor U398 (N_398,In_191,In_578);
and U399 (N_399,In_144,In_180);
xor U400 (N_400,In_883,In_417);
nor U401 (N_401,In_598,In_600);
or U402 (N_402,In_623,In_958);
and U403 (N_403,In_514,In_985);
nor U404 (N_404,In_101,In_88);
and U405 (N_405,In_345,In_539);
or U406 (N_406,In_322,In_481);
nand U407 (N_407,In_657,In_92);
xor U408 (N_408,In_663,In_400);
nor U409 (N_409,In_354,In_509);
or U410 (N_410,In_325,In_490);
nand U411 (N_411,In_782,In_586);
nand U412 (N_412,In_153,In_457);
and U413 (N_413,In_552,In_635);
and U414 (N_414,In_324,In_287);
nand U415 (N_415,In_456,In_427);
nor U416 (N_416,In_972,In_781);
nand U417 (N_417,In_356,In_451);
or U418 (N_418,In_303,In_851);
or U419 (N_419,In_686,In_615);
nor U420 (N_420,In_335,In_878);
or U421 (N_421,In_597,In_59);
and U422 (N_422,In_511,In_482);
and U423 (N_423,In_945,In_82);
nand U424 (N_424,In_251,In_307);
or U425 (N_425,In_575,In_558);
or U426 (N_426,In_971,In_186);
nand U427 (N_427,In_551,In_729);
or U428 (N_428,In_798,In_642);
nor U429 (N_429,In_676,In_440);
and U430 (N_430,In_556,In_25);
nor U431 (N_431,In_267,In_125);
nor U432 (N_432,In_814,In_160);
and U433 (N_433,In_133,In_706);
nor U434 (N_434,In_143,In_487);
nand U435 (N_435,In_272,In_194);
and U436 (N_436,In_754,In_612);
or U437 (N_437,In_609,In_636);
nand U438 (N_438,In_537,In_973);
nand U439 (N_439,In_966,In_98);
and U440 (N_440,In_712,In_709);
or U441 (N_441,In_387,In_193);
nand U442 (N_442,In_220,In_555);
and U443 (N_443,In_26,In_929);
or U444 (N_444,In_916,In_632);
nand U445 (N_445,In_4,In_42);
and U446 (N_446,In_550,In_271);
nand U447 (N_447,In_78,In_812);
and U448 (N_448,In_529,In_793);
nor U449 (N_449,In_185,In_290);
or U450 (N_450,In_321,In_292);
xor U451 (N_451,In_991,In_941);
nor U452 (N_452,In_599,In_462);
or U453 (N_453,In_543,In_29);
or U454 (N_454,In_291,In_777);
or U455 (N_455,In_620,In_50);
nand U456 (N_456,In_507,In_530);
nand U457 (N_457,In_16,In_721);
nand U458 (N_458,In_835,In_569);
or U459 (N_459,In_357,In_630);
nor U460 (N_460,In_495,In_667);
and U461 (N_461,In_1,In_301);
or U462 (N_462,In_28,In_205);
nand U463 (N_463,In_841,In_519);
and U464 (N_464,In_252,In_588);
nor U465 (N_465,In_108,In_429);
nand U466 (N_466,In_177,In_87);
xor U467 (N_467,In_369,In_373);
nand U468 (N_468,In_876,In_910);
or U469 (N_469,In_873,In_584);
nor U470 (N_470,In_768,In_106);
nor U471 (N_471,In_535,In_215);
or U472 (N_472,In_11,In_166);
and U473 (N_473,In_540,In_704);
nand U474 (N_474,In_6,In_631);
nor U475 (N_475,In_764,In_137);
or U476 (N_476,In_266,In_165);
or U477 (N_477,In_827,In_35);
or U478 (N_478,In_342,In_684);
and U479 (N_479,In_261,In_350);
or U480 (N_480,In_197,In_769);
and U481 (N_481,In_257,In_47);
nor U482 (N_482,In_202,In_85);
nand U483 (N_483,In_241,In_131);
nor U484 (N_484,In_411,In_836);
nor U485 (N_485,In_10,In_925);
nand U486 (N_486,In_455,In_249);
nor U487 (N_487,In_3,In_739);
nand U488 (N_488,In_834,In_62);
and U489 (N_489,In_698,In_331);
nor U490 (N_490,In_235,In_379);
or U491 (N_491,In_226,In_932);
nor U492 (N_492,In_508,In_696);
nor U493 (N_493,In_699,In_806);
or U494 (N_494,In_20,In_758);
and U495 (N_495,In_474,In_259);
and U496 (N_496,In_752,In_904);
or U497 (N_497,In_154,In_250);
and U498 (N_498,In_900,In_776);
nor U499 (N_499,In_216,In_439);
nor U500 (N_500,In_481,In_419);
and U501 (N_501,In_631,In_108);
and U502 (N_502,In_349,In_581);
and U503 (N_503,In_94,In_848);
nor U504 (N_504,In_14,In_881);
nand U505 (N_505,In_43,In_677);
and U506 (N_506,In_353,In_715);
nor U507 (N_507,In_330,In_3);
nor U508 (N_508,In_691,In_157);
nor U509 (N_509,In_862,In_166);
nor U510 (N_510,In_777,In_910);
or U511 (N_511,In_395,In_402);
or U512 (N_512,In_629,In_56);
or U513 (N_513,In_789,In_406);
xnor U514 (N_514,In_668,In_773);
nand U515 (N_515,In_158,In_291);
nand U516 (N_516,In_242,In_366);
and U517 (N_517,In_762,In_832);
or U518 (N_518,In_796,In_190);
and U519 (N_519,In_834,In_824);
or U520 (N_520,In_575,In_78);
or U521 (N_521,In_703,In_644);
nand U522 (N_522,In_896,In_941);
or U523 (N_523,In_369,In_278);
and U524 (N_524,In_148,In_55);
and U525 (N_525,In_314,In_838);
or U526 (N_526,In_623,In_927);
and U527 (N_527,In_252,In_358);
or U528 (N_528,In_283,In_655);
or U529 (N_529,In_180,In_620);
nand U530 (N_530,In_348,In_280);
nand U531 (N_531,In_97,In_762);
nand U532 (N_532,In_368,In_852);
nor U533 (N_533,In_618,In_183);
and U534 (N_534,In_943,In_21);
nand U535 (N_535,In_779,In_979);
and U536 (N_536,In_430,In_507);
and U537 (N_537,In_978,In_91);
nor U538 (N_538,In_285,In_70);
nor U539 (N_539,In_758,In_787);
and U540 (N_540,In_896,In_111);
nand U541 (N_541,In_795,In_878);
nand U542 (N_542,In_564,In_435);
nand U543 (N_543,In_764,In_196);
nand U544 (N_544,In_417,In_787);
and U545 (N_545,In_33,In_622);
or U546 (N_546,In_314,In_237);
nor U547 (N_547,In_293,In_206);
nor U548 (N_548,In_938,In_16);
nand U549 (N_549,In_449,In_222);
and U550 (N_550,In_173,In_454);
nand U551 (N_551,In_117,In_668);
and U552 (N_552,In_444,In_972);
nand U553 (N_553,In_945,In_330);
and U554 (N_554,In_627,In_643);
or U555 (N_555,In_997,In_326);
or U556 (N_556,In_442,In_886);
or U557 (N_557,In_977,In_255);
or U558 (N_558,In_846,In_669);
and U559 (N_559,In_435,In_464);
nor U560 (N_560,In_762,In_499);
nor U561 (N_561,In_336,In_255);
or U562 (N_562,In_355,In_379);
nor U563 (N_563,In_530,In_37);
nor U564 (N_564,In_918,In_973);
and U565 (N_565,In_2,In_853);
and U566 (N_566,In_71,In_937);
nor U567 (N_567,In_435,In_913);
nand U568 (N_568,In_738,In_169);
and U569 (N_569,In_143,In_875);
nor U570 (N_570,In_273,In_203);
or U571 (N_571,In_116,In_724);
nor U572 (N_572,In_16,In_942);
nand U573 (N_573,In_504,In_324);
nand U574 (N_574,In_805,In_297);
and U575 (N_575,In_860,In_958);
xor U576 (N_576,In_757,In_204);
nand U577 (N_577,In_542,In_83);
or U578 (N_578,In_274,In_812);
nand U579 (N_579,In_969,In_31);
nor U580 (N_580,In_500,In_164);
nand U581 (N_581,In_436,In_261);
or U582 (N_582,In_970,In_671);
and U583 (N_583,In_176,In_766);
nor U584 (N_584,In_828,In_833);
and U585 (N_585,In_959,In_246);
and U586 (N_586,In_830,In_44);
nand U587 (N_587,In_325,In_106);
and U588 (N_588,In_436,In_333);
or U589 (N_589,In_990,In_892);
or U590 (N_590,In_881,In_801);
or U591 (N_591,In_62,In_297);
and U592 (N_592,In_942,In_23);
nand U593 (N_593,In_688,In_452);
and U594 (N_594,In_149,In_371);
or U595 (N_595,In_811,In_206);
xnor U596 (N_596,In_511,In_661);
nor U597 (N_597,In_950,In_946);
nor U598 (N_598,In_487,In_837);
nand U599 (N_599,In_282,In_924);
nor U600 (N_600,In_810,In_352);
nand U601 (N_601,In_630,In_995);
or U602 (N_602,In_279,In_544);
nand U603 (N_603,In_46,In_253);
and U604 (N_604,In_773,In_677);
nor U605 (N_605,In_762,In_373);
or U606 (N_606,In_223,In_422);
and U607 (N_607,In_79,In_170);
nand U608 (N_608,In_41,In_471);
nor U609 (N_609,In_225,In_661);
nor U610 (N_610,In_458,In_794);
nand U611 (N_611,In_246,In_764);
or U612 (N_612,In_741,In_281);
nand U613 (N_613,In_533,In_114);
and U614 (N_614,In_812,In_855);
or U615 (N_615,In_866,In_185);
nand U616 (N_616,In_961,In_192);
nor U617 (N_617,In_274,In_418);
or U618 (N_618,In_938,In_127);
or U619 (N_619,In_796,In_801);
and U620 (N_620,In_527,In_178);
and U621 (N_621,In_804,In_865);
or U622 (N_622,In_332,In_336);
and U623 (N_623,In_91,In_15);
and U624 (N_624,In_557,In_838);
nand U625 (N_625,In_795,In_242);
and U626 (N_626,In_788,In_789);
nand U627 (N_627,In_171,In_150);
nand U628 (N_628,In_230,In_269);
nor U629 (N_629,In_825,In_775);
nand U630 (N_630,In_186,In_434);
nor U631 (N_631,In_893,In_595);
nor U632 (N_632,In_293,In_94);
and U633 (N_633,In_341,In_708);
nand U634 (N_634,In_339,In_65);
nand U635 (N_635,In_309,In_658);
and U636 (N_636,In_590,In_477);
and U637 (N_637,In_618,In_855);
nand U638 (N_638,In_398,In_829);
nor U639 (N_639,In_834,In_490);
nor U640 (N_640,In_774,In_292);
or U641 (N_641,In_418,In_255);
nor U642 (N_642,In_303,In_929);
nand U643 (N_643,In_428,In_839);
or U644 (N_644,In_750,In_753);
or U645 (N_645,In_554,In_497);
and U646 (N_646,In_150,In_817);
nand U647 (N_647,In_255,In_589);
nand U648 (N_648,In_151,In_524);
nand U649 (N_649,In_764,In_47);
nor U650 (N_650,In_953,In_137);
nand U651 (N_651,In_607,In_690);
nand U652 (N_652,In_103,In_964);
nor U653 (N_653,In_905,In_828);
nor U654 (N_654,In_474,In_678);
and U655 (N_655,In_476,In_133);
nand U656 (N_656,In_224,In_580);
nand U657 (N_657,In_594,In_595);
nand U658 (N_658,In_872,In_4);
nand U659 (N_659,In_152,In_213);
and U660 (N_660,In_450,In_433);
nand U661 (N_661,In_97,In_105);
or U662 (N_662,In_228,In_553);
xnor U663 (N_663,In_170,In_858);
and U664 (N_664,In_251,In_630);
and U665 (N_665,In_20,In_80);
xnor U666 (N_666,In_985,In_905);
and U667 (N_667,In_406,In_364);
or U668 (N_668,In_856,In_420);
and U669 (N_669,In_48,In_456);
or U670 (N_670,In_470,In_81);
nand U671 (N_671,In_672,In_290);
nand U672 (N_672,In_663,In_159);
or U673 (N_673,In_752,In_412);
nor U674 (N_674,In_287,In_291);
or U675 (N_675,In_683,In_693);
and U676 (N_676,In_358,In_199);
nand U677 (N_677,In_71,In_744);
nand U678 (N_678,In_513,In_657);
and U679 (N_679,In_300,In_5);
nor U680 (N_680,In_505,In_387);
and U681 (N_681,In_84,In_902);
and U682 (N_682,In_186,In_190);
xnor U683 (N_683,In_575,In_494);
and U684 (N_684,In_514,In_507);
or U685 (N_685,In_187,In_359);
or U686 (N_686,In_783,In_86);
nand U687 (N_687,In_295,In_46);
nand U688 (N_688,In_583,In_549);
and U689 (N_689,In_191,In_106);
and U690 (N_690,In_11,In_41);
nor U691 (N_691,In_209,In_434);
and U692 (N_692,In_367,In_234);
nor U693 (N_693,In_482,In_399);
xnor U694 (N_694,In_581,In_215);
nand U695 (N_695,In_969,In_90);
nand U696 (N_696,In_243,In_196);
nand U697 (N_697,In_893,In_996);
nor U698 (N_698,In_812,In_999);
nor U699 (N_699,In_131,In_804);
and U700 (N_700,In_594,In_530);
or U701 (N_701,In_312,In_148);
and U702 (N_702,In_817,In_718);
and U703 (N_703,In_112,In_528);
and U704 (N_704,In_994,In_256);
nand U705 (N_705,In_100,In_886);
and U706 (N_706,In_556,In_219);
nand U707 (N_707,In_69,In_75);
and U708 (N_708,In_301,In_351);
and U709 (N_709,In_574,In_56);
and U710 (N_710,In_505,In_130);
nand U711 (N_711,In_464,In_439);
or U712 (N_712,In_88,In_771);
and U713 (N_713,In_309,In_70);
nor U714 (N_714,In_653,In_42);
or U715 (N_715,In_426,In_18);
or U716 (N_716,In_601,In_575);
nor U717 (N_717,In_665,In_149);
nor U718 (N_718,In_700,In_181);
nor U719 (N_719,In_44,In_20);
nand U720 (N_720,In_866,In_444);
nand U721 (N_721,In_116,In_268);
or U722 (N_722,In_172,In_546);
or U723 (N_723,In_783,In_785);
nor U724 (N_724,In_493,In_180);
xnor U725 (N_725,In_526,In_604);
or U726 (N_726,In_897,In_412);
or U727 (N_727,In_893,In_990);
or U728 (N_728,In_992,In_590);
nand U729 (N_729,In_124,In_262);
and U730 (N_730,In_818,In_968);
or U731 (N_731,In_776,In_179);
and U732 (N_732,In_714,In_915);
or U733 (N_733,In_939,In_393);
or U734 (N_734,In_592,In_623);
or U735 (N_735,In_230,In_603);
nor U736 (N_736,In_431,In_962);
or U737 (N_737,In_998,In_972);
and U738 (N_738,In_255,In_552);
and U739 (N_739,In_640,In_836);
nor U740 (N_740,In_781,In_72);
or U741 (N_741,In_71,In_799);
nor U742 (N_742,In_763,In_947);
nor U743 (N_743,In_979,In_526);
xor U744 (N_744,In_481,In_563);
xnor U745 (N_745,In_173,In_726);
nor U746 (N_746,In_974,In_42);
nand U747 (N_747,In_962,In_999);
and U748 (N_748,In_105,In_197);
nor U749 (N_749,In_669,In_649);
nor U750 (N_750,In_981,In_780);
nand U751 (N_751,In_839,In_777);
or U752 (N_752,In_386,In_749);
and U753 (N_753,In_513,In_19);
or U754 (N_754,In_924,In_598);
or U755 (N_755,In_716,In_148);
and U756 (N_756,In_17,In_827);
nor U757 (N_757,In_167,In_256);
and U758 (N_758,In_734,In_963);
or U759 (N_759,In_422,In_863);
nand U760 (N_760,In_130,In_888);
or U761 (N_761,In_115,In_896);
or U762 (N_762,In_667,In_0);
nand U763 (N_763,In_329,In_77);
and U764 (N_764,In_725,In_595);
or U765 (N_765,In_519,In_560);
or U766 (N_766,In_470,In_593);
or U767 (N_767,In_895,In_856);
and U768 (N_768,In_518,In_289);
and U769 (N_769,In_817,In_41);
and U770 (N_770,In_383,In_237);
and U771 (N_771,In_133,In_490);
or U772 (N_772,In_50,In_203);
nand U773 (N_773,In_807,In_270);
or U774 (N_774,In_855,In_621);
or U775 (N_775,In_227,In_418);
nor U776 (N_776,In_378,In_465);
nand U777 (N_777,In_622,In_710);
nand U778 (N_778,In_73,In_49);
nor U779 (N_779,In_944,In_977);
or U780 (N_780,In_551,In_51);
or U781 (N_781,In_518,In_50);
and U782 (N_782,In_608,In_210);
or U783 (N_783,In_836,In_620);
and U784 (N_784,In_290,In_643);
or U785 (N_785,In_417,In_952);
and U786 (N_786,In_581,In_676);
nor U787 (N_787,In_359,In_736);
or U788 (N_788,In_772,In_123);
nand U789 (N_789,In_784,In_134);
nand U790 (N_790,In_499,In_58);
and U791 (N_791,In_941,In_690);
and U792 (N_792,In_443,In_138);
nand U793 (N_793,In_200,In_968);
or U794 (N_794,In_82,In_83);
nand U795 (N_795,In_699,In_886);
and U796 (N_796,In_280,In_362);
or U797 (N_797,In_988,In_885);
and U798 (N_798,In_608,In_350);
or U799 (N_799,In_314,In_520);
nand U800 (N_800,In_91,In_333);
and U801 (N_801,In_306,In_637);
nor U802 (N_802,In_859,In_727);
nand U803 (N_803,In_832,In_964);
and U804 (N_804,In_423,In_786);
nand U805 (N_805,In_971,In_53);
or U806 (N_806,In_889,In_331);
nor U807 (N_807,In_440,In_992);
nand U808 (N_808,In_163,In_507);
nand U809 (N_809,In_990,In_391);
nor U810 (N_810,In_739,In_265);
and U811 (N_811,In_598,In_835);
and U812 (N_812,In_108,In_505);
nand U813 (N_813,In_634,In_777);
or U814 (N_814,In_104,In_455);
and U815 (N_815,In_290,In_694);
or U816 (N_816,In_520,In_666);
or U817 (N_817,In_753,In_995);
xnor U818 (N_818,In_320,In_281);
nand U819 (N_819,In_597,In_745);
nor U820 (N_820,In_228,In_965);
nand U821 (N_821,In_35,In_691);
and U822 (N_822,In_105,In_677);
xor U823 (N_823,In_485,In_171);
or U824 (N_824,In_144,In_264);
nand U825 (N_825,In_847,In_403);
nand U826 (N_826,In_783,In_603);
and U827 (N_827,In_40,In_455);
nand U828 (N_828,In_271,In_905);
nand U829 (N_829,In_892,In_42);
nor U830 (N_830,In_808,In_614);
or U831 (N_831,In_820,In_34);
nand U832 (N_832,In_993,In_280);
xor U833 (N_833,In_784,In_612);
and U834 (N_834,In_502,In_418);
or U835 (N_835,In_487,In_966);
nor U836 (N_836,In_806,In_222);
nand U837 (N_837,In_708,In_956);
and U838 (N_838,In_615,In_542);
or U839 (N_839,In_22,In_689);
xor U840 (N_840,In_534,In_658);
nor U841 (N_841,In_114,In_429);
and U842 (N_842,In_854,In_189);
nor U843 (N_843,In_343,In_500);
and U844 (N_844,In_131,In_520);
nor U845 (N_845,In_718,In_51);
and U846 (N_846,In_63,In_161);
nor U847 (N_847,In_182,In_631);
and U848 (N_848,In_727,In_841);
and U849 (N_849,In_831,In_929);
nand U850 (N_850,In_552,In_401);
nand U851 (N_851,In_903,In_689);
or U852 (N_852,In_780,In_543);
nor U853 (N_853,In_225,In_984);
and U854 (N_854,In_191,In_315);
or U855 (N_855,In_302,In_253);
and U856 (N_856,In_539,In_218);
nand U857 (N_857,In_811,In_28);
and U858 (N_858,In_40,In_44);
nand U859 (N_859,In_320,In_845);
or U860 (N_860,In_841,In_718);
or U861 (N_861,In_714,In_993);
nor U862 (N_862,In_618,In_818);
nor U863 (N_863,In_782,In_541);
nor U864 (N_864,In_817,In_833);
or U865 (N_865,In_906,In_374);
and U866 (N_866,In_419,In_980);
nand U867 (N_867,In_782,In_998);
or U868 (N_868,In_76,In_571);
and U869 (N_869,In_285,In_807);
nor U870 (N_870,In_598,In_728);
nand U871 (N_871,In_112,In_49);
or U872 (N_872,In_959,In_473);
nand U873 (N_873,In_123,In_68);
and U874 (N_874,In_983,In_121);
xor U875 (N_875,In_175,In_860);
or U876 (N_876,In_293,In_498);
and U877 (N_877,In_997,In_179);
nor U878 (N_878,In_602,In_948);
or U879 (N_879,In_380,In_489);
and U880 (N_880,In_764,In_916);
nand U881 (N_881,In_335,In_547);
nand U882 (N_882,In_471,In_379);
xor U883 (N_883,In_393,In_337);
nand U884 (N_884,In_522,In_920);
nand U885 (N_885,In_945,In_508);
or U886 (N_886,In_424,In_866);
and U887 (N_887,In_363,In_382);
or U888 (N_888,In_74,In_695);
or U889 (N_889,In_468,In_419);
and U890 (N_890,In_38,In_48);
or U891 (N_891,In_974,In_128);
and U892 (N_892,In_960,In_72);
nor U893 (N_893,In_18,In_724);
nor U894 (N_894,In_846,In_38);
or U895 (N_895,In_133,In_46);
and U896 (N_896,In_965,In_171);
and U897 (N_897,In_923,In_185);
xnor U898 (N_898,In_443,In_968);
and U899 (N_899,In_619,In_206);
nand U900 (N_900,In_30,In_697);
or U901 (N_901,In_474,In_4);
or U902 (N_902,In_741,In_802);
xnor U903 (N_903,In_797,In_337);
nand U904 (N_904,In_530,In_953);
and U905 (N_905,In_397,In_809);
or U906 (N_906,In_846,In_607);
nor U907 (N_907,In_107,In_755);
or U908 (N_908,In_230,In_193);
and U909 (N_909,In_838,In_879);
nand U910 (N_910,In_589,In_939);
and U911 (N_911,In_878,In_297);
or U912 (N_912,In_576,In_432);
or U913 (N_913,In_94,In_896);
nand U914 (N_914,In_453,In_357);
xor U915 (N_915,In_989,In_861);
nor U916 (N_916,In_371,In_716);
xor U917 (N_917,In_176,In_497);
nor U918 (N_918,In_558,In_140);
and U919 (N_919,In_655,In_582);
nand U920 (N_920,In_280,In_947);
and U921 (N_921,In_689,In_310);
nor U922 (N_922,In_210,In_495);
nand U923 (N_923,In_800,In_276);
nand U924 (N_924,In_375,In_703);
and U925 (N_925,In_665,In_475);
and U926 (N_926,In_247,In_49);
nand U927 (N_927,In_525,In_442);
and U928 (N_928,In_930,In_655);
or U929 (N_929,In_954,In_369);
and U930 (N_930,In_879,In_750);
nand U931 (N_931,In_22,In_490);
or U932 (N_932,In_472,In_624);
or U933 (N_933,In_930,In_994);
nand U934 (N_934,In_413,In_245);
and U935 (N_935,In_697,In_50);
nand U936 (N_936,In_240,In_571);
and U937 (N_937,In_272,In_937);
and U938 (N_938,In_860,In_742);
nand U939 (N_939,In_292,In_634);
nand U940 (N_940,In_435,In_416);
nand U941 (N_941,In_924,In_45);
and U942 (N_942,In_783,In_188);
and U943 (N_943,In_233,In_113);
or U944 (N_944,In_353,In_647);
nor U945 (N_945,In_801,In_516);
nand U946 (N_946,In_260,In_140);
and U947 (N_947,In_132,In_516);
nor U948 (N_948,In_227,In_510);
nor U949 (N_949,In_893,In_184);
nand U950 (N_950,In_161,In_762);
nor U951 (N_951,In_751,In_979);
nor U952 (N_952,In_36,In_988);
and U953 (N_953,In_482,In_437);
and U954 (N_954,In_621,In_771);
nand U955 (N_955,In_351,In_938);
or U956 (N_956,In_219,In_766);
nand U957 (N_957,In_158,In_908);
nand U958 (N_958,In_977,In_19);
nand U959 (N_959,In_537,In_954);
nor U960 (N_960,In_972,In_269);
nor U961 (N_961,In_622,In_391);
and U962 (N_962,In_566,In_66);
or U963 (N_963,In_575,In_444);
nor U964 (N_964,In_469,In_369);
and U965 (N_965,In_184,In_219);
and U966 (N_966,In_60,In_213);
or U967 (N_967,In_436,In_362);
nand U968 (N_968,In_221,In_800);
and U969 (N_969,In_746,In_24);
and U970 (N_970,In_925,In_87);
nand U971 (N_971,In_94,In_262);
and U972 (N_972,In_580,In_407);
or U973 (N_973,In_512,In_489);
or U974 (N_974,In_191,In_652);
or U975 (N_975,In_30,In_59);
and U976 (N_976,In_333,In_881);
or U977 (N_977,In_746,In_312);
nand U978 (N_978,In_890,In_816);
nand U979 (N_979,In_198,In_919);
or U980 (N_980,In_607,In_283);
nor U981 (N_981,In_819,In_13);
nor U982 (N_982,In_917,In_439);
nor U983 (N_983,In_387,In_820);
nand U984 (N_984,In_566,In_856);
nor U985 (N_985,In_909,In_391);
or U986 (N_986,In_268,In_300);
nor U987 (N_987,In_76,In_215);
or U988 (N_988,In_954,In_29);
nor U989 (N_989,In_374,In_99);
or U990 (N_990,In_893,In_301);
or U991 (N_991,In_722,In_451);
nand U992 (N_992,In_597,In_696);
and U993 (N_993,In_667,In_306);
nand U994 (N_994,In_372,In_565);
nor U995 (N_995,In_765,In_105);
nor U996 (N_996,In_396,In_426);
and U997 (N_997,In_921,In_875);
and U998 (N_998,In_930,In_686);
and U999 (N_999,In_337,In_943);
nand U1000 (N_1000,In_320,In_39);
nor U1001 (N_1001,In_854,In_28);
nor U1002 (N_1002,In_217,In_519);
and U1003 (N_1003,In_189,In_638);
nand U1004 (N_1004,In_834,In_913);
or U1005 (N_1005,In_351,In_972);
nor U1006 (N_1006,In_417,In_440);
and U1007 (N_1007,In_203,In_265);
or U1008 (N_1008,In_828,In_807);
or U1009 (N_1009,In_49,In_829);
and U1010 (N_1010,In_371,In_918);
and U1011 (N_1011,In_514,In_656);
and U1012 (N_1012,In_333,In_194);
nor U1013 (N_1013,In_349,In_390);
or U1014 (N_1014,In_538,In_944);
and U1015 (N_1015,In_716,In_418);
nor U1016 (N_1016,In_474,In_735);
nor U1017 (N_1017,In_614,In_629);
nor U1018 (N_1018,In_429,In_988);
and U1019 (N_1019,In_944,In_834);
and U1020 (N_1020,In_335,In_2);
or U1021 (N_1021,In_275,In_30);
xor U1022 (N_1022,In_669,In_880);
nor U1023 (N_1023,In_161,In_248);
nand U1024 (N_1024,In_602,In_375);
and U1025 (N_1025,In_892,In_772);
and U1026 (N_1026,In_147,In_727);
nor U1027 (N_1027,In_219,In_610);
nor U1028 (N_1028,In_562,In_712);
nor U1029 (N_1029,In_839,In_128);
nand U1030 (N_1030,In_851,In_191);
nor U1031 (N_1031,In_870,In_81);
nor U1032 (N_1032,In_126,In_640);
and U1033 (N_1033,In_133,In_906);
nand U1034 (N_1034,In_857,In_276);
or U1035 (N_1035,In_726,In_436);
and U1036 (N_1036,In_62,In_377);
or U1037 (N_1037,In_58,In_311);
and U1038 (N_1038,In_745,In_882);
nand U1039 (N_1039,In_824,In_120);
nor U1040 (N_1040,In_264,In_460);
nor U1041 (N_1041,In_458,In_611);
or U1042 (N_1042,In_448,In_552);
and U1043 (N_1043,In_33,In_804);
nand U1044 (N_1044,In_279,In_269);
nor U1045 (N_1045,In_700,In_663);
and U1046 (N_1046,In_387,In_70);
and U1047 (N_1047,In_655,In_519);
and U1048 (N_1048,In_998,In_221);
and U1049 (N_1049,In_424,In_388);
and U1050 (N_1050,In_255,In_355);
nand U1051 (N_1051,In_703,In_38);
nor U1052 (N_1052,In_948,In_381);
nand U1053 (N_1053,In_611,In_7);
nor U1054 (N_1054,In_462,In_362);
or U1055 (N_1055,In_970,In_704);
nand U1056 (N_1056,In_481,In_336);
or U1057 (N_1057,In_526,In_424);
or U1058 (N_1058,In_942,In_105);
and U1059 (N_1059,In_263,In_8);
or U1060 (N_1060,In_842,In_60);
and U1061 (N_1061,In_729,In_28);
nor U1062 (N_1062,In_584,In_595);
or U1063 (N_1063,In_202,In_613);
nor U1064 (N_1064,In_326,In_356);
nor U1065 (N_1065,In_506,In_15);
or U1066 (N_1066,In_745,In_708);
xor U1067 (N_1067,In_24,In_233);
nand U1068 (N_1068,In_404,In_445);
nand U1069 (N_1069,In_381,In_300);
or U1070 (N_1070,In_642,In_701);
and U1071 (N_1071,In_251,In_383);
nand U1072 (N_1072,In_722,In_155);
and U1073 (N_1073,In_527,In_5);
nor U1074 (N_1074,In_770,In_725);
and U1075 (N_1075,In_757,In_939);
nand U1076 (N_1076,In_786,In_373);
nand U1077 (N_1077,In_647,In_272);
nor U1078 (N_1078,In_879,In_505);
and U1079 (N_1079,In_136,In_798);
or U1080 (N_1080,In_922,In_892);
nor U1081 (N_1081,In_406,In_163);
and U1082 (N_1082,In_579,In_810);
nor U1083 (N_1083,In_674,In_205);
and U1084 (N_1084,In_859,In_220);
or U1085 (N_1085,In_198,In_527);
nand U1086 (N_1086,In_568,In_744);
and U1087 (N_1087,In_702,In_984);
or U1088 (N_1088,In_382,In_20);
and U1089 (N_1089,In_855,In_6);
and U1090 (N_1090,In_214,In_371);
nand U1091 (N_1091,In_674,In_595);
nand U1092 (N_1092,In_150,In_220);
or U1093 (N_1093,In_466,In_10);
and U1094 (N_1094,In_891,In_466);
nor U1095 (N_1095,In_217,In_548);
and U1096 (N_1096,In_375,In_338);
nor U1097 (N_1097,In_283,In_516);
or U1098 (N_1098,In_298,In_613);
nor U1099 (N_1099,In_389,In_454);
or U1100 (N_1100,In_574,In_960);
and U1101 (N_1101,In_992,In_756);
and U1102 (N_1102,In_940,In_336);
nor U1103 (N_1103,In_598,In_268);
and U1104 (N_1104,In_871,In_759);
nand U1105 (N_1105,In_997,In_990);
and U1106 (N_1106,In_613,In_619);
or U1107 (N_1107,In_665,In_404);
nand U1108 (N_1108,In_715,In_146);
or U1109 (N_1109,In_8,In_433);
or U1110 (N_1110,In_61,In_552);
nand U1111 (N_1111,In_928,In_325);
and U1112 (N_1112,In_128,In_758);
nor U1113 (N_1113,In_761,In_59);
nand U1114 (N_1114,In_239,In_964);
nand U1115 (N_1115,In_620,In_219);
nor U1116 (N_1116,In_364,In_694);
and U1117 (N_1117,In_289,In_357);
or U1118 (N_1118,In_910,In_875);
nand U1119 (N_1119,In_31,In_777);
and U1120 (N_1120,In_908,In_335);
or U1121 (N_1121,In_756,In_241);
and U1122 (N_1122,In_116,In_255);
or U1123 (N_1123,In_7,In_984);
nand U1124 (N_1124,In_356,In_669);
nor U1125 (N_1125,In_901,In_221);
nand U1126 (N_1126,In_597,In_823);
nand U1127 (N_1127,In_797,In_53);
nor U1128 (N_1128,In_382,In_595);
or U1129 (N_1129,In_433,In_18);
xor U1130 (N_1130,In_729,In_592);
nor U1131 (N_1131,In_486,In_372);
nor U1132 (N_1132,In_298,In_296);
and U1133 (N_1133,In_401,In_151);
nand U1134 (N_1134,In_633,In_14);
xnor U1135 (N_1135,In_75,In_507);
nor U1136 (N_1136,In_487,In_984);
xnor U1137 (N_1137,In_541,In_411);
nor U1138 (N_1138,In_558,In_50);
or U1139 (N_1139,In_202,In_837);
or U1140 (N_1140,In_716,In_389);
nor U1141 (N_1141,In_194,In_867);
and U1142 (N_1142,In_301,In_775);
and U1143 (N_1143,In_613,In_730);
nand U1144 (N_1144,In_100,In_884);
or U1145 (N_1145,In_498,In_660);
and U1146 (N_1146,In_142,In_729);
or U1147 (N_1147,In_407,In_149);
nor U1148 (N_1148,In_930,In_668);
nor U1149 (N_1149,In_695,In_209);
nor U1150 (N_1150,In_537,In_6);
or U1151 (N_1151,In_832,In_803);
nor U1152 (N_1152,In_476,In_552);
and U1153 (N_1153,In_894,In_636);
and U1154 (N_1154,In_604,In_323);
nor U1155 (N_1155,In_208,In_423);
or U1156 (N_1156,In_936,In_95);
nand U1157 (N_1157,In_333,In_466);
nor U1158 (N_1158,In_522,In_992);
and U1159 (N_1159,In_637,In_585);
and U1160 (N_1160,In_513,In_979);
xor U1161 (N_1161,In_203,In_83);
nand U1162 (N_1162,In_71,In_266);
nand U1163 (N_1163,In_172,In_738);
and U1164 (N_1164,In_714,In_27);
and U1165 (N_1165,In_863,In_692);
or U1166 (N_1166,In_813,In_311);
xnor U1167 (N_1167,In_447,In_690);
nor U1168 (N_1168,In_497,In_527);
or U1169 (N_1169,In_663,In_520);
and U1170 (N_1170,In_705,In_509);
or U1171 (N_1171,In_475,In_87);
and U1172 (N_1172,In_868,In_245);
or U1173 (N_1173,In_884,In_321);
or U1174 (N_1174,In_30,In_522);
nand U1175 (N_1175,In_517,In_55);
or U1176 (N_1176,In_145,In_919);
nor U1177 (N_1177,In_801,In_770);
nor U1178 (N_1178,In_62,In_336);
or U1179 (N_1179,In_22,In_32);
nor U1180 (N_1180,In_453,In_168);
and U1181 (N_1181,In_892,In_534);
xor U1182 (N_1182,In_664,In_876);
or U1183 (N_1183,In_98,In_261);
nor U1184 (N_1184,In_710,In_443);
or U1185 (N_1185,In_359,In_934);
or U1186 (N_1186,In_488,In_98);
nor U1187 (N_1187,In_129,In_876);
nor U1188 (N_1188,In_797,In_545);
or U1189 (N_1189,In_364,In_645);
xnor U1190 (N_1190,In_954,In_348);
nor U1191 (N_1191,In_152,In_851);
nand U1192 (N_1192,In_16,In_601);
and U1193 (N_1193,In_322,In_701);
nand U1194 (N_1194,In_748,In_218);
nor U1195 (N_1195,In_49,In_529);
nor U1196 (N_1196,In_67,In_518);
and U1197 (N_1197,In_405,In_872);
or U1198 (N_1198,In_774,In_97);
nand U1199 (N_1199,In_70,In_315);
or U1200 (N_1200,In_195,In_54);
and U1201 (N_1201,In_942,In_543);
or U1202 (N_1202,In_534,In_191);
nor U1203 (N_1203,In_428,In_80);
and U1204 (N_1204,In_816,In_154);
or U1205 (N_1205,In_367,In_228);
nand U1206 (N_1206,In_276,In_70);
and U1207 (N_1207,In_322,In_588);
or U1208 (N_1208,In_302,In_710);
and U1209 (N_1209,In_808,In_193);
nand U1210 (N_1210,In_219,In_325);
or U1211 (N_1211,In_342,In_66);
nor U1212 (N_1212,In_515,In_198);
or U1213 (N_1213,In_60,In_71);
nor U1214 (N_1214,In_33,In_283);
and U1215 (N_1215,In_729,In_672);
nor U1216 (N_1216,In_36,In_131);
nand U1217 (N_1217,In_583,In_904);
nand U1218 (N_1218,In_703,In_856);
nor U1219 (N_1219,In_378,In_643);
or U1220 (N_1220,In_655,In_249);
nand U1221 (N_1221,In_629,In_623);
and U1222 (N_1222,In_18,In_950);
xnor U1223 (N_1223,In_524,In_107);
nand U1224 (N_1224,In_837,In_375);
or U1225 (N_1225,In_33,In_513);
and U1226 (N_1226,In_451,In_270);
nor U1227 (N_1227,In_338,In_256);
nand U1228 (N_1228,In_871,In_327);
or U1229 (N_1229,In_111,In_952);
or U1230 (N_1230,In_285,In_289);
or U1231 (N_1231,In_638,In_770);
and U1232 (N_1232,In_327,In_379);
nand U1233 (N_1233,In_355,In_73);
nand U1234 (N_1234,In_728,In_212);
and U1235 (N_1235,In_604,In_263);
nand U1236 (N_1236,In_247,In_770);
nand U1237 (N_1237,In_404,In_482);
nor U1238 (N_1238,In_955,In_394);
nand U1239 (N_1239,In_286,In_832);
and U1240 (N_1240,In_475,In_241);
and U1241 (N_1241,In_697,In_886);
or U1242 (N_1242,In_129,In_476);
or U1243 (N_1243,In_865,In_174);
or U1244 (N_1244,In_269,In_855);
nand U1245 (N_1245,In_222,In_310);
nand U1246 (N_1246,In_22,In_715);
and U1247 (N_1247,In_423,In_141);
nand U1248 (N_1248,In_546,In_13);
and U1249 (N_1249,In_61,In_620);
or U1250 (N_1250,In_234,In_726);
or U1251 (N_1251,In_527,In_181);
nor U1252 (N_1252,In_135,In_232);
nor U1253 (N_1253,In_804,In_443);
nor U1254 (N_1254,In_696,In_328);
xor U1255 (N_1255,In_783,In_113);
nor U1256 (N_1256,In_545,In_612);
or U1257 (N_1257,In_189,In_646);
nor U1258 (N_1258,In_232,In_645);
nand U1259 (N_1259,In_256,In_739);
nor U1260 (N_1260,In_535,In_766);
nand U1261 (N_1261,In_670,In_796);
nor U1262 (N_1262,In_842,In_930);
nor U1263 (N_1263,In_377,In_532);
or U1264 (N_1264,In_930,In_484);
nor U1265 (N_1265,In_153,In_58);
nand U1266 (N_1266,In_431,In_618);
nand U1267 (N_1267,In_855,In_820);
nand U1268 (N_1268,In_488,In_683);
and U1269 (N_1269,In_472,In_238);
nor U1270 (N_1270,In_298,In_426);
nand U1271 (N_1271,In_990,In_822);
and U1272 (N_1272,In_533,In_124);
or U1273 (N_1273,In_65,In_473);
or U1274 (N_1274,In_962,In_26);
and U1275 (N_1275,In_165,In_281);
nor U1276 (N_1276,In_907,In_33);
nand U1277 (N_1277,In_616,In_913);
and U1278 (N_1278,In_606,In_593);
xnor U1279 (N_1279,In_488,In_432);
or U1280 (N_1280,In_216,In_64);
or U1281 (N_1281,In_544,In_686);
nor U1282 (N_1282,In_255,In_976);
and U1283 (N_1283,In_447,In_643);
and U1284 (N_1284,In_802,In_889);
nor U1285 (N_1285,In_376,In_915);
or U1286 (N_1286,In_937,In_607);
nand U1287 (N_1287,In_559,In_196);
or U1288 (N_1288,In_240,In_634);
nor U1289 (N_1289,In_340,In_285);
nand U1290 (N_1290,In_913,In_275);
nor U1291 (N_1291,In_91,In_916);
or U1292 (N_1292,In_269,In_976);
or U1293 (N_1293,In_193,In_651);
or U1294 (N_1294,In_456,In_936);
xnor U1295 (N_1295,In_605,In_524);
nand U1296 (N_1296,In_674,In_574);
nand U1297 (N_1297,In_657,In_686);
nor U1298 (N_1298,In_24,In_881);
nor U1299 (N_1299,In_762,In_506);
nor U1300 (N_1300,In_503,In_116);
and U1301 (N_1301,In_349,In_499);
nand U1302 (N_1302,In_35,In_310);
nor U1303 (N_1303,In_596,In_178);
and U1304 (N_1304,In_384,In_357);
and U1305 (N_1305,In_915,In_993);
and U1306 (N_1306,In_747,In_818);
nand U1307 (N_1307,In_905,In_377);
or U1308 (N_1308,In_899,In_492);
and U1309 (N_1309,In_493,In_30);
nor U1310 (N_1310,In_658,In_516);
nor U1311 (N_1311,In_516,In_491);
nand U1312 (N_1312,In_636,In_294);
xor U1313 (N_1313,In_255,In_41);
or U1314 (N_1314,In_454,In_705);
and U1315 (N_1315,In_525,In_234);
or U1316 (N_1316,In_806,In_150);
nor U1317 (N_1317,In_793,In_31);
or U1318 (N_1318,In_823,In_248);
nor U1319 (N_1319,In_316,In_905);
nand U1320 (N_1320,In_738,In_236);
or U1321 (N_1321,In_384,In_1);
nand U1322 (N_1322,In_262,In_163);
nor U1323 (N_1323,In_337,In_786);
nor U1324 (N_1324,In_454,In_953);
and U1325 (N_1325,In_681,In_679);
and U1326 (N_1326,In_35,In_895);
and U1327 (N_1327,In_529,In_838);
nor U1328 (N_1328,In_796,In_422);
and U1329 (N_1329,In_850,In_92);
nor U1330 (N_1330,In_988,In_51);
nand U1331 (N_1331,In_110,In_489);
nor U1332 (N_1332,In_340,In_490);
or U1333 (N_1333,In_98,In_571);
or U1334 (N_1334,In_506,In_825);
and U1335 (N_1335,In_447,In_502);
xnor U1336 (N_1336,In_392,In_588);
nand U1337 (N_1337,In_331,In_855);
nor U1338 (N_1338,In_26,In_263);
or U1339 (N_1339,In_21,In_625);
nand U1340 (N_1340,In_420,In_925);
and U1341 (N_1341,In_869,In_732);
and U1342 (N_1342,In_835,In_933);
or U1343 (N_1343,In_526,In_605);
and U1344 (N_1344,In_978,In_485);
or U1345 (N_1345,In_117,In_895);
nand U1346 (N_1346,In_269,In_721);
or U1347 (N_1347,In_880,In_705);
nor U1348 (N_1348,In_598,In_269);
or U1349 (N_1349,In_546,In_603);
and U1350 (N_1350,In_859,In_110);
and U1351 (N_1351,In_974,In_697);
or U1352 (N_1352,In_672,In_53);
nor U1353 (N_1353,In_450,In_752);
and U1354 (N_1354,In_959,In_223);
nand U1355 (N_1355,In_857,In_523);
or U1356 (N_1356,In_912,In_742);
nor U1357 (N_1357,In_508,In_338);
nand U1358 (N_1358,In_739,In_131);
nand U1359 (N_1359,In_128,In_368);
or U1360 (N_1360,In_419,In_926);
nor U1361 (N_1361,In_501,In_341);
xnor U1362 (N_1362,In_124,In_156);
and U1363 (N_1363,In_862,In_500);
nor U1364 (N_1364,In_657,In_269);
nor U1365 (N_1365,In_365,In_394);
nand U1366 (N_1366,In_149,In_718);
or U1367 (N_1367,In_735,In_841);
nand U1368 (N_1368,In_627,In_307);
or U1369 (N_1369,In_985,In_959);
and U1370 (N_1370,In_522,In_490);
nor U1371 (N_1371,In_680,In_455);
nor U1372 (N_1372,In_113,In_436);
and U1373 (N_1373,In_673,In_412);
nor U1374 (N_1374,In_750,In_898);
nand U1375 (N_1375,In_812,In_539);
nand U1376 (N_1376,In_34,In_748);
nand U1377 (N_1377,In_903,In_525);
or U1378 (N_1378,In_295,In_840);
nand U1379 (N_1379,In_866,In_751);
or U1380 (N_1380,In_660,In_606);
or U1381 (N_1381,In_791,In_103);
xor U1382 (N_1382,In_352,In_50);
or U1383 (N_1383,In_489,In_481);
and U1384 (N_1384,In_795,In_98);
or U1385 (N_1385,In_688,In_664);
nor U1386 (N_1386,In_25,In_169);
nor U1387 (N_1387,In_571,In_858);
nand U1388 (N_1388,In_25,In_644);
nand U1389 (N_1389,In_301,In_93);
or U1390 (N_1390,In_408,In_581);
nor U1391 (N_1391,In_385,In_43);
nor U1392 (N_1392,In_784,In_727);
nor U1393 (N_1393,In_825,In_373);
nand U1394 (N_1394,In_804,In_945);
nand U1395 (N_1395,In_540,In_517);
nor U1396 (N_1396,In_718,In_408);
or U1397 (N_1397,In_306,In_180);
nor U1398 (N_1398,In_952,In_558);
or U1399 (N_1399,In_948,In_212);
and U1400 (N_1400,In_671,In_518);
or U1401 (N_1401,In_193,In_576);
or U1402 (N_1402,In_714,In_603);
and U1403 (N_1403,In_994,In_44);
or U1404 (N_1404,In_948,In_350);
nor U1405 (N_1405,In_133,In_256);
nor U1406 (N_1406,In_857,In_433);
xor U1407 (N_1407,In_724,In_757);
nor U1408 (N_1408,In_967,In_352);
nand U1409 (N_1409,In_958,In_57);
nor U1410 (N_1410,In_743,In_944);
or U1411 (N_1411,In_174,In_748);
nand U1412 (N_1412,In_971,In_758);
nand U1413 (N_1413,In_171,In_999);
or U1414 (N_1414,In_775,In_397);
nor U1415 (N_1415,In_46,In_923);
nor U1416 (N_1416,In_737,In_710);
and U1417 (N_1417,In_523,In_781);
nor U1418 (N_1418,In_432,In_517);
nand U1419 (N_1419,In_859,In_342);
and U1420 (N_1420,In_363,In_75);
nor U1421 (N_1421,In_663,In_580);
nor U1422 (N_1422,In_56,In_898);
nor U1423 (N_1423,In_334,In_232);
nand U1424 (N_1424,In_615,In_618);
xnor U1425 (N_1425,In_938,In_651);
and U1426 (N_1426,In_158,In_776);
and U1427 (N_1427,In_523,In_509);
nor U1428 (N_1428,In_974,In_364);
or U1429 (N_1429,In_415,In_756);
or U1430 (N_1430,In_152,In_531);
nand U1431 (N_1431,In_623,In_868);
and U1432 (N_1432,In_752,In_552);
and U1433 (N_1433,In_765,In_758);
nor U1434 (N_1434,In_892,In_626);
or U1435 (N_1435,In_370,In_931);
and U1436 (N_1436,In_285,In_79);
nor U1437 (N_1437,In_280,In_568);
nor U1438 (N_1438,In_816,In_507);
or U1439 (N_1439,In_462,In_6);
and U1440 (N_1440,In_701,In_804);
or U1441 (N_1441,In_38,In_603);
and U1442 (N_1442,In_362,In_760);
or U1443 (N_1443,In_968,In_807);
and U1444 (N_1444,In_115,In_811);
nor U1445 (N_1445,In_977,In_153);
nand U1446 (N_1446,In_22,In_306);
nor U1447 (N_1447,In_290,In_59);
nand U1448 (N_1448,In_954,In_874);
nor U1449 (N_1449,In_869,In_53);
nor U1450 (N_1450,In_131,In_437);
nor U1451 (N_1451,In_556,In_373);
or U1452 (N_1452,In_752,In_21);
nand U1453 (N_1453,In_378,In_66);
nor U1454 (N_1454,In_195,In_945);
nand U1455 (N_1455,In_298,In_565);
and U1456 (N_1456,In_987,In_465);
or U1457 (N_1457,In_682,In_300);
or U1458 (N_1458,In_17,In_786);
nor U1459 (N_1459,In_739,In_491);
nor U1460 (N_1460,In_848,In_359);
nor U1461 (N_1461,In_173,In_382);
or U1462 (N_1462,In_588,In_994);
and U1463 (N_1463,In_766,In_668);
or U1464 (N_1464,In_68,In_582);
nand U1465 (N_1465,In_6,In_87);
nand U1466 (N_1466,In_266,In_306);
nand U1467 (N_1467,In_647,In_251);
and U1468 (N_1468,In_998,In_90);
and U1469 (N_1469,In_144,In_459);
nand U1470 (N_1470,In_275,In_66);
or U1471 (N_1471,In_267,In_142);
or U1472 (N_1472,In_4,In_763);
nor U1473 (N_1473,In_51,In_291);
and U1474 (N_1474,In_103,In_96);
or U1475 (N_1475,In_764,In_749);
nor U1476 (N_1476,In_930,In_419);
nor U1477 (N_1477,In_898,In_781);
nor U1478 (N_1478,In_65,In_83);
or U1479 (N_1479,In_996,In_680);
nor U1480 (N_1480,In_112,In_738);
or U1481 (N_1481,In_923,In_247);
and U1482 (N_1482,In_93,In_753);
nand U1483 (N_1483,In_153,In_988);
and U1484 (N_1484,In_705,In_357);
and U1485 (N_1485,In_660,In_850);
and U1486 (N_1486,In_632,In_368);
or U1487 (N_1487,In_330,In_427);
and U1488 (N_1488,In_712,In_881);
nor U1489 (N_1489,In_708,In_173);
or U1490 (N_1490,In_269,In_42);
or U1491 (N_1491,In_249,In_997);
nor U1492 (N_1492,In_171,In_87);
and U1493 (N_1493,In_832,In_643);
nor U1494 (N_1494,In_327,In_127);
nor U1495 (N_1495,In_862,In_657);
or U1496 (N_1496,In_497,In_357);
nor U1497 (N_1497,In_611,In_190);
and U1498 (N_1498,In_448,In_884);
nor U1499 (N_1499,In_368,In_617);
xnor U1500 (N_1500,In_806,In_716);
and U1501 (N_1501,In_772,In_261);
or U1502 (N_1502,In_764,In_894);
nor U1503 (N_1503,In_201,In_55);
and U1504 (N_1504,In_931,In_635);
or U1505 (N_1505,In_290,In_649);
and U1506 (N_1506,In_866,In_274);
nor U1507 (N_1507,In_711,In_831);
nand U1508 (N_1508,In_467,In_113);
nand U1509 (N_1509,In_711,In_594);
nor U1510 (N_1510,In_592,In_956);
and U1511 (N_1511,In_149,In_973);
nand U1512 (N_1512,In_493,In_753);
and U1513 (N_1513,In_328,In_777);
nor U1514 (N_1514,In_791,In_414);
or U1515 (N_1515,In_571,In_878);
nor U1516 (N_1516,In_813,In_722);
and U1517 (N_1517,In_84,In_558);
and U1518 (N_1518,In_166,In_97);
or U1519 (N_1519,In_614,In_761);
and U1520 (N_1520,In_695,In_399);
and U1521 (N_1521,In_933,In_857);
or U1522 (N_1522,In_194,In_812);
or U1523 (N_1523,In_430,In_79);
nor U1524 (N_1524,In_722,In_350);
nor U1525 (N_1525,In_2,In_448);
nor U1526 (N_1526,In_894,In_835);
nand U1527 (N_1527,In_8,In_463);
nand U1528 (N_1528,In_78,In_508);
xnor U1529 (N_1529,In_85,In_350);
nand U1530 (N_1530,In_479,In_364);
nand U1531 (N_1531,In_468,In_6);
nor U1532 (N_1532,In_178,In_790);
or U1533 (N_1533,In_115,In_771);
nand U1534 (N_1534,In_701,In_730);
nor U1535 (N_1535,In_683,In_922);
and U1536 (N_1536,In_867,In_837);
nand U1537 (N_1537,In_982,In_62);
and U1538 (N_1538,In_614,In_830);
and U1539 (N_1539,In_783,In_733);
or U1540 (N_1540,In_473,In_78);
xor U1541 (N_1541,In_952,In_981);
or U1542 (N_1542,In_327,In_305);
nor U1543 (N_1543,In_456,In_600);
and U1544 (N_1544,In_254,In_408);
and U1545 (N_1545,In_106,In_363);
and U1546 (N_1546,In_506,In_752);
xor U1547 (N_1547,In_293,In_415);
or U1548 (N_1548,In_698,In_195);
nand U1549 (N_1549,In_591,In_634);
or U1550 (N_1550,In_86,In_736);
nor U1551 (N_1551,In_627,In_260);
or U1552 (N_1552,In_942,In_230);
nor U1553 (N_1553,In_844,In_661);
and U1554 (N_1554,In_247,In_22);
nand U1555 (N_1555,In_492,In_845);
nand U1556 (N_1556,In_463,In_503);
nor U1557 (N_1557,In_435,In_796);
and U1558 (N_1558,In_188,In_707);
or U1559 (N_1559,In_162,In_169);
nor U1560 (N_1560,In_429,In_779);
nand U1561 (N_1561,In_113,In_459);
and U1562 (N_1562,In_937,In_637);
nor U1563 (N_1563,In_475,In_239);
and U1564 (N_1564,In_210,In_322);
nor U1565 (N_1565,In_558,In_971);
nand U1566 (N_1566,In_682,In_728);
nor U1567 (N_1567,In_934,In_140);
nand U1568 (N_1568,In_62,In_444);
and U1569 (N_1569,In_6,In_884);
and U1570 (N_1570,In_835,In_719);
and U1571 (N_1571,In_851,In_528);
xor U1572 (N_1572,In_727,In_234);
nor U1573 (N_1573,In_533,In_457);
or U1574 (N_1574,In_150,In_804);
nor U1575 (N_1575,In_616,In_289);
and U1576 (N_1576,In_888,In_629);
nand U1577 (N_1577,In_270,In_682);
or U1578 (N_1578,In_517,In_419);
nor U1579 (N_1579,In_924,In_115);
and U1580 (N_1580,In_231,In_913);
or U1581 (N_1581,In_81,In_397);
and U1582 (N_1582,In_331,In_518);
nand U1583 (N_1583,In_488,In_561);
or U1584 (N_1584,In_867,In_950);
nor U1585 (N_1585,In_302,In_849);
xnor U1586 (N_1586,In_645,In_129);
nand U1587 (N_1587,In_705,In_245);
and U1588 (N_1588,In_199,In_331);
and U1589 (N_1589,In_427,In_716);
nand U1590 (N_1590,In_407,In_67);
nand U1591 (N_1591,In_860,In_344);
and U1592 (N_1592,In_598,In_372);
nor U1593 (N_1593,In_446,In_107);
and U1594 (N_1594,In_962,In_549);
and U1595 (N_1595,In_467,In_414);
nor U1596 (N_1596,In_490,In_644);
and U1597 (N_1597,In_382,In_335);
nor U1598 (N_1598,In_646,In_845);
or U1599 (N_1599,In_529,In_72);
nand U1600 (N_1600,In_649,In_199);
and U1601 (N_1601,In_662,In_469);
and U1602 (N_1602,In_467,In_34);
nor U1603 (N_1603,In_329,In_157);
or U1604 (N_1604,In_324,In_12);
or U1605 (N_1605,In_354,In_524);
or U1606 (N_1606,In_11,In_449);
or U1607 (N_1607,In_889,In_32);
nand U1608 (N_1608,In_583,In_469);
or U1609 (N_1609,In_538,In_967);
nor U1610 (N_1610,In_543,In_437);
nor U1611 (N_1611,In_362,In_659);
and U1612 (N_1612,In_959,In_734);
nand U1613 (N_1613,In_184,In_315);
nand U1614 (N_1614,In_619,In_333);
and U1615 (N_1615,In_333,In_582);
nand U1616 (N_1616,In_409,In_132);
nor U1617 (N_1617,In_630,In_218);
nand U1618 (N_1618,In_701,In_942);
and U1619 (N_1619,In_90,In_390);
nand U1620 (N_1620,In_986,In_536);
nor U1621 (N_1621,In_304,In_195);
and U1622 (N_1622,In_235,In_7);
nand U1623 (N_1623,In_369,In_328);
and U1624 (N_1624,In_437,In_961);
and U1625 (N_1625,In_447,In_639);
nor U1626 (N_1626,In_210,In_193);
or U1627 (N_1627,In_887,In_894);
and U1628 (N_1628,In_796,In_823);
nor U1629 (N_1629,In_954,In_875);
xnor U1630 (N_1630,In_34,In_575);
xor U1631 (N_1631,In_869,In_957);
and U1632 (N_1632,In_710,In_607);
nor U1633 (N_1633,In_136,In_640);
and U1634 (N_1634,In_568,In_160);
nand U1635 (N_1635,In_205,In_682);
nor U1636 (N_1636,In_826,In_348);
nand U1637 (N_1637,In_523,In_868);
and U1638 (N_1638,In_762,In_595);
nand U1639 (N_1639,In_878,In_501);
and U1640 (N_1640,In_184,In_974);
and U1641 (N_1641,In_749,In_407);
nand U1642 (N_1642,In_103,In_195);
nand U1643 (N_1643,In_538,In_352);
or U1644 (N_1644,In_831,In_521);
nor U1645 (N_1645,In_358,In_797);
and U1646 (N_1646,In_843,In_582);
and U1647 (N_1647,In_932,In_183);
or U1648 (N_1648,In_32,In_195);
and U1649 (N_1649,In_26,In_181);
nand U1650 (N_1650,In_333,In_175);
and U1651 (N_1651,In_926,In_36);
or U1652 (N_1652,In_60,In_671);
or U1653 (N_1653,In_924,In_816);
nor U1654 (N_1654,In_805,In_347);
nor U1655 (N_1655,In_744,In_946);
nand U1656 (N_1656,In_269,In_155);
nor U1657 (N_1657,In_504,In_306);
nand U1658 (N_1658,In_414,In_133);
nor U1659 (N_1659,In_108,In_442);
or U1660 (N_1660,In_285,In_933);
nand U1661 (N_1661,In_972,In_906);
or U1662 (N_1662,In_26,In_111);
nor U1663 (N_1663,In_684,In_986);
and U1664 (N_1664,In_527,In_331);
and U1665 (N_1665,In_115,In_371);
nor U1666 (N_1666,In_252,In_317);
and U1667 (N_1667,In_242,In_166);
nand U1668 (N_1668,In_728,In_923);
nand U1669 (N_1669,In_240,In_646);
or U1670 (N_1670,In_895,In_102);
nand U1671 (N_1671,In_716,In_582);
or U1672 (N_1672,In_817,In_725);
and U1673 (N_1673,In_890,In_258);
nand U1674 (N_1674,In_266,In_861);
and U1675 (N_1675,In_269,In_708);
nor U1676 (N_1676,In_832,In_145);
or U1677 (N_1677,In_463,In_35);
nand U1678 (N_1678,In_355,In_206);
and U1679 (N_1679,In_200,In_674);
nand U1680 (N_1680,In_19,In_850);
nor U1681 (N_1681,In_406,In_122);
nor U1682 (N_1682,In_119,In_654);
or U1683 (N_1683,In_30,In_901);
nor U1684 (N_1684,In_141,In_565);
or U1685 (N_1685,In_818,In_879);
nor U1686 (N_1686,In_222,In_805);
or U1687 (N_1687,In_602,In_315);
xnor U1688 (N_1688,In_856,In_518);
or U1689 (N_1689,In_872,In_758);
nand U1690 (N_1690,In_583,In_417);
nand U1691 (N_1691,In_49,In_282);
or U1692 (N_1692,In_126,In_655);
and U1693 (N_1693,In_659,In_797);
or U1694 (N_1694,In_615,In_46);
nand U1695 (N_1695,In_346,In_374);
or U1696 (N_1696,In_15,In_613);
nand U1697 (N_1697,In_943,In_922);
or U1698 (N_1698,In_913,In_567);
or U1699 (N_1699,In_63,In_716);
and U1700 (N_1700,In_394,In_903);
and U1701 (N_1701,In_229,In_222);
or U1702 (N_1702,In_629,In_106);
nand U1703 (N_1703,In_286,In_312);
nor U1704 (N_1704,In_13,In_552);
nand U1705 (N_1705,In_467,In_182);
and U1706 (N_1706,In_955,In_17);
nor U1707 (N_1707,In_433,In_926);
and U1708 (N_1708,In_83,In_840);
nor U1709 (N_1709,In_446,In_106);
or U1710 (N_1710,In_259,In_309);
and U1711 (N_1711,In_524,In_890);
and U1712 (N_1712,In_859,In_497);
nor U1713 (N_1713,In_301,In_724);
and U1714 (N_1714,In_279,In_283);
or U1715 (N_1715,In_411,In_846);
nand U1716 (N_1716,In_8,In_556);
and U1717 (N_1717,In_266,In_166);
or U1718 (N_1718,In_491,In_263);
and U1719 (N_1719,In_295,In_881);
or U1720 (N_1720,In_959,In_142);
nor U1721 (N_1721,In_361,In_108);
nor U1722 (N_1722,In_86,In_855);
nor U1723 (N_1723,In_327,In_845);
or U1724 (N_1724,In_498,In_799);
nor U1725 (N_1725,In_339,In_944);
and U1726 (N_1726,In_479,In_978);
and U1727 (N_1727,In_902,In_791);
and U1728 (N_1728,In_631,In_905);
nor U1729 (N_1729,In_88,In_727);
nand U1730 (N_1730,In_366,In_944);
nand U1731 (N_1731,In_337,In_18);
nand U1732 (N_1732,In_279,In_347);
or U1733 (N_1733,In_480,In_875);
nand U1734 (N_1734,In_869,In_655);
and U1735 (N_1735,In_217,In_212);
or U1736 (N_1736,In_309,In_499);
or U1737 (N_1737,In_992,In_93);
nand U1738 (N_1738,In_749,In_84);
and U1739 (N_1739,In_513,In_204);
or U1740 (N_1740,In_121,In_458);
nand U1741 (N_1741,In_498,In_831);
nand U1742 (N_1742,In_707,In_211);
and U1743 (N_1743,In_961,In_851);
nand U1744 (N_1744,In_828,In_202);
nor U1745 (N_1745,In_72,In_391);
and U1746 (N_1746,In_631,In_676);
or U1747 (N_1747,In_799,In_962);
and U1748 (N_1748,In_995,In_680);
nand U1749 (N_1749,In_435,In_109);
nand U1750 (N_1750,In_551,In_786);
and U1751 (N_1751,In_379,In_503);
nand U1752 (N_1752,In_759,In_915);
nor U1753 (N_1753,In_318,In_198);
nand U1754 (N_1754,In_840,In_448);
or U1755 (N_1755,In_451,In_16);
and U1756 (N_1756,In_2,In_217);
and U1757 (N_1757,In_320,In_135);
nand U1758 (N_1758,In_756,In_487);
or U1759 (N_1759,In_275,In_743);
xnor U1760 (N_1760,In_249,In_686);
and U1761 (N_1761,In_10,In_258);
nor U1762 (N_1762,In_839,In_747);
or U1763 (N_1763,In_437,In_255);
and U1764 (N_1764,In_108,In_285);
nor U1765 (N_1765,In_110,In_896);
and U1766 (N_1766,In_539,In_601);
nand U1767 (N_1767,In_842,In_479);
nor U1768 (N_1768,In_590,In_792);
or U1769 (N_1769,In_893,In_883);
nand U1770 (N_1770,In_807,In_974);
nor U1771 (N_1771,In_780,In_976);
nor U1772 (N_1772,In_678,In_527);
nor U1773 (N_1773,In_227,In_784);
nor U1774 (N_1774,In_336,In_197);
or U1775 (N_1775,In_972,In_896);
nor U1776 (N_1776,In_406,In_498);
or U1777 (N_1777,In_15,In_723);
or U1778 (N_1778,In_642,In_121);
nor U1779 (N_1779,In_262,In_219);
and U1780 (N_1780,In_464,In_84);
or U1781 (N_1781,In_230,In_280);
nor U1782 (N_1782,In_734,In_403);
nor U1783 (N_1783,In_865,In_797);
and U1784 (N_1784,In_475,In_339);
nand U1785 (N_1785,In_487,In_948);
nor U1786 (N_1786,In_239,In_676);
nand U1787 (N_1787,In_512,In_819);
nand U1788 (N_1788,In_179,In_219);
or U1789 (N_1789,In_740,In_434);
nor U1790 (N_1790,In_720,In_987);
nand U1791 (N_1791,In_171,In_136);
nor U1792 (N_1792,In_987,In_446);
or U1793 (N_1793,In_728,In_268);
and U1794 (N_1794,In_489,In_986);
nor U1795 (N_1795,In_692,In_713);
nand U1796 (N_1796,In_326,In_794);
nand U1797 (N_1797,In_858,In_835);
nand U1798 (N_1798,In_902,In_146);
xor U1799 (N_1799,In_65,In_290);
nor U1800 (N_1800,In_79,In_440);
nor U1801 (N_1801,In_285,In_201);
nor U1802 (N_1802,In_269,In_610);
nor U1803 (N_1803,In_778,In_65);
and U1804 (N_1804,In_112,In_302);
xnor U1805 (N_1805,In_314,In_463);
or U1806 (N_1806,In_23,In_464);
or U1807 (N_1807,In_685,In_781);
nor U1808 (N_1808,In_273,In_463);
nor U1809 (N_1809,In_651,In_416);
nor U1810 (N_1810,In_789,In_36);
nand U1811 (N_1811,In_488,In_10);
nand U1812 (N_1812,In_612,In_442);
nor U1813 (N_1813,In_860,In_115);
nor U1814 (N_1814,In_328,In_338);
and U1815 (N_1815,In_713,In_372);
nand U1816 (N_1816,In_986,In_582);
or U1817 (N_1817,In_685,In_427);
nor U1818 (N_1818,In_378,In_141);
nor U1819 (N_1819,In_31,In_373);
and U1820 (N_1820,In_182,In_14);
and U1821 (N_1821,In_452,In_275);
or U1822 (N_1822,In_791,In_256);
and U1823 (N_1823,In_752,In_989);
or U1824 (N_1824,In_710,In_510);
or U1825 (N_1825,In_409,In_184);
or U1826 (N_1826,In_95,In_339);
and U1827 (N_1827,In_184,In_111);
and U1828 (N_1828,In_390,In_246);
nor U1829 (N_1829,In_86,In_699);
or U1830 (N_1830,In_941,In_971);
and U1831 (N_1831,In_655,In_422);
xnor U1832 (N_1832,In_784,In_819);
nand U1833 (N_1833,In_622,In_457);
and U1834 (N_1834,In_156,In_749);
nor U1835 (N_1835,In_292,In_825);
nand U1836 (N_1836,In_853,In_360);
and U1837 (N_1837,In_99,In_443);
nand U1838 (N_1838,In_370,In_421);
nand U1839 (N_1839,In_132,In_637);
or U1840 (N_1840,In_50,In_681);
or U1841 (N_1841,In_845,In_467);
and U1842 (N_1842,In_80,In_264);
xnor U1843 (N_1843,In_196,In_44);
or U1844 (N_1844,In_677,In_429);
and U1845 (N_1845,In_646,In_543);
nand U1846 (N_1846,In_73,In_350);
and U1847 (N_1847,In_423,In_931);
or U1848 (N_1848,In_829,In_582);
or U1849 (N_1849,In_190,In_555);
nand U1850 (N_1850,In_898,In_30);
and U1851 (N_1851,In_703,In_94);
or U1852 (N_1852,In_822,In_211);
xor U1853 (N_1853,In_175,In_764);
or U1854 (N_1854,In_583,In_6);
or U1855 (N_1855,In_597,In_187);
or U1856 (N_1856,In_569,In_42);
xnor U1857 (N_1857,In_512,In_412);
and U1858 (N_1858,In_867,In_563);
or U1859 (N_1859,In_254,In_78);
or U1860 (N_1860,In_346,In_967);
nor U1861 (N_1861,In_920,In_545);
or U1862 (N_1862,In_760,In_999);
xor U1863 (N_1863,In_822,In_89);
or U1864 (N_1864,In_774,In_542);
nor U1865 (N_1865,In_645,In_567);
nor U1866 (N_1866,In_815,In_580);
and U1867 (N_1867,In_516,In_933);
nor U1868 (N_1868,In_100,In_831);
nand U1869 (N_1869,In_42,In_870);
nor U1870 (N_1870,In_473,In_268);
nor U1871 (N_1871,In_631,In_513);
nor U1872 (N_1872,In_95,In_703);
nand U1873 (N_1873,In_52,In_727);
nor U1874 (N_1874,In_983,In_702);
and U1875 (N_1875,In_806,In_835);
nor U1876 (N_1876,In_34,In_586);
and U1877 (N_1877,In_213,In_566);
or U1878 (N_1878,In_782,In_607);
nand U1879 (N_1879,In_425,In_967);
and U1880 (N_1880,In_615,In_765);
nor U1881 (N_1881,In_265,In_657);
nor U1882 (N_1882,In_946,In_655);
and U1883 (N_1883,In_840,In_874);
and U1884 (N_1884,In_183,In_230);
or U1885 (N_1885,In_386,In_479);
nor U1886 (N_1886,In_967,In_340);
nor U1887 (N_1887,In_449,In_606);
xor U1888 (N_1888,In_340,In_588);
or U1889 (N_1889,In_484,In_853);
or U1890 (N_1890,In_494,In_142);
nand U1891 (N_1891,In_294,In_917);
nand U1892 (N_1892,In_585,In_697);
nor U1893 (N_1893,In_429,In_676);
nor U1894 (N_1894,In_279,In_373);
or U1895 (N_1895,In_254,In_526);
nand U1896 (N_1896,In_912,In_263);
nand U1897 (N_1897,In_362,In_555);
nand U1898 (N_1898,In_871,In_812);
nand U1899 (N_1899,In_74,In_802);
or U1900 (N_1900,In_292,In_293);
nor U1901 (N_1901,In_465,In_444);
nand U1902 (N_1902,In_113,In_614);
nor U1903 (N_1903,In_18,In_807);
or U1904 (N_1904,In_487,In_176);
and U1905 (N_1905,In_933,In_455);
nor U1906 (N_1906,In_50,In_546);
and U1907 (N_1907,In_233,In_91);
nand U1908 (N_1908,In_480,In_144);
or U1909 (N_1909,In_629,In_687);
nor U1910 (N_1910,In_883,In_115);
nand U1911 (N_1911,In_725,In_792);
or U1912 (N_1912,In_598,In_213);
and U1913 (N_1913,In_334,In_739);
or U1914 (N_1914,In_224,In_297);
and U1915 (N_1915,In_894,In_399);
nand U1916 (N_1916,In_822,In_325);
nand U1917 (N_1917,In_924,In_756);
nand U1918 (N_1918,In_302,In_552);
nor U1919 (N_1919,In_289,In_693);
nand U1920 (N_1920,In_67,In_515);
and U1921 (N_1921,In_623,In_969);
and U1922 (N_1922,In_595,In_35);
and U1923 (N_1923,In_866,In_454);
or U1924 (N_1924,In_89,In_965);
nand U1925 (N_1925,In_734,In_88);
nand U1926 (N_1926,In_185,In_27);
nand U1927 (N_1927,In_354,In_550);
nand U1928 (N_1928,In_882,In_773);
and U1929 (N_1929,In_294,In_185);
and U1930 (N_1930,In_580,In_242);
nand U1931 (N_1931,In_33,In_336);
nand U1932 (N_1932,In_12,In_978);
nand U1933 (N_1933,In_13,In_497);
and U1934 (N_1934,In_557,In_776);
xnor U1935 (N_1935,In_939,In_698);
or U1936 (N_1936,In_844,In_822);
nor U1937 (N_1937,In_483,In_492);
xor U1938 (N_1938,In_476,In_447);
nand U1939 (N_1939,In_435,In_720);
nor U1940 (N_1940,In_769,In_379);
nor U1941 (N_1941,In_127,In_622);
or U1942 (N_1942,In_294,In_852);
nand U1943 (N_1943,In_773,In_320);
nor U1944 (N_1944,In_189,In_289);
nand U1945 (N_1945,In_165,In_835);
or U1946 (N_1946,In_999,In_992);
or U1947 (N_1947,In_980,In_240);
nor U1948 (N_1948,In_523,In_92);
and U1949 (N_1949,In_975,In_679);
or U1950 (N_1950,In_137,In_746);
nand U1951 (N_1951,In_70,In_273);
nor U1952 (N_1952,In_13,In_192);
or U1953 (N_1953,In_881,In_438);
and U1954 (N_1954,In_704,In_552);
xnor U1955 (N_1955,In_819,In_866);
nand U1956 (N_1956,In_225,In_49);
and U1957 (N_1957,In_191,In_91);
or U1958 (N_1958,In_871,In_117);
and U1959 (N_1959,In_427,In_699);
nand U1960 (N_1960,In_805,In_491);
nor U1961 (N_1961,In_467,In_636);
and U1962 (N_1962,In_69,In_951);
or U1963 (N_1963,In_347,In_195);
xnor U1964 (N_1964,In_949,In_668);
nand U1965 (N_1965,In_903,In_937);
or U1966 (N_1966,In_676,In_436);
or U1967 (N_1967,In_371,In_610);
and U1968 (N_1968,In_322,In_333);
or U1969 (N_1969,In_74,In_323);
nand U1970 (N_1970,In_114,In_518);
nor U1971 (N_1971,In_660,In_855);
and U1972 (N_1972,In_472,In_668);
and U1973 (N_1973,In_984,In_988);
or U1974 (N_1974,In_330,In_597);
or U1975 (N_1975,In_904,In_328);
or U1976 (N_1976,In_824,In_300);
or U1977 (N_1977,In_704,In_452);
xor U1978 (N_1978,In_699,In_404);
nand U1979 (N_1979,In_0,In_757);
nor U1980 (N_1980,In_68,In_702);
nor U1981 (N_1981,In_625,In_703);
or U1982 (N_1982,In_146,In_798);
nor U1983 (N_1983,In_749,In_970);
and U1984 (N_1984,In_754,In_271);
nor U1985 (N_1985,In_88,In_480);
nand U1986 (N_1986,In_167,In_139);
nor U1987 (N_1987,In_650,In_852);
and U1988 (N_1988,In_928,In_287);
nand U1989 (N_1989,In_12,In_883);
nor U1990 (N_1990,In_6,In_274);
or U1991 (N_1991,In_230,In_188);
nand U1992 (N_1992,In_305,In_997);
nand U1993 (N_1993,In_250,In_470);
nor U1994 (N_1994,In_195,In_497);
nor U1995 (N_1995,In_332,In_696);
nand U1996 (N_1996,In_292,In_509);
nor U1997 (N_1997,In_142,In_128);
or U1998 (N_1998,In_779,In_513);
nor U1999 (N_1999,In_680,In_803);
and U2000 (N_2000,N_564,N_545);
and U2001 (N_2001,N_1049,N_1989);
and U2002 (N_2002,N_1520,N_361);
and U2003 (N_2003,N_83,N_493);
and U2004 (N_2004,N_771,N_1125);
or U2005 (N_2005,N_1205,N_72);
or U2006 (N_2006,N_1339,N_427);
nor U2007 (N_2007,N_196,N_1206);
nand U2008 (N_2008,N_1383,N_1760);
nand U2009 (N_2009,N_1578,N_277);
nand U2010 (N_2010,N_1755,N_1690);
nand U2011 (N_2011,N_218,N_1374);
and U2012 (N_2012,N_1447,N_654);
or U2013 (N_2013,N_1421,N_579);
nand U2014 (N_2014,N_1695,N_1112);
nor U2015 (N_2015,N_1918,N_517);
nand U2016 (N_2016,N_942,N_1614);
and U2017 (N_2017,N_1845,N_1319);
and U2018 (N_2018,N_115,N_323);
nand U2019 (N_2019,N_1917,N_1671);
or U2020 (N_2020,N_1435,N_1192);
nor U2021 (N_2021,N_630,N_1854);
nand U2022 (N_2022,N_1764,N_421);
nand U2023 (N_2023,N_1281,N_743);
nor U2024 (N_2024,N_242,N_293);
and U2025 (N_2025,N_643,N_718);
and U2026 (N_2026,N_300,N_442);
nand U2027 (N_2027,N_375,N_145);
and U2028 (N_2028,N_1804,N_749);
or U2029 (N_2029,N_711,N_1636);
or U2030 (N_2030,N_1083,N_1911);
nand U2031 (N_2031,N_1489,N_169);
or U2032 (N_2032,N_1219,N_1343);
or U2033 (N_2033,N_719,N_1066);
nand U2034 (N_2034,N_338,N_1922);
nand U2035 (N_2035,N_156,N_129);
and U2036 (N_2036,N_27,N_1229);
nand U2037 (N_2037,N_456,N_287);
nor U2038 (N_2038,N_1036,N_127);
and U2039 (N_2039,N_366,N_1617);
nand U2040 (N_2040,N_316,N_922);
nand U2041 (N_2041,N_1752,N_486);
nand U2042 (N_2042,N_1446,N_1988);
or U2043 (N_2043,N_617,N_987);
and U2044 (N_2044,N_755,N_1580);
and U2045 (N_2045,N_1373,N_921);
nor U2046 (N_2046,N_1579,N_1562);
and U2047 (N_2047,N_931,N_932);
or U2048 (N_2048,N_1660,N_820);
nand U2049 (N_2049,N_346,N_822);
and U2050 (N_2050,N_32,N_1960);
and U2051 (N_2051,N_1784,N_143);
or U2052 (N_2052,N_1358,N_1728);
nor U2053 (N_2053,N_1789,N_933);
nor U2054 (N_2054,N_62,N_702);
nor U2055 (N_2055,N_529,N_886);
nor U2056 (N_2056,N_31,N_867);
or U2057 (N_2057,N_1001,N_237);
or U2058 (N_2058,N_1443,N_109);
nor U2059 (N_2059,N_1243,N_451);
nand U2060 (N_2060,N_1076,N_123);
xor U2061 (N_2061,N_190,N_289);
nor U2062 (N_2062,N_1424,N_1089);
or U2063 (N_2063,N_312,N_21);
xor U2064 (N_2064,N_1283,N_1927);
or U2065 (N_2065,N_495,N_1821);
nor U2066 (N_2066,N_1277,N_1770);
or U2067 (N_2067,N_86,N_211);
or U2068 (N_2068,N_1890,N_843);
nand U2069 (N_2069,N_432,N_849);
nand U2070 (N_2070,N_1148,N_1590);
nor U2071 (N_2071,N_393,N_1663);
and U2072 (N_2072,N_1965,N_1893);
nor U2073 (N_2073,N_446,N_1644);
or U2074 (N_2074,N_1384,N_118);
or U2075 (N_2075,N_675,N_496);
nand U2076 (N_2076,N_518,N_982);
nor U2077 (N_2077,N_1753,N_1892);
or U2078 (N_2078,N_176,N_317);
and U2079 (N_2079,N_1322,N_126);
or U2080 (N_2080,N_725,N_1492);
and U2081 (N_2081,N_1667,N_1244);
and U2082 (N_2082,N_833,N_204);
and U2083 (N_2083,N_816,N_1838);
nand U2084 (N_2084,N_175,N_1315);
nor U2085 (N_2085,N_1907,N_618);
nand U2086 (N_2086,N_1070,N_923);
nand U2087 (N_2087,N_917,N_1682);
and U2088 (N_2088,N_508,N_796);
or U2089 (N_2089,N_1003,N_340);
nor U2090 (N_2090,N_908,N_25);
nor U2091 (N_2091,N_459,N_436);
nand U2092 (N_2092,N_983,N_1844);
or U2093 (N_2093,N_1510,N_1296);
nor U2094 (N_2094,N_1805,N_504);
or U2095 (N_2095,N_1883,N_1146);
nor U2096 (N_2096,N_1596,N_1938);
and U2097 (N_2097,N_756,N_798);
nor U2098 (N_2098,N_305,N_1295);
nor U2099 (N_2099,N_1956,N_23);
nor U2100 (N_2100,N_851,N_1191);
nand U2101 (N_2101,N_708,N_1937);
and U2102 (N_2102,N_1353,N_65);
or U2103 (N_2103,N_1109,N_871);
nor U2104 (N_2104,N_1400,N_1376);
or U2105 (N_2105,N_360,N_195);
and U2106 (N_2106,N_882,N_863);
nor U2107 (N_2107,N_542,N_1891);
nor U2108 (N_2108,N_1778,N_1952);
nor U2109 (N_2109,N_552,N_1055);
or U2110 (N_2110,N_1847,N_160);
or U2111 (N_2111,N_1857,N_1173);
and U2112 (N_2112,N_1002,N_434);
nand U2113 (N_2113,N_995,N_888);
or U2114 (N_2114,N_1433,N_1203);
nand U2115 (N_2115,N_980,N_993);
and U2116 (N_2116,N_1889,N_154);
or U2117 (N_2117,N_532,N_1265);
nor U2118 (N_2118,N_1272,N_1439);
nor U2119 (N_2119,N_536,N_868);
nand U2120 (N_2120,N_1485,N_153);
nand U2121 (N_2121,N_1618,N_945);
and U2122 (N_2122,N_1680,N_331);
and U2123 (N_2123,N_74,N_584);
and U2124 (N_2124,N_824,N_230);
and U2125 (N_2125,N_207,N_117);
or U2126 (N_2126,N_1042,N_597);
nand U2127 (N_2127,N_150,N_59);
and U2128 (N_2128,N_1628,N_1862);
and U2129 (N_2129,N_120,N_1454);
nor U2130 (N_2130,N_1311,N_1121);
and U2131 (N_2131,N_979,N_779);
or U2132 (N_2132,N_678,N_1067);
nor U2133 (N_2133,N_1739,N_314);
or U2134 (N_2134,N_1422,N_138);
nand U2135 (N_2135,N_813,N_620);
or U2136 (N_2136,N_1887,N_1776);
xnor U2137 (N_2137,N_1334,N_1233);
and U2138 (N_2138,N_1387,N_498);
or U2139 (N_2139,N_1954,N_1758);
xor U2140 (N_2140,N_1250,N_1405);
and U2141 (N_2141,N_477,N_114);
nand U2142 (N_2142,N_1713,N_1584);
nand U2143 (N_2143,N_531,N_1585);
nand U2144 (N_2144,N_1060,N_1212);
nand U2145 (N_2145,N_1084,N_1073);
nor U2146 (N_2146,N_406,N_1503);
and U2147 (N_2147,N_170,N_927);
or U2148 (N_2148,N_834,N_958);
or U2149 (N_2149,N_232,N_1249);
and U2150 (N_2150,N_919,N_1106);
nand U2151 (N_2151,N_844,N_119);
or U2152 (N_2152,N_1831,N_497);
and U2153 (N_2153,N_1327,N_1882);
nand U2154 (N_2154,N_1855,N_1210);
nor U2155 (N_2155,N_1341,N_1472);
nand U2156 (N_2156,N_94,N_180);
nand U2157 (N_2157,N_914,N_954);
and U2158 (N_2158,N_1523,N_227);
and U2159 (N_2159,N_1627,N_152);
nor U2160 (N_2160,N_1525,N_1412);
nand U2161 (N_2161,N_1709,N_1289);
nand U2162 (N_2162,N_609,N_1043);
xnor U2163 (N_2163,N_44,N_805);
and U2164 (N_2164,N_861,N_1701);
or U2165 (N_2165,N_135,N_836);
and U2166 (N_2166,N_371,N_694);
nor U2167 (N_2167,N_9,N_774);
nand U2168 (N_2168,N_1589,N_1615);
nor U2169 (N_2169,N_281,N_1732);
and U2170 (N_2170,N_1325,N_1624);
and U2171 (N_2171,N_1564,N_1087);
or U2172 (N_2172,N_296,N_1669);
or U2173 (N_2173,N_1587,N_350);
and U2174 (N_2174,N_1340,N_487);
nor U2175 (N_2175,N_381,N_348);
nand U2176 (N_2176,N_1824,N_972);
and U2177 (N_2177,N_193,N_1631);
or U2178 (N_2178,N_1519,N_869);
or U2179 (N_2179,N_918,N_409);
and U2180 (N_2180,N_1874,N_1176);
nand U2181 (N_2181,N_1330,N_158);
and U2182 (N_2182,N_1939,N_1116);
and U2183 (N_2183,N_1639,N_373);
or U2184 (N_2184,N_1186,N_234);
and U2185 (N_2185,N_500,N_61);
and U2186 (N_2186,N_1885,N_194);
and U2187 (N_2187,N_627,N_1935);
nand U2188 (N_2188,N_261,N_644);
nor U2189 (N_2189,N_971,N_1720);
nor U2190 (N_2190,N_677,N_1015);
nor U2191 (N_2191,N_1946,N_1910);
nor U2192 (N_2192,N_1021,N_470);
or U2193 (N_2193,N_1724,N_191);
nand U2194 (N_2194,N_550,N_1393);
and U2195 (N_2195,N_1127,N_872);
and U2196 (N_2196,N_1287,N_1829);
or U2197 (N_2197,N_580,N_377);
nand U2198 (N_2198,N_1098,N_857);
or U2199 (N_2199,N_853,N_947);
nand U2200 (N_2200,N_1275,N_1773);
or U2201 (N_2201,N_997,N_1529);
or U2202 (N_2202,N_1128,N_174);
nand U2203 (N_2203,N_99,N_1411);
xor U2204 (N_2204,N_1375,N_262);
and U2205 (N_2205,N_670,N_1687);
nand U2206 (N_2206,N_1135,N_359);
or U2207 (N_2207,N_1511,N_826);
and U2208 (N_2208,N_765,N_1350);
nor U2209 (N_2209,N_353,N_511);
nor U2210 (N_2210,N_1553,N_610);
and U2211 (N_2211,N_848,N_327);
and U2212 (N_2212,N_1572,N_1533);
or U2213 (N_2213,N_1793,N_1574);
and U2214 (N_2214,N_1011,N_1198);
and U2215 (N_2215,N_1715,N_1050);
and U2216 (N_2216,N_1561,N_1502);
or U2217 (N_2217,N_1969,N_1677);
and U2218 (N_2218,N_1994,N_1924);
nor U2219 (N_2219,N_852,N_1936);
and U2220 (N_2220,N_769,N_267);
and U2221 (N_2221,N_1896,N_683);
or U2222 (N_2222,N_611,N_1547);
nor U2223 (N_2223,N_422,N_854);
or U2224 (N_2224,N_1783,N_659);
or U2225 (N_2225,N_587,N_619);
nor U2226 (N_2226,N_1966,N_1072);
nor U2227 (N_2227,N_468,N_786);
nor U2228 (N_2228,N_315,N_516);
and U2229 (N_2229,N_1710,N_1257);
nor U2230 (N_2230,N_593,N_1575);
or U2231 (N_2231,N_1286,N_132);
nand U2232 (N_2232,N_271,N_548);
nor U2233 (N_2233,N_1174,N_1745);
nand U2234 (N_2234,N_1723,N_162);
nand U2235 (N_2235,N_1200,N_624);
nor U2236 (N_2236,N_900,N_808);
and U2237 (N_2237,N_60,N_1095);
nand U2238 (N_2238,N_103,N_1056);
or U2239 (N_2239,N_1497,N_777);
nor U2240 (N_2240,N_530,N_1306);
or U2241 (N_2241,N_1879,N_159);
and U2242 (N_2242,N_1856,N_1241);
nand U2243 (N_2243,N_1679,N_33);
nand U2244 (N_2244,N_490,N_1288);
nand U2245 (N_2245,N_1674,N_576);
nor U2246 (N_2246,N_1461,N_806);
nor U2247 (N_2247,N_1803,N_1538);
and U2248 (N_2248,N_622,N_669);
or U2249 (N_2249,N_151,N_450);
and U2250 (N_2250,N_326,N_915);
nand U2251 (N_2251,N_1208,N_1901);
nor U2252 (N_2252,N_1651,N_286);
and U2253 (N_2253,N_387,N_1977);
nand U2254 (N_2254,N_1835,N_1023);
nand U2255 (N_2255,N_1704,N_1594);
nand U2256 (N_2256,N_841,N_36);
or U2257 (N_2257,N_1657,N_946);
xor U2258 (N_2258,N_1133,N_819);
nand U2259 (N_2259,N_1762,N_653);
or U2260 (N_2260,N_1419,N_686);
nor U2261 (N_2261,N_1025,N_607);
nor U2262 (N_2262,N_1742,N_1649);
nor U2263 (N_2263,N_181,N_344);
nor U2264 (N_2264,N_1157,N_462);
xor U2265 (N_2265,N_423,N_832);
nor U2266 (N_2266,N_1534,N_1779);
nand U2267 (N_2267,N_512,N_1386);
nand U2268 (N_2268,N_95,N_288);
or U2269 (N_2269,N_1973,N_1221);
nor U2270 (N_2270,N_1873,N_429);
nor U2271 (N_2271,N_1491,N_538);
nor U2272 (N_2272,N_229,N_1979);
nor U2273 (N_2273,N_1138,N_1389);
nor U2274 (N_2274,N_524,N_1708);
nand U2275 (N_2275,N_1160,N_1569);
nand U2276 (N_2276,N_1550,N_1217);
nor U2277 (N_2277,N_1749,N_1766);
or U2278 (N_2278,N_10,N_1848);
nor U2279 (N_2279,N_829,N_628);
nand U2280 (N_2280,N_1817,N_1787);
or U2281 (N_2281,N_457,N_664);
and U2282 (N_2282,N_1344,N_1797);
nand U2283 (N_2283,N_105,N_673);
nor U2284 (N_2284,N_1494,N_1512);
nand U2285 (N_2285,N_727,N_1134);
nand U2286 (N_2286,N_471,N_1466);
xor U2287 (N_2287,N_292,N_1171);
nor U2288 (N_2288,N_1888,N_1189);
and U2289 (N_2289,N_1456,N_1031);
and U2290 (N_2290,N_1482,N_173);
and U2291 (N_2291,N_934,N_1366);
or U2292 (N_2292,N_1030,N_1463);
or U2293 (N_2293,N_1634,N_122);
nor U2294 (N_2294,N_1744,N_986);
nor U2295 (N_2295,N_108,N_325);
nand U2296 (N_2296,N_1111,N_1273);
and U2297 (N_2297,N_1961,N_1409);
xnor U2298 (N_2298,N_163,N_726);
nor U2299 (N_2299,N_45,N_1788);
and U2300 (N_2300,N_1396,N_284);
or U2301 (N_2301,N_1323,N_825);
and U2302 (N_2302,N_1640,N_944);
nor U2303 (N_2303,N_1434,N_793);
nand U2304 (N_2304,N_1402,N_1673);
nand U2305 (N_2305,N_1140,N_1798);
or U2306 (N_2306,N_1555,N_655);
nand U2307 (N_2307,N_1602,N_1459);
xor U2308 (N_2308,N_1790,N_662);
and U2309 (N_2309,N_1242,N_1354);
or U2310 (N_2310,N_910,N_1501);
and U2311 (N_2311,N_125,N_41);
and U2312 (N_2312,N_1702,N_263);
and U2313 (N_2313,N_1582,N_1239);
nor U2314 (N_2314,N_341,N_1488);
nand U2315 (N_2315,N_1761,N_887);
nor U2316 (N_2316,N_370,N_1302);
and U2317 (N_2317,N_689,N_1825);
xnor U2318 (N_2318,N_1567,N_1577);
and U2319 (N_2319,N_328,N_911);
nand U2320 (N_2320,N_959,N_623);
and U2321 (N_2321,N_1841,N_715);
and U2322 (N_2322,N_555,N_551);
or U2323 (N_2323,N_404,N_364);
and U2324 (N_2324,N_713,N_978);
or U2325 (N_2325,N_894,N_144);
nor U2326 (N_2326,N_948,N_909);
and U2327 (N_2327,N_684,N_710);
and U2328 (N_2328,N_1253,N_385);
nor U2329 (N_2329,N_1655,N_1871);
or U2330 (N_2330,N_951,N_1780);
and U2331 (N_2331,N_1981,N_301);
or U2332 (N_2332,N_68,N_1929);
nor U2333 (N_2333,N_697,N_772);
nand U2334 (N_2334,N_1291,N_881);
nor U2335 (N_2335,N_1132,N_1000);
or U2336 (N_2336,N_828,N_7);
nor U2337 (N_2337,N_403,N_401);
nor U2338 (N_2338,N_1899,N_1863);
and U2339 (N_2339,N_509,N_294);
nand U2340 (N_2340,N_56,N_112);
nand U2341 (N_2341,N_554,N_840);
or U2342 (N_2342,N_443,N_1734);
nor U2343 (N_2343,N_1612,N_1107);
or U2344 (N_2344,N_1490,N_397);
and U2345 (N_2345,N_1545,N_202);
nor U2346 (N_2346,N_1448,N_313);
nand U2347 (N_2347,N_1451,N_811);
nand U2348 (N_2348,N_330,N_896);
nor U2349 (N_2349,N_592,N_924);
nand U2350 (N_2350,N_636,N_148);
nand U2351 (N_2351,N_11,N_562);
and U2352 (N_2352,N_1041,N_1062);
and U2353 (N_2353,N_753,N_1364);
nand U2354 (N_2354,N_311,N_795);
or U2355 (N_2355,N_1033,N_342);
nor U2356 (N_2356,N_1026,N_1183);
nand U2357 (N_2357,N_1395,N_19);
and U2358 (N_2358,N_437,N_791);
and U2359 (N_2359,N_809,N_320);
or U2360 (N_2360,N_1775,N_1641);
nand U2361 (N_2361,N_1006,N_1867);
and U2362 (N_2362,N_994,N_560);
nand U2363 (N_2363,N_950,N_1818);
or U2364 (N_2364,N_258,N_801);
nand U2365 (N_2365,N_735,N_380);
and U2366 (N_2366,N_378,N_415);
or U2367 (N_2367,N_1260,N_615);
and U2368 (N_2368,N_1093,N_1811);
nand U2369 (N_2369,N_693,N_1007);
and U2370 (N_2370,N_939,N_501);
nor U2371 (N_2371,N_1057,N_1986);
or U2372 (N_2372,N_1096,N_1933);
and U2373 (N_2373,N_1470,N_39);
or U2374 (N_2374,N_1182,N_147);
or U2375 (N_2375,N_20,N_667);
or U2376 (N_2376,N_1207,N_570);
and U2377 (N_2377,N_155,N_1843);
and U2378 (N_2378,N_1086,N_1630);
or U2379 (N_2379,N_859,N_40);
xor U2380 (N_2380,N_1931,N_778);
and U2381 (N_2381,N_1638,N_186);
nand U2382 (N_2382,N_1591,N_598);
and U2383 (N_2383,N_1968,N_249);
or U2384 (N_2384,N_601,N_177);
nand U2385 (N_2385,N_1997,N_799);
and U2386 (N_2386,N_1371,N_210);
and U2387 (N_2387,N_585,N_1201);
or U2388 (N_2388,N_1022,N_784);
and U2389 (N_2389,N_1149,N_1165);
xor U2390 (N_2390,N_1683,N_1763);
nor U2391 (N_2391,N_969,N_974);
nor U2392 (N_2392,N_1970,N_803);
nor U2393 (N_2393,N_321,N_876);
and U2394 (N_2394,N_637,N_57);
nor U2395 (N_2395,N_722,N_463);
nor U2396 (N_2396,N_1204,N_1609);
and U2397 (N_2397,N_533,N_503);
nand U2398 (N_2398,N_1916,N_566);
nor U2399 (N_2399,N_1934,N_1278);
xor U2400 (N_2400,N_187,N_740);
or U2401 (N_2401,N_221,N_873);
xnor U2402 (N_2402,N_1832,N_407);
nand U2403 (N_2403,N_1958,N_1849);
or U2404 (N_2404,N_304,N_1996);
or U2405 (N_2405,N_362,N_1484);
nor U2406 (N_2406,N_1750,N_1468);
nor U2407 (N_2407,N_812,N_890);
or U2408 (N_2408,N_981,N_671);
or U2409 (N_2409,N_431,N_233);
and U2410 (N_2410,N_64,N_426);
or U2411 (N_2411,N_1263,N_704);
or U2412 (N_2412,N_131,N_1228);
and U2413 (N_2413,N_439,N_775);
xor U2414 (N_2414,N_1279,N_1114);
nor U2415 (N_2415,N_1016,N_1508);
nor U2416 (N_2416,N_1372,N_1799);
xnor U2417 (N_2417,N_1622,N_1450);
and U2418 (N_2418,N_1517,N_1008);
nor U2419 (N_2419,N_1842,N_514);
nor U2420 (N_2420,N_741,N_1215);
and U2421 (N_2421,N_382,N_1426);
nor U2422 (N_2422,N_124,N_1046);
nor U2423 (N_2423,N_1202,N_213);
and U2424 (N_2424,N_738,N_1542);
or U2425 (N_2425,N_817,N_1188);
nand U2426 (N_2426,N_821,N_1403);
or U2427 (N_2427,N_1665,N_50);
nand U2428 (N_2428,N_1880,N_690);
or U2429 (N_2429,N_640,N_557);
nor U2430 (N_2430,N_51,N_238);
and U2431 (N_2431,N_1051,N_395);
and U2432 (N_2432,N_1531,N_192);
and U2433 (N_2433,N_502,N_225);
nor U2434 (N_2434,N_188,N_16);
and U2435 (N_2435,N_4,N_1606);
or U2436 (N_2436,N_1180,N_334);
and U2437 (N_2437,N_680,N_63);
nor U2438 (N_2438,N_1052,N_49);
nand U2439 (N_2439,N_1115,N_1099);
nand U2440 (N_2440,N_1676,N_413);
or U2441 (N_2441,N_1347,N_1987);
and U2442 (N_2442,N_1978,N_641);
and U2443 (N_2443,N_1356,N_1126);
nor U2444 (N_2444,N_1297,N_265);
nor U2445 (N_2445,N_1616,N_206);
xor U2446 (N_2446,N_1020,N_1474);
nand U2447 (N_2447,N_345,N_1795);
nor U2448 (N_2448,N_1740,N_556);
and U2449 (N_2449,N_1355,N_1568);
nand U2450 (N_2450,N_748,N_133);
or U2451 (N_2451,N_157,N_770);
and U2452 (N_2452,N_319,N_492);
or U2453 (N_2453,N_1159,N_1172);
nor U2454 (N_2454,N_1993,N_1707);
nor U2455 (N_2455,N_1427,N_855);
nand U2456 (N_2456,N_1091,N_1619);
and U2457 (N_2457,N_1689,N_1082);
and U2458 (N_2458,N_69,N_1156);
nor U2459 (N_2459,N_48,N_1626);
and U2460 (N_2460,N_1394,N_1876);
nor U2461 (N_2461,N_1471,N_106);
nand U2462 (N_2462,N_605,N_466);
nand U2463 (N_2463,N_303,N_1809);
and U2464 (N_2464,N_1223,N_12);
or U2465 (N_2465,N_838,N_898);
or U2466 (N_2466,N_1187,N_569);
nor U2467 (N_2467,N_365,N_14);
nand U2468 (N_2468,N_200,N_1342);
or U2469 (N_2469,N_789,N_573);
nand U2470 (N_2470,N_1436,N_52);
or U2471 (N_2471,N_467,N_252);
nand U2472 (N_2472,N_1919,N_1566);
and U2473 (N_2473,N_101,N_1620);
nand U2474 (N_2474,N_767,N_1706);
nor U2475 (N_2475,N_1236,N_1028);
or U2476 (N_2476,N_1741,N_1559);
nand U2477 (N_2477,N_1774,N_639);
or U2478 (N_2478,N_1772,N_1310);
and U2479 (N_2479,N_571,N_484);
nor U2480 (N_2480,N_878,N_102);
nor U2481 (N_2481,N_754,N_629);
or U2482 (N_2482,N_998,N_1633);
nand U2483 (N_2483,N_480,N_1059);
nand U2484 (N_2484,N_130,N_13);
nor U2485 (N_2485,N_1711,N_77);
xor U2486 (N_2486,N_136,N_269);
nand U2487 (N_2487,N_583,N_1230);
nor U2488 (N_2488,N_482,N_1943);
nor U2489 (N_2489,N_43,N_1248);
and U2490 (N_2490,N_1833,N_510);
and U2491 (N_2491,N_219,N_1232);
nand U2492 (N_2492,N_1332,N_651);
nand U2493 (N_2493,N_245,N_1816);
and U2494 (N_2494,N_790,N_1635);
nand U2495 (N_2495,N_961,N_1320);
nor U2496 (N_2496,N_1407,N_1352);
and U2497 (N_2497,N_1331,N_1826);
nor U2498 (N_2498,N_1827,N_1653);
and U2499 (N_2499,N_1012,N_860);
or U2500 (N_2500,N_706,N_374);
or U2501 (N_2501,N_1768,N_1869);
or U2502 (N_2502,N_438,N_241);
nand U2503 (N_2503,N_1019,N_613);
nand U2504 (N_2504,N_260,N_1398);
nor U2505 (N_2505,N_1040,N_1326);
or U2506 (N_2506,N_1369,N_299);
nand U2507 (N_2507,N_110,N_534);
xnor U2508 (N_2508,N_247,N_634);
or U2509 (N_2509,N_1336,N_561);
nand U2510 (N_2510,N_1558,N_540);
nor U2511 (N_2511,N_985,N_696);
nand U2512 (N_2512,N_1736,N_97);
nand U2513 (N_2513,N_1851,N_76);
or U2514 (N_2514,N_214,N_1264);
and U2515 (N_2515,N_1444,N_604);
nor U2516 (N_2516,N_1539,N_67);
nor U2517 (N_2517,N_1077,N_441);
or U2518 (N_2518,N_1925,N_322);
nor U2519 (N_2519,N_308,N_1101);
nor U2520 (N_2520,N_1800,N_1048);
nor U2521 (N_2521,N_1581,N_15);
or U2522 (N_2522,N_1654,N_1377);
nand U2523 (N_2523,N_42,N_537);
nand U2524 (N_2524,N_1840,N_999);
nand U2525 (N_2525,N_473,N_818);
and U2526 (N_2526,N_400,N_167);
nand U2527 (N_2527,N_1153,N_1467);
or U2528 (N_2528,N_1625,N_329);
or U2529 (N_2529,N_757,N_412);
nand U2530 (N_2530,N_1613,N_383);
and U2531 (N_2531,N_1004,N_96);
or U2532 (N_2532,N_1449,N_476);
xnor U2533 (N_2533,N_1014,N_1068);
or U2534 (N_2534,N_22,N_1054);
or U2535 (N_2535,N_746,N_1413);
and U2536 (N_2536,N_522,N_926);
nor U2537 (N_2537,N_417,N_1786);
nand U2538 (N_2538,N_1659,N_1820);
or U2539 (N_2539,N_1573,N_1166);
nand U2540 (N_2540,N_1211,N_1237);
xnor U2541 (N_2541,N_1791,N_787);
and U2542 (N_2542,N_730,N_559);
and U2543 (N_2543,N_1143,N_309);
or U2544 (N_2544,N_73,N_1487);
nand U2545 (N_2545,N_1304,N_668);
or U2546 (N_2546,N_897,N_1493);
and U2547 (N_2547,N_850,N_1765);
and U2548 (N_2548,N_720,N_1131);
nand U2549 (N_2549,N_1465,N_862);
nand U2550 (N_2550,N_1853,N_835);
nand U2551 (N_2551,N_600,N_989);
nor U2552 (N_2552,N_1175,N_392);
or U2553 (N_2553,N_1861,N_433);
and U2554 (N_2554,N_1906,N_100);
nor U2555 (N_2555,N_250,N_591);
or U2556 (N_2556,N_588,N_665);
xnor U2557 (N_2557,N_1746,N_257);
nor U2558 (N_2558,N_707,N_1144);
nor U2559 (N_2559,N_256,N_391);
and U2560 (N_2560,N_606,N_208);
and U2561 (N_2561,N_1318,N_714);
or U2562 (N_2562,N_682,N_447);
and U2563 (N_2563,N_1399,N_425);
nand U2564 (N_2564,N_343,N_631);
and U2565 (N_2565,N_692,N_679);
nand U2566 (N_2566,N_788,N_92);
nand U2567 (N_2567,N_259,N_235);
or U2568 (N_2568,N_405,N_535);
nand U2569 (N_2569,N_1338,N_1962);
or U2570 (N_2570,N_1822,N_1610);
nand U2571 (N_2571,N_1570,N_1945);
xor U2572 (N_2572,N_98,N_1837);
nor U2573 (N_2573,N_402,N_1694);
and U2574 (N_2574,N_546,N_1866);
or U2575 (N_2575,N_1604,N_390);
nand U2576 (N_2576,N_224,N_705);
nor U2577 (N_2577,N_1796,N_1170);
nand U2578 (N_2578,N_676,N_1894);
nand U2579 (N_2579,N_1540,N_121);
or U2580 (N_2580,N_783,N_276);
nand U2581 (N_2581,N_1308,N_920);
nor U2582 (N_2582,N_596,N_291);
or U2583 (N_2583,N_1592,N_1361);
or U2584 (N_2584,N_283,N_761);
and U2585 (N_2585,N_87,N_408);
nor U2586 (N_2586,N_1337,N_1193);
nand U2587 (N_2587,N_1717,N_469);
and U2588 (N_2588,N_1357,N_603);
nor U2589 (N_2589,N_1716,N_1346);
and U2590 (N_2590,N_1607,N_1045);
nor U2591 (N_2591,N_53,N_528);
and U2592 (N_2592,N_1392,N_310);
or U2593 (N_2593,N_1163,N_1420);
and U2594 (N_2594,N_1013,N_1431);
nor U2595 (N_2595,N_750,N_297);
nor U2596 (N_2596,N_1509,N_1909);
or U2597 (N_2597,N_657,N_650);
and U2598 (N_2598,N_992,N_1268);
nor U2599 (N_2599,N_963,N_166);
nand U2600 (N_2600,N_30,N_1276);
and U2601 (N_2601,N_184,N_1256);
or U2602 (N_2602,N_744,N_411);
or U2603 (N_2603,N_1675,N_1152);
nand U2604 (N_2604,N_1549,N_515);
nand U2605 (N_2605,N_1974,N_1950);
nor U2606 (N_2606,N_590,N_1932);
and U2607 (N_2607,N_625,N_1464);
nand U2608 (N_2608,N_481,N_1269);
nand U2609 (N_2609,N_810,N_1063);
and U2610 (N_2610,N_1902,N_1522);
nor U2611 (N_2611,N_1226,N_1266);
nor U2612 (N_2612,N_912,N_752);
and U2613 (N_2613,N_1759,N_1729);
and U2614 (N_2614,N_539,N_695);
nor U2615 (N_2615,N_168,N_1100);
nand U2616 (N_2616,N_1860,N_782);
and U2617 (N_2617,N_1782,N_1080);
or U2618 (N_2618,N_17,N_1944);
or U2619 (N_2619,N_1991,N_231);
nand U2620 (N_2620,N_903,N_1094);
nand U2621 (N_2621,N_574,N_577);
nor U2622 (N_2622,N_646,N_1971);
and U2623 (N_2623,N_728,N_544);
nor U2624 (N_2624,N_541,N_1865);
and U2625 (N_2625,N_1298,N_203);
nor U2626 (N_2626,N_226,N_845);
nor U2627 (N_2627,N_1104,N_357);
and U2628 (N_2628,N_1599,N_1884);
and U2629 (N_2629,N_355,N_479);
nor U2630 (N_2630,N_178,N_1983);
or U2631 (N_2631,N_1957,N_488);
nand U2632 (N_2632,N_1551,N_1418);
nand U2633 (N_2633,N_970,N_614);
xnor U2634 (N_2634,N_1767,N_0);
and U2635 (N_2635,N_324,N_1458);
or U2636 (N_2636,N_1998,N_1222);
nand U2637 (N_2637,N_1586,N_1500);
nor U2638 (N_2638,N_973,N_1812);
nor U2639 (N_2639,N_1324,N_1605);
and U2640 (N_2640,N_1496,N_399);
and U2641 (N_2641,N_685,N_1719);
or U2642 (N_2642,N_1379,N_1092);
nor U2643 (N_2643,N_1251,N_1481);
xor U2644 (N_2644,N_937,N_895);
and U2645 (N_2645,N_1603,N_1417);
and U2646 (N_2646,N_1452,N_240);
nand U2647 (N_2647,N_1696,N_1141);
or U2648 (N_2648,N_1136,N_430);
and U2649 (N_2649,N_1670,N_1238);
nand U2650 (N_2650,N_1351,N_632);
nand U2651 (N_2651,N_1097,N_472);
and U2652 (N_2652,N_91,N_608);
and U2653 (N_2653,N_478,N_75);
nand U2654 (N_2654,N_1560,N_582);
nor U2655 (N_2655,N_1565,N_1546);
or U2656 (N_2656,N_1926,N_1391);
nand U2657 (N_2657,N_253,N_1317);
nand U2658 (N_2658,N_1808,N_5);
and U2659 (N_2659,N_984,N_732);
and U2660 (N_2660,N_171,N_1541);
nand U2661 (N_2661,N_1930,N_1661);
nor U2662 (N_2662,N_889,N_1769);
or U2663 (N_2663,N_1984,N_266);
nand U2664 (N_2664,N_1697,N_747);
nor U2665 (N_2665,N_633,N_85);
nor U2666 (N_2666,N_1678,N_674);
and U2667 (N_2667,N_901,N_879);
nand U2668 (N_2668,N_902,N_90);
or U2669 (N_2669,N_1810,N_1074);
or U2670 (N_2670,N_228,N_435);
nand U2671 (N_2671,N_1151,N_1498);
and U2672 (N_2672,N_1985,N_721);
and U2673 (N_2673,N_282,N_525);
nor U2674 (N_2674,N_494,N_1735);
and U2675 (N_2675,N_1190,N_688);
or U2676 (N_2676,N_1771,N_660);
or U2677 (N_2677,N_47,N_1576);
nor U2678 (N_2678,N_578,N_398);
nand U2679 (N_2679,N_616,N_1872);
nor U2680 (N_2680,N_1363,N_1495);
or U2681 (N_2681,N_567,N_1378);
or U2682 (N_2682,N_1194,N_642);
or U2683 (N_2683,N_440,N_724);
or U2684 (N_2684,N_621,N_1595);
nand U2685 (N_2685,N_712,N_1515);
nand U2686 (N_2686,N_768,N_1478);
nor U2687 (N_2687,N_1839,N_140);
and U2688 (N_2688,N_1010,N_165);
and U2689 (N_2689,N_666,N_1686);
nand U2690 (N_2690,N_1118,N_24);
nor U2691 (N_2691,N_182,N_1557);
or U2692 (N_2692,N_916,N_763);
nand U2693 (N_2693,N_905,N_1721);
and U2694 (N_2694,N_766,N_1666);
nand U2695 (N_2695,N_475,N_290);
and U2696 (N_2696,N_1980,N_1457);
nor U2697 (N_2697,N_1313,N_239);
or U2698 (N_2698,N_1185,N_209);
and U2699 (N_2699,N_991,N_141);
or U2700 (N_2700,N_723,N_1693);
or U2701 (N_2701,N_1124,N_58);
or U2702 (N_2702,N_1908,N_1629);
nor U2703 (N_2703,N_1027,N_830);
and U2704 (N_2704,N_1823,N_458);
or U2705 (N_2705,N_1053,N_37);
nor U2706 (N_2706,N_1285,N_419);
nand U2707 (N_2707,N_814,N_1216);
and U2708 (N_2708,N_1105,N_1316);
nor U2709 (N_2709,N_71,N_1601);
nor U2710 (N_2710,N_1637,N_1875);
nor U2711 (N_2711,N_1524,N_410);
and U2712 (N_2712,N_1672,N_1044);
nand U2713 (N_2713,N_846,N_1445);
and U2714 (N_2714,N_866,N_1571);
nand U2715 (N_2715,N_1700,N_875);
or U2716 (N_2716,N_794,N_1982);
nand U2717 (N_2717,N_137,N_565);
nand U2718 (N_2718,N_1328,N_960);
or U2719 (N_2719,N_1479,N_837);
nor U2720 (N_2720,N_1460,N_1913);
and U2721 (N_2721,N_1245,N_1751);
nand U2722 (N_2722,N_1563,N_185);
nand U2723 (N_2723,N_464,N_938);
and U2724 (N_2724,N_1877,N_699);
nor U2725 (N_2725,N_521,N_449);
xnor U2726 (N_2726,N_1881,N_1293);
nor U2727 (N_2727,N_1360,N_1597);
or U2728 (N_2728,N_388,N_1085);
or U2729 (N_2729,N_1598,N_248);
nor U2730 (N_2730,N_563,N_1362);
or U2731 (N_2731,N_18,N_222);
and U2732 (N_2732,N_1486,N_1455);
nand U2733 (N_2733,N_1018,N_1017);
nor U2734 (N_2734,N_1815,N_349);
nor U2735 (N_2735,N_1380,N_1382);
or U2736 (N_2736,N_189,N_1959);
nor U2737 (N_2737,N_142,N_1912);
or U2738 (N_2738,N_369,N_1554);
nor U2739 (N_2739,N_448,N_1348);
and U2740 (N_2740,N_198,N_1920);
nand U2741 (N_2741,N_652,N_736);
or U2742 (N_2742,N_1718,N_594);
nand U2743 (N_2743,N_1441,N_474);
nor U2744 (N_2744,N_1743,N_1513);
nand U2745 (N_2745,N_1164,N_205);
or U2746 (N_2746,N_1662,N_89);
nor U2747 (N_2747,N_1199,N_1103);
nand U2748 (N_2748,N_1440,N_1367);
and U2749 (N_2749,N_1300,N_1814);
nand U2750 (N_2750,N_28,N_3);
nand U2751 (N_2751,N_1240,N_734);
and U2752 (N_2752,N_988,N_792);
and U2753 (N_2753,N_823,N_1307);
nand U2754 (N_2754,N_996,N_1213);
nor U2755 (N_2755,N_967,N_1544);
xor U2756 (N_2756,N_483,N_264);
nand U2757 (N_2757,N_964,N_1556);
or U2758 (N_2758,N_444,N_558);
and U2759 (N_2759,N_1408,N_1499);
and U2760 (N_2760,N_1819,N_1681);
or U2761 (N_2761,N_975,N_648);
xnor U2762 (N_2762,N_1949,N_376);
nor U2763 (N_2763,N_647,N_807);
or U2764 (N_2764,N_575,N_1600);
nor U2765 (N_2765,N_1504,N_941);
nand U2766 (N_2766,N_104,N_333);
and U2767 (N_2767,N_1528,N_1218);
nor U2768 (N_2768,N_966,N_1684);
nor U2769 (N_2769,N_1951,N_1349);
or U2770 (N_2770,N_1801,N_79);
nor U2771 (N_2771,N_1169,N_1828);
nor U2772 (N_2772,N_1370,N_1065);
nor U2773 (N_2773,N_88,N_461);
and U2774 (N_2774,N_1058,N_201);
nand U2775 (N_2775,N_1321,N_1521);
nand U2776 (N_2776,N_1731,N_215);
nor U2777 (N_2777,N_831,N_26);
or U2778 (N_2778,N_1037,N_197);
and U2779 (N_2779,N_384,N_1475);
and U2780 (N_2780,N_519,N_1915);
nand U2781 (N_2781,N_1254,N_1261);
nand U2782 (N_2782,N_1196,N_1415);
nor U2783 (N_2783,N_1271,N_572);
nand U2784 (N_2784,N_1365,N_1964);
nor U2785 (N_2785,N_764,N_1224);
or U2786 (N_2786,N_589,N_739);
nand U2787 (N_2787,N_1785,N_1548);
nand U2788 (N_2788,N_279,N_880);
nand U2789 (N_2789,N_1,N_1532);
or U2790 (N_2790,N_1423,N_70);
nand U2791 (N_2791,N_80,N_1852);
or U2792 (N_2792,N_1658,N_1102);
nand U2793 (N_2793,N_1161,N_687);
nor U2794 (N_2794,N_892,N_1878);
nand U2795 (N_2795,N_773,N_776);
or U2796 (N_2796,N_1483,N_990);
nand U2797 (N_2797,N_1309,N_936);
nand U2798 (N_2798,N_1220,N_864);
or U2799 (N_2799,N_1830,N_513);
or U2800 (N_2800,N_460,N_306);
nand U2801 (N_2801,N_38,N_1335);
and U2802 (N_2802,N_1792,N_865);
nand U2803 (N_2803,N_6,N_298);
or U2804 (N_2804,N_368,N_759);
nand U2805 (N_2805,N_268,N_146);
nor U2806 (N_2806,N_1035,N_1647);
nor U2807 (N_2807,N_1868,N_1142);
and U2808 (N_2808,N_1507,N_1806);
xor U2809 (N_2809,N_568,N_1303);
nor U2810 (N_2810,N_1381,N_672);
nand U2811 (N_2811,N_1802,N_1255);
nor U2812 (N_2812,N_1145,N_1162);
and U2813 (N_2813,N_717,N_351);
nor U2814 (N_2814,N_953,N_874);
nand U2815 (N_2815,N_1122,N_1685);
and U2816 (N_2816,N_1038,N_827);
or U2817 (N_2817,N_1292,N_1859);
nand U2818 (N_2818,N_1227,N_1990);
or U2819 (N_2819,N_278,N_1643);
or U2820 (N_2820,N_1733,N_1137);
or U2821 (N_2821,N_1703,N_1397);
nand U2822 (N_2822,N_251,N_1621);
or U2823 (N_2823,N_78,N_804);
nor U2824 (N_2824,N_762,N_1948);
nor U2825 (N_2825,N_1274,N_1147);
nand U2826 (N_2826,N_394,N_1726);
or U2827 (N_2827,N_543,N_1955);
nand U2828 (N_2828,N_1928,N_1234);
or U2829 (N_2829,N_1075,N_505);
and U2830 (N_2830,N_1813,N_1656);
nand U2831 (N_2831,N_455,N_414);
nor U2832 (N_2832,N_760,N_949);
nor U2833 (N_2833,N_396,N_870);
and U2834 (N_2834,N_1406,N_1975);
nand U2835 (N_2835,N_1247,N_1897);
and U2836 (N_2836,N_1747,N_199);
or U2837 (N_2837,N_1850,N_1738);
and U2838 (N_2838,N_1009,N_1069);
nor U2839 (N_2839,N_1757,N_856);
nor U2840 (N_2840,N_737,N_595);
nand U2841 (N_2841,N_489,N_2);
nor U2842 (N_2842,N_1129,N_930);
or U2843 (N_2843,N_907,N_626);
nor U2844 (N_2844,N_1588,N_1476);
and U2845 (N_2845,N_1836,N_1777);
nand U2846 (N_2846,N_295,N_957);
and U2847 (N_2847,N_1314,N_929);
and U2848 (N_2848,N_1425,N_1410);
nand U2849 (N_2849,N_1552,N_356);
or U2850 (N_2850,N_1691,N_1722);
and U2851 (N_2851,N_1299,N_161);
and U2852 (N_2852,N_29,N_733);
or U2853 (N_2853,N_1905,N_1940);
nor U2854 (N_2854,N_1312,N_1453);
nand U2855 (N_2855,N_354,N_1469);
nand U2856 (N_2856,N_81,N_663);
nand U2857 (N_2857,N_389,N_904);
or U2858 (N_2858,N_928,N_885);
nor U2859 (N_2859,N_1781,N_424);
nor U2860 (N_2860,N_1110,N_893);
and U2861 (N_2861,N_499,N_272);
or U2862 (N_2862,N_1167,N_273);
or U2863 (N_2863,N_1526,N_1177);
or U2864 (N_2864,N_661,N_55);
or U2865 (N_2865,N_1705,N_1039);
xor U2866 (N_2866,N_1130,N_1168);
nand U2867 (N_2867,N_1537,N_1388);
nor U2868 (N_2868,N_1611,N_700);
or U2869 (N_2869,N_913,N_1593);
nor U2870 (N_2870,N_729,N_1437);
nand U2871 (N_2871,N_453,N_1947);
or U2872 (N_2872,N_802,N_1645);
or U2873 (N_2873,N_1992,N_302);
nand U2874 (N_2874,N_54,N_491);
or U2875 (N_2875,N_681,N_1807);
nand U2876 (N_2876,N_952,N_1390);
and U2877 (N_2877,N_899,N_1262);
or U2878 (N_2878,N_553,N_1688);
nor U2879 (N_2879,N_1535,N_742);
or U2880 (N_2880,N_1432,N_1632);
nand U2881 (N_2881,N_1270,N_1900);
nor U2882 (N_2882,N_1282,N_1506);
nor U2883 (N_2883,N_842,N_1953);
nor U2884 (N_2884,N_386,N_139);
nand U2885 (N_2885,N_336,N_93);
nand U2886 (N_2886,N_1252,N_1385);
or U2887 (N_2887,N_1231,N_658);
nor U2888 (N_2888,N_1079,N_940);
and U2889 (N_2889,N_1301,N_691);
and U2890 (N_2890,N_1047,N_107);
nand U2891 (N_2891,N_318,N_1117);
and U2892 (N_2892,N_445,N_1081);
and U2893 (N_2893,N_858,N_1514);
nand U2894 (N_2894,N_1179,N_800);
or U2895 (N_2895,N_1650,N_1259);
and U2896 (N_2896,N_956,N_1652);
nand U2897 (N_2897,N_216,N_243);
or U2898 (N_2898,N_1536,N_797);
nor U2899 (N_2899,N_1155,N_1642);
or U2900 (N_2900,N_1438,N_339);
or U2901 (N_2901,N_1181,N_454);
nor U2902 (N_2902,N_82,N_46);
nand U2903 (N_2903,N_1368,N_1430);
or U2904 (N_2904,N_244,N_1120);
xor U2905 (N_2905,N_179,N_1280);
nand U2906 (N_2906,N_581,N_1290);
nor U2907 (N_2907,N_217,N_507);
nor U2908 (N_2908,N_1108,N_1333);
nor U2909 (N_2909,N_1692,N_34);
xor U2910 (N_2910,N_1209,N_337);
and U2911 (N_2911,N_367,N_452);
and U2912 (N_2912,N_1995,N_1623);
and U2913 (N_2913,N_172,N_236);
xnor U2914 (N_2914,N_1178,N_128);
nand U2915 (N_2915,N_164,N_1886);
nand U2916 (N_2916,N_307,N_891);
nor U2917 (N_2917,N_255,N_428);
or U2918 (N_2918,N_1756,N_1914);
nor U2919 (N_2919,N_1139,N_113);
nand U2920 (N_2920,N_1473,N_1195);
nand U2921 (N_2921,N_1972,N_1921);
or U2922 (N_2922,N_1527,N_149);
and U2923 (N_2923,N_701,N_638);
or U2924 (N_2924,N_1064,N_285);
and U2925 (N_2925,N_1530,N_35);
nor U2926 (N_2926,N_1516,N_1088);
or U2927 (N_2927,N_962,N_1029);
nand U2928 (N_2928,N_358,N_84);
nor U2929 (N_2929,N_372,N_847);
and U2930 (N_2930,N_612,N_1024);
or U2931 (N_2931,N_1428,N_523);
and U2932 (N_2932,N_506,N_418);
and U2933 (N_2933,N_815,N_1942);
and U2934 (N_2934,N_599,N_703);
or U2935 (N_2935,N_547,N_877);
nand U2936 (N_2936,N_1668,N_1727);
xor U2937 (N_2937,N_1034,N_246);
and U2938 (N_2938,N_977,N_275);
nor U2939 (N_2939,N_1664,N_780);
nand U2940 (N_2940,N_1480,N_781);
and U2941 (N_2941,N_549,N_1477);
and U2942 (N_2942,N_925,N_906);
nand U2943 (N_2943,N_111,N_1754);
nor U2944 (N_2944,N_1090,N_1794);
nand U2945 (N_2945,N_955,N_965);
nand U2946 (N_2946,N_134,N_416);
or U2947 (N_2947,N_1698,N_1903);
nand U2948 (N_2948,N_1518,N_709);
nand U2949 (N_2949,N_1284,N_1858);
or U2950 (N_2950,N_1864,N_1714);
and U2951 (N_2951,N_839,N_1999);
nand U2952 (N_2952,N_485,N_1246);
or U2953 (N_2953,N_649,N_527);
nand U2954 (N_2954,N_220,N_1294);
and U2955 (N_2955,N_420,N_1184);
nand U2956 (N_2956,N_1543,N_335);
and U2957 (N_2957,N_379,N_1462);
and U2958 (N_2958,N_883,N_751);
and U2959 (N_2959,N_1359,N_745);
or U2960 (N_2960,N_785,N_1305);
nor U2961 (N_2961,N_1699,N_1345);
and U2962 (N_2962,N_1235,N_116);
and U2963 (N_2963,N_1923,N_1941);
nor U2964 (N_2964,N_1648,N_1834);
nor U2965 (N_2965,N_1895,N_1429);
nor U2966 (N_2966,N_1414,N_520);
or U2967 (N_2967,N_1258,N_968);
or U2968 (N_2968,N_223,N_976);
xor U2969 (N_2969,N_1725,N_1158);
and U2970 (N_2970,N_1061,N_363);
nor U2971 (N_2971,N_1608,N_1154);
and U2972 (N_2972,N_1005,N_935);
nor U2973 (N_2973,N_1748,N_716);
or U2974 (N_2974,N_1119,N_1898);
nand U2975 (N_2975,N_66,N_1150);
or U2976 (N_2976,N_1225,N_352);
nand U2977 (N_2977,N_731,N_332);
and U2978 (N_2978,N_1113,N_698);
or U2979 (N_2979,N_1976,N_1846);
and U2980 (N_2980,N_586,N_1730);
nor U2981 (N_2981,N_1904,N_1214);
nand U2982 (N_2982,N_656,N_635);
nor U2983 (N_2983,N_1712,N_1401);
nand U2984 (N_2984,N_1404,N_1329);
and U2985 (N_2985,N_1078,N_8);
nand U2986 (N_2986,N_526,N_270);
or U2987 (N_2987,N_212,N_1963);
nor U2988 (N_2988,N_1032,N_1646);
and U2989 (N_2989,N_1416,N_1197);
nor U2990 (N_2990,N_1267,N_1442);
xor U2991 (N_2991,N_183,N_645);
nor U2992 (N_2992,N_1967,N_602);
and U2993 (N_2993,N_465,N_280);
nand U2994 (N_2994,N_884,N_1737);
nor U2995 (N_2995,N_274,N_943);
nand U2996 (N_2996,N_1505,N_758);
nor U2997 (N_2997,N_1583,N_1071);
nor U2998 (N_2998,N_254,N_347);
or U2999 (N_2999,N_1870,N_1123);
nor U3000 (N_3000,N_873,N_1572);
nor U3001 (N_3001,N_1250,N_943);
or U3002 (N_3002,N_1370,N_429);
nor U3003 (N_3003,N_89,N_1997);
nand U3004 (N_3004,N_39,N_57);
and U3005 (N_3005,N_201,N_1057);
nand U3006 (N_3006,N_150,N_932);
or U3007 (N_3007,N_1750,N_991);
or U3008 (N_3008,N_971,N_889);
and U3009 (N_3009,N_140,N_1313);
nand U3010 (N_3010,N_322,N_202);
nand U3011 (N_3011,N_915,N_325);
nor U3012 (N_3012,N_1372,N_688);
nand U3013 (N_3013,N_1465,N_447);
or U3014 (N_3014,N_1189,N_1985);
and U3015 (N_3015,N_941,N_1125);
or U3016 (N_3016,N_1742,N_61);
or U3017 (N_3017,N_1185,N_318);
nand U3018 (N_3018,N_1853,N_386);
nand U3019 (N_3019,N_1332,N_1945);
or U3020 (N_3020,N_1360,N_1102);
and U3021 (N_3021,N_886,N_1091);
nand U3022 (N_3022,N_1273,N_217);
nor U3023 (N_3023,N_129,N_686);
and U3024 (N_3024,N_1269,N_1545);
and U3025 (N_3025,N_1208,N_1512);
and U3026 (N_3026,N_1272,N_1010);
nand U3027 (N_3027,N_1826,N_1024);
or U3028 (N_3028,N_1555,N_355);
nor U3029 (N_3029,N_878,N_202);
nand U3030 (N_3030,N_558,N_1936);
nand U3031 (N_3031,N_1,N_320);
nand U3032 (N_3032,N_957,N_1475);
nor U3033 (N_3033,N_1901,N_229);
nor U3034 (N_3034,N_206,N_909);
and U3035 (N_3035,N_1897,N_177);
and U3036 (N_3036,N_1222,N_822);
nor U3037 (N_3037,N_1683,N_1014);
nand U3038 (N_3038,N_868,N_1239);
nor U3039 (N_3039,N_1639,N_628);
or U3040 (N_3040,N_1940,N_724);
nor U3041 (N_3041,N_1930,N_855);
nand U3042 (N_3042,N_564,N_1164);
or U3043 (N_3043,N_65,N_993);
or U3044 (N_3044,N_1632,N_648);
xnor U3045 (N_3045,N_1131,N_358);
or U3046 (N_3046,N_1148,N_1829);
and U3047 (N_3047,N_1641,N_1593);
nand U3048 (N_3048,N_928,N_487);
and U3049 (N_3049,N_1924,N_879);
nand U3050 (N_3050,N_1543,N_1242);
nand U3051 (N_3051,N_383,N_1393);
or U3052 (N_3052,N_509,N_319);
nand U3053 (N_3053,N_55,N_200);
or U3054 (N_3054,N_1628,N_1243);
and U3055 (N_3055,N_746,N_1087);
nor U3056 (N_3056,N_484,N_649);
xor U3057 (N_3057,N_1174,N_1707);
nor U3058 (N_3058,N_1167,N_1958);
nor U3059 (N_3059,N_1266,N_1830);
nand U3060 (N_3060,N_100,N_1384);
nand U3061 (N_3061,N_1946,N_442);
nand U3062 (N_3062,N_693,N_226);
or U3063 (N_3063,N_1166,N_1812);
or U3064 (N_3064,N_544,N_1318);
and U3065 (N_3065,N_804,N_1423);
nor U3066 (N_3066,N_1358,N_91);
and U3067 (N_3067,N_1079,N_1214);
nand U3068 (N_3068,N_1429,N_102);
or U3069 (N_3069,N_385,N_1691);
nand U3070 (N_3070,N_1699,N_658);
or U3071 (N_3071,N_911,N_1741);
nand U3072 (N_3072,N_309,N_150);
nor U3073 (N_3073,N_1088,N_1659);
or U3074 (N_3074,N_7,N_1543);
and U3075 (N_3075,N_787,N_1977);
nor U3076 (N_3076,N_300,N_545);
or U3077 (N_3077,N_1784,N_556);
nor U3078 (N_3078,N_931,N_854);
and U3079 (N_3079,N_1599,N_1140);
nand U3080 (N_3080,N_1118,N_1467);
nand U3081 (N_3081,N_811,N_1156);
or U3082 (N_3082,N_1800,N_880);
or U3083 (N_3083,N_194,N_1141);
nand U3084 (N_3084,N_1401,N_1066);
or U3085 (N_3085,N_1251,N_10);
and U3086 (N_3086,N_1385,N_1111);
nand U3087 (N_3087,N_1577,N_105);
or U3088 (N_3088,N_122,N_293);
nand U3089 (N_3089,N_875,N_1216);
and U3090 (N_3090,N_1163,N_1241);
or U3091 (N_3091,N_469,N_1273);
nor U3092 (N_3092,N_561,N_130);
nor U3093 (N_3093,N_353,N_1648);
nand U3094 (N_3094,N_1648,N_26);
and U3095 (N_3095,N_1652,N_1501);
or U3096 (N_3096,N_1966,N_60);
nand U3097 (N_3097,N_1894,N_1607);
or U3098 (N_3098,N_974,N_341);
nor U3099 (N_3099,N_692,N_172);
nand U3100 (N_3100,N_84,N_1280);
nand U3101 (N_3101,N_738,N_140);
nand U3102 (N_3102,N_1609,N_1405);
nor U3103 (N_3103,N_1652,N_1756);
and U3104 (N_3104,N_1567,N_140);
and U3105 (N_3105,N_59,N_1414);
and U3106 (N_3106,N_650,N_109);
nor U3107 (N_3107,N_1400,N_1283);
nand U3108 (N_3108,N_205,N_1370);
nand U3109 (N_3109,N_12,N_1321);
or U3110 (N_3110,N_213,N_1481);
or U3111 (N_3111,N_1954,N_1872);
or U3112 (N_3112,N_1772,N_1765);
nand U3113 (N_3113,N_1708,N_1713);
nor U3114 (N_3114,N_1278,N_1305);
nand U3115 (N_3115,N_1895,N_1032);
nor U3116 (N_3116,N_1893,N_177);
nor U3117 (N_3117,N_500,N_83);
or U3118 (N_3118,N_1758,N_228);
nor U3119 (N_3119,N_1057,N_1219);
and U3120 (N_3120,N_21,N_745);
or U3121 (N_3121,N_1551,N_1828);
or U3122 (N_3122,N_839,N_897);
and U3123 (N_3123,N_367,N_979);
and U3124 (N_3124,N_775,N_1301);
nor U3125 (N_3125,N_1831,N_1288);
or U3126 (N_3126,N_360,N_225);
and U3127 (N_3127,N_417,N_1843);
and U3128 (N_3128,N_286,N_215);
nor U3129 (N_3129,N_1677,N_285);
nand U3130 (N_3130,N_1271,N_1280);
nor U3131 (N_3131,N_1566,N_735);
nor U3132 (N_3132,N_1803,N_512);
and U3133 (N_3133,N_277,N_1389);
or U3134 (N_3134,N_1605,N_1492);
and U3135 (N_3135,N_704,N_717);
nor U3136 (N_3136,N_1833,N_1398);
and U3137 (N_3137,N_881,N_389);
nor U3138 (N_3138,N_1757,N_1861);
xnor U3139 (N_3139,N_1761,N_167);
or U3140 (N_3140,N_1516,N_182);
nand U3141 (N_3141,N_1061,N_544);
or U3142 (N_3142,N_569,N_7);
nand U3143 (N_3143,N_1443,N_1731);
nand U3144 (N_3144,N_1377,N_1069);
or U3145 (N_3145,N_787,N_1165);
or U3146 (N_3146,N_411,N_1146);
or U3147 (N_3147,N_1209,N_279);
nand U3148 (N_3148,N_1779,N_296);
or U3149 (N_3149,N_486,N_1212);
and U3150 (N_3150,N_560,N_1085);
nand U3151 (N_3151,N_1401,N_345);
nor U3152 (N_3152,N_1326,N_1423);
nor U3153 (N_3153,N_434,N_786);
nand U3154 (N_3154,N_1376,N_1961);
or U3155 (N_3155,N_720,N_347);
and U3156 (N_3156,N_232,N_1489);
nor U3157 (N_3157,N_1837,N_153);
nor U3158 (N_3158,N_1418,N_770);
nor U3159 (N_3159,N_1412,N_993);
nand U3160 (N_3160,N_139,N_1288);
nor U3161 (N_3161,N_1095,N_1921);
nand U3162 (N_3162,N_384,N_1975);
and U3163 (N_3163,N_1069,N_1133);
nor U3164 (N_3164,N_1746,N_1340);
nor U3165 (N_3165,N_1930,N_331);
nor U3166 (N_3166,N_243,N_1585);
xor U3167 (N_3167,N_917,N_386);
nor U3168 (N_3168,N_603,N_1150);
nand U3169 (N_3169,N_1432,N_788);
nand U3170 (N_3170,N_490,N_1891);
and U3171 (N_3171,N_1055,N_799);
and U3172 (N_3172,N_1663,N_609);
and U3173 (N_3173,N_731,N_1520);
nor U3174 (N_3174,N_670,N_1878);
nor U3175 (N_3175,N_250,N_15);
nor U3176 (N_3176,N_806,N_286);
nor U3177 (N_3177,N_1517,N_1234);
or U3178 (N_3178,N_1419,N_212);
or U3179 (N_3179,N_1845,N_1785);
nand U3180 (N_3180,N_1124,N_223);
and U3181 (N_3181,N_292,N_373);
nor U3182 (N_3182,N_1506,N_1132);
nor U3183 (N_3183,N_1489,N_1028);
nand U3184 (N_3184,N_1044,N_1639);
nand U3185 (N_3185,N_1036,N_606);
and U3186 (N_3186,N_1036,N_1190);
or U3187 (N_3187,N_1740,N_1143);
or U3188 (N_3188,N_1960,N_1681);
or U3189 (N_3189,N_1543,N_1082);
nor U3190 (N_3190,N_1134,N_153);
xnor U3191 (N_3191,N_975,N_336);
and U3192 (N_3192,N_358,N_1464);
nor U3193 (N_3193,N_169,N_1008);
or U3194 (N_3194,N_929,N_760);
and U3195 (N_3195,N_474,N_624);
and U3196 (N_3196,N_1510,N_70);
and U3197 (N_3197,N_849,N_1542);
and U3198 (N_3198,N_1288,N_389);
nand U3199 (N_3199,N_1898,N_270);
or U3200 (N_3200,N_1214,N_1384);
and U3201 (N_3201,N_530,N_402);
or U3202 (N_3202,N_794,N_919);
nor U3203 (N_3203,N_1681,N_391);
nand U3204 (N_3204,N_378,N_1081);
nor U3205 (N_3205,N_1067,N_1208);
or U3206 (N_3206,N_1972,N_579);
or U3207 (N_3207,N_279,N_1042);
or U3208 (N_3208,N_856,N_1713);
nand U3209 (N_3209,N_1858,N_246);
and U3210 (N_3210,N_463,N_1660);
and U3211 (N_3211,N_1813,N_837);
nor U3212 (N_3212,N_1068,N_374);
and U3213 (N_3213,N_1447,N_642);
or U3214 (N_3214,N_1332,N_1435);
and U3215 (N_3215,N_300,N_1102);
nand U3216 (N_3216,N_1198,N_322);
and U3217 (N_3217,N_1083,N_807);
or U3218 (N_3218,N_531,N_576);
and U3219 (N_3219,N_107,N_1555);
or U3220 (N_3220,N_559,N_632);
and U3221 (N_3221,N_1376,N_1766);
nand U3222 (N_3222,N_1128,N_1986);
and U3223 (N_3223,N_422,N_1193);
or U3224 (N_3224,N_1653,N_69);
or U3225 (N_3225,N_181,N_817);
xor U3226 (N_3226,N_1894,N_1188);
or U3227 (N_3227,N_1702,N_100);
nor U3228 (N_3228,N_244,N_1478);
nand U3229 (N_3229,N_1208,N_1174);
or U3230 (N_3230,N_346,N_1596);
or U3231 (N_3231,N_349,N_1061);
nor U3232 (N_3232,N_355,N_1091);
xor U3233 (N_3233,N_1691,N_1148);
and U3234 (N_3234,N_1546,N_864);
nand U3235 (N_3235,N_960,N_862);
nor U3236 (N_3236,N_1400,N_595);
and U3237 (N_3237,N_1055,N_776);
and U3238 (N_3238,N_1489,N_1098);
nor U3239 (N_3239,N_1417,N_1141);
nor U3240 (N_3240,N_119,N_1423);
nor U3241 (N_3241,N_1378,N_1769);
or U3242 (N_3242,N_1789,N_1908);
and U3243 (N_3243,N_181,N_1364);
or U3244 (N_3244,N_566,N_1561);
nand U3245 (N_3245,N_631,N_620);
and U3246 (N_3246,N_1529,N_1361);
nor U3247 (N_3247,N_0,N_490);
or U3248 (N_3248,N_365,N_145);
and U3249 (N_3249,N_1330,N_800);
nor U3250 (N_3250,N_816,N_1007);
nor U3251 (N_3251,N_1714,N_1220);
nor U3252 (N_3252,N_1240,N_1198);
or U3253 (N_3253,N_125,N_1325);
and U3254 (N_3254,N_346,N_1901);
and U3255 (N_3255,N_1266,N_19);
nand U3256 (N_3256,N_1075,N_1025);
nor U3257 (N_3257,N_191,N_1208);
or U3258 (N_3258,N_131,N_190);
nor U3259 (N_3259,N_1269,N_587);
nor U3260 (N_3260,N_311,N_1809);
nand U3261 (N_3261,N_1688,N_174);
and U3262 (N_3262,N_365,N_327);
nand U3263 (N_3263,N_746,N_912);
nor U3264 (N_3264,N_1473,N_294);
nand U3265 (N_3265,N_817,N_1917);
or U3266 (N_3266,N_374,N_649);
and U3267 (N_3267,N_336,N_1581);
nand U3268 (N_3268,N_1068,N_795);
and U3269 (N_3269,N_424,N_29);
and U3270 (N_3270,N_280,N_1484);
nand U3271 (N_3271,N_399,N_707);
and U3272 (N_3272,N_1881,N_238);
and U3273 (N_3273,N_681,N_1180);
or U3274 (N_3274,N_57,N_753);
nand U3275 (N_3275,N_415,N_1550);
nand U3276 (N_3276,N_119,N_28);
nor U3277 (N_3277,N_403,N_81);
and U3278 (N_3278,N_46,N_2);
nand U3279 (N_3279,N_1663,N_789);
nand U3280 (N_3280,N_1719,N_848);
xor U3281 (N_3281,N_1864,N_415);
or U3282 (N_3282,N_1439,N_212);
or U3283 (N_3283,N_2,N_1133);
and U3284 (N_3284,N_31,N_653);
and U3285 (N_3285,N_713,N_1370);
or U3286 (N_3286,N_1329,N_383);
nand U3287 (N_3287,N_1158,N_1643);
or U3288 (N_3288,N_1648,N_1503);
nand U3289 (N_3289,N_434,N_970);
nor U3290 (N_3290,N_416,N_1774);
or U3291 (N_3291,N_209,N_1193);
and U3292 (N_3292,N_1801,N_1626);
nand U3293 (N_3293,N_1056,N_136);
and U3294 (N_3294,N_462,N_938);
nor U3295 (N_3295,N_1366,N_1611);
nor U3296 (N_3296,N_1038,N_422);
or U3297 (N_3297,N_867,N_1938);
nor U3298 (N_3298,N_990,N_734);
nand U3299 (N_3299,N_807,N_1128);
or U3300 (N_3300,N_746,N_374);
or U3301 (N_3301,N_1824,N_1309);
or U3302 (N_3302,N_1262,N_952);
or U3303 (N_3303,N_425,N_557);
or U3304 (N_3304,N_541,N_1515);
nor U3305 (N_3305,N_1437,N_468);
xnor U3306 (N_3306,N_479,N_752);
and U3307 (N_3307,N_1801,N_897);
nand U3308 (N_3308,N_1216,N_1376);
and U3309 (N_3309,N_1518,N_1725);
nor U3310 (N_3310,N_1644,N_684);
nor U3311 (N_3311,N_1979,N_1757);
and U3312 (N_3312,N_335,N_342);
and U3313 (N_3313,N_623,N_1573);
and U3314 (N_3314,N_534,N_1169);
or U3315 (N_3315,N_116,N_1117);
nand U3316 (N_3316,N_1996,N_1926);
or U3317 (N_3317,N_1668,N_1239);
nand U3318 (N_3318,N_1908,N_989);
and U3319 (N_3319,N_997,N_1285);
xor U3320 (N_3320,N_46,N_519);
nor U3321 (N_3321,N_80,N_772);
nor U3322 (N_3322,N_258,N_822);
and U3323 (N_3323,N_925,N_1967);
nor U3324 (N_3324,N_160,N_743);
or U3325 (N_3325,N_1102,N_678);
nor U3326 (N_3326,N_1591,N_1559);
nand U3327 (N_3327,N_43,N_1280);
and U3328 (N_3328,N_513,N_334);
or U3329 (N_3329,N_625,N_457);
and U3330 (N_3330,N_1825,N_1748);
or U3331 (N_3331,N_1022,N_783);
nor U3332 (N_3332,N_501,N_1825);
and U3333 (N_3333,N_437,N_59);
nor U3334 (N_3334,N_1273,N_1947);
or U3335 (N_3335,N_422,N_1015);
and U3336 (N_3336,N_63,N_323);
xor U3337 (N_3337,N_1082,N_1713);
nand U3338 (N_3338,N_549,N_679);
nand U3339 (N_3339,N_417,N_1121);
and U3340 (N_3340,N_1125,N_1838);
and U3341 (N_3341,N_1314,N_989);
and U3342 (N_3342,N_1368,N_1183);
or U3343 (N_3343,N_568,N_1663);
or U3344 (N_3344,N_1244,N_622);
and U3345 (N_3345,N_1974,N_1661);
nand U3346 (N_3346,N_862,N_1851);
or U3347 (N_3347,N_1866,N_690);
and U3348 (N_3348,N_1439,N_141);
nor U3349 (N_3349,N_1892,N_691);
or U3350 (N_3350,N_511,N_1778);
nor U3351 (N_3351,N_1734,N_105);
or U3352 (N_3352,N_1139,N_1833);
nand U3353 (N_3353,N_419,N_1326);
nand U3354 (N_3354,N_1,N_1390);
and U3355 (N_3355,N_1748,N_314);
nor U3356 (N_3356,N_1896,N_1359);
nand U3357 (N_3357,N_1731,N_1789);
nand U3358 (N_3358,N_1026,N_1741);
nor U3359 (N_3359,N_884,N_354);
and U3360 (N_3360,N_91,N_1994);
and U3361 (N_3361,N_1826,N_1034);
nand U3362 (N_3362,N_254,N_330);
nor U3363 (N_3363,N_829,N_1681);
nand U3364 (N_3364,N_289,N_1906);
and U3365 (N_3365,N_1030,N_1967);
nand U3366 (N_3366,N_1977,N_984);
and U3367 (N_3367,N_570,N_1332);
and U3368 (N_3368,N_590,N_376);
xnor U3369 (N_3369,N_660,N_1990);
nand U3370 (N_3370,N_1116,N_1483);
nor U3371 (N_3371,N_490,N_1537);
nand U3372 (N_3372,N_1603,N_1880);
or U3373 (N_3373,N_841,N_1056);
nor U3374 (N_3374,N_1674,N_1401);
and U3375 (N_3375,N_1914,N_694);
nor U3376 (N_3376,N_261,N_1949);
and U3377 (N_3377,N_639,N_696);
nor U3378 (N_3378,N_382,N_1550);
nand U3379 (N_3379,N_496,N_999);
nand U3380 (N_3380,N_1495,N_1827);
and U3381 (N_3381,N_665,N_773);
and U3382 (N_3382,N_1433,N_736);
or U3383 (N_3383,N_946,N_1668);
or U3384 (N_3384,N_1883,N_1105);
nor U3385 (N_3385,N_1503,N_1620);
xor U3386 (N_3386,N_1868,N_953);
or U3387 (N_3387,N_635,N_565);
nor U3388 (N_3388,N_1772,N_1838);
and U3389 (N_3389,N_1628,N_1608);
nor U3390 (N_3390,N_1622,N_888);
and U3391 (N_3391,N_525,N_997);
or U3392 (N_3392,N_1997,N_597);
nor U3393 (N_3393,N_1157,N_776);
and U3394 (N_3394,N_159,N_3);
and U3395 (N_3395,N_1708,N_1914);
and U3396 (N_3396,N_746,N_868);
nor U3397 (N_3397,N_1498,N_1327);
nor U3398 (N_3398,N_323,N_1351);
nand U3399 (N_3399,N_1824,N_1960);
and U3400 (N_3400,N_138,N_847);
or U3401 (N_3401,N_1106,N_909);
nand U3402 (N_3402,N_1395,N_1377);
and U3403 (N_3403,N_1445,N_477);
and U3404 (N_3404,N_95,N_760);
nor U3405 (N_3405,N_802,N_1507);
nor U3406 (N_3406,N_567,N_832);
or U3407 (N_3407,N_100,N_693);
or U3408 (N_3408,N_1330,N_952);
and U3409 (N_3409,N_181,N_1141);
nor U3410 (N_3410,N_1508,N_1859);
and U3411 (N_3411,N_1158,N_1611);
and U3412 (N_3412,N_806,N_1781);
and U3413 (N_3413,N_1865,N_1003);
nor U3414 (N_3414,N_959,N_765);
nor U3415 (N_3415,N_1842,N_397);
and U3416 (N_3416,N_676,N_1311);
and U3417 (N_3417,N_990,N_561);
and U3418 (N_3418,N_898,N_1396);
nor U3419 (N_3419,N_1236,N_397);
and U3420 (N_3420,N_843,N_534);
nor U3421 (N_3421,N_711,N_1929);
nand U3422 (N_3422,N_534,N_1723);
nor U3423 (N_3423,N_1544,N_1829);
and U3424 (N_3424,N_727,N_1315);
or U3425 (N_3425,N_720,N_80);
or U3426 (N_3426,N_660,N_811);
nand U3427 (N_3427,N_1261,N_1898);
nand U3428 (N_3428,N_3,N_678);
nand U3429 (N_3429,N_74,N_1337);
or U3430 (N_3430,N_997,N_243);
and U3431 (N_3431,N_23,N_1180);
nand U3432 (N_3432,N_206,N_724);
or U3433 (N_3433,N_809,N_77);
nand U3434 (N_3434,N_1323,N_1106);
or U3435 (N_3435,N_529,N_1627);
and U3436 (N_3436,N_1103,N_1390);
or U3437 (N_3437,N_1862,N_1782);
nand U3438 (N_3438,N_1852,N_912);
or U3439 (N_3439,N_355,N_1462);
and U3440 (N_3440,N_844,N_87);
and U3441 (N_3441,N_1224,N_269);
nand U3442 (N_3442,N_32,N_1657);
and U3443 (N_3443,N_1608,N_914);
nor U3444 (N_3444,N_11,N_1349);
nand U3445 (N_3445,N_1480,N_1);
nand U3446 (N_3446,N_1263,N_468);
and U3447 (N_3447,N_651,N_1947);
and U3448 (N_3448,N_1737,N_544);
or U3449 (N_3449,N_549,N_1311);
nor U3450 (N_3450,N_338,N_120);
or U3451 (N_3451,N_1685,N_1740);
or U3452 (N_3452,N_892,N_543);
or U3453 (N_3453,N_101,N_878);
or U3454 (N_3454,N_453,N_1896);
or U3455 (N_3455,N_470,N_316);
nor U3456 (N_3456,N_961,N_1097);
nor U3457 (N_3457,N_1420,N_39);
and U3458 (N_3458,N_152,N_720);
nor U3459 (N_3459,N_135,N_1312);
nand U3460 (N_3460,N_101,N_19);
xor U3461 (N_3461,N_1308,N_1335);
nor U3462 (N_3462,N_517,N_160);
or U3463 (N_3463,N_32,N_506);
and U3464 (N_3464,N_475,N_291);
nor U3465 (N_3465,N_229,N_863);
nor U3466 (N_3466,N_1475,N_1721);
nand U3467 (N_3467,N_1169,N_620);
nand U3468 (N_3468,N_1287,N_1319);
nand U3469 (N_3469,N_1783,N_1930);
or U3470 (N_3470,N_497,N_310);
or U3471 (N_3471,N_240,N_1338);
and U3472 (N_3472,N_406,N_1250);
or U3473 (N_3473,N_580,N_1312);
and U3474 (N_3474,N_254,N_152);
xnor U3475 (N_3475,N_1347,N_1894);
nor U3476 (N_3476,N_32,N_1988);
nand U3477 (N_3477,N_1637,N_639);
or U3478 (N_3478,N_1154,N_1566);
xnor U3479 (N_3479,N_1906,N_1000);
or U3480 (N_3480,N_192,N_0);
nor U3481 (N_3481,N_323,N_1168);
or U3482 (N_3482,N_1697,N_1013);
and U3483 (N_3483,N_607,N_1534);
and U3484 (N_3484,N_1291,N_1854);
nor U3485 (N_3485,N_328,N_1465);
or U3486 (N_3486,N_1565,N_63);
nor U3487 (N_3487,N_1487,N_27);
and U3488 (N_3488,N_535,N_1189);
nor U3489 (N_3489,N_1719,N_188);
or U3490 (N_3490,N_531,N_1754);
or U3491 (N_3491,N_782,N_488);
and U3492 (N_3492,N_523,N_428);
and U3493 (N_3493,N_1481,N_445);
and U3494 (N_3494,N_1446,N_889);
or U3495 (N_3495,N_536,N_129);
nor U3496 (N_3496,N_1499,N_61);
or U3497 (N_3497,N_13,N_263);
nand U3498 (N_3498,N_466,N_822);
and U3499 (N_3499,N_390,N_498);
and U3500 (N_3500,N_1543,N_772);
nand U3501 (N_3501,N_1157,N_228);
nor U3502 (N_3502,N_1423,N_1327);
and U3503 (N_3503,N_1103,N_1635);
nand U3504 (N_3504,N_155,N_231);
nor U3505 (N_3505,N_1973,N_438);
and U3506 (N_3506,N_1659,N_689);
or U3507 (N_3507,N_1585,N_276);
or U3508 (N_3508,N_430,N_1799);
nand U3509 (N_3509,N_175,N_1621);
or U3510 (N_3510,N_1543,N_1114);
nor U3511 (N_3511,N_357,N_1242);
nand U3512 (N_3512,N_526,N_253);
nor U3513 (N_3513,N_149,N_1671);
nand U3514 (N_3514,N_349,N_699);
nand U3515 (N_3515,N_248,N_1660);
or U3516 (N_3516,N_1631,N_562);
and U3517 (N_3517,N_1945,N_382);
or U3518 (N_3518,N_1266,N_1373);
and U3519 (N_3519,N_1678,N_377);
nand U3520 (N_3520,N_273,N_1432);
nor U3521 (N_3521,N_384,N_1749);
or U3522 (N_3522,N_1690,N_1094);
nand U3523 (N_3523,N_1026,N_1410);
and U3524 (N_3524,N_484,N_354);
nor U3525 (N_3525,N_422,N_1832);
nor U3526 (N_3526,N_575,N_1843);
nand U3527 (N_3527,N_1621,N_1696);
and U3528 (N_3528,N_904,N_401);
or U3529 (N_3529,N_1299,N_17);
nand U3530 (N_3530,N_949,N_660);
and U3531 (N_3531,N_1903,N_993);
nand U3532 (N_3532,N_858,N_1873);
nand U3533 (N_3533,N_326,N_536);
and U3534 (N_3534,N_877,N_211);
nand U3535 (N_3535,N_1733,N_1214);
nand U3536 (N_3536,N_791,N_1646);
and U3537 (N_3537,N_836,N_651);
nor U3538 (N_3538,N_1701,N_254);
nor U3539 (N_3539,N_1781,N_1942);
or U3540 (N_3540,N_910,N_1379);
and U3541 (N_3541,N_1083,N_1534);
and U3542 (N_3542,N_1408,N_1173);
or U3543 (N_3543,N_1288,N_1849);
nor U3544 (N_3544,N_1471,N_565);
or U3545 (N_3545,N_886,N_1869);
nor U3546 (N_3546,N_678,N_9);
nand U3547 (N_3547,N_900,N_1435);
xor U3548 (N_3548,N_1691,N_1132);
nor U3549 (N_3549,N_750,N_636);
nand U3550 (N_3550,N_1813,N_1816);
nor U3551 (N_3551,N_1988,N_30);
or U3552 (N_3552,N_736,N_370);
or U3553 (N_3553,N_1706,N_254);
and U3554 (N_3554,N_691,N_1420);
or U3555 (N_3555,N_1008,N_1266);
nand U3556 (N_3556,N_996,N_136);
and U3557 (N_3557,N_1959,N_1039);
and U3558 (N_3558,N_1669,N_278);
or U3559 (N_3559,N_1967,N_1669);
or U3560 (N_3560,N_392,N_26);
nand U3561 (N_3561,N_1166,N_585);
xnor U3562 (N_3562,N_1425,N_1460);
or U3563 (N_3563,N_619,N_90);
and U3564 (N_3564,N_493,N_1442);
nor U3565 (N_3565,N_1867,N_455);
and U3566 (N_3566,N_427,N_1120);
or U3567 (N_3567,N_1443,N_956);
and U3568 (N_3568,N_1918,N_1428);
nand U3569 (N_3569,N_773,N_372);
nand U3570 (N_3570,N_673,N_724);
nand U3571 (N_3571,N_481,N_1722);
or U3572 (N_3572,N_1597,N_690);
nor U3573 (N_3573,N_1939,N_898);
nand U3574 (N_3574,N_1448,N_863);
nand U3575 (N_3575,N_851,N_1757);
or U3576 (N_3576,N_250,N_582);
nand U3577 (N_3577,N_1165,N_1002);
or U3578 (N_3578,N_1242,N_52);
or U3579 (N_3579,N_1722,N_1048);
or U3580 (N_3580,N_731,N_289);
and U3581 (N_3581,N_864,N_1086);
nor U3582 (N_3582,N_75,N_324);
nor U3583 (N_3583,N_1156,N_234);
or U3584 (N_3584,N_890,N_1050);
or U3585 (N_3585,N_1807,N_1535);
or U3586 (N_3586,N_1813,N_649);
or U3587 (N_3587,N_207,N_965);
or U3588 (N_3588,N_1702,N_812);
and U3589 (N_3589,N_1290,N_445);
nand U3590 (N_3590,N_1160,N_605);
or U3591 (N_3591,N_794,N_1669);
nand U3592 (N_3592,N_1901,N_1548);
or U3593 (N_3593,N_1503,N_700);
or U3594 (N_3594,N_1708,N_616);
nor U3595 (N_3595,N_755,N_1030);
and U3596 (N_3596,N_630,N_1914);
nand U3597 (N_3597,N_1167,N_1648);
nand U3598 (N_3598,N_391,N_548);
nand U3599 (N_3599,N_670,N_368);
and U3600 (N_3600,N_274,N_1519);
and U3601 (N_3601,N_168,N_828);
and U3602 (N_3602,N_1295,N_165);
or U3603 (N_3603,N_200,N_1142);
or U3604 (N_3604,N_1945,N_1745);
nand U3605 (N_3605,N_99,N_1957);
and U3606 (N_3606,N_1298,N_1076);
and U3607 (N_3607,N_1934,N_487);
nor U3608 (N_3608,N_873,N_691);
nor U3609 (N_3609,N_1783,N_1377);
or U3610 (N_3610,N_1627,N_1675);
nor U3611 (N_3611,N_1895,N_1501);
nor U3612 (N_3612,N_1130,N_1527);
and U3613 (N_3613,N_1395,N_1455);
and U3614 (N_3614,N_1045,N_110);
nand U3615 (N_3615,N_1078,N_1800);
nor U3616 (N_3616,N_1274,N_759);
or U3617 (N_3617,N_1789,N_604);
and U3618 (N_3618,N_65,N_1319);
or U3619 (N_3619,N_1588,N_1974);
and U3620 (N_3620,N_1333,N_1649);
or U3621 (N_3621,N_1291,N_908);
nand U3622 (N_3622,N_790,N_1141);
nand U3623 (N_3623,N_1434,N_152);
nor U3624 (N_3624,N_67,N_317);
and U3625 (N_3625,N_168,N_987);
xor U3626 (N_3626,N_929,N_1738);
nand U3627 (N_3627,N_1484,N_613);
or U3628 (N_3628,N_649,N_933);
nor U3629 (N_3629,N_879,N_812);
and U3630 (N_3630,N_1563,N_655);
nor U3631 (N_3631,N_802,N_666);
or U3632 (N_3632,N_1103,N_109);
nand U3633 (N_3633,N_1305,N_1919);
nor U3634 (N_3634,N_957,N_525);
or U3635 (N_3635,N_895,N_1947);
nor U3636 (N_3636,N_590,N_119);
nor U3637 (N_3637,N_465,N_634);
or U3638 (N_3638,N_411,N_923);
nand U3639 (N_3639,N_1657,N_1632);
or U3640 (N_3640,N_269,N_79);
nor U3641 (N_3641,N_1598,N_1066);
xor U3642 (N_3642,N_656,N_750);
nand U3643 (N_3643,N_1615,N_1176);
or U3644 (N_3644,N_1514,N_1692);
or U3645 (N_3645,N_14,N_241);
nand U3646 (N_3646,N_454,N_1873);
or U3647 (N_3647,N_1264,N_517);
or U3648 (N_3648,N_258,N_1259);
nor U3649 (N_3649,N_899,N_1740);
and U3650 (N_3650,N_194,N_1657);
nand U3651 (N_3651,N_247,N_869);
nand U3652 (N_3652,N_1794,N_648);
nor U3653 (N_3653,N_8,N_1066);
nand U3654 (N_3654,N_1143,N_1544);
and U3655 (N_3655,N_1305,N_712);
or U3656 (N_3656,N_1801,N_261);
and U3657 (N_3657,N_779,N_710);
and U3658 (N_3658,N_1777,N_1552);
nor U3659 (N_3659,N_1143,N_533);
and U3660 (N_3660,N_387,N_843);
and U3661 (N_3661,N_1614,N_1972);
nand U3662 (N_3662,N_1434,N_255);
and U3663 (N_3663,N_1983,N_1470);
and U3664 (N_3664,N_1362,N_1731);
or U3665 (N_3665,N_269,N_816);
nor U3666 (N_3666,N_412,N_187);
and U3667 (N_3667,N_296,N_1094);
or U3668 (N_3668,N_1890,N_1373);
xnor U3669 (N_3669,N_1639,N_425);
nand U3670 (N_3670,N_149,N_1910);
or U3671 (N_3671,N_1568,N_1268);
or U3672 (N_3672,N_779,N_1364);
nor U3673 (N_3673,N_319,N_1399);
nor U3674 (N_3674,N_318,N_718);
or U3675 (N_3675,N_205,N_776);
nand U3676 (N_3676,N_541,N_242);
and U3677 (N_3677,N_200,N_756);
or U3678 (N_3678,N_841,N_1441);
nand U3679 (N_3679,N_481,N_657);
nand U3680 (N_3680,N_1721,N_1582);
nor U3681 (N_3681,N_0,N_481);
or U3682 (N_3682,N_1475,N_341);
and U3683 (N_3683,N_1709,N_1291);
or U3684 (N_3684,N_1697,N_73);
or U3685 (N_3685,N_1577,N_579);
nor U3686 (N_3686,N_1326,N_329);
nor U3687 (N_3687,N_446,N_1742);
or U3688 (N_3688,N_1563,N_239);
xnor U3689 (N_3689,N_1034,N_33);
or U3690 (N_3690,N_1517,N_1513);
nand U3691 (N_3691,N_955,N_1935);
or U3692 (N_3692,N_714,N_1876);
or U3693 (N_3693,N_1314,N_781);
nor U3694 (N_3694,N_1690,N_1655);
nand U3695 (N_3695,N_939,N_208);
nor U3696 (N_3696,N_1078,N_145);
and U3697 (N_3697,N_1471,N_1648);
nor U3698 (N_3698,N_704,N_83);
and U3699 (N_3699,N_1704,N_1821);
or U3700 (N_3700,N_1522,N_1546);
xor U3701 (N_3701,N_286,N_1576);
xnor U3702 (N_3702,N_1998,N_131);
nand U3703 (N_3703,N_1425,N_784);
nand U3704 (N_3704,N_560,N_1027);
nand U3705 (N_3705,N_1481,N_387);
or U3706 (N_3706,N_1101,N_1173);
nor U3707 (N_3707,N_1004,N_629);
nor U3708 (N_3708,N_1282,N_1762);
nor U3709 (N_3709,N_329,N_1956);
nor U3710 (N_3710,N_1468,N_1054);
nand U3711 (N_3711,N_1188,N_1764);
or U3712 (N_3712,N_1188,N_1419);
nor U3713 (N_3713,N_1914,N_53);
or U3714 (N_3714,N_332,N_1902);
nand U3715 (N_3715,N_523,N_406);
or U3716 (N_3716,N_38,N_1813);
nand U3717 (N_3717,N_118,N_1179);
nor U3718 (N_3718,N_1289,N_1121);
nor U3719 (N_3719,N_1197,N_584);
and U3720 (N_3720,N_1023,N_1471);
nor U3721 (N_3721,N_1147,N_1577);
and U3722 (N_3722,N_819,N_132);
and U3723 (N_3723,N_368,N_338);
nand U3724 (N_3724,N_687,N_916);
nor U3725 (N_3725,N_699,N_603);
or U3726 (N_3726,N_549,N_7);
and U3727 (N_3727,N_790,N_1591);
and U3728 (N_3728,N_1257,N_120);
or U3729 (N_3729,N_136,N_1501);
nand U3730 (N_3730,N_445,N_1078);
nand U3731 (N_3731,N_1519,N_387);
and U3732 (N_3732,N_731,N_1231);
and U3733 (N_3733,N_991,N_1741);
xnor U3734 (N_3734,N_1375,N_1112);
or U3735 (N_3735,N_631,N_1942);
nor U3736 (N_3736,N_348,N_723);
and U3737 (N_3737,N_1773,N_101);
xor U3738 (N_3738,N_850,N_1307);
and U3739 (N_3739,N_470,N_897);
and U3740 (N_3740,N_251,N_230);
nor U3741 (N_3741,N_423,N_1916);
nand U3742 (N_3742,N_1449,N_97);
nor U3743 (N_3743,N_79,N_382);
nor U3744 (N_3744,N_167,N_1255);
or U3745 (N_3745,N_1779,N_586);
or U3746 (N_3746,N_1029,N_850);
or U3747 (N_3747,N_308,N_845);
and U3748 (N_3748,N_281,N_223);
or U3749 (N_3749,N_1567,N_1290);
or U3750 (N_3750,N_994,N_457);
nand U3751 (N_3751,N_1794,N_1187);
nand U3752 (N_3752,N_1956,N_282);
and U3753 (N_3753,N_479,N_1806);
and U3754 (N_3754,N_411,N_395);
and U3755 (N_3755,N_1565,N_1963);
or U3756 (N_3756,N_1331,N_1629);
or U3757 (N_3757,N_50,N_1970);
or U3758 (N_3758,N_755,N_513);
nor U3759 (N_3759,N_1400,N_1486);
nand U3760 (N_3760,N_1992,N_847);
nand U3761 (N_3761,N_942,N_1452);
nand U3762 (N_3762,N_1646,N_513);
or U3763 (N_3763,N_1197,N_1055);
and U3764 (N_3764,N_1212,N_1487);
nand U3765 (N_3765,N_668,N_290);
or U3766 (N_3766,N_889,N_318);
nor U3767 (N_3767,N_722,N_958);
or U3768 (N_3768,N_1871,N_812);
or U3769 (N_3769,N_852,N_1052);
nand U3770 (N_3770,N_1232,N_768);
nand U3771 (N_3771,N_567,N_1514);
nor U3772 (N_3772,N_264,N_1300);
and U3773 (N_3773,N_1349,N_1306);
or U3774 (N_3774,N_1801,N_450);
nand U3775 (N_3775,N_667,N_1598);
or U3776 (N_3776,N_1056,N_1523);
or U3777 (N_3777,N_1693,N_638);
and U3778 (N_3778,N_443,N_123);
nand U3779 (N_3779,N_383,N_417);
or U3780 (N_3780,N_200,N_693);
nor U3781 (N_3781,N_1845,N_1823);
or U3782 (N_3782,N_730,N_1523);
nor U3783 (N_3783,N_975,N_474);
nor U3784 (N_3784,N_145,N_1416);
or U3785 (N_3785,N_673,N_378);
nor U3786 (N_3786,N_1007,N_1342);
and U3787 (N_3787,N_1713,N_718);
nor U3788 (N_3788,N_1444,N_1359);
nand U3789 (N_3789,N_1934,N_762);
nor U3790 (N_3790,N_1056,N_763);
or U3791 (N_3791,N_1063,N_507);
or U3792 (N_3792,N_785,N_970);
or U3793 (N_3793,N_197,N_1179);
or U3794 (N_3794,N_844,N_1649);
or U3795 (N_3795,N_814,N_1801);
nand U3796 (N_3796,N_1004,N_740);
or U3797 (N_3797,N_1732,N_598);
nand U3798 (N_3798,N_561,N_740);
or U3799 (N_3799,N_560,N_1458);
and U3800 (N_3800,N_1396,N_839);
nand U3801 (N_3801,N_10,N_660);
xor U3802 (N_3802,N_859,N_687);
nor U3803 (N_3803,N_1992,N_1179);
nand U3804 (N_3804,N_467,N_730);
nand U3805 (N_3805,N_101,N_1960);
nand U3806 (N_3806,N_1203,N_1090);
or U3807 (N_3807,N_513,N_350);
and U3808 (N_3808,N_1672,N_1924);
and U3809 (N_3809,N_1211,N_1384);
nor U3810 (N_3810,N_1608,N_1836);
nand U3811 (N_3811,N_1310,N_1812);
and U3812 (N_3812,N_883,N_1785);
and U3813 (N_3813,N_1366,N_1521);
nand U3814 (N_3814,N_933,N_491);
nor U3815 (N_3815,N_494,N_850);
nand U3816 (N_3816,N_1531,N_417);
nand U3817 (N_3817,N_1942,N_1145);
xnor U3818 (N_3818,N_765,N_1014);
or U3819 (N_3819,N_1809,N_762);
and U3820 (N_3820,N_1882,N_983);
or U3821 (N_3821,N_353,N_843);
or U3822 (N_3822,N_656,N_1148);
and U3823 (N_3823,N_1987,N_332);
and U3824 (N_3824,N_1244,N_1524);
or U3825 (N_3825,N_164,N_1795);
and U3826 (N_3826,N_1674,N_864);
nor U3827 (N_3827,N_773,N_812);
and U3828 (N_3828,N_1220,N_958);
or U3829 (N_3829,N_1214,N_277);
and U3830 (N_3830,N_459,N_387);
xor U3831 (N_3831,N_1459,N_241);
or U3832 (N_3832,N_1136,N_1254);
nand U3833 (N_3833,N_1816,N_567);
nand U3834 (N_3834,N_267,N_1496);
and U3835 (N_3835,N_1598,N_66);
nand U3836 (N_3836,N_1066,N_611);
and U3837 (N_3837,N_1937,N_1521);
or U3838 (N_3838,N_625,N_928);
or U3839 (N_3839,N_643,N_654);
nor U3840 (N_3840,N_522,N_1374);
and U3841 (N_3841,N_1364,N_1817);
nor U3842 (N_3842,N_1826,N_82);
and U3843 (N_3843,N_1250,N_1450);
nor U3844 (N_3844,N_1459,N_211);
or U3845 (N_3845,N_426,N_1536);
nand U3846 (N_3846,N_652,N_250);
nor U3847 (N_3847,N_1565,N_1705);
nor U3848 (N_3848,N_16,N_807);
and U3849 (N_3849,N_1508,N_995);
and U3850 (N_3850,N_1680,N_41);
or U3851 (N_3851,N_400,N_352);
nand U3852 (N_3852,N_344,N_1958);
or U3853 (N_3853,N_1750,N_988);
or U3854 (N_3854,N_313,N_470);
nor U3855 (N_3855,N_1896,N_884);
nand U3856 (N_3856,N_1341,N_1212);
nor U3857 (N_3857,N_1479,N_399);
and U3858 (N_3858,N_534,N_1124);
nand U3859 (N_3859,N_631,N_1766);
nor U3860 (N_3860,N_180,N_217);
or U3861 (N_3861,N_1768,N_272);
xnor U3862 (N_3862,N_834,N_926);
nand U3863 (N_3863,N_1141,N_1655);
or U3864 (N_3864,N_1779,N_98);
nand U3865 (N_3865,N_1432,N_809);
or U3866 (N_3866,N_1985,N_569);
or U3867 (N_3867,N_1991,N_758);
nand U3868 (N_3868,N_511,N_1845);
and U3869 (N_3869,N_23,N_38);
nand U3870 (N_3870,N_620,N_301);
and U3871 (N_3871,N_1312,N_808);
and U3872 (N_3872,N_542,N_1873);
or U3873 (N_3873,N_896,N_1817);
and U3874 (N_3874,N_141,N_142);
and U3875 (N_3875,N_736,N_887);
or U3876 (N_3876,N_1915,N_317);
or U3877 (N_3877,N_1552,N_1765);
nand U3878 (N_3878,N_1835,N_1849);
nand U3879 (N_3879,N_1678,N_546);
nand U3880 (N_3880,N_1411,N_496);
nor U3881 (N_3881,N_1932,N_671);
and U3882 (N_3882,N_220,N_1652);
or U3883 (N_3883,N_1122,N_209);
nand U3884 (N_3884,N_88,N_1576);
and U3885 (N_3885,N_239,N_1365);
and U3886 (N_3886,N_151,N_1866);
or U3887 (N_3887,N_994,N_291);
and U3888 (N_3888,N_686,N_979);
nor U3889 (N_3889,N_314,N_1057);
or U3890 (N_3890,N_1264,N_467);
or U3891 (N_3891,N_473,N_744);
and U3892 (N_3892,N_1371,N_14);
and U3893 (N_3893,N_1255,N_390);
nor U3894 (N_3894,N_1435,N_352);
nand U3895 (N_3895,N_1823,N_587);
and U3896 (N_3896,N_1906,N_209);
nand U3897 (N_3897,N_8,N_1654);
xnor U3898 (N_3898,N_707,N_1561);
nand U3899 (N_3899,N_1504,N_441);
and U3900 (N_3900,N_1444,N_1126);
nand U3901 (N_3901,N_421,N_1554);
nor U3902 (N_3902,N_259,N_1451);
nand U3903 (N_3903,N_417,N_1899);
nor U3904 (N_3904,N_523,N_808);
or U3905 (N_3905,N_1441,N_737);
or U3906 (N_3906,N_191,N_307);
and U3907 (N_3907,N_723,N_1367);
nor U3908 (N_3908,N_1288,N_1949);
and U3909 (N_3909,N_84,N_1655);
or U3910 (N_3910,N_47,N_120);
nand U3911 (N_3911,N_926,N_1216);
nand U3912 (N_3912,N_577,N_105);
and U3913 (N_3913,N_327,N_1707);
or U3914 (N_3914,N_412,N_1196);
or U3915 (N_3915,N_1214,N_247);
nand U3916 (N_3916,N_1424,N_1023);
or U3917 (N_3917,N_7,N_339);
or U3918 (N_3918,N_698,N_89);
and U3919 (N_3919,N_1066,N_1067);
xor U3920 (N_3920,N_477,N_151);
and U3921 (N_3921,N_1370,N_1130);
and U3922 (N_3922,N_1396,N_1825);
or U3923 (N_3923,N_49,N_1526);
and U3924 (N_3924,N_1028,N_241);
nand U3925 (N_3925,N_453,N_1340);
and U3926 (N_3926,N_1382,N_1836);
nor U3927 (N_3927,N_1100,N_360);
nand U3928 (N_3928,N_956,N_52);
nor U3929 (N_3929,N_1529,N_459);
and U3930 (N_3930,N_125,N_159);
or U3931 (N_3931,N_423,N_673);
nor U3932 (N_3932,N_1740,N_693);
and U3933 (N_3933,N_1358,N_1727);
and U3934 (N_3934,N_1322,N_203);
or U3935 (N_3935,N_1143,N_1713);
nor U3936 (N_3936,N_500,N_835);
nor U3937 (N_3937,N_793,N_794);
or U3938 (N_3938,N_549,N_1362);
nand U3939 (N_3939,N_148,N_76);
and U3940 (N_3940,N_464,N_10);
or U3941 (N_3941,N_1218,N_220);
and U3942 (N_3942,N_1950,N_852);
or U3943 (N_3943,N_322,N_1053);
nand U3944 (N_3944,N_1860,N_1880);
nand U3945 (N_3945,N_696,N_1509);
or U3946 (N_3946,N_1502,N_419);
nand U3947 (N_3947,N_505,N_1134);
xnor U3948 (N_3948,N_1552,N_354);
nor U3949 (N_3949,N_1769,N_671);
nand U3950 (N_3950,N_1709,N_58);
nor U3951 (N_3951,N_1799,N_337);
nor U3952 (N_3952,N_667,N_968);
xnor U3953 (N_3953,N_1090,N_1892);
nor U3954 (N_3954,N_278,N_291);
and U3955 (N_3955,N_955,N_919);
or U3956 (N_3956,N_699,N_936);
and U3957 (N_3957,N_995,N_669);
or U3958 (N_3958,N_1945,N_117);
nand U3959 (N_3959,N_636,N_1688);
or U3960 (N_3960,N_818,N_173);
or U3961 (N_3961,N_740,N_370);
nand U3962 (N_3962,N_781,N_1133);
or U3963 (N_3963,N_1525,N_684);
and U3964 (N_3964,N_938,N_1434);
and U3965 (N_3965,N_1547,N_653);
or U3966 (N_3966,N_343,N_50);
nor U3967 (N_3967,N_1892,N_303);
nand U3968 (N_3968,N_66,N_1490);
nand U3969 (N_3969,N_1697,N_1909);
nor U3970 (N_3970,N_261,N_1398);
xnor U3971 (N_3971,N_783,N_1071);
nor U3972 (N_3972,N_1437,N_389);
xor U3973 (N_3973,N_74,N_1879);
or U3974 (N_3974,N_1652,N_190);
nor U3975 (N_3975,N_1893,N_522);
nand U3976 (N_3976,N_1841,N_680);
nand U3977 (N_3977,N_421,N_1844);
or U3978 (N_3978,N_812,N_730);
or U3979 (N_3979,N_454,N_736);
nor U3980 (N_3980,N_1518,N_1607);
and U3981 (N_3981,N_1570,N_1965);
nand U3982 (N_3982,N_774,N_1760);
or U3983 (N_3983,N_1523,N_391);
or U3984 (N_3984,N_951,N_1115);
nand U3985 (N_3985,N_978,N_1999);
and U3986 (N_3986,N_725,N_1601);
xnor U3987 (N_3987,N_296,N_1020);
nand U3988 (N_3988,N_754,N_197);
nor U3989 (N_3989,N_1117,N_272);
nor U3990 (N_3990,N_680,N_98);
nand U3991 (N_3991,N_1031,N_1229);
or U3992 (N_3992,N_110,N_1375);
or U3993 (N_3993,N_343,N_1616);
or U3994 (N_3994,N_1363,N_1728);
nand U3995 (N_3995,N_314,N_948);
and U3996 (N_3996,N_1731,N_1706);
or U3997 (N_3997,N_1633,N_286);
and U3998 (N_3998,N_228,N_1857);
nor U3999 (N_3999,N_1520,N_372);
or U4000 (N_4000,N_3501,N_2317);
nand U4001 (N_4001,N_3367,N_2798);
nand U4002 (N_4002,N_2514,N_2587);
nand U4003 (N_4003,N_2996,N_3092);
nand U4004 (N_4004,N_3914,N_2816);
nand U4005 (N_4005,N_2336,N_2190);
nand U4006 (N_4006,N_2539,N_2402);
or U4007 (N_4007,N_3513,N_2745);
xnor U4008 (N_4008,N_3894,N_3647);
nor U4009 (N_4009,N_2167,N_2557);
nand U4010 (N_4010,N_3899,N_2691);
nand U4011 (N_4011,N_3742,N_3630);
and U4012 (N_4012,N_3849,N_3814);
nand U4013 (N_4013,N_2796,N_3182);
and U4014 (N_4014,N_3911,N_3981);
nand U4015 (N_4015,N_3836,N_2156);
nand U4016 (N_4016,N_2791,N_2563);
or U4017 (N_4017,N_3681,N_3714);
nor U4018 (N_4018,N_3290,N_2312);
nor U4019 (N_4019,N_2401,N_2723);
and U4020 (N_4020,N_3403,N_3080);
and U4021 (N_4021,N_3005,N_2582);
nand U4022 (N_4022,N_2934,N_2201);
nor U4023 (N_4023,N_3793,N_3198);
and U4024 (N_4024,N_2044,N_2846);
and U4025 (N_4025,N_2345,N_2565);
nor U4026 (N_4026,N_3078,N_2133);
and U4027 (N_4027,N_3248,N_2763);
and U4028 (N_4028,N_3517,N_3750);
or U4029 (N_4029,N_2154,N_3328);
nor U4030 (N_4030,N_3510,N_2307);
or U4031 (N_4031,N_3229,N_3283);
nor U4032 (N_4032,N_2130,N_3075);
or U4033 (N_4033,N_2486,N_2525);
or U4034 (N_4034,N_2021,N_2974);
and U4035 (N_4035,N_3208,N_2131);
nor U4036 (N_4036,N_2781,N_3994);
nor U4037 (N_4037,N_2544,N_3298);
nor U4038 (N_4038,N_2939,N_2794);
nand U4039 (N_4039,N_2792,N_2387);
nor U4040 (N_4040,N_3842,N_3418);
or U4041 (N_4041,N_2249,N_3292);
or U4042 (N_4042,N_3712,N_3378);
nand U4043 (N_4043,N_2170,N_3325);
and U4044 (N_4044,N_3048,N_2032);
nand U4045 (N_4045,N_3760,N_2024);
nand U4046 (N_4046,N_2164,N_3875);
nor U4047 (N_4047,N_3779,N_2162);
or U4048 (N_4048,N_2653,N_2177);
xnor U4049 (N_4049,N_2208,N_2376);
and U4050 (N_4050,N_3905,N_2166);
nor U4051 (N_4051,N_3958,N_2385);
nor U4052 (N_4052,N_2528,N_2997);
and U4053 (N_4053,N_2219,N_3550);
and U4054 (N_4054,N_2921,N_2398);
or U4055 (N_4055,N_3168,N_3929);
nand U4056 (N_4056,N_2982,N_2589);
or U4057 (N_4057,N_3172,N_3096);
nor U4058 (N_4058,N_2260,N_3205);
and U4059 (N_4059,N_3044,N_3424);
or U4060 (N_4060,N_2835,N_2574);
nand U4061 (N_4061,N_2606,N_2408);
or U4062 (N_4062,N_2603,N_3727);
and U4063 (N_4063,N_2004,N_2183);
nor U4064 (N_4064,N_2901,N_3968);
and U4065 (N_4065,N_3640,N_2947);
or U4066 (N_4066,N_2225,N_2141);
or U4067 (N_4067,N_2071,N_3040);
nand U4068 (N_4068,N_2025,N_2082);
or U4069 (N_4069,N_2296,N_3269);
nor U4070 (N_4070,N_2909,N_3938);
nor U4071 (N_4071,N_3568,N_3989);
or U4072 (N_4072,N_2590,N_3065);
nand U4073 (N_4073,N_3865,N_2553);
or U4074 (N_4074,N_3210,N_2185);
nand U4075 (N_4075,N_3536,N_3434);
and U4076 (N_4076,N_3617,N_2833);
nor U4077 (N_4077,N_2628,N_3333);
and U4078 (N_4078,N_3547,N_3670);
and U4079 (N_4079,N_2019,N_3058);
nand U4080 (N_4080,N_2168,N_2262);
and U4081 (N_4081,N_2878,N_2330);
nand U4082 (N_4082,N_2320,N_3483);
nor U4083 (N_4083,N_2832,N_3680);
nor U4084 (N_4084,N_2028,N_3456);
and U4085 (N_4085,N_3847,N_3488);
and U4086 (N_4086,N_3982,N_2046);
or U4087 (N_4087,N_2567,N_2991);
and U4088 (N_4088,N_3996,N_2418);
or U4089 (N_4089,N_2963,N_3857);
xor U4090 (N_4090,N_2403,N_2124);
and U4091 (N_4091,N_2661,N_3344);
nand U4092 (N_4092,N_3533,N_2783);
and U4093 (N_4093,N_3618,N_2689);
and U4094 (N_4094,N_3913,N_2441);
nand U4095 (N_4095,N_2456,N_2643);
and U4096 (N_4096,N_3338,N_2365);
nand U4097 (N_4097,N_3294,N_2920);
nand U4098 (N_4098,N_2862,N_3309);
and U4099 (N_4099,N_3498,N_2522);
or U4100 (N_4100,N_2186,N_2984);
nor U4101 (N_4101,N_2093,N_2849);
nor U4102 (N_4102,N_3464,N_2622);
and U4103 (N_4103,N_2710,N_2586);
and U4104 (N_4104,N_3976,N_2102);
and U4105 (N_4105,N_2207,N_2298);
and U4106 (N_4106,N_2142,N_3851);
nand U4107 (N_4107,N_2944,N_3861);
nand U4108 (N_4108,N_2638,N_3348);
nor U4109 (N_4109,N_3364,N_2613);
nor U4110 (N_4110,N_3113,N_3770);
and U4111 (N_4111,N_2072,N_2989);
nand U4112 (N_4112,N_2516,N_3329);
or U4113 (N_4113,N_2550,N_2425);
nand U4114 (N_4114,N_2226,N_2075);
nor U4115 (N_4115,N_3305,N_3937);
and U4116 (N_4116,N_2200,N_2034);
nor U4117 (N_4117,N_3500,N_3060);
nor U4118 (N_4118,N_3398,N_2632);
or U4119 (N_4119,N_3232,N_2147);
and U4120 (N_4120,N_3869,N_2578);
or U4121 (N_4121,N_3628,N_3451);
xor U4122 (N_4122,N_2035,N_2520);
or U4123 (N_4123,N_2535,N_2502);
or U4124 (N_4124,N_2378,N_2434);
xnor U4125 (N_4125,N_2374,N_3320);
and U4126 (N_4126,N_2874,N_3763);
or U4127 (N_4127,N_3186,N_3528);
nor U4128 (N_4128,N_2679,N_2955);
nand U4129 (N_4129,N_2845,N_2828);
or U4130 (N_4130,N_2411,N_3773);
or U4131 (N_4131,N_3392,N_3735);
nand U4132 (N_4132,N_2671,N_3357);
or U4133 (N_4133,N_3459,N_3184);
nor U4134 (N_4134,N_3031,N_3682);
or U4135 (N_4135,N_2990,N_2198);
nor U4136 (N_4136,N_2615,N_2364);
nor U4137 (N_4137,N_3771,N_2000);
nand U4138 (N_4138,N_3543,N_2526);
nor U4139 (N_4139,N_3702,N_2215);
nor U4140 (N_4140,N_3455,N_3067);
or U4141 (N_4141,N_3446,N_3175);
nor U4142 (N_4142,N_2419,N_3070);
and U4143 (N_4143,N_3594,N_3073);
nand U4144 (N_4144,N_3002,N_2209);
nor U4145 (N_4145,N_3605,N_2962);
nor U4146 (N_4146,N_3970,N_2258);
nand U4147 (N_4147,N_2158,N_2477);
nor U4148 (N_4148,N_2736,N_3672);
and U4149 (N_4149,N_2057,N_3752);
or U4150 (N_4150,N_3537,N_2961);
or U4151 (N_4151,N_3188,N_3711);
nand U4152 (N_4152,N_3127,N_2692);
or U4153 (N_4153,N_2308,N_2125);
nor U4154 (N_4154,N_2808,N_2029);
and U4155 (N_4155,N_2211,N_3634);
nor U4156 (N_4156,N_2337,N_3153);
and U4157 (N_4157,N_3164,N_2016);
or U4158 (N_4158,N_3614,N_2700);
or U4159 (N_4159,N_3107,N_2457);
or U4160 (N_4160,N_2150,N_3878);
or U4161 (N_4161,N_2667,N_3017);
nor U4162 (N_4162,N_2817,N_2455);
nand U4163 (N_4163,N_3792,N_3947);
nor U4164 (N_4164,N_3926,N_3102);
and U4165 (N_4165,N_3803,N_3924);
nor U4166 (N_4166,N_2357,N_3915);
and U4167 (N_4167,N_3038,N_2511);
nand U4168 (N_4168,N_3918,N_2316);
and U4169 (N_4169,N_3016,N_2508);
or U4170 (N_4170,N_2439,N_3962);
nor U4171 (N_4171,N_2136,N_2888);
and U4172 (N_4172,N_3995,N_2304);
nand U4173 (N_4173,N_3748,N_3492);
nor U4174 (N_4174,N_3419,N_3293);
nor U4175 (N_4175,N_3006,N_2840);
or U4176 (N_4176,N_2759,N_3693);
nand U4177 (N_4177,N_2863,N_2010);
and U4178 (N_4178,N_2640,N_3971);
nand U4179 (N_4179,N_3809,N_2468);
and U4180 (N_4180,N_2246,N_3595);
nand U4181 (N_4181,N_2799,N_3093);
or U4182 (N_4182,N_2730,N_2814);
xnor U4183 (N_4183,N_3588,N_2804);
and U4184 (N_4184,N_2726,N_3241);
nor U4185 (N_4185,N_3395,N_3355);
and U4186 (N_4186,N_2676,N_2519);
or U4187 (N_4187,N_2875,N_2255);
or U4188 (N_4188,N_3219,N_2732);
nor U4189 (N_4189,N_2197,N_2143);
and U4190 (N_4190,N_3405,N_3237);
and U4191 (N_4191,N_3432,N_2279);
nor U4192 (N_4192,N_2916,N_2424);
nor U4193 (N_4193,N_3389,N_2543);
nor U4194 (N_4194,N_2980,N_3105);
nand U4195 (N_4195,N_2534,N_2678);
and U4196 (N_4196,N_2247,N_3146);
and U4197 (N_4197,N_2076,N_3068);
nand U4198 (N_4198,N_3375,N_3558);
and U4199 (N_4199,N_2275,N_3648);
or U4200 (N_4200,N_2104,N_2503);
nand U4201 (N_4201,N_3445,N_3694);
and U4202 (N_4202,N_2105,N_2447);
and U4203 (N_4203,N_2889,N_2416);
nor U4204 (N_4204,N_3804,N_3521);
and U4205 (N_4205,N_2490,N_3365);
and U4206 (N_4206,N_3291,N_3766);
nor U4207 (N_4207,N_2524,N_2070);
nand U4208 (N_4208,N_2639,N_3725);
xor U4209 (N_4209,N_3719,N_2002);
nand U4210 (N_4210,N_2542,N_3585);
nor U4211 (N_4211,N_3930,N_3281);
or U4212 (N_4212,N_2406,N_3271);
nand U4213 (N_4213,N_2039,N_3011);
and U4214 (N_4214,N_2435,N_3362);
nor U4215 (N_4215,N_2810,N_2687);
or U4216 (N_4216,N_2785,N_2851);
nor U4217 (N_4217,N_2668,N_3360);
and U4218 (N_4218,N_2096,N_2634);
or U4219 (N_4219,N_2397,N_3575);
nand U4220 (N_4220,N_2952,N_2940);
or U4221 (N_4221,N_3907,N_3977);
nand U4222 (N_4222,N_2560,N_2054);
nor U4223 (N_4223,N_3654,N_3676);
nor U4224 (N_4224,N_2256,N_3114);
nand U4225 (N_4225,N_3235,N_2517);
or U4226 (N_4226,N_3313,N_3255);
nor U4227 (N_4227,N_2829,N_2263);
and U4228 (N_4228,N_2472,N_3862);
and U4229 (N_4229,N_2857,N_3593);
nor U4230 (N_4230,N_3579,N_2273);
nand U4231 (N_4231,N_3003,N_2344);
nor U4232 (N_4232,N_2965,N_3508);
or U4233 (N_4233,N_3191,N_3484);
or U4234 (N_4234,N_2098,N_3826);
nor U4235 (N_4235,N_2975,N_2598);
and U4236 (N_4236,N_3376,N_2015);
nand U4237 (N_4237,N_2051,N_2248);
and U4238 (N_4238,N_2487,N_3876);
or U4239 (N_4239,N_2338,N_3904);
or U4240 (N_4240,N_2068,N_3877);
or U4241 (N_4241,N_2847,N_2079);
and U4242 (N_4242,N_3286,N_2876);
or U4243 (N_4243,N_2631,N_2972);
or U4244 (N_4244,N_3317,N_2719);
or U4245 (N_4245,N_3984,N_3729);
and U4246 (N_4246,N_2351,N_3731);
nand U4247 (N_4247,N_2770,N_3589);
nand U4248 (N_4248,N_2746,N_2358);
or U4249 (N_4249,N_2196,N_3131);
or U4250 (N_4250,N_3134,N_2549);
or U4251 (N_4251,N_2592,N_2795);
nor U4252 (N_4252,N_3300,N_2103);
or U4253 (N_4253,N_3124,N_3870);
nor U4254 (N_4254,N_2427,N_3987);
nor U4255 (N_4255,N_3156,N_2652);
xor U4256 (N_4256,N_2891,N_3202);
nand U4257 (N_4257,N_2930,N_3110);
nor U4258 (N_4258,N_3025,N_2937);
or U4259 (N_4259,N_2957,N_2465);
and U4260 (N_4260,N_3468,N_3920);
or U4261 (N_4261,N_3089,N_2766);
and U4262 (N_4262,N_3385,N_3753);
nand U4263 (N_4263,N_3334,N_2698);
nor U4264 (N_4264,N_3452,N_2777);
or U4265 (N_4265,N_2844,N_2265);
or U4266 (N_4266,N_2742,N_2484);
nand U4267 (N_4267,N_2033,N_2393);
or U4268 (N_4268,N_3580,N_3326);
or U4269 (N_4269,N_2165,N_2601);
and U4270 (N_4270,N_3206,N_2738);
and U4271 (N_4271,N_3497,N_3145);
nand U4272 (N_4272,N_3509,N_2116);
xor U4273 (N_4273,N_2101,N_2675);
nand U4274 (N_4274,N_2390,N_3336);
and U4275 (N_4275,N_2917,N_3544);
and U4276 (N_4276,N_2548,N_2080);
and U4277 (N_4277,N_2161,N_2827);
nor U4278 (N_4278,N_3252,N_2762);
or U4279 (N_4279,N_2359,N_2681);
or U4280 (N_4280,N_2340,N_2043);
and U4281 (N_4281,N_2556,N_3043);
or U4282 (N_4282,N_3627,N_2064);
or U4283 (N_4283,N_2581,N_2893);
nor U4284 (N_4284,N_3413,N_3975);
nor U4285 (N_4285,N_3626,N_3493);
or U4286 (N_4286,N_3820,N_2491);
or U4287 (N_4287,N_3688,N_2597);
or U4288 (N_4288,N_2266,N_3928);
nor U4289 (N_4289,N_2583,N_2212);
nor U4290 (N_4290,N_3077,N_3399);
nand U4291 (N_4291,N_2721,N_3858);
xor U4292 (N_4292,N_3155,N_2600);
and U4293 (N_4293,N_3289,N_2464);
and U4294 (N_4294,N_3382,N_3474);
nand U4295 (N_4295,N_2053,N_3757);
or U4296 (N_4296,N_3818,N_2836);
nor U4297 (N_4297,N_3679,N_3176);
nor U4298 (N_4298,N_3658,N_2280);
and U4299 (N_4299,N_2869,N_2530);
or U4300 (N_4300,N_3505,N_3549);
or U4301 (N_4301,N_3236,N_2091);
nand U4302 (N_4302,N_2914,N_3400);
nor U4303 (N_4303,N_2967,N_2645);
xor U4304 (N_4304,N_3957,N_3366);
nor U4305 (N_4305,N_2752,N_2690);
nor U4306 (N_4306,N_2110,N_2321);
nor U4307 (N_4307,N_3925,N_2291);
nand U4308 (N_4308,N_3353,N_3657);
or U4309 (N_4309,N_3311,N_2483);
and U4310 (N_4310,N_3120,N_3577);
or U4311 (N_4311,N_3966,N_2189);
nor U4312 (N_4312,N_3039,N_2174);
xor U4313 (N_4313,N_2271,N_3087);
xnor U4314 (N_4314,N_2129,N_3986);
xor U4315 (N_4315,N_2325,N_2117);
nor U4316 (N_4316,N_3101,N_3169);
and U4317 (N_4317,N_3374,N_2218);
nand U4318 (N_4318,N_3377,N_3216);
nor U4319 (N_4319,N_3897,N_2228);
or U4320 (N_4320,N_2445,N_2669);
or U4321 (N_4321,N_3121,N_3831);
nand U4322 (N_4322,N_2148,N_2361);
and U4323 (N_4323,N_2782,N_2970);
and U4324 (N_4324,N_2459,N_3586);
nor U4325 (N_4325,N_2239,N_3460);
or U4326 (N_4326,N_2405,N_3838);
and U4327 (N_4327,N_3029,N_2078);
nand U4328 (N_4328,N_3481,N_3007);
nor U4329 (N_4329,N_3785,N_3499);
and U4330 (N_4330,N_2612,N_3447);
and U4331 (N_4331,N_2538,N_2444);
nor U4332 (N_4332,N_3931,N_2335);
and U4333 (N_4333,N_2910,N_3284);
and U4334 (N_4334,N_3906,N_2205);
nand U4335 (N_4335,N_3224,N_3581);
or U4336 (N_4336,N_3250,N_3315);
or U4337 (N_4337,N_2929,N_3462);
or U4338 (N_4338,N_3213,N_2496);
nand U4339 (N_4339,N_3154,N_3428);
nand U4340 (N_4340,N_2059,N_2060);
nand U4341 (N_4341,N_2062,N_3453);
and U4342 (N_4342,N_3222,N_2918);
nor U4343 (N_4343,N_2134,N_2146);
or U4344 (N_4344,N_2008,N_2480);
and U4345 (N_4345,N_3636,N_2813);
and U4346 (N_4346,N_3884,N_3754);
or U4347 (N_4347,N_2003,N_2693);
and U4348 (N_4348,N_3276,N_3787);
or U4349 (N_4349,N_3069,N_2949);
nand U4350 (N_4350,N_2153,N_3062);
nand U4351 (N_4351,N_2584,N_3346);
nor U4352 (N_4352,N_3525,N_2727);
nor U4353 (N_4353,N_3567,N_3018);
or U4354 (N_4354,N_3123,N_2386);
or U4355 (N_4355,N_3431,N_2452);
nor U4356 (N_4356,N_2287,N_3912);
nand U4357 (N_4357,N_2831,N_2518);
or U4358 (N_4358,N_2718,N_3845);
or U4359 (N_4359,N_3072,N_2780);
nor U4360 (N_4360,N_2540,N_3324);
or U4361 (N_4361,N_3259,N_2111);
and U4362 (N_4362,N_3756,N_3992);
or U4363 (N_4363,N_3337,N_2436);
or U4364 (N_4364,N_2728,N_3883);
and U4365 (N_4365,N_3279,N_3843);
or U4366 (N_4366,N_2194,N_2521);
and U4367 (N_4367,N_2801,N_3162);
or U4368 (N_4368,N_2213,N_3590);
and U4369 (N_4369,N_3523,N_3303);
nor U4370 (N_4370,N_2284,N_2375);
nor U4371 (N_4371,N_2904,N_2011);
nand U4372 (N_4372,N_3893,N_2686);
nand U4373 (N_4373,N_2013,N_3444);
nor U4374 (N_4374,N_3584,N_3821);
nand U4375 (N_4375,N_3437,N_2716);
nand U4376 (N_4376,N_3265,N_3192);
nor U4377 (N_4377,N_3314,N_2865);
or U4378 (N_4378,N_3258,N_3529);
and U4379 (N_4379,N_2356,N_3502);
nand U4380 (N_4380,N_2466,N_3319);
and U4381 (N_4381,N_3408,N_3530);
nor U4382 (N_4382,N_3383,N_3106);
nor U4383 (N_4383,N_3495,N_2115);
and U4384 (N_4384,N_2811,N_2908);
or U4385 (N_4385,N_2175,N_2095);
and U4386 (N_4386,N_3713,N_3220);
nor U4387 (N_4387,N_3637,N_2802);
or U4388 (N_4388,N_3012,N_2928);
nor U4389 (N_4389,N_2506,N_3323);
nand U4390 (N_4390,N_2259,N_3592);
nand U4391 (N_4391,N_2031,N_3243);
or U4392 (N_4392,N_2772,N_2709);
nor U4393 (N_4393,N_3420,N_2654);
nor U4394 (N_4394,N_2237,N_3936);
or U4395 (N_4395,N_3624,N_2712);
nand U4396 (N_4396,N_2852,N_3457);
or U4397 (N_4397,N_2463,N_2277);
nand U4398 (N_4398,N_3004,N_2343);
or U4399 (N_4399,N_3350,N_2683);
nand U4400 (N_4400,N_2417,N_2552);
or U4401 (N_4401,N_2887,N_2090);
and U4402 (N_4402,N_3489,N_2069);
or U4403 (N_4403,N_3433,N_3997);
nor U4404 (N_4404,N_3935,N_2896);
and U4405 (N_4405,N_3301,N_3496);
nand U4406 (N_4406,N_2642,N_2707);
nand U4407 (N_4407,N_3136,N_3504);
nor U4408 (N_4408,N_3978,N_2482);
and U4409 (N_4409,N_2339,N_3778);
nor U4410 (N_4410,N_2559,N_2276);
and U4411 (N_4411,N_2658,N_3387);
xor U4412 (N_4412,N_3562,N_3532);
nand U4413 (N_4413,N_3769,N_2058);
nand U4414 (N_4414,N_2446,N_3183);
and U4415 (N_4415,N_2244,N_2569);
and U4416 (N_4416,N_3764,N_3369);
nor U4417 (N_4417,N_3223,N_3703);
and U4418 (N_4418,N_3767,N_2608);
and U4419 (N_4419,N_2779,N_2925);
and U4420 (N_4420,N_2720,N_2301);
nand U4421 (N_4421,N_2555,N_2854);
nand U4422 (N_4422,N_3972,N_3638);
or U4423 (N_4423,N_3879,N_2510);
nand U4424 (N_4424,N_3867,N_3909);
nand U4425 (N_4425,N_2743,N_2903);
xor U4426 (N_4426,N_3860,N_3094);
nor U4427 (N_4427,N_2722,N_2531);
or U4428 (N_4428,N_2036,N_3086);
nand U4429 (N_4429,N_3921,N_2674);
nand U4430 (N_4430,N_3540,N_2853);
or U4431 (N_4431,N_3559,N_2206);
nand U4432 (N_4432,N_3221,N_3185);
or U4433 (N_4433,N_3274,N_3479);
nand U4434 (N_4434,N_2856,N_2089);
nor U4435 (N_4435,N_2270,N_3442);
or U4436 (N_4436,N_2030,N_3242);
and U4437 (N_4437,N_2257,N_3755);
nor U4438 (N_4438,N_2366,N_3143);
or U4439 (N_4439,N_3218,N_2094);
nor U4440 (N_4440,N_3422,N_2665);
or U4441 (N_4441,N_3841,N_3545);
and U4442 (N_4442,N_3611,N_3800);
or U4443 (N_4443,N_3449,N_3045);
nand U4444 (N_4444,N_3204,N_2380);
nor U4445 (N_4445,N_3844,N_2733);
nand U4446 (N_4446,N_3079,N_3049);
nor U4447 (N_4447,N_2987,N_3228);
nand U4448 (N_4448,N_2969,N_3850);
nand U4449 (N_4449,N_3423,N_3116);
nor U4450 (N_4450,N_2753,N_2670);
or U4451 (N_4451,N_3631,N_2907);
or U4452 (N_4452,N_3687,N_2655);
nor U4453 (N_4453,N_2498,N_2993);
nand U4454 (N_4454,N_3167,N_3660);
or U4455 (N_4455,N_2773,N_3349);
and U4456 (N_4456,N_3339,N_2610);
and U4457 (N_4457,N_3076,N_2122);
and U4458 (N_4458,N_2803,N_2221);
nand U4459 (N_4459,N_3587,N_3612);
or U4460 (N_4460,N_2572,N_3010);
nor U4461 (N_4461,N_2106,N_2493);
nand U4462 (N_4462,N_3356,N_3901);
nand U4463 (N_4463,N_2768,N_3028);
nor U4464 (N_4464,N_2859,N_2573);
nand U4465 (N_4465,N_2571,N_3190);
and U4466 (N_4466,N_3715,N_3788);
nand U4467 (N_4467,N_3129,N_2602);
nor U4468 (N_4468,N_2360,N_3209);
nand U4469 (N_4469,N_3370,N_3700);
nor U4470 (N_4470,N_3699,N_2625);
or U4471 (N_4471,N_3665,N_2651);
xor U4472 (N_4472,N_3784,N_2354);
nor U4473 (N_4473,N_3015,N_3014);
or U4474 (N_4474,N_2714,N_2604);
nand U4475 (N_4475,N_3885,N_3063);
and U4476 (N_4476,N_2245,N_3616);
nand U4477 (N_4477,N_2191,N_3759);
nand U4478 (N_4478,N_2353,N_3263);
or U4479 (N_4479,N_3761,N_2755);
and U4480 (N_4480,N_2898,N_2850);
nand U4481 (N_4481,N_2440,N_3494);
and U4482 (N_4482,N_2229,N_3601);
and U4483 (N_4483,N_2951,N_3762);
and U4484 (N_4484,N_2243,N_3623);
nor U4485 (N_4485,N_3606,N_3846);
nand U4486 (N_4486,N_2927,N_3109);
and U4487 (N_4487,N_3946,N_2877);
and U4488 (N_4488,N_2858,N_3082);
or U4489 (N_4489,N_3934,N_3280);
and U4490 (N_4490,N_3684,N_2985);
nor U4491 (N_4491,N_3022,N_2160);
nor U4492 (N_4492,N_3629,N_2793);
or U4493 (N_4493,N_3151,N_3193);
nor U4494 (N_4494,N_2178,N_2163);
or U4495 (N_4495,N_3066,N_3417);
nor U4496 (N_4496,N_2389,N_3917);
nor U4497 (N_4497,N_3194,N_3030);
nor U4498 (N_4498,N_2839,N_3371);
nor U4499 (N_4499,N_2217,N_3476);
nor U4500 (N_4500,N_3824,N_3683);
nand U4501 (N_4501,N_3572,N_3669);
or U4502 (N_4502,N_2254,N_2172);
nor U4503 (N_4503,N_2108,N_3932);
nand U4504 (N_4504,N_2626,N_2040);
nand U4505 (N_4505,N_3874,N_2494);
and U4506 (N_4506,N_2293,N_2334);
nand U4507 (N_4507,N_2038,N_3564);
and U4508 (N_4508,N_2328,N_3868);
nand U4509 (N_4509,N_2193,N_2861);
and U4510 (N_4510,N_2541,N_3083);
nand U4511 (N_4511,N_3013,N_2055);
nor U4512 (N_4512,N_3573,N_3643);
nand U4513 (N_4513,N_2577,N_2495);
and U4514 (N_4514,N_2757,N_2660);
or U4515 (N_4515,N_2294,N_2789);
and U4516 (N_4516,N_3384,N_2764);
or U4517 (N_4517,N_3535,N_3960);
xor U4518 (N_4518,N_3751,N_3179);
nand U4519 (N_4519,N_2536,N_2537);
nand U4520 (N_4520,N_2956,N_3864);
nor U4521 (N_4521,N_2066,N_3359);
or U4522 (N_4522,N_2157,N_2699);
nor U4523 (N_4523,N_3217,N_3983);
or U4524 (N_4524,N_2906,N_3873);
nand U4525 (N_4525,N_2462,N_3565);
xor U4526 (N_4526,N_3855,N_3827);
or U4527 (N_4527,N_3342,N_2314);
nor U4528 (N_4528,N_3717,N_2945);
or U4529 (N_4529,N_2926,N_2554);
or U4530 (N_4530,N_3282,N_3645);
or U4531 (N_4531,N_3507,N_2635);
or U4532 (N_4532,N_3686,N_3882);
and U4533 (N_4533,N_3429,N_2629);
nand U4534 (N_4534,N_2744,N_3563);
or U4535 (N_4535,N_2074,N_3569);
or U4536 (N_4536,N_2713,N_2421);
nor U4537 (N_4537,N_2007,N_2771);
or U4538 (N_4538,N_3436,N_2232);
or U4539 (N_4539,N_3830,N_2703);
or U4540 (N_4540,N_3227,N_3388);
or U4541 (N_4541,N_3659,N_3777);
nand U4542 (N_4542,N_3620,N_3173);
nor U4543 (N_4543,N_2825,N_3368);
nor U4544 (N_4544,N_2085,N_2501);
and U4545 (N_4545,N_3790,N_3231);
or U4546 (N_4546,N_2290,N_3091);
or U4547 (N_4547,N_2009,N_3187);
nand U4548 (N_4548,N_3740,N_3738);
or U4549 (N_4549,N_2740,N_3991);
nand U4550 (N_4550,N_3490,N_3570);
nand U4551 (N_4551,N_2885,N_3152);
and U4552 (N_4552,N_2529,N_2837);
or U4553 (N_4553,N_3226,N_3352);
and U4554 (N_4554,N_2621,N_3695);
nor U4555 (N_4555,N_3561,N_2152);
nor U4556 (N_4556,N_3622,N_2729);
nand U4557 (N_4557,N_2138,N_2048);
nor U4558 (N_4558,N_3652,N_2841);
nand U4559 (N_4559,N_3942,N_2299);
nor U4560 (N_4560,N_2313,N_3961);
and U4561 (N_4561,N_2609,N_2512);
nor U4562 (N_4562,N_2119,N_2018);
nor U4563 (N_4563,N_3287,N_3240);
and U4564 (N_4564,N_3122,N_3852);
or U4565 (N_4565,N_2735,N_2633);
nand U4566 (N_4566,N_3197,N_3599);
nor U4567 (N_4567,N_3948,N_3919);
nand U4568 (N_4568,N_2545,N_2943);
and U4569 (N_4569,N_2881,N_3653);
or U4570 (N_4570,N_2747,N_3985);
nand U4571 (N_4571,N_2333,N_2523);
nor U4572 (N_4572,N_2352,N_2139);
nand U4573 (N_4573,N_3212,N_3035);
nor U4574 (N_4574,N_3632,N_2426);
nand U4575 (N_4575,N_2868,N_3071);
or U4576 (N_4576,N_2919,N_3607);
or U4577 (N_4577,N_3794,N_2192);
nand U4578 (N_4578,N_2843,N_3288);
nand U4579 (N_4579,N_3677,N_3393);
nor U4580 (N_4580,N_3707,N_2968);
or U4581 (N_4581,N_2050,N_2127);
nor U4582 (N_4582,N_2149,N_3142);
nor U4583 (N_4583,N_2020,N_3160);
and U4584 (N_4584,N_2409,N_2588);
and U4585 (N_4585,N_2347,N_2924);
nor U4586 (N_4586,N_3421,N_3514);
nand U4587 (N_4587,N_2666,N_2725);
nor U4588 (N_4588,N_3988,N_2504);
xor U4589 (N_4589,N_3511,N_3741);
or U4590 (N_4590,N_2694,N_2045);
or U4591 (N_4591,N_2056,N_3140);
and U4592 (N_4592,N_2911,N_2145);
nor U4593 (N_4593,N_2902,N_3786);
nand U4594 (N_4594,N_2662,N_3180);
nand U4595 (N_4595,N_2761,N_2236);
or U4596 (N_4596,N_3697,N_2214);
and U4597 (N_4597,N_2499,N_3552);
nor U4598 (N_4598,N_2037,N_2900);
and U4599 (N_4599,N_3891,N_3394);
and U4600 (N_4600,N_3840,N_3927);
nor U4601 (N_4601,N_2123,N_3450);
nand U4602 (N_4602,N_2659,N_3472);
nor U4603 (N_4603,N_2179,N_3597);
nor U4604 (N_4604,N_2619,N_2734);
nor U4605 (N_4605,N_3522,N_3949);
or U4606 (N_4606,N_3404,N_2318);
nor U4607 (N_4607,N_2188,N_2306);
nor U4608 (N_4608,N_2216,N_3736);
and U4609 (N_4609,N_3430,N_3650);
nand U4610 (N_4610,N_2870,N_2289);
nor U4611 (N_4611,N_3829,N_3239);
and U4612 (N_4612,N_2332,N_2894);
nand U4613 (N_4613,N_3268,N_2935);
xnor U4614 (N_4614,N_2818,N_2591);
and U4615 (N_4615,N_2121,N_3443);
nor U4616 (N_4616,N_2605,N_3886);
nand U4617 (N_4617,N_3033,N_2994);
and U4618 (N_4618,N_2269,N_3796);
and U4619 (N_4619,N_3576,N_3486);
nor U4620 (N_4620,N_3853,N_2395);
or U4621 (N_4621,N_3866,N_3343);
and U4622 (N_4622,N_2758,N_3207);
or U4623 (N_4623,N_3137,N_2315);
nor U4624 (N_4624,N_3651,N_3396);
nor U4625 (N_4625,N_3835,N_2151);
and U4626 (N_4626,N_3415,N_3519);
nor U4627 (N_4627,N_2756,N_2527);
xnor U4628 (N_4628,N_3118,N_3888);
nand U4629 (N_4629,N_2371,N_3999);
nand U4630 (N_4630,N_3161,N_2492);
and U4631 (N_4631,N_2041,N_2251);
and U4632 (N_4632,N_3126,N_2824);
nand U4633 (N_4633,N_2933,N_3663);
and U4634 (N_4634,N_3008,N_3264);
nor U4635 (N_4635,N_2391,N_2327);
nor U4636 (N_4636,N_2181,N_3705);
nor U4637 (N_4637,N_3251,N_3482);
or U4638 (N_4638,N_3726,N_2497);
nand U4639 (N_4639,N_2724,N_2697);
nand U4640 (N_4640,N_2656,N_3908);
nand U4641 (N_4641,N_3956,N_2302);
and U4642 (N_4642,N_2561,N_2739);
nor U4643 (N_4643,N_2872,N_3747);
or U4644 (N_4644,N_3990,N_3034);
nand U4645 (N_4645,N_2180,N_2855);
or U4646 (N_4646,N_2617,N_2648);
nand U4647 (N_4647,N_2099,N_3438);
or U4648 (N_4648,N_3469,N_2005);
nand U4649 (N_4649,N_3801,N_3144);
or U4650 (N_4650,N_2883,N_3828);
nand U4651 (N_4651,N_3557,N_2017);
and U4652 (N_4652,N_2309,N_3487);
nand U4653 (N_4653,N_3454,N_2220);
nor U4654 (N_4654,N_2475,N_3733);
nor U4655 (N_4655,N_3461,N_3898);
nand U4656 (N_4656,N_2805,N_3621);
nor U4657 (N_4657,N_2372,N_2884);
or U4658 (N_4658,N_3655,N_2282);
nor U4659 (N_4659,N_2049,N_2941);
and U4660 (N_4660,N_3520,N_3189);
or U4661 (N_4661,N_3199,N_2964);
and U4662 (N_4662,N_2310,N_2381);
and U4663 (N_4663,N_2748,N_2500);
nand U4664 (N_4664,N_2442,N_3887);
nand U4665 (N_4665,N_3690,N_2731);
nor U4666 (N_4666,N_3644,N_3598);
nand U4667 (N_4667,N_3119,N_2912);
or U4668 (N_4668,N_2341,N_2437);
nor U4669 (N_4669,N_2261,N_3296);
nand U4670 (N_4670,N_2430,N_2614);
and U4671 (N_4671,N_2088,N_3608);
nand U4672 (N_4672,N_3174,N_3147);
and U4673 (N_4673,N_3625,N_3057);
nor U4674 (N_4674,N_3117,N_2750);
or U4675 (N_4675,N_3051,N_3299);
and U4676 (N_4676,N_2073,N_2864);
nand U4677 (N_4677,N_3635,N_3295);
nor U4678 (N_4678,N_3361,N_3307);
or U4679 (N_4679,N_3097,N_2815);
nor U4680 (N_4680,N_3791,N_3306);
nor U4681 (N_4681,N_2182,N_3467);
or U4682 (N_4682,N_2367,N_2599);
and U4683 (N_4683,N_3980,N_2706);
and U4684 (N_4684,N_3416,N_2224);
nand U4685 (N_4685,N_2551,N_3411);
or U4686 (N_4686,N_2303,N_2087);
nand U4687 (N_4687,N_3024,N_3673);
or U4688 (N_4688,N_2388,N_2558);
nor U4689 (N_4689,N_2240,N_3541);
nand U4690 (N_4690,N_2368,N_3822);
nand U4691 (N_4691,N_3085,N_3863);
nand U4692 (N_4692,N_3571,N_3678);
nor U4693 (N_4693,N_2394,N_3238);
and U4694 (N_4694,N_2478,N_2618);
or U4695 (N_4695,N_3475,N_3799);
nor U4696 (N_4696,N_3685,N_2042);
nor U4697 (N_4697,N_3554,N_3425);
nor U4698 (N_4698,N_3610,N_2171);
nand U4699 (N_4699,N_3407,N_2410);
nand U4700 (N_4700,N_3689,N_2450);
nor U4701 (N_4701,N_2717,N_2252);
and U4702 (N_4702,N_3163,N_2936);
or U4703 (N_4703,N_2324,N_2250);
and U4704 (N_4704,N_3098,N_2790);
nor U4705 (N_4705,N_3397,N_3485);
and U4706 (N_4706,N_3582,N_2532);
nor U4707 (N_4707,N_2715,N_2283);
and U4708 (N_4708,N_3710,N_3746);
nor U4709 (N_4709,N_3178,N_2067);
or U4710 (N_4710,N_3603,N_3345);
or U4711 (N_4711,N_3234,N_3133);
or U4712 (N_4712,N_2774,N_3132);
or U4713 (N_4713,N_2677,N_2923);
nor U4714 (N_4714,N_2077,N_2580);
nor U4715 (N_4715,N_3775,N_2998);
or U4716 (N_4716,N_2006,N_2438);
and U4717 (N_4717,N_2204,N_3410);
and U4718 (N_4718,N_2684,N_3774);
nor U4719 (N_4719,N_2593,N_3721);
nor U4720 (N_4720,N_2942,N_2471);
xor U4721 (N_4721,N_2489,N_3401);
xor U4722 (N_4722,N_3171,N_2413);
nor U4723 (N_4723,N_3890,N_3944);
nor U4724 (N_4724,N_3253,N_3103);
nor U4725 (N_4725,N_3661,N_3090);
nand U4726 (N_4726,N_3166,N_3619);
xor U4727 (N_4727,N_3112,N_2882);
nand U4728 (N_4728,N_3027,N_2806);
and U4729 (N_4729,N_3379,N_2346);
nor U4730 (N_4730,N_2132,N_2807);
and U4731 (N_4731,N_2778,N_3941);
and U4732 (N_4732,N_2931,N_3409);
nor U4733 (N_4733,N_2741,N_3059);
nand U4734 (N_4734,N_3959,N_2369);
nand U4735 (N_4735,N_2485,N_3526);
and U4736 (N_4736,N_3130,N_3902);
nand U4737 (N_4737,N_2922,N_3722);
nand U4738 (N_4738,N_2607,N_2234);
and U4739 (N_4739,N_2830,N_3275);
nor U4740 (N_4740,N_3805,N_3157);
and U4741 (N_4741,N_3322,N_2513);
and U4742 (N_4742,N_3923,N_2820);
and U4743 (N_4743,N_3477,N_2159);
or U4744 (N_4744,N_3203,N_2809);
nand U4745 (N_4745,N_2173,N_3745);
and U4746 (N_4746,N_2084,N_3331);
or U4747 (N_4747,N_2026,N_2890);
or U4748 (N_4748,N_2144,N_2137);
and U4749 (N_4749,N_2414,N_2140);
or U4750 (N_4750,N_3534,N_2300);
nand U4751 (N_4751,N_3466,N_3308);
and U4752 (N_4752,N_2199,N_2295);
and U4753 (N_4753,N_3285,N_3262);
and U4754 (N_4754,N_2231,N_2507);
and U4755 (N_4755,N_2657,N_3839);
nor U4756 (N_4756,N_2797,N_2326);
and U4757 (N_4757,N_3270,N_3054);
nand U4758 (N_4758,N_3854,N_2114);
nor U4759 (N_4759,N_3807,N_2451);
nand U4760 (N_4760,N_3402,N_3667);
or U4761 (N_4761,N_2169,N_2467);
or U4762 (N_4762,N_2749,N_2210);
or U4763 (N_4763,N_2751,N_2195);
nor U4764 (N_4764,N_3373,N_3940);
or U4765 (N_4765,N_3165,N_3050);
nand U4766 (N_4766,N_3074,N_3435);
and U4767 (N_4767,N_2420,N_3159);
nor U4768 (N_4768,N_3542,N_3950);
and U4769 (N_4769,N_2899,N_3215);
or U4770 (N_4770,N_3516,N_2776);
or U4771 (N_4771,N_3889,N_2754);
nor U4772 (N_4772,N_2562,N_2377);
nand U4773 (N_4773,N_3723,N_3233);
and U4774 (N_4774,N_2688,N_2867);
nand U4775 (N_4775,N_2382,N_2999);
or U4776 (N_4776,N_2787,N_2272);
nand U4777 (N_4777,N_2433,N_3448);
nand U4778 (N_4778,N_3053,N_3668);
nor U4779 (N_4779,N_3081,N_2616);
nor U4780 (N_4780,N_3412,N_3278);
nor U4781 (N_4781,N_2092,N_3953);
nor U4782 (N_4782,N_3609,N_2267);
nor U4783 (N_4783,N_2784,N_2473);
and U4784 (N_4784,N_3023,N_2109);
or U4785 (N_4785,N_2449,N_3798);
nand U4786 (N_4786,N_3052,N_3903);
nand U4787 (N_4787,N_3555,N_3641);
nor U4788 (N_4788,N_3811,N_3813);
nor U4789 (N_4789,N_3556,N_2065);
and U4790 (N_4790,N_3473,N_3524);
nor U4791 (N_4791,N_2819,N_2932);
and U4792 (N_4792,N_2568,N_2786);
or U4793 (N_4793,N_2460,N_3128);
nor U4794 (N_4794,N_2187,N_3111);
or U4795 (N_4795,N_2995,N_3546);
nor U4796 (N_4796,N_3020,N_2570);
nor U4797 (N_4797,N_3297,N_2047);
nand U4798 (N_4798,N_3414,N_3104);
or U4799 (N_4799,N_2509,N_2311);
and U4800 (N_4800,N_3718,N_2954);
nand U4801 (N_4801,N_2624,N_2705);
nand U4802 (N_4802,N_3302,N_3125);
nor U4803 (N_4803,N_3969,N_3965);
and U4804 (N_4804,N_3518,N_2331);
and U4805 (N_4805,N_2649,N_3463);
and U4806 (N_4806,N_2285,N_2611);
nand U4807 (N_4807,N_2423,N_3566);
or U4808 (N_4808,N_2685,N_3358);
nand U4809 (N_4809,N_3084,N_3583);
nor U4810 (N_4810,N_3426,N_2821);
nor U4811 (N_4811,N_3115,N_2959);
nor U4812 (N_4812,N_3749,N_3692);
nand U4813 (N_4813,N_3709,N_2988);
or U4814 (N_4814,N_3046,N_2322);
nand U4815 (N_4815,N_3100,N_2107);
and U4816 (N_4816,N_3815,N_3856);
nand U4817 (N_4817,N_3808,N_2242);
or U4818 (N_4818,N_3200,N_3267);
nand U4819 (N_4819,N_3427,N_3744);
nor U4820 (N_4820,N_3596,N_3354);
nor U4821 (N_4821,N_3728,N_3327);
nor U4822 (N_4822,N_2319,N_3261);
nor U4823 (N_4823,N_3734,N_3706);
nor U4824 (N_4824,N_3797,N_2488);
nand U4825 (N_4825,N_3691,N_2083);
and U4826 (N_4826,N_3372,N_2866);
or U4827 (N_4827,N_3021,N_3806);
and U4828 (N_4828,N_3260,N_2620);
nand U4829 (N_4829,N_2973,N_2086);
nand U4830 (N_4830,N_2399,N_2848);
and U4831 (N_4831,N_3979,N_3812);
and U4832 (N_4832,N_2233,N_2913);
nor U4833 (N_4833,N_3574,N_3639);
and U4834 (N_4834,N_2505,N_2392);
nand U4835 (N_4835,N_2576,N_3506);
nand U4836 (N_4836,N_2415,N_3055);
nor U4837 (N_4837,N_3974,N_3633);
xnor U4838 (N_4838,N_2429,N_3380);
and U4839 (N_4839,N_3880,N_3150);
and U4840 (N_4840,N_3704,N_3036);
or U4841 (N_4841,N_2842,N_3257);
or U4842 (N_4842,N_2453,N_2230);
nand U4843 (N_4843,N_3386,N_3256);
nand U4844 (N_4844,N_3042,N_2348);
and U4845 (N_4845,N_2383,N_2547);
xor U4846 (N_4846,N_2155,N_3817);
nor U4847 (N_4847,N_2227,N_3272);
nor U4848 (N_4848,N_3553,N_3277);
and U4849 (N_4849,N_2469,N_3515);
and U4850 (N_4850,N_3832,N_3716);
and U4851 (N_4851,N_2286,N_2176);
or U4852 (N_4852,N_2014,N_2120);
or U4853 (N_4853,N_2292,N_3781);
and U4854 (N_4854,N_3795,N_2223);
nand U4855 (N_4855,N_3061,N_3881);
nand U4856 (N_4856,N_2012,N_2915);
nor U4857 (N_4857,N_2948,N_2479);
nand U4858 (N_4858,N_2672,N_2481);
nand U4859 (N_4859,N_2128,N_3341);
nand U4860 (N_4860,N_2767,N_3312);
or U4861 (N_4861,N_3244,N_3602);
or U4862 (N_4862,N_2443,N_2097);
nand U4863 (N_4863,N_3675,N_2873);
nor U4864 (N_4864,N_3724,N_3381);
nand U4865 (N_4865,N_3730,N_3214);
and U4866 (N_4866,N_3548,N_3964);
nor U4867 (N_4867,N_2363,N_3249);
and U4868 (N_4868,N_2135,N_2268);
nand U4869 (N_4869,N_3470,N_3026);
xnor U4870 (N_4870,N_3560,N_2052);
or U4871 (N_4871,N_3304,N_2428);
nor U4872 (N_4872,N_2222,N_3088);
nand U4873 (N_4873,N_3772,N_3776);
or U4874 (N_4874,N_2412,N_2323);
and U4875 (N_4875,N_2470,N_2400);
or U4876 (N_4876,N_3743,N_2112);
and U4877 (N_4877,N_2585,N_2594);
nor U4878 (N_4878,N_2769,N_3254);
nor U4879 (N_4879,N_3538,N_3833);
nand U4880 (N_4880,N_3335,N_3671);
or U4881 (N_4881,N_3196,N_3872);
and U4882 (N_4882,N_2860,N_3095);
or U4883 (N_4883,N_3656,N_2977);
nor U4884 (N_4884,N_3758,N_2946);
and U4885 (N_4885,N_2476,N_3802);
or U4886 (N_4886,N_3591,N_3896);
and U4887 (N_4887,N_3765,N_2379);
or U4888 (N_4888,N_2431,N_2880);
nor U4889 (N_4889,N_2278,N_3211);
nand U4890 (N_4890,N_3019,N_3149);
or U4891 (N_4891,N_2579,N_3539);
and U4892 (N_4892,N_3998,N_2238);
or U4893 (N_4893,N_2978,N_2905);
nor U4894 (N_4894,N_3720,N_2596);
and U4895 (N_4895,N_2384,N_3139);
or U4896 (N_4896,N_3649,N_3225);
nand U4897 (N_4897,N_2708,N_3604);
or U4898 (N_4898,N_3247,N_2533);
xnor U4899 (N_4899,N_3041,N_3441);
or U4900 (N_4900,N_3064,N_2644);
nor U4901 (N_4901,N_2695,N_2288);
and U4902 (N_4902,N_2274,N_2448);
nand U4903 (N_4903,N_2253,N_3973);
nor U4904 (N_4904,N_3848,N_2432);
and U4905 (N_4905,N_3531,N_2701);
and U4906 (N_4906,N_3892,N_2711);
nand U4907 (N_4907,N_2897,N_2938);
and U4908 (N_4908,N_2636,N_2373);
or U4909 (N_4909,N_3834,N_2664);
or U4910 (N_4910,N_3001,N_3825);
nand U4911 (N_4911,N_2281,N_3922);
nand U4912 (N_4912,N_3666,N_3230);
nor U4913 (N_4913,N_3859,N_3945);
nand U4914 (N_4914,N_3955,N_2983);
nor U4915 (N_4915,N_2100,N_3600);
nor U4916 (N_4916,N_2650,N_3138);
xnor U4917 (N_4917,N_3316,N_3662);
nor U4918 (N_4918,N_3458,N_2113);
nand U4919 (N_4919,N_3181,N_3332);
nand U4920 (N_4920,N_2981,N_3810);
nand U4921 (N_4921,N_2404,N_3491);
nor U4922 (N_4922,N_2641,N_2800);
or U4923 (N_4923,N_3141,N_2458);
and U4924 (N_4924,N_2023,N_3478);
nand U4925 (N_4925,N_2126,N_3440);
or U4926 (N_4926,N_3512,N_3943);
nor U4927 (N_4927,N_3390,N_3708);
nand U4928 (N_4928,N_3871,N_3266);
and U4929 (N_4929,N_3318,N_3780);
nand U4930 (N_4930,N_2329,N_3646);
or U4931 (N_4931,N_2953,N_2546);
nor U4932 (N_4932,N_3642,N_3351);
and U4933 (N_4933,N_2407,N_2081);
or U4934 (N_4934,N_2680,N_3406);
and U4935 (N_4935,N_2564,N_2627);
nand U4936 (N_4936,N_2349,N_3330);
nand U4937 (N_4937,N_2297,N_3739);
and U4938 (N_4938,N_3321,N_2950);
nand U4939 (N_4939,N_3837,N_2986);
and U4940 (N_4940,N_3939,N_2595);
xnor U4941 (N_4941,N_2958,N_3170);
or U4942 (N_4942,N_3037,N_3363);
xnor U4943 (N_4943,N_2822,N_3099);
nand U4944 (N_4944,N_2682,N_2886);
or U4945 (N_4945,N_3480,N_2454);
nand U4946 (N_4946,N_3195,N_2892);
or U4947 (N_4947,N_2022,N_2871);
and U4948 (N_4948,N_3273,N_2765);
nor U4949 (N_4949,N_3967,N_3135);
nand U4950 (N_4950,N_2992,N_2879);
and U4951 (N_4951,N_2826,N_2235);
nor U4952 (N_4952,N_3674,N_3201);
or U4953 (N_4953,N_3578,N_2063);
and U4954 (N_4954,N_2960,N_2370);
nor U4955 (N_4955,N_3698,N_2118);
and U4956 (N_4956,N_2566,N_3177);
or U4957 (N_4957,N_2737,N_3148);
and U4958 (N_4958,N_3952,N_3503);
nand U4959 (N_4959,N_3000,N_2422);
and U4960 (N_4960,N_3768,N_2264);
nand U4961 (N_4961,N_2461,N_2396);
or U4962 (N_4962,N_3900,N_3696);
nor U4963 (N_4963,N_3823,N_3245);
nand U4964 (N_4964,N_2812,N_2976);
nand U4965 (N_4965,N_3615,N_2305);
nor U4966 (N_4966,N_3465,N_2663);
nand U4967 (N_4967,N_3819,N_2788);
nor U4968 (N_4968,N_3108,N_3816);
or U4969 (N_4969,N_3613,N_2704);
nand U4970 (N_4970,N_2673,N_2355);
or U4971 (N_4971,N_2971,N_2203);
nand U4972 (N_4972,N_2702,N_2515);
or U4973 (N_4973,N_3310,N_3963);
or U4974 (N_4974,N_2575,N_3782);
or U4975 (N_4975,N_2623,N_3933);
nor U4976 (N_4976,N_2838,N_3895);
nand U4977 (N_4977,N_3910,N_2647);
nor U4978 (N_4978,N_2474,N_2362);
or U4979 (N_4979,N_3009,N_2646);
or U4980 (N_4980,N_3527,N_3047);
nand U4981 (N_4981,N_3032,N_3664);
nor U4982 (N_4982,N_3783,N_3340);
and U4983 (N_4983,N_3056,N_2241);
nor U4984 (N_4984,N_3391,N_3951);
and U4985 (N_4985,N_3158,N_2760);
nand U4986 (N_4986,N_2184,N_3789);
and U4987 (N_4987,N_3246,N_2630);
nand U4988 (N_4988,N_2637,N_3347);
nor U4989 (N_4989,N_2834,N_2202);
or U4990 (N_4990,N_2823,N_3954);
nand U4991 (N_4991,N_2350,N_3993);
and U4992 (N_4992,N_2895,N_2342);
nand U4993 (N_4993,N_2001,N_3551);
nand U4994 (N_4994,N_2027,N_2775);
nand U4995 (N_4995,N_2696,N_3737);
and U4996 (N_4996,N_3732,N_3701);
or U4997 (N_4997,N_2061,N_2966);
and U4998 (N_4998,N_3439,N_3471);
or U4999 (N_4999,N_2979,N_3916);
nor U5000 (N_5000,N_2694,N_2303);
nand U5001 (N_5001,N_3722,N_3569);
and U5002 (N_5002,N_3891,N_3139);
or U5003 (N_5003,N_3122,N_3692);
and U5004 (N_5004,N_3011,N_2715);
or U5005 (N_5005,N_3066,N_3554);
nand U5006 (N_5006,N_3119,N_3785);
and U5007 (N_5007,N_3721,N_3508);
and U5008 (N_5008,N_2903,N_3604);
and U5009 (N_5009,N_3960,N_2432);
xnor U5010 (N_5010,N_2855,N_3438);
and U5011 (N_5011,N_2973,N_3615);
nand U5012 (N_5012,N_3300,N_3420);
nor U5013 (N_5013,N_3145,N_3862);
nor U5014 (N_5014,N_2895,N_3158);
nor U5015 (N_5015,N_3993,N_2405);
nand U5016 (N_5016,N_2706,N_3090);
nor U5017 (N_5017,N_3065,N_3114);
nand U5018 (N_5018,N_2412,N_3508);
nor U5019 (N_5019,N_2802,N_2393);
or U5020 (N_5020,N_3550,N_2035);
and U5021 (N_5021,N_3949,N_3962);
and U5022 (N_5022,N_2808,N_2929);
nand U5023 (N_5023,N_2901,N_3413);
or U5024 (N_5024,N_2042,N_3152);
or U5025 (N_5025,N_3531,N_2359);
and U5026 (N_5026,N_3833,N_2661);
nor U5027 (N_5027,N_3588,N_2303);
or U5028 (N_5028,N_3556,N_3748);
nand U5029 (N_5029,N_3558,N_3721);
nand U5030 (N_5030,N_2282,N_2884);
nand U5031 (N_5031,N_2692,N_2837);
nor U5032 (N_5032,N_3582,N_3187);
nor U5033 (N_5033,N_3100,N_2593);
nand U5034 (N_5034,N_2819,N_3344);
or U5035 (N_5035,N_3990,N_3248);
or U5036 (N_5036,N_3978,N_2128);
and U5037 (N_5037,N_3827,N_2672);
or U5038 (N_5038,N_3420,N_2182);
or U5039 (N_5039,N_3253,N_3282);
or U5040 (N_5040,N_2876,N_3705);
xor U5041 (N_5041,N_3505,N_3903);
or U5042 (N_5042,N_2598,N_2550);
and U5043 (N_5043,N_2882,N_3590);
nand U5044 (N_5044,N_2565,N_3211);
nor U5045 (N_5045,N_2113,N_2659);
and U5046 (N_5046,N_2514,N_2188);
or U5047 (N_5047,N_3976,N_2380);
nand U5048 (N_5048,N_3974,N_3456);
or U5049 (N_5049,N_3196,N_3418);
nor U5050 (N_5050,N_2296,N_2206);
and U5051 (N_5051,N_3874,N_3113);
or U5052 (N_5052,N_2758,N_2500);
nand U5053 (N_5053,N_3919,N_2896);
nor U5054 (N_5054,N_2501,N_2308);
and U5055 (N_5055,N_3710,N_3008);
and U5056 (N_5056,N_2988,N_3967);
and U5057 (N_5057,N_2553,N_2836);
or U5058 (N_5058,N_2199,N_3474);
nand U5059 (N_5059,N_2156,N_3753);
and U5060 (N_5060,N_2812,N_2489);
or U5061 (N_5061,N_3015,N_3313);
nor U5062 (N_5062,N_2342,N_2400);
nor U5063 (N_5063,N_2750,N_3623);
nor U5064 (N_5064,N_3955,N_3642);
or U5065 (N_5065,N_3463,N_3272);
nor U5066 (N_5066,N_3300,N_2820);
or U5067 (N_5067,N_3848,N_2173);
nor U5068 (N_5068,N_2557,N_3694);
xnor U5069 (N_5069,N_3043,N_3095);
nand U5070 (N_5070,N_2590,N_2283);
or U5071 (N_5071,N_3223,N_3631);
or U5072 (N_5072,N_3601,N_3689);
nand U5073 (N_5073,N_3629,N_2404);
and U5074 (N_5074,N_2305,N_3773);
and U5075 (N_5075,N_2588,N_3568);
nor U5076 (N_5076,N_2638,N_2645);
nand U5077 (N_5077,N_2166,N_2255);
and U5078 (N_5078,N_2171,N_2178);
or U5079 (N_5079,N_3621,N_2196);
nor U5080 (N_5080,N_2008,N_3003);
or U5081 (N_5081,N_3427,N_2578);
nor U5082 (N_5082,N_2928,N_2836);
nand U5083 (N_5083,N_3659,N_3532);
nor U5084 (N_5084,N_3191,N_2967);
nor U5085 (N_5085,N_3904,N_2949);
and U5086 (N_5086,N_2398,N_2793);
or U5087 (N_5087,N_3289,N_2920);
or U5088 (N_5088,N_3828,N_3442);
and U5089 (N_5089,N_2644,N_2297);
nor U5090 (N_5090,N_2623,N_3889);
and U5091 (N_5091,N_2440,N_3647);
nor U5092 (N_5092,N_2382,N_2706);
and U5093 (N_5093,N_3416,N_2020);
and U5094 (N_5094,N_3142,N_2507);
nor U5095 (N_5095,N_3305,N_2499);
nand U5096 (N_5096,N_2303,N_3425);
xnor U5097 (N_5097,N_2948,N_3260);
nor U5098 (N_5098,N_3021,N_3370);
xor U5099 (N_5099,N_3262,N_3590);
or U5100 (N_5100,N_3738,N_2727);
nand U5101 (N_5101,N_2403,N_3175);
nand U5102 (N_5102,N_3417,N_3138);
or U5103 (N_5103,N_3799,N_3269);
and U5104 (N_5104,N_2025,N_2449);
nor U5105 (N_5105,N_3813,N_2256);
nand U5106 (N_5106,N_3735,N_2564);
nor U5107 (N_5107,N_2478,N_2906);
nor U5108 (N_5108,N_2875,N_2238);
nor U5109 (N_5109,N_3918,N_3437);
nand U5110 (N_5110,N_2499,N_2665);
and U5111 (N_5111,N_3056,N_2897);
xor U5112 (N_5112,N_2489,N_2916);
nor U5113 (N_5113,N_2246,N_2939);
or U5114 (N_5114,N_3457,N_2167);
nand U5115 (N_5115,N_2334,N_2472);
nor U5116 (N_5116,N_2434,N_3229);
nand U5117 (N_5117,N_3448,N_2326);
and U5118 (N_5118,N_2175,N_3982);
and U5119 (N_5119,N_2351,N_3484);
nor U5120 (N_5120,N_3904,N_2019);
and U5121 (N_5121,N_2480,N_2695);
nand U5122 (N_5122,N_2354,N_3280);
nand U5123 (N_5123,N_2096,N_2564);
and U5124 (N_5124,N_2644,N_2629);
and U5125 (N_5125,N_2060,N_2809);
xnor U5126 (N_5126,N_2441,N_3693);
nand U5127 (N_5127,N_2766,N_3587);
or U5128 (N_5128,N_3367,N_3351);
nand U5129 (N_5129,N_2293,N_3009);
and U5130 (N_5130,N_3909,N_3212);
nand U5131 (N_5131,N_3334,N_3452);
or U5132 (N_5132,N_2238,N_2063);
or U5133 (N_5133,N_3170,N_3703);
nor U5134 (N_5134,N_3967,N_2915);
nand U5135 (N_5135,N_2451,N_3729);
or U5136 (N_5136,N_2919,N_2881);
nand U5137 (N_5137,N_2298,N_3941);
xnor U5138 (N_5138,N_3080,N_3528);
or U5139 (N_5139,N_2440,N_3691);
and U5140 (N_5140,N_3931,N_3490);
nor U5141 (N_5141,N_2745,N_2764);
and U5142 (N_5142,N_3706,N_3710);
nand U5143 (N_5143,N_2538,N_2127);
nand U5144 (N_5144,N_3236,N_2017);
nor U5145 (N_5145,N_3012,N_2229);
nor U5146 (N_5146,N_3336,N_2773);
nand U5147 (N_5147,N_3516,N_2227);
nand U5148 (N_5148,N_3255,N_3405);
nor U5149 (N_5149,N_3893,N_3355);
nor U5150 (N_5150,N_3405,N_3632);
nand U5151 (N_5151,N_2172,N_2260);
nand U5152 (N_5152,N_2994,N_3908);
nand U5153 (N_5153,N_2215,N_2147);
and U5154 (N_5154,N_3119,N_2395);
and U5155 (N_5155,N_2299,N_2048);
nor U5156 (N_5156,N_2852,N_3654);
and U5157 (N_5157,N_2098,N_3270);
nor U5158 (N_5158,N_3676,N_2187);
nor U5159 (N_5159,N_3599,N_3210);
and U5160 (N_5160,N_3757,N_3477);
nand U5161 (N_5161,N_2502,N_3563);
or U5162 (N_5162,N_2439,N_3559);
nand U5163 (N_5163,N_3713,N_2154);
nand U5164 (N_5164,N_3343,N_3896);
and U5165 (N_5165,N_3783,N_2161);
nor U5166 (N_5166,N_2148,N_3632);
nor U5167 (N_5167,N_2041,N_3695);
and U5168 (N_5168,N_3300,N_2662);
nor U5169 (N_5169,N_3156,N_3555);
and U5170 (N_5170,N_3426,N_2008);
nand U5171 (N_5171,N_3898,N_2696);
and U5172 (N_5172,N_3097,N_2154);
and U5173 (N_5173,N_3576,N_3577);
and U5174 (N_5174,N_3829,N_2762);
and U5175 (N_5175,N_2952,N_2930);
nand U5176 (N_5176,N_2970,N_3447);
nor U5177 (N_5177,N_3270,N_3157);
nand U5178 (N_5178,N_3709,N_2785);
and U5179 (N_5179,N_2388,N_2203);
xnor U5180 (N_5180,N_2137,N_3821);
nand U5181 (N_5181,N_2495,N_3175);
or U5182 (N_5182,N_3779,N_2021);
or U5183 (N_5183,N_2297,N_2152);
or U5184 (N_5184,N_3873,N_2971);
or U5185 (N_5185,N_2679,N_3503);
and U5186 (N_5186,N_2041,N_3457);
nor U5187 (N_5187,N_2695,N_2740);
or U5188 (N_5188,N_2437,N_2758);
or U5189 (N_5189,N_2100,N_3563);
and U5190 (N_5190,N_2700,N_2826);
or U5191 (N_5191,N_2859,N_2923);
nor U5192 (N_5192,N_2776,N_3866);
or U5193 (N_5193,N_3606,N_3461);
or U5194 (N_5194,N_3031,N_2654);
or U5195 (N_5195,N_2670,N_2570);
or U5196 (N_5196,N_2179,N_2950);
and U5197 (N_5197,N_2310,N_2146);
and U5198 (N_5198,N_3538,N_2962);
and U5199 (N_5199,N_2823,N_3792);
nand U5200 (N_5200,N_2643,N_2345);
or U5201 (N_5201,N_2381,N_3430);
or U5202 (N_5202,N_2333,N_3662);
and U5203 (N_5203,N_3204,N_3996);
nand U5204 (N_5204,N_3454,N_3050);
and U5205 (N_5205,N_2179,N_3485);
nor U5206 (N_5206,N_3926,N_2247);
and U5207 (N_5207,N_2552,N_3390);
and U5208 (N_5208,N_3780,N_3931);
nand U5209 (N_5209,N_3166,N_2805);
nand U5210 (N_5210,N_2732,N_3396);
nor U5211 (N_5211,N_2875,N_2559);
and U5212 (N_5212,N_3383,N_3072);
or U5213 (N_5213,N_2419,N_3336);
nand U5214 (N_5214,N_2060,N_3622);
nand U5215 (N_5215,N_3507,N_2345);
nor U5216 (N_5216,N_2882,N_2987);
nor U5217 (N_5217,N_2738,N_3667);
nand U5218 (N_5218,N_3204,N_2423);
nand U5219 (N_5219,N_3826,N_3661);
or U5220 (N_5220,N_2073,N_3821);
and U5221 (N_5221,N_3066,N_3505);
xnor U5222 (N_5222,N_3317,N_2049);
or U5223 (N_5223,N_3811,N_2263);
and U5224 (N_5224,N_2372,N_2572);
or U5225 (N_5225,N_2137,N_3305);
or U5226 (N_5226,N_3142,N_3487);
xnor U5227 (N_5227,N_3220,N_3131);
and U5228 (N_5228,N_2793,N_3146);
nor U5229 (N_5229,N_2075,N_2767);
and U5230 (N_5230,N_2880,N_3289);
nor U5231 (N_5231,N_2009,N_2325);
nor U5232 (N_5232,N_2283,N_2418);
and U5233 (N_5233,N_2867,N_2692);
or U5234 (N_5234,N_2106,N_3163);
nor U5235 (N_5235,N_3847,N_3803);
or U5236 (N_5236,N_2798,N_2832);
nor U5237 (N_5237,N_3224,N_2571);
nor U5238 (N_5238,N_3367,N_2543);
or U5239 (N_5239,N_2638,N_3050);
nor U5240 (N_5240,N_2117,N_2655);
nand U5241 (N_5241,N_2371,N_2896);
and U5242 (N_5242,N_2593,N_3033);
nand U5243 (N_5243,N_2754,N_3209);
nand U5244 (N_5244,N_2784,N_3089);
nand U5245 (N_5245,N_2192,N_2282);
and U5246 (N_5246,N_2867,N_3119);
nand U5247 (N_5247,N_3864,N_3704);
or U5248 (N_5248,N_3079,N_3080);
nor U5249 (N_5249,N_3844,N_2022);
and U5250 (N_5250,N_2291,N_3222);
or U5251 (N_5251,N_2789,N_3641);
or U5252 (N_5252,N_2829,N_2483);
and U5253 (N_5253,N_3337,N_2226);
or U5254 (N_5254,N_3394,N_3513);
nand U5255 (N_5255,N_3477,N_3220);
or U5256 (N_5256,N_3870,N_2787);
and U5257 (N_5257,N_2697,N_3168);
and U5258 (N_5258,N_2632,N_2034);
or U5259 (N_5259,N_3158,N_2457);
or U5260 (N_5260,N_2959,N_2374);
nor U5261 (N_5261,N_2407,N_2822);
or U5262 (N_5262,N_2979,N_2678);
nand U5263 (N_5263,N_3976,N_2547);
or U5264 (N_5264,N_2377,N_2778);
nor U5265 (N_5265,N_2921,N_3098);
nand U5266 (N_5266,N_2246,N_3585);
nor U5267 (N_5267,N_3908,N_3983);
nand U5268 (N_5268,N_3323,N_3669);
nor U5269 (N_5269,N_3376,N_2150);
and U5270 (N_5270,N_3718,N_3908);
or U5271 (N_5271,N_3614,N_3887);
nor U5272 (N_5272,N_2773,N_2563);
nand U5273 (N_5273,N_2626,N_2074);
or U5274 (N_5274,N_2273,N_3998);
nor U5275 (N_5275,N_2743,N_3427);
nor U5276 (N_5276,N_3936,N_2890);
and U5277 (N_5277,N_3846,N_2159);
nand U5278 (N_5278,N_2399,N_3883);
nor U5279 (N_5279,N_3980,N_2744);
nand U5280 (N_5280,N_2889,N_3913);
nor U5281 (N_5281,N_3908,N_2899);
and U5282 (N_5282,N_2628,N_3369);
nand U5283 (N_5283,N_2338,N_2929);
or U5284 (N_5284,N_3548,N_3186);
nor U5285 (N_5285,N_3813,N_3549);
nor U5286 (N_5286,N_3365,N_2870);
xnor U5287 (N_5287,N_3430,N_2116);
and U5288 (N_5288,N_2728,N_2697);
nand U5289 (N_5289,N_3266,N_2427);
and U5290 (N_5290,N_3070,N_2272);
nor U5291 (N_5291,N_2383,N_2171);
and U5292 (N_5292,N_3606,N_3119);
xnor U5293 (N_5293,N_3295,N_3190);
or U5294 (N_5294,N_2471,N_2914);
nor U5295 (N_5295,N_2130,N_3908);
and U5296 (N_5296,N_2663,N_3654);
nor U5297 (N_5297,N_2429,N_3581);
and U5298 (N_5298,N_2285,N_2843);
nand U5299 (N_5299,N_3773,N_2111);
xnor U5300 (N_5300,N_3019,N_2232);
nand U5301 (N_5301,N_3871,N_3289);
nand U5302 (N_5302,N_3701,N_3220);
nand U5303 (N_5303,N_3918,N_2836);
nand U5304 (N_5304,N_3854,N_3007);
nand U5305 (N_5305,N_3871,N_3922);
and U5306 (N_5306,N_2463,N_3337);
nor U5307 (N_5307,N_2233,N_3917);
or U5308 (N_5308,N_3268,N_2567);
nand U5309 (N_5309,N_3391,N_3944);
or U5310 (N_5310,N_2795,N_3165);
nand U5311 (N_5311,N_3750,N_3606);
nor U5312 (N_5312,N_3700,N_3573);
or U5313 (N_5313,N_2534,N_3219);
or U5314 (N_5314,N_2224,N_2989);
or U5315 (N_5315,N_2342,N_3886);
nand U5316 (N_5316,N_3881,N_3551);
nand U5317 (N_5317,N_3134,N_3768);
and U5318 (N_5318,N_2308,N_2339);
and U5319 (N_5319,N_2447,N_2070);
nand U5320 (N_5320,N_3638,N_2938);
and U5321 (N_5321,N_3980,N_2350);
nand U5322 (N_5322,N_3889,N_3178);
or U5323 (N_5323,N_3338,N_2243);
nand U5324 (N_5324,N_3746,N_3651);
nand U5325 (N_5325,N_3642,N_2861);
or U5326 (N_5326,N_3530,N_3610);
nand U5327 (N_5327,N_3317,N_3629);
or U5328 (N_5328,N_3988,N_3914);
nand U5329 (N_5329,N_2976,N_3587);
and U5330 (N_5330,N_3122,N_3088);
nand U5331 (N_5331,N_2899,N_2189);
nand U5332 (N_5332,N_2382,N_2600);
nand U5333 (N_5333,N_2561,N_2220);
or U5334 (N_5334,N_3876,N_2553);
and U5335 (N_5335,N_2541,N_3858);
xnor U5336 (N_5336,N_2982,N_3257);
and U5337 (N_5337,N_2785,N_2915);
nand U5338 (N_5338,N_3054,N_2050);
nor U5339 (N_5339,N_2987,N_2818);
and U5340 (N_5340,N_2636,N_2908);
nand U5341 (N_5341,N_3921,N_3586);
nor U5342 (N_5342,N_2013,N_2681);
xor U5343 (N_5343,N_2711,N_2643);
and U5344 (N_5344,N_2431,N_3153);
or U5345 (N_5345,N_2095,N_3224);
nand U5346 (N_5346,N_3823,N_3099);
and U5347 (N_5347,N_2627,N_2558);
nor U5348 (N_5348,N_2808,N_3669);
and U5349 (N_5349,N_2976,N_2983);
nor U5350 (N_5350,N_3767,N_2017);
xor U5351 (N_5351,N_2265,N_3064);
nand U5352 (N_5352,N_2130,N_3007);
and U5353 (N_5353,N_3617,N_3055);
nor U5354 (N_5354,N_3874,N_3630);
or U5355 (N_5355,N_3358,N_3460);
or U5356 (N_5356,N_2928,N_3891);
nand U5357 (N_5357,N_3249,N_3692);
and U5358 (N_5358,N_2617,N_3793);
and U5359 (N_5359,N_3339,N_3805);
or U5360 (N_5360,N_3848,N_2658);
nand U5361 (N_5361,N_2942,N_2281);
nor U5362 (N_5362,N_2793,N_2724);
or U5363 (N_5363,N_2061,N_2309);
or U5364 (N_5364,N_2154,N_3980);
nand U5365 (N_5365,N_3635,N_3762);
or U5366 (N_5366,N_3685,N_3073);
or U5367 (N_5367,N_2168,N_2130);
nand U5368 (N_5368,N_3028,N_2539);
nand U5369 (N_5369,N_3119,N_3668);
nand U5370 (N_5370,N_2482,N_2652);
and U5371 (N_5371,N_2636,N_2004);
or U5372 (N_5372,N_3369,N_2309);
or U5373 (N_5373,N_3556,N_3384);
and U5374 (N_5374,N_3974,N_3145);
nand U5375 (N_5375,N_2904,N_2261);
and U5376 (N_5376,N_2051,N_2901);
nand U5377 (N_5377,N_2073,N_3049);
xnor U5378 (N_5378,N_2495,N_3336);
or U5379 (N_5379,N_2018,N_3589);
and U5380 (N_5380,N_3313,N_3431);
nor U5381 (N_5381,N_3056,N_3303);
nand U5382 (N_5382,N_3445,N_2749);
or U5383 (N_5383,N_3988,N_3001);
xnor U5384 (N_5384,N_3469,N_2765);
and U5385 (N_5385,N_3435,N_2123);
nand U5386 (N_5386,N_3876,N_2522);
or U5387 (N_5387,N_2847,N_2926);
nand U5388 (N_5388,N_2815,N_3052);
or U5389 (N_5389,N_3671,N_2691);
nand U5390 (N_5390,N_3988,N_2716);
or U5391 (N_5391,N_2196,N_2946);
and U5392 (N_5392,N_2275,N_2756);
and U5393 (N_5393,N_3682,N_3950);
nand U5394 (N_5394,N_2774,N_2942);
xnor U5395 (N_5395,N_3322,N_2945);
and U5396 (N_5396,N_3165,N_3009);
and U5397 (N_5397,N_3881,N_3737);
nand U5398 (N_5398,N_3229,N_2339);
nor U5399 (N_5399,N_2704,N_2194);
nand U5400 (N_5400,N_3616,N_3229);
nand U5401 (N_5401,N_2294,N_3131);
or U5402 (N_5402,N_2175,N_2926);
nand U5403 (N_5403,N_3949,N_3137);
nor U5404 (N_5404,N_3861,N_3441);
nor U5405 (N_5405,N_3372,N_3724);
or U5406 (N_5406,N_2845,N_2519);
nand U5407 (N_5407,N_3454,N_3057);
or U5408 (N_5408,N_2799,N_3907);
and U5409 (N_5409,N_2357,N_3659);
and U5410 (N_5410,N_2287,N_2710);
nand U5411 (N_5411,N_3725,N_3991);
nand U5412 (N_5412,N_2726,N_3141);
nor U5413 (N_5413,N_2885,N_2005);
or U5414 (N_5414,N_2666,N_3317);
and U5415 (N_5415,N_2441,N_3222);
nor U5416 (N_5416,N_3792,N_2442);
and U5417 (N_5417,N_3920,N_2108);
and U5418 (N_5418,N_2071,N_2787);
and U5419 (N_5419,N_2345,N_3242);
or U5420 (N_5420,N_2208,N_2719);
or U5421 (N_5421,N_2902,N_2303);
xor U5422 (N_5422,N_2222,N_2464);
nor U5423 (N_5423,N_3248,N_3846);
nor U5424 (N_5424,N_2838,N_3848);
nand U5425 (N_5425,N_2003,N_2136);
nand U5426 (N_5426,N_2472,N_3032);
nor U5427 (N_5427,N_2116,N_3644);
nand U5428 (N_5428,N_3052,N_2284);
or U5429 (N_5429,N_2991,N_3246);
or U5430 (N_5430,N_2654,N_3575);
and U5431 (N_5431,N_2170,N_2221);
or U5432 (N_5432,N_2759,N_2667);
nor U5433 (N_5433,N_2819,N_2492);
or U5434 (N_5434,N_3020,N_3461);
and U5435 (N_5435,N_3648,N_3529);
or U5436 (N_5436,N_2096,N_3919);
or U5437 (N_5437,N_2010,N_2387);
and U5438 (N_5438,N_3017,N_3376);
nor U5439 (N_5439,N_2227,N_2764);
or U5440 (N_5440,N_3456,N_3150);
nor U5441 (N_5441,N_3850,N_3985);
and U5442 (N_5442,N_3322,N_3924);
or U5443 (N_5443,N_2995,N_3435);
nand U5444 (N_5444,N_2059,N_3377);
nand U5445 (N_5445,N_2495,N_2443);
nand U5446 (N_5446,N_2861,N_3266);
nand U5447 (N_5447,N_3082,N_3851);
or U5448 (N_5448,N_3533,N_3299);
and U5449 (N_5449,N_3345,N_3175);
or U5450 (N_5450,N_2417,N_2944);
xnor U5451 (N_5451,N_2742,N_3198);
and U5452 (N_5452,N_2365,N_2859);
or U5453 (N_5453,N_2003,N_2128);
and U5454 (N_5454,N_3570,N_2241);
and U5455 (N_5455,N_2447,N_3310);
nand U5456 (N_5456,N_2563,N_2050);
nor U5457 (N_5457,N_3393,N_3009);
nor U5458 (N_5458,N_3823,N_2914);
and U5459 (N_5459,N_3841,N_3248);
and U5460 (N_5460,N_3280,N_2021);
nand U5461 (N_5461,N_2550,N_2110);
nand U5462 (N_5462,N_2742,N_3906);
nand U5463 (N_5463,N_3728,N_3373);
nand U5464 (N_5464,N_3953,N_2872);
nand U5465 (N_5465,N_3463,N_3215);
and U5466 (N_5466,N_3278,N_2805);
or U5467 (N_5467,N_2848,N_2577);
nor U5468 (N_5468,N_2876,N_2463);
nand U5469 (N_5469,N_3149,N_2991);
nor U5470 (N_5470,N_2511,N_2082);
nor U5471 (N_5471,N_2980,N_3057);
nor U5472 (N_5472,N_2741,N_2594);
and U5473 (N_5473,N_2384,N_3639);
or U5474 (N_5474,N_3187,N_2934);
and U5475 (N_5475,N_3654,N_2505);
and U5476 (N_5476,N_3057,N_3389);
nor U5477 (N_5477,N_2868,N_3700);
nand U5478 (N_5478,N_2760,N_2580);
and U5479 (N_5479,N_2334,N_3343);
nand U5480 (N_5480,N_3496,N_3559);
nor U5481 (N_5481,N_3601,N_3264);
nand U5482 (N_5482,N_2521,N_3957);
nand U5483 (N_5483,N_2598,N_3714);
nand U5484 (N_5484,N_3722,N_3561);
nor U5485 (N_5485,N_3549,N_3758);
nor U5486 (N_5486,N_2772,N_3249);
or U5487 (N_5487,N_2252,N_3914);
nand U5488 (N_5488,N_3704,N_3638);
nand U5489 (N_5489,N_2553,N_3413);
nor U5490 (N_5490,N_2450,N_3483);
nand U5491 (N_5491,N_2485,N_3316);
nand U5492 (N_5492,N_3317,N_3652);
nor U5493 (N_5493,N_2954,N_3530);
nor U5494 (N_5494,N_3768,N_2775);
nand U5495 (N_5495,N_2965,N_3956);
nand U5496 (N_5496,N_2610,N_3584);
or U5497 (N_5497,N_2153,N_2596);
and U5498 (N_5498,N_3667,N_3846);
or U5499 (N_5499,N_2039,N_2195);
nor U5500 (N_5500,N_2000,N_2581);
xor U5501 (N_5501,N_2136,N_2038);
nor U5502 (N_5502,N_2094,N_3093);
nand U5503 (N_5503,N_2282,N_3123);
and U5504 (N_5504,N_2766,N_2648);
nand U5505 (N_5505,N_3610,N_3342);
xnor U5506 (N_5506,N_3937,N_2466);
nor U5507 (N_5507,N_3143,N_2611);
nand U5508 (N_5508,N_2702,N_3684);
nand U5509 (N_5509,N_3766,N_3364);
and U5510 (N_5510,N_2064,N_2297);
xor U5511 (N_5511,N_2468,N_3238);
nand U5512 (N_5512,N_2395,N_3831);
or U5513 (N_5513,N_3531,N_3223);
nand U5514 (N_5514,N_3057,N_3850);
nand U5515 (N_5515,N_3023,N_3366);
or U5516 (N_5516,N_3119,N_3506);
nor U5517 (N_5517,N_3970,N_2703);
or U5518 (N_5518,N_2694,N_2951);
nand U5519 (N_5519,N_2956,N_3493);
or U5520 (N_5520,N_2309,N_2446);
nor U5521 (N_5521,N_3364,N_2228);
nor U5522 (N_5522,N_3184,N_3117);
and U5523 (N_5523,N_2826,N_3671);
nor U5524 (N_5524,N_3711,N_3584);
nand U5525 (N_5525,N_3069,N_3186);
or U5526 (N_5526,N_2537,N_3436);
and U5527 (N_5527,N_2796,N_3237);
and U5528 (N_5528,N_3539,N_2251);
or U5529 (N_5529,N_2460,N_2050);
nor U5530 (N_5530,N_2622,N_3183);
or U5531 (N_5531,N_2173,N_2865);
or U5532 (N_5532,N_2979,N_3007);
or U5533 (N_5533,N_3912,N_3061);
or U5534 (N_5534,N_2032,N_2859);
nand U5535 (N_5535,N_2218,N_3869);
and U5536 (N_5536,N_2544,N_2297);
nor U5537 (N_5537,N_2007,N_3253);
and U5538 (N_5538,N_2759,N_2612);
nand U5539 (N_5539,N_2931,N_2939);
xor U5540 (N_5540,N_3816,N_2557);
or U5541 (N_5541,N_2048,N_2774);
nor U5542 (N_5542,N_3765,N_2264);
nand U5543 (N_5543,N_2889,N_3118);
or U5544 (N_5544,N_3341,N_2953);
nand U5545 (N_5545,N_3281,N_2633);
or U5546 (N_5546,N_2346,N_3626);
or U5547 (N_5547,N_3625,N_3578);
nand U5548 (N_5548,N_3840,N_2555);
nor U5549 (N_5549,N_2329,N_3462);
or U5550 (N_5550,N_3153,N_2831);
or U5551 (N_5551,N_2014,N_2556);
or U5552 (N_5552,N_2981,N_3187);
or U5553 (N_5553,N_2807,N_3886);
nand U5554 (N_5554,N_2958,N_3899);
and U5555 (N_5555,N_2188,N_3619);
nand U5556 (N_5556,N_2535,N_2312);
nor U5557 (N_5557,N_3295,N_2074);
xnor U5558 (N_5558,N_3216,N_2294);
or U5559 (N_5559,N_2063,N_2056);
nand U5560 (N_5560,N_2157,N_2397);
and U5561 (N_5561,N_2163,N_2929);
nand U5562 (N_5562,N_3464,N_3808);
or U5563 (N_5563,N_2659,N_3869);
and U5564 (N_5564,N_3709,N_2939);
or U5565 (N_5565,N_3270,N_2254);
nand U5566 (N_5566,N_2809,N_3284);
or U5567 (N_5567,N_2689,N_2632);
and U5568 (N_5568,N_3274,N_2553);
nand U5569 (N_5569,N_3526,N_2895);
nand U5570 (N_5570,N_3119,N_2184);
nor U5571 (N_5571,N_3460,N_3676);
nor U5572 (N_5572,N_2341,N_3854);
nand U5573 (N_5573,N_3799,N_2583);
or U5574 (N_5574,N_2364,N_3889);
nor U5575 (N_5575,N_3113,N_3958);
nand U5576 (N_5576,N_3221,N_3609);
nor U5577 (N_5577,N_2790,N_2796);
or U5578 (N_5578,N_2642,N_3357);
nor U5579 (N_5579,N_2711,N_3046);
nor U5580 (N_5580,N_2650,N_3595);
nor U5581 (N_5581,N_2027,N_3658);
and U5582 (N_5582,N_2905,N_3426);
and U5583 (N_5583,N_3101,N_2417);
and U5584 (N_5584,N_3633,N_3492);
nand U5585 (N_5585,N_3781,N_3385);
or U5586 (N_5586,N_2496,N_2806);
or U5587 (N_5587,N_3069,N_3679);
or U5588 (N_5588,N_2709,N_3636);
and U5589 (N_5589,N_2646,N_3842);
nand U5590 (N_5590,N_3077,N_3101);
nor U5591 (N_5591,N_2769,N_3535);
or U5592 (N_5592,N_3697,N_3463);
nor U5593 (N_5593,N_2425,N_3793);
nand U5594 (N_5594,N_3710,N_2162);
nor U5595 (N_5595,N_3274,N_3839);
and U5596 (N_5596,N_3910,N_3228);
and U5597 (N_5597,N_2092,N_2219);
and U5598 (N_5598,N_3081,N_3912);
nor U5599 (N_5599,N_3126,N_2417);
nand U5600 (N_5600,N_2583,N_2468);
nor U5601 (N_5601,N_3821,N_2450);
nor U5602 (N_5602,N_3282,N_3986);
or U5603 (N_5603,N_2564,N_2698);
and U5604 (N_5604,N_3772,N_3680);
or U5605 (N_5605,N_3522,N_2936);
xnor U5606 (N_5606,N_2072,N_3005);
and U5607 (N_5607,N_2386,N_2358);
and U5608 (N_5608,N_3375,N_3427);
nand U5609 (N_5609,N_2981,N_3034);
and U5610 (N_5610,N_2546,N_3868);
nor U5611 (N_5611,N_3437,N_3719);
or U5612 (N_5612,N_2386,N_3256);
nand U5613 (N_5613,N_2917,N_2968);
or U5614 (N_5614,N_2850,N_2893);
and U5615 (N_5615,N_2100,N_3851);
nand U5616 (N_5616,N_3925,N_3166);
xnor U5617 (N_5617,N_3631,N_2108);
or U5618 (N_5618,N_2649,N_2949);
and U5619 (N_5619,N_3846,N_2695);
nor U5620 (N_5620,N_3365,N_3203);
and U5621 (N_5621,N_2639,N_3196);
nand U5622 (N_5622,N_2041,N_3875);
xnor U5623 (N_5623,N_3340,N_3027);
nor U5624 (N_5624,N_3727,N_2274);
nand U5625 (N_5625,N_3866,N_3814);
nor U5626 (N_5626,N_2754,N_3885);
and U5627 (N_5627,N_2298,N_2741);
and U5628 (N_5628,N_2592,N_3754);
nor U5629 (N_5629,N_3787,N_2109);
or U5630 (N_5630,N_3375,N_3131);
and U5631 (N_5631,N_2478,N_3287);
and U5632 (N_5632,N_2777,N_3828);
or U5633 (N_5633,N_3419,N_3103);
or U5634 (N_5634,N_2728,N_2938);
and U5635 (N_5635,N_3007,N_3255);
and U5636 (N_5636,N_2603,N_2518);
and U5637 (N_5637,N_3674,N_3143);
xnor U5638 (N_5638,N_3757,N_2815);
and U5639 (N_5639,N_2286,N_3131);
or U5640 (N_5640,N_2547,N_3707);
xor U5641 (N_5641,N_2036,N_2735);
nand U5642 (N_5642,N_2722,N_3953);
nor U5643 (N_5643,N_3337,N_3129);
or U5644 (N_5644,N_3797,N_2431);
nand U5645 (N_5645,N_3449,N_3918);
nand U5646 (N_5646,N_2975,N_2011);
nand U5647 (N_5647,N_3885,N_2745);
nand U5648 (N_5648,N_2338,N_3866);
or U5649 (N_5649,N_2380,N_3109);
nor U5650 (N_5650,N_2887,N_3750);
and U5651 (N_5651,N_3813,N_2675);
and U5652 (N_5652,N_2299,N_3183);
nor U5653 (N_5653,N_2355,N_3060);
nor U5654 (N_5654,N_3756,N_2724);
and U5655 (N_5655,N_3131,N_2938);
nor U5656 (N_5656,N_3849,N_3175);
or U5657 (N_5657,N_3817,N_2698);
or U5658 (N_5658,N_2661,N_2554);
and U5659 (N_5659,N_2656,N_3263);
nand U5660 (N_5660,N_2011,N_2330);
and U5661 (N_5661,N_3088,N_3235);
nand U5662 (N_5662,N_2868,N_3486);
nor U5663 (N_5663,N_3568,N_3433);
or U5664 (N_5664,N_2554,N_3496);
nor U5665 (N_5665,N_3871,N_3165);
and U5666 (N_5666,N_2692,N_3401);
or U5667 (N_5667,N_2175,N_2966);
and U5668 (N_5668,N_2112,N_2168);
or U5669 (N_5669,N_3988,N_3222);
and U5670 (N_5670,N_3411,N_3866);
and U5671 (N_5671,N_3888,N_2169);
nand U5672 (N_5672,N_3133,N_3818);
and U5673 (N_5673,N_2099,N_3372);
xor U5674 (N_5674,N_2067,N_3611);
and U5675 (N_5675,N_2444,N_2946);
nand U5676 (N_5676,N_2349,N_2475);
and U5677 (N_5677,N_2907,N_2119);
and U5678 (N_5678,N_3585,N_2869);
nor U5679 (N_5679,N_3014,N_3045);
nor U5680 (N_5680,N_3200,N_2684);
or U5681 (N_5681,N_2336,N_2741);
and U5682 (N_5682,N_3206,N_2177);
or U5683 (N_5683,N_2151,N_3063);
or U5684 (N_5684,N_3290,N_2940);
or U5685 (N_5685,N_2521,N_2219);
or U5686 (N_5686,N_3255,N_3345);
or U5687 (N_5687,N_2570,N_2380);
or U5688 (N_5688,N_3013,N_3415);
and U5689 (N_5689,N_3216,N_2952);
nand U5690 (N_5690,N_3863,N_3237);
and U5691 (N_5691,N_3582,N_2088);
or U5692 (N_5692,N_3376,N_3864);
nand U5693 (N_5693,N_2113,N_3562);
and U5694 (N_5694,N_3302,N_2859);
and U5695 (N_5695,N_2716,N_3688);
nor U5696 (N_5696,N_3728,N_3337);
nand U5697 (N_5697,N_2838,N_2173);
or U5698 (N_5698,N_2041,N_2431);
nor U5699 (N_5699,N_3407,N_3806);
or U5700 (N_5700,N_2815,N_3527);
nor U5701 (N_5701,N_3462,N_2303);
xnor U5702 (N_5702,N_3101,N_2341);
and U5703 (N_5703,N_3622,N_2833);
nand U5704 (N_5704,N_3185,N_2118);
and U5705 (N_5705,N_2666,N_2896);
nor U5706 (N_5706,N_3120,N_3221);
xor U5707 (N_5707,N_2296,N_2531);
or U5708 (N_5708,N_3363,N_2362);
nand U5709 (N_5709,N_3830,N_3203);
nand U5710 (N_5710,N_2765,N_3584);
or U5711 (N_5711,N_2020,N_2599);
nor U5712 (N_5712,N_2458,N_3385);
nor U5713 (N_5713,N_2726,N_2315);
or U5714 (N_5714,N_2478,N_3605);
or U5715 (N_5715,N_2635,N_3670);
nor U5716 (N_5716,N_3870,N_2349);
and U5717 (N_5717,N_2695,N_3771);
nand U5718 (N_5718,N_2351,N_2100);
and U5719 (N_5719,N_3490,N_3300);
or U5720 (N_5720,N_2446,N_3959);
nand U5721 (N_5721,N_3727,N_3407);
or U5722 (N_5722,N_3893,N_3171);
nand U5723 (N_5723,N_2195,N_3919);
xnor U5724 (N_5724,N_2387,N_2694);
and U5725 (N_5725,N_3439,N_2126);
nor U5726 (N_5726,N_2713,N_3304);
nand U5727 (N_5727,N_3815,N_2235);
nor U5728 (N_5728,N_2942,N_3404);
nand U5729 (N_5729,N_3452,N_3307);
or U5730 (N_5730,N_2743,N_2887);
nand U5731 (N_5731,N_3714,N_3285);
and U5732 (N_5732,N_3129,N_2711);
nand U5733 (N_5733,N_3862,N_3982);
nor U5734 (N_5734,N_2507,N_3310);
nand U5735 (N_5735,N_3953,N_2180);
or U5736 (N_5736,N_3429,N_2935);
and U5737 (N_5737,N_3249,N_2052);
nor U5738 (N_5738,N_3454,N_2748);
nand U5739 (N_5739,N_2602,N_2163);
or U5740 (N_5740,N_3946,N_2991);
nand U5741 (N_5741,N_3798,N_2901);
and U5742 (N_5742,N_3609,N_2307);
nor U5743 (N_5743,N_3688,N_3261);
and U5744 (N_5744,N_2814,N_2820);
and U5745 (N_5745,N_2192,N_3300);
xnor U5746 (N_5746,N_2639,N_2484);
nand U5747 (N_5747,N_3189,N_2566);
and U5748 (N_5748,N_3380,N_2735);
nor U5749 (N_5749,N_2350,N_3203);
nand U5750 (N_5750,N_3268,N_2336);
nand U5751 (N_5751,N_2218,N_2574);
or U5752 (N_5752,N_3430,N_3054);
nand U5753 (N_5753,N_3982,N_2594);
or U5754 (N_5754,N_3942,N_3320);
nor U5755 (N_5755,N_3125,N_2501);
xnor U5756 (N_5756,N_3809,N_2834);
nor U5757 (N_5757,N_3062,N_2639);
and U5758 (N_5758,N_2444,N_2810);
nor U5759 (N_5759,N_2165,N_3366);
nor U5760 (N_5760,N_2287,N_2727);
nor U5761 (N_5761,N_2357,N_2326);
nor U5762 (N_5762,N_2745,N_3855);
xnor U5763 (N_5763,N_3360,N_3284);
nor U5764 (N_5764,N_2287,N_3775);
nand U5765 (N_5765,N_3837,N_3947);
nor U5766 (N_5766,N_2779,N_2540);
and U5767 (N_5767,N_3049,N_2088);
nor U5768 (N_5768,N_2743,N_2121);
or U5769 (N_5769,N_3873,N_2065);
nand U5770 (N_5770,N_2759,N_2023);
and U5771 (N_5771,N_3963,N_3000);
and U5772 (N_5772,N_3343,N_3255);
nor U5773 (N_5773,N_3994,N_3173);
and U5774 (N_5774,N_3854,N_3813);
or U5775 (N_5775,N_2782,N_2031);
and U5776 (N_5776,N_2501,N_2999);
nor U5777 (N_5777,N_3053,N_2610);
nand U5778 (N_5778,N_3163,N_2719);
nor U5779 (N_5779,N_2063,N_3204);
and U5780 (N_5780,N_3843,N_3504);
or U5781 (N_5781,N_3279,N_3028);
nand U5782 (N_5782,N_2550,N_3174);
or U5783 (N_5783,N_3829,N_2126);
nand U5784 (N_5784,N_2871,N_2651);
nor U5785 (N_5785,N_2730,N_3573);
or U5786 (N_5786,N_3519,N_2720);
nor U5787 (N_5787,N_2944,N_2109);
nand U5788 (N_5788,N_3754,N_2459);
or U5789 (N_5789,N_2218,N_3617);
or U5790 (N_5790,N_2580,N_3903);
nor U5791 (N_5791,N_3110,N_3003);
nor U5792 (N_5792,N_3492,N_3937);
xor U5793 (N_5793,N_2659,N_2175);
or U5794 (N_5794,N_2191,N_2719);
or U5795 (N_5795,N_2520,N_3507);
or U5796 (N_5796,N_3560,N_3876);
and U5797 (N_5797,N_2747,N_3070);
nand U5798 (N_5798,N_3854,N_3484);
nor U5799 (N_5799,N_2484,N_3910);
nand U5800 (N_5800,N_3292,N_2744);
nand U5801 (N_5801,N_3786,N_3738);
xor U5802 (N_5802,N_2860,N_2142);
nor U5803 (N_5803,N_3135,N_2935);
or U5804 (N_5804,N_3137,N_2855);
nor U5805 (N_5805,N_2936,N_2962);
nand U5806 (N_5806,N_3842,N_2353);
or U5807 (N_5807,N_2333,N_2974);
or U5808 (N_5808,N_2657,N_3645);
or U5809 (N_5809,N_3220,N_2905);
or U5810 (N_5810,N_2377,N_3383);
nor U5811 (N_5811,N_3539,N_2804);
nand U5812 (N_5812,N_2255,N_2768);
nor U5813 (N_5813,N_2983,N_2282);
or U5814 (N_5814,N_3298,N_2927);
or U5815 (N_5815,N_3834,N_2387);
and U5816 (N_5816,N_2308,N_2658);
nand U5817 (N_5817,N_2393,N_3038);
nor U5818 (N_5818,N_3977,N_2183);
nand U5819 (N_5819,N_3317,N_2663);
nand U5820 (N_5820,N_3227,N_2951);
nor U5821 (N_5821,N_3757,N_2108);
nor U5822 (N_5822,N_2231,N_3720);
and U5823 (N_5823,N_3617,N_2643);
and U5824 (N_5824,N_3576,N_2432);
and U5825 (N_5825,N_2221,N_2118);
and U5826 (N_5826,N_2612,N_2888);
nor U5827 (N_5827,N_2400,N_2972);
xnor U5828 (N_5828,N_2284,N_2100);
nor U5829 (N_5829,N_2921,N_3927);
nand U5830 (N_5830,N_2371,N_2247);
nand U5831 (N_5831,N_2273,N_3513);
and U5832 (N_5832,N_3586,N_2906);
or U5833 (N_5833,N_2611,N_2311);
nor U5834 (N_5834,N_2740,N_2384);
nor U5835 (N_5835,N_2218,N_3531);
or U5836 (N_5836,N_3430,N_3612);
nor U5837 (N_5837,N_3778,N_3271);
and U5838 (N_5838,N_2360,N_2657);
or U5839 (N_5839,N_3771,N_3346);
nor U5840 (N_5840,N_2735,N_2864);
nor U5841 (N_5841,N_3484,N_2805);
and U5842 (N_5842,N_2402,N_3929);
nand U5843 (N_5843,N_3188,N_3505);
nor U5844 (N_5844,N_2163,N_2936);
nor U5845 (N_5845,N_3657,N_3238);
nor U5846 (N_5846,N_2938,N_3189);
or U5847 (N_5847,N_2850,N_3326);
or U5848 (N_5848,N_2382,N_2148);
or U5849 (N_5849,N_3354,N_2133);
nor U5850 (N_5850,N_3772,N_2842);
nor U5851 (N_5851,N_3172,N_3588);
nor U5852 (N_5852,N_2125,N_3651);
and U5853 (N_5853,N_2712,N_2969);
or U5854 (N_5854,N_2111,N_3765);
or U5855 (N_5855,N_3722,N_2877);
or U5856 (N_5856,N_3592,N_3683);
or U5857 (N_5857,N_2964,N_2956);
nor U5858 (N_5858,N_2966,N_2228);
and U5859 (N_5859,N_2090,N_2369);
or U5860 (N_5860,N_2390,N_2618);
nor U5861 (N_5861,N_2215,N_2232);
nor U5862 (N_5862,N_2904,N_2034);
nand U5863 (N_5863,N_2966,N_3987);
or U5864 (N_5864,N_2609,N_3527);
or U5865 (N_5865,N_2189,N_2185);
or U5866 (N_5866,N_2075,N_2611);
nor U5867 (N_5867,N_3612,N_3812);
or U5868 (N_5868,N_3780,N_2719);
nand U5869 (N_5869,N_2467,N_2047);
xnor U5870 (N_5870,N_2934,N_3883);
and U5871 (N_5871,N_2316,N_3948);
or U5872 (N_5872,N_3005,N_2631);
nor U5873 (N_5873,N_2514,N_3894);
nor U5874 (N_5874,N_3104,N_2209);
and U5875 (N_5875,N_2766,N_2572);
or U5876 (N_5876,N_2246,N_3358);
nand U5877 (N_5877,N_2254,N_2145);
nor U5878 (N_5878,N_3527,N_3173);
nor U5879 (N_5879,N_3850,N_2843);
and U5880 (N_5880,N_3050,N_3877);
nand U5881 (N_5881,N_2051,N_2576);
nor U5882 (N_5882,N_2681,N_3076);
or U5883 (N_5883,N_2524,N_2303);
or U5884 (N_5884,N_2686,N_2382);
and U5885 (N_5885,N_3770,N_3864);
nand U5886 (N_5886,N_2657,N_2115);
nand U5887 (N_5887,N_2239,N_2860);
or U5888 (N_5888,N_3986,N_2439);
xor U5889 (N_5889,N_3411,N_3828);
nand U5890 (N_5890,N_3201,N_3880);
nand U5891 (N_5891,N_2949,N_3149);
nand U5892 (N_5892,N_2867,N_2868);
nand U5893 (N_5893,N_3792,N_2847);
nand U5894 (N_5894,N_2638,N_2651);
nor U5895 (N_5895,N_3896,N_2250);
or U5896 (N_5896,N_2373,N_3046);
or U5897 (N_5897,N_2440,N_2223);
nor U5898 (N_5898,N_2127,N_3635);
nand U5899 (N_5899,N_3615,N_3531);
and U5900 (N_5900,N_3553,N_2345);
or U5901 (N_5901,N_3205,N_3998);
nor U5902 (N_5902,N_3621,N_3903);
xnor U5903 (N_5903,N_3779,N_3517);
xnor U5904 (N_5904,N_3376,N_2623);
nor U5905 (N_5905,N_2982,N_2393);
and U5906 (N_5906,N_3829,N_2651);
and U5907 (N_5907,N_3854,N_2054);
nor U5908 (N_5908,N_3594,N_2212);
nand U5909 (N_5909,N_2491,N_3467);
nor U5910 (N_5910,N_2796,N_2379);
or U5911 (N_5911,N_3215,N_2996);
nor U5912 (N_5912,N_3207,N_2131);
nor U5913 (N_5913,N_2618,N_3875);
nor U5914 (N_5914,N_2000,N_2080);
nand U5915 (N_5915,N_2445,N_2002);
nand U5916 (N_5916,N_3684,N_2815);
or U5917 (N_5917,N_2604,N_3092);
or U5918 (N_5918,N_3932,N_3458);
or U5919 (N_5919,N_2848,N_2775);
nand U5920 (N_5920,N_2028,N_2167);
and U5921 (N_5921,N_2335,N_3961);
or U5922 (N_5922,N_3731,N_3297);
or U5923 (N_5923,N_3566,N_2049);
and U5924 (N_5924,N_2994,N_2859);
nor U5925 (N_5925,N_2927,N_2401);
or U5926 (N_5926,N_2137,N_2573);
nor U5927 (N_5927,N_2045,N_3425);
nand U5928 (N_5928,N_2164,N_3258);
nand U5929 (N_5929,N_3462,N_3046);
nand U5930 (N_5930,N_3449,N_3489);
nor U5931 (N_5931,N_3365,N_2937);
nor U5932 (N_5932,N_3384,N_2947);
nand U5933 (N_5933,N_2419,N_3291);
nand U5934 (N_5934,N_2356,N_2389);
nor U5935 (N_5935,N_3285,N_2567);
nor U5936 (N_5936,N_2007,N_2822);
xor U5937 (N_5937,N_3275,N_2073);
nor U5938 (N_5938,N_2702,N_3467);
nor U5939 (N_5939,N_3105,N_3635);
or U5940 (N_5940,N_3442,N_2043);
and U5941 (N_5941,N_2638,N_2141);
nor U5942 (N_5942,N_3242,N_3593);
and U5943 (N_5943,N_2394,N_2683);
or U5944 (N_5944,N_3793,N_2748);
nor U5945 (N_5945,N_3220,N_3752);
nand U5946 (N_5946,N_2113,N_3745);
or U5947 (N_5947,N_3969,N_2025);
or U5948 (N_5948,N_3289,N_3520);
nor U5949 (N_5949,N_2701,N_2763);
or U5950 (N_5950,N_2744,N_3752);
or U5951 (N_5951,N_2677,N_3852);
nand U5952 (N_5952,N_3516,N_3005);
xnor U5953 (N_5953,N_2353,N_2017);
nor U5954 (N_5954,N_3201,N_2317);
nand U5955 (N_5955,N_2443,N_3594);
or U5956 (N_5956,N_3804,N_2278);
nor U5957 (N_5957,N_3705,N_3474);
nand U5958 (N_5958,N_2148,N_2748);
and U5959 (N_5959,N_2602,N_2070);
or U5960 (N_5960,N_3045,N_3154);
and U5961 (N_5961,N_3967,N_3321);
nor U5962 (N_5962,N_2908,N_3558);
and U5963 (N_5963,N_3396,N_2743);
and U5964 (N_5964,N_3401,N_3571);
or U5965 (N_5965,N_2290,N_3441);
nor U5966 (N_5966,N_2269,N_2590);
and U5967 (N_5967,N_3973,N_2004);
nor U5968 (N_5968,N_2328,N_2220);
nor U5969 (N_5969,N_2129,N_2019);
nand U5970 (N_5970,N_3617,N_3745);
nand U5971 (N_5971,N_3590,N_3455);
or U5972 (N_5972,N_3252,N_2320);
or U5973 (N_5973,N_3910,N_2732);
nand U5974 (N_5974,N_2169,N_2474);
nor U5975 (N_5975,N_3920,N_3906);
nand U5976 (N_5976,N_3547,N_3381);
nor U5977 (N_5977,N_3338,N_3668);
or U5978 (N_5978,N_2958,N_3909);
and U5979 (N_5979,N_2134,N_2837);
or U5980 (N_5980,N_2513,N_2810);
nor U5981 (N_5981,N_2491,N_2901);
nor U5982 (N_5982,N_3525,N_3740);
nand U5983 (N_5983,N_3684,N_2347);
nor U5984 (N_5984,N_3232,N_3986);
or U5985 (N_5985,N_3583,N_3258);
or U5986 (N_5986,N_2314,N_2128);
nor U5987 (N_5987,N_2792,N_3824);
and U5988 (N_5988,N_2609,N_2691);
nand U5989 (N_5989,N_3087,N_3170);
or U5990 (N_5990,N_3645,N_2231);
and U5991 (N_5991,N_2168,N_3988);
nor U5992 (N_5992,N_2341,N_3366);
nor U5993 (N_5993,N_3471,N_2995);
and U5994 (N_5994,N_3721,N_2397);
xor U5995 (N_5995,N_2048,N_2578);
and U5996 (N_5996,N_3557,N_3181);
or U5997 (N_5997,N_3052,N_3668);
nand U5998 (N_5998,N_3850,N_2361);
or U5999 (N_5999,N_2111,N_2937);
nand U6000 (N_6000,N_5602,N_5225);
or U6001 (N_6001,N_5134,N_4777);
and U6002 (N_6002,N_4882,N_4952);
or U6003 (N_6003,N_4159,N_4119);
or U6004 (N_6004,N_5715,N_5125);
or U6005 (N_6005,N_5524,N_4359);
nor U6006 (N_6006,N_4708,N_5728);
nor U6007 (N_6007,N_4475,N_4205);
nand U6008 (N_6008,N_4805,N_5086);
nand U6009 (N_6009,N_4265,N_5238);
and U6010 (N_6010,N_5351,N_5488);
nor U6011 (N_6011,N_4567,N_4076);
nor U6012 (N_6012,N_5635,N_4393);
and U6013 (N_6013,N_5271,N_5423);
nor U6014 (N_6014,N_5142,N_5419);
nor U6015 (N_6015,N_5667,N_5081);
and U6016 (N_6016,N_4761,N_4150);
and U6017 (N_6017,N_4658,N_4572);
or U6018 (N_6018,N_5124,N_5992);
nor U6019 (N_6019,N_5076,N_5658);
and U6020 (N_6020,N_5820,N_5362);
nand U6021 (N_6021,N_5607,N_4970);
nand U6022 (N_6022,N_4257,N_4997);
nand U6023 (N_6023,N_5983,N_5449);
nor U6024 (N_6024,N_5815,N_4547);
and U6025 (N_6025,N_5630,N_5769);
or U6026 (N_6026,N_4017,N_4370);
and U6027 (N_6027,N_4538,N_4378);
nand U6028 (N_6028,N_4812,N_4142);
nor U6029 (N_6029,N_5850,N_5755);
nor U6030 (N_6030,N_4508,N_5916);
nor U6031 (N_6031,N_4587,N_4958);
nor U6032 (N_6032,N_5822,N_4908);
and U6033 (N_6033,N_4451,N_5382);
nand U6034 (N_6034,N_5054,N_5513);
or U6035 (N_6035,N_5539,N_5463);
nor U6036 (N_6036,N_5313,N_5447);
and U6037 (N_6037,N_5892,N_5115);
xnor U6038 (N_6038,N_5029,N_5442);
or U6039 (N_6039,N_5034,N_5026);
or U6040 (N_6040,N_4801,N_5915);
or U6041 (N_6041,N_5632,N_5089);
or U6042 (N_6042,N_5101,N_5179);
and U6043 (N_6043,N_4629,N_5523);
nor U6044 (N_6044,N_4395,N_5138);
nor U6045 (N_6045,N_5944,N_4480);
or U6046 (N_6046,N_4627,N_5074);
and U6047 (N_6047,N_4756,N_5876);
and U6048 (N_6048,N_4273,N_5923);
xor U6049 (N_6049,N_5230,N_4774);
or U6050 (N_6050,N_5192,N_5098);
and U6051 (N_6051,N_5891,N_5512);
nor U6052 (N_6052,N_4862,N_5814);
and U6053 (N_6053,N_4876,N_5527);
and U6054 (N_6054,N_4576,N_5147);
nand U6055 (N_6055,N_5218,N_4710);
and U6056 (N_6056,N_5614,N_5304);
and U6057 (N_6057,N_4900,N_4580);
and U6058 (N_6058,N_4157,N_5993);
nand U6059 (N_6059,N_4069,N_4137);
and U6060 (N_6060,N_5253,N_5032);
nor U6061 (N_6061,N_4481,N_5693);
or U6062 (N_6062,N_4975,N_5918);
nor U6063 (N_6063,N_5795,N_5590);
or U6064 (N_6064,N_5484,N_4248);
or U6065 (N_6065,N_5152,N_4221);
or U6066 (N_6066,N_5331,N_4051);
and U6067 (N_6067,N_5399,N_4376);
nand U6068 (N_6068,N_4985,N_5033);
or U6069 (N_6069,N_5652,N_5121);
and U6070 (N_6070,N_4637,N_5063);
or U6071 (N_6071,N_5057,N_5754);
or U6072 (N_6072,N_5178,N_5831);
nand U6073 (N_6073,N_4957,N_5546);
and U6074 (N_6074,N_5500,N_4793);
xor U6075 (N_6075,N_4063,N_4836);
and U6076 (N_6076,N_5520,N_4660);
nand U6077 (N_6077,N_4094,N_4235);
nand U6078 (N_6078,N_5256,N_5269);
nand U6079 (N_6079,N_4798,N_5196);
or U6080 (N_6080,N_5401,N_5429);
or U6081 (N_6081,N_4476,N_5112);
nand U6082 (N_6082,N_4187,N_4670);
and U6083 (N_6083,N_4531,N_4542);
xor U6084 (N_6084,N_5722,N_5565);
nor U6085 (N_6085,N_5438,N_5244);
nand U6086 (N_6086,N_5422,N_4494);
and U6087 (N_6087,N_5837,N_4281);
or U6088 (N_6088,N_4607,N_5702);
or U6089 (N_6089,N_4739,N_4690);
and U6090 (N_6090,N_5002,N_4417);
nand U6091 (N_6091,N_5100,N_5267);
and U6092 (N_6092,N_4737,N_4227);
and U6093 (N_6093,N_5928,N_4114);
xor U6094 (N_6094,N_5289,N_4408);
and U6095 (N_6095,N_4244,N_5069);
nor U6096 (N_6096,N_4707,N_4055);
or U6097 (N_6097,N_4672,N_5986);
and U6098 (N_6098,N_4180,N_5622);
nor U6099 (N_6099,N_5644,N_5185);
nand U6100 (N_6100,N_4079,N_5227);
nand U6101 (N_6101,N_5593,N_5249);
nand U6102 (N_6102,N_5670,N_5566);
nor U6103 (N_6103,N_5296,N_4288);
and U6104 (N_6104,N_5330,N_5472);
and U6105 (N_6105,N_5941,N_5353);
nor U6106 (N_6106,N_4401,N_5301);
nand U6107 (N_6107,N_5273,N_5221);
or U6108 (N_6108,N_4655,N_5369);
or U6109 (N_6109,N_4458,N_5131);
or U6110 (N_6110,N_4215,N_5490);
and U6111 (N_6111,N_5260,N_4038);
nand U6112 (N_6112,N_5970,N_4392);
nand U6113 (N_6113,N_4694,N_4047);
nor U6114 (N_6114,N_5215,N_4930);
and U6115 (N_6115,N_5344,N_5777);
nand U6116 (N_6116,N_5698,N_4861);
and U6117 (N_6117,N_5174,N_5028);
nand U6118 (N_6118,N_4977,N_5339);
and U6119 (N_6119,N_5586,N_4746);
and U6120 (N_6120,N_5001,N_5551);
xor U6121 (N_6121,N_5024,N_5507);
and U6122 (N_6122,N_4754,N_5428);
and U6123 (N_6123,N_4034,N_4695);
nand U6124 (N_6124,N_5794,N_4551);
and U6125 (N_6125,N_4610,N_5924);
nand U6126 (N_6126,N_4742,N_5333);
or U6127 (N_6127,N_5917,N_5396);
nor U6128 (N_6128,N_5276,N_5655);
nor U6129 (N_6129,N_4251,N_4799);
and U6130 (N_6130,N_4546,N_5875);
nor U6131 (N_6131,N_5035,N_5025);
nor U6132 (N_6132,N_4220,N_5467);
nor U6133 (N_6133,N_5038,N_5342);
or U6134 (N_6134,N_5424,N_5716);
xnor U6135 (N_6135,N_4693,N_4686);
nor U6136 (N_6136,N_5621,N_5688);
or U6137 (N_6137,N_4816,N_4771);
nand U6138 (N_6138,N_5293,N_4425);
and U6139 (N_6139,N_5390,N_4571);
nand U6140 (N_6140,N_5842,N_4125);
nand U6141 (N_6141,N_4699,N_5020);
nand U6142 (N_6142,N_4734,N_4825);
or U6143 (N_6143,N_5677,N_4716);
and U6144 (N_6144,N_4441,N_4222);
nand U6145 (N_6145,N_5995,N_5625);
nand U6146 (N_6146,N_5361,N_5768);
nor U6147 (N_6147,N_4712,N_5400);
and U6148 (N_6148,N_5184,N_4644);
nor U6149 (N_6149,N_5937,N_4782);
nand U6150 (N_6150,N_4361,N_5783);
nand U6151 (N_6151,N_4999,N_4826);
nand U6152 (N_6152,N_4618,N_5407);
and U6153 (N_6153,N_4258,N_4520);
nand U6154 (N_6154,N_4138,N_4267);
nand U6155 (N_6155,N_5735,N_5654);
nor U6156 (N_6156,N_5833,N_4880);
and U6157 (N_6157,N_4250,N_4489);
nor U6158 (N_6158,N_5170,N_4131);
and U6159 (N_6159,N_4337,N_5933);
or U6160 (N_6160,N_5056,N_4843);
and U6161 (N_6161,N_5136,N_4200);
nor U6162 (N_6162,N_4926,N_5936);
or U6163 (N_6163,N_5263,N_4657);
nor U6164 (N_6164,N_4133,N_5019);
or U6165 (N_6165,N_4402,N_5542);
and U6166 (N_6166,N_5562,N_5886);
or U6167 (N_6167,N_4462,N_5480);
nand U6168 (N_6168,N_4356,N_4307);
nand U6169 (N_6169,N_4024,N_4647);
nand U6170 (N_6170,N_4340,N_4355);
nor U6171 (N_6171,N_4072,N_4078);
or U6172 (N_6172,N_4797,N_4332);
nor U6173 (N_6173,N_5307,N_5888);
or U6174 (N_6174,N_5058,N_4788);
or U6175 (N_6175,N_4562,N_4866);
or U6176 (N_6176,N_4775,N_4169);
nor U6177 (N_6177,N_4113,N_4285);
or U6178 (N_6178,N_4140,N_4469);
or U6179 (N_6179,N_4488,N_5869);
nand U6180 (N_6180,N_4852,N_5912);
and U6181 (N_6181,N_4559,N_4988);
nand U6182 (N_6182,N_5234,N_5990);
nand U6183 (N_6183,N_4101,N_5648);
or U6184 (N_6184,N_5650,N_4949);
nor U6185 (N_6185,N_5753,N_4887);
and U6186 (N_6186,N_4535,N_5270);
and U6187 (N_6187,N_5280,N_4236);
nand U6188 (N_6188,N_4075,N_4297);
nor U6189 (N_6189,N_4346,N_4490);
nor U6190 (N_6190,N_4036,N_5398);
nor U6191 (N_6191,N_5219,N_4884);
or U6192 (N_6192,N_4396,N_4192);
or U6193 (N_6193,N_4706,N_4185);
and U6194 (N_6194,N_5859,N_5096);
nor U6195 (N_6195,N_5976,N_5211);
nand U6196 (N_6196,N_4158,N_4147);
and U6197 (N_6197,N_5914,N_4642);
nand U6198 (N_6198,N_5105,N_4023);
nor U6199 (N_6199,N_4060,N_5853);
and U6200 (N_6200,N_4696,N_4522);
nand U6201 (N_6201,N_4615,N_4280);
nor U6202 (N_6202,N_5931,N_4633);
nand U6203 (N_6203,N_5092,N_5816);
nand U6204 (N_6204,N_4173,N_5727);
and U6205 (N_6205,N_4681,N_5909);
or U6206 (N_6206,N_5363,N_5903);
or U6207 (N_6207,N_4374,N_4423);
or U6208 (N_6208,N_4683,N_4011);
and U6209 (N_6209,N_5459,N_4726);
nor U6210 (N_6210,N_4904,N_4440);
nand U6211 (N_6211,N_5750,N_5160);
nand U6212 (N_6212,N_4599,N_5247);
nor U6213 (N_6213,N_4065,N_5127);
nor U6214 (N_6214,N_5445,N_4473);
or U6215 (N_6215,N_4561,N_5511);
nand U6216 (N_6216,N_5987,N_5656);
or U6217 (N_6217,N_4500,N_4713);
nand U6218 (N_6218,N_4093,N_5380);
and U6219 (N_6219,N_5981,N_5515);
nand U6220 (N_6220,N_4776,N_4045);
nor U6221 (N_6221,N_4584,N_4783);
and U6222 (N_6222,N_5505,N_4299);
nor U6223 (N_6223,N_4962,N_5871);
and U6224 (N_6224,N_4936,N_5682);
nor U6225 (N_6225,N_5763,N_5714);
nor U6226 (N_6226,N_4565,N_5126);
or U6227 (N_6227,N_4730,N_5486);
and U6228 (N_6228,N_4558,N_4006);
nand U6229 (N_6229,N_4426,N_4444);
and U6230 (N_6230,N_5953,N_5139);
nor U6231 (N_6231,N_5984,N_4089);
and U6232 (N_6232,N_5526,N_4806);
nand U6233 (N_6233,N_4953,N_5636);
and U6234 (N_6234,N_4564,N_5575);
or U6235 (N_6235,N_4669,N_4819);
nor U6236 (N_6236,N_4207,N_4530);
nand U6237 (N_6237,N_4759,N_5278);
or U6238 (N_6238,N_5141,N_5010);
and U6239 (N_6239,N_5379,N_4588);
or U6240 (N_6240,N_5952,N_5696);
nand U6241 (N_6241,N_4947,N_4027);
nand U6242 (N_6242,N_4301,N_4100);
or U6243 (N_6243,N_4684,N_4049);
nand U6244 (N_6244,N_5347,N_5994);
nand U6245 (N_6245,N_5319,N_5724);
or U6246 (N_6246,N_4829,N_4243);
nor U6247 (N_6247,N_4780,N_4501);
nor U6248 (N_6248,N_4868,N_5355);
and U6249 (N_6249,N_4019,N_4303);
and U6250 (N_6250,N_5675,N_4973);
and U6251 (N_6251,N_4925,N_5907);
nor U6252 (N_6252,N_4808,N_4581);
and U6253 (N_6253,N_4550,N_5574);
nor U6254 (N_6254,N_4966,N_4569);
and U6255 (N_6255,N_4008,N_5600);
nor U6256 (N_6256,N_4362,N_4418);
nand U6257 (N_6257,N_4659,N_5229);
nor U6258 (N_6258,N_4189,N_4083);
nor U6259 (N_6259,N_4330,N_4357);
nor U6260 (N_6260,N_4311,N_4116);
nor U6261 (N_6261,N_4172,N_4096);
or U6262 (N_6262,N_5543,N_5545);
and U6263 (N_6263,N_4081,N_4711);
nor U6264 (N_6264,N_4278,N_4616);
nand U6265 (N_6265,N_4430,N_5773);
nor U6266 (N_6266,N_5199,N_5881);
nor U6267 (N_6267,N_5938,N_4056);
or U6268 (N_6268,N_5797,N_5491);
nor U6269 (N_6269,N_4653,N_5746);
nand U6270 (N_6270,N_4928,N_5767);
nor U6271 (N_6271,N_4933,N_5665);
and U6272 (N_6272,N_4478,N_4692);
or U6273 (N_6273,N_4283,N_4463);
nor U6274 (N_6274,N_5308,N_5796);
nand U6275 (N_6275,N_5083,N_4807);
and U6276 (N_6276,N_4913,N_5188);
or U6277 (N_6277,N_4604,N_4032);
and U6278 (N_6278,N_4135,N_5341);
nor U6279 (N_6279,N_5427,N_5821);
nand U6280 (N_6280,N_4468,N_5294);
nand U6281 (N_6281,N_4838,N_5712);
or U6282 (N_6282,N_4557,N_4948);
and U6283 (N_6283,N_5062,N_5373);
and U6284 (N_6284,N_5645,N_5177);
nor U6285 (N_6285,N_5169,N_4287);
or U6286 (N_6286,N_5452,N_4968);
nor U6287 (N_6287,N_5320,N_4025);
or U6288 (N_6288,N_5252,N_5504);
or U6289 (N_6289,N_5734,N_5246);
nand U6290 (N_6290,N_4573,N_5956);
nand U6291 (N_6291,N_5388,N_4934);
or U6292 (N_6292,N_4316,N_5298);
or U6293 (N_6293,N_4160,N_4390);
nand U6294 (N_6294,N_4245,N_4578);
nand U6295 (N_6295,N_4817,N_4020);
nand U6296 (N_6296,N_5884,N_5774);
and U6297 (N_6297,N_5921,N_5672);
nand U6298 (N_6298,N_5477,N_4967);
and U6299 (N_6299,N_5552,N_4087);
nor U6300 (N_6300,N_5167,N_4086);
nor U6301 (N_6301,N_5966,N_5826);
and U6302 (N_6302,N_4612,N_5759);
nand U6303 (N_6303,N_5860,N_5159);
and U6304 (N_6304,N_5947,N_4994);
nand U6305 (N_6305,N_4464,N_5037);
xor U6306 (N_6306,N_4136,N_4269);
and U6307 (N_6307,N_5535,N_5474);
nand U6308 (N_6308,N_4398,N_5902);
and U6309 (N_6309,N_4784,N_5782);
and U6310 (N_6310,N_4132,N_5779);
nor U6311 (N_6311,N_4859,N_4733);
and U6312 (N_6312,N_5288,N_5883);
nand U6313 (N_6313,N_4422,N_4354);
nor U6314 (N_6314,N_4146,N_5343);
and U6315 (N_6315,N_4661,N_4750);
xor U6316 (N_6316,N_4989,N_5402);
nor U6317 (N_6317,N_5806,N_4896);
nor U6318 (N_6318,N_4082,N_4529);
nand U6319 (N_6319,N_5528,N_4613);
and U6320 (N_6320,N_5999,N_5075);
and U6321 (N_6321,N_4645,N_4638);
and U6322 (N_6322,N_5664,N_4911);
or U6323 (N_6323,N_5581,N_4184);
and U6324 (N_6324,N_5241,N_5908);
nor U6325 (N_6325,N_4343,N_4595);
or U6326 (N_6326,N_4831,N_5786);
or U6327 (N_6327,N_5945,N_5691);
nand U6328 (N_6328,N_4912,N_4366);
nor U6329 (N_6329,N_4971,N_4104);
nor U6330 (N_6330,N_5157,N_4106);
nor U6331 (N_6331,N_5877,N_5070);
or U6332 (N_6332,N_5117,N_4103);
or U6333 (N_6333,N_5023,N_5619);
nand U6334 (N_6334,N_5760,N_4141);
and U6335 (N_6335,N_5317,N_4855);
xnor U6336 (N_6336,N_4731,N_4648);
or U6337 (N_6337,N_5482,N_4001);
or U6338 (N_6338,N_4667,N_5613);
or U6339 (N_6339,N_5149,N_5872);
nor U6340 (N_6340,N_5186,N_4495);
and U6341 (N_6341,N_4519,N_4850);
or U6342 (N_6342,N_5766,N_4993);
nand U6343 (N_6343,N_4446,N_5564);
or U6344 (N_6344,N_5102,N_5761);
or U6345 (N_6345,N_5485,N_5109);
and U6346 (N_6346,N_5110,N_4409);
or U6347 (N_6347,N_4149,N_5444);
nand U6348 (N_6348,N_4715,N_5748);
or U6349 (N_6349,N_5775,N_4677);
or U6350 (N_6350,N_5757,N_4407);
or U6351 (N_6351,N_4260,N_4460);
nand U6352 (N_6352,N_5687,N_5996);
and U6353 (N_6353,N_5228,N_4411);
nand U6354 (N_6354,N_5740,N_4676);
and U6355 (N_6355,N_4996,N_4099);
and U6356 (N_6356,N_4515,N_4620);
or U6357 (N_6357,N_5541,N_4840);
and U6358 (N_6358,N_5873,N_5948);
nand U6359 (N_6359,N_4981,N_5053);
nand U6360 (N_6360,N_4275,N_5018);
and U6361 (N_6361,N_5466,N_4810);
nor U6362 (N_6362,N_5749,N_5925);
xor U6363 (N_6363,N_5303,N_4511);
nor U6364 (N_6364,N_5509,N_4214);
xnor U6365 (N_6365,N_4323,N_4091);
nor U6366 (N_6366,N_4129,N_4188);
nand U6367 (N_6367,N_4767,N_4582);
and U6368 (N_6368,N_4641,N_4624);
or U6369 (N_6369,N_5222,N_4540);
or U6370 (N_6370,N_4689,N_4074);
and U6371 (N_6371,N_5164,N_5325);
or U6372 (N_6372,N_5408,N_5906);
or U6373 (N_6373,N_5591,N_5846);
nand U6374 (N_6374,N_5660,N_4537);
nor U6375 (N_6375,N_5878,N_5699);
or U6376 (N_6376,N_5437,N_4745);
nand U6377 (N_6377,N_5310,N_4014);
or U6378 (N_6378,N_4679,N_4791);
nor U6379 (N_6379,N_5071,N_4154);
and U6380 (N_6380,N_5412,N_5961);
nor U6381 (N_6381,N_5974,N_5108);
and U6382 (N_6382,N_4552,N_5627);
and U6383 (N_6383,N_5803,N_4510);
nand U6384 (N_6384,N_4371,N_4853);
or U6385 (N_6385,N_4987,N_4268);
nand U6386 (N_6386,N_5243,N_5455);
nor U6387 (N_6387,N_5231,N_5744);
nor U6388 (N_6388,N_5697,N_4955);
xor U6389 (N_6389,N_5604,N_4951);
or U6390 (N_6390,N_5060,N_5251);
nand U6391 (N_6391,N_5723,N_4084);
nor U6392 (N_6392,N_4212,N_5791);
nor U6393 (N_6393,N_5095,N_4143);
or U6394 (N_6394,N_5493,N_4654);
and U6395 (N_6395,N_4673,N_4111);
and U6396 (N_6396,N_5371,N_5559);
or U6397 (N_6397,N_5003,N_5977);
and U6398 (N_6398,N_5299,N_4863);
or U6399 (N_6399,N_5854,N_5762);
nor U6400 (N_6400,N_5348,N_5879);
and U6401 (N_6401,N_4961,N_4211);
or U6402 (N_6402,N_4972,N_5862);
nor U6403 (N_6403,N_4424,N_5140);
or U6404 (N_6404,N_5690,N_5680);
nand U6405 (N_6405,N_5262,N_4246);
nand U6406 (N_6406,N_4702,N_5726);
or U6407 (N_6407,N_5129,N_4964);
or U6408 (N_6408,N_4272,N_5181);
and U6409 (N_6409,N_4773,N_5066);
or U6410 (N_6410,N_5856,N_5237);
nand U6411 (N_6411,N_5316,N_4168);
and U6412 (N_6412,N_4899,N_5898);
nand U6413 (N_6413,N_4445,N_5730);
and U6414 (N_6414,N_4284,N_5957);
xor U6415 (N_6415,N_4929,N_4685);
nor U6416 (N_6416,N_4443,N_5823);
nor U6417 (N_6417,N_4874,N_4636);
xnor U6418 (N_6418,N_5106,N_5599);
and U6419 (N_6419,N_5819,N_5250);
and U6420 (N_6420,N_4623,N_4650);
nor U6421 (N_6421,N_4218,N_4066);
and U6422 (N_6422,N_4050,N_5700);
xor U6423 (N_6423,N_5224,N_4639);
or U6424 (N_6424,N_5649,N_5587);
nor U6425 (N_6425,N_4005,N_5703);
nand U6426 (N_6426,N_4318,N_4198);
nor U6427 (N_6427,N_4107,N_5537);
and U6428 (N_6428,N_5397,N_5261);
and U6429 (N_6429,N_4313,N_4544);
nor U6430 (N_6430,N_5805,N_4419);
nor U6431 (N_6431,N_4902,N_5804);
nand U6432 (N_6432,N_4940,N_4379);
or U6433 (N_6433,N_4643,N_4593);
nor U6434 (N_6434,N_4932,N_4845);
nor U6435 (N_6435,N_5557,N_4252);
nor U6436 (N_6436,N_4353,N_4886);
and U6437 (N_6437,N_5415,N_5616);
nor U6438 (N_6438,N_4282,N_4735);
xnor U6439 (N_6439,N_4437,N_4090);
and U6440 (N_6440,N_5501,N_5838);
or U6441 (N_6441,N_5352,N_5284);
nor U6442 (N_6442,N_4178,N_4484);
nand U6443 (N_6443,N_4487,N_4504);
and U6444 (N_6444,N_5571,N_4892);
or U6445 (N_6445,N_4007,N_5830);
nor U6446 (N_6446,N_5824,N_5052);
nand U6447 (N_6447,N_4814,N_5356);
nand U6448 (N_6448,N_4873,N_5579);
nor U6449 (N_6449,N_5084,N_5817);
nor U6450 (N_6450,N_5764,N_5306);
xor U6451 (N_6451,N_4170,N_4339);
and U6452 (N_6452,N_5836,N_5420);
or U6453 (N_6453,N_4059,N_4786);
nand U6454 (N_6454,N_5114,N_4021);
nand U6455 (N_6455,N_4291,N_5686);
nor U6456 (N_6456,N_4503,N_5738);
nand U6457 (N_6457,N_5404,N_4796);
and U6458 (N_6458,N_4848,N_5360);
or U6459 (N_6459,N_5416,N_5475);
or U6460 (N_6460,N_4858,N_5272);
nand U6461 (N_6461,N_4483,N_5922);
or U6462 (N_6462,N_4678,N_5671);
and U6463 (N_6463,N_4255,N_4450);
nor U6464 (N_6464,N_5171,N_5132);
nand U6465 (N_6465,N_5499,N_5737);
or U6466 (N_6466,N_4941,N_5643);
and U6467 (N_6467,N_5770,N_4319);
or U6468 (N_6468,N_4219,N_4950);
or U6469 (N_6469,N_5802,N_5409);
or U6470 (N_6470,N_4763,N_4867);
nor U6471 (N_6471,N_5030,N_4322);
nand U6472 (N_6472,N_5413,N_5538);
nor U6473 (N_6473,N_4037,N_5311);
and U6474 (N_6474,N_4671,N_4592);
and U6475 (N_6475,N_4556,N_4474);
or U6476 (N_6476,N_4338,N_4175);
and U6477 (N_6477,N_5865,N_5161);
nor U6478 (N_6478,N_5022,N_5573);
or U6479 (N_6479,N_4583,N_4839);
and U6480 (N_6480,N_5258,N_4331);
and U6481 (N_6481,N_4271,N_4864);
nor U6482 (N_6482,N_4691,N_4732);
and U6483 (N_6483,N_4415,N_5732);
or U6484 (N_6484,N_4109,N_5067);
and U6485 (N_6485,N_5971,N_5277);
or U6486 (N_6486,N_4760,N_5560);
nor U6487 (N_6487,N_5531,N_5784);
nand U6488 (N_6488,N_5930,N_5099);
nor U6489 (N_6489,N_5955,N_5741);
nor U6490 (N_6490,N_4598,N_5997);
nor U6491 (N_6491,N_4309,N_5495);
nor U6492 (N_6492,N_5618,N_5979);
xnor U6493 (N_6493,N_5041,N_5631);
nand U6494 (N_6494,N_4498,N_4959);
nor U6495 (N_6495,N_5213,N_4924);
and U6496 (N_6496,N_5265,N_4206);
nand U6497 (N_6497,N_5611,N_5895);
nand U6498 (N_6498,N_4609,N_4202);
and U6499 (N_6499,N_4071,N_4982);
and U6500 (N_6500,N_5612,N_4196);
nand U6501 (N_6501,N_4665,N_4491);
or U6502 (N_6502,N_5489,N_5812);
and U6503 (N_6503,N_5676,N_4765);
and U6504 (N_6504,N_4177,N_5935);
or U6505 (N_6505,N_4589,N_5701);
or U6506 (N_6506,N_5940,N_5122);
and U6507 (N_6507,N_5080,N_5745);
nand U6508 (N_6508,N_5006,N_4028);
nand U6509 (N_6509,N_4296,N_4115);
or U6510 (N_6510,N_5845,N_5346);
nor U6511 (N_6511,N_4879,N_5255);
or U6512 (N_6512,N_4105,N_4563);
and U6513 (N_6513,N_4431,N_4939);
nand U6514 (N_6514,N_5487,N_5297);
and U6515 (N_6515,N_5926,N_4747);
nand U6516 (N_6516,N_4375,N_5336);
nor U6517 (N_6517,N_4854,N_4470);
or U6518 (N_6518,N_5889,N_4523);
or U6519 (N_6519,N_5322,N_5692);
nand U6520 (N_6520,N_5350,N_5799);
nand U6521 (N_6521,N_4410,N_4216);
or U6522 (N_6522,N_5354,N_5532);
or U6523 (N_6523,N_4148,N_4594);
or U6524 (N_6524,N_4223,N_5608);
nand U6525 (N_6525,N_5291,N_4978);
or U6526 (N_6526,N_4822,N_4811);
and U6527 (N_6527,N_4719,N_5448);
xor U6528 (N_6528,N_4485,N_4514);
nand U6529 (N_6529,N_4605,N_5684);
and U6530 (N_6530,N_5329,N_5951);
and U6531 (N_6531,N_5998,N_4897);
and U6532 (N_6532,N_5282,N_4389);
and U6533 (N_6533,N_4603,N_4770);
nand U6534 (N_6534,N_4261,N_5248);
or U6535 (N_6535,N_5633,N_4888);
nor U6536 (N_6536,N_5440,N_5162);
nand U6537 (N_6537,N_5332,N_4012);
nand U6538 (N_6538,N_5426,N_5954);
or U6539 (N_6539,N_5040,N_5364);
and U6540 (N_6540,N_4516,N_5852);
nand U6541 (N_6541,N_4802,N_4058);
or U6542 (N_6542,N_4914,N_5318);
xor U6543 (N_6543,N_4203,N_4555);
or U6544 (N_6544,N_5666,N_4048);
nand U6545 (N_6545,N_5456,N_4197);
and U6546 (N_6546,N_4031,N_4035);
and U6547 (N_6547,N_5969,N_5357);
nand U6548 (N_6548,N_5148,N_4984);
nand U6549 (N_6549,N_5647,N_4352);
nor U6550 (N_6550,N_4429,N_4865);
nor U6551 (N_6551,N_4976,N_4813);
and U6552 (N_6552,N_4320,N_4404);
nand U6553 (N_6553,N_5207,N_4518);
or U6554 (N_6554,N_4327,N_4823);
or U6555 (N_6555,N_4764,N_4600);
nand U6556 (N_6556,N_5156,N_4310);
or U6557 (N_6557,N_4536,N_5778);
or U6558 (N_6558,N_4472,N_4640);
and U6559 (N_6559,N_4217,N_5610);
or U6560 (N_6560,N_5497,N_5481);
and U6561 (N_6561,N_4714,N_4092);
and U6562 (N_6562,N_4946,N_4314);
or U6563 (N_6563,N_5093,N_5494);
or U6564 (N_6564,N_4209,N_5868);
nand U6565 (N_6565,N_4664,N_5433);
and U6566 (N_6566,N_5240,N_4768);
and U6567 (N_6567,N_5042,N_5468);
and U6568 (N_6568,N_5626,N_5772);
or U6569 (N_6569,N_4698,N_4586);
or U6570 (N_6570,N_4980,N_5725);
nand U6571 (N_6571,N_5742,N_5536);
nor U6572 (N_6572,N_4351,N_5800);
nand U6573 (N_6573,N_4030,N_5385);
or U6574 (N_6574,N_4883,N_4723);
nor U6575 (N_6575,N_4386,N_4161);
nand U6576 (N_6576,N_4834,N_5638);
and U6577 (N_6577,N_4905,N_5717);
xnor U6578 (N_6578,N_4270,N_4724);
nand U6579 (N_6579,N_5751,N_5788);
nor U6580 (N_6580,N_4334,N_4266);
and U6581 (N_6581,N_4042,N_5939);
or U6582 (N_6582,N_4513,N_5340);
nand U6583 (N_6583,N_4875,N_5197);
nand U6584 (N_6584,N_4080,N_5965);
and U6585 (N_6585,N_5393,N_4675);
nor U6586 (N_6586,N_5606,N_5000);
or U6587 (N_6587,N_5887,N_5048);
and U6588 (N_6588,N_4729,N_4720);
and U6589 (N_6589,N_5128,N_5789);
nand U6590 (N_6590,N_4878,N_5103);
and U6591 (N_6591,N_5036,N_4242);
nor U6592 (N_6592,N_5568,N_4302);
nor U6593 (N_6593,N_4979,N_5988);
and U6594 (N_6594,N_5835,N_4800);
nand U6595 (N_6595,N_4348,N_4766);
or U6596 (N_6596,N_5810,N_4532);
nor U6597 (N_6597,N_5055,N_5785);
nand U6598 (N_6598,N_5300,N_4088);
nand U6599 (N_6599,N_4728,N_4794);
or U6600 (N_6600,N_5450,N_5464);
nand U6601 (N_6601,N_4341,N_4881);
nor U6602 (N_6602,N_4632,N_4434);
and U6603 (N_6603,N_5418,N_4043);
nor U6604 (N_6604,N_4960,N_4004);
nand U6605 (N_6605,N_4139,N_4380);
nand U6606 (N_6606,N_4891,N_5829);
and U6607 (N_6607,N_4439,N_4682);
or U6608 (N_6608,N_4917,N_5519);
and U6609 (N_6609,N_4986,N_5163);
nor U6610 (N_6610,N_5808,N_5479);
nor U6611 (N_6611,N_5894,N_4098);
or U6612 (N_6612,N_4492,N_5044);
nand U6613 (N_6613,N_4234,N_4804);
and U6614 (N_6614,N_4412,N_5257);
nor U6615 (N_6615,N_5719,N_5384);
or U6616 (N_6616,N_4145,N_4626);
and U6617 (N_6617,N_5629,N_4231);
nand U6618 (N_6618,N_4608,N_5432);
or U6619 (N_6619,N_5203,N_5597);
nand U6620 (N_6620,N_5292,N_5694);
or U6621 (N_6621,N_5135,N_5798);
xor U6622 (N_6622,N_4435,N_5217);
and U6623 (N_6623,N_5904,N_4877);
and U6624 (N_6624,N_4579,N_4772);
nor U6625 (N_6625,N_5882,N_5946);
or U6626 (N_6626,N_5386,N_5403);
and U6627 (N_6627,N_5890,N_5978);
nor U6628 (N_6628,N_5825,N_4898);
and U6629 (N_6629,N_5502,N_5790);
or U6630 (N_6630,N_5314,N_5743);
nand U6631 (N_6631,N_4000,N_5039);
or U6632 (N_6632,N_5078,N_4183);
and U6633 (N_6633,N_4945,N_4350);
nor U6634 (N_6634,N_5792,N_4363);
nor U6635 (N_6635,N_5378,N_4321);
and U6636 (N_6636,N_4787,N_4889);
nand U6637 (N_6637,N_5668,N_4022);
and U6638 (N_6638,N_5046,N_4029);
or U6639 (N_6639,N_4164,N_5787);
nor U6640 (N_6640,N_5483,N_4837);
and U6641 (N_6641,N_5462,N_5268);
or U6642 (N_6642,N_4403,N_5077);
or U6643 (N_6643,N_4449,N_5843);
nand U6644 (N_6644,N_4026,N_4053);
and U6645 (N_6645,N_4420,N_5620);
nor U6646 (N_6646,N_4009,N_4300);
and U6647 (N_6647,N_4457,N_5596);
nor U6648 (N_6648,N_4315,N_4870);
nor U6649 (N_6649,N_5577,N_5661);
nor U6650 (N_6650,N_4039,N_4117);
nand U6651 (N_6651,N_4406,N_4628);
nand U6652 (N_6652,N_4479,N_4545);
and U6653 (N_6653,N_4851,N_4385);
or U6654 (N_6654,N_5601,N_4849);
nand U6655 (N_6655,N_4630,N_5216);
and U6656 (N_6656,N_4174,N_4741);
or U6657 (N_6657,N_4688,N_4921);
or U6658 (N_6658,N_5473,N_4575);
nand U6659 (N_6659,N_5173,N_4381);
nor U6660 (N_6660,N_5841,N_5855);
nand U6661 (N_6661,N_4818,N_4128);
and U6662 (N_6662,N_4611,N_5045);
nor U6663 (N_6663,N_5189,N_4279);
nand U6664 (N_6664,N_5368,N_4828);
or U6665 (N_6665,N_5212,N_5123);
or U6666 (N_6666,N_5870,N_4130);
xnor U6667 (N_6667,N_5017,N_5043);
and U6668 (N_6668,N_4727,N_4305);
or U6669 (N_6669,N_4869,N_5375);
or U6670 (N_6670,N_5832,N_5430);
or U6671 (N_6671,N_4256,N_5534);
or U6672 (N_6672,N_5585,N_4068);
nand U6673 (N_6673,N_4349,N_5338);
and U6674 (N_6674,N_4195,N_4345);
or U6675 (N_6675,N_4910,N_5439);
nor U6676 (N_6676,N_4482,N_4163);
nor U6677 (N_6677,N_4992,N_4748);
nand U6678 (N_6678,N_4438,N_4162);
nand U6679 (N_6679,N_4738,N_5972);
nand U6680 (N_6680,N_5864,N_5107);
nand U6681 (N_6681,N_4121,N_5651);
nor U6682 (N_6682,N_5781,N_4326);
or U6683 (N_6683,N_5309,N_4602);
and U6684 (N_6684,N_4517,N_5370);
nor U6685 (N_6685,N_5465,N_4276);
nor U6686 (N_6686,N_4453,N_4596);
and U6687 (N_6687,N_4452,N_4264);
and U6688 (N_6688,N_4237,N_5049);
nor U6689 (N_6689,N_5540,N_4015);
and U6690 (N_6690,N_5175,N_4901);
or U6691 (N_6691,N_4991,N_5583);
or U6692 (N_6692,N_4938,N_4606);
and U6693 (N_6693,N_4466,N_5210);
and U6694 (N_6694,N_5013,N_4709);
or U6695 (N_6695,N_5793,N_5461);
nor U6696 (N_6696,N_5195,N_4725);
nand U6697 (N_6697,N_4856,N_4789);
nand U6698 (N_6698,N_5857,N_5009);
xor U6699 (N_6699,N_5434,N_5572);
or U6700 (N_6700,N_5960,N_4064);
nand U6701 (N_6701,N_5544,N_5756);
or U6702 (N_6702,N_4792,N_5266);
or U6703 (N_6703,N_5866,N_5150);
nand U6704 (N_6704,N_5594,N_4312);
and U6705 (N_6705,N_5707,N_4505);
nand U6706 (N_6706,N_5555,N_5014);
or U6707 (N_6707,N_4394,N_5365);
or U6708 (N_6708,N_4477,N_4033);
nand U6709 (N_6709,N_5451,N_4553);
and U6710 (N_6710,N_4920,N_4274);
nor U6711 (N_6711,N_4974,N_4666);
and U6712 (N_6712,N_5718,N_4803);
nor U6713 (N_6713,N_5153,N_4827);
or U6714 (N_6714,N_4965,N_5942);
and U6715 (N_6715,N_5595,N_5061);
xor U6716 (N_6716,N_4740,N_4333);
or U6717 (N_6717,N_4290,N_4182);
nand U6718 (N_6718,N_5359,N_5425);
nand U6719 (N_6719,N_4317,N_4903);
nand U6720 (N_6720,N_4367,N_5685);
nand U6721 (N_6721,N_5963,N_5695);
and U6722 (N_6722,N_4751,N_4368);
nand U6723 (N_6723,N_5962,N_4833);
or U6724 (N_6724,N_5807,N_5899);
nand U6725 (N_6725,N_4815,N_4204);
or U6726 (N_6726,N_5245,N_5897);
nand U6727 (N_6727,N_5047,N_5811);
and U6728 (N_6728,N_5120,N_4062);
nand U6729 (N_6729,N_4841,N_4414);
and U6730 (N_6730,N_4229,N_5506);
and U6731 (N_6731,N_5198,N_5839);
and U6732 (N_6732,N_4718,N_5050);
nor U6733 (N_6733,N_5844,N_5669);
nor U6734 (N_6734,N_4176,N_4663);
nand U6735 (N_6735,N_4541,N_5548);
nor U6736 (N_6736,N_5958,N_4943);
nor U6737 (N_6737,N_5068,N_5235);
xor U6738 (N_6738,N_4549,N_5705);
nor U6739 (N_6739,N_5905,N_5834);
and U6740 (N_6740,N_4289,N_5021);
and U6741 (N_6741,N_5980,N_5435);
nand U6742 (N_6742,N_4459,N_5421);
and U6743 (N_6743,N_5016,N_4365);
and U6744 (N_6744,N_4253,N_4832);
nand U6745 (N_6745,N_4687,N_5476);
or U6746 (N_6746,N_4895,N_5662);
and U6747 (N_6747,N_4342,N_5176);
and U6748 (N_6748,N_4526,N_4442);
nor U6749 (N_6749,N_5780,N_4230);
nand U6750 (N_6750,N_4554,N_5849);
nand U6751 (N_6751,N_4779,N_5964);
and U6752 (N_6752,N_5617,N_5335);
or U6753 (N_6753,N_4167,N_5283);
and U6754 (N_6754,N_4649,N_5950);
nor U6755 (N_6755,N_4016,N_5518);
nor U6756 (N_6756,N_5982,N_5460);
or U6757 (N_6757,N_5529,N_5337);
xor U6758 (N_6758,N_5137,N_4830);
and U6759 (N_6759,N_4755,N_4397);
nor U6760 (N_6760,N_4304,N_5927);
and U6761 (N_6761,N_5312,N_5733);
nand U6762 (N_6762,N_5508,N_4907);
nand U6763 (N_6763,N_5517,N_4166);
or U6764 (N_6764,N_4388,N_4743);
nor U6765 (N_6765,N_5328,N_4040);
nor U6766 (N_6766,N_5598,N_5469);
nor U6767 (N_6767,N_5327,N_5580);
or U6768 (N_6768,N_4634,N_5943);
and U6769 (N_6769,N_5315,N_4871);
nor U6770 (N_6770,N_5801,N_5326);
or U6771 (N_6771,N_4369,N_4155);
or U6772 (N_6772,N_5592,N_4447);
and U6773 (N_6773,N_4306,N_5729);
nand U6774 (N_6774,N_4954,N_5008);
nand U6775 (N_6775,N_5209,N_4860);
xor U6776 (N_6776,N_5183,N_5496);
nor U6777 (N_6777,N_5323,N_4585);
nor U6778 (N_6778,N_4239,N_4224);
nor U6779 (N_6779,N_5366,N_5254);
and U6780 (N_6780,N_5383,N_5279);
and U6781 (N_6781,N_5776,N_5901);
and U6782 (N_6782,N_5287,N_5007);
nor U6783 (N_6783,N_4110,N_4674);
or U6784 (N_6784,N_4118,N_4108);
and U6785 (N_6785,N_5233,N_5848);
nor U6786 (N_6786,N_4969,N_5094);
or U6787 (N_6787,N_5405,N_4232);
or U6788 (N_6788,N_4124,N_5031);
nor U6789 (N_6789,N_5985,N_4927);
and U6790 (N_6790,N_5454,N_4795);
and U6791 (N_6791,N_5200,N_4344);
nor U6792 (N_6792,N_5201,N_4456);
or U6793 (N_6793,N_4471,N_5012);
or U6794 (N_6794,N_5005,N_4433);
xnor U6795 (N_6795,N_5194,N_4697);
nand U6796 (N_6796,N_4120,N_4335);
or U6797 (N_6797,N_5713,N_4454);
or U6798 (N_6798,N_4590,N_5392);
nand U6799 (N_6799,N_4428,N_5569);
and U6800 (N_6800,N_4277,N_5588);
nand U6801 (N_6801,N_5959,N_5208);
or U6802 (N_6802,N_4186,N_5582);
nor U6803 (N_6803,N_4656,N_5919);
nor U6804 (N_6804,N_4543,N_5968);
or U6805 (N_6805,N_5880,N_5893);
and U6806 (N_6806,N_5158,N_5190);
nand U6807 (N_6807,N_5372,N_4286);
nand U6808 (N_6808,N_5453,N_4560);
nor U6809 (N_6809,N_4384,N_4391);
and U6810 (N_6810,N_5721,N_4790);
and U6811 (N_6811,N_4210,N_5867);
or U6812 (N_6812,N_5478,N_5949);
nand U6813 (N_6813,N_4651,N_5731);
or U6814 (N_6814,N_5295,N_4003);
or U6815 (N_6815,N_5736,N_4057);
nor U6816 (N_6816,N_5431,N_5530);
and U6817 (N_6817,N_4497,N_5498);
or U6818 (N_6818,N_5334,N_4347);
or U6819 (N_6819,N_5851,N_4915);
nor U6820 (N_6820,N_4528,N_4919);
nand U6821 (N_6821,N_5514,N_5097);
nor U6822 (N_6822,N_4413,N_4527);
or U6823 (N_6823,N_5165,N_4002);
and U6824 (N_6824,N_4512,N_4990);
nand U6825 (N_6825,N_4372,N_4680);
nand U6826 (N_6826,N_4533,N_4134);
and U6827 (N_6827,N_5683,N_4298);
nand U6828 (N_6828,N_5863,N_4191);
xor U6829 (N_6829,N_5264,N_5637);
or U6830 (N_6830,N_4360,N_4931);
and U6831 (N_6831,N_4700,N_4156);
nand U6832 (N_6832,N_5085,N_4018);
nor U6833 (N_6833,N_4601,N_4399);
nand U6834 (N_6834,N_5091,N_5133);
and U6835 (N_6835,N_5679,N_5417);
or U6836 (N_6836,N_5145,N_4364);
or U6837 (N_6837,N_4427,N_4171);
or U6838 (N_6838,N_4294,N_4292);
or U6839 (N_6839,N_4387,N_5065);
xor U6840 (N_6840,N_5510,N_5004);
and U6841 (N_6841,N_4382,N_5239);
or U6842 (N_6842,N_5706,N_4194);
nand U6843 (N_6843,N_5226,N_4077);
or U6844 (N_6844,N_4942,N_4944);
or U6845 (N_6845,N_4846,N_5547);
and U6846 (N_6846,N_4486,N_5166);
nand U6847 (N_6847,N_4885,N_5653);
or U6848 (N_6848,N_5642,N_5920);
nand U6849 (N_6849,N_5681,N_5710);
xor U6850 (N_6850,N_4112,N_5204);
and U6851 (N_6851,N_4521,N_4566);
nor U6852 (N_6852,N_5259,N_5274);
nand U6853 (N_6853,N_5242,N_4377);
nand U6854 (N_6854,N_5503,N_5151);
nand U6855 (N_6855,N_4179,N_5563);
or U6856 (N_6856,N_4752,N_5553);
and U6857 (N_6857,N_4835,N_4923);
nor U6858 (N_6858,N_4625,N_4646);
nor U6859 (N_6859,N_4293,N_5874);
nor U6860 (N_6860,N_5911,N_5395);
nor U6861 (N_6861,N_5064,N_5967);
and U6862 (N_6862,N_4844,N_4983);
and U6863 (N_6863,N_5674,N_5367);
and U6864 (N_6864,N_4506,N_4328);
and U6865 (N_6865,N_4568,N_4631);
nand U6866 (N_6866,N_4013,N_4054);
nand U6867 (N_6867,N_4785,N_5202);
nor U6868 (N_6868,N_5411,N_4956);
nand U6869 (N_6869,N_4916,N_4233);
or U6870 (N_6870,N_5991,N_5765);
nor U6871 (N_6871,N_4263,N_4507);
nor U6872 (N_6872,N_4652,N_5549);
nor U6873 (N_6873,N_5214,N_5578);
nor U6874 (N_6874,N_4703,N_5704);
and U6875 (N_6875,N_5191,N_5989);
and U6876 (N_6876,N_5657,N_5809);
nor U6877 (N_6877,N_5556,N_5286);
or U6878 (N_6878,N_5576,N_4574);
nor U6879 (N_6879,N_4421,N_4635);
and U6880 (N_6880,N_5522,N_5913);
or U6881 (N_6881,N_5236,N_4123);
and U6882 (N_6882,N_4295,N_4213);
and U6883 (N_6883,N_4102,N_5232);
or U6884 (N_6884,N_4405,N_5840);
nor U6885 (N_6885,N_4525,N_5059);
or U6886 (N_6886,N_5827,N_5206);
nor U6887 (N_6887,N_4165,N_5305);
nor U6888 (N_6888,N_5154,N_5090);
nand U6889 (N_6889,N_5758,N_5623);
nand U6890 (N_6890,N_4909,N_4201);
or U6891 (N_6891,N_4324,N_5861);
nor U6892 (N_6892,N_4127,N_5646);
or U6893 (N_6893,N_4151,N_4193);
nor U6894 (N_6894,N_5088,N_4662);
nor U6895 (N_6895,N_4509,N_4254);
or U6896 (N_6896,N_5441,N_5436);
and U6897 (N_6897,N_4722,N_5689);
nand U6898 (N_6898,N_5119,N_4614);
and U6899 (N_6899,N_5609,N_4668);
or U6900 (N_6900,N_5302,N_5752);
or U6901 (N_6901,N_4621,N_5847);
xor U6902 (N_6902,N_4241,N_4247);
nor U6903 (N_6903,N_4922,N_4570);
nor U6904 (N_6904,N_4208,N_5414);
and U6905 (N_6905,N_4238,N_5275);
nand U6906 (N_6906,N_5634,N_5446);
nor U6907 (N_6907,N_5910,N_4493);
or U6908 (N_6908,N_5321,N_5628);
nand U6909 (N_6909,N_5567,N_4085);
nor U6910 (N_6910,N_4757,N_5570);
nor U6911 (N_6911,N_4769,N_5376);
and U6912 (N_6912,N_5932,N_5709);
or U6913 (N_6913,N_5858,N_4998);
nor U6914 (N_6914,N_4190,N_4199);
and U6915 (N_6915,N_5155,N_5975);
or U6916 (N_6916,N_4890,N_4857);
and U6917 (N_6917,N_4432,N_4995);
or U6918 (N_6918,N_5443,N_5168);
nor U6919 (N_6919,N_5900,N_5104);
or U6920 (N_6920,N_4918,N_5471);
or U6921 (N_6921,N_5828,N_4144);
and U6922 (N_6922,N_5708,N_4534);
or U6923 (N_6923,N_5324,N_4847);
nor U6924 (N_6924,N_4383,N_5111);
or U6925 (N_6925,N_5558,N_5051);
or U6926 (N_6926,N_5406,N_4622);
and U6927 (N_6927,N_4373,N_5285);
and U6928 (N_6928,N_5673,N_5349);
or U6929 (N_6929,N_5144,N_4758);
and U6930 (N_6930,N_4436,N_4502);
nor U6931 (N_6931,N_5516,N_5603);
xor U6932 (N_6932,N_5470,N_4336);
or U6933 (N_6933,N_4052,N_4762);
or U6934 (N_6934,N_5896,N_5143);
nand U6935 (N_6935,N_5659,N_5525);
nand U6936 (N_6936,N_4749,N_5747);
or U6937 (N_6937,N_4893,N_4126);
nand U6938 (N_6938,N_4228,N_5584);
nor U6939 (N_6939,N_5187,N_5220);
nor U6940 (N_6940,N_4496,N_4577);
or U6941 (N_6941,N_5615,N_5130);
nand U6942 (N_6942,N_5389,N_5358);
or U6943 (N_6943,N_4781,N_5410);
nand U6944 (N_6944,N_4448,N_4704);
or U6945 (N_6945,N_5205,N_5027);
xor U6946 (N_6946,N_4937,N_5818);
nor U6947 (N_6947,N_4061,N_4591);
or U6948 (N_6948,N_5973,N_5739);
or U6949 (N_6949,N_5457,N_4465);
nor U6950 (N_6950,N_5641,N_4358);
nor U6951 (N_6951,N_4325,N_4963);
or U6952 (N_6952,N_4499,N_4809);
and U6953 (N_6953,N_4097,N_5281);
or U6954 (N_6954,N_5072,N_4240);
nand U6955 (N_6955,N_4524,N_5605);
nor U6956 (N_6956,N_4778,N_4539);
nand U6957 (N_6957,N_5387,N_5391);
nor U6958 (N_6958,N_4820,N_5290);
and U6959 (N_6959,N_4461,N_5118);
nor U6960 (N_6960,N_4935,N_4705);
nand U6961 (N_6961,N_5180,N_4872);
or U6962 (N_6962,N_4249,N_4821);
nand U6963 (N_6963,N_4073,N_5079);
nor U6964 (N_6964,N_5116,N_5533);
nor U6965 (N_6965,N_4226,N_4046);
nand U6966 (N_6966,N_4308,N_5015);
and U6967 (N_6967,N_5711,N_5663);
or U6968 (N_6968,N_4721,N_4894);
and U6969 (N_6969,N_4455,N_5172);
or U6970 (N_6970,N_4906,N_5550);
and U6971 (N_6971,N_5771,N_4467);
xnor U6972 (N_6972,N_5193,N_4153);
nand U6973 (N_6973,N_4701,N_5521);
nor U6974 (N_6974,N_4744,N_5087);
or U6975 (N_6975,N_5073,N_4095);
or U6976 (N_6976,N_5720,N_5934);
nand U6977 (N_6977,N_5589,N_5554);
and U6978 (N_6978,N_5374,N_4617);
nor U6979 (N_6979,N_5345,N_4753);
nor U6980 (N_6980,N_4152,N_4824);
or U6981 (N_6981,N_5929,N_4044);
nand U6982 (N_6982,N_5223,N_5492);
or U6983 (N_6983,N_5813,N_5394);
nand U6984 (N_6984,N_4181,N_4067);
nor U6985 (N_6985,N_4619,N_4070);
nor U6986 (N_6986,N_5624,N_4010);
nor U6987 (N_6987,N_5113,N_5082);
nor U6988 (N_6988,N_5011,N_5458);
nand U6989 (N_6989,N_4736,N_4122);
nand U6990 (N_6990,N_4717,N_4597);
nand U6991 (N_6991,N_4262,N_4225);
nor U6992 (N_6992,N_5639,N_4259);
nand U6993 (N_6993,N_5377,N_4329);
nor U6994 (N_6994,N_5678,N_4548);
and U6995 (N_6995,N_4842,N_4041);
nor U6996 (N_6996,N_5561,N_4400);
and U6997 (N_6997,N_4416,N_5182);
and U6998 (N_6998,N_5381,N_5146);
or U6999 (N_6999,N_5640,N_5885);
nor U7000 (N_7000,N_4711,N_5378);
and U7001 (N_7001,N_4819,N_5949);
or U7002 (N_7002,N_5333,N_4250);
and U7003 (N_7003,N_5743,N_5277);
or U7004 (N_7004,N_5328,N_4425);
nor U7005 (N_7005,N_5590,N_5353);
nor U7006 (N_7006,N_4921,N_5610);
or U7007 (N_7007,N_4886,N_5764);
and U7008 (N_7008,N_4097,N_4016);
or U7009 (N_7009,N_5794,N_5346);
nor U7010 (N_7010,N_4712,N_4626);
nand U7011 (N_7011,N_4243,N_4071);
or U7012 (N_7012,N_5719,N_5032);
nand U7013 (N_7013,N_5771,N_5093);
nor U7014 (N_7014,N_4425,N_4462);
nor U7015 (N_7015,N_4263,N_5209);
or U7016 (N_7016,N_5734,N_5355);
and U7017 (N_7017,N_5805,N_4238);
and U7018 (N_7018,N_4881,N_5585);
nor U7019 (N_7019,N_5275,N_5356);
nand U7020 (N_7020,N_5922,N_5967);
or U7021 (N_7021,N_5188,N_5750);
nor U7022 (N_7022,N_4763,N_4720);
nor U7023 (N_7023,N_4219,N_4247);
and U7024 (N_7024,N_4113,N_5947);
nand U7025 (N_7025,N_4976,N_4611);
nand U7026 (N_7026,N_5283,N_4551);
nand U7027 (N_7027,N_4315,N_5945);
and U7028 (N_7028,N_4823,N_4032);
and U7029 (N_7029,N_4641,N_5272);
nor U7030 (N_7030,N_4536,N_4045);
or U7031 (N_7031,N_5220,N_4718);
nand U7032 (N_7032,N_4605,N_4690);
or U7033 (N_7033,N_4338,N_5518);
nor U7034 (N_7034,N_5907,N_5281);
or U7035 (N_7035,N_4758,N_4270);
nand U7036 (N_7036,N_5702,N_4333);
and U7037 (N_7037,N_5247,N_4204);
or U7038 (N_7038,N_4307,N_4977);
and U7039 (N_7039,N_5694,N_4063);
nand U7040 (N_7040,N_5013,N_5159);
nand U7041 (N_7041,N_4509,N_5305);
nor U7042 (N_7042,N_4635,N_5929);
or U7043 (N_7043,N_5502,N_4960);
or U7044 (N_7044,N_5438,N_4234);
and U7045 (N_7045,N_4442,N_4489);
and U7046 (N_7046,N_4492,N_5029);
nand U7047 (N_7047,N_5494,N_5586);
nand U7048 (N_7048,N_4134,N_4682);
and U7049 (N_7049,N_4855,N_5680);
and U7050 (N_7050,N_4660,N_5290);
nor U7051 (N_7051,N_5680,N_5473);
and U7052 (N_7052,N_5424,N_5132);
nor U7053 (N_7053,N_4897,N_4574);
nand U7054 (N_7054,N_4863,N_5170);
and U7055 (N_7055,N_5492,N_4443);
xor U7056 (N_7056,N_5175,N_4694);
nor U7057 (N_7057,N_5015,N_4193);
nor U7058 (N_7058,N_5676,N_4426);
nor U7059 (N_7059,N_4644,N_4789);
or U7060 (N_7060,N_5119,N_5391);
or U7061 (N_7061,N_5501,N_5764);
and U7062 (N_7062,N_5629,N_4919);
or U7063 (N_7063,N_4973,N_4409);
nand U7064 (N_7064,N_4986,N_5506);
nand U7065 (N_7065,N_5578,N_4076);
xnor U7066 (N_7066,N_5639,N_5685);
or U7067 (N_7067,N_5028,N_4991);
and U7068 (N_7068,N_4480,N_5501);
or U7069 (N_7069,N_5665,N_4135);
nand U7070 (N_7070,N_5500,N_5145);
or U7071 (N_7071,N_4657,N_5159);
nand U7072 (N_7072,N_4077,N_4588);
and U7073 (N_7073,N_5818,N_5384);
and U7074 (N_7074,N_5219,N_4708);
nand U7075 (N_7075,N_4104,N_5454);
nor U7076 (N_7076,N_4053,N_4356);
and U7077 (N_7077,N_5323,N_5664);
or U7078 (N_7078,N_4364,N_5162);
or U7079 (N_7079,N_4868,N_4494);
and U7080 (N_7080,N_4882,N_4184);
nand U7081 (N_7081,N_5241,N_5396);
nand U7082 (N_7082,N_5140,N_4325);
nand U7083 (N_7083,N_4819,N_4373);
nand U7084 (N_7084,N_5033,N_5769);
nand U7085 (N_7085,N_5655,N_5884);
nand U7086 (N_7086,N_5659,N_5356);
nor U7087 (N_7087,N_5238,N_5668);
nand U7088 (N_7088,N_4669,N_5792);
nor U7089 (N_7089,N_4441,N_5141);
and U7090 (N_7090,N_4869,N_4515);
nor U7091 (N_7091,N_5797,N_5815);
or U7092 (N_7092,N_5894,N_5449);
nand U7093 (N_7093,N_4572,N_4688);
and U7094 (N_7094,N_4893,N_5188);
nor U7095 (N_7095,N_4793,N_4384);
or U7096 (N_7096,N_4575,N_5075);
nand U7097 (N_7097,N_4582,N_4810);
or U7098 (N_7098,N_5039,N_4643);
or U7099 (N_7099,N_4422,N_4506);
nand U7100 (N_7100,N_4674,N_4285);
nor U7101 (N_7101,N_4309,N_4742);
and U7102 (N_7102,N_5315,N_5178);
or U7103 (N_7103,N_4563,N_4133);
nand U7104 (N_7104,N_4814,N_4803);
or U7105 (N_7105,N_4637,N_5979);
or U7106 (N_7106,N_5163,N_4162);
nor U7107 (N_7107,N_5626,N_4430);
or U7108 (N_7108,N_5847,N_5726);
nand U7109 (N_7109,N_5204,N_5408);
or U7110 (N_7110,N_4137,N_5409);
nor U7111 (N_7111,N_5251,N_4327);
and U7112 (N_7112,N_5128,N_5051);
or U7113 (N_7113,N_5072,N_5951);
nand U7114 (N_7114,N_4758,N_5560);
and U7115 (N_7115,N_4545,N_5199);
and U7116 (N_7116,N_5411,N_4109);
nand U7117 (N_7117,N_5501,N_4508);
and U7118 (N_7118,N_4408,N_5132);
or U7119 (N_7119,N_4688,N_5969);
nor U7120 (N_7120,N_5215,N_5669);
or U7121 (N_7121,N_5920,N_4751);
nor U7122 (N_7122,N_4251,N_4661);
nor U7123 (N_7123,N_5038,N_4199);
and U7124 (N_7124,N_4159,N_4270);
xnor U7125 (N_7125,N_5287,N_5414);
nor U7126 (N_7126,N_5918,N_5331);
nand U7127 (N_7127,N_5001,N_5160);
and U7128 (N_7128,N_4030,N_5436);
and U7129 (N_7129,N_5935,N_4508);
nand U7130 (N_7130,N_4164,N_5229);
and U7131 (N_7131,N_5904,N_4455);
or U7132 (N_7132,N_5734,N_4328);
or U7133 (N_7133,N_5683,N_5653);
nor U7134 (N_7134,N_5838,N_4091);
nand U7135 (N_7135,N_4140,N_5446);
or U7136 (N_7136,N_4573,N_4747);
nand U7137 (N_7137,N_4692,N_4058);
or U7138 (N_7138,N_5500,N_4168);
or U7139 (N_7139,N_4680,N_5312);
nand U7140 (N_7140,N_4319,N_4075);
nor U7141 (N_7141,N_5462,N_5188);
and U7142 (N_7142,N_4358,N_5751);
nand U7143 (N_7143,N_5137,N_4964);
or U7144 (N_7144,N_5675,N_5737);
or U7145 (N_7145,N_4149,N_5686);
or U7146 (N_7146,N_5389,N_5804);
or U7147 (N_7147,N_4654,N_5388);
and U7148 (N_7148,N_5077,N_5453);
or U7149 (N_7149,N_5701,N_5655);
nor U7150 (N_7150,N_4456,N_5747);
nor U7151 (N_7151,N_5460,N_4261);
nand U7152 (N_7152,N_4017,N_5472);
nand U7153 (N_7153,N_5778,N_5979);
and U7154 (N_7154,N_5160,N_4993);
nand U7155 (N_7155,N_5769,N_5348);
and U7156 (N_7156,N_5013,N_5691);
or U7157 (N_7157,N_5430,N_4446);
and U7158 (N_7158,N_4887,N_4570);
or U7159 (N_7159,N_5425,N_4862);
nand U7160 (N_7160,N_5308,N_5516);
nor U7161 (N_7161,N_4697,N_4357);
nor U7162 (N_7162,N_4139,N_4470);
or U7163 (N_7163,N_5492,N_4646);
and U7164 (N_7164,N_5404,N_5691);
or U7165 (N_7165,N_4798,N_4815);
nor U7166 (N_7166,N_4800,N_4242);
nand U7167 (N_7167,N_5627,N_5526);
nand U7168 (N_7168,N_5538,N_4775);
nor U7169 (N_7169,N_5147,N_5072);
nor U7170 (N_7170,N_4488,N_5842);
nor U7171 (N_7171,N_4767,N_4400);
nor U7172 (N_7172,N_5237,N_4834);
nor U7173 (N_7173,N_4893,N_4371);
nand U7174 (N_7174,N_4735,N_4342);
or U7175 (N_7175,N_5355,N_4224);
or U7176 (N_7176,N_4746,N_5337);
or U7177 (N_7177,N_5922,N_4607);
nand U7178 (N_7178,N_5841,N_4534);
or U7179 (N_7179,N_4112,N_4057);
nor U7180 (N_7180,N_4222,N_4276);
and U7181 (N_7181,N_5443,N_5742);
nand U7182 (N_7182,N_5357,N_5366);
nor U7183 (N_7183,N_5076,N_4485);
xor U7184 (N_7184,N_4082,N_5552);
or U7185 (N_7185,N_5365,N_5854);
nand U7186 (N_7186,N_4787,N_5242);
nand U7187 (N_7187,N_4442,N_4556);
or U7188 (N_7188,N_4139,N_4885);
xnor U7189 (N_7189,N_4771,N_5402);
nor U7190 (N_7190,N_4576,N_4126);
nand U7191 (N_7191,N_4447,N_4415);
or U7192 (N_7192,N_5093,N_5281);
nand U7193 (N_7193,N_4205,N_4819);
or U7194 (N_7194,N_4609,N_4321);
and U7195 (N_7195,N_5131,N_5106);
nor U7196 (N_7196,N_4306,N_5545);
xnor U7197 (N_7197,N_4320,N_5804);
and U7198 (N_7198,N_5094,N_5005);
nand U7199 (N_7199,N_4587,N_5137);
or U7200 (N_7200,N_4971,N_4739);
and U7201 (N_7201,N_5265,N_5898);
nor U7202 (N_7202,N_5086,N_4024);
and U7203 (N_7203,N_4136,N_4606);
and U7204 (N_7204,N_4088,N_5391);
nor U7205 (N_7205,N_4729,N_5280);
and U7206 (N_7206,N_4552,N_5579);
nor U7207 (N_7207,N_4221,N_4309);
or U7208 (N_7208,N_4920,N_4974);
nor U7209 (N_7209,N_5528,N_4387);
and U7210 (N_7210,N_4014,N_4257);
or U7211 (N_7211,N_5095,N_5047);
nand U7212 (N_7212,N_4405,N_4663);
nand U7213 (N_7213,N_4188,N_5253);
nand U7214 (N_7214,N_5471,N_4571);
and U7215 (N_7215,N_4865,N_4182);
or U7216 (N_7216,N_4592,N_4125);
or U7217 (N_7217,N_5733,N_4131);
xor U7218 (N_7218,N_5767,N_4046);
and U7219 (N_7219,N_4370,N_4357);
nor U7220 (N_7220,N_4539,N_4775);
and U7221 (N_7221,N_4717,N_5996);
and U7222 (N_7222,N_4590,N_4880);
or U7223 (N_7223,N_4391,N_5092);
nand U7224 (N_7224,N_4428,N_5099);
or U7225 (N_7225,N_5872,N_4826);
or U7226 (N_7226,N_4658,N_4827);
or U7227 (N_7227,N_4920,N_4307);
nand U7228 (N_7228,N_5778,N_5844);
nand U7229 (N_7229,N_5347,N_4384);
and U7230 (N_7230,N_5647,N_4236);
and U7231 (N_7231,N_4113,N_4893);
nor U7232 (N_7232,N_5674,N_4188);
xor U7233 (N_7233,N_5172,N_5688);
or U7234 (N_7234,N_5512,N_5162);
and U7235 (N_7235,N_5567,N_5780);
nand U7236 (N_7236,N_4349,N_4298);
nand U7237 (N_7237,N_5391,N_5071);
or U7238 (N_7238,N_5988,N_4301);
nor U7239 (N_7239,N_5115,N_5088);
and U7240 (N_7240,N_4148,N_4451);
nor U7241 (N_7241,N_5661,N_5293);
and U7242 (N_7242,N_4391,N_4382);
or U7243 (N_7243,N_4135,N_5459);
or U7244 (N_7244,N_5623,N_5567);
and U7245 (N_7245,N_4425,N_5579);
or U7246 (N_7246,N_5553,N_5175);
and U7247 (N_7247,N_4189,N_4192);
nor U7248 (N_7248,N_5331,N_5538);
or U7249 (N_7249,N_4280,N_5395);
nor U7250 (N_7250,N_5942,N_4635);
xnor U7251 (N_7251,N_4838,N_4795);
nor U7252 (N_7252,N_4267,N_4789);
nand U7253 (N_7253,N_4088,N_5121);
and U7254 (N_7254,N_5268,N_5406);
and U7255 (N_7255,N_5266,N_4237);
nor U7256 (N_7256,N_4834,N_5536);
nand U7257 (N_7257,N_5057,N_4463);
and U7258 (N_7258,N_4428,N_4787);
nand U7259 (N_7259,N_4053,N_4965);
nor U7260 (N_7260,N_5300,N_5464);
and U7261 (N_7261,N_4516,N_5917);
nor U7262 (N_7262,N_5913,N_4885);
and U7263 (N_7263,N_5563,N_5339);
or U7264 (N_7264,N_4475,N_5159);
and U7265 (N_7265,N_5326,N_4978);
nor U7266 (N_7266,N_4315,N_4732);
nand U7267 (N_7267,N_5784,N_5790);
nor U7268 (N_7268,N_5166,N_5244);
or U7269 (N_7269,N_4654,N_4855);
nor U7270 (N_7270,N_4459,N_5136);
nand U7271 (N_7271,N_5353,N_5872);
nand U7272 (N_7272,N_5181,N_5369);
nor U7273 (N_7273,N_4662,N_5599);
nor U7274 (N_7274,N_4105,N_5492);
and U7275 (N_7275,N_4776,N_5020);
or U7276 (N_7276,N_4904,N_5625);
nor U7277 (N_7277,N_4937,N_5404);
and U7278 (N_7278,N_4321,N_5743);
or U7279 (N_7279,N_4331,N_4884);
xnor U7280 (N_7280,N_5034,N_5873);
nand U7281 (N_7281,N_4221,N_5837);
or U7282 (N_7282,N_5491,N_4614);
xor U7283 (N_7283,N_4469,N_4691);
and U7284 (N_7284,N_4216,N_5564);
nand U7285 (N_7285,N_5753,N_4575);
nand U7286 (N_7286,N_4715,N_5797);
nand U7287 (N_7287,N_5787,N_5349);
or U7288 (N_7288,N_5306,N_4519);
and U7289 (N_7289,N_4804,N_4507);
nand U7290 (N_7290,N_5145,N_5261);
xor U7291 (N_7291,N_5082,N_4840);
nor U7292 (N_7292,N_4247,N_4648);
nor U7293 (N_7293,N_4764,N_5514);
and U7294 (N_7294,N_5526,N_5162);
nor U7295 (N_7295,N_4339,N_5812);
nor U7296 (N_7296,N_4475,N_5134);
nor U7297 (N_7297,N_4089,N_5521);
or U7298 (N_7298,N_5302,N_5715);
nand U7299 (N_7299,N_4856,N_4719);
nor U7300 (N_7300,N_5822,N_5837);
or U7301 (N_7301,N_4201,N_4088);
nand U7302 (N_7302,N_4602,N_4417);
or U7303 (N_7303,N_5892,N_4478);
or U7304 (N_7304,N_4402,N_4667);
nand U7305 (N_7305,N_4559,N_4364);
nand U7306 (N_7306,N_5564,N_5500);
nand U7307 (N_7307,N_5685,N_4961);
nand U7308 (N_7308,N_5236,N_5123);
or U7309 (N_7309,N_4519,N_5546);
nand U7310 (N_7310,N_4693,N_4807);
or U7311 (N_7311,N_4840,N_5456);
xnor U7312 (N_7312,N_4094,N_4099);
nand U7313 (N_7313,N_5523,N_4824);
nand U7314 (N_7314,N_4173,N_5782);
and U7315 (N_7315,N_5198,N_5171);
nor U7316 (N_7316,N_4739,N_5378);
and U7317 (N_7317,N_4747,N_4553);
and U7318 (N_7318,N_4318,N_4768);
nor U7319 (N_7319,N_4594,N_5086);
and U7320 (N_7320,N_4146,N_5467);
and U7321 (N_7321,N_4652,N_5699);
and U7322 (N_7322,N_4221,N_4822);
nor U7323 (N_7323,N_4743,N_4049);
and U7324 (N_7324,N_5580,N_4213);
nand U7325 (N_7325,N_5100,N_4995);
nand U7326 (N_7326,N_4292,N_5602);
nand U7327 (N_7327,N_5590,N_4230);
nand U7328 (N_7328,N_4802,N_4841);
or U7329 (N_7329,N_5981,N_4643);
nand U7330 (N_7330,N_5931,N_4723);
nor U7331 (N_7331,N_4030,N_4450);
or U7332 (N_7332,N_4044,N_4733);
and U7333 (N_7333,N_4584,N_4049);
and U7334 (N_7334,N_4776,N_4842);
nor U7335 (N_7335,N_5847,N_5885);
nand U7336 (N_7336,N_4151,N_5324);
nand U7337 (N_7337,N_5598,N_5357);
and U7338 (N_7338,N_5191,N_5291);
nor U7339 (N_7339,N_5332,N_4568);
nand U7340 (N_7340,N_4191,N_5729);
nor U7341 (N_7341,N_4109,N_5591);
nor U7342 (N_7342,N_5021,N_5605);
nand U7343 (N_7343,N_5698,N_5882);
or U7344 (N_7344,N_5507,N_5862);
or U7345 (N_7345,N_4125,N_4290);
nand U7346 (N_7346,N_4688,N_4800);
nand U7347 (N_7347,N_4010,N_5882);
nor U7348 (N_7348,N_4164,N_5468);
nor U7349 (N_7349,N_5844,N_5681);
or U7350 (N_7350,N_5719,N_4874);
and U7351 (N_7351,N_4817,N_5411);
or U7352 (N_7352,N_5057,N_5160);
or U7353 (N_7353,N_5718,N_5632);
nand U7354 (N_7354,N_5681,N_4765);
and U7355 (N_7355,N_4297,N_5576);
nand U7356 (N_7356,N_5428,N_4467);
nand U7357 (N_7357,N_5882,N_4402);
nor U7358 (N_7358,N_5620,N_4363);
or U7359 (N_7359,N_4913,N_5880);
nor U7360 (N_7360,N_5362,N_4622);
or U7361 (N_7361,N_4254,N_4848);
nor U7362 (N_7362,N_5054,N_4015);
nor U7363 (N_7363,N_5866,N_4240);
nand U7364 (N_7364,N_4562,N_4667);
and U7365 (N_7365,N_4931,N_4571);
nor U7366 (N_7366,N_4112,N_5980);
and U7367 (N_7367,N_4648,N_5875);
nor U7368 (N_7368,N_5135,N_5802);
nand U7369 (N_7369,N_4340,N_5049);
or U7370 (N_7370,N_4145,N_5202);
and U7371 (N_7371,N_4979,N_5852);
nand U7372 (N_7372,N_4074,N_4591);
and U7373 (N_7373,N_5166,N_4785);
nor U7374 (N_7374,N_4751,N_4235);
nand U7375 (N_7375,N_4131,N_5293);
nor U7376 (N_7376,N_5056,N_4767);
nor U7377 (N_7377,N_5494,N_4635);
nand U7378 (N_7378,N_4290,N_5780);
or U7379 (N_7379,N_4588,N_5011);
nand U7380 (N_7380,N_5560,N_4542);
nand U7381 (N_7381,N_5188,N_4141);
nor U7382 (N_7382,N_4907,N_5256);
xor U7383 (N_7383,N_4872,N_4579);
and U7384 (N_7384,N_5529,N_4413);
or U7385 (N_7385,N_4026,N_5550);
and U7386 (N_7386,N_5642,N_5135);
nor U7387 (N_7387,N_5951,N_5349);
and U7388 (N_7388,N_5731,N_4914);
and U7389 (N_7389,N_4489,N_5839);
or U7390 (N_7390,N_4492,N_4100);
and U7391 (N_7391,N_4052,N_5645);
or U7392 (N_7392,N_5822,N_5595);
or U7393 (N_7393,N_4630,N_5938);
nand U7394 (N_7394,N_5026,N_4698);
nand U7395 (N_7395,N_5267,N_5318);
nand U7396 (N_7396,N_4661,N_4929);
and U7397 (N_7397,N_5316,N_5477);
nand U7398 (N_7398,N_4694,N_4194);
or U7399 (N_7399,N_4539,N_5316);
nand U7400 (N_7400,N_5878,N_4441);
and U7401 (N_7401,N_5214,N_5539);
nand U7402 (N_7402,N_5650,N_4932);
nand U7403 (N_7403,N_5968,N_5797);
nor U7404 (N_7404,N_5840,N_5036);
nor U7405 (N_7405,N_4572,N_4119);
or U7406 (N_7406,N_5171,N_5356);
or U7407 (N_7407,N_4545,N_4560);
and U7408 (N_7408,N_5888,N_4615);
nor U7409 (N_7409,N_4735,N_4590);
xor U7410 (N_7410,N_5273,N_4161);
or U7411 (N_7411,N_5686,N_5318);
or U7412 (N_7412,N_5491,N_4523);
and U7413 (N_7413,N_4565,N_4101);
nand U7414 (N_7414,N_5883,N_5880);
nand U7415 (N_7415,N_4930,N_4594);
and U7416 (N_7416,N_5828,N_4863);
nand U7417 (N_7417,N_4665,N_5074);
nand U7418 (N_7418,N_4231,N_5285);
nor U7419 (N_7419,N_4326,N_4458);
nor U7420 (N_7420,N_5494,N_5580);
and U7421 (N_7421,N_5063,N_5365);
xnor U7422 (N_7422,N_5389,N_4132);
or U7423 (N_7423,N_4732,N_4906);
and U7424 (N_7424,N_5477,N_5913);
nor U7425 (N_7425,N_5190,N_5379);
or U7426 (N_7426,N_5363,N_4829);
nor U7427 (N_7427,N_5427,N_5892);
and U7428 (N_7428,N_4948,N_4422);
nor U7429 (N_7429,N_4887,N_4879);
nand U7430 (N_7430,N_5731,N_5723);
nand U7431 (N_7431,N_4066,N_5052);
and U7432 (N_7432,N_5987,N_5302);
nor U7433 (N_7433,N_4546,N_4994);
and U7434 (N_7434,N_4106,N_5833);
and U7435 (N_7435,N_4319,N_4748);
nand U7436 (N_7436,N_4997,N_4785);
and U7437 (N_7437,N_5674,N_4478);
nor U7438 (N_7438,N_5108,N_5697);
or U7439 (N_7439,N_4981,N_5370);
nor U7440 (N_7440,N_4008,N_5307);
nand U7441 (N_7441,N_5307,N_5863);
or U7442 (N_7442,N_5740,N_5810);
or U7443 (N_7443,N_4936,N_4606);
nand U7444 (N_7444,N_5551,N_5845);
or U7445 (N_7445,N_4308,N_4790);
nor U7446 (N_7446,N_4034,N_4948);
or U7447 (N_7447,N_5643,N_4990);
nor U7448 (N_7448,N_4009,N_4662);
and U7449 (N_7449,N_5514,N_4589);
nand U7450 (N_7450,N_5345,N_4184);
nand U7451 (N_7451,N_4557,N_5784);
nor U7452 (N_7452,N_5179,N_4948);
or U7453 (N_7453,N_4241,N_5210);
or U7454 (N_7454,N_4195,N_4511);
nor U7455 (N_7455,N_5608,N_4278);
and U7456 (N_7456,N_5090,N_5243);
and U7457 (N_7457,N_5354,N_4975);
and U7458 (N_7458,N_5770,N_4769);
and U7459 (N_7459,N_5240,N_4234);
and U7460 (N_7460,N_5413,N_5942);
and U7461 (N_7461,N_5027,N_4827);
nor U7462 (N_7462,N_5974,N_5506);
or U7463 (N_7463,N_5937,N_4883);
or U7464 (N_7464,N_5358,N_4893);
or U7465 (N_7465,N_4227,N_4018);
nand U7466 (N_7466,N_4202,N_5624);
and U7467 (N_7467,N_5186,N_5987);
and U7468 (N_7468,N_4559,N_5011);
nand U7469 (N_7469,N_5808,N_5370);
nor U7470 (N_7470,N_5897,N_4103);
or U7471 (N_7471,N_5456,N_4297);
or U7472 (N_7472,N_5319,N_4712);
nand U7473 (N_7473,N_5234,N_4275);
or U7474 (N_7474,N_4323,N_5531);
nand U7475 (N_7475,N_5693,N_5738);
and U7476 (N_7476,N_4613,N_4990);
or U7477 (N_7477,N_4518,N_5617);
or U7478 (N_7478,N_4023,N_4453);
nor U7479 (N_7479,N_5889,N_4681);
or U7480 (N_7480,N_5865,N_4406);
and U7481 (N_7481,N_4737,N_5706);
and U7482 (N_7482,N_4284,N_5717);
and U7483 (N_7483,N_5834,N_4019);
nor U7484 (N_7484,N_4676,N_5088);
nor U7485 (N_7485,N_5656,N_5457);
nor U7486 (N_7486,N_5716,N_5394);
nor U7487 (N_7487,N_4663,N_4351);
and U7488 (N_7488,N_5535,N_4798);
or U7489 (N_7489,N_5619,N_5432);
or U7490 (N_7490,N_5796,N_4227);
nand U7491 (N_7491,N_5787,N_5266);
or U7492 (N_7492,N_4338,N_4979);
nor U7493 (N_7493,N_4338,N_5780);
and U7494 (N_7494,N_4639,N_4047);
nor U7495 (N_7495,N_4173,N_5471);
nand U7496 (N_7496,N_4141,N_4683);
and U7497 (N_7497,N_4765,N_5127);
or U7498 (N_7498,N_4507,N_5152);
nor U7499 (N_7499,N_5213,N_4521);
nor U7500 (N_7500,N_4849,N_5612);
or U7501 (N_7501,N_4724,N_5611);
nand U7502 (N_7502,N_4196,N_4860);
nor U7503 (N_7503,N_4027,N_5388);
nand U7504 (N_7504,N_4835,N_4954);
nor U7505 (N_7505,N_5002,N_4412);
and U7506 (N_7506,N_5577,N_5976);
and U7507 (N_7507,N_5773,N_4457);
or U7508 (N_7508,N_5400,N_4849);
nor U7509 (N_7509,N_4030,N_4923);
nor U7510 (N_7510,N_4738,N_4650);
nand U7511 (N_7511,N_5006,N_5036);
and U7512 (N_7512,N_5773,N_5686);
nand U7513 (N_7513,N_4016,N_5469);
nor U7514 (N_7514,N_5151,N_4981);
xor U7515 (N_7515,N_4308,N_4787);
and U7516 (N_7516,N_4006,N_4267);
nor U7517 (N_7517,N_4231,N_5452);
and U7518 (N_7518,N_5754,N_5544);
or U7519 (N_7519,N_4830,N_5683);
nand U7520 (N_7520,N_4079,N_5129);
or U7521 (N_7521,N_4367,N_4448);
or U7522 (N_7522,N_4617,N_5016);
and U7523 (N_7523,N_5018,N_5930);
nand U7524 (N_7524,N_4808,N_5567);
or U7525 (N_7525,N_5738,N_5962);
or U7526 (N_7526,N_5561,N_5823);
and U7527 (N_7527,N_5157,N_5146);
or U7528 (N_7528,N_5025,N_4883);
nand U7529 (N_7529,N_4047,N_5496);
nor U7530 (N_7530,N_5309,N_4823);
nor U7531 (N_7531,N_4235,N_5195);
and U7532 (N_7532,N_5348,N_4239);
nand U7533 (N_7533,N_4388,N_4053);
nand U7534 (N_7534,N_5994,N_5760);
and U7535 (N_7535,N_5813,N_5646);
or U7536 (N_7536,N_5038,N_5738);
nor U7537 (N_7537,N_5676,N_4246);
nor U7538 (N_7538,N_5035,N_4420);
nand U7539 (N_7539,N_4284,N_5000);
and U7540 (N_7540,N_4938,N_4898);
or U7541 (N_7541,N_4783,N_5821);
nor U7542 (N_7542,N_4622,N_4226);
nor U7543 (N_7543,N_4090,N_4369);
and U7544 (N_7544,N_4633,N_5550);
nand U7545 (N_7545,N_4520,N_5075);
or U7546 (N_7546,N_5828,N_4444);
nand U7547 (N_7547,N_5160,N_5987);
nor U7548 (N_7548,N_4068,N_5167);
or U7549 (N_7549,N_4064,N_4123);
nor U7550 (N_7550,N_5293,N_4364);
nor U7551 (N_7551,N_4646,N_5967);
nand U7552 (N_7552,N_5809,N_5051);
or U7553 (N_7553,N_4986,N_5037);
and U7554 (N_7554,N_5311,N_4379);
or U7555 (N_7555,N_4721,N_5881);
and U7556 (N_7556,N_5587,N_5677);
and U7557 (N_7557,N_4905,N_4495);
and U7558 (N_7558,N_4842,N_5951);
nor U7559 (N_7559,N_4961,N_4114);
and U7560 (N_7560,N_5142,N_5979);
or U7561 (N_7561,N_5718,N_5478);
xnor U7562 (N_7562,N_4631,N_5549);
xor U7563 (N_7563,N_5400,N_5353);
and U7564 (N_7564,N_4233,N_5219);
and U7565 (N_7565,N_4865,N_5999);
and U7566 (N_7566,N_4504,N_4193);
and U7567 (N_7567,N_5283,N_4128);
nand U7568 (N_7568,N_4886,N_4435);
and U7569 (N_7569,N_4056,N_4654);
xor U7570 (N_7570,N_4056,N_5531);
and U7571 (N_7571,N_5465,N_4941);
or U7572 (N_7572,N_4764,N_4532);
nand U7573 (N_7573,N_4949,N_5163);
nor U7574 (N_7574,N_5006,N_5991);
and U7575 (N_7575,N_5944,N_5830);
and U7576 (N_7576,N_5304,N_4946);
nand U7577 (N_7577,N_4753,N_5728);
and U7578 (N_7578,N_5596,N_4523);
nor U7579 (N_7579,N_5194,N_5891);
nand U7580 (N_7580,N_5190,N_5835);
nor U7581 (N_7581,N_4553,N_4612);
or U7582 (N_7582,N_5645,N_5269);
nand U7583 (N_7583,N_4371,N_4677);
and U7584 (N_7584,N_4766,N_4627);
nand U7585 (N_7585,N_4295,N_5625);
or U7586 (N_7586,N_5020,N_5799);
nor U7587 (N_7587,N_4276,N_4995);
nor U7588 (N_7588,N_5983,N_5593);
nor U7589 (N_7589,N_4173,N_5312);
nor U7590 (N_7590,N_4052,N_5271);
xnor U7591 (N_7591,N_5935,N_5419);
and U7592 (N_7592,N_4281,N_4649);
or U7593 (N_7593,N_5588,N_4441);
and U7594 (N_7594,N_5675,N_5257);
and U7595 (N_7595,N_4066,N_5937);
or U7596 (N_7596,N_5002,N_5594);
nor U7597 (N_7597,N_5816,N_5263);
nor U7598 (N_7598,N_4716,N_5513);
and U7599 (N_7599,N_4892,N_5569);
nand U7600 (N_7600,N_4655,N_5016);
nand U7601 (N_7601,N_5769,N_4322);
or U7602 (N_7602,N_5962,N_5993);
nand U7603 (N_7603,N_4650,N_4409);
nor U7604 (N_7604,N_4929,N_4881);
and U7605 (N_7605,N_4561,N_4209);
and U7606 (N_7606,N_5278,N_4997);
and U7607 (N_7607,N_5599,N_5104);
or U7608 (N_7608,N_4959,N_5028);
and U7609 (N_7609,N_5440,N_4368);
and U7610 (N_7610,N_5989,N_5061);
xor U7611 (N_7611,N_4828,N_5545);
and U7612 (N_7612,N_4461,N_5682);
and U7613 (N_7613,N_5043,N_4416);
and U7614 (N_7614,N_4875,N_5541);
and U7615 (N_7615,N_4880,N_5484);
nor U7616 (N_7616,N_5224,N_5684);
nor U7617 (N_7617,N_5214,N_4453);
or U7618 (N_7618,N_4863,N_5241);
nor U7619 (N_7619,N_4082,N_5864);
and U7620 (N_7620,N_5225,N_5266);
or U7621 (N_7621,N_4855,N_4052);
xnor U7622 (N_7622,N_4823,N_5562);
nor U7623 (N_7623,N_5086,N_4035);
xor U7624 (N_7624,N_4849,N_5356);
nor U7625 (N_7625,N_5932,N_5395);
and U7626 (N_7626,N_4215,N_4979);
or U7627 (N_7627,N_4195,N_4359);
or U7628 (N_7628,N_5234,N_4496);
or U7629 (N_7629,N_4776,N_5186);
nand U7630 (N_7630,N_5678,N_4856);
and U7631 (N_7631,N_5477,N_5268);
and U7632 (N_7632,N_4215,N_5714);
nand U7633 (N_7633,N_4119,N_4221);
nand U7634 (N_7634,N_5512,N_5306);
nor U7635 (N_7635,N_4992,N_5050);
nor U7636 (N_7636,N_4903,N_4340);
and U7637 (N_7637,N_5037,N_5743);
and U7638 (N_7638,N_4019,N_5022);
or U7639 (N_7639,N_4072,N_5064);
nand U7640 (N_7640,N_4715,N_4874);
or U7641 (N_7641,N_5650,N_4224);
and U7642 (N_7642,N_4304,N_5849);
or U7643 (N_7643,N_4955,N_5075);
and U7644 (N_7644,N_5276,N_5811);
and U7645 (N_7645,N_4334,N_5118);
nor U7646 (N_7646,N_4824,N_5701);
nand U7647 (N_7647,N_4737,N_4437);
or U7648 (N_7648,N_5390,N_5100);
or U7649 (N_7649,N_4118,N_4262);
or U7650 (N_7650,N_5522,N_4096);
nand U7651 (N_7651,N_4487,N_4570);
or U7652 (N_7652,N_5758,N_4566);
nor U7653 (N_7653,N_4316,N_5469);
and U7654 (N_7654,N_4659,N_4024);
nor U7655 (N_7655,N_4634,N_4222);
or U7656 (N_7656,N_4769,N_5026);
nand U7657 (N_7657,N_4006,N_5491);
nor U7658 (N_7658,N_5498,N_5089);
nand U7659 (N_7659,N_4835,N_4885);
nand U7660 (N_7660,N_5782,N_5357);
or U7661 (N_7661,N_4216,N_5643);
and U7662 (N_7662,N_5859,N_4046);
nor U7663 (N_7663,N_5262,N_5524);
nand U7664 (N_7664,N_5651,N_5174);
or U7665 (N_7665,N_5673,N_5392);
nor U7666 (N_7666,N_4410,N_4603);
nor U7667 (N_7667,N_4632,N_5751);
nand U7668 (N_7668,N_5719,N_5773);
and U7669 (N_7669,N_5572,N_4212);
or U7670 (N_7670,N_5311,N_5905);
nand U7671 (N_7671,N_5245,N_5831);
nand U7672 (N_7672,N_4094,N_5549);
and U7673 (N_7673,N_4052,N_4069);
and U7674 (N_7674,N_5018,N_5214);
nand U7675 (N_7675,N_4031,N_4742);
and U7676 (N_7676,N_5622,N_5165);
or U7677 (N_7677,N_5848,N_5821);
nand U7678 (N_7678,N_5120,N_5339);
nor U7679 (N_7679,N_5143,N_5965);
nand U7680 (N_7680,N_4879,N_4304);
nor U7681 (N_7681,N_5499,N_5672);
nor U7682 (N_7682,N_4489,N_5591);
and U7683 (N_7683,N_5272,N_5166);
or U7684 (N_7684,N_5739,N_4060);
and U7685 (N_7685,N_4606,N_4903);
and U7686 (N_7686,N_5015,N_4980);
nand U7687 (N_7687,N_5785,N_5299);
nor U7688 (N_7688,N_4924,N_4099);
nand U7689 (N_7689,N_4811,N_4050);
xor U7690 (N_7690,N_4277,N_4611);
nor U7691 (N_7691,N_5634,N_5469);
and U7692 (N_7692,N_5018,N_5112);
and U7693 (N_7693,N_5206,N_5909);
xor U7694 (N_7694,N_4781,N_5509);
nand U7695 (N_7695,N_5577,N_4821);
and U7696 (N_7696,N_4711,N_4492);
nor U7697 (N_7697,N_5189,N_5933);
nand U7698 (N_7698,N_4741,N_5204);
and U7699 (N_7699,N_5417,N_5861);
or U7700 (N_7700,N_4440,N_4591);
nand U7701 (N_7701,N_4488,N_5141);
nor U7702 (N_7702,N_4477,N_4883);
nand U7703 (N_7703,N_4656,N_5898);
nor U7704 (N_7704,N_4392,N_4011);
or U7705 (N_7705,N_5997,N_4737);
nand U7706 (N_7706,N_4684,N_4553);
nor U7707 (N_7707,N_5427,N_5865);
nand U7708 (N_7708,N_5320,N_5398);
nor U7709 (N_7709,N_5496,N_5404);
and U7710 (N_7710,N_5803,N_5024);
nand U7711 (N_7711,N_4051,N_4973);
nor U7712 (N_7712,N_4484,N_5864);
nand U7713 (N_7713,N_5983,N_5713);
or U7714 (N_7714,N_4925,N_5432);
nand U7715 (N_7715,N_4886,N_4369);
and U7716 (N_7716,N_4574,N_5461);
nand U7717 (N_7717,N_4063,N_4781);
and U7718 (N_7718,N_5266,N_5335);
nor U7719 (N_7719,N_4359,N_4227);
nand U7720 (N_7720,N_5216,N_5562);
or U7721 (N_7721,N_5172,N_5073);
nor U7722 (N_7722,N_4781,N_5590);
or U7723 (N_7723,N_5478,N_5953);
or U7724 (N_7724,N_4633,N_4231);
and U7725 (N_7725,N_5583,N_5239);
and U7726 (N_7726,N_5354,N_5309);
nor U7727 (N_7727,N_4252,N_4450);
nand U7728 (N_7728,N_5657,N_5345);
and U7729 (N_7729,N_4936,N_4932);
nand U7730 (N_7730,N_5806,N_5524);
nand U7731 (N_7731,N_4091,N_5163);
and U7732 (N_7732,N_5681,N_4660);
or U7733 (N_7733,N_4965,N_5689);
nand U7734 (N_7734,N_5762,N_4685);
nor U7735 (N_7735,N_4283,N_4279);
and U7736 (N_7736,N_5740,N_5002);
nand U7737 (N_7737,N_4137,N_4376);
and U7738 (N_7738,N_4235,N_4044);
nor U7739 (N_7739,N_4418,N_5579);
nor U7740 (N_7740,N_5311,N_5993);
nor U7741 (N_7741,N_5981,N_5049);
and U7742 (N_7742,N_5390,N_5462);
or U7743 (N_7743,N_4218,N_5641);
or U7744 (N_7744,N_5722,N_5060);
nor U7745 (N_7745,N_4751,N_4554);
or U7746 (N_7746,N_4201,N_5056);
or U7747 (N_7747,N_5633,N_4090);
and U7748 (N_7748,N_4044,N_4175);
nand U7749 (N_7749,N_5792,N_4416);
and U7750 (N_7750,N_5444,N_4212);
or U7751 (N_7751,N_5098,N_4077);
and U7752 (N_7752,N_4800,N_4149);
xor U7753 (N_7753,N_4720,N_5559);
or U7754 (N_7754,N_5933,N_5505);
nor U7755 (N_7755,N_5934,N_4095);
nand U7756 (N_7756,N_4497,N_5295);
nand U7757 (N_7757,N_5989,N_5051);
and U7758 (N_7758,N_5412,N_5975);
and U7759 (N_7759,N_4465,N_5043);
and U7760 (N_7760,N_4912,N_5799);
nor U7761 (N_7761,N_4441,N_4957);
nand U7762 (N_7762,N_5504,N_4361);
nor U7763 (N_7763,N_4133,N_4861);
and U7764 (N_7764,N_5121,N_5808);
or U7765 (N_7765,N_4930,N_4752);
nor U7766 (N_7766,N_4923,N_5880);
nor U7767 (N_7767,N_4233,N_5648);
or U7768 (N_7768,N_4320,N_4736);
nand U7769 (N_7769,N_5307,N_5342);
or U7770 (N_7770,N_4522,N_4432);
nor U7771 (N_7771,N_5439,N_5873);
nor U7772 (N_7772,N_4621,N_5483);
nand U7773 (N_7773,N_4741,N_5679);
nor U7774 (N_7774,N_4610,N_4269);
nand U7775 (N_7775,N_5715,N_5893);
and U7776 (N_7776,N_5749,N_5812);
nand U7777 (N_7777,N_5178,N_5238);
nor U7778 (N_7778,N_5331,N_5225);
nand U7779 (N_7779,N_4016,N_5417);
nor U7780 (N_7780,N_5823,N_4671);
nand U7781 (N_7781,N_4346,N_5861);
nand U7782 (N_7782,N_4767,N_5361);
nand U7783 (N_7783,N_5140,N_5559);
nor U7784 (N_7784,N_4720,N_4846);
nand U7785 (N_7785,N_4307,N_5437);
nand U7786 (N_7786,N_5048,N_4474);
and U7787 (N_7787,N_4176,N_4991);
and U7788 (N_7788,N_4537,N_4025);
nand U7789 (N_7789,N_5013,N_5470);
nand U7790 (N_7790,N_4433,N_4616);
or U7791 (N_7791,N_4215,N_4865);
or U7792 (N_7792,N_5563,N_4567);
or U7793 (N_7793,N_5721,N_5458);
nand U7794 (N_7794,N_4680,N_4404);
or U7795 (N_7795,N_4261,N_4787);
nand U7796 (N_7796,N_5987,N_5131);
nand U7797 (N_7797,N_5048,N_5613);
nand U7798 (N_7798,N_5410,N_5863);
or U7799 (N_7799,N_5962,N_4973);
or U7800 (N_7800,N_4027,N_5526);
or U7801 (N_7801,N_5697,N_5139);
and U7802 (N_7802,N_5458,N_4239);
or U7803 (N_7803,N_4866,N_5888);
nor U7804 (N_7804,N_4516,N_5242);
and U7805 (N_7805,N_5773,N_4686);
or U7806 (N_7806,N_4254,N_4707);
or U7807 (N_7807,N_5653,N_5930);
nand U7808 (N_7808,N_4613,N_4124);
nor U7809 (N_7809,N_4019,N_4863);
and U7810 (N_7810,N_5992,N_5012);
xor U7811 (N_7811,N_5470,N_5727);
nor U7812 (N_7812,N_5764,N_5400);
nand U7813 (N_7813,N_5317,N_4410);
or U7814 (N_7814,N_4133,N_5607);
and U7815 (N_7815,N_5967,N_4604);
or U7816 (N_7816,N_4739,N_5459);
and U7817 (N_7817,N_4792,N_4150);
and U7818 (N_7818,N_5128,N_4723);
nand U7819 (N_7819,N_5559,N_5694);
nor U7820 (N_7820,N_4447,N_5450);
nor U7821 (N_7821,N_4264,N_5654);
nor U7822 (N_7822,N_4201,N_4293);
nand U7823 (N_7823,N_4817,N_5223);
nor U7824 (N_7824,N_4350,N_5912);
nor U7825 (N_7825,N_5446,N_4847);
nand U7826 (N_7826,N_5838,N_5458);
and U7827 (N_7827,N_5201,N_5563);
or U7828 (N_7828,N_5061,N_5528);
or U7829 (N_7829,N_5878,N_4058);
nand U7830 (N_7830,N_4608,N_5782);
and U7831 (N_7831,N_4899,N_4983);
nor U7832 (N_7832,N_4565,N_4172);
and U7833 (N_7833,N_4670,N_4683);
nand U7834 (N_7834,N_5480,N_5203);
nand U7835 (N_7835,N_4794,N_5157);
nand U7836 (N_7836,N_4288,N_5956);
nand U7837 (N_7837,N_4983,N_4037);
nand U7838 (N_7838,N_5554,N_5083);
or U7839 (N_7839,N_4639,N_5625);
nand U7840 (N_7840,N_4607,N_5649);
nor U7841 (N_7841,N_5321,N_4582);
or U7842 (N_7842,N_5331,N_4313);
nor U7843 (N_7843,N_4088,N_4355);
and U7844 (N_7844,N_4475,N_4084);
nor U7845 (N_7845,N_4896,N_5618);
nand U7846 (N_7846,N_4025,N_5170);
nor U7847 (N_7847,N_5535,N_5096);
nand U7848 (N_7848,N_5733,N_5653);
nor U7849 (N_7849,N_5514,N_4766);
nand U7850 (N_7850,N_5847,N_5222);
or U7851 (N_7851,N_4244,N_4653);
and U7852 (N_7852,N_5182,N_4579);
or U7853 (N_7853,N_4321,N_5331);
and U7854 (N_7854,N_4657,N_4655);
or U7855 (N_7855,N_5423,N_5701);
or U7856 (N_7856,N_4354,N_5894);
nor U7857 (N_7857,N_5201,N_4761);
nor U7858 (N_7858,N_5829,N_5536);
or U7859 (N_7859,N_5603,N_5853);
nor U7860 (N_7860,N_5731,N_5771);
or U7861 (N_7861,N_5949,N_4809);
and U7862 (N_7862,N_4993,N_4054);
or U7863 (N_7863,N_4059,N_4254);
and U7864 (N_7864,N_5416,N_4733);
or U7865 (N_7865,N_5558,N_5053);
and U7866 (N_7866,N_4054,N_5425);
or U7867 (N_7867,N_4706,N_5874);
nand U7868 (N_7868,N_5336,N_5928);
nand U7869 (N_7869,N_5471,N_4360);
and U7870 (N_7870,N_5378,N_4798);
nor U7871 (N_7871,N_5199,N_5356);
nand U7872 (N_7872,N_5062,N_4925);
nor U7873 (N_7873,N_5195,N_4631);
nand U7874 (N_7874,N_5720,N_5733);
nor U7875 (N_7875,N_5114,N_4048);
and U7876 (N_7876,N_5153,N_4915);
or U7877 (N_7877,N_4721,N_5461);
nand U7878 (N_7878,N_5221,N_5226);
nor U7879 (N_7879,N_5016,N_4637);
nor U7880 (N_7880,N_5892,N_5825);
or U7881 (N_7881,N_4048,N_5166);
nor U7882 (N_7882,N_5528,N_5981);
or U7883 (N_7883,N_5087,N_4138);
nand U7884 (N_7884,N_4496,N_4484);
or U7885 (N_7885,N_4456,N_5798);
nor U7886 (N_7886,N_5699,N_5707);
nor U7887 (N_7887,N_4611,N_4151);
nand U7888 (N_7888,N_4954,N_4041);
and U7889 (N_7889,N_5745,N_5967);
or U7890 (N_7890,N_4694,N_5059);
and U7891 (N_7891,N_5142,N_4332);
nand U7892 (N_7892,N_5633,N_4870);
or U7893 (N_7893,N_5916,N_5712);
or U7894 (N_7894,N_4568,N_5452);
nor U7895 (N_7895,N_5410,N_4254);
and U7896 (N_7896,N_4741,N_5800);
or U7897 (N_7897,N_4205,N_4971);
or U7898 (N_7898,N_5235,N_4508);
nand U7899 (N_7899,N_4401,N_5813);
and U7900 (N_7900,N_4938,N_5331);
nand U7901 (N_7901,N_4431,N_5313);
nand U7902 (N_7902,N_4412,N_5213);
and U7903 (N_7903,N_4711,N_4750);
and U7904 (N_7904,N_4849,N_5696);
and U7905 (N_7905,N_5054,N_4425);
and U7906 (N_7906,N_4420,N_4015);
and U7907 (N_7907,N_5134,N_5303);
nand U7908 (N_7908,N_4997,N_4453);
and U7909 (N_7909,N_4847,N_4472);
nand U7910 (N_7910,N_5048,N_4478);
nor U7911 (N_7911,N_5954,N_4450);
or U7912 (N_7912,N_5627,N_5255);
or U7913 (N_7913,N_5602,N_5664);
nor U7914 (N_7914,N_5391,N_4156);
nand U7915 (N_7915,N_5861,N_5598);
nand U7916 (N_7916,N_5486,N_5679);
or U7917 (N_7917,N_4110,N_4387);
nor U7918 (N_7918,N_5640,N_4309);
or U7919 (N_7919,N_4486,N_4658);
xnor U7920 (N_7920,N_4643,N_4075);
nand U7921 (N_7921,N_5941,N_4428);
or U7922 (N_7922,N_5304,N_5290);
or U7923 (N_7923,N_4066,N_4074);
nor U7924 (N_7924,N_5771,N_4883);
and U7925 (N_7925,N_5181,N_5087);
nand U7926 (N_7926,N_4522,N_4076);
or U7927 (N_7927,N_4072,N_4399);
nand U7928 (N_7928,N_5605,N_4581);
nand U7929 (N_7929,N_4677,N_4341);
nand U7930 (N_7930,N_5555,N_5229);
and U7931 (N_7931,N_4793,N_5635);
or U7932 (N_7932,N_5337,N_5819);
and U7933 (N_7933,N_4620,N_5228);
or U7934 (N_7934,N_5912,N_5135);
xnor U7935 (N_7935,N_5916,N_5862);
nand U7936 (N_7936,N_4955,N_5806);
xor U7937 (N_7937,N_5174,N_5995);
and U7938 (N_7938,N_4887,N_4743);
nor U7939 (N_7939,N_4204,N_4035);
or U7940 (N_7940,N_5296,N_4199);
or U7941 (N_7941,N_5396,N_4446);
nor U7942 (N_7942,N_4093,N_4538);
or U7943 (N_7943,N_4064,N_4914);
and U7944 (N_7944,N_5386,N_5551);
nor U7945 (N_7945,N_5062,N_4792);
or U7946 (N_7946,N_4431,N_5347);
nand U7947 (N_7947,N_4888,N_4625);
nor U7948 (N_7948,N_5374,N_5620);
or U7949 (N_7949,N_5286,N_4458);
nor U7950 (N_7950,N_5921,N_5293);
nand U7951 (N_7951,N_5944,N_4186);
nand U7952 (N_7952,N_4984,N_4523);
nor U7953 (N_7953,N_4147,N_5738);
and U7954 (N_7954,N_5098,N_5188);
or U7955 (N_7955,N_4729,N_5176);
and U7956 (N_7956,N_5079,N_5628);
and U7957 (N_7957,N_4761,N_5456);
nand U7958 (N_7958,N_5961,N_4236);
and U7959 (N_7959,N_5074,N_5392);
nor U7960 (N_7960,N_4497,N_5101);
nand U7961 (N_7961,N_5234,N_5806);
nor U7962 (N_7962,N_4586,N_5748);
or U7963 (N_7963,N_5494,N_5343);
nor U7964 (N_7964,N_4049,N_4011);
and U7965 (N_7965,N_5846,N_5877);
or U7966 (N_7966,N_5556,N_5127);
nor U7967 (N_7967,N_5154,N_5057);
nor U7968 (N_7968,N_5824,N_4882);
nand U7969 (N_7969,N_4938,N_4994);
nand U7970 (N_7970,N_4122,N_5121);
xnor U7971 (N_7971,N_5247,N_4095);
and U7972 (N_7972,N_5424,N_4466);
and U7973 (N_7973,N_5670,N_4968);
nor U7974 (N_7974,N_4615,N_4266);
and U7975 (N_7975,N_5144,N_5460);
or U7976 (N_7976,N_4893,N_5958);
and U7977 (N_7977,N_5123,N_4077);
nor U7978 (N_7978,N_5432,N_5674);
nor U7979 (N_7979,N_4179,N_4432);
or U7980 (N_7980,N_5799,N_5234);
nand U7981 (N_7981,N_5684,N_4091);
nand U7982 (N_7982,N_5942,N_5318);
or U7983 (N_7983,N_5942,N_4602);
nor U7984 (N_7984,N_5475,N_5310);
nand U7985 (N_7985,N_5249,N_5887);
xor U7986 (N_7986,N_4815,N_5430);
nor U7987 (N_7987,N_5961,N_5470);
or U7988 (N_7988,N_4386,N_5690);
or U7989 (N_7989,N_5241,N_5570);
and U7990 (N_7990,N_5302,N_4648);
or U7991 (N_7991,N_5654,N_5584);
nor U7992 (N_7992,N_5706,N_5753);
or U7993 (N_7993,N_4943,N_4631);
nor U7994 (N_7994,N_4799,N_5111);
xor U7995 (N_7995,N_5602,N_5414);
and U7996 (N_7996,N_4394,N_4967);
or U7997 (N_7997,N_4523,N_5090);
nand U7998 (N_7998,N_4768,N_4522);
nor U7999 (N_7999,N_5062,N_4549);
and U8000 (N_8000,N_7816,N_6813);
or U8001 (N_8001,N_6981,N_6221);
xor U8002 (N_8002,N_7369,N_7104);
and U8003 (N_8003,N_6868,N_7487);
nand U8004 (N_8004,N_7960,N_6685);
nand U8005 (N_8005,N_6734,N_7761);
nand U8006 (N_8006,N_7825,N_6012);
nand U8007 (N_8007,N_7490,N_6722);
or U8008 (N_8008,N_6992,N_7562);
nand U8009 (N_8009,N_6637,N_6146);
and U8010 (N_8010,N_6015,N_6927);
nor U8011 (N_8011,N_6307,N_6894);
nor U8012 (N_8012,N_6457,N_7869);
or U8013 (N_8013,N_7031,N_6484);
or U8014 (N_8014,N_7343,N_6787);
and U8015 (N_8015,N_7096,N_7258);
or U8016 (N_8016,N_7147,N_6036);
nor U8017 (N_8017,N_6585,N_7935);
or U8018 (N_8018,N_6429,N_6797);
nor U8019 (N_8019,N_6958,N_6501);
or U8020 (N_8020,N_7182,N_7297);
nor U8021 (N_8021,N_7447,N_7330);
or U8022 (N_8022,N_7113,N_6643);
nor U8023 (N_8023,N_7638,N_7098);
and U8024 (N_8024,N_7344,N_6961);
and U8025 (N_8025,N_7668,N_6354);
nor U8026 (N_8026,N_6343,N_7066);
or U8027 (N_8027,N_6963,N_7386);
or U8028 (N_8028,N_6728,N_7662);
nor U8029 (N_8029,N_7630,N_7223);
xor U8030 (N_8030,N_7524,N_6274);
nand U8031 (N_8031,N_7106,N_7900);
or U8032 (N_8032,N_6268,N_6127);
and U8033 (N_8033,N_7008,N_7578);
nand U8034 (N_8034,N_6910,N_7418);
or U8035 (N_8035,N_7733,N_6892);
or U8036 (N_8036,N_6672,N_6689);
and U8037 (N_8037,N_6114,N_6737);
or U8038 (N_8038,N_7174,N_7639);
and U8039 (N_8039,N_7160,N_6575);
or U8040 (N_8040,N_6009,N_7795);
and U8041 (N_8041,N_6162,N_6627);
nor U8042 (N_8042,N_7671,N_6432);
or U8043 (N_8043,N_6356,N_6298);
or U8044 (N_8044,N_7005,N_7050);
or U8045 (N_8045,N_7323,N_6156);
nand U8046 (N_8046,N_7924,N_6548);
and U8047 (N_8047,N_7191,N_6111);
nand U8048 (N_8048,N_7666,N_7209);
and U8049 (N_8049,N_7566,N_7695);
nor U8050 (N_8050,N_7164,N_7043);
nand U8051 (N_8051,N_7644,N_7509);
nand U8052 (N_8052,N_6362,N_7052);
and U8053 (N_8053,N_6906,N_7067);
or U8054 (N_8054,N_6522,N_6412);
and U8055 (N_8055,N_6302,N_7457);
or U8056 (N_8056,N_6173,N_7593);
nand U8057 (N_8057,N_7797,N_6203);
and U8058 (N_8058,N_6665,N_6855);
and U8059 (N_8059,N_6789,N_6245);
and U8060 (N_8060,N_7440,N_7766);
nor U8061 (N_8061,N_7173,N_7119);
xnor U8062 (N_8062,N_6092,N_7423);
nor U8063 (N_8063,N_6443,N_6025);
or U8064 (N_8064,N_6396,N_7422);
nor U8065 (N_8065,N_7726,N_6810);
or U8066 (N_8066,N_6930,N_6014);
and U8067 (N_8067,N_6380,N_7821);
or U8068 (N_8068,N_7632,N_6107);
nand U8069 (N_8069,N_6512,N_7988);
nand U8070 (N_8070,N_6932,N_6044);
nor U8071 (N_8071,N_6509,N_6612);
or U8072 (N_8072,N_7047,N_6229);
nor U8073 (N_8073,N_6066,N_6914);
nand U8074 (N_8074,N_6346,N_7388);
or U8075 (N_8075,N_7450,N_6902);
nor U8076 (N_8076,N_6675,N_6969);
nor U8077 (N_8077,N_7517,N_6397);
nor U8078 (N_8078,N_7172,N_6453);
and U8079 (N_8079,N_7401,N_7499);
nor U8080 (N_8080,N_6843,N_6350);
and U8081 (N_8081,N_6985,N_6223);
nor U8082 (N_8082,N_7221,N_7959);
xnor U8083 (N_8083,N_7244,N_6254);
nand U8084 (N_8084,N_6149,N_7790);
and U8085 (N_8085,N_6986,N_6565);
or U8086 (N_8086,N_7482,N_6285);
or U8087 (N_8087,N_6742,N_6904);
xor U8088 (N_8088,N_6060,N_7583);
or U8089 (N_8089,N_6681,N_7990);
and U8090 (N_8090,N_7702,N_6803);
nand U8091 (N_8091,N_7617,N_7302);
and U8092 (N_8092,N_7218,N_6760);
nor U8093 (N_8093,N_7828,N_7765);
nand U8094 (N_8094,N_6401,N_6308);
nor U8095 (N_8095,N_6937,N_6845);
nor U8096 (N_8096,N_6122,N_7186);
nor U8097 (N_8097,N_7560,N_6409);
or U8098 (N_8098,N_7752,N_7851);
or U8099 (N_8099,N_6574,N_6326);
nor U8100 (N_8100,N_7940,N_7549);
or U8101 (N_8101,N_6204,N_7425);
nand U8102 (N_8102,N_6069,N_6387);
or U8103 (N_8103,N_7925,N_7670);
and U8104 (N_8104,N_7272,N_6151);
or U8105 (N_8105,N_7682,N_7460);
or U8106 (N_8106,N_7192,N_7262);
and U8107 (N_8107,N_6253,N_7352);
nand U8108 (N_8108,N_7212,N_7665);
nand U8109 (N_8109,N_6535,N_7946);
nand U8110 (N_8110,N_6070,N_6506);
nor U8111 (N_8111,N_6200,N_6622);
and U8112 (N_8112,N_6365,N_7839);
and U8113 (N_8113,N_6828,N_7928);
or U8114 (N_8114,N_7219,N_6440);
and U8115 (N_8115,N_7176,N_7242);
nor U8116 (N_8116,N_6018,N_6135);
and U8117 (N_8117,N_7916,N_6246);
nand U8118 (N_8118,N_6849,N_6936);
nand U8119 (N_8119,N_6048,N_7781);
or U8120 (N_8120,N_6090,N_6376);
nand U8121 (N_8121,N_7166,N_7601);
nand U8122 (N_8122,N_7290,N_7546);
nor U8123 (N_8123,N_7226,N_7021);
and U8124 (N_8124,N_6481,N_7918);
nand U8125 (N_8125,N_6418,N_7110);
and U8126 (N_8126,N_7235,N_6664);
nand U8127 (N_8127,N_6769,N_7124);
nand U8128 (N_8128,N_6693,N_6402);
xor U8129 (N_8129,N_6613,N_7729);
nand U8130 (N_8130,N_7372,N_7194);
nor U8131 (N_8131,N_7348,N_7334);
nand U8132 (N_8132,N_7328,N_7347);
and U8133 (N_8133,N_7971,N_6464);
nand U8134 (N_8134,N_7070,N_7148);
nand U8135 (N_8135,N_6931,N_7999);
nand U8136 (N_8136,N_6997,N_7199);
and U8137 (N_8137,N_7234,N_6544);
nor U8138 (N_8138,N_6852,N_6820);
nand U8139 (N_8139,N_6407,N_7397);
nand U8140 (N_8140,N_7806,N_7986);
or U8141 (N_8141,N_6252,N_7462);
or U8142 (N_8142,N_7492,N_7609);
nor U8143 (N_8143,N_6141,N_6004);
nor U8144 (N_8144,N_6392,N_6829);
or U8145 (N_8145,N_7286,N_7956);
nand U8146 (N_8146,N_7108,N_6578);
nand U8147 (N_8147,N_6194,N_7970);
nor U8148 (N_8148,N_7202,N_7133);
nand U8149 (N_8149,N_7684,N_7154);
and U8150 (N_8150,N_6469,N_7426);
or U8151 (N_8151,N_7834,N_7003);
xor U8152 (N_8152,N_6877,N_7786);
xnor U8153 (N_8153,N_6287,N_7405);
and U8154 (N_8154,N_7544,N_6272);
and U8155 (N_8155,N_6752,N_7449);
nor U8156 (N_8156,N_6152,N_7421);
and U8157 (N_8157,N_7461,N_7365);
nor U8158 (N_8158,N_7255,N_6555);
or U8159 (N_8159,N_7819,N_6792);
or U8160 (N_8160,N_7149,N_7303);
or U8161 (N_8161,N_6269,N_6404);
and U8162 (N_8162,N_7811,N_6697);
nand U8163 (N_8163,N_7068,N_7929);
nand U8164 (N_8164,N_6707,N_7804);
nand U8165 (N_8165,N_7979,N_7785);
or U8166 (N_8166,N_6510,N_7885);
and U8167 (N_8167,N_6125,N_6919);
xor U8168 (N_8168,N_7884,N_7132);
nand U8169 (N_8169,N_6041,N_6026);
and U8170 (N_8170,N_6461,N_7467);
or U8171 (N_8171,N_7871,N_6130);
nor U8172 (N_8172,N_6115,N_7687);
nand U8173 (N_8173,N_7399,N_6498);
or U8174 (N_8174,N_7585,N_6449);
or U8175 (N_8175,N_7216,N_7769);
nor U8176 (N_8176,N_7139,N_7126);
and U8177 (N_8177,N_7056,N_6043);
nand U8178 (N_8178,N_7350,N_7211);
and U8179 (N_8179,N_7832,N_7553);
or U8180 (N_8180,N_6291,N_7101);
or U8181 (N_8181,N_7845,N_7650);
or U8182 (N_8182,N_7075,N_7958);
nor U8183 (N_8183,N_6772,N_6743);
nor U8184 (N_8184,N_6879,N_6732);
or U8185 (N_8185,N_6977,N_6591);
nor U8186 (N_8186,N_7739,N_7927);
xor U8187 (N_8187,N_7902,N_6933);
or U8188 (N_8188,N_6870,N_7897);
nand U8189 (N_8189,N_6867,N_7342);
nand U8190 (N_8190,N_6106,N_6242);
nand U8191 (N_8191,N_6639,N_6507);
or U8192 (N_8192,N_7531,N_7859);
nand U8193 (N_8193,N_6284,N_6875);
and U8194 (N_8194,N_6480,N_7432);
xor U8195 (N_8195,N_6206,N_6128);
and U8196 (N_8196,N_6196,N_6620);
or U8197 (N_8197,N_7952,N_7019);
nand U8198 (N_8198,N_6010,N_7510);
or U8199 (N_8199,N_7493,N_7150);
nor U8200 (N_8200,N_6995,N_6860);
nand U8201 (N_8201,N_6395,N_7264);
or U8202 (N_8202,N_6279,N_7151);
nand U8203 (N_8203,N_7146,N_6880);
or U8204 (N_8204,N_7805,N_6052);
and U8205 (N_8205,N_7201,N_7868);
nor U8206 (N_8206,N_6975,N_6465);
and U8207 (N_8207,N_6640,N_6726);
and U8208 (N_8208,N_6993,N_7308);
and U8209 (N_8209,N_6646,N_6554);
and U8210 (N_8210,N_6027,N_6598);
nor U8211 (N_8211,N_6935,N_7187);
nor U8212 (N_8212,N_7094,N_7294);
and U8213 (N_8213,N_6816,N_6372);
nor U8214 (N_8214,N_7635,N_7317);
and U8215 (N_8215,N_7236,N_6295);
or U8216 (N_8216,N_6355,N_6373);
nor U8217 (N_8217,N_7316,N_7957);
nand U8218 (N_8218,N_6609,N_6901);
and U8219 (N_8219,N_6562,N_6884);
nand U8220 (N_8220,N_7471,N_7747);
nand U8221 (N_8221,N_6594,N_6520);
nand U8222 (N_8222,N_7818,N_6065);
nor U8223 (N_8223,N_6718,N_6842);
or U8224 (N_8224,N_6164,N_7496);
nand U8225 (N_8225,N_6383,N_6903);
and U8226 (N_8226,N_7391,N_6227);
nor U8227 (N_8227,N_7331,N_7773);
and U8228 (N_8228,N_7995,N_6192);
or U8229 (N_8229,N_7200,N_6806);
nand U8230 (N_8230,N_6489,N_6228);
nand U8231 (N_8231,N_7534,N_7329);
nand U8232 (N_8232,N_7518,N_7319);
nand U8233 (N_8233,N_6034,N_7824);
and U8234 (N_8234,N_6037,N_6360);
or U8235 (N_8235,N_6629,N_7207);
or U8236 (N_8236,N_6944,N_6016);
nand U8237 (N_8237,N_6633,N_7459);
or U8238 (N_8238,N_6116,N_6299);
and U8239 (N_8239,N_6485,N_6900);
nor U8240 (N_8240,N_7587,N_7774);
and U8241 (N_8241,N_6739,N_7812);
and U8242 (N_8242,N_7972,N_7760);
or U8243 (N_8243,N_7413,N_6344);
nor U8244 (N_8244,N_7500,N_7091);
or U8245 (N_8245,N_6825,N_7469);
nand U8246 (N_8246,N_6815,N_7872);
and U8247 (N_8247,N_7646,N_7610);
and U8248 (N_8248,N_7521,N_6754);
nand U8249 (N_8249,N_6042,N_7810);
nand U8250 (N_8250,N_6193,N_7782);
nor U8251 (N_8251,N_7105,N_7455);
or U8252 (N_8252,N_7842,N_6332);
and U8253 (N_8253,N_7963,N_7919);
and U8254 (N_8254,N_7757,N_7168);
and U8255 (N_8255,N_7196,N_7243);
and U8256 (N_8256,N_7748,N_7380);
or U8257 (N_8257,N_6918,N_6165);
nor U8258 (N_8258,N_6095,N_7948);
or U8259 (N_8259,N_6329,N_7197);
and U8260 (N_8260,N_7083,N_7436);
nand U8261 (N_8261,N_7968,N_7994);
nor U8262 (N_8262,N_6100,N_6233);
nor U8263 (N_8263,N_7771,N_6865);
or U8264 (N_8264,N_6945,N_7896);
nand U8265 (N_8265,N_7131,N_6839);
nor U8266 (N_8266,N_6801,N_6478);
or U8267 (N_8267,N_7220,N_7836);
nand U8268 (N_8268,N_6539,N_7307);
and U8269 (N_8269,N_6148,N_6327);
or U8270 (N_8270,N_7820,N_6924);
nor U8271 (N_8271,N_7442,N_6922);
nor U8272 (N_8272,N_6784,N_7356);
nand U8273 (N_8273,N_6955,N_6124);
or U8274 (N_8274,N_7627,N_6369);
and U8275 (N_8275,N_6261,N_7273);
nor U8276 (N_8276,N_7177,N_7858);
nor U8277 (N_8277,N_7511,N_7720);
or U8278 (N_8278,N_6776,N_7306);
and U8279 (N_8279,N_7557,N_6790);
or U8280 (N_8280,N_7345,N_7975);
nand U8281 (N_8281,N_7370,N_6800);
or U8282 (N_8282,N_7336,N_7606);
or U8283 (N_8283,N_7964,N_7679);
nand U8284 (N_8284,N_6998,N_6911);
nand U8285 (N_8285,N_7338,N_6439);
nor U8286 (N_8286,N_7826,N_6972);
nor U8287 (N_8287,N_6292,N_6472);
nand U8288 (N_8288,N_7983,N_7530);
nand U8289 (N_8289,N_7980,N_6731);
and U8290 (N_8290,N_7755,N_6405);
xor U8291 (N_8291,N_6526,N_7374);
or U8292 (N_8292,N_7167,N_7522);
or U8293 (N_8293,N_7115,N_7751);
nor U8294 (N_8294,N_7414,N_7038);
or U8295 (N_8295,N_7894,N_7802);
and U8296 (N_8296,N_7574,N_7570);
nor U8297 (N_8297,N_6808,N_7508);
nand U8298 (N_8298,N_7181,N_7248);
and U8299 (N_8299,N_6802,N_6436);
nor U8300 (N_8300,N_7830,N_6452);
nor U8301 (N_8301,N_6729,N_7822);
nand U8302 (N_8302,N_7602,N_6331);
nor U8303 (N_8303,N_7238,N_6202);
or U8304 (N_8304,N_6798,N_7387);
and U8305 (N_8305,N_6614,N_6420);
and U8306 (N_8306,N_6305,N_6477);
nand U8307 (N_8307,N_7920,N_7034);
xor U8308 (N_8308,N_7799,N_7892);
nor U8309 (N_8309,N_6517,N_6736);
or U8310 (N_8310,N_6278,N_6753);
nand U8311 (N_8311,N_6414,N_7018);
nor U8312 (N_8312,N_7648,N_7366);
nor U8313 (N_8313,N_6750,N_7295);
and U8314 (N_8314,N_7375,N_6866);
or U8315 (N_8315,N_6471,N_7520);
nand U8316 (N_8316,N_6965,N_6167);
nor U8317 (N_8317,N_6530,N_6231);
or U8318 (N_8318,N_6851,N_7502);
nand U8319 (N_8319,N_7180,N_7441);
and U8320 (N_8320,N_7603,N_7853);
or U8321 (N_8321,N_7077,N_7228);
nor U8322 (N_8322,N_7984,N_6210);
nor U8323 (N_8323,N_7481,N_6301);
nor U8324 (N_8324,N_7667,N_7762);
nor U8325 (N_8325,N_6078,N_6213);
nand U8326 (N_8326,N_6119,N_7656);
and U8327 (N_8327,N_7850,N_7783);
nand U8328 (N_8328,N_7128,N_7582);
nor U8329 (N_8329,N_7663,N_7398);
and U8330 (N_8330,N_6054,N_6692);
nor U8331 (N_8331,N_6938,N_7277);
and U8332 (N_8332,N_7183,N_7363);
nand U8333 (N_8333,N_6764,N_7099);
nand U8334 (N_8334,N_6438,N_7753);
and U8335 (N_8335,N_7867,N_7296);
or U8336 (N_8336,N_6207,N_6602);
nand U8337 (N_8337,N_7358,N_6593);
or U8338 (N_8338,N_7476,N_7558);
nor U8339 (N_8339,N_7246,N_6641);
nand U8340 (N_8340,N_6587,N_6701);
or U8341 (N_8341,N_6616,N_7614);
nor U8342 (N_8342,N_7905,N_7835);
nand U8343 (N_8343,N_7263,N_6031);
or U8344 (N_8344,N_6670,N_6170);
or U8345 (N_8345,N_6759,N_7093);
or U8346 (N_8346,N_6072,N_7324);
nand U8347 (N_8347,N_7592,N_6059);
nand U8348 (N_8348,N_7179,N_6183);
nand U8349 (N_8349,N_7643,N_7672);
nand U8350 (N_8350,N_6774,N_6419);
nor U8351 (N_8351,N_6497,N_6184);
nor U8352 (N_8352,N_6131,N_7410);
nand U8353 (N_8353,N_6710,N_6628);
or U8354 (N_8354,N_7655,N_6094);
or U8355 (N_8355,N_7694,N_6493);
nand U8356 (N_8356,N_7225,N_7775);
or U8357 (N_8357,N_7749,N_6767);
nor U8358 (N_8358,N_6294,N_6896);
or U8359 (N_8359,N_7991,N_6603);
and U8360 (N_8360,N_7466,N_6428);
or U8361 (N_8361,N_7784,N_6573);
and U8362 (N_8362,N_6123,N_6046);
or U8363 (N_8363,N_7210,N_7256);
nand U8364 (N_8364,N_6596,N_6775);
nor U8365 (N_8365,N_7321,N_6260);
nor U8366 (N_8366,N_7675,N_7379);
nor U8367 (N_8367,N_7727,N_6656);
nor U8368 (N_8368,N_7163,N_6385);
and U8369 (N_8369,N_6290,N_6926);
nor U8370 (N_8370,N_6258,N_7333);
nor U8371 (N_8371,N_6818,N_6198);
or U8372 (N_8372,N_7116,N_7454);
or U8373 (N_8373,N_6540,N_7477);
nor U8374 (N_8374,N_7923,N_7962);
nand U8375 (N_8375,N_7605,N_6721);
and U8376 (N_8376,N_6674,N_6177);
and U8377 (N_8377,N_6495,N_6608);
nand U8378 (N_8378,N_6964,N_6543);
and U8379 (N_8379,N_7580,N_6623);
or U8380 (N_8380,N_6248,N_7322);
nand U8381 (N_8381,N_6516,N_7910);
nand U8382 (N_8382,N_6921,N_7428);
nor U8383 (N_8383,N_7504,N_6869);
and U8384 (N_8384,N_6878,N_7063);
or U8385 (N_8385,N_6545,N_6306);
xor U8386 (N_8386,N_6661,N_7898);
nand U8387 (N_8387,N_7184,N_7584);
nand U8388 (N_8388,N_7542,N_7165);
nand U8389 (N_8389,N_6474,N_6057);
nand U8390 (N_8390,N_7082,N_6102);
or U8391 (N_8391,N_7230,N_6142);
and U8392 (N_8392,N_6197,N_6342);
nor U8393 (N_8393,N_7190,N_6503);
nor U8394 (N_8394,N_6804,N_6208);
nor U8395 (N_8395,N_7848,N_6886);
nand U8396 (N_8396,N_6368,N_7171);
nor U8397 (N_8397,N_6505,N_7152);
nor U8398 (N_8398,N_6617,N_7373);
or U8399 (N_8399,N_6479,N_6834);
nand U8400 (N_8400,N_7059,N_7028);
nor U8401 (N_8401,N_6652,N_6099);
and U8402 (N_8402,N_6833,N_7301);
and U8403 (N_8403,N_6442,N_7114);
xor U8404 (N_8404,N_6864,N_7621);
nor U8405 (N_8405,N_6606,N_7046);
nor U8406 (N_8406,N_6755,N_7976);
or U8407 (N_8407,N_6630,N_6668);
and U8408 (N_8408,N_6393,N_6984);
nor U8409 (N_8409,N_6648,N_7393);
or U8410 (N_8410,N_7376,N_7279);
nor U8411 (N_8411,N_7710,N_6313);
nor U8412 (N_8412,N_7268,N_7887);
nor U8413 (N_8413,N_7705,N_6741);
nand U8414 (N_8414,N_7536,N_7862);
or U8415 (N_8415,N_7483,N_7943);
or U8416 (N_8416,N_7314,N_7161);
nor U8417 (N_8417,N_6348,N_7416);
nor U8418 (N_8418,N_7793,N_6882);
and U8419 (N_8419,N_6421,N_7299);
or U8420 (N_8420,N_7657,N_7291);
or U8421 (N_8421,N_7117,N_7178);
or U8422 (N_8422,N_7355,N_6255);
and U8423 (N_8423,N_6605,N_7403);
and U8424 (N_8424,N_7275,N_7654);
nor U8425 (N_8425,N_7844,N_7876);
xnor U8426 (N_8426,N_6377,N_6055);
and U8427 (N_8427,N_6595,N_6973);
or U8428 (N_8428,N_7882,N_7915);
nor U8429 (N_8429,N_7516,N_6336);
and U8430 (N_8430,N_6688,N_7776);
or U8431 (N_8431,N_6399,N_7563);
or U8432 (N_8432,N_6347,N_6422);
nand U8433 (N_8433,N_6270,N_6607);
nor U8434 (N_8434,N_6067,N_7554);
and U8435 (N_8435,N_6007,N_6045);
nand U8436 (N_8436,N_7057,N_6660);
nor U8437 (N_8437,N_7037,N_6653);
nor U8438 (N_8438,N_6858,N_7015);
nand U8439 (N_8439,N_7458,N_6424);
nand U8440 (N_8440,N_7633,N_7852);
xnor U8441 (N_8441,N_6638,N_6013);
nor U8442 (N_8442,N_6243,N_7326);
or U8443 (N_8443,N_6691,N_6035);
nand U8444 (N_8444,N_7907,N_7287);
nor U8445 (N_8445,N_6188,N_6083);
or U8446 (N_8446,N_6618,N_7445);
or U8447 (N_8447,N_7332,N_6887);
nor U8448 (N_8448,N_6039,N_7266);
nand U8449 (N_8449,N_6462,N_7588);
and U8450 (N_8450,N_6564,N_7860);
nor U8451 (N_8451,N_6657,N_6658);
or U8452 (N_8452,N_7026,N_7719);
and U8453 (N_8453,N_6058,N_6821);
nor U8454 (N_8454,N_6671,N_6502);
nor U8455 (N_8455,N_7764,N_7788);
and U8456 (N_8456,N_6236,N_7661);
nor U8457 (N_8457,N_6021,N_6030);
and U8458 (N_8458,N_6650,N_7722);
nand U8459 (N_8459,N_6724,N_7559);
nor U8460 (N_8460,N_7740,N_7505);
and U8461 (N_8461,N_7974,N_7489);
nor U8462 (N_8462,N_6987,N_6020);
nand U8463 (N_8463,N_6073,N_7660);
or U8464 (N_8464,N_6435,N_7224);
nand U8465 (N_8465,N_7807,N_7053);
nor U8466 (N_8466,N_6777,N_6703);
and U8467 (N_8467,N_7889,N_6160);
nor U8468 (N_8468,N_6029,N_7817);
nor U8469 (N_8469,N_7080,N_6704);
nor U8470 (N_8470,N_6735,N_7311);
or U8471 (N_8471,N_6154,N_7042);
nor U8472 (N_8472,N_6430,N_6000);
nand U8473 (N_8473,N_7261,N_7515);
nand U8474 (N_8474,N_6621,N_6256);
or U8475 (N_8475,N_6238,N_7231);
and U8476 (N_8476,N_6956,N_7615);
xnor U8477 (N_8477,N_7512,N_6928);
nor U8478 (N_8478,N_6071,N_6216);
nor U8479 (N_8479,N_6444,N_7404);
or U8480 (N_8480,N_7253,N_6455);
or U8481 (N_8481,N_7598,N_7006);
or U8482 (N_8482,N_7170,N_6168);
nand U8483 (N_8483,N_6979,N_7407);
and U8484 (N_8484,N_7020,N_7427);
nand U8485 (N_8485,N_6615,N_7125);
or U8486 (N_8486,N_7434,N_6276);
or U8487 (N_8487,N_6143,N_7881);
nor U8488 (N_8488,N_7745,N_7547);
nor U8489 (N_8489,N_6230,N_7589);
and U8490 (N_8490,N_7215,N_7550);
or U8491 (N_8491,N_7137,N_7129);
nand U8492 (N_8492,N_6224,N_6683);
or U8493 (N_8493,N_6853,N_7641);
nor U8494 (N_8494,N_7967,N_6569);
and U8495 (N_8495,N_6163,N_6913);
and U8496 (N_8496,N_7686,N_6050);
or U8497 (N_8497,N_7856,N_6323);
nor U8498 (N_8498,N_6239,N_6219);
and U8499 (N_8499,N_6631,N_7634);
and U8500 (N_8500,N_7778,N_6716);
nor U8501 (N_8501,N_7362,N_6001);
nand U8502 (N_8502,N_6996,N_7913);
and U8503 (N_8503,N_6171,N_6519);
or U8504 (N_8504,N_7051,N_7613);
nor U8505 (N_8505,N_6725,N_6680);
nand U8506 (N_8506,N_6390,N_6179);
and U8507 (N_8507,N_6780,N_7541);
and U8508 (N_8508,N_6838,N_7250);
or U8509 (N_8509,N_7346,N_7855);
or U8510 (N_8510,N_7864,N_7877);
or U8511 (N_8511,N_7402,N_6335);
and U8512 (N_8512,N_6571,N_6632);
and U8513 (N_8513,N_7010,N_6642);
or U8514 (N_8514,N_6304,N_7313);
and U8515 (N_8515,N_6317,N_7624);
and U8516 (N_8516,N_6488,N_7870);
nand U8517 (N_8517,N_7140,N_7936);
or U8518 (N_8518,N_7280,N_7750);
nor U8519 (N_8519,N_6706,N_7744);
and U8520 (N_8520,N_7696,N_6002);
nand U8521 (N_8521,N_7120,N_7941);
xnor U8522 (N_8522,N_7829,N_7188);
and U8523 (N_8523,N_6720,N_6563);
or U8524 (N_8524,N_6133,N_6403);
nand U8525 (N_8525,N_7136,N_7770);
nor U8526 (N_8526,N_6281,N_7861);
or U8527 (N_8527,N_6110,N_6244);
or U8528 (N_8528,N_6592,N_6051);
or U8529 (N_8529,N_6983,N_6582);
nand U8530 (N_8530,N_6134,N_6482);
or U8531 (N_8531,N_6822,N_7939);
or U8532 (N_8532,N_7596,N_6263);
xor U8533 (N_8533,N_6600,N_6320);
nor U8534 (N_8534,N_6881,N_6651);
nand U8535 (N_8535,N_7001,N_7697);
nand U8536 (N_8536,N_6425,N_7049);
nand U8537 (N_8537,N_6534,N_6340);
nor U8538 (N_8538,N_7446,N_6819);
or U8539 (N_8539,N_7645,N_6361);
or U8540 (N_8540,N_6889,N_6586);
nor U8541 (N_8541,N_6676,N_6771);
and U8542 (N_8542,N_6084,N_7304);
and U8543 (N_8543,N_6169,N_7618);
and U8544 (N_8544,N_6490,N_6195);
nand U8545 (N_8545,N_6747,N_6859);
and U8546 (N_8546,N_6458,N_6500);
nor U8547 (N_8547,N_7480,N_7341);
nor U8548 (N_8548,N_7608,N_7060);
nand U8549 (N_8549,N_7568,N_7789);
and U8550 (N_8550,N_6912,N_6536);
or U8551 (N_8551,N_6139,N_7746);
nand U8552 (N_8552,N_6538,N_7123);
or U8553 (N_8553,N_6559,N_6063);
and U8554 (N_8554,N_6844,N_7495);
or U8555 (N_8555,N_6314,N_6277);
and U8556 (N_8556,N_6768,N_7353);
nor U8557 (N_8557,N_6024,N_7899);
and U8558 (N_8558,N_7078,N_6450);
or U8559 (N_8559,N_6841,N_6781);
nand U8560 (N_8560,N_7439,N_7071);
or U8561 (N_8561,N_7361,N_7573);
xor U8562 (N_8562,N_7742,N_7419);
and U8563 (N_8563,N_6730,N_7652);
and U8564 (N_8564,N_6518,N_7293);
nand U8565 (N_8565,N_7158,N_7843);
and U8566 (N_8566,N_7525,N_6920);
and U8567 (N_8567,N_7274,N_6666);
or U8568 (N_8568,N_6515,N_7926);
nand U8569 (N_8569,N_6417,N_6991);
and U8570 (N_8570,N_7412,N_6527);
nor U8571 (N_8571,N_7247,N_7491);
nor U8572 (N_8572,N_7711,N_6546);
or U8573 (N_8573,N_7571,N_6959);
nor U8574 (N_8574,N_6189,N_6566);
or U8575 (N_8575,N_6406,N_7048);
or U8576 (N_8576,N_6282,N_6636);
xnor U8577 (N_8577,N_7683,N_7572);
or U8578 (N_8578,N_7987,N_6283);
nand U8579 (N_8579,N_7977,N_6275);
and U8580 (N_8580,N_7269,N_7443);
nor U8581 (N_8581,N_6074,N_6962);
or U8582 (N_8582,N_7527,N_6740);
and U8583 (N_8583,N_7600,N_6663);
and U8584 (N_8584,N_6126,N_7408);
or U8585 (N_8585,N_7854,N_6909);
nor U8586 (N_8586,N_7590,N_6702);
nor U8587 (N_8587,N_6408,N_6561);
or U8588 (N_8588,N_6850,N_7704);
or U8589 (N_8589,N_7886,N_7203);
and U8590 (N_8590,N_6187,N_7095);
or U8591 (N_8591,N_7523,N_6467);
or U8592 (N_8592,N_7036,N_6068);
or U8593 (N_8593,N_7259,N_6883);
nor U8594 (N_8594,N_6040,N_6976);
nor U8595 (N_8595,N_7134,N_6303);
and U8596 (N_8596,N_6240,N_6357);
nor U8597 (N_8597,N_7193,N_7382);
xor U8598 (N_8598,N_7024,N_6686);
or U8599 (N_8599,N_6150,N_7488);
and U8600 (N_8600,N_7714,N_6374);
or U8601 (N_8601,N_6807,N_6109);
or U8602 (N_8602,N_6486,N_6744);
and U8603 (N_8603,N_6757,N_6056);
and U8604 (N_8604,N_6634,N_7827);
and U8605 (N_8605,N_7878,N_7847);
nor U8606 (N_8606,N_7846,N_6091);
and U8607 (N_8607,N_6567,N_6293);
or U8608 (N_8608,N_7716,N_6942);
or U8609 (N_8609,N_7392,N_6971);
or U8610 (N_8610,N_6398,N_7463);
nor U8611 (N_8611,N_7415,N_7961);
or U8612 (N_8612,N_6709,N_6645);
or U8613 (N_8613,N_7548,N_6779);
or U8614 (N_8614,N_7791,N_6599);
and U8615 (N_8615,N_7312,N_6840);
nor U8616 (N_8616,N_6719,N_6316);
or U8617 (N_8617,N_6990,N_6445);
or U8618 (N_8618,N_6836,N_7339);
nand U8619 (N_8619,N_6654,N_7175);
nand U8620 (N_8620,N_6118,N_6006);
nor U8621 (N_8621,N_7625,N_7400);
nor U8622 (N_8622,N_7814,N_6093);
nand U8623 (N_8623,N_6968,N_6289);
xor U8624 (N_8624,N_7949,N_7611);
xnor U8625 (N_8625,N_6019,N_7938);
and U8626 (N_8626,N_7431,N_7130);
nor U8627 (N_8627,N_7448,N_7062);
or U8628 (N_8628,N_6049,N_7283);
or U8629 (N_8629,N_6923,N_6738);
nand U8630 (N_8630,N_6960,N_7430);
xnor U8631 (N_8631,N_7813,N_7700);
nor U8632 (N_8632,N_7429,N_7647);
nor U8633 (N_8633,N_7270,N_6446);
and U8634 (N_8634,N_7681,N_6325);
and U8635 (N_8635,N_7945,N_7241);
nor U8636 (N_8636,N_6028,N_7088);
nand U8637 (N_8637,N_6644,N_6047);
nand U8638 (N_8638,N_6934,N_7367);
and U8639 (N_8639,N_7285,N_6711);
nor U8640 (N_8640,N_7044,N_6264);
or U8641 (N_8641,N_6677,N_7628);
nor U8642 (N_8642,N_7685,N_6951);
and U8643 (N_8643,N_7013,N_7498);
nand U8644 (N_8644,N_7497,N_7035);
and U8645 (N_8645,N_6076,N_7501);
nor U8646 (N_8646,N_6835,N_7767);
nand U8647 (N_8647,N_7377,N_6713);
nand U8648 (N_8648,N_6762,N_6339);
nor U8649 (N_8649,N_7631,N_7718);
nor U8650 (N_8650,N_7073,N_7389);
nor U8651 (N_8651,N_6121,N_6081);
nor U8652 (N_8652,N_6312,N_6831);
or U8653 (N_8653,N_6717,N_7737);
nand U8654 (N_8654,N_7237,N_7736);
or U8655 (N_8655,N_6416,N_7721);
nor U8656 (N_8656,N_6345,N_7622);
and U8657 (N_8657,N_7636,N_7109);
and U8658 (N_8658,N_7232,N_7837);
nand U8659 (N_8659,N_6856,N_6394);
nor U8660 (N_8660,N_6626,N_6766);
or U8661 (N_8661,N_6359,N_7908);
or U8662 (N_8662,N_6723,N_6364);
and U8663 (N_8663,N_7734,N_6694);
or U8664 (N_8664,N_7709,N_7552);
nor U8665 (N_8665,N_7676,N_6837);
nor U8666 (N_8666,N_7252,N_6415);
nand U8667 (N_8667,N_7849,N_6832);
and U8668 (N_8668,N_6053,N_7724);
xnor U8669 (N_8669,N_7282,N_6468);
and U8670 (N_8670,N_7922,N_6667);
or U8671 (N_8671,N_7768,N_7438);
and U8672 (N_8672,N_6328,N_7738);
nor U8673 (N_8673,N_7741,N_7514);
nor U8674 (N_8674,N_6241,N_7260);
xnor U8675 (N_8675,N_6655,N_6925);
or U8676 (N_8676,N_7451,N_6528);
nor U8677 (N_8677,N_6064,N_7917);
or U8678 (N_8678,N_6300,N_7688);
nand U8679 (N_8679,N_7528,N_7337);
or U8680 (N_8680,N_7658,N_6916);
nand U8681 (N_8681,N_6580,N_6448);
or U8682 (N_8682,N_6915,N_6475);
nor U8683 (N_8683,N_7653,N_7831);
nand U8684 (N_8684,N_7100,N_6266);
nor U8685 (N_8685,N_6939,N_6978);
or U8686 (N_8686,N_6032,N_6948);
nor U8687 (N_8687,N_6552,N_6363);
and U8688 (N_8688,N_6181,N_7555);
nor U8689 (N_8689,N_6008,N_6378);
and U8690 (N_8690,N_7620,N_7659);
and U8691 (N_8691,N_6161,N_6451);
and U8692 (N_8692,N_6898,N_6136);
nor U8693 (N_8693,N_6542,N_7227);
and U8694 (N_8694,N_6098,N_6103);
nand U8695 (N_8695,N_6315,N_6310);
or U8696 (N_8696,N_7086,N_7435);
nor U8697 (N_8697,N_7543,N_6745);
or U8698 (N_8698,N_7978,N_7931);
nand U8699 (N_8699,N_6296,N_7779);
and U8700 (N_8700,N_6549,N_7111);
and U8701 (N_8701,N_7561,N_7673);
or U8702 (N_8702,N_7539,N_7298);
nor U8703 (N_8703,N_7484,N_7950);
and U8704 (N_8704,N_6597,N_7903);
and U8705 (N_8705,N_7135,N_7619);
nor U8706 (N_8706,N_6218,N_6799);
and U8707 (N_8707,N_7792,N_6678);
or U8708 (N_8708,N_7623,N_7406);
or U8709 (N_8709,N_6433,N_7039);
nor U8710 (N_8710,N_6318,N_7707);
or U8711 (N_8711,N_7801,N_7315);
nand U8712 (N_8712,N_7107,N_6581);
nor U8713 (N_8713,N_6684,N_6185);
nand U8714 (N_8714,N_6097,N_6967);
or U8715 (N_8715,N_6201,N_7642);
nand U8716 (N_8716,N_6431,N_6384);
nand U8717 (N_8717,N_7996,N_7022);
nor U8718 (N_8718,N_7551,N_6523);
nand U8719 (N_8719,N_6411,N_6553);
nor U8720 (N_8720,N_6604,N_7198);
nand U8721 (N_8721,N_6949,N_6547);
or U8722 (N_8722,N_6953,N_6349);
nor U8723 (N_8723,N_6297,N_7089);
nand U8724 (N_8724,N_7076,N_7061);
and U8725 (N_8725,N_6682,N_7437);
and U8726 (N_8726,N_6531,N_6137);
nand U8727 (N_8727,N_6249,N_7267);
nor U8728 (N_8728,N_6794,N_7532);
or U8729 (N_8729,N_6205,N_7478);
nand U8730 (N_8730,N_7674,N_7384);
and U8731 (N_8731,N_6584,N_7649);
nor U8732 (N_8732,N_7743,N_7932);
nor U8733 (N_8733,N_6286,N_6257);
nand U8734 (N_8734,N_6237,N_7371);
nand U8735 (N_8735,N_6391,N_7955);
and U8736 (N_8736,N_7626,N_7934);
and U8737 (N_8737,N_7465,N_7381);
and U8738 (N_8738,N_6700,N_7815);
and U8739 (N_8739,N_6309,N_6525);
nor U8740 (N_8740,N_7157,N_7103);
nand U8741 (N_8741,N_6496,N_6215);
or U8742 (N_8742,N_6358,N_6908);
and U8743 (N_8743,N_6619,N_6508);
nor U8744 (N_8744,N_7360,N_6714);
or U8745 (N_8745,N_7914,N_6273);
or U8746 (N_8746,N_7545,N_6982);
or U8747 (N_8747,N_6947,N_6893);
nand U8748 (N_8748,N_6782,N_6062);
nand U8749 (N_8749,N_7901,N_6814);
nand U8750 (N_8750,N_6625,N_7468);
and U8751 (N_8751,N_7030,N_7787);
or U8752 (N_8752,N_7874,N_7349);
or U8753 (N_8753,N_7009,N_7616);
or U8754 (N_8754,N_6166,N_7214);
and U8755 (N_8755,N_6830,N_7863);
nor U8756 (N_8756,N_6727,N_6761);
nor U8757 (N_8757,N_6966,N_7540);
and U8758 (N_8758,N_7599,N_7189);
or U8759 (N_8759,N_7479,N_6635);
nand U8760 (N_8760,N_7033,N_7708);
and U8761 (N_8761,N_6499,N_7526);
nand U8762 (N_8762,N_7586,N_7944);
nand U8763 (N_8763,N_6235,N_7390);
and U8764 (N_8764,N_7912,N_7141);
nand U8765 (N_8765,N_7763,N_6212);
and U8766 (N_8766,N_7411,N_7240);
nor U8767 (N_8767,N_6082,N_7065);
nor U8768 (N_8768,N_6447,N_6941);
and U8769 (N_8769,N_7982,N_7156);
xor U8770 (N_8770,N_7875,N_7102);
nand U8771 (N_8771,N_6138,N_6005);
nand U8772 (N_8772,N_6382,N_7470);
or U8773 (N_8773,N_6075,N_6568);
and U8774 (N_8774,N_6765,N_6817);
and U8775 (N_8775,N_7699,N_7594);
xor U8776 (N_8776,N_6857,N_6558);
or U8777 (N_8777,N_6601,N_6338);
or U8778 (N_8778,N_6120,N_7890);
nand U8779 (N_8779,N_6324,N_6504);
nand U8780 (N_8780,N_7327,N_7565);
nor U8781 (N_8781,N_6577,N_7452);
and U8782 (N_8782,N_7254,N_6466);
or U8783 (N_8783,N_7325,N_7591);
nor U8784 (N_8784,N_6259,N_7288);
or U8785 (N_8785,N_6262,N_7072);
or U8786 (N_8786,N_7143,N_7007);
nand U8787 (N_8787,N_7595,N_7965);
nor U8788 (N_8788,N_7690,N_7014);
or U8789 (N_8789,N_7092,N_7064);
nor U8790 (N_8790,N_7420,N_6708);
nand U8791 (N_8791,N_6017,N_7651);
or U8792 (N_8792,N_6929,N_6105);
nand U8793 (N_8793,N_6529,N_7701);
xor U8794 (N_8794,N_7879,N_7997);
nand U8795 (N_8795,N_6080,N_7780);
or U8796 (N_8796,N_6456,N_7564);
or U8797 (N_8797,N_7310,N_7357);
or U8798 (N_8798,N_7385,N_6687);
and U8799 (N_8799,N_6974,N_6353);
or U8800 (N_8800,N_6888,N_6537);
and U8801 (N_8801,N_7803,N_6795);
nand U8802 (N_8802,N_7474,N_7464);
and U8803 (N_8803,N_6410,N_6389);
nor U8804 (N_8804,N_6182,N_6158);
and U8805 (N_8805,N_6698,N_6521);
or U8806 (N_8806,N_7581,N_7217);
nor U8807 (N_8807,N_6096,N_7213);
nor U8808 (N_8808,N_6895,N_6492);
nand U8809 (N_8809,N_6989,N_6890);
or U8810 (N_8810,N_6088,N_7698);
nor U8811 (N_8811,N_7993,N_6970);
or U8812 (N_8812,N_6473,N_6366);
and U8813 (N_8813,N_7069,N_7278);
nor U8814 (N_8814,N_6379,N_7084);
and U8815 (N_8815,N_7579,N_7041);
and U8816 (N_8816,N_7989,N_6003);
or U8817 (N_8817,N_7045,N_7664);
nor U8818 (N_8818,N_6226,N_6733);
or U8819 (N_8819,N_7058,N_6423);
nor U8820 (N_8820,N_7992,N_7485);
nand U8821 (N_8821,N_7364,N_7678);
or U8822 (N_8822,N_6351,N_6952);
nand U8823 (N_8823,N_6876,N_7351);
or U8824 (N_8824,N_6788,N_7204);
nor U8825 (N_8825,N_7155,N_6381);
xnor U8826 (N_8826,N_7906,N_6557);
and U8827 (N_8827,N_6863,N_6132);
or U8828 (N_8828,N_6117,N_6234);
or U8829 (N_8829,N_7731,N_7717);
nor U8830 (N_8830,N_7023,N_6513);
nand U8831 (N_8831,N_7424,N_6854);
nor U8832 (N_8832,N_7637,N_6796);
nor U8833 (N_8833,N_6999,N_7759);
and U8834 (N_8834,N_6191,N_6061);
and U8835 (N_8835,N_7276,N_6427);
or U8836 (N_8836,N_6751,N_7249);
nor U8837 (N_8837,N_6271,N_7016);
nand U8838 (N_8838,N_6550,N_7693);
nor U8839 (N_8839,N_6155,N_7025);
and U8840 (N_8840,N_6649,N_7305);
and U8841 (N_8841,N_7607,N_6211);
nor U8842 (N_8842,N_6673,N_7289);
and U8843 (N_8843,N_6232,N_7354);
and U8844 (N_8844,N_6153,N_6085);
and U8845 (N_8845,N_7567,N_6812);
nand U8846 (N_8846,N_6899,N_7145);
nand U8847 (N_8847,N_7953,N_7669);
and U8848 (N_8848,N_7735,N_7809);
nand U8849 (N_8849,N_7284,N_7713);
nand U8850 (N_8850,N_6494,N_6669);
nand U8851 (N_8851,N_7185,N_7823);
and U8852 (N_8852,N_6588,N_6763);
nor U8853 (N_8853,N_7973,N_6690);
nand U8854 (N_8854,N_6954,N_6089);
nand U8855 (N_8855,N_7841,N_7074);
and U8856 (N_8856,N_7085,N_7233);
or U8857 (N_8857,N_7703,N_7873);
nor U8858 (N_8858,N_7394,N_6805);
nand U8859 (N_8859,N_6532,N_6413);
or U8860 (N_8860,N_6321,N_6011);
and U8861 (N_8861,N_7000,N_6590);
and U8862 (N_8862,N_7229,N_6441);
and U8863 (N_8863,N_7966,N_7951);
nand U8864 (N_8864,N_7706,N_7756);
xor U8865 (N_8865,N_7138,N_6217);
nand U8866 (N_8866,N_7998,N_7629);
nand U8867 (N_8867,N_6145,N_6280);
nor U8868 (N_8868,N_7245,N_7838);
nor U8869 (N_8869,N_6288,N_6087);
or U8870 (N_8870,N_6610,N_6367);
and U8871 (N_8871,N_6570,N_6334);
nor U8872 (N_8872,N_7732,N_6463);
and U8873 (N_8873,N_6758,N_7097);
nor U8874 (N_8874,N_7292,N_7453);
nor U8875 (N_8875,N_7640,N_7142);
nor U8876 (N_8876,N_6209,N_7691);
or U8877 (N_8877,N_6101,N_7933);
nor U8878 (N_8878,N_7378,N_7604);
and U8879 (N_8879,N_6225,N_6874);
and U8880 (N_8880,N_7395,N_7122);
nand U8881 (N_8881,N_7730,N_6178);
or U8882 (N_8882,N_7027,N_6190);
or U8883 (N_8883,N_6746,N_7271);
nor U8884 (N_8884,N_7597,N_6551);
or U8885 (N_8885,N_6917,N_6679);
nand U8886 (N_8886,N_6524,N_7159);
or U8887 (N_8887,N_7320,N_6647);
and U8888 (N_8888,N_6576,N_6659);
or U8889 (N_8889,N_6897,N_6756);
and U8890 (N_8890,N_6129,N_6400);
or U8891 (N_8891,N_7144,N_6388);
and U8892 (N_8892,N_6265,N_7475);
or U8893 (N_8893,N_6579,N_7121);
and U8894 (N_8894,N_6176,N_7368);
or U8895 (N_8895,N_6846,N_7937);
and U8896 (N_8896,N_7507,N_7090);
nand U8897 (N_8897,N_7396,N_6038);
nor U8898 (N_8898,N_6699,N_6872);
nor U8899 (N_8899,N_7433,N_7715);
nor U8900 (N_8900,N_6871,N_6222);
nor U8901 (N_8901,N_6220,N_6319);
nor U8902 (N_8902,N_7055,N_7239);
nand U8903 (N_8903,N_7911,N_7891);
and U8904 (N_8904,N_7880,N_7758);
nand U8905 (N_8905,N_7954,N_6491);
and U8906 (N_8906,N_7040,N_7904);
and U8907 (N_8907,N_6483,N_7265);
nand U8908 (N_8908,N_7529,N_6514);
nor U8909 (N_8909,N_6891,N_7712);
or U8910 (N_8910,N_6250,N_7895);
or U8911 (N_8911,N_6487,N_7883);
or U8912 (N_8912,N_6624,N_7533);
and U8913 (N_8913,N_6470,N_6023);
nor U8914 (N_8914,N_7383,N_7206);
nor U8915 (N_8915,N_7575,N_6386);
and U8916 (N_8916,N_6946,N_6370);
nand U8917 (N_8917,N_7251,N_6144);
nor U8918 (N_8918,N_7162,N_6770);
or U8919 (N_8919,N_7728,N_6994);
or U8920 (N_8920,N_7865,N_6159);
or U8921 (N_8921,N_6957,N_6426);
and U8922 (N_8922,N_6791,N_7012);
or U8923 (N_8923,N_7840,N_6748);
or U8924 (N_8924,N_6214,N_7208);
nand U8925 (N_8925,N_7359,N_7692);
and U8926 (N_8926,N_7112,N_7754);
or U8927 (N_8927,N_7538,N_7794);
or U8928 (N_8928,N_7335,N_6175);
and U8929 (N_8929,N_7494,N_6454);
and U8930 (N_8930,N_7087,N_6352);
nor U8931 (N_8931,N_7222,N_7537);
nor U8932 (N_8932,N_6827,N_6511);
and U8933 (N_8933,N_6696,N_7798);
nand U8934 (N_8934,N_6077,N_7409);
nand U8935 (N_8935,N_6459,N_7417);
and U8936 (N_8936,N_6322,N_6022);
and U8937 (N_8937,N_6785,N_6104);
or U8938 (N_8938,N_7772,N_7506);
nor U8939 (N_8939,N_7195,N_6862);
and U8940 (N_8940,N_6980,N_7153);
or U8941 (N_8941,N_7800,N_6186);
nand U8942 (N_8942,N_6079,N_7011);
nor U8943 (N_8943,N_7081,N_6943);
nand U8944 (N_8944,N_7472,N_7969);
and U8945 (N_8945,N_7723,N_6611);
and U8946 (N_8946,N_7893,N_6108);
nand U8947 (N_8947,N_6861,N_6905);
or U8948 (N_8948,N_6174,N_7169);
nor U8949 (N_8949,N_6251,N_6824);
nor U8950 (N_8950,N_6988,N_6556);
nand U8951 (N_8951,N_6333,N_7118);
nand U8952 (N_8952,N_7677,N_7029);
nor U8953 (N_8953,N_7985,N_7017);
or U8954 (N_8954,N_7300,N_6907);
or U8955 (N_8955,N_6560,N_6147);
nand U8956 (N_8956,N_6786,N_6715);
and U8957 (N_8957,N_6793,N_6950);
or U8958 (N_8958,N_6033,N_7556);
and U8959 (N_8959,N_6172,N_6705);
or U8960 (N_8960,N_7921,N_7888);
and U8961 (N_8961,N_6885,N_6086);
nor U8962 (N_8962,N_7004,N_6695);
or U8963 (N_8963,N_7833,N_7909);
and U8964 (N_8964,N_6199,N_6337);
nand U8965 (N_8965,N_7777,N_7689);
nor U8966 (N_8966,N_6113,N_7947);
nor U8967 (N_8967,N_6330,N_6749);
nor U8968 (N_8968,N_6140,N_6873);
and U8969 (N_8969,N_6778,N_6940);
nand U8970 (N_8970,N_6826,N_6589);
nor U8971 (N_8971,N_7577,N_6847);
nor U8972 (N_8972,N_6112,N_7680);
nand U8973 (N_8973,N_7519,N_6157);
nand U8974 (N_8974,N_7866,N_7535);
or U8975 (N_8975,N_6662,N_7002);
or U8976 (N_8976,N_6848,N_7725);
nand U8977 (N_8977,N_6460,N_6712);
or U8978 (N_8978,N_7281,N_7808);
and U8979 (N_8979,N_7054,N_7942);
or U8980 (N_8980,N_6247,N_6267);
nor U8981 (N_8981,N_7309,N_7257);
and U8982 (N_8982,N_6476,N_7032);
or U8983 (N_8983,N_7796,N_7127);
nor U8984 (N_8984,N_6773,N_7473);
or U8985 (N_8985,N_6572,N_6811);
and U8986 (N_8986,N_7456,N_7503);
or U8987 (N_8987,N_6823,N_6809);
nor U8988 (N_8988,N_6311,N_6434);
and U8989 (N_8989,N_7612,N_6533);
or U8990 (N_8990,N_7569,N_7857);
and U8991 (N_8991,N_7205,N_7513);
and U8992 (N_8992,N_6437,N_7340);
nand U8993 (N_8993,N_7981,N_6583);
nor U8994 (N_8994,N_6180,N_6341);
or U8995 (N_8995,N_6541,N_6371);
nor U8996 (N_8996,N_6375,N_7079);
or U8997 (N_8997,N_7444,N_7486);
nor U8998 (N_8998,N_7576,N_7318);
or U8999 (N_8999,N_7930,N_6783);
and U9000 (N_9000,N_7933,N_6463);
or U9001 (N_9001,N_7013,N_7877);
nand U9002 (N_9002,N_7353,N_6083);
and U9003 (N_9003,N_7923,N_6605);
nand U9004 (N_9004,N_6654,N_7783);
or U9005 (N_9005,N_6317,N_7465);
or U9006 (N_9006,N_7425,N_6881);
or U9007 (N_9007,N_6865,N_6552);
nor U9008 (N_9008,N_7038,N_7818);
nor U9009 (N_9009,N_7549,N_6044);
nand U9010 (N_9010,N_6298,N_6944);
and U9011 (N_9011,N_7473,N_7244);
and U9012 (N_9012,N_7885,N_7979);
and U9013 (N_9013,N_7457,N_6010);
nor U9014 (N_9014,N_7462,N_7237);
nand U9015 (N_9015,N_7557,N_7089);
nor U9016 (N_9016,N_6906,N_6295);
and U9017 (N_9017,N_6566,N_7858);
or U9018 (N_9018,N_7309,N_7858);
or U9019 (N_9019,N_6198,N_7565);
or U9020 (N_9020,N_6430,N_7880);
or U9021 (N_9021,N_6835,N_7812);
and U9022 (N_9022,N_6612,N_7683);
and U9023 (N_9023,N_6654,N_7557);
and U9024 (N_9024,N_6430,N_6041);
nand U9025 (N_9025,N_7889,N_6164);
nand U9026 (N_9026,N_6703,N_6840);
or U9027 (N_9027,N_7099,N_7016);
nand U9028 (N_9028,N_6424,N_7934);
or U9029 (N_9029,N_6352,N_7375);
nand U9030 (N_9030,N_6437,N_7041);
nor U9031 (N_9031,N_7707,N_7174);
or U9032 (N_9032,N_7380,N_6891);
nand U9033 (N_9033,N_6848,N_7205);
or U9034 (N_9034,N_7600,N_7891);
nand U9035 (N_9035,N_6205,N_7004);
nor U9036 (N_9036,N_7262,N_7552);
and U9037 (N_9037,N_7688,N_6480);
xnor U9038 (N_9038,N_7993,N_6262);
nor U9039 (N_9039,N_7944,N_7983);
nor U9040 (N_9040,N_7633,N_6057);
nor U9041 (N_9041,N_6561,N_6061);
nor U9042 (N_9042,N_6103,N_7155);
nor U9043 (N_9043,N_7571,N_6295);
nand U9044 (N_9044,N_7050,N_7678);
nor U9045 (N_9045,N_7481,N_6676);
nand U9046 (N_9046,N_7200,N_7184);
nor U9047 (N_9047,N_7078,N_6531);
and U9048 (N_9048,N_7349,N_6146);
or U9049 (N_9049,N_7441,N_6412);
or U9050 (N_9050,N_6171,N_7186);
and U9051 (N_9051,N_7763,N_6983);
nand U9052 (N_9052,N_7913,N_7140);
nor U9053 (N_9053,N_6347,N_7007);
nand U9054 (N_9054,N_6132,N_6814);
nand U9055 (N_9055,N_6315,N_6973);
nand U9056 (N_9056,N_6747,N_6953);
xnor U9057 (N_9057,N_7584,N_7923);
or U9058 (N_9058,N_6967,N_7826);
nor U9059 (N_9059,N_7462,N_6423);
and U9060 (N_9060,N_6014,N_6522);
and U9061 (N_9061,N_7243,N_7524);
nand U9062 (N_9062,N_6242,N_6547);
or U9063 (N_9063,N_6947,N_7636);
and U9064 (N_9064,N_6532,N_7697);
or U9065 (N_9065,N_6468,N_6056);
or U9066 (N_9066,N_7159,N_6355);
nor U9067 (N_9067,N_6097,N_7920);
nor U9068 (N_9068,N_7036,N_6413);
and U9069 (N_9069,N_6121,N_7959);
nor U9070 (N_9070,N_6540,N_6789);
nor U9071 (N_9071,N_7224,N_6866);
or U9072 (N_9072,N_6179,N_6766);
or U9073 (N_9073,N_6103,N_7731);
nor U9074 (N_9074,N_7836,N_7007);
and U9075 (N_9075,N_7266,N_7260);
nor U9076 (N_9076,N_7579,N_7000);
and U9077 (N_9077,N_7007,N_7877);
nand U9078 (N_9078,N_7842,N_7769);
and U9079 (N_9079,N_7841,N_6113);
and U9080 (N_9080,N_7518,N_6246);
nand U9081 (N_9081,N_7949,N_6199);
and U9082 (N_9082,N_7301,N_6568);
nand U9083 (N_9083,N_6825,N_7678);
or U9084 (N_9084,N_6086,N_7909);
and U9085 (N_9085,N_7013,N_7097);
nand U9086 (N_9086,N_7085,N_6040);
or U9087 (N_9087,N_6589,N_6242);
or U9088 (N_9088,N_6142,N_6755);
and U9089 (N_9089,N_7430,N_7871);
nor U9090 (N_9090,N_7357,N_6108);
and U9091 (N_9091,N_6822,N_6674);
or U9092 (N_9092,N_7110,N_6256);
xor U9093 (N_9093,N_7083,N_6564);
or U9094 (N_9094,N_6314,N_7390);
xor U9095 (N_9095,N_7500,N_6224);
and U9096 (N_9096,N_6307,N_6614);
nand U9097 (N_9097,N_6378,N_6396);
nand U9098 (N_9098,N_7649,N_6150);
and U9099 (N_9099,N_7857,N_6926);
nand U9100 (N_9100,N_6399,N_6006);
nor U9101 (N_9101,N_6403,N_7765);
and U9102 (N_9102,N_7784,N_7264);
or U9103 (N_9103,N_7225,N_7917);
nor U9104 (N_9104,N_6871,N_7048);
or U9105 (N_9105,N_6753,N_7219);
nand U9106 (N_9106,N_6220,N_6033);
nor U9107 (N_9107,N_7303,N_6880);
nor U9108 (N_9108,N_6169,N_6599);
nor U9109 (N_9109,N_7192,N_6317);
or U9110 (N_9110,N_7780,N_7090);
or U9111 (N_9111,N_6247,N_6481);
nor U9112 (N_9112,N_6772,N_7706);
or U9113 (N_9113,N_7243,N_7433);
or U9114 (N_9114,N_6228,N_6002);
nand U9115 (N_9115,N_7520,N_6226);
nor U9116 (N_9116,N_7725,N_6560);
nand U9117 (N_9117,N_6419,N_7530);
and U9118 (N_9118,N_7497,N_6807);
nand U9119 (N_9119,N_7468,N_6005);
nor U9120 (N_9120,N_6775,N_6276);
nor U9121 (N_9121,N_6572,N_6446);
and U9122 (N_9122,N_6334,N_6852);
or U9123 (N_9123,N_7719,N_7031);
or U9124 (N_9124,N_6137,N_6311);
and U9125 (N_9125,N_6349,N_6337);
nor U9126 (N_9126,N_6800,N_6936);
or U9127 (N_9127,N_7681,N_6632);
xor U9128 (N_9128,N_7238,N_6192);
nand U9129 (N_9129,N_7984,N_6486);
nand U9130 (N_9130,N_6618,N_6270);
or U9131 (N_9131,N_6358,N_6460);
nor U9132 (N_9132,N_6591,N_6311);
xor U9133 (N_9133,N_6635,N_7664);
nand U9134 (N_9134,N_7101,N_6246);
or U9135 (N_9135,N_6276,N_6498);
or U9136 (N_9136,N_6279,N_6217);
nand U9137 (N_9137,N_7500,N_6743);
or U9138 (N_9138,N_6174,N_6253);
or U9139 (N_9139,N_6982,N_6731);
and U9140 (N_9140,N_6732,N_7542);
and U9141 (N_9141,N_6931,N_7459);
or U9142 (N_9142,N_6687,N_6586);
xnor U9143 (N_9143,N_6980,N_6053);
and U9144 (N_9144,N_6209,N_6028);
nor U9145 (N_9145,N_6394,N_7994);
and U9146 (N_9146,N_6395,N_7320);
or U9147 (N_9147,N_6549,N_6933);
nand U9148 (N_9148,N_7979,N_6249);
xnor U9149 (N_9149,N_6622,N_7500);
nand U9150 (N_9150,N_7664,N_6530);
nand U9151 (N_9151,N_6808,N_6003);
and U9152 (N_9152,N_7760,N_6299);
or U9153 (N_9153,N_6864,N_7487);
nor U9154 (N_9154,N_7944,N_6149);
nor U9155 (N_9155,N_6526,N_6421);
nor U9156 (N_9156,N_7916,N_7365);
nor U9157 (N_9157,N_7287,N_7316);
and U9158 (N_9158,N_6955,N_7917);
nand U9159 (N_9159,N_7806,N_6958);
xnor U9160 (N_9160,N_7108,N_7232);
or U9161 (N_9161,N_6946,N_7039);
nand U9162 (N_9162,N_7320,N_7369);
nand U9163 (N_9163,N_6639,N_6885);
or U9164 (N_9164,N_7189,N_7900);
and U9165 (N_9165,N_6199,N_6547);
xnor U9166 (N_9166,N_6380,N_6954);
nand U9167 (N_9167,N_6571,N_6492);
and U9168 (N_9168,N_7754,N_6276);
nand U9169 (N_9169,N_7316,N_6740);
or U9170 (N_9170,N_6938,N_7544);
or U9171 (N_9171,N_6728,N_7210);
nand U9172 (N_9172,N_7167,N_7034);
nor U9173 (N_9173,N_6561,N_7615);
or U9174 (N_9174,N_7821,N_6071);
nand U9175 (N_9175,N_6606,N_7505);
nor U9176 (N_9176,N_6514,N_7434);
and U9177 (N_9177,N_6045,N_6708);
or U9178 (N_9178,N_7687,N_6988);
and U9179 (N_9179,N_6207,N_6130);
xnor U9180 (N_9180,N_7692,N_6954);
and U9181 (N_9181,N_6454,N_6924);
xor U9182 (N_9182,N_7620,N_7922);
nor U9183 (N_9183,N_6782,N_7770);
nor U9184 (N_9184,N_7652,N_7851);
and U9185 (N_9185,N_7535,N_6285);
and U9186 (N_9186,N_7091,N_7284);
or U9187 (N_9187,N_6370,N_6142);
nor U9188 (N_9188,N_7878,N_6715);
and U9189 (N_9189,N_7445,N_6695);
nor U9190 (N_9190,N_7599,N_6212);
nand U9191 (N_9191,N_6522,N_7070);
nand U9192 (N_9192,N_6977,N_7794);
or U9193 (N_9193,N_6686,N_7946);
and U9194 (N_9194,N_7124,N_7797);
nor U9195 (N_9195,N_6538,N_7993);
nand U9196 (N_9196,N_6857,N_6950);
nand U9197 (N_9197,N_7639,N_6441);
or U9198 (N_9198,N_6040,N_6094);
nor U9199 (N_9199,N_6211,N_7737);
or U9200 (N_9200,N_6206,N_7822);
or U9201 (N_9201,N_7782,N_7467);
and U9202 (N_9202,N_6218,N_6817);
or U9203 (N_9203,N_6450,N_7093);
nand U9204 (N_9204,N_7453,N_7811);
or U9205 (N_9205,N_7675,N_6202);
nor U9206 (N_9206,N_7434,N_7187);
or U9207 (N_9207,N_7645,N_7584);
nand U9208 (N_9208,N_6971,N_7279);
or U9209 (N_9209,N_6698,N_7459);
or U9210 (N_9210,N_7905,N_7770);
nor U9211 (N_9211,N_7511,N_7359);
and U9212 (N_9212,N_7915,N_7516);
nand U9213 (N_9213,N_7233,N_7048);
nand U9214 (N_9214,N_7460,N_7716);
nand U9215 (N_9215,N_6442,N_7850);
and U9216 (N_9216,N_7838,N_7705);
and U9217 (N_9217,N_6115,N_6187);
nor U9218 (N_9218,N_6086,N_6889);
or U9219 (N_9219,N_7037,N_7023);
nand U9220 (N_9220,N_6658,N_6685);
and U9221 (N_9221,N_7729,N_7123);
or U9222 (N_9222,N_7499,N_6644);
nor U9223 (N_9223,N_7350,N_7788);
nand U9224 (N_9224,N_6036,N_7555);
or U9225 (N_9225,N_7846,N_7007);
nand U9226 (N_9226,N_6763,N_7790);
nor U9227 (N_9227,N_6655,N_6541);
nor U9228 (N_9228,N_7250,N_6434);
nand U9229 (N_9229,N_7157,N_6829);
nand U9230 (N_9230,N_7369,N_7491);
nand U9231 (N_9231,N_6019,N_6680);
nor U9232 (N_9232,N_7812,N_7496);
nor U9233 (N_9233,N_7767,N_6237);
or U9234 (N_9234,N_6467,N_7064);
nand U9235 (N_9235,N_6427,N_7917);
nor U9236 (N_9236,N_7572,N_7414);
or U9237 (N_9237,N_7763,N_6696);
nor U9238 (N_9238,N_6493,N_6462);
and U9239 (N_9239,N_7296,N_6562);
or U9240 (N_9240,N_7627,N_7988);
or U9241 (N_9241,N_6349,N_6701);
xor U9242 (N_9242,N_6060,N_7278);
nor U9243 (N_9243,N_7508,N_7674);
nand U9244 (N_9244,N_6504,N_7430);
nor U9245 (N_9245,N_7280,N_6148);
nand U9246 (N_9246,N_6686,N_7193);
nor U9247 (N_9247,N_7210,N_7293);
nand U9248 (N_9248,N_6217,N_6444);
or U9249 (N_9249,N_7641,N_7339);
and U9250 (N_9250,N_6932,N_6342);
nand U9251 (N_9251,N_7752,N_7589);
nand U9252 (N_9252,N_7871,N_6350);
and U9253 (N_9253,N_7755,N_7004);
nand U9254 (N_9254,N_6451,N_6980);
nand U9255 (N_9255,N_7693,N_6736);
nand U9256 (N_9256,N_7515,N_7010);
nand U9257 (N_9257,N_7600,N_7569);
nor U9258 (N_9258,N_6049,N_7560);
and U9259 (N_9259,N_7299,N_7824);
nor U9260 (N_9260,N_7015,N_7451);
and U9261 (N_9261,N_6401,N_7027);
and U9262 (N_9262,N_7792,N_6819);
nor U9263 (N_9263,N_6828,N_7055);
nor U9264 (N_9264,N_7882,N_7267);
nor U9265 (N_9265,N_7692,N_7360);
or U9266 (N_9266,N_6641,N_6487);
nor U9267 (N_9267,N_6198,N_6592);
nand U9268 (N_9268,N_6348,N_6446);
and U9269 (N_9269,N_6223,N_7528);
and U9270 (N_9270,N_6729,N_6934);
xor U9271 (N_9271,N_7051,N_6471);
and U9272 (N_9272,N_6754,N_7242);
nor U9273 (N_9273,N_6497,N_6917);
nand U9274 (N_9274,N_6074,N_7806);
or U9275 (N_9275,N_7041,N_7288);
and U9276 (N_9276,N_7029,N_6459);
xnor U9277 (N_9277,N_6458,N_7290);
nand U9278 (N_9278,N_7694,N_7451);
nor U9279 (N_9279,N_6216,N_6109);
and U9280 (N_9280,N_7452,N_6925);
or U9281 (N_9281,N_6853,N_7475);
and U9282 (N_9282,N_7456,N_7030);
nand U9283 (N_9283,N_6680,N_7798);
and U9284 (N_9284,N_7046,N_6502);
or U9285 (N_9285,N_7322,N_7672);
or U9286 (N_9286,N_6488,N_7938);
and U9287 (N_9287,N_7394,N_6841);
nand U9288 (N_9288,N_7486,N_6057);
and U9289 (N_9289,N_6641,N_7035);
and U9290 (N_9290,N_7962,N_7129);
and U9291 (N_9291,N_6865,N_6903);
nor U9292 (N_9292,N_6265,N_6355);
or U9293 (N_9293,N_6138,N_6997);
nor U9294 (N_9294,N_6572,N_7417);
nor U9295 (N_9295,N_7383,N_6841);
or U9296 (N_9296,N_6788,N_7894);
nand U9297 (N_9297,N_7346,N_7370);
or U9298 (N_9298,N_7934,N_7025);
or U9299 (N_9299,N_6960,N_6227);
or U9300 (N_9300,N_7022,N_7505);
and U9301 (N_9301,N_7531,N_7046);
and U9302 (N_9302,N_7382,N_6389);
or U9303 (N_9303,N_6619,N_6169);
nor U9304 (N_9304,N_7920,N_7502);
nand U9305 (N_9305,N_6938,N_6358);
or U9306 (N_9306,N_6463,N_7830);
nand U9307 (N_9307,N_6226,N_7528);
xnor U9308 (N_9308,N_6934,N_6514);
nor U9309 (N_9309,N_7918,N_6201);
nor U9310 (N_9310,N_6242,N_7582);
or U9311 (N_9311,N_6979,N_7055);
nand U9312 (N_9312,N_6963,N_6669);
or U9313 (N_9313,N_6075,N_6375);
nor U9314 (N_9314,N_6437,N_6788);
or U9315 (N_9315,N_7333,N_7494);
nor U9316 (N_9316,N_7111,N_6371);
nand U9317 (N_9317,N_7295,N_6961);
or U9318 (N_9318,N_6559,N_6459);
nand U9319 (N_9319,N_7834,N_7261);
xnor U9320 (N_9320,N_6574,N_7979);
nand U9321 (N_9321,N_6710,N_6255);
or U9322 (N_9322,N_6573,N_7096);
nor U9323 (N_9323,N_6448,N_6445);
and U9324 (N_9324,N_6021,N_6678);
nor U9325 (N_9325,N_7020,N_7304);
nor U9326 (N_9326,N_6119,N_7972);
nor U9327 (N_9327,N_7896,N_7890);
nor U9328 (N_9328,N_6038,N_7712);
and U9329 (N_9329,N_6908,N_7469);
nand U9330 (N_9330,N_6718,N_6399);
and U9331 (N_9331,N_6331,N_6804);
or U9332 (N_9332,N_7899,N_7785);
nand U9333 (N_9333,N_7899,N_7807);
and U9334 (N_9334,N_6745,N_6755);
and U9335 (N_9335,N_7470,N_6704);
nand U9336 (N_9336,N_7799,N_7625);
nand U9337 (N_9337,N_7797,N_7778);
and U9338 (N_9338,N_7253,N_7826);
nor U9339 (N_9339,N_6965,N_6316);
and U9340 (N_9340,N_6180,N_7926);
nand U9341 (N_9341,N_6008,N_7564);
nand U9342 (N_9342,N_6078,N_6354);
nor U9343 (N_9343,N_7163,N_6732);
nor U9344 (N_9344,N_6928,N_7765);
or U9345 (N_9345,N_6232,N_7864);
nand U9346 (N_9346,N_7415,N_6979);
nand U9347 (N_9347,N_7268,N_6030);
nand U9348 (N_9348,N_6666,N_6094);
nand U9349 (N_9349,N_7977,N_7078);
and U9350 (N_9350,N_6336,N_7604);
nand U9351 (N_9351,N_6662,N_6884);
and U9352 (N_9352,N_7721,N_7259);
nor U9353 (N_9353,N_6477,N_6845);
and U9354 (N_9354,N_7491,N_7987);
or U9355 (N_9355,N_7272,N_6535);
and U9356 (N_9356,N_7000,N_7632);
nand U9357 (N_9357,N_7745,N_7868);
nand U9358 (N_9358,N_6902,N_6655);
xnor U9359 (N_9359,N_6851,N_7315);
nor U9360 (N_9360,N_6227,N_6089);
or U9361 (N_9361,N_7262,N_7898);
nor U9362 (N_9362,N_7672,N_6266);
nand U9363 (N_9363,N_6114,N_6151);
and U9364 (N_9364,N_6351,N_7810);
xor U9365 (N_9365,N_6134,N_7757);
nand U9366 (N_9366,N_7984,N_6743);
nand U9367 (N_9367,N_6702,N_7579);
or U9368 (N_9368,N_6284,N_7653);
or U9369 (N_9369,N_7469,N_7384);
and U9370 (N_9370,N_7514,N_6528);
and U9371 (N_9371,N_7836,N_7734);
or U9372 (N_9372,N_6088,N_6609);
nand U9373 (N_9373,N_7095,N_7183);
and U9374 (N_9374,N_6924,N_6453);
nor U9375 (N_9375,N_7727,N_7745);
and U9376 (N_9376,N_7086,N_6908);
nand U9377 (N_9377,N_6788,N_7448);
nand U9378 (N_9378,N_6376,N_7930);
nor U9379 (N_9379,N_7073,N_7752);
and U9380 (N_9380,N_7300,N_6126);
nor U9381 (N_9381,N_6071,N_6547);
nand U9382 (N_9382,N_7615,N_6226);
and U9383 (N_9383,N_7298,N_6303);
and U9384 (N_9384,N_7116,N_6316);
nor U9385 (N_9385,N_6692,N_6507);
and U9386 (N_9386,N_6832,N_6117);
or U9387 (N_9387,N_6611,N_7318);
and U9388 (N_9388,N_6182,N_6492);
or U9389 (N_9389,N_7966,N_6695);
nand U9390 (N_9390,N_7071,N_7654);
nor U9391 (N_9391,N_7189,N_7880);
or U9392 (N_9392,N_6020,N_7210);
or U9393 (N_9393,N_6983,N_6174);
nand U9394 (N_9394,N_7880,N_7993);
nand U9395 (N_9395,N_6788,N_6561);
nor U9396 (N_9396,N_7958,N_6402);
nand U9397 (N_9397,N_6505,N_6881);
nor U9398 (N_9398,N_6990,N_7169);
or U9399 (N_9399,N_6480,N_6270);
nand U9400 (N_9400,N_7338,N_6189);
or U9401 (N_9401,N_6889,N_6227);
and U9402 (N_9402,N_6344,N_7435);
or U9403 (N_9403,N_7346,N_6861);
and U9404 (N_9404,N_6464,N_7086);
nand U9405 (N_9405,N_7895,N_6302);
nor U9406 (N_9406,N_6062,N_7716);
nand U9407 (N_9407,N_7358,N_6272);
and U9408 (N_9408,N_7233,N_7260);
nand U9409 (N_9409,N_6297,N_7059);
nor U9410 (N_9410,N_7916,N_6484);
xnor U9411 (N_9411,N_6806,N_7755);
or U9412 (N_9412,N_7165,N_6777);
nor U9413 (N_9413,N_7692,N_7056);
and U9414 (N_9414,N_7430,N_6305);
nand U9415 (N_9415,N_6638,N_6988);
and U9416 (N_9416,N_6176,N_6912);
and U9417 (N_9417,N_7120,N_6160);
and U9418 (N_9418,N_6290,N_7761);
nor U9419 (N_9419,N_6190,N_6071);
nand U9420 (N_9420,N_7184,N_6343);
nor U9421 (N_9421,N_6947,N_7960);
or U9422 (N_9422,N_7055,N_6866);
or U9423 (N_9423,N_7942,N_7380);
and U9424 (N_9424,N_7496,N_6089);
nand U9425 (N_9425,N_6113,N_7248);
nand U9426 (N_9426,N_7828,N_6479);
or U9427 (N_9427,N_6895,N_7181);
nand U9428 (N_9428,N_6692,N_6281);
nor U9429 (N_9429,N_7263,N_7314);
and U9430 (N_9430,N_7798,N_6673);
nor U9431 (N_9431,N_6751,N_7858);
nand U9432 (N_9432,N_7889,N_6226);
nand U9433 (N_9433,N_6792,N_7712);
or U9434 (N_9434,N_7498,N_6628);
or U9435 (N_9435,N_7221,N_6740);
or U9436 (N_9436,N_7341,N_6921);
nor U9437 (N_9437,N_6176,N_7608);
or U9438 (N_9438,N_6724,N_7068);
nand U9439 (N_9439,N_7019,N_7780);
and U9440 (N_9440,N_6173,N_6165);
nand U9441 (N_9441,N_6283,N_7698);
nor U9442 (N_9442,N_6883,N_7454);
and U9443 (N_9443,N_7119,N_7189);
nor U9444 (N_9444,N_7172,N_7859);
nor U9445 (N_9445,N_7186,N_7066);
nand U9446 (N_9446,N_6057,N_7514);
or U9447 (N_9447,N_6147,N_6950);
and U9448 (N_9448,N_7156,N_7470);
nand U9449 (N_9449,N_7360,N_7498);
and U9450 (N_9450,N_6853,N_6140);
nor U9451 (N_9451,N_7708,N_6499);
and U9452 (N_9452,N_6432,N_7231);
and U9453 (N_9453,N_6919,N_6573);
nand U9454 (N_9454,N_6732,N_6289);
and U9455 (N_9455,N_7302,N_6292);
nand U9456 (N_9456,N_6453,N_7632);
nor U9457 (N_9457,N_6006,N_7131);
nand U9458 (N_9458,N_6675,N_6502);
nor U9459 (N_9459,N_7643,N_7412);
nor U9460 (N_9460,N_7019,N_7782);
or U9461 (N_9461,N_7454,N_6460);
nor U9462 (N_9462,N_6537,N_7102);
and U9463 (N_9463,N_7046,N_6125);
nand U9464 (N_9464,N_6628,N_6509);
nand U9465 (N_9465,N_7409,N_6703);
and U9466 (N_9466,N_6727,N_6336);
nor U9467 (N_9467,N_7174,N_6361);
nor U9468 (N_9468,N_7213,N_7794);
nor U9469 (N_9469,N_7518,N_7098);
nor U9470 (N_9470,N_7917,N_7476);
or U9471 (N_9471,N_7186,N_7216);
or U9472 (N_9472,N_6157,N_7946);
nor U9473 (N_9473,N_6238,N_6596);
nand U9474 (N_9474,N_7673,N_7939);
or U9475 (N_9475,N_7185,N_7612);
and U9476 (N_9476,N_6879,N_6931);
nand U9477 (N_9477,N_6066,N_7147);
nor U9478 (N_9478,N_6236,N_7169);
or U9479 (N_9479,N_6377,N_7657);
and U9480 (N_9480,N_6027,N_6381);
nor U9481 (N_9481,N_7849,N_6013);
nand U9482 (N_9482,N_6015,N_6656);
nor U9483 (N_9483,N_6808,N_7178);
and U9484 (N_9484,N_7712,N_7302);
or U9485 (N_9485,N_6242,N_7139);
or U9486 (N_9486,N_7564,N_7430);
nor U9487 (N_9487,N_6499,N_7543);
nor U9488 (N_9488,N_6008,N_6392);
and U9489 (N_9489,N_6037,N_7373);
nand U9490 (N_9490,N_7444,N_7451);
and U9491 (N_9491,N_7077,N_6745);
nor U9492 (N_9492,N_6787,N_7985);
and U9493 (N_9493,N_7103,N_6210);
and U9494 (N_9494,N_6196,N_6719);
and U9495 (N_9495,N_6044,N_7299);
nand U9496 (N_9496,N_6065,N_7340);
nor U9497 (N_9497,N_7490,N_7735);
nor U9498 (N_9498,N_6453,N_7576);
or U9499 (N_9499,N_6600,N_6141);
or U9500 (N_9500,N_6606,N_6438);
nor U9501 (N_9501,N_7764,N_7741);
nand U9502 (N_9502,N_6073,N_6351);
and U9503 (N_9503,N_7649,N_7680);
and U9504 (N_9504,N_6852,N_7887);
nor U9505 (N_9505,N_6118,N_7000);
nand U9506 (N_9506,N_6788,N_7218);
or U9507 (N_9507,N_7573,N_7443);
or U9508 (N_9508,N_7752,N_6928);
and U9509 (N_9509,N_7844,N_6766);
and U9510 (N_9510,N_6342,N_7072);
nand U9511 (N_9511,N_7881,N_7873);
nor U9512 (N_9512,N_6842,N_6894);
and U9513 (N_9513,N_7771,N_7724);
and U9514 (N_9514,N_6111,N_7788);
or U9515 (N_9515,N_6190,N_6054);
nand U9516 (N_9516,N_6936,N_6523);
nor U9517 (N_9517,N_7517,N_6779);
nor U9518 (N_9518,N_7973,N_7703);
and U9519 (N_9519,N_6886,N_7377);
nand U9520 (N_9520,N_6293,N_7368);
and U9521 (N_9521,N_6420,N_7327);
nand U9522 (N_9522,N_7336,N_7759);
nand U9523 (N_9523,N_6390,N_7123);
nor U9524 (N_9524,N_7870,N_7987);
nor U9525 (N_9525,N_6489,N_7619);
nand U9526 (N_9526,N_6960,N_7002);
nand U9527 (N_9527,N_7578,N_7581);
nor U9528 (N_9528,N_7686,N_6960);
nand U9529 (N_9529,N_7998,N_7341);
and U9530 (N_9530,N_6528,N_6306);
nor U9531 (N_9531,N_6044,N_7003);
nand U9532 (N_9532,N_7628,N_7209);
or U9533 (N_9533,N_7734,N_6756);
nor U9534 (N_9534,N_7332,N_6265);
nand U9535 (N_9535,N_7401,N_7821);
or U9536 (N_9536,N_6995,N_7944);
nand U9537 (N_9537,N_6067,N_6524);
or U9538 (N_9538,N_7668,N_6406);
nor U9539 (N_9539,N_6281,N_6472);
or U9540 (N_9540,N_7180,N_6121);
or U9541 (N_9541,N_7435,N_6335);
or U9542 (N_9542,N_6183,N_7831);
or U9543 (N_9543,N_6396,N_6515);
nor U9544 (N_9544,N_6553,N_6339);
and U9545 (N_9545,N_7666,N_7502);
and U9546 (N_9546,N_6509,N_6345);
nand U9547 (N_9547,N_7029,N_6366);
and U9548 (N_9548,N_6054,N_7100);
nor U9549 (N_9549,N_6668,N_6087);
nor U9550 (N_9550,N_7709,N_6640);
and U9551 (N_9551,N_6097,N_6968);
or U9552 (N_9552,N_7869,N_7175);
nand U9553 (N_9553,N_7189,N_7070);
nor U9554 (N_9554,N_6729,N_6120);
and U9555 (N_9555,N_6545,N_6087);
or U9556 (N_9556,N_7296,N_7935);
or U9557 (N_9557,N_7390,N_7459);
or U9558 (N_9558,N_6160,N_7182);
and U9559 (N_9559,N_7325,N_7674);
or U9560 (N_9560,N_7935,N_7147);
and U9561 (N_9561,N_6090,N_6756);
or U9562 (N_9562,N_6987,N_7900);
nor U9563 (N_9563,N_7032,N_7129);
and U9564 (N_9564,N_7945,N_7359);
and U9565 (N_9565,N_6488,N_7955);
and U9566 (N_9566,N_6111,N_6236);
nand U9567 (N_9567,N_6029,N_7893);
and U9568 (N_9568,N_6067,N_6959);
nand U9569 (N_9569,N_7904,N_7977);
or U9570 (N_9570,N_7199,N_6189);
or U9571 (N_9571,N_6892,N_6926);
nand U9572 (N_9572,N_6637,N_6883);
nand U9573 (N_9573,N_7485,N_6050);
nand U9574 (N_9574,N_6240,N_7970);
nor U9575 (N_9575,N_6108,N_7370);
or U9576 (N_9576,N_7600,N_7923);
or U9577 (N_9577,N_6288,N_6306);
nand U9578 (N_9578,N_7875,N_6998);
nor U9579 (N_9579,N_6329,N_7610);
nand U9580 (N_9580,N_6414,N_6133);
nor U9581 (N_9581,N_6409,N_6953);
nor U9582 (N_9582,N_7504,N_6438);
and U9583 (N_9583,N_7798,N_6913);
or U9584 (N_9584,N_7549,N_7383);
nand U9585 (N_9585,N_6503,N_6841);
xor U9586 (N_9586,N_6637,N_7789);
and U9587 (N_9587,N_7637,N_7791);
nor U9588 (N_9588,N_7341,N_7530);
nor U9589 (N_9589,N_6394,N_7684);
xnor U9590 (N_9590,N_6046,N_7561);
or U9591 (N_9591,N_7829,N_6040);
nor U9592 (N_9592,N_7757,N_6955);
or U9593 (N_9593,N_6239,N_7374);
or U9594 (N_9594,N_7545,N_7058);
and U9595 (N_9595,N_6841,N_7732);
and U9596 (N_9596,N_7294,N_7641);
nand U9597 (N_9597,N_7928,N_6573);
or U9598 (N_9598,N_7347,N_6158);
nor U9599 (N_9599,N_6365,N_6967);
or U9600 (N_9600,N_6767,N_6063);
nand U9601 (N_9601,N_7176,N_6109);
nand U9602 (N_9602,N_6665,N_7996);
or U9603 (N_9603,N_7285,N_7449);
xor U9604 (N_9604,N_6913,N_7658);
nor U9605 (N_9605,N_7896,N_7689);
or U9606 (N_9606,N_6617,N_6327);
and U9607 (N_9607,N_6150,N_7776);
nor U9608 (N_9608,N_7060,N_7563);
or U9609 (N_9609,N_6268,N_6430);
nand U9610 (N_9610,N_7736,N_6659);
or U9611 (N_9611,N_6086,N_7186);
or U9612 (N_9612,N_6809,N_7390);
and U9613 (N_9613,N_7538,N_6624);
nor U9614 (N_9614,N_6847,N_6840);
and U9615 (N_9615,N_6690,N_7481);
nand U9616 (N_9616,N_7438,N_7056);
and U9617 (N_9617,N_6023,N_6695);
or U9618 (N_9618,N_7903,N_7601);
or U9619 (N_9619,N_7542,N_6805);
nand U9620 (N_9620,N_7637,N_7888);
nand U9621 (N_9621,N_6302,N_7458);
and U9622 (N_9622,N_6410,N_6786);
or U9623 (N_9623,N_7753,N_6295);
nand U9624 (N_9624,N_6506,N_7343);
and U9625 (N_9625,N_7106,N_6693);
nor U9626 (N_9626,N_6829,N_7878);
nand U9627 (N_9627,N_7819,N_6883);
nand U9628 (N_9628,N_6703,N_6310);
or U9629 (N_9629,N_7142,N_7423);
nor U9630 (N_9630,N_7750,N_7695);
and U9631 (N_9631,N_7561,N_7655);
nor U9632 (N_9632,N_6675,N_6136);
and U9633 (N_9633,N_6394,N_7544);
nor U9634 (N_9634,N_7866,N_7920);
nand U9635 (N_9635,N_7193,N_7125);
nor U9636 (N_9636,N_6287,N_7179);
nand U9637 (N_9637,N_6961,N_6395);
nor U9638 (N_9638,N_7622,N_6073);
or U9639 (N_9639,N_7106,N_6654);
and U9640 (N_9640,N_6931,N_6733);
nand U9641 (N_9641,N_6015,N_7271);
or U9642 (N_9642,N_6460,N_6134);
and U9643 (N_9643,N_7166,N_7464);
or U9644 (N_9644,N_6598,N_7764);
nor U9645 (N_9645,N_7767,N_7139);
and U9646 (N_9646,N_7688,N_6702);
nand U9647 (N_9647,N_6429,N_7602);
nand U9648 (N_9648,N_6001,N_6424);
nand U9649 (N_9649,N_6681,N_6033);
or U9650 (N_9650,N_6940,N_7178);
nand U9651 (N_9651,N_6993,N_6438);
nor U9652 (N_9652,N_7748,N_7674);
and U9653 (N_9653,N_6857,N_6074);
or U9654 (N_9654,N_7445,N_7808);
or U9655 (N_9655,N_6132,N_6700);
and U9656 (N_9656,N_6756,N_7658);
nand U9657 (N_9657,N_7335,N_7066);
or U9658 (N_9658,N_6307,N_6243);
nor U9659 (N_9659,N_6647,N_7185);
nand U9660 (N_9660,N_7439,N_7543);
nor U9661 (N_9661,N_6179,N_7744);
or U9662 (N_9662,N_6066,N_6518);
xnor U9663 (N_9663,N_6637,N_6491);
nand U9664 (N_9664,N_7233,N_6024);
and U9665 (N_9665,N_6603,N_7312);
nand U9666 (N_9666,N_7567,N_6585);
and U9667 (N_9667,N_6342,N_7918);
and U9668 (N_9668,N_6704,N_6001);
and U9669 (N_9669,N_7996,N_7422);
nand U9670 (N_9670,N_6742,N_6582);
nand U9671 (N_9671,N_6229,N_6697);
nor U9672 (N_9672,N_7543,N_6307);
and U9673 (N_9673,N_7693,N_6312);
nand U9674 (N_9674,N_7675,N_6349);
nor U9675 (N_9675,N_7478,N_6555);
nor U9676 (N_9676,N_7066,N_6840);
nor U9677 (N_9677,N_7336,N_6625);
and U9678 (N_9678,N_7374,N_7364);
nor U9679 (N_9679,N_7417,N_7078);
or U9680 (N_9680,N_6679,N_6267);
or U9681 (N_9681,N_6148,N_6226);
nand U9682 (N_9682,N_7275,N_6673);
and U9683 (N_9683,N_7968,N_6343);
nand U9684 (N_9684,N_7146,N_7339);
or U9685 (N_9685,N_6329,N_6497);
nor U9686 (N_9686,N_6744,N_6114);
and U9687 (N_9687,N_7434,N_6196);
nor U9688 (N_9688,N_6910,N_7632);
nor U9689 (N_9689,N_7267,N_6070);
nor U9690 (N_9690,N_7811,N_7726);
and U9691 (N_9691,N_7598,N_6184);
or U9692 (N_9692,N_7404,N_6121);
and U9693 (N_9693,N_7886,N_6841);
nor U9694 (N_9694,N_7433,N_6077);
and U9695 (N_9695,N_6098,N_6482);
xor U9696 (N_9696,N_6473,N_6854);
nand U9697 (N_9697,N_7045,N_6562);
nor U9698 (N_9698,N_6933,N_7958);
nand U9699 (N_9699,N_7823,N_6129);
nor U9700 (N_9700,N_6228,N_6777);
or U9701 (N_9701,N_6282,N_6522);
nand U9702 (N_9702,N_6640,N_6963);
nand U9703 (N_9703,N_7870,N_7302);
or U9704 (N_9704,N_6010,N_6081);
xor U9705 (N_9705,N_6041,N_6812);
nor U9706 (N_9706,N_7918,N_6270);
or U9707 (N_9707,N_6184,N_7702);
nand U9708 (N_9708,N_6223,N_6228);
nor U9709 (N_9709,N_7308,N_6327);
nor U9710 (N_9710,N_7996,N_7011);
nand U9711 (N_9711,N_6223,N_7920);
nor U9712 (N_9712,N_6163,N_6034);
and U9713 (N_9713,N_6752,N_6477);
or U9714 (N_9714,N_6855,N_7124);
nand U9715 (N_9715,N_6569,N_7737);
nor U9716 (N_9716,N_7012,N_6407);
nor U9717 (N_9717,N_7769,N_6750);
nor U9718 (N_9718,N_6952,N_6005);
and U9719 (N_9719,N_6643,N_7808);
nor U9720 (N_9720,N_6272,N_6259);
nand U9721 (N_9721,N_7705,N_7897);
nor U9722 (N_9722,N_6782,N_7745);
xnor U9723 (N_9723,N_6275,N_7108);
nand U9724 (N_9724,N_6763,N_7141);
or U9725 (N_9725,N_7686,N_7606);
and U9726 (N_9726,N_7348,N_7987);
nand U9727 (N_9727,N_7768,N_7681);
and U9728 (N_9728,N_7240,N_7770);
nand U9729 (N_9729,N_7506,N_7646);
xnor U9730 (N_9730,N_6390,N_6628);
nor U9731 (N_9731,N_7415,N_6917);
and U9732 (N_9732,N_6894,N_7365);
and U9733 (N_9733,N_6882,N_6854);
nand U9734 (N_9734,N_6086,N_6924);
or U9735 (N_9735,N_7453,N_6758);
and U9736 (N_9736,N_7038,N_6991);
nor U9737 (N_9737,N_6635,N_7727);
nand U9738 (N_9738,N_7839,N_7546);
xor U9739 (N_9739,N_6924,N_6478);
or U9740 (N_9740,N_7761,N_7241);
nor U9741 (N_9741,N_6667,N_7968);
and U9742 (N_9742,N_6875,N_6433);
nor U9743 (N_9743,N_7225,N_6437);
and U9744 (N_9744,N_6049,N_7703);
nor U9745 (N_9745,N_6387,N_6311);
nand U9746 (N_9746,N_7701,N_7640);
nand U9747 (N_9747,N_6999,N_7435);
or U9748 (N_9748,N_6938,N_6246);
nand U9749 (N_9749,N_6961,N_6056);
nand U9750 (N_9750,N_7571,N_7594);
and U9751 (N_9751,N_6139,N_7449);
and U9752 (N_9752,N_6548,N_6530);
nor U9753 (N_9753,N_7066,N_6317);
nor U9754 (N_9754,N_6016,N_6170);
or U9755 (N_9755,N_7548,N_7859);
and U9756 (N_9756,N_7217,N_6159);
and U9757 (N_9757,N_7042,N_6637);
nor U9758 (N_9758,N_7621,N_7060);
nand U9759 (N_9759,N_6467,N_6615);
and U9760 (N_9760,N_6902,N_7691);
nor U9761 (N_9761,N_7660,N_6913);
nand U9762 (N_9762,N_6102,N_7437);
nor U9763 (N_9763,N_7853,N_6996);
nand U9764 (N_9764,N_6447,N_6304);
or U9765 (N_9765,N_6061,N_6327);
and U9766 (N_9766,N_6405,N_7559);
and U9767 (N_9767,N_6274,N_6170);
or U9768 (N_9768,N_6440,N_6149);
or U9769 (N_9769,N_6731,N_7194);
and U9770 (N_9770,N_6191,N_6013);
and U9771 (N_9771,N_6461,N_7954);
and U9772 (N_9772,N_7901,N_6176);
nor U9773 (N_9773,N_6197,N_7955);
nand U9774 (N_9774,N_7278,N_6153);
or U9775 (N_9775,N_7302,N_6093);
and U9776 (N_9776,N_6298,N_7975);
or U9777 (N_9777,N_6455,N_6270);
nor U9778 (N_9778,N_7206,N_6035);
nand U9779 (N_9779,N_6207,N_6350);
or U9780 (N_9780,N_6799,N_7382);
and U9781 (N_9781,N_7298,N_7455);
or U9782 (N_9782,N_7789,N_6500);
nand U9783 (N_9783,N_7447,N_6661);
and U9784 (N_9784,N_6775,N_7104);
nor U9785 (N_9785,N_6434,N_6267);
or U9786 (N_9786,N_6471,N_7427);
nand U9787 (N_9787,N_7045,N_6782);
or U9788 (N_9788,N_7614,N_7814);
nor U9789 (N_9789,N_6904,N_6582);
nor U9790 (N_9790,N_6568,N_7721);
nor U9791 (N_9791,N_7950,N_6277);
and U9792 (N_9792,N_7204,N_6193);
nand U9793 (N_9793,N_7575,N_6408);
xor U9794 (N_9794,N_7056,N_6365);
and U9795 (N_9795,N_6755,N_6558);
or U9796 (N_9796,N_6622,N_7170);
or U9797 (N_9797,N_6328,N_7865);
nor U9798 (N_9798,N_6232,N_7184);
and U9799 (N_9799,N_7184,N_7074);
or U9800 (N_9800,N_7833,N_7487);
nand U9801 (N_9801,N_7217,N_7692);
or U9802 (N_9802,N_6601,N_6922);
nor U9803 (N_9803,N_7602,N_7899);
xnor U9804 (N_9804,N_7311,N_7172);
nand U9805 (N_9805,N_7602,N_6417);
xnor U9806 (N_9806,N_7674,N_6782);
and U9807 (N_9807,N_6842,N_7715);
or U9808 (N_9808,N_7813,N_6673);
or U9809 (N_9809,N_6333,N_6172);
or U9810 (N_9810,N_7811,N_6773);
or U9811 (N_9811,N_6689,N_7500);
nand U9812 (N_9812,N_6553,N_6472);
nor U9813 (N_9813,N_6051,N_6758);
or U9814 (N_9814,N_6575,N_7476);
xor U9815 (N_9815,N_7607,N_7681);
nor U9816 (N_9816,N_7112,N_6179);
and U9817 (N_9817,N_7981,N_7324);
and U9818 (N_9818,N_6340,N_7446);
xor U9819 (N_9819,N_7530,N_7129);
or U9820 (N_9820,N_7162,N_6581);
nor U9821 (N_9821,N_6970,N_6908);
and U9822 (N_9822,N_6937,N_7506);
nand U9823 (N_9823,N_6426,N_7076);
or U9824 (N_9824,N_7550,N_6034);
or U9825 (N_9825,N_6568,N_6685);
or U9826 (N_9826,N_7529,N_7616);
nand U9827 (N_9827,N_6624,N_7434);
nand U9828 (N_9828,N_7187,N_7386);
and U9829 (N_9829,N_6088,N_6671);
nor U9830 (N_9830,N_7084,N_7585);
xnor U9831 (N_9831,N_7218,N_6585);
nand U9832 (N_9832,N_6245,N_7258);
or U9833 (N_9833,N_7235,N_6642);
nor U9834 (N_9834,N_6682,N_6085);
nand U9835 (N_9835,N_7788,N_6926);
and U9836 (N_9836,N_6747,N_6720);
and U9837 (N_9837,N_7532,N_6062);
or U9838 (N_9838,N_7448,N_7920);
nor U9839 (N_9839,N_7276,N_7144);
or U9840 (N_9840,N_7021,N_6628);
nand U9841 (N_9841,N_6081,N_7071);
nor U9842 (N_9842,N_6312,N_6214);
nand U9843 (N_9843,N_6951,N_7776);
nand U9844 (N_9844,N_7698,N_6431);
nor U9845 (N_9845,N_6382,N_6889);
and U9846 (N_9846,N_6630,N_6168);
and U9847 (N_9847,N_6658,N_7856);
nand U9848 (N_9848,N_6603,N_7693);
and U9849 (N_9849,N_7596,N_7912);
and U9850 (N_9850,N_7435,N_6953);
or U9851 (N_9851,N_6429,N_7382);
and U9852 (N_9852,N_7491,N_7252);
nor U9853 (N_9853,N_7756,N_6820);
nand U9854 (N_9854,N_7138,N_6641);
nor U9855 (N_9855,N_6376,N_6540);
nor U9856 (N_9856,N_6143,N_7663);
or U9857 (N_9857,N_6993,N_6014);
nand U9858 (N_9858,N_7154,N_6092);
and U9859 (N_9859,N_6103,N_6559);
and U9860 (N_9860,N_7608,N_7669);
nor U9861 (N_9861,N_6183,N_6094);
nor U9862 (N_9862,N_6344,N_6299);
and U9863 (N_9863,N_6517,N_7824);
or U9864 (N_9864,N_6942,N_7444);
and U9865 (N_9865,N_7470,N_7115);
and U9866 (N_9866,N_7100,N_6162);
and U9867 (N_9867,N_6943,N_7456);
nor U9868 (N_9868,N_6481,N_6525);
or U9869 (N_9869,N_7521,N_7947);
nor U9870 (N_9870,N_6581,N_6371);
nor U9871 (N_9871,N_7991,N_6823);
or U9872 (N_9872,N_7425,N_7808);
nor U9873 (N_9873,N_7427,N_7920);
or U9874 (N_9874,N_7040,N_6579);
or U9875 (N_9875,N_6038,N_7042);
and U9876 (N_9876,N_7098,N_7212);
nor U9877 (N_9877,N_7889,N_6032);
or U9878 (N_9878,N_7056,N_6420);
nor U9879 (N_9879,N_6978,N_7802);
or U9880 (N_9880,N_7546,N_6363);
nor U9881 (N_9881,N_6333,N_7765);
nor U9882 (N_9882,N_7189,N_6138);
nand U9883 (N_9883,N_7063,N_6124);
or U9884 (N_9884,N_6358,N_7352);
xor U9885 (N_9885,N_7052,N_7886);
xor U9886 (N_9886,N_7274,N_7624);
and U9887 (N_9887,N_7752,N_7637);
and U9888 (N_9888,N_6897,N_6240);
nor U9889 (N_9889,N_6415,N_7642);
and U9890 (N_9890,N_6606,N_6450);
or U9891 (N_9891,N_7840,N_7519);
or U9892 (N_9892,N_7219,N_7025);
or U9893 (N_9893,N_6487,N_7609);
nor U9894 (N_9894,N_7732,N_6529);
nand U9895 (N_9895,N_7214,N_6122);
and U9896 (N_9896,N_7327,N_6359);
xnor U9897 (N_9897,N_6812,N_7138);
or U9898 (N_9898,N_6656,N_7757);
or U9899 (N_9899,N_6537,N_7228);
or U9900 (N_9900,N_6879,N_7912);
or U9901 (N_9901,N_6889,N_6412);
and U9902 (N_9902,N_6818,N_6106);
or U9903 (N_9903,N_6619,N_7089);
and U9904 (N_9904,N_7225,N_7933);
or U9905 (N_9905,N_6108,N_6209);
nor U9906 (N_9906,N_6950,N_6191);
and U9907 (N_9907,N_6369,N_7721);
or U9908 (N_9908,N_7501,N_6641);
nor U9909 (N_9909,N_7785,N_6034);
and U9910 (N_9910,N_7721,N_6335);
nor U9911 (N_9911,N_6977,N_6784);
and U9912 (N_9912,N_6248,N_6206);
nor U9913 (N_9913,N_6306,N_6277);
and U9914 (N_9914,N_6649,N_6053);
or U9915 (N_9915,N_6801,N_6121);
nor U9916 (N_9916,N_7855,N_6939);
nor U9917 (N_9917,N_6730,N_6084);
nor U9918 (N_9918,N_6605,N_6739);
and U9919 (N_9919,N_7182,N_6105);
or U9920 (N_9920,N_6358,N_7101);
nor U9921 (N_9921,N_6100,N_6163);
nor U9922 (N_9922,N_6315,N_7904);
or U9923 (N_9923,N_6584,N_6592);
or U9924 (N_9924,N_7500,N_6419);
or U9925 (N_9925,N_6435,N_6832);
nand U9926 (N_9926,N_7493,N_7442);
nor U9927 (N_9927,N_7659,N_7843);
or U9928 (N_9928,N_7728,N_7264);
nand U9929 (N_9929,N_7455,N_6909);
and U9930 (N_9930,N_7793,N_7825);
and U9931 (N_9931,N_6577,N_7292);
nor U9932 (N_9932,N_6135,N_6909);
nor U9933 (N_9933,N_6505,N_6990);
or U9934 (N_9934,N_7519,N_7311);
xor U9935 (N_9935,N_7516,N_6970);
and U9936 (N_9936,N_6292,N_6581);
nand U9937 (N_9937,N_6604,N_7351);
or U9938 (N_9938,N_6174,N_7267);
and U9939 (N_9939,N_7302,N_7115);
nor U9940 (N_9940,N_7291,N_6002);
nand U9941 (N_9941,N_7028,N_7114);
nor U9942 (N_9942,N_6480,N_7060);
nand U9943 (N_9943,N_6673,N_7210);
xnor U9944 (N_9944,N_7971,N_7735);
nor U9945 (N_9945,N_6856,N_7790);
and U9946 (N_9946,N_6904,N_6995);
and U9947 (N_9947,N_6710,N_7453);
or U9948 (N_9948,N_7659,N_6032);
or U9949 (N_9949,N_7899,N_7704);
or U9950 (N_9950,N_7134,N_7421);
or U9951 (N_9951,N_6335,N_7518);
or U9952 (N_9952,N_6202,N_6904);
or U9953 (N_9953,N_6667,N_7031);
or U9954 (N_9954,N_6016,N_7637);
or U9955 (N_9955,N_7642,N_7999);
or U9956 (N_9956,N_6297,N_6496);
and U9957 (N_9957,N_6806,N_7082);
or U9958 (N_9958,N_7726,N_6797);
or U9959 (N_9959,N_6974,N_6670);
or U9960 (N_9960,N_6933,N_6323);
nand U9961 (N_9961,N_6836,N_7307);
and U9962 (N_9962,N_7140,N_6261);
nand U9963 (N_9963,N_7427,N_7474);
or U9964 (N_9964,N_6642,N_7323);
or U9965 (N_9965,N_7595,N_7895);
nand U9966 (N_9966,N_6283,N_7980);
and U9967 (N_9967,N_7542,N_6209);
and U9968 (N_9968,N_6676,N_7444);
and U9969 (N_9969,N_6638,N_6789);
and U9970 (N_9970,N_6668,N_6533);
or U9971 (N_9971,N_7066,N_6206);
and U9972 (N_9972,N_7940,N_7682);
or U9973 (N_9973,N_6780,N_7311);
nand U9974 (N_9974,N_7075,N_6167);
nor U9975 (N_9975,N_7959,N_7794);
nor U9976 (N_9976,N_6365,N_6692);
nor U9977 (N_9977,N_7640,N_6231);
nor U9978 (N_9978,N_6968,N_6545);
or U9979 (N_9979,N_6816,N_7167);
and U9980 (N_9980,N_6679,N_6268);
nor U9981 (N_9981,N_6146,N_6540);
or U9982 (N_9982,N_7359,N_6081);
nor U9983 (N_9983,N_7488,N_6288);
and U9984 (N_9984,N_6614,N_6529);
or U9985 (N_9985,N_6209,N_7897);
nand U9986 (N_9986,N_6450,N_7593);
nor U9987 (N_9987,N_6189,N_7224);
nand U9988 (N_9988,N_6303,N_7963);
nand U9989 (N_9989,N_7399,N_7396);
nor U9990 (N_9990,N_6600,N_7304);
nor U9991 (N_9991,N_6119,N_6105);
and U9992 (N_9992,N_6502,N_6827);
nand U9993 (N_9993,N_7164,N_6467);
nor U9994 (N_9994,N_7252,N_7945);
and U9995 (N_9995,N_6910,N_7150);
and U9996 (N_9996,N_7214,N_7192);
xor U9997 (N_9997,N_7808,N_7743);
nor U9998 (N_9998,N_7823,N_6861);
or U9999 (N_9999,N_7943,N_6617);
nor UO_0 (O_0,N_8350,N_9835);
nand UO_1 (O_1,N_8582,N_8965);
and UO_2 (O_2,N_9787,N_8378);
nand UO_3 (O_3,N_9903,N_9964);
nand UO_4 (O_4,N_8995,N_8941);
or UO_5 (O_5,N_9064,N_8442);
nand UO_6 (O_6,N_9797,N_8414);
and UO_7 (O_7,N_8118,N_8905);
and UO_8 (O_8,N_8474,N_8654);
nor UO_9 (O_9,N_8263,N_8741);
or UO_10 (O_10,N_8675,N_8178);
nor UO_11 (O_11,N_9949,N_9522);
or UO_12 (O_12,N_8503,N_9307);
nand UO_13 (O_13,N_9709,N_8469);
or UO_14 (O_14,N_9326,N_8816);
nand UO_15 (O_15,N_8725,N_8008);
and UO_16 (O_16,N_9673,N_8598);
nand UO_17 (O_17,N_9228,N_9707);
and UO_18 (O_18,N_9267,N_8628);
nand UO_19 (O_19,N_9285,N_9985);
and UO_20 (O_20,N_8748,N_8964);
nand UO_21 (O_21,N_8116,N_9584);
and UO_22 (O_22,N_8298,N_8190);
nor UO_23 (O_23,N_9593,N_9183);
or UO_24 (O_24,N_9448,N_9234);
nor UO_25 (O_25,N_9099,N_9209);
nor UO_26 (O_26,N_9864,N_8092);
and UO_27 (O_27,N_8493,N_9640);
or UO_28 (O_28,N_9339,N_9194);
nand UO_29 (O_29,N_8956,N_9116);
nor UO_30 (O_30,N_8841,N_8291);
nor UO_31 (O_31,N_8904,N_9679);
nand UO_32 (O_32,N_8030,N_9033);
nor UO_33 (O_33,N_8184,N_9669);
nor UO_34 (O_34,N_9893,N_8988);
nand UO_35 (O_35,N_8089,N_9443);
xor UO_36 (O_36,N_9541,N_8990);
nor UO_37 (O_37,N_9352,N_8659);
or UO_38 (O_38,N_9534,N_8874);
nand UO_39 (O_39,N_8785,N_9906);
nand UO_40 (O_40,N_8788,N_9966);
nor UO_41 (O_41,N_8061,N_9042);
nor UO_42 (O_42,N_9856,N_9999);
and UO_43 (O_43,N_8633,N_8399);
or UO_44 (O_44,N_9926,N_9716);
and UO_45 (O_45,N_8819,N_9970);
nand UO_46 (O_46,N_8739,N_9508);
nor UO_47 (O_47,N_9585,N_8865);
nor UO_48 (O_48,N_9426,N_8609);
or UO_49 (O_49,N_9420,N_8193);
nand UO_50 (O_50,N_9582,N_9745);
nand UO_51 (O_51,N_9989,N_9629);
nand UO_52 (O_52,N_9177,N_9337);
or UO_53 (O_53,N_9325,N_9370);
xor UO_54 (O_54,N_8219,N_9625);
nor UO_55 (O_55,N_9773,N_8637);
and UO_56 (O_56,N_8806,N_8880);
nor UO_57 (O_57,N_9273,N_9134);
nor UO_58 (O_58,N_9184,N_8954);
and UO_59 (O_59,N_9176,N_9768);
or UO_60 (O_60,N_8171,N_8370);
and UO_61 (O_61,N_9609,N_8820);
nand UO_62 (O_62,N_8516,N_8967);
or UO_63 (O_63,N_9652,N_8685);
nor UO_64 (O_64,N_8472,N_9857);
nand UO_65 (O_65,N_8492,N_8374);
nand UO_66 (O_66,N_8159,N_8925);
nor UO_67 (O_67,N_8071,N_9535);
and UO_68 (O_68,N_9061,N_8188);
nand UO_69 (O_69,N_9761,N_8680);
nand UO_70 (O_70,N_9688,N_9168);
or UO_71 (O_71,N_8626,N_8405);
or UO_72 (O_72,N_9904,N_8424);
or UO_73 (O_73,N_8362,N_9675);
or UO_74 (O_74,N_8120,N_8556);
and UO_75 (O_75,N_8643,N_9065);
nor UO_76 (O_76,N_8569,N_9023);
nor UO_77 (O_77,N_9715,N_8936);
and UO_78 (O_78,N_9338,N_9586);
nand UO_79 (O_79,N_8307,N_8288);
nand UO_80 (O_80,N_8194,N_9252);
nand UO_81 (O_81,N_9552,N_9263);
and UO_82 (O_82,N_8529,N_8349);
or UO_83 (O_83,N_8638,N_9705);
or UO_84 (O_84,N_9692,N_8890);
nand UO_85 (O_85,N_9427,N_8133);
nor UO_86 (O_86,N_8713,N_9548);
nor UO_87 (O_87,N_8729,N_8804);
nand UO_88 (O_88,N_8999,N_8044);
nor UO_89 (O_89,N_9386,N_8496);
xnor UO_90 (O_90,N_9305,N_8220);
or UO_91 (O_91,N_9462,N_9380);
nor UO_92 (O_92,N_8100,N_8153);
nor UO_93 (O_93,N_9026,N_9980);
nand UO_94 (O_94,N_8591,N_9332);
or UO_95 (O_95,N_9765,N_9001);
nand UO_96 (O_96,N_9555,N_9727);
and UO_97 (O_97,N_9588,N_9400);
or UO_98 (O_98,N_8286,N_8982);
nor UO_99 (O_99,N_9938,N_8302);
nor UO_100 (O_100,N_8850,N_8580);
nand UO_101 (O_101,N_9284,N_9862);
nor UO_102 (O_102,N_9217,N_9747);
nor UO_103 (O_103,N_8687,N_9054);
or UO_104 (O_104,N_9934,N_9786);
and UO_105 (O_105,N_8005,N_9892);
nand UO_106 (O_106,N_9068,N_8952);
or UO_107 (O_107,N_9082,N_9684);
or UO_108 (O_108,N_9847,N_8473);
and UO_109 (O_109,N_9936,N_9073);
nor UO_110 (O_110,N_9411,N_8028);
or UO_111 (O_111,N_9930,N_9324);
xnor UO_112 (O_112,N_9662,N_9471);
nor UO_113 (O_113,N_9363,N_8484);
nand UO_114 (O_114,N_8674,N_8355);
or UO_115 (O_115,N_9851,N_8660);
and UO_116 (O_116,N_8119,N_8105);
or UO_117 (O_117,N_8782,N_9683);
nand UO_118 (O_118,N_9240,N_8017);
nor UO_119 (O_119,N_8131,N_8397);
nand UO_120 (O_120,N_9371,N_8199);
nor UO_121 (O_121,N_8755,N_8331);
nand UO_122 (O_122,N_8146,N_8692);
and UO_123 (O_123,N_9170,N_8267);
nor UO_124 (O_124,N_9825,N_9416);
nand UO_125 (O_125,N_9923,N_8848);
and UO_126 (O_126,N_9405,N_9458);
or UO_127 (O_127,N_8210,N_9137);
and UO_128 (O_128,N_9150,N_8610);
or UO_129 (O_129,N_8588,N_9104);
nand UO_130 (O_130,N_9476,N_8024);
nand UO_131 (O_131,N_8336,N_8137);
and UO_132 (O_132,N_8832,N_9986);
and UO_133 (O_133,N_9464,N_8018);
and UO_134 (O_134,N_9900,N_9699);
and UO_135 (O_135,N_9646,N_9084);
or UO_136 (O_136,N_9293,N_9823);
nor UO_137 (O_137,N_8415,N_9800);
and UO_138 (O_138,N_9093,N_8651);
nand UO_139 (O_139,N_8808,N_8549);
or UO_140 (O_140,N_8517,N_9838);
and UO_141 (O_141,N_9556,N_8553);
or UO_142 (O_142,N_8753,N_8047);
nor UO_143 (O_143,N_8666,N_8619);
nand UO_144 (O_144,N_8854,N_9627);
or UO_145 (O_145,N_8211,N_8106);
or UO_146 (O_146,N_8984,N_8132);
nor UO_147 (O_147,N_9025,N_9869);
or UO_148 (O_148,N_8949,N_9622);
nand UO_149 (O_149,N_8677,N_9329);
nor UO_150 (O_150,N_8974,N_9497);
or UO_151 (O_151,N_8770,N_9811);
nor UO_152 (O_152,N_9051,N_8101);
nand UO_153 (O_153,N_9706,N_8640);
and UO_154 (O_154,N_8877,N_9179);
or UO_155 (O_155,N_8515,N_9136);
nand UO_156 (O_156,N_8090,N_8143);
and UO_157 (O_157,N_9920,N_8987);
and UO_158 (O_158,N_8420,N_9603);
nor UO_159 (O_159,N_8325,N_9839);
nor UO_160 (O_160,N_8766,N_9613);
or UO_161 (O_161,N_8879,N_8324);
xnor UO_162 (O_162,N_8707,N_8292);
nand UO_163 (O_163,N_9660,N_9830);
nand UO_164 (O_164,N_8720,N_8617);
nand UO_165 (O_165,N_8125,N_8130);
or UO_166 (O_166,N_8096,N_9347);
or UO_167 (O_167,N_8606,N_9218);
or UO_168 (O_168,N_8466,N_9384);
nor UO_169 (O_169,N_9100,N_9083);
nand UO_170 (O_170,N_8903,N_8479);
or UO_171 (O_171,N_9124,N_8306);
or UO_172 (O_172,N_9062,N_8966);
or UO_173 (O_173,N_9712,N_8909);
or UO_174 (O_174,N_8215,N_9265);
and UO_175 (O_175,N_9475,N_8142);
nand UO_176 (O_176,N_8695,N_9882);
and UO_177 (O_177,N_9597,N_9049);
nand UO_178 (O_178,N_9147,N_9560);
and UO_179 (O_179,N_8597,N_8311);
nor UO_180 (O_180,N_9867,N_9279);
xnor UO_181 (O_181,N_9000,N_9089);
nand UO_182 (O_182,N_9860,N_8250);
xor UO_183 (O_183,N_9578,N_8551);
xor UO_184 (O_184,N_9395,N_8803);
nor UO_185 (O_185,N_8682,N_8570);
nor UO_186 (O_186,N_8076,N_9342);
or UO_187 (O_187,N_8161,N_9200);
nand UO_188 (O_188,N_8321,N_8351);
and UO_189 (O_189,N_9212,N_8165);
nor UO_190 (O_190,N_9636,N_8462);
nand UO_191 (O_191,N_8391,N_8658);
nand UO_192 (O_192,N_8299,N_9898);
nand UO_193 (O_193,N_8392,N_9780);
or UO_194 (O_194,N_9658,N_8022);
and UO_195 (O_195,N_9292,N_8846);
and UO_196 (O_196,N_9301,N_8227);
and UO_197 (O_197,N_8140,N_9998);
and UO_198 (O_198,N_9071,N_8077);
nor UO_199 (O_199,N_9872,N_8475);
and UO_200 (O_200,N_9058,N_9808);
and UO_201 (O_201,N_8151,N_9929);
or UO_202 (O_202,N_9160,N_8947);
and UO_203 (O_203,N_8272,N_8114);
nand UO_204 (O_204,N_8775,N_8585);
or UO_205 (O_205,N_9059,N_8656);
and UO_206 (O_206,N_8412,N_8274);
or UO_207 (O_207,N_8579,N_9897);
or UO_208 (O_208,N_9852,N_8858);
nand UO_209 (O_209,N_9782,N_9630);
or UO_210 (O_210,N_8812,N_9511);
and UO_211 (O_211,N_8972,N_8786);
nor UO_212 (O_212,N_8430,N_8704);
and UO_213 (O_213,N_9742,N_9169);
nand UO_214 (O_214,N_9086,N_8700);
nand UO_215 (O_215,N_9583,N_8086);
nor UO_216 (O_216,N_8026,N_8636);
or UO_217 (O_217,N_8754,N_8231);
nand UO_218 (O_218,N_9608,N_8544);
nor UO_219 (O_219,N_8814,N_8867);
or UO_220 (O_220,N_9121,N_8110);
xnor UO_221 (O_221,N_9990,N_9264);
nor UO_222 (O_222,N_9087,N_8724);
nor UO_223 (O_223,N_9385,N_9971);
nand UO_224 (O_224,N_9317,N_9878);
or UO_225 (O_225,N_9663,N_8236);
nor UO_226 (O_226,N_8507,N_9070);
nand UO_227 (O_227,N_8940,N_8962);
nor UO_228 (O_228,N_8975,N_8917);
nand UO_229 (O_229,N_8148,N_8094);
or UO_230 (O_230,N_9127,N_9047);
and UO_231 (O_231,N_9820,N_9312);
or UO_232 (O_232,N_9912,N_9398);
and UO_233 (O_233,N_9817,N_8514);
nor UO_234 (O_234,N_8872,N_8357);
or UO_235 (O_235,N_8064,N_9557);
or UO_236 (O_236,N_9007,N_9422);
nor UO_237 (O_237,N_9291,N_8627);
nor UO_238 (O_238,N_9813,N_9554);
nand UO_239 (O_239,N_8287,N_8543);
or UO_240 (O_240,N_9965,N_8953);
nor UO_241 (O_241,N_8657,N_8891);
or UO_242 (O_242,N_8407,N_9055);
or UO_243 (O_243,N_9710,N_9972);
or UO_244 (O_244,N_9197,N_9784);
and UO_245 (O_245,N_8310,N_9014);
nand UO_246 (O_246,N_9298,N_8482);
nand UO_247 (O_247,N_9592,N_8584);
and UO_248 (O_248,N_9114,N_9199);
and UO_249 (O_249,N_9655,N_8678);
and UO_250 (O_250,N_8300,N_8383);
nand UO_251 (O_251,N_8871,N_9802);
or UO_252 (O_252,N_8513,N_9547);
nor UO_253 (O_253,N_9175,N_9902);
nand UO_254 (O_254,N_8526,N_8422);
or UO_255 (O_255,N_8634,N_8266);
nand UO_256 (O_256,N_9503,N_9565);
nor UO_257 (O_257,N_8552,N_8013);
xor UO_258 (O_258,N_9696,N_9632);
or UO_259 (O_259,N_8981,N_8670);
nand UO_260 (O_260,N_8779,N_8115);
nand UO_261 (O_261,N_9732,N_9163);
or UO_262 (O_262,N_9573,N_9571);
or UO_263 (O_263,N_8075,N_9079);
or UO_264 (O_264,N_8326,N_9506);
or UO_265 (O_265,N_9446,N_8837);
and UO_266 (O_266,N_8452,N_8445);
or UO_267 (O_267,N_8260,N_8817);
and UO_268 (O_268,N_8168,N_8180);
or UO_269 (O_269,N_8856,N_9360);
or UO_270 (O_270,N_9246,N_9726);
or UO_271 (O_271,N_8453,N_9138);
or UO_272 (O_272,N_8979,N_9602);
and UO_273 (O_273,N_9203,N_8058);
and UO_274 (O_274,N_9479,N_9181);
nor UO_275 (O_275,N_8961,N_9762);
nor UO_276 (O_276,N_9243,N_8581);
and UO_277 (O_277,N_9048,N_9204);
nor UO_278 (O_278,N_8328,N_9271);
or UO_279 (O_279,N_8530,N_9610);
nand UO_280 (O_280,N_8170,N_8971);
and UO_281 (O_281,N_9656,N_9978);
nor UO_282 (O_282,N_9392,N_9502);
or UO_283 (O_283,N_9453,N_8041);
or UO_284 (O_284,N_8270,N_8358);
and UO_285 (O_285,N_8200,N_8093);
nand UO_286 (O_286,N_9946,N_8135);
or UO_287 (O_287,N_8278,N_9076);
and UO_288 (O_288,N_8986,N_8344);
nor UO_289 (O_289,N_8489,N_9269);
or UO_290 (O_290,N_8611,N_9222);
xnor UO_291 (O_291,N_8346,N_9957);
and UO_292 (O_292,N_8485,N_9477);
nor UO_293 (O_293,N_9935,N_9533);
and UO_294 (O_294,N_8379,N_9235);
nand UO_295 (O_295,N_9031,N_8341);
nor UO_296 (O_296,N_8511,N_8107);
and UO_297 (O_297,N_8059,N_9117);
and UO_298 (O_298,N_9532,N_9909);
and UO_299 (O_299,N_8538,N_8122);
and UO_300 (O_300,N_9649,N_9377);
nand UO_301 (O_301,N_9249,N_8365);
or UO_302 (O_302,N_8461,N_9341);
nor UO_303 (O_303,N_9539,N_8589);
nor UO_304 (O_304,N_8767,N_9146);
and UO_305 (O_305,N_9956,N_9159);
or UO_306 (O_306,N_8918,N_8304);
nand UO_307 (O_307,N_9974,N_9188);
nor UO_308 (O_308,N_8467,N_8983);
xor UO_309 (O_309,N_8312,N_9135);
nor UO_310 (O_310,N_8934,N_8446);
and UO_311 (O_311,N_9225,N_9361);
and UO_312 (O_312,N_8884,N_9939);
and UO_313 (O_313,N_8062,N_8175);
nor UO_314 (O_314,N_9517,N_8053);
or UO_315 (O_315,N_8727,N_8388);
or UO_316 (O_316,N_8376,N_9202);
and UO_317 (O_317,N_8883,N_9733);
nor UO_318 (O_318,N_8046,N_9091);
or UO_319 (O_319,N_9098,N_9343);
and UO_320 (O_320,N_8969,N_9242);
nand UO_321 (O_321,N_9155,N_9357);
nor UO_322 (O_322,N_8242,N_9703);
or UO_323 (O_323,N_8875,N_8978);
nor UO_324 (O_324,N_8932,N_9685);
and UO_325 (O_325,N_9429,N_9485);
or UO_326 (O_326,N_9858,N_9090);
nand UO_327 (O_327,N_8016,N_9460);
nor UO_328 (O_328,N_9807,N_8989);
nor UO_329 (O_329,N_8946,N_8333);
nand UO_330 (O_330,N_8916,N_9589);
or UO_331 (O_331,N_8547,N_8824);
and UO_332 (O_332,N_9987,N_9433);
nand UO_333 (O_333,N_8523,N_9101);
nor UO_334 (O_334,N_8000,N_9372);
and UO_335 (O_335,N_8012,N_8778);
or UO_336 (O_336,N_9689,N_9111);
and UO_337 (O_337,N_8620,N_8011);
or UO_338 (O_338,N_9428,N_8691);
nor UO_339 (O_339,N_8531,N_8718);
nand UO_340 (O_340,N_9748,N_8679);
or UO_341 (O_341,N_8323,N_9650);
and UO_342 (O_342,N_9538,N_9468);
nand UO_343 (O_343,N_8839,N_8253);
nand UO_344 (O_344,N_8542,N_9907);
or UO_345 (O_345,N_8400,N_9319);
and UO_346 (O_346,N_9483,N_8512);
nor UO_347 (O_347,N_8758,N_9013);
or UO_348 (O_348,N_8738,N_9604);
and UO_349 (O_349,N_8191,N_9948);
xnor UO_350 (O_350,N_9621,N_9018);
xnor UO_351 (O_351,N_8375,N_8010);
or UO_352 (O_352,N_9407,N_9382);
or UO_353 (O_353,N_8676,N_9299);
nor UO_354 (O_354,N_8750,N_8160);
nor UO_355 (O_355,N_9691,N_9296);
nand UO_356 (O_356,N_8404,N_9873);
and UO_357 (O_357,N_8082,N_9178);
and UO_358 (O_358,N_8719,N_8443);
nand UO_359 (O_359,N_9596,N_9527);
xor UO_360 (O_360,N_9828,N_9172);
and UO_361 (O_361,N_9558,N_9043);
or UO_362 (O_362,N_8481,N_8237);
nand UO_363 (O_363,N_8863,N_8744);
and UO_364 (O_364,N_8829,N_9067);
and UO_365 (O_365,N_8478,N_8280);
and UO_366 (O_366,N_8394,N_9697);
and UO_367 (O_367,N_9313,N_8124);
and UO_368 (O_368,N_9180,N_8888);
nor UO_369 (O_369,N_8217,N_9066);
nor UO_370 (O_370,N_8463,N_8623);
nor UO_371 (O_371,N_8761,N_8483);
or UO_372 (O_372,N_8795,N_8600);
and UO_373 (O_373,N_8590,N_9525);
and UO_374 (O_374,N_9886,N_9568);
nor UO_375 (O_375,N_9566,N_9327);
and UO_376 (O_376,N_8545,N_9600);
and UO_377 (O_377,N_8866,N_8395);
nor UO_378 (O_378,N_9102,N_9676);
or UO_379 (O_379,N_9053,N_9801);
or UO_380 (O_380,N_8639,N_9781);
or UO_381 (O_381,N_9431,N_9275);
or UO_382 (O_382,N_8337,N_8246);
or UO_383 (O_383,N_8743,N_8223);
and UO_384 (O_384,N_8403,N_9766);
or UO_385 (O_385,N_9754,N_8487);
or UO_386 (O_386,N_8799,N_8275);
or UO_387 (O_387,N_9257,N_8693);
or UO_388 (O_388,N_8285,N_8413);
and UO_389 (O_389,N_9729,N_8838);
nor UO_390 (O_390,N_8360,N_9481);
or UO_391 (O_391,N_9606,N_9919);
and UO_392 (O_392,N_9221,N_8586);
or UO_393 (O_393,N_8813,N_8732);
or UO_394 (O_394,N_9010,N_9598);
and UO_395 (O_395,N_8836,N_9931);
and UO_396 (O_396,N_9736,N_9916);
and UO_397 (O_397,N_9115,N_8189);
or UO_398 (O_398,N_9303,N_9859);
and UO_399 (O_399,N_8673,N_8497);
nand UO_400 (O_400,N_9278,N_9545);
and UO_401 (O_401,N_9799,N_9414);
and UO_402 (O_402,N_9666,N_9328);
nand UO_403 (O_403,N_9616,N_9383);
and UO_404 (O_404,N_9871,N_8894);
and UO_405 (O_405,N_9247,N_9988);
nand UO_406 (O_406,N_9186,N_8613);
nor UO_407 (O_407,N_8709,N_9868);
or UO_408 (O_408,N_9861,N_8476);
nor UO_409 (O_409,N_8282,N_8038);
nand UO_410 (O_410,N_8243,N_9148);
nand UO_411 (O_411,N_8575,N_9196);
nor UO_412 (O_412,N_9977,N_8083);
or UO_413 (O_413,N_9157,N_8330);
or UO_414 (O_414,N_8396,N_8776);
and UO_415 (O_415,N_9962,N_9624);
nor UO_416 (O_416,N_9394,N_9698);
or UO_417 (O_417,N_8235,N_9671);
nor UO_418 (O_418,N_8334,N_8652);
or UO_419 (O_419,N_8759,N_9848);
and UO_420 (O_420,N_9816,N_8923);
nand UO_421 (O_421,N_8491,N_9495);
and UO_422 (O_422,N_9192,N_9693);
nand UO_423 (O_423,N_9145,N_8248);
nor UO_424 (O_424,N_9826,N_8035);
nor UO_425 (O_425,N_8958,N_8921);
nor UO_426 (O_426,N_8714,N_8845);
or UO_427 (O_427,N_9306,N_8056);
or UO_428 (O_428,N_9272,N_8807);
or UO_429 (O_429,N_8134,N_8710);
or UO_430 (O_430,N_8810,N_8342);
nand UO_431 (O_431,N_9760,N_9277);
or UO_432 (O_432,N_9143,N_8157);
and UO_433 (O_433,N_8162,N_8173);
xnor UO_434 (O_434,N_9152,N_8631);
or UO_435 (O_435,N_8825,N_8564);
nor UO_436 (O_436,N_8149,N_9419);
nor UO_437 (O_437,N_9953,N_9144);
nand UO_438 (O_438,N_9261,N_8212);
nor UO_439 (O_439,N_9519,N_8070);
nand UO_440 (O_440,N_8668,N_9738);
nand UO_441 (O_441,N_9330,N_8749);
nand UO_442 (O_442,N_8960,N_9772);
and UO_443 (O_443,N_9375,N_9810);
and UO_444 (O_444,N_8169,N_9258);
or UO_445 (O_445,N_9833,N_8976);
and UO_446 (O_446,N_9913,N_9300);
and UO_447 (O_447,N_8258,N_9028);
and UO_448 (O_448,N_8835,N_8108);
nand UO_449 (O_449,N_8733,N_8554);
nor UO_450 (O_450,N_9499,N_9425);
or UO_451 (O_451,N_8464,N_8632);
nor UO_452 (O_452,N_8273,N_9259);
nor UO_453 (O_453,N_8920,N_9173);
or UO_454 (O_454,N_9465,N_8889);
and UO_455 (O_455,N_9256,N_9129);
nor UO_456 (O_456,N_9110,N_8811);
or UO_457 (O_457,N_9737,N_8508);
and UO_458 (O_458,N_8645,N_9132);
and UO_459 (O_459,N_9036,N_9286);
and UO_460 (O_460,N_8208,N_9198);
nor UO_461 (O_461,N_8686,N_9647);
and UO_462 (O_462,N_9992,N_8821);
nand UO_463 (O_463,N_8195,N_9351);
xor UO_464 (O_464,N_8801,N_8045);
nor UO_465 (O_465,N_8906,N_9415);
nand UO_466 (O_466,N_9954,N_9947);
nor UO_467 (O_467,N_9943,N_9870);
nand UO_468 (O_468,N_8356,N_8295);
or UO_469 (O_469,N_9982,N_9883);
or UO_470 (O_470,N_9409,N_8773);
and UO_471 (O_471,N_9829,N_8241);
nor UO_472 (O_472,N_8103,N_8926);
or UO_473 (O_473,N_8897,N_8706);
nand UO_474 (O_474,N_8648,N_9501);
nor UO_475 (O_475,N_8655,N_9680);
or UO_476 (O_476,N_9167,N_9876);
or UO_477 (O_477,N_8091,N_8723);
and UO_478 (O_478,N_9678,N_9165);
or UO_479 (O_479,N_9027,N_8283);
nand UO_480 (O_480,N_8158,N_8389);
nor UO_481 (O_481,N_9412,N_8572);
nand UO_482 (O_482,N_8931,N_8339);
nor UO_483 (O_483,N_9855,N_9777);
nand UO_484 (O_484,N_9030,N_8762);
and UO_485 (O_485,N_9791,N_8576);
nor UO_486 (O_486,N_9454,N_9491);
nand UO_487 (O_487,N_9182,N_9940);
and UO_488 (O_488,N_9320,N_9997);
nand UO_489 (O_489,N_8329,N_9390);
nor UO_490 (O_490,N_9498,N_9723);
or UO_491 (O_491,N_9365,N_8138);
and UO_492 (O_492,N_9623,N_9518);
and UO_493 (O_493,N_9374,N_9576);
and UO_494 (O_494,N_9120,N_8247);
and UO_495 (O_495,N_9174,N_9232);
nand UO_496 (O_496,N_9887,N_9309);
nor UO_497 (O_497,N_9759,N_8279);
xor UO_498 (O_498,N_8534,N_8933);
nand UO_499 (O_499,N_8121,N_8271);
nand UO_500 (O_500,N_9993,N_8444);
nand UO_501 (O_501,N_9254,N_8646);
nand UO_502 (O_502,N_8893,N_8276);
or UO_503 (O_503,N_9125,N_8500);
or UO_504 (O_504,N_9119,N_8608);
nor UO_505 (O_505,N_9387,N_8313);
and UO_506 (O_506,N_9543,N_9908);
and UO_507 (O_507,N_9034,N_9628);
nor UO_508 (O_508,N_8519,N_8428);
nor UO_509 (O_509,N_8774,N_9896);
nand UO_510 (O_510,N_9735,N_8031);
nor UO_511 (O_511,N_8155,N_9366);
or UO_512 (O_512,N_9778,N_8099);
and UO_513 (O_513,N_8533,N_8459);
nand UO_514 (O_514,N_9482,N_9469);
and UO_515 (O_515,N_9004,N_9149);
nor UO_516 (O_516,N_9290,N_8849);
or UO_517 (O_517,N_9480,N_8577);
nor UO_518 (O_518,N_8562,N_9911);
nand UO_519 (O_519,N_9665,N_8177);
nor UO_520 (O_520,N_9346,N_9044);
or UO_521 (O_521,N_9657,N_8805);
nand UO_522 (O_522,N_8264,N_9770);
or UO_523 (O_523,N_8705,N_8616);
and UO_524 (O_524,N_9223,N_8080);
and UO_525 (O_525,N_8063,N_9515);
or UO_526 (O_526,N_9077,N_8072);
nor UO_527 (O_527,N_9003,N_8546);
nand UO_528 (O_528,N_8793,N_9574);
or UO_529 (O_529,N_9785,N_9635);
or UO_530 (O_530,N_9350,N_8698);
or UO_531 (O_531,N_8912,N_9752);
and UO_532 (O_532,N_8232,N_8343);
nor UO_533 (O_533,N_9507,N_9107);
nor UO_534 (O_534,N_9952,N_9019);
and UO_535 (O_535,N_9331,N_9281);
xor UO_536 (O_536,N_8521,N_9245);
nor UO_537 (O_537,N_8363,N_8289);
or UO_538 (O_538,N_9740,N_8992);
or UO_539 (O_539,N_9057,N_8922);
or UO_540 (O_540,N_8084,N_9473);
nor UO_541 (O_541,N_9056,N_8387);
or UO_542 (O_542,N_9717,N_8112);
nor UO_543 (O_543,N_9753,N_9315);
and UO_544 (O_544,N_8385,N_8014);
and UO_545 (O_545,N_9526,N_9016);
nor UO_546 (O_546,N_8843,N_8878);
or UO_547 (O_547,N_8910,N_8206);
or UO_548 (O_548,N_8683,N_8139);
xor UO_549 (O_549,N_8861,N_9641);
and UO_550 (O_550,N_9744,N_8352);
and UO_551 (O_551,N_9227,N_8181);
and UO_552 (O_552,N_9790,N_9681);
nand UO_553 (O_553,N_9756,N_8502);
or UO_554 (O_554,N_8001,N_9108);
nor UO_555 (O_555,N_9345,N_9105);
and UO_556 (O_556,N_8587,N_9151);
nand UO_557 (O_557,N_9973,N_8176);
or UO_558 (O_558,N_9441,N_9094);
nor UO_559 (O_559,N_8166,N_8876);
and UO_560 (O_560,N_9021,N_8558);
and UO_561 (O_561,N_8844,N_9945);
and UO_562 (O_562,N_9417,N_9206);
or UO_563 (O_563,N_9490,N_9504);
nor UO_564 (O_564,N_8221,N_9643);
and UO_565 (O_565,N_9403,N_9336);
and UO_566 (O_566,N_9827,N_9963);
nor UO_567 (O_567,N_9396,N_8065);
nor UO_568 (O_568,N_8416,N_8834);
or UO_569 (O_569,N_9397,N_8772);
nand UO_570 (O_570,N_8688,N_9850);
and UO_571 (O_571,N_8167,N_8822);
nor UO_572 (O_572,N_9158,N_8527);
or UO_573 (O_573,N_8629,N_9373);
nor UO_574 (O_574,N_8060,N_9701);
and UO_575 (O_575,N_8225,N_9335);
or UO_576 (O_576,N_8573,N_8605);
and UO_577 (O_577,N_9216,N_9559);
and UO_578 (O_578,N_8367,N_8293);
or UO_579 (O_579,N_8187,N_9274);
nor UO_580 (O_580,N_8163,N_9941);
nor UO_581 (O_581,N_9620,N_8535);
or UO_582 (O_582,N_9804,N_8621);
and UO_583 (O_583,N_8745,N_8109);
and UO_584 (O_584,N_9739,N_9544);
nand UO_585 (O_585,N_8661,N_8340);
nand UO_586 (O_586,N_8039,N_9310);
nand UO_587 (O_587,N_8650,N_9459);
and UO_588 (O_588,N_9670,N_9520);
nor UO_589 (O_589,N_9845,N_8985);
nor UO_590 (O_590,N_9052,N_9060);
nor UO_591 (O_591,N_9391,N_8996);
or UO_592 (O_592,N_9750,N_9022);
or UO_593 (O_593,N_9208,N_8401);
or UO_594 (O_594,N_9219,N_9521);
or UO_595 (O_595,N_9611,N_8624);
nand UO_596 (O_596,N_8477,N_8870);
nor UO_597 (O_597,N_9832,N_8736);
nor UO_598 (O_598,N_9445,N_8381);
nand UO_599 (O_599,N_9788,N_9844);
or UO_600 (O_600,N_9722,N_9720);
or UO_601 (O_601,N_9834,N_8887);
nand UO_602 (O_602,N_8043,N_8555);
or UO_603 (O_603,N_9109,N_8037);
or UO_604 (O_604,N_9487,N_8129);
nor UO_605 (O_605,N_9260,N_8261);
or UO_606 (O_606,N_9612,N_8284);
or UO_607 (O_607,N_8930,N_8251);
nor UO_608 (O_608,N_9631,N_8800);
xnor UO_609 (O_609,N_9615,N_9432);
or UO_610 (O_610,N_8882,N_9187);
nor UO_611 (O_611,N_8252,N_8520);
nand UO_612 (O_612,N_9915,N_9921);
and UO_613 (O_613,N_9783,N_8297);
nor UO_614 (O_614,N_8411,N_9721);
nand UO_615 (O_615,N_9579,N_8255);
and UO_616 (O_616,N_9191,N_8384);
and UO_617 (O_617,N_9645,N_9819);
and UO_618 (O_618,N_8864,N_8183);
nor UO_619 (O_619,N_9424,N_9156);
nand UO_620 (O_620,N_8033,N_9078);
nor UO_621 (O_621,N_8504,N_9253);
nor UO_622 (O_622,N_8127,N_8945);
nor UO_623 (O_623,N_9805,N_9895);
nor UO_624 (O_624,N_8386,N_9755);
nand UO_625 (O_625,N_8784,N_8644);
xnor UO_626 (O_626,N_9979,N_9577);
nand UO_627 (O_627,N_9139,N_8345);
nand UO_628 (O_628,N_8048,N_8207);
nand UO_629 (O_629,N_9250,N_8815);
nand UO_630 (O_630,N_8997,N_9379);
nand UO_631 (O_631,N_9719,N_9080);
nand UO_632 (O_632,N_8398,N_8368);
or UO_633 (O_633,N_9510,N_8635);
nor UO_634 (O_634,N_9575,N_9297);
or UO_635 (O_635,N_8615,N_9354);
and UO_636 (O_636,N_9128,N_8823);
and UO_637 (O_637,N_8557,N_9478);
or UO_638 (O_638,N_8382,N_8440);
or UO_639 (O_639,N_9467,N_8447);
nand UO_640 (O_640,N_9779,N_8410);
and UO_641 (O_641,N_8204,N_8417);
nor UO_642 (O_642,N_8537,N_8402);
or UO_643 (O_643,N_8787,N_8994);
nand UO_644 (O_644,N_8740,N_8441);
nor UO_645 (O_645,N_8040,N_8361);
or UO_646 (O_646,N_8641,N_9457);
nand UO_647 (O_647,N_8794,N_9853);
nand UO_648 (O_648,N_9006,N_9282);
and UO_649 (O_649,N_8599,N_8664);
nor UO_650 (O_650,N_8332,N_9388);
or UO_651 (O_651,N_8831,N_8604);
or UO_652 (O_652,N_9029,N_9040);
nand UO_653 (O_653,N_8603,N_9549);
and UO_654 (O_654,N_9524,N_9512);
and UO_655 (O_655,N_8448,N_8338);
nand UO_656 (O_656,N_8164,N_8006);
nor UO_657 (O_657,N_8373,N_9815);
nand UO_658 (O_658,N_8366,N_9456);
xor UO_659 (O_659,N_9270,N_8751);
and UO_660 (O_660,N_8959,N_9540);
nand UO_661 (O_661,N_9814,N_9639);
and UO_662 (O_662,N_9776,N_8980);
and UO_663 (O_663,N_8136,N_8663);
and UO_664 (O_664,N_8752,N_9451);
or UO_665 (O_665,N_9633,N_9461);
xnor UO_666 (O_666,N_9711,N_9381);
nand UO_667 (O_667,N_8073,N_8088);
nand UO_668 (O_668,N_9449,N_8057);
nand UO_669 (O_669,N_8662,N_8068);
and UO_670 (O_670,N_9268,N_9436);
nor UO_671 (O_671,N_9849,N_9505);
and UO_672 (O_672,N_9664,N_9311);
nand UO_673 (O_673,N_8528,N_8213);
or UO_674 (O_674,N_9634,N_9032);
and UO_675 (O_675,N_9438,N_9995);
nand UO_676 (O_676,N_9466,N_9841);
or UO_677 (O_677,N_9251,N_8009);
nor UO_678 (O_678,N_9546,N_8320);
and UO_679 (O_679,N_8421,N_8908);
nand UO_680 (O_680,N_8004,N_9763);
and UO_681 (O_681,N_8647,N_9961);
nand UO_682 (O_682,N_8470,N_9924);
nand UO_683 (O_683,N_8672,N_9287);
nor UO_684 (O_684,N_9531,N_9580);
nand UO_685 (O_685,N_8929,N_8826);
nand UO_686 (O_686,N_8571,N_8316);
nand UO_687 (O_687,N_9207,N_8152);
or UO_688 (O_688,N_9189,N_9950);
nor UO_689 (O_689,N_9423,N_8050);
nand UO_690 (O_690,N_9185,N_9702);
nor UO_691 (O_691,N_8239,N_9447);
and UO_692 (O_692,N_9734,N_9553);
or UO_693 (O_693,N_9955,N_8007);
nand UO_694 (O_694,N_8901,N_9937);
and UO_695 (O_695,N_8852,N_9651);
nand UO_696 (O_696,N_9063,N_8290);
nand UO_697 (O_697,N_9843,N_8681);
and UO_698 (O_698,N_9123,N_9444);
or UO_699 (O_699,N_8592,N_8942);
or UO_700 (O_700,N_8172,N_9595);
and UO_701 (O_701,N_9213,N_9046);
nor UO_702 (O_702,N_8265,N_8684);
or UO_703 (O_703,N_9803,N_8425);
and UO_704 (O_704,N_8951,N_9648);
and UO_705 (O_705,N_8436,N_9321);
nor UO_706 (O_706,N_8439,N_8771);
nor UO_707 (O_707,N_8490,N_9767);
nor UO_708 (O_708,N_8886,N_8480);
and UO_709 (O_709,N_8294,N_9333);
and UO_710 (O_710,N_8566,N_9358);
or UO_711 (O_711,N_8192,N_9378);
nand UO_712 (O_712,N_8054,N_8431);
and UO_713 (O_713,N_9401,N_9983);
nand UO_714 (O_714,N_8087,N_9968);
nor UO_715 (O_715,N_8228,N_9741);
and UO_716 (O_716,N_8653,N_8712);
nand UO_717 (O_717,N_8023,N_9118);
xor UO_718 (O_718,N_8614,N_8102);
and UO_719 (O_719,N_9215,N_9960);
nor UO_720 (O_720,N_8881,N_9725);
or UO_721 (O_721,N_9951,N_8833);
or UO_722 (O_722,N_9009,N_8550);
and UO_723 (O_723,N_8095,N_9523);
nand UO_724 (O_724,N_8885,N_8602);
or UO_725 (O_725,N_8468,N_9607);
nand UO_726 (O_726,N_9792,N_8842);
and UO_727 (O_727,N_8240,N_8977);
nor UO_728 (O_728,N_8907,N_8353);
nand UO_729 (O_729,N_8561,N_8730);
nand UO_730 (O_730,N_8281,N_9095);
nand UO_731 (O_731,N_9340,N_8869);
or UO_732 (O_732,N_8578,N_9567);
and UO_733 (O_733,N_8437,N_9106);
and UO_734 (O_734,N_8224,N_8541);
nor UO_735 (O_735,N_8731,N_8902);
nor UO_736 (O_736,N_9914,N_9131);
nand UO_737 (O_737,N_9840,N_8760);
and UO_738 (O_738,N_8318,N_8111);
nand UO_739 (O_739,N_8268,N_8372);
nor UO_740 (O_740,N_9500,N_9226);
nor UO_741 (O_741,N_9743,N_9528);
nand UO_742 (O_742,N_9474,N_9694);
nand UO_743 (O_743,N_8198,N_8450);
xor UO_744 (O_744,N_8715,N_9536);
xnor UO_745 (O_745,N_8141,N_9901);
and UO_746 (O_746,N_9359,N_9193);
nand UO_747 (O_747,N_9563,N_8499);
nand UO_748 (O_748,N_8218,N_8756);
or UO_749 (O_749,N_9237,N_9368);
or UO_750 (O_750,N_9617,N_9642);
or UO_751 (O_751,N_9879,N_8699);
nor UO_752 (O_752,N_8256,N_9122);
or UO_753 (O_753,N_9230,N_8764);
nor UO_754 (O_754,N_9677,N_9088);
nor UO_755 (O_755,N_9542,N_8601);
or UO_756 (O_756,N_8567,N_9418);
nand UO_757 (O_757,N_8765,N_9302);
nor UO_758 (O_758,N_8532,N_9700);
nand UO_759 (O_759,N_9011,N_8069);
nor UO_760 (O_760,N_8214,N_8938);
nor UO_761 (O_761,N_8563,N_8898);
or UO_762 (O_762,N_9316,N_8694);
or UO_763 (O_763,N_9161,N_8126);
or UO_764 (O_764,N_9041,N_9884);
nand UO_765 (O_765,N_9572,N_9818);
nor UO_766 (O_766,N_8911,N_9141);
and UO_767 (O_767,N_8380,N_8669);
or UO_768 (O_768,N_9280,N_8406);
or UO_769 (O_769,N_8734,N_8408);
nand UO_770 (O_770,N_9015,N_8900);
nand UO_771 (O_771,N_9024,N_8359);
nor UO_772 (O_772,N_9255,N_8098);
nand UO_773 (O_773,N_9399,N_9421);
nor UO_774 (O_774,N_9605,N_9836);
nand UO_775 (O_775,N_9238,N_8303);
or UO_776 (O_776,N_8203,N_9440);
or UO_777 (O_777,N_8862,N_8728);
xnor UO_778 (O_778,N_9334,N_9283);
nand UO_779 (O_779,N_9686,N_8937);
nor UO_780 (O_780,N_9231,N_8847);
or UO_781 (O_781,N_8002,N_9393);
and UO_782 (O_782,N_8970,N_9323);
and UO_783 (O_783,N_9214,N_8703);
nand UO_784 (O_784,N_9667,N_9236);
or UO_785 (O_785,N_8593,N_8501);
or UO_786 (O_786,N_8855,N_9012);
nand UO_787 (O_787,N_9890,N_8797);
xnor UO_788 (O_788,N_8085,N_9590);
and UO_789 (O_789,N_9244,N_9891);
and UO_790 (O_790,N_9430,N_9846);
nand UO_791 (O_791,N_9486,N_9806);
nor UO_792 (O_792,N_8963,N_8671);
or UO_793 (O_793,N_9537,N_8737);
and UO_794 (O_794,N_8642,N_9881);
and UO_795 (O_795,N_9513,N_8717);
or UO_796 (O_796,N_9822,N_9017);
and UO_797 (O_797,N_9933,N_9865);
or UO_798 (O_798,N_9618,N_9668);
nand UO_799 (O_799,N_8433,N_8209);
or UO_800 (O_800,N_9494,N_8244);
nor UO_801 (O_801,N_8055,N_9404);
and UO_802 (O_802,N_8780,N_8234);
or UO_803 (O_803,N_8859,N_9928);
and UO_804 (O_804,N_9262,N_8257);
or UO_805 (O_805,N_8222,N_9434);
nor UO_806 (O_806,N_8460,N_9874);
or UO_807 (O_807,N_8711,N_8229);
nor UO_808 (O_808,N_9353,N_9587);
nand UO_809 (O_809,N_8015,N_9344);
and UO_810 (O_810,N_8828,N_9166);
nor UO_811 (O_811,N_8182,N_9349);
or UO_812 (O_812,N_9248,N_9981);
or UO_813 (O_813,N_8079,N_9614);
and UO_814 (O_814,N_8049,N_8144);
and UO_815 (O_815,N_8154,N_9224);
xnor UO_816 (O_816,N_8438,N_8667);
nor UO_817 (O_817,N_8913,N_9644);
nor UO_818 (O_818,N_9889,N_9758);
nor UO_819 (O_819,N_9672,N_8560);
nor UO_820 (O_820,N_9304,N_9154);
nand UO_821 (O_821,N_8216,N_9619);
and UO_822 (O_822,N_9369,N_8104);
and UO_823 (O_823,N_8036,N_9406);
or UO_824 (O_824,N_8721,N_9364);
nand UO_825 (O_825,N_8791,N_8128);
and UO_826 (O_826,N_9133,N_9408);
nand UO_827 (O_827,N_9837,N_8205);
nor UO_828 (O_828,N_9097,N_9674);
or UO_829 (O_829,N_8197,N_9452);
nor UO_830 (O_830,N_8458,N_9812);
nand UO_831 (O_831,N_9654,N_9038);
nand UO_832 (O_832,N_9035,N_8019);
or UO_833 (O_833,N_9437,N_9927);
and UO_834 (O_834,N_8147,N_9932);
and UO_835 (O_835,N_9439,N_8830);
or UO_836 (O_836,N_9205,N_9854);
and UO_837 (O_837,N_8456,N_8768);
nor UO_838 (O_838,N_8409,N_9562);
nand UO_839 (O_839,N_9570,N_9769);
and UO_840 (O_840,N_9211,N_9724);
nand UO_841 (O_841,N_8522,N_8309);
or UO_842 (O_842,N_8777,N_9455);
nand UO_843 (O_843,N_8746,N_9092);
or UO_844 (O_844,N_8818,N_9757);
and UO_845 (O_845,N_9599,N_8032);
and UO_846 (O_846,N_9659,N_9967);
or UO_847 (O_847,N_8524,N_8763);
nor UO_848 (O_848,N_8432,N_9153);
nand UO_849 (O_849,N_9276,N_9514);
and UO_850 (O_850,N_8021,N_9162);
and UO_851 (O_851,N_8583,N_8003);
xnor UO_852 (O_852,N_8305,N_9322);
and UO_853 (O_853,N_9821,N_9435);
nand UO_854 (O_854,N_8796,N_8020);
nand UO_855 (O_855,N_8701,N_8051);
nor UO_856 (O_856,N_8296,N_8783);
nor UO_857 (O_857,N_9126,N_8319);
or UO_858 (O_858,N_8029,N_9638);
nand UO_859 (O_859,N_8423,N_9749);
nand UO_860 (O_860,N_8393,N_9130);
and UO_861 (O_861,N_8067,N_8186);
nand UO_862 (O_862,N_9796,N_8892);
nor UO_863 (O_863,N_8449,N_8113);
nand UO_864 (O_864,N_8078,N_8230);
nor UO_865 (O_865,N_8548,N_9831);
nand UO_866 (O_866,N_8612,N_8277);
nand UO_867 (O_867,N_8249,N_9713);
or UO_868 (O_868,N_8769,N_9045);
or UO_869 (O_869,N_8924,N_8509);
or UO_870 (O_870,N_9695,N_9233);
and UO_871 (O_871,N_8518,N_9450);
xor UO_872 (O_872,N_9037,N_9866);
nand UO_873 (O_873,N_8991,N_8993);
nor UO_874 (O_874,N_8052,N_9318);
and UO_875 (O_875,N_9958,N_9842);
nor UO_876 (O_876,N_8665,N_9241);
nand UO_877 (O_877,N_9008,N_8789);
nor UO_878 (O_878,N_8262,N_8935);
nor UO_879 (O_879,N_9509,N_9637);
and UO_880 (O_880,N_8269,N_8998);
or UO_881 (O_881,N_9994,N_8630);
and UO_882 (O_882,N_8742,N_8622);
nand UO_883 (O_883,N_9069,N_8957);
nor UO_884 (O_884,N_8690,N_9885);
nand UO_885 (O_885,N_9942,N_8426);
nand UO_886 (O_886,N_9944,N_9072);
or UO_887 (O_887,N_8827,N_8540);
xor UO_888 (O_888,N_9771,N_9530);
nor UO_889 (O_889,N_8944,N_8596);
nor UO_890 (O_890,N_8042,N_8327);
or UO_891 (O_891,N_8747,N_8429);
nor UO_892 (O_892,N_9470,N_8950);
or UO_893 (O_893,N_8081,N_8781);
and UO_894 (O_894,N_9516,N_9718);
or UO_895 (O_895,N_9969,N_8860);
or UO_896 (O_896,N_8498,N_8928);
and UO_897 (O_897,N_9113,N_9002);
xnor UO_898 (O_898,N_9751,N_8174);
nand UO_899 (O_899,N_8097,N_8792);
nand UO_900 (O_900,N_8455,N_8322);
or UO_901 (O_901,N_8494,N_8117);
or UO_902 (O_902,N_9314,N_9463);
nor UO_903 (O_903,N_8525,N_9229);
or UO_904 (O_904,N_8196,N_9039);
nand UO_905 (O_905,N_8618,N_9731);
and UO_906 (O_906,N_9239,N_8565);
nor UO_907 (O_907,N_8308,N_8348);
nand UO_908 (O_908,N_8179,N_8201);
or UO_909 (O_909,N_9308,N_8702);
nor UO_910 (O_910,N_8716,N_8696);
or UO_911 (O_911,N_9561,N_9877);
or UO_912 (O_912,N_8914,N_8156);
nand UO_913 (O_913,N_9488,N_9794);
nor UO_914 (O_914,N_8943,N_9005);
and UO_915 (O_915,N_8919,N_9905);
or UO_916 (O_916,N_8435,N_9626);
and UO_917 (O_917,N_8238,N_8896);
nand UO_918 (O_918,N_9984,N_8390);
xor UO_919 (O_919,N_9918,N_9355);
and UO_920 (O_920,N_9708,N_9496);
nor UO_921 (O_921,N_8505,N_9551);
and UO_922 (O_922,N_8809,N_8025);
nand UO_923 (O_923,N_8968,N_9690);
and UO_924 (O_924,N_8735,N_9081);
nand UO_925 (O_925,N_8840,N_9195);
nand UO_926 (O_926,N_9687,N_9389);
nor UO_927 (O_927,N_9795,N_9489);
or UO_928 (O_928,N_9140,N_9594);
nand UO_929 (O_929,N_9774,N_8434);
nand UO_930 (O_930,N_9550,N_8259);
xnor UO_931 (O_931,N_9289,N_9075);
nand UO_932 (O_932,N_8145,N_9103);
nand UO_933 (O_933,N_9917,N_9809);
nor UO_934 (O_934,N_8427,N_9764);
xnor UO_935 (O_935,N_8722,N_8927);
nand UO_936 (O_936,N_9402,N_8034);
nor UO_937 (O_937,N_9142,N_8254);
and UO_938 (O_938,N_9653,N_8226);
and UO_939 (O_939,N_9190,N_8371);
or UO_940 (O_940,N_8314,N_9288);
nor UO_941 (O_941,N_9959,N_8536);
nor UO_942 (O_942,N_9714,N_8726);
and UO_943 (O_943,N_8506,N_9294);
and UO_944 (O_944,N_8027,N_9922);
or UO_945 (O_945,N_8595,N_9201);
and UO_946 (O_946,N_9356,N_8301);
or UO_947 (O_947,N_9975,N_8202);
nor UO_948 (O_948,N_9295,N_9910);
nor UO_949 (O_949,N_8419,N_9050);
xnor UO_950 (O_950,N_9367,N_9164);
or UO_951 (O_951,N_8510,N_8955);
or UO_952 (O_952,N_9484,N_8488);
and UO_953 (O_953,N_9410,N_8471);
or UO_954 (O_954,N_8559,N_9793);
and UO_955 (O_955,N_9210,N_8354);
and UO_956 (O_956,N_8899,N_8451);
nor UO_957 (O_957,N_9085,N_8790);
nand UO_958 (O_958,N_8486,N_8123);
or UO_959 (O_959,N_8574,N_9925);
and UO_960 (O_960,N_8066,N_8649);
and UO_961 (O_961,N_8851,N_8315);
nand UO_962 (O_962,N_9661,N_9348);
nand UO_963 (O_963,N_9899,N_9728);
nand UO_964 (O_964,N_8697,N_8798);
and UO_965 (O_965,N_8689,N_9996);
nand UO_966 (O_966,N_8347,N_8245);
and UO_967 (O_967,N_8074,N_8607);
nor UO_968 (O_968,N_8948,N_9220);
nor UO_969 (O_969,N_9564,N_9704);
nand UO_970 (O_970,N_9746,N_9492);
nand UO_971 (O_971,N_9824,N_8233);
nand UO_972 (O_972,N_9096,N_8369);
and UO_973 (O_973,N_9362,N_9888);
nor UO_974 (O_974,N_9376,N_8895);
nor UO_975 (O_975,N_8317,N_9863);
nor UO_976 (O_976,N_8868,N_9442);
and UO_977 (O_977,N_8457,N_8802);
and UO_978 (O_978,N_9730,N_8708);
nand UO_979 (O_979,N_8335,N_9171);
and UO_980 (O_980,N_9413,N_9682);
xor UO_981 (O_981,N_9581,N_9789);
nor UO_982 (O_982,N_9775,N_8418);
or UO_983 (O_983,N_9266,N_8873);
nor UO_984 (O_984,N_9798,N_9472);
nand UO_985 (O_985,N_8150,N_9493);
or UO_986 (O_986,N_9569,N_8857);
or UO_987 (O_987,N_9601,N_8757);
nor UO_988 (O_988,N_8973,N_8539);
or UO_989 (O_989,N_9529,N_8185);
or UO_990 (O_990,N_8853,N_9880);
nand UO_991 (O_991,N_9991,N_8377);
nand UO_992 (O_992,N_8364,N_9894);
and UO_993 (O_993,N_9074,N_8495);
xnor UO_994 (O_994,N_9976,N_9591);
nand UO_995 (O_995,N_9020,N_8915);
xor UO_996 (O_996,N_8568,N_8939);
nor UO_997 (O_997,N_9112,N_8625);
and UO_998 (O_998,N_9875,N_8465);
nor UO_999 (O_999,N_8454,N_8594);
or UO_1000 (O_1000,N_8314,N_8626);
or UO_1001 (O_1001,N_8894,N_8376);
and UO_1002 (O_1002,N_9005,N_8767);
or UO_1003 (O_1003,N_9183,N_9801);
or UO_1004 (O_1004,N_8202,N_8040);
or UO_1005 (O_1005,N_9513,N_8910);
or UO_1006 (O_1006,N_9391,N_8268);
nand UO_1007 (O_1007,N_9786,N_9379);
and UO_1008 (O_1008,N_8776,N_9267);
and UO_1009 (O_1009,N_8632,N_9641);
nand UO_1010 (O_1010,N_8191,N_9668);
and UO_1011 (O_1011,N_8004,N_9289);
and UO_1012 (O_1012,N_9054,N_8927);
and UO_1013 (O_1013,N_8297,N_9387);
or UO_1014 (O_1014,N_9034,N_8234);
and UO_1015 (O_1015,N_9222,N_9122);
nand UO_1016 (O_1016,N_9172,N_8917);
nand UO_1017 (O_1017,N_9366,N_9637);
nand UO_1018 (O_1018,N_9932,N_9808);
or UO_1019 (O_1019,N_9441,N_8363);
and UO_1020 (O_1020,N_9726,N_9293);
or UO_1021 (O_1021,N_9438,N_8736);
and UO_1022 (O_1022,N_8013,N_9516);
and UO_1023 (O_1023,N_9457,N_8634);
xnor UO_1024 (O_1024,N_9086,N_8270);
nor UO_1025 (O_1025,N_9323,N_9085);
nor UO_1026 (O_1026,N_8750,N_9177);
nor UO_1027 (O_1027,N_9096,N_9804);
nor UO_1028 (O_1028,N_8138,N_9635);
or UO_1029 (O_1029,N_9267,N_9133);
or UO_1030 (O_1030,N_8202,N_9730);
and UO_1031 (O_1031,N_8653,N_8098);
or UO_1032 (O_1032,N_9581,N_8526);
nor UO_1033 (O_1033,N_8594,N_9209);
nor UO_1034 (O_1034,N_8172,N_8571);
or UO_1035 (O_1035,N_8134,N_9396);
nand UO_1036 (O_1036,N_9314,N_8054);
and UO_1037 (O_1037,N_9369,N_8474);
xnor UO_1038 (O_1038,N_9265,N_9011);
nor UO_1039 (O_1039,N_9782,N_9298);
and UO_1040 (O_1040,N_8551,N_8663);
and UO_1041 (O_1041,N_8887,N_9064);
and UO_1042 (O_1042,N_9362,N_9033);
xor UO_1043 (O_1043,N_9199,N_8584);
or UO_1044 (O_1044,N_8901,N_8799);
or UO_1045 (O_1045,N_8849,N_8941);
nor UO_1046 (O_1046,N_8635,N_8195);
and UO_1047 (O_1047,N_8757,N_8578);
or UO_1048 (O_1048,N_9689,N_8024);
and UO_1049 (O_1049,N_8944,N_8103);
and UO_1050 (O_1050,N_8789,N_8471);
nor UO_1051 (O_1051,N_8154,N_9820);
nor UO_1052 (O_1052,N_9229,N_9895);
or UO_1053 (O_1053,N_8583,N_9498);
or UO_1054 (O_1054,N_8566,N_8516);
or UO_1055 (O_1055,N_9446,N_8437);
or UO_1056 (O_1056,N_8723,N_9460);
nand UO_1057 (O_1057,N_9007,N_9368);
and UO_1058 (O_1058,N_8728,N_8822);
nor UO_1059 (O_1059,N_9071,N_8571);
and UO_1060 (O_1060,N_9584,N_9238);
or UO_1061 (O_1061,N_9588,N_9161);
nand UO_1062 (O_1062,N_9719,N_9392);
nor UO_1063 (O_1063,N_8729,N_8860);
and UO_1064 (O_1064,N_9659,N_9507);
nor UO_1065 (O_1065,N_9319,N_8730);
or UO_1066 (O_1066,N_8300,N_9235);
and UO_1067 (O_1067,N_8424,N_8727);
and UO_1068 (O_1068,N_9937,N_8859);
nor UO_1069 (O_1069,N_8511,N_9111);
or UO_1070 (O_1070,N_8927,N_9370);
nor UO_1071 (O_1071,N_8838,N_8722);
nand UO_1072 (O_1072,N_8362,N_9362);
nor UO_1073 (O_1073,N_9618,N_9609);
nand UO_1074 (O_1074,N_8329,N_9856);
or UO_1075 (O_1075,N_9559,N_8327);
nand UO_1076 (O_1076,N_9249,N_9369);
or UO_1077 (O_1077,N_9606,N_8682);
nor UO_1078 (O_1078,N_8243,N_8706);
nor UO_1079 (O_1079,N_8891,N_9756);
or UO_1080 (O_1080,N_8702,N_8445);
nand UO_1081 (O_1081,N_9473,N_8069);
nor UO_1082 (O_1082,N_8055,N_9088);
or UO_1083 (O_1083,N_9887,N_9657);
or UO_1084 (O_1084,N_8451,N_9057);
nand UO_1085 (O_1085,N_9164,N_8357);
and UO_1086 (O_1086,N_8727,N_8833);
nand UO_1087 (O_1087,N_8941,N_8434);
nand UO_1088 (O_1088,N_9497,N_8404);
or UO_1089 (O_1089,N_9717,N_9905);
nand UO_1090 (O_1090,N_9882,N_8080);
nand UO_1091 (O_1091,N_8683,N_9599);
and UO_1092 (O_1092,N_9963,N_8330);
xnor UO_1093 (O_1093,N_8781,N_8208);
nand UO_1094 (O_1094,N_8535,N_9407);
nand UO_1095 (O_1095,N_9779,N_9161);
nand UO_1096 (O_1096,N_8573,N_9229);
nand UO_1097 (O_1097,N_8646,N_9904);
and UO_1098 (O_1098,N_8917,N_9521);
or UO_1099 (O_1099,N_8197,N_8393);
and UO_1100 (O_1100,N_9149,N_8448);
or UO_1101 (O_1101,N_8595,N_9912);
xor UO_1102 (O_1102,N_8944,N_8163);
xor UO_1103 (O_1103,N_9856,N_8746);
and UO_1104 (O_1104,N_9554,N_9115);
and UO_1105 (O_1105,N_8914,N_8493);
or UO_1106 (O_1106,N_8729,N_8294);
nor UO_1107 (O_1107,N_8544,N_8584);
or UO_1108 (O_1108,N_9435,N_8325);
and UO_1109 (O_1109,N_9692,N_9541);
or UO_1110 (O_1110,N_8856,N_8837);
nor UO_1111 (O_1111,N_9860,N_8407);
and UO_1112 (O_1112,N_9460,N_9234);
nand UO_1113 (O_1113,N_8861,N_8264);
nor UO_1114 (O_1114,N_9970,N_9927);
nand UO_1115 (O_1115,N_9315,N_8432);
nand UO_1116 (O_1116,N_8434,N_9877);
xor UO_1117 (O_1117,N_8539,N_8415);
nor UO_1118 (O_1118,N_8513,N_9984);
nor UO_1119 (O_1119,N_8139,N_8704);
and UO_1120 (O_1120,N_8605,N_9025);
nor UO_1121 (O_1121,N_9794,N_8763);
or UO_1122 (O_1122,N_9720,N_9747);
or UO_1123 (O_1123,N_8810,N_9160);
nor UO_1124 (O_1124,N_9758,N_9894);
and UO_1125 (O_1125,N_9701,N_9778);
nor UO_1126 (O_1126,N_8687,N_8521);
nand UO_1127 (O_1127,N_9821,N_8525);
or UO_1128 (O_1128,N_8126,N_9597);
and UO_1129 (O_1129,N_9424,N_9594);
or UO_1130 (O_1130,N_8064,N_9709);
and UO_1131 (O_1131,N_9705,N_8175);
or UO_1132 (O_1132,N_9325,N_9501);
nand UO_1133 (O_1133,N_9658,N_9472);
nor UO_1134 (O_1134,N_8719,N_8167);
or UO_1135 (O_1135,N_8532,N_8303);
nand UO_1136 (O_1136,N_9864,N_9229);
or UO_1137 (O_1137,N_8167,N_8349);
nand UO_1138 (O_1138,N_8077,N_9445);
nor UO_1139 (O_1139,N_9568,N_8297);
nand UO_1140 (O_1140,N_8492,N_9881);
nor UO_1141 (O_1141,N_8202,N_8312);
nor UO_1142 (O_1142,N_8534,N_8436);
or UO_1143 (O_1143,N_9672,N_9449);
xnor UO_1144 (O_1144,N_8182,N_8991);
and UO_1145 (O_1145,N_9303,N_9005);
or UO_1146 (O_1146,N_9823,N_8329);
nand UO_1147 (O_1147,N_9783,N_9231);
or UO_1148 (O_1148,N_8715,N_8570);
nor UO_1149 (O_1149,N_8170,N_8672);
nor UO_1150 (O_1150,N_9886,N_8620);
nand UO_1151 (O_1151,N_8966,N_9462);
nor UO_1152 (O_1152,N_8834,N_8763);
nand UO_1153 (O_1153,N_8619,N_9823);
nand UO_1154 (O_1154,N_8471,N_9720);
nor UO_1155 (O_1155,N_9803,N_8463);
and UO_1156 (O_1156,N_9443,N_9347);
nor UO_1157 (O_1157,N_9137,N_9341);
nor UO_1158 (O_1158,N_8393,N_8934);
or UO_1159 (O_1159,N_8259,N_9658);
or UO_1160 (O_1160,N_8018,N_9822);
or UO_1161 (O_1161,N_8077,N_9679);
or UO_1162 (O_1162,N_8102,N_8574);
or UO_1163 (O_1163,N_9648,N_8832);
and UO_1164 (O_1164,N_8439,N_9757);
or UO_1165 (O_1165,N_9739,N_9914);
or UO_1166 (O_1166,N_8126,N_9036);
nand UO_1167 (O_1167,N_8325,N_9113);
and UO_1168 (O_1168,N_8222,N_9343);
nand UO_1169 (O_1169,N_9349,N_8113);
nand UO_1170 (O_1170,N_9972,N_9241);
or UO_1171 (O_1171,N_9606,N_9037);
xnor UO_1172 (O_1172,N_9111,N_8972);
xnor UO_1173 (O_1173,N_8352,N_9291);
nor UO_1174 (O_1174,N_9465,N_8522);
nor UO_1175 (O_1175,N_9556,N_9045);
nor UO_1176 (O_1176,N_9736,N_8923);
xor UO_1177 (O_1177,N_8196,N_8176);
and UO_1178 (O_1178,N_8187,N_8638);
nor UO_1179 (O_1179,N_9198,N_9781);
nor UO_1180 (O_1180,N_8997,N_9899);
or UO_1181 (O_1181,N_8044,N_8715);
nor UO_1182 (O_1182,N_9895,N_9627);
or UO_1183 (O_1183,N_8686,N_8272);
nor UO_1184 (O_1184,N_9484,N_8898);
or UO_1185 (O_1185,N_9249,N_9607);
nand UO_1186 (O_1186,N_9906,N_9830);
nor UO_1187 (O_1187,N_9558,N_8314);
nor UO_1188 (O_1188,N_8318,N_9524);
or UO_1189 (O_1189,N_8916,N_8719);
and UO_1190 (O_1190,N_8610,N_9656);
and UO_1191 (O_1191,N_9714,N_9548);
nand UO_1192 (O_1192,N_9675,N_9537);
and UO_1193 (O_1193,N_9395,N_8570);
or UO_1194 (O_1194,N_9782,N_9713);
nor UO_1195 (O_1195,N_9030,N_8840);
and UO_1196 (O_1196,N_9374,N_9543);
or UO_1197 (O_1197,N_8931,N_9070);
and UO_1198 (O_1198,N_8950,N_9517);
and UO_1199 (O_1199,N_9480,N_8648);
or UO_1200 (O_1200,N_9754,N_9588);
and UO_1201 (O_1201,N_8549,N_9030);
and UO_1202 (O_1202,N_9910,N_8073);
nand UO_1203 (O_1203,N_8531,N_8046);
nor UO_1204 (O_1204,N_9426,N_9327);
nor UO_1205 (O_1205,N_8473,N_8799);
and UO_1206 (O_1206,N_9577,N_8055);
nand UO_1207 (O_1207,N_8538,N_8890);
nand UO_1208 (O_1208,N_8136,N_9007);
or UO_1209 (O_1209,N_9220,N_9320);
and UO_1210 (O_1210,N_8148,N_8186);
and UO_1211 (O_1211,N_8365,N_8983);
or UO_1212 (O_1212,N_8338,N_8022);
nor UO_1213 (O_1213,N_8570,N_9020);
nor UO_1214 (O_1214,N_8230,N_9951);
and UO_1215 (O_1215,N_9077,N_8271);
nor UO_1216 (O_1216,N_9758,N_8161);
or UO_1217 (O_1217,N_8687,N_9748);
xnor UO_1218 (O_1218,N_9237,N_8974);
or UO_1219 (O_1219,N_8333,N_9561);
nand UO_1220 (O_1220,N_8635,N_8291);
and UO_1221 (O_1221,N_9825,N_9585);
nand UO_1222 (O_1222,N_9852,N_9550);
or UO_1223 (O_1223,N_8398,N_9892);
or UO_1224 (O_1224,N_8725,N_9980);
and UO_1225 (O_1225,N_8089,N_8185);
nand UO_1226 (O_1226,N_8613,N_8359);
or UO_1227 (O_1227,N_9515,N_9972);
or UO_1228 (O_1228,N_8717,N_8275);
nand UO_1229 (O_1229,N_8569,N_9691);
nor UO_1230 (O_1230,N_9258,N_9361);
or UO_1231 (O_1231,N_9558,N_8506);
or UO_1232 (O_1232,N_9833,N_8375);
nand UO_1233 (O_1233,N_8573,N_9499);
or UO_1234 (O_1234,N_8812,N_9572);
or UO_1235 (O_1235,N_8659,N_9442);
nor UO_1236 (O_1236,N_9237,N_9561);
nor UO_1237 (O_1237,N_8892,N_8739);
nand UO_1238 (O_1238,N_8915,N_8859);
and UO_1239 (O_1239,N_8809,N_9537);
nand UO_1240 (O_1240,N_8191,N_8643);
or UO_1241 (O_1241,N_8745,N_8458);
nor UO_1242 (O_1242,N_9960,N_8853);
nor UO_1243 (O_1243,N_9557,N_9414);
or UO_1244 (O_1244,N_8687,N_8288);
nand UO_1245 (O_1245,N_9041,N_9389);
nand UO_1246 (O_1246,N_9401,N_9395);
nor UO_1247 (O_1247,N_8557,N_8810);
or UO_1248 (O_1248,N_8503,N_8251);
nand UO_1249 (O_1249,N_9667,N_9561);
nand UO_1250 (O_1250,N_9486,N_9824);
and UO_1251 (O_1251,N_8826,N_9336);
or UO_1252 (O_1252,N_9042,N_8122);
nor UO_1253 (O_1253,N_8635,N_8789);
or UO_1254 (O_1254,N_9516,N_8642);
and UO_1255 (O_1255,N_8349,N_8563);
or UO_1256 (O_1256,N_8149,N_8113);
nor UO_1257 (O_1257,N_9031,N_9675);
and UO_1258 (O_1258,N_8132,N_8627);
nor UO_1259 (O_1259,N_9902,N_8723);
and UO_1260 (O_1260,N_9020,N_8717);
nand UO_1261 (O_1261,N_8482,N_8525);
or UO_1262 (O_1262,N_9194,N_8596);
and UO_1263 (O_1263,N_9553,N_9684);
nor UO_1264 (O_1264,N_8116,N_9477);
or UO_1265 (O_1265,N_9363,N_8939);
nor UO_1266 (O_1266,N_8983,N_8988);
or UO_1267 (O_1267,N_8796,N_9987);
and UO_1268 (O_1268,N_9361,N_8373);
and UO_1269 (O_1269,N_9373,N_8417);
xnor UO_1270 (O_1270,N_9339,N_8528);
or UO_1271 (O_1271,N_9514,N_9918);
nand UO_1272 (O_1272,N_9100,N_8846);
or UO_1273 (O_1273,N_9387,N_9072);
and UO_1274 (O_1274,N_8656,N_8321);
nand UO_1275 (O_1275,N_8143,N_9652);
nand UO_1276 (O_1276,N_8758,N_8464);
or UO_1277 (O_1277,N_9562,N_9590);
and UO_1278 (O_1278,N_8159,N_9547);
xor UO_1279 (O_1279,N_8218,N_8452);
or UO_1280 (O_1280,N_9917,N_9257);
nor UO_1281 (O_1281,N_8665,N_9984);
xor UO_1282 (O_1282,N_9912,N_9482);
or UO_1283 (O_1283,N_8376,N_9564);
nand UO_1284 (O_1284,N_9198,N_8470);
nor UO_1285 (O_1285,N_8407,N_8242);
xor UO_1286 (O_1286,N_8428,N_8903);
nand UO_1287 (O_1287,N_9039,N_9059);
and UO_1288 (O_1288,N_8122,N_9915);
or UO_1289 (O_1289,N_8737,N_8554);
and UO_1290 (O_1290,N_9096,N_8589);
nor UO_1291 (O_1291,N_8356,N_9473);
nand UO_1292 (O_1292,N_9194,N_9368);
nand UO_1293 (O_1293,N_9254,N_9955);
and UO_1294 (O_1294,N_8461,N_9343);
nand UO_1295 (O_1295,N_8947,N_9940);
or UO_1296 (O_1296,N_8828,N_9130);
and UO_1297 (O_1297,N_8304,N_9354);
or UO_1298 (O_1298,N_8382,N_9419);
nand UO_1299 (O_1299,N_9936,N_9353);
nand UO_1300 (O_1300,N_9286,N_9543);
nor UO_1301 (O_1301,N_9449,N_8852);
nand UO_1302 (O_1302,N_9703,N_8513);
nand UO_1303 (O_1303,N_8935,N_8514);
nor UO_1304 (O_1304,N_8979,N_8329);
nand UO_1305 (O_1305,N_8262,N_9129);
nand UO_1306 (O_1306,N_8696,N_8465);
or UO_1307 (O_1307,N_9688,N_9298);
nor UO_1308 (O_1308,N_9543,N_9827);
nand UO_1309 (O_1309,N_9213,N_9968);
and UO_1310 (O_1310,N_9158,N_8491);
nor UO_1311 (O_1311,N_9419,N_8394);
and UO_1312 (O_1312,N_9943,N_9066);
nor UO_1313 (O_1313,N_8483,N_8948);
nand UO_1314 (O_1314,N_8888,N_9247);
or UO_1315 (O_1315,N_9368,N_9145);
nor UO_1316 (O_1316,N_9905,N_8169);
or UO_1317 (O_1317,N_8217,N_9125);
or UO_1318 (O_1318,N_9948,N_9136);
xor UO_1319 (O_1319,N_8580,N_9010);
nand UO_1320 (O_1320,N_8447,N_9906);
and UO_1321 (O_1321,N_8310,N_8744);
or UO_1322 (O_1322,N_8306,N_9426);
or UO_1323 (O_1323,N_9947,N_8964);
nor UO_1324 (O_1324,N_9676,N_9877);
xnor UO_1325 (O_1325,N_9869,N_8276);
nor UO_1326 (O_1326,N_8794,N_9110);
or UO_1327 (O_1327,N_8459,N_8066);
nand UO_1328 (O_1328,N_9354,N_9439);
or UO_1329 (O_1329,N_9478,N_9310);
or UO_1330 (O_1330,N_8807,N_8084);
nand UO_1331 (O_1331,N_9291,N_8111);
and UO_1332 (O_1332,N_9335,N_8899);
nand UO_1333 (O_1333,N_9913,N_8478);
and UO_1334 (O_1334,N_9464,N_8213);
nor UO_1335 (O_1335,N_9524,N_8878);
or UO_1336 (O_1336,N_8897,N_8683);
nand UO_1337 (O_1337,N_8732,N_9124);
and UO_1338 (O_1338,N_8015,N_8473);
and UO_1339 (O_1339,N_9381,N_8757);
and UO_1340 (O_1340,N_8290,N_8532);
nand UO_1341 (O_1341,N_9366,N_8369);
or UO_1342 (O_1342,N_9800,N_8692);
xor UO_1343 (O_1343,N_8706,N_8235);
nand UO_1344 (O_1344,N_8274,N_8342);
or UO_1345 (O_1345,N_9921,N_9911);
or UO_1346 (O_1346,N_8701,N_9482);
and UO_1347 (O_1347,N_8132,N_9528);
nand UO_1348 (O_1348,N_8598,N_8417);
or UO_1349 (O_1349,N_9616,N_9787);
or UO_1350 (O_1350,N_9513,N_8266);
nor UO_1351 (O_1351,N_8745,N_9484);
nand UO_1352 (O_1352,N_9007,N_8549);
nor UO_1353 (O_1353,N_8582,N_9956);
and UO_1354 (O_1354,N_8738,N_9043);
nand UO_1355 (O_1355,N_9689,N_9602);
or UO_1356 (O_1356,N_9989,N_8433);
and UO_1357 (O_1357,N_9581,N_9916);
and UO_1358 (O_1358,N_8662,N_8788);
and UO_1359 (O_1359,N_9230,N_9506);
and UO_1360 (O_1360,N_8311,N_8549);
and UO_1361 (O_1361,N_9008,N_8442);
and UO_1362 (O_1362,N_9888,N_8051);
and UO_1363 (O_1363,N_9927,N_8750);
nor UO_1364 (O_1364,N_8626,N_8735);
or UO_1365 (O_1365,N_8174,N_8481);
and UO_1366 (O_1366,N_8593,N_9373);
and UO_1367 (O_1367,N_8500,N_8707);
nor UO_1368 (O_1368,N_9344,N_8222);
nor UO_1369 (O_1369,N_8701,N_8695);
nand UO_1370 (O_1370,N_9914,N_9748);
nor UO_1371 (O_1371,N_8542,N_8902);
or UO_1372 (O_1372,N_9005,N_9978);
xor UO_1373 (O_1373,N_8634,N_9492);
or UO_1374 (O_1374,N_9253,N_9712);
or UO_1375 (O_1375,N_9024,N_9207);
or UO_1376 (O_1376,N_9354,N_8375);
nor UO_1377 (O_1377,N_8193,N_8956);
xnor UO_1378 (O_1378,N_8790,N_9923);
or UO_1379 (O_1379,N_9860,N_9415);
nand UO_1380 (O_1380,N_9733,N_8721);
or UO_1381 (O_1381,N_8077,N_9201);
or UO_1382 (O_1382,N_9409,N_9865);
nand UO_1383 (O_1383,N_8567,N_9693);
nor UO_1384 (O_1384,N_9120,N_8479);
nand UO_1385 (O_1385,N_9915,N_8092);
or UO_1386 (O_1386,N_9944,N_9856);
or UO_1387 (O_1387,N_9624,N_8292);
and UO_1388 (O_1388,N_8095,N_8869);
nand UO_1389 (O_1389,N_8650,N_9104);
nor UO_1390 (O_1390,N_9599,N_9439);
nor UO_1391 (O_1391,N_8380,N_8122);
nor UO_1392 (O_1392,N_9283,N_9221);
nand UO_1393 (O_1393,N_9659,N_9813);
xnor UO_1394 (O_1394,N_8696,N_8532);
xor UO_1395 (O_1395,N_8194,N_9557);
nand UO_1396 (O_1396,N_9115,N_9660);
nor UO_1397 (O_1397,N_9735,N_8206);
or UO_1398 (O_1398,N_9780,N_9872);
nand UO_1399 (O_1399,N_9282,N_9343);
nand UO_1400 (O_1400,N_8403,N_9329);
or UO_1401 (O_1401,N_9352,N_8053);
and UO_1402 (O_1402,N_8877,N_9313);
nor UO_1403 (O_1403,N_9567,N_8679);
nand UO_1404 (O_1404,N_8166,N_9433);
and UO_1405 (O_1405,N_8175,N_8561);
and UO_1406 (O_1406,N_8831,N_9680);
nor UO_1407 (O_1407,N_9487,N_8335);
nor UO_1408 (O_1408,N_9388,N_9297);
and UO_1409 (O_1409,N_8425,N_9679);
and UO_1410 (O_1410,N_9444,N_9080);
and UO_1411 (O_1411,N_8493,N_9030);
nand UO_1412 (O_1412,N_8543,N_9006);
nand UO_1413 (O_1413,N_8789,N_9806);
nor UO_1414 (O_1414,N_9965,N_8522);
nor UO_1415 (O_1415,N_9176,N_9549);
nand UO_1416 (O_1416,N_9349,N_8854);
or UO_1417 (O_1417,N_8493,N_8281);
nor UO_1418 (O_1418,N_9408,N_9180);
nor UO_1419 (O_1419,N_9448,N_9458);
nand UO_1420 (O_1420,N_9611,N_9567);
or UO_1421 (O_1421,N_9204,N_8787);
or UO_1422 (O_1422,N_9098,N_9728);
nand UO_1423 (O_1423,N_8479,N_8853);
nor UO_1424 (O_1424,N_9264,N_9376);
and UO_1425 (O_1425,N_9028,N_9482);
and UO_1426 (O_1426,N_8838,N_9029);
and UO_1427 (O_1427,N_8734,N_8290);
xor UO_1428 (O_1428,N_9230,N_8311);
nor UO_1429 (O_1429,N_9535,N_8069);
and UO_1430 (O_1430,N_8586,N_9903);
or UO_1431 (O_1431,N_9210,N_8215);
nor UO_1432 (O_1432,N_9343,N_8771);
nor UO_1433 (O_1433,N_9243,N_8590);
xor UO_1434 (O_1434,N_9844,N_9170);
nand UO_1435 (O_1435,N_8772,N_9084);
nand UO_1436 (O_1436,N_9321,N_8121);
or UO_1437 (O_1437,N_8932,N_8719);
nor UO_1438 (O_1438,N_8692,N_8077);
nand UO_1439 (O_1439,N_9142,N_8120);
nor UO_1440 (O_1440,N_8063,N_8041);
or UO_1441 (O_1441,N_9475,N_9712);
and UO_1442 (O_1442,N_8767,N_9745);
xnor UO_1443 (O_1443,N_8163,N_9848);
and UO_1444 (O_1444,N_8792,N_9617);
nor UO_1445 (O_1445,N_9432,N_8619);
and UO_1446 (O_1446,N_9271,N_9854);
and UO_1447 (O_1447,N_9225,N_9884);
nand UO_1448 (O_1448,N_8612,N_8389);
and UO_1449 (O_1449,N_8065,N_9038);
nor UO_1450 (O_1450,N_9611,N_8566);
and UO_1451 (O_1451,N_8023,N_8052);
and UO_1452 (O_1452,N_9944,N_8321);
nor UO_1453 (O_1453,N_9823,N_8998);
nor UO_1454 (O_1454,N_9298,N_9370);
and UO_1455 (O_1455,N_9783,N_9723);
nand UO_1456 (O_1456,N_9303,N_8028);
or UO_1457 (O_1457,N_8922,N_9975);
nor UO_1458 (O_1458,N_8652,N_9171);
nand UO_1459 (O_1459,N_9200,N_8077);
nor UO_1460 (O_1460,N_9500,N_9459);
or UO_1461 (O_1461,N_8305,N_8259);
nand UO_1462 (O_1462,N_8806,N_9095);
nor UO_1463 (O_1463,N_9161,N_8488);
nor UO_1464 (O_1464,N_9128,N_8737);
nand UO_1465 (O_1465,N_8069,N_9725);
nor UO_1466 (O_1466,N_9138,N_8008);
and UO_1467 (O_1467,N_8960,N_8331);
nand UO_1468 (O_1468,N_9343,N_8486);
and UO_1469 (O_1469,N_8265,N_9286);
or UO_1470 (O_1470,N_9676,N_9068);
nand UO_1471 (O_1471,N_9452,N_8220);
or UO_1472 (O_1472,N_8372,N_8192);
or UO_1473 (O_1473,N_9987,N_9265);
or UO_1474 (O_1474,N_8521,N_9321);
nor UO_1475 (O_1475,N_8214,N_8837);
xor UO_1476 (O_1476,N_8277,N_8043);
and UO_1477 (O_1477,N_8885,N_8995);
or UO_1478 (O_1478,N_8710,N_9224);
nand UO_1479 (O_1479,N_8477,N_9542);
nor UO_1480 (O_1480,N_9373,N_8854);
nand UO_1481 (O_1481,N_9073,N_9295);
nand UO_1482 (O_1482,N_8326,N_9252);
or UO_1483 (O_1483,N_8383,N_9975);
nand UO_1484 (O_1484,N_8345,N_9226);
and UO_1485 (O_1485,N_9732,N_8999);
or UO_1486 (O_1486,N_9378,N_9330);
nor UO_1487 (O_1487,N_8339,N_9307);
or UO_1488 (O_1488,N_9883,N_9534);
nand UO_1489 (O_1489,N_8079,N_9863);
nor UO_1490 (O_1490,N_9858,N_9272);
or UO_1491 (O_1491,N_8124,N_9292);
and UO_1492 (O_1492,N_8214,N_8246);
and UO_1493 (O_1493,N_8763,N_8878);
nand UO_1494 (O_1494,N_9005,N_8219);
nor UO_1495 (O_1495,N_9502,N_9296);
nand UO_1496 (O_1496,N_8028,N_8966);
or UO_1497 (O_1497,N_9136,N_8375);
nand UO_1498 (O_1498,N_8530,N_8584);
or UO_1499 (O_1499,N_8392,N_9517);
endmodule