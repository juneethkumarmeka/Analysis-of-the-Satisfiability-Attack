module basic_750_5000_1000_25_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_320,In_545);
nand U1 (N_1,In_508,In_187);
nor U2 (N_2,In_33,In_182);
and U3 (N_3,In_408,In_624);
or U4 (N_4,In_691,In_150);
nand U5 (N_5,In_319,In_701);
and U6 (N_6,In_711,In_232);
nor U7 (N_7,In_642,In_0);
xnor U8 (N_8,In_739,In_548);
and U9 (N_9,In_269,In_174);
and U10 (N_10,In_335,In_189);
or U11 (N_11,In_442,In_564);
nor U12 (N_12,In_213,In_115);
or U13 (N_13,In_70,In_585);
nand U14 (N_14,In_374,In_126);
nor U15 (N_15,In_721,In_541);
or U16 (N_16,In_388,In_26);
and U17 (N_17,In_741,In_121);
nor U18 (N_18,In_162,In_521);
or U19 (N_19,In_295,In_418);
nor U20 (N_20,In_119,In_364);
nor U21 (N_21,In_127,In_202);
nor U22 (N_22,In_568,In_567);
and U23 (N_23,In_192,In_78);
or U24 (N_24,In_230,In_738);
or U25 (N_25,In_608,In_594);
nand U26 (N_26,In_318,In_358);
xor U27 (N_27,In_407,In_484);
xnor U28 (N_28,In_98,In_490);
or U29 (N_29,In_460,In_373);
xor U30 (N_30,In_720,In_402);
xor U31 (N_31,In_307,In_493);
nor U32 (N_32,In_625,In_728);
xnor U33 (N_33,In_404,In_241);
or U34 (N_34,In_11,In_497);
nand U35 (N_35,In_570,In_532);
or U36 (N_36,In_592,In_433);
or U37 (N_37,In_539,In_468);
xnor U38 (N_38,In_535,In_392);
xnor U39 (N_39,In_399,In_76);
nor U40 (N_40,In_572,In_324);
xor U41 (N_41,In_540,In_247);
and U42 (N_42,In_130,In_748);
xor U43 (N_43,In_124,In_429);
and U44 (N_44,In_84,In_195);
xnor U45 (N_45,In_657,In_290);
and U46 (N_46,In_176,In_527);
and U47 (N_47,In_149,In_282);
xnor U48 (N_48,In_467,In_495);
nor U49 (N_49,In_59,In_743);
nor U50 (N_50,In_310,In_737);
nand U51 (N_51,In_466,In_219);
nor U52 (N_52,In_113,In_89);
or U53 (N_53,In_57,In_574);
nor U54 (N_54,In_185,In_413);
xnor U55 (N_55,In_622,In_357);
and U56 (N_56,In_38,In_41);
nor U57 (N_57,In_469,In_365);
nand U58 (N_58,In_306,In_681);
or U59 (N_59,In_552,In_370);
xor U60 (N_60,In_414,In_639);
xor U61 (N_61,In_44,In_675);
or U62 (N_62,In_734,In_516);
nand U63 (N_63,In_291,In_557);
and U64 (N_64,In_278,In_673);
and U65 (N_65,In_401,In_501);
and U66 (N_66,In_361,In_560);
nor U67 (N_67,In_139,In_30);
xnor U68 (N_68,In_104,In_117);
nand U69 (N_69,In_666,In_338);
nor U70 (N_70,In_252,In_607);
and U71 (N_71,In_313,In_415);
xnor U72 (N_72,In_280,In_668);
nor U73 (N_73,In_156,In_746);
nand U74 (N_74,In_679,In_27);
or U75 (N_75,In_707,In_91);
nor U76 (N_76,In_366,In_43);
xnor U77 (N_77,In_393,In_647);
nand U78 (N_78,In_284,In_118);
nor U79 (N_79,In_458,In_183);
and U80 (N_80,In_444,In_268);
xor U81 (N_81,In_641,In_287);
nand U82 (N_82,In_491,In_312);
nand U83 (N_83,In_224,In_193);
and U84 (N_84,In_346,In_7);
and U85 (N_85,In_194,In_598);
nor U86 (N_86,In_656,In_729);
or U87 (N_87,In_169,In_222);
nor U88 (N_88,In_64,In_396);
nand U89 (N_89,In_631,In_311);
nand U90 (N_90,In_724,In_201);
nand U91 (N_91,In_671,In_745);
nand U92 (N_92,In_217,In_163);
and U93 (N_93,In_723,In_12);
nor U94 (N_94,In_47,In_582);
nand U95 (N_95,In_29,In_680);
nand U96 (N_96,In_299,In_6);
or U97 (N_97,In_276,In_496);
and U98 (N_98,In_690,In_638);
or U99 (N_99,In_81,In_661);
nor U100 (N_100,In_604,In_561);
nor U101 (N_101,In_615,In_24);
nor U102 (N_102,In_479,In_520);
nand U103 (N_103,In_660,In_101);
nor U104 (N_104,In_472,In_97);
and U105 (N_105,In_428,In_733);
or U106 (N_106,In_102,In_328);
nand U107 (N_107,In_504,In_505);
nor U108 (N_108,In_713,In_630);
and U109 (N_109,In_152,In_612);
and U110 (N_110,In_134,In_403);
and U111 (N_111,In_227,In_556);
nor U112 (N_112,In_355,In_191);
xor U113 (N_113,In_674,In_305);
xor U114 (N_114,In_209,In_250);
or U115 (N_115,In_553,In_390);
nand U116 (N_116,In_712,In_480);
and U117 (N_117,In_292,In_275);
nand U118 (N_118,In_456,In_459);
or U119 (N_119,In_212,In_451);
or U120 (N_120,In_112,In_649);
or U121 (N_121,In_159,In_670);
xnor U122 (N_122,In_482,In_236);
xor U123 (N_123,In_92,In_643);
nor U124 (N_124,In_161,In_147);
xnor U125 (N_125,In_455,In_270);
nand U126 (N_126,In_709,In_315);
or U127 (N_127,In_283,In_636);
or U128 (N_128,In_61,In_135);
or U129 (N_129,In_144,In_543);
nand U130 (N_130,In_386,In_462);
nand U131 (N_131,In_42,In_143);
xnor U132 (N_132,In_699,In_231);
or U133 (N_133,In_544,In_88);
nor U134 (N_134,In_389,In_181);
nand U135 (N_135,In_533,In_411);
or U136 (N_136,In_378,In_277);
and U137 (N_137,In_345,In_63);
or U138 (N_138,In_199,In_547);
or U139 (N_139,In_317,In_175);
nand U140 (N_140,In_448,In_529);
and U141 (N_141,In_581,In_648);
and U142 (N_142,In_715,In_37);
and U143 (N_143,In_279,In_445);
or U144 (N_144,In_31,In_613);
xnor U145 (N_145,In_116,In_90);
xnor U146 (N_146,In_589,In_500);
nor U147 (N_147,In_34,In_294);
nand U148 (N_148,In_260,In_372);
xnor U149 (N_149,In_184,In_749);
or U150 (N_150,In_423,In_473);
xnor U151 (N_151,In_524,In_196);
xor U152 (N_152,In_457,In_137);
nand U153 (N_153,In_66,In_190);
nor U154 (N_154,In_710,In_129);
and U155 (N_155,In_575,In_629);
and U156 (N_156,In_512,In_39);
and U157 (N_157,In_281,In_293);
or U158 (N_158,In_329,In_515);
and U159 (N_159,In_301,In_410);
or U160 (N_160,In_421,In_453);
nand U161 (N_161,In_628,In_341);
nor U162 (N_162,In_700,In_172);
nand U163 (N_163,In_464,In_447);
xnor U164 (N_164,In_449,In_171);
nor U165 (N_165,In_46,In_157);
nand U166 (N_166,In_702,In_214);
xnor U167 (N_167,In_461,In_611);
and U168 (N_168,In_22,In_667);
or U169 (N_169,In_375,In_228);
and U170 (N_170,In_593,In_634);
and U171 (N_171,In_158,In_692);
and U172 (N_172,In_71,In_85);
and U173 (N_173,In_651,In_166);
nor U174 (N_174,In_371,In_237);
nor U175 (N_175,In_337,In_110);
nor U176 (N_176,In_258,In_600);
or U177 (N_177,In_331,In_587);
nand U178 (N_178,In_332,In_207);
xor U179 (N_179,In_736,In_554);
xor U180 (N_180,In_2,In_488);
and U181 (N_181,In_506,In_694);
nor U182 (N_182,In_94,In_417);
or U183 (N_183,In_99,In_597);
xnor U184 (N_184,In_36,In_610);
or U185 (N_185,In_669,In_528);
nand U186 (N_186,In_640,In_48);
nor U187 (N_187,In_206,In_717);
xor U188 (N_188,In_369,In_264);
xnor U189 (N_189,In_87,In_664);
or U190 (N_190,In_632,In_436);
and U191 (N_191,In_503,In_507);
xor U192 (N_192,In_525,In_186);
nor U193 (N_193,In_510,In_398);
xor U194 (N_194,In_16,In_606);
or U195 (N_195,In_77,In_427);
or U196 (N_196,In_443,In_492);
nor U197 (N_197,In_165,In_246);
or U198 (N_198,In_49,In_83);
nor U199 (N_199,In_602,In_19);
nand U200 (N_200,In_153,N_104);
nand U201 (N_201,In_1,In_558);
and U202 (N_202,N_11,N_33);
xnor U203 (N_203,N_58,N_181);
and U204 (N_204,In_54,In_40);
and U205 (N_205,In_140,N_121);
nand U206 (N_206,In_573,In_578);
nand U207 (N_207,In_617,N_101);
or U208 (N_208,In_477,N_138);
nand U209 (N_209,N_142,N_32);
nand U210 (N_210,N_197,In_550);
and U211 (N_211,In_590,In_367);
or U212 (N_212,In_383,In_204);
or U213 (N_213,N_51,In_684);
or U214 (N_214,In_714,In_652);
and U215 (N_215,In_619,In_15);
or U216 (N_216,In_425,N_196);
xnor U217 (N_217,In_321,N_114);
nor U218 (N_218,N_30,In_327);
xnor U219 (N_219,N_157,In_385);
nand U220 (N_220,In_256,In_576);
nor U221 (N_221,In_314,N_69);
nand U222 (N_222,In_359,In_266);
xor U223 (N_223,In_435,In_405);
nand U224 (N_224,In_122,In_689);
xor U225 (N_225,N_98,In_654);
xor U226 (N_226,In_526,N_49);
or U227 (N_227,In_218,N_74);
xor U228 (N_228,N_131,In_376);
and U229 (N_229,In_303,In_391);
nor U230 (N_230,N_174,In_722);
and U231 (N_231,N_110,In_397);
nor U232 (N_232,In_420,In_719);
xnor U233 (N_233,In_518,In_562);
nor U234 (N_234,N_40,N_7);
nor U235 (N_235,In_55,In_551);
nor U236 (N_236,In_123,In_434);
and U237 (N_237,In_253,N_171);
and U238 (N_238,N_0,N_77);
nand U239 (N_239,In_586,N_168);
and U240 (N_240,N_128,In_426);
nor U241 (N_241,In_718,In_180);
nand U242 (N_242,N_78,In_229);
xnor U243 (N_243,In_234,In_200);
nand U244 (N_244,N_141,In_693);
xnor U245 (N_245,In_5,In_394);
xnor U246 (N_246,In_580,In_211);
nor U247 (N_247,In_716,N_154);
xor U248 (N_248,N_45,In_72);
nand U249 (N_249,In_45,N_14);
xor U250 (N_250,In_485,N_107);
or U251 (N_251,In_441,In_537);
and U252 (N_252,N_34,N_184);
nor U253 (N_253,N_10,In_62);
or U254 (N_254,In_571,N_54);
and U255 (N_255,N_190,In_514);
nand U256 (N_256,In_463,In_340);
and U257 (N_257,In_164,N_70);
and U258 (N_258,N_28,In_4);
or U259 (N_259,N_176,In_170);
xnor U260 (N_260,In_381,N_115);
or U261 (N_261,N_80,N_135);
xnor U262 (N_262,In_637,In_254);
nor U263 (N_263,N_130,N_60);
xnor U264 (N_264,N_66,In_744);
or U265 (N_265,In_142,N_47);
and U266 (N_266,In_614,In_646);
nand U267 (N_267,In_265,N_59);
xnor U268 (N_268,In_82,N_136);
nor U269 (N_269,In_730,In_263);
or U270 (N_270,In_95,N_170);
nor U271 (N_271,In_659,N_3);
nor U272 (N_272,N_86,N_120);
xor U273 (N_273,In_687,In_644);
nor U274 (N_274,N_188,N_93);
nand U275 (N_275,N_162,In_430);
or U276 (N_276,In_395,In_297);
nor U277 (N_277,In_523,N_84);
or U278 (N_278,N_29,In_96);
and U279 (N_279,In_167,In_347);
or U280 (N_280,N_56,In_356);
xnor U281 (N_281,N_38,In_555);
nor U282 (N_282,In_145,N_92);
nand U283 (N_283,In_618,N_22);
nor U284 (N_284,In_616,In_216);
xnor U285 (N_285,N_106,In_242);
and U286 (N_286,In_563,In_498);
nor U287 (N_287,In_56,In_353);
nand U288 (N_288,In_584,In_665);
nor U289 (N_289,In_363,N_150);
or U290 (N_290,In_79,In_698);
and U291 (N_291,In_261,N_76);
nand U292 (N_292,In_50,In_133);
and U293 (N_293,In_706,N_52);
and U294 (N_294,In_128,In_678);
and U295 (N_295,In_362,In_316);
nand U296 (N_296,In_352,In_682);
or U297 (N_297,In_522,N_159);
and U298 (N_298,N_20,In_65);
nor U299 (N_299,N_177,In_400);
nor U300 (N_300,In_267,In_742);
and U301 (N_301,In_705,N_12);
and U302 (N_302,In_138,In_304);
and U303 (N_303,In_330,In_18);
xnor U304 (N_304,In_703,In_245);
nand U305 (N_305,N_102,In_596);
and U306 (N_306,N_36,N_149);
xor U307 (N_307,In_454,In_499);
xor U308 (N_308,In_273,In_422);
or U309 (N_309,In_146,In_536);
nand U310 (N_310,In_565,In_534);
nand U311 (N_311,N_193,In_662);
nor U312 (N_312,In_549,N_25);
nand U313 (N_313,N_160,In_188);
and U314 (N_314,In_296,In_380);
xnor U315 (N_315,In_697,In_348);
nor U316 (N_316,N_48,In_141);
xnor U317 (N_317,In_308,N_180);
nor U318 (N_318,N_17,In_259);
xor U319 (N_319,In_302,In_178);
or U320 (N_320,N_97,N_195);
and U321 (N_321,In_384,In_708);
nor U322 (N_322,In_148,In_255);
and U323 (N_323,In_620,In_120);
nand U324 (N_324,N_63,In_579);
nand U325 (N_325,In_559,N_155);
nor U326 (N_326,In_354,In_603);
xor U327 (N_327,In_334,In_272);
or U328 (N_328,In_645,N_26);
and U329 (N_329,In_197,In_676);
nor U330 (N_330,In_75,In_475);
or U331 (N_331,In_609,N_89);
and U332 (N_332,In_650,In_233);
or U333 (N_333,In_271,In_151);
xnor U334 (N_334,In_368,N_82);
and U335 (N_335,N_143,In_221);
nand U336 (N_336,N_140,In_731);
nor U337 (N_337,N_39,In_203);
xnor U338 (N_338,In_223,N_153);
or U339 (N_339,N_178,In_309);
or U340 (N_340,In_235,In_106);
xor U341 (N_341,N_173,N_116);
and U342 (N_342,In_10,N_156);
and U343 (N_343,N_88,N_112);
nor U344 (N_344,In_238,N_1);
nor U345 (N_345,N_182,In_226);
xor U346 (N_346,N_132,In_595);
nor U347 (N_347,In_215,In_300);
xnor U348 (N_348,In_350,N_194);
or U349 (N_349,N_43,N_44);
xnor U350 (N_350,In_80,N_64);
and U351 (N_351,In_74,N_172);
or U352 (N_352,In_20,N_175);
or U353 (N_353,In_546,In_726);
and U354 (N_354,In_32,In_377);
and U355 (N_355,In_68,In_73);
or U356 (N_356,In_591,N_105);
or U357 (N_357,N_13,N_109);
nor U358 (N_358,In_406,In_9);
nand U359 (N_359,N_161,In_132);
xnor U360 (N_360,In_530,In_439);
nand U361 (N_361,N_96,In_509);
nor U362 (N_362,In_538,In_288);
or U363 (N_363,In_735,In_623);
nor U364 (N_364,In_257,In_704);
or U365 (N_365,N_15,N_99);
nand U366 (N_366,N_133,N_152);
and U367 (N_367,In_173,In_239);
nand U368 (N_368,N_53,In_360);
nor U369 (N_369,In_322,In_683);
nand U370 (N_370,In_740,In_732);
nand U371 (N_371,In_379,In_519);
xor U372 (N_372,In_489,In_569);
xnor U373 (N_373,In_105,N_124);
and U374 (N_374,In_225,In_67);
or U375 (N_375,In_494,N_179);
xnor U376 (N_376,In_663,In_107);
nor U377 (N_377,N_147,In_243);
xor U378 (N_378,In_13,N_166);
nand U379 (N_379,In_285,N_24);
or U380 (N_380,In_446,In_53);
nor U381 (N_381,N_119,N_91);
nor U382 (N_382,N_55,In_111);
nor U383 (N_383,In_382,In_695);
xnor U384 (N_384,In_517,In_688);
and U385 (N_385,N_95,N_35);
xor U386 (N_386,In_653,N_8);
xnor U387 (N_387,In_344,In_100);
xor U388 (N_388,In_160,In_601);
or U389 (N_389,N_163,N_169);
or U390 (N_390,In_424,N_31);
nand U391 (N_391,In_325,In_205);
nor U392 (N_392,In_60,N_62);
and U393 (N_393,N_73,N_61);
xor U394 (N_394,In_437,In_511);
nand U395 (N_395,N_94,N_118);
xor U396 (N_396,In_251,In_685);
and U397 (N_397,In_23,In_481);
or U398 (N_398,N_192,N_125);
or U399 (N_399,In_262,N_71);
and U400 (N_400,N_275,In_633);
xnor U401 (N_401,In_419,N_222);
nand U402 (N_402,N_364,N_151);
nand U403 (N_403,In_21,N_282);
xnor U404 (N_404,N_234,In_109);
xnor U405 (N_405,In_513,N_388);
xor U406 (N_406,N_345,N_23);
nand U407 (N_407,N_271,N_341);
nor U408 (N_408,N_200,N_272);
and U409 (N_409,N_268,In_8);
nand U410 (N_410,N_42,N_185);
xor U411 (N_411,In_452,N_209);
and U412 (N_412,N_90,N_122);
xnor U413 (N_413,N_329,In_696);
or U414 (N_414,In_655,N_238);
nand U415 (N_415,N_321,N_219);
xnor U416 (N_416,N_213,N_251);
and U417 (N_417,N_214,N_318);
and U418 (N_418,N_376,In_409);
nor U419 (N_419,In_58,N_306);
and U420 (N_420,N_396,N_134);
nor U421 (N_421,N_87,N_229);
nand U422 (N_422,N_385,N_370);
nand U423 (N_423,In_531,N_375);
or U424 (N_424,In_470,N_242);
nand U425 (N_425,N_41,In_349);
xor U426 (N_426,N_247,N_239);
nand U427 (N_427,N_303,N_146);
nand U428 (N_428,In_431,In_438);
xnor U429 (N_429,N_381,In_465);
nand U430 (N_430,In_69,N_354);
and U431 (N_431,N_46,N_338);
nand U432 (N_432,In_333,N_186);
and U433 (N_433,N_85,N_217);
and U434 (N_434,N_260,In_487);
xnor U435 (N_435,N_313,In_25);
nand U436 (N_436,N_395,N_212);
or U437 (N_437,N_108,N_248);
nor U438 (N_438,N_391,N_335);
and U439 (N_439,N_337,N_202);
nand U440 (N_440,In_208,N_397);
or U441 (N_441,In_198,In_566);
xnor U442 (N_442,N_349,In_626);
and U443 (N_443,N_334,N_252);
nor U444 (N_444,N_231,N_283);
nor U445 (N_445,N_264,N_265);
and U446 (N_446,N_286,N_294);
xor U447 (N_447,N_358,N_75);
nor U448 (N_448,In_339,N_355);
nand U449 (N_449,N_123,In_727);
and U450 (N_450,In_131,N_368);
nor U451 (N_451,N_399,N_220);
or U452 (N_452,N_332,N_333);
nand U453 (N_453,N_81,N_386);
nand U454 (N_454,N_393,In_635);
or U455 (N_455,N_317,N_221);
or U456 (N_456,N_280,N_266);
nor U457 (N_457,In_125,N_79);
nand U458 (N_458,N_249,N_372);
nand U459 (N_459,N_225,N_244);
xnor U460 (N_460,N_320,N_201);
xor U461 (N_461,N_274,In_342);
nor U462 (N_462,N_256,N_276);
or U463 (N_463,In_17,N_206);
nor U464 (N_464,N_339,N_346);
nand U465 (N_465,In_476,N_218);
and U466 (N_466,N_211,In_154);
or U467 (N_467,N_293,N_309);
nor U468 (N_468,N_316,In_478);
nand U469 (N_469,N_240,N_191);
nand U470 (N_470,In_114,N_285);
nor U471 (N_471,In_179,N_351);
and U472 (N_472,N_67,N_258);
nor U473 (N_473,In_168,N_279);
xnor U474 (N_474,In_432,In_577);
and U475 (N_475,N_224,N_288);
xor U476 (N_476,N_254,N_137);
nand U477 (N_477,In_210,N_352);
nand U478 (N_478,N_127,N_227);
or U479 (N_479,In_725,N_6);
and U480 (N_480,In_240,N_284);
xor U481 (N_481,In_542,In_177);
or U482 (N_482,N_362,In_605);
and U483 (N_483,N_199,N_148);
or U484 (N_484,N_325,N_232);
nand U485 (N_485,In_220,N_365);
or U486 (N_486,N_322,N_374);
nand U487 (N_487,N_295,N_298);
xor U488 (N_488,N_366,N_236);
or U489 (N_489,In_336,N_72);
and U490 (N_490,In_627,In_658);
or U491 (N_491,N_257,N_287);
or U492 (N_492,N_237,In_52);
or U493 (N_493,N_111,N_245);
or U494 (N_494,In_136,In_588);
xnor U495 (N_495,N_347,In_3);
nor U496 (N_496,In_298,N_331);
xnor U497 (N_497,N_302,N_378);
nor U498 (N_498,N_367,N_83);
and U499 (N_499,N_241,N_19);
xnor U500 (N_500,In_155,N_126);
xor U501 (N_501,In_108,N_304);
or U502 (N_502,In_28,N_319);
or U503 (N_503,N_198,N_246);
or U504 (N_504,N_360,N_250);
and U505 (N_505,N_369,In_483);
and U506 (N_506,N_259,N_330);
xor U507 (N_507,In_486,N_139);
or U508 (N_508,N_310,N_103);
nand U509 (N_509,N_327,N_216);
or U510 (N_510,N_363,N_357);
xnor U511 (N_511,N_394,N_392);
and U512 (N_512,N_299,N_314);
nor U513 (N_513,N_340,N_183);
xor U514 (N_514,N_300,N_65);
xnor U515 (N_515,N_380,In_450);
xnor U516 (N_516,In_440,N_223);
and U517 (N_517,N_27,N_379);
nand U518 (N_518,N_292,N_50);
nand U519 (N_519,N_16,In_672);
nor U520 (N_520,N_113,N_291);
nand U521 (N_521,N_297,N_4);
nor U522 (N_522,N_9,N_311);
or U523 (N_523,N_312,In_248);
or U524 (N_524,In_583,N_117);
or U525 (N_525,In_103,N_208);
nor U526 (N_526,N_371,In_249);
nand U527 (N_527,N_289,In_677);
or U528 (N_528,In_326,In_621);
nand U529 (N_529,N_144,N_305);
nor U530 (N_530,N_384,N_390);
nor U531 (N_531,N_145,N_187);
nor U532 (N_532,N_315,N_307);
or U533 (N_533,In_599,N_129);
nor U534 (N_534,N_255,N_207);
nor U535 (N_535,In_244,N_205);
xor U536 (N_536,N_100,N_344);
or U537 (N_537,N_57,N_210);
xor U538 (N_538,N_228,N_164);
and U539 (N_539,N_204,N_353);
nor U540 (N_540,In_412,N_262);
nor U541 (N_541,N_203,N_243);
or U542 (N_542,N_382,N_267);
nand U543 (N_543,N_270,In_14);
and U544 (N_544,N_281,In_86);
xnor U545 (N_545,N_373,N_278);
or U546 (N_546,N_2,In_387);
and U547 (N_547,N_308,N_273);
nand U548 (N_548,In_474,N_359);
and U549 (N_549,In_289,In_323);
xor U550 (N_550,In_35,N_389);
nor U551 (N_551,In_502,N_167);
nor U552 (N_552,N_68,N_324);
nor U553 (N_553,N_277,N_230);
nor U554 (N_554,N_165,N_253);
nand U555 (N_555,N_343,N_328);
nand U556 (N_556,In_51,N_5);
xor U557 (N_557,N_37,In_686);
nor U558 (N_558,N_356,N_377);
xnor U559 (N_559,N_21,In_286);
or U560 (N_560,N_301,In_416);
or U561 (N_561,N_233,N_158);
xnor U562 (N_562,N_323,N_269);
and U563 (N_563,N_235,In_471);
and U564 (N_564,N_226,N_350);
nor U565 (N_565,N_348,In_274);
nand U566 (N_566,N_290,In_747);
and U567 (N_567,In_351,N_215);
nor U568 (N_568,N_261,N_18);
nor U569 (N_569,N_336,N_383);
nand U570 (N_570,In_93,N_387);
nand U571 (N_571,N_342,N_398);
nand U572 (N_572,N_296,N_361);
and U573 (N_573,N_189,In_343);
xnor U574 (N_574,N_326,N_263);
and U575 (N_575,N_200,N_288);
xnor U576 (N_576,In_696,In_621);
or U577 (N_577,N_252,N_211);
and U578 (N_578,N_340,N_284);
nand U579 (N_579,N_351,N_238);
or U580 (N_580,N_325,N_240);
nand U581 (N_581,In_486,N_90);
and U582 (N_582,In_93,In_412);
or U583 (N_583,N_398,N_284);
and U584 (N_584,N_307,N_267);
xor U585 (N_585,N_392,In_336);
nand U586 (N_586,N_277,N_385);
or U587 (N_587,N_293,N_367);
or U588 (N_588,N_368,N_233);
and U589 (N_589,N_348,In_513);
nor U590 (N_590,N_286,N_382);
or U591 (N_591,N_258,In_471);
nand U592 (N_592,N_228,N_295);
and U593 (N_593,N_198,N_226);
or U594 (N_594,N_372,N_343);
xnor U595 (N_595,In_432,N_240);
nand U596 (N_596,In_339,In_483);
xnor U597 (N_597,In_108,N_301);
and U598 (N_598,N_83,In_583);
nand U599 (N_599,N_376,N_335);
xnor U600 (N_600,N_419,N_463);
nor U601 (N_601,N_543,N_451);
and U602 (N_602,N_412,N_559);
xnor U603 (N_603,N_465,N_420);
or U604 (N_604,N_525,N_539);
nor U605 (N_605,N_427,N_480);
nor U606 (N_606,N_566,N_404);
and U607 (N_607,N_552,N_501);
or U608 (N_608,N_514,N_584);
or U609 (N_609,N_569,N_400);
nand U610 (N_610,N_577,N_503);
and U611 (N_611,N_493,N_567);
xor U612 (N_612,N_578,N_441);
nor U613 (N_613,N_547,N_401);
xnor U614 (N_614,N_479,N_452);
nand U615 (N_615,N_505,N_496);
xnor U616 (N_616,N_495,N_408);
xnor U617 (N_617,N_599,N_423);
xor U618 (N_618,N_548,N_529);
or U619 (N_619,N_520,N_435);
xnor U620 (N_620,N_518,N_580);
nand U621 (N_621,N_475,N_593);
nor U622 (N_622,N_524,N_522);
nor U623 (N_623,N_574,N_464);
and U624 (N_624,N_512,N_424);
nor U625 (N_625,N_414,N_570);
and U626 (N_626,N_575,N_540);
xnor U627 (N_627,N_489,N_516);
xnor U628 (N_628,N_447,N_549);
xor U629 (N_629,N_571,N_486);
or U630 (N_630,N_587,N_532);
nor U631 (N_631,N_487,N_418);
nor U632 (N_632,N_494,N_429);
and U633 (N_633,N_530,N_483);
xor U634 (N_634,N_541,N_588);
and U635 (N_635,N_519,N_406);
nor U636 (N_636,N_572,N_476);
and U637 (N_637,N_582,N_568);
or U638 (N_638,N_513,N_542);
or U639 (N_639,N_498,N_473);
nor U640 (N_640,N_500,N_443);
and U641 (N_641,N_597,N_554);
nor U642 (N_642,N_407,N_560);
nor U643 (N_643,N_477,N_523);
and U644 (N_644,N_482,N_453);
nor U645 (N_645,N_478,N_573);
or U646 (N_646,N_491,N_507);
xor U647 (N_647,N_576,N_590);
or U648 (N_648,N_426,N_425);
or U649 (N_649,N_469,N_508);
xor U650 (N_650,N_490,N_434);
or U651 (N_651,N_460,N_448);
xnor U652 (N_652,N_504,N_485);
xnor U653 (N_653,N_545,N_416);
xnor U654 (N_654,N_538,N_413);
and U655 (N_655,N_563,N_442);
nand U656 (N_656,N_446,N_585);
nor U657 (N_657,N_517,N_431);
nand U658 (N_658,N_594,N_555);
and U659 (N_659,N_468,N_439);
xnor U660 (N_660,N_484,N_449);
or U661 (N_661,N_546,N_428);
nand U662 (N_662,N_564,N_565);
nand U663 (N_663,N_461,N_438);
and U664 (N_664,N_402,N_528);
nand U665 (N_665,N_596,N_430);
nor U666 (N_666,N_506,N_492);
nor U667 (N_667,N_561,N_415);
xnor U668 (N_668,N_527,N_422);
nand U669 (N_669,N_433,N_474);
nor U670 (N_670,N_445,N_531);
nor U671 (N_671,N_511,N_456);
nand U672 (N_672,N_437,N_544);
and U673 (N_673,N_521,N_470);
nor U674 (N_674,N_455,N_450);
nand U675 (N_675,N_466,N_497);
or U676 (N_676,N_592,N_579);
or U677 (N_677,N_556,N_515);
nor U678 (N_678,N_410,N_403);
and U679 (N_679,N_467,N_454);
nor U680 (N_680,N_509,N_499);
nand U681 (N_681,N_583,N_589);
nor U682 (N_682,N_457,N_458);
xor U683 (N_683,N_502,N_472);
nor U684 (N_684,N_510,N_421);
nor U685 (N_685,N_586,N_411);
and U686 (N_686,N_440,N_536);
xor U687 (N_687,N_558,N_591);
and U688 (N_688,N_557,N_459);
or U689 (N_689,N_534,N_551);
nor U690 (N_690,N_444,N_595);
nand U691 (N_691,N_417,N_488);
nand U692 (N_692,N_553,N_436);
nor U693 (N_693,N_526,N_432);
and U694 (N_694,N_405,N_550);
nor U695 (N_695,N_462,N_471);
xnor U696 (N_696,N_537,N_409);
and U697 (N_697,N_598,N_481);
nand U698 (N_698,N_535,N_562);
nand U699 (N_699,N_533,N_581);
xnor U700 (N_700,N_491,N_419);
nor U701 (N_701,N_567,N_424);
xor U702 (N_702,N_561,N_485);
or U703 (N_703,N_591,N_429);
nor U704 (N_704,N_454,N_571);
nand U705 (N_705,N_561,N_490);
and U706 (N_706,N_523,N_575);
nor U707 (N_707,N_400,N_461);
nor U708 (N_708,N_559,N_405);
and U709 (N_709,N_454,N_551);
and U710 (N_710,N_447,N_561);
nand U711 (N_711,N_549,N_455);
nand U712 (N_712,N_523,N_433);
nor U713 (N_713,N_406,N_517);
xnor U714 (N_714,N_472,N_546);
or U715 (N_715,N_530,N_403);
and U716 (N_716,N_460,N_471);
nand U717 (N_717,N_467,N_428);
and U718 (N_718,N_526,N_454);
nand U719 (N_719,N_501,N_492);
nand U720 (N_720,N_569,N_537);
and U721 (N_721,N_564,N_450);
xnor U722 (N_722,N_439,N_465);
nor U723 (N_723,N_519,N_427);
nor U724 (N_724,N_481,N_412);
or U725 (N_725,N_436,N_536);
nand U726 (N_726,N_491,N_476);
nor U727 (N_727,N_458,N_427);
or U728 (N_728,N_465,N_539);
and U729 (N_729,N_512,N_568);
nand U730 (N_730,N_505,N_519);
or U731 (N_731,N_573,N_493);
nand U732 (N_732,N_570,N_448);
nand U733 (N_733,N_450,N_460);
or U734 (N_734,N_426,N_489);
or U735 (N_735,N_425,N_565);
and U736 (N_736,N_557,N_400);
nand U737 (N_737,N_415,N_516);
and U738 (N_738,N_448,N_528);
nor U739 (N_739,N_496,N_405);
or U740 (N_740,N_441,N_579);
or U741 (N_741,N_584,N_427);
nor U742 (N_742,N_458,N_476);
xor U743 (N_743,N_509,N_429);
xor U744 (N_744,N_482,N_418);
xor U745 (N_745,N_490,N_533);
and U746 (N_746,N_556,N_485);
or U747 (N_747,N_412,N_443);
xnor U748 (N_748,N_451,N_489);
or U749 (N_749,N_500,N_433);
xnor U750 (N_750,N_528,N_574);
xor U751 (N_751,N_557,N_513);
and U752 (N_752,N_409,N_527);
nor U753 (N_753,N_594,N_465);
and U754 (N_754,N_484,N_587);
xnor U755 (N_755,N_425,N_400);
nor U756 (N_756,N_405,N_519);
nor U757 (N_757,N_536,N_435);
nand U758 (N_758,N_469,N_491);
nand U759 (N_759,N_484,N_573);
nor U760 (N_760,N_448,N_462);
nor U761 (N_761,N_415,N_403);
and U762 (N_762,N_482,N_425);
or U763 (N_763,N_578,N_486);
and U764 (N_764,N_509,N_425);
or U765 (N_765,N_558,N_462);
and U766 (N_766,N_497,N_567);
nor U767 (N_767,N_572,N_539);
and U768 (N_768,N_478,N_428);
or U769 (N_769,N_404,N_553);
xnor U770 (N_770,N_486,N_549);
nor U771 (N_771,N_572,N_485);
nand U772 (N_772,N_527,N_504);
and U773 (N_773,N_538,N_483);
or U774 (N_774,N_479,N_418);
or U775 (N_775,N_419,N_598);
nand U776 (N_776,N_553,N_502);
or U777 (N_777,N_515,N_462);
nor U778 (N_778,N_458,N_510);
nor U779 (N_779,N_569,N_452);
xor U780 (N_780,N_588,N_409);
nor U781 (N_781,N_575,N_425);
xor U782 (N_782,N_454,N_490);
xnor U783 (N_783,N_522,N_433);
xor U784 (N_784,N_533,N_465);
or U785 (N_785,N_439,N_448);
xor U786 (N_786,N_523,N_423);
or U787 (N_787,N_573,N_477);
or U788 (N_788,N_527,N_480);
and U789 (N_789,N_506,N_451);
nand U790 (N_790,N_486,N_454);
and U791 (N_791,N_516,N_544);
or U792 (N_792,N_525,N_535);
xnor U793 (N_793,N_596,N_553);
nand U794 (N_794,N_430,N_553);
xor U795 (N_795,N_506,N_586);
nand U796 (N_796,N_556,N_449);
and U797 (N_797,N_554,N_483);
nand U798 (N_798,N_426,N_473);
and U799 (N_799,N_538,N_514);
nand U800 (N_800,N_682,N_742);
xor U801 (N_801,N_782,N_781);
and U802 (N_802,N_620,N_777);
nor U803 (N_803,N_731,N_791);
or U804 (N_804,N_656,N_732);
xor U805 (N_805,N_765,N_679);
xor U806 (N_806,N_717,N_683);
xnor U807 (N_807,N_621,N_726);
nand U808 (N_808,N_737,N_647);
nand U809 (N_809,N_667,N_658);
and U810 (N_810,N_728,N_660);
nand U811 (N_811,N_626,N_624);
or U812 (N_812,N_652,N_609);
nor U813 (N_813,N_629,N_794);
nor U814 (N_814,N_696,N_670);
or U815 (N_815,N_720,N_604);
nand U816 (N_816,N_659,N_723);
or U817 (N_817,N_741,N_648);
or U818 (N_818,N_778,N_740);
or U819 (N_819,N_730,N_617);
and U820 (N_820,N_774,N_603);
and U821 (N_821,N_691,N_719);
or U822 (N_822,N_722,N_690);
or U823 (N_823,N_702,N_795);
nor U824 (N_824,N_637,N_650);
and U825 (N_825,N_628,N_661);
or U826 (N_826,N_779,N_693);
xnor U827 (N_827,N_642,N_640);
nor U828 (N_828,N_615,N_664);
nand U829 (N_829,N_789,N_706);
nand U830 (N_830,N_799,N_767);
and U831 (N_831,N_770,N_733);
xor U832 (N_832,N_766,N_668);
xor U833 (N_833,N_713,N_738);
and U834 (N_834,N_694,N_687);
xor U835 (N_835,N_748,N_669);
nor U836 (N_836,N_712,N_688);
nor U837 (N_837,N_707,N_635);
xnor U838 (N_838,N_752,N_747);
xor U839 (N_839,N_716,N_756);
xnor U840 (N_840,N_769,N_797);
xnor U841 (N_841,N_784,N_763);
nor U842 (N_842,N_704,N_677);
and U843 (N_843,N_714,N_721);
nor U844 (N_844,N_735,N_689);
nor U845 (N_845,N_655,N_753);
nand U846 (N_846,N_708,N_645);
and U847 (N_847,N_783,N_773);
and U848 (N_848,N_625,N_649);
and U849 (N_849,N_772,N_798);
or U850 (N_850,N_644,N_618);
or U851 (N_851,N_684,N_725);
nand U852 (N_852,N_760,N_759);
nand U853 (N_853,N_605,N_703);
or U854 (N_854,N_715,N_698);
xor U855 (N_855,N_646,N_602);
and U856 (N_856,N_734,N_608);
nor U857 (N_857,N_768,N_739);
nand U858 (N_858,N_600,N_744);
and U859 (N_859,N_622,N_710);
nor U860 (N_860,N_787,N_727);
nand U861 (N_861,N_671,N_699);
xor U862 (N_862,N_627,N_654);
nor U863 (N_863,N_750,N_662);
or U864 (N_864,N_641,N_672);
nor U865 (N_865,N_634,N_745);
xor U866 (N_866,N_754,N_631);
nor U867 (N_867,N_709,N_610);
nor U868 (N_868,N_638,N_601);
and U869 (N_869,N_633,N_729);
and U870 (N_870,N_632,N_607);
and U871 (N_871,N_757,N_743);
nor U872 (N_872,N_780,N_612);
nand U873 (N_873,N_705,N_619);
xnor U874 (N_874,N_636,N_674);
nand U875 (N_875,N_630,N_724);
xnor U876 (N_876,N_786,N_746);
nor U877 (N_877,N_758,N_790);
nand U878 (N_878,N_675,N_685);
nor U879 (N_879,N_695,N_749);
or U880 (N_880,N_711,N_614);
xnor U881 (N_881,N_616,N_657);
nor U882 (N_882,N_764,N_611);
nor U883 (N_883,N_623,N_775);
or U884 (N_884,N_686,N_736);
nand U885 (N_885,N_613,N_681);
xnor U886 (N_886,N_663,N_701);
and U887 (N_887,N_792,N_665);
or U888 (N_888,N_776,N_697);
xnor U889 (N_889,N_751,N_678);
nand U890 (N_890,N_606,N_666);
nor U891 (N_891,N_762,N_643);
nor U892 (N_892,N_761,N_718);
nand U893 (N_893,N_651,N_700);
and U894 (N_894,N_673,N_793);
or U895 (N_895,N_785,N_788);
and U896 (N_896,N_680,N_692);
xnor U897 (N_897,N_639,N_653);
nor U898 (N_898,N_676,N_796);
xor U899 (N_899,N_771,N_755);
and U900 (N_900,N_779,N_753);
nor U901 (N_901,N_655,N_799);
nor U902 (N_902,N_756,N_670);
nor U903 (N_903,N_652,N_650);
or U904 (N_904,N_757,N_734);
xor U905 (N_905,N_636,N_782);
nor U906 (N_906,N_696,N_788);
xnor U907 (N_907,N_650,N_717);
nor U908 (N_908,N_658,N_681);
nand U909 (N_909,N_602,N_708);
xnor U910 (N_910,N_602,N_719);
xnor U911 (N_911,N_650,N_606);
xnor U912 (N_912,N_692,N_641);
or U913 (N_913,N_636,N_756);
or U914 (N_914,N_794,N_703);
and U915 (N_915,N_618,N_702);
or U916 (N_916,N_795,N_676);
and U917 (N_917,N_687,N_654);
and U918 (N_918,N_719,N_775);
nand U919 (N_919,N_701,N_665);
nor U920 (N_920,N_629,N_718);
and U921 (N_921,N_694,N_708);
nor U922 (N_922,N_772,N_633);
and U923 (N_923,N_736,N_637);
or U924 (N_924,N_693,N_627);
nor U925 (N_925,N_603,N_634);
or U926 (N_926,N_647,N_744);
and U927 (N_927,N_605,N_676);
or U928 (N_928,N_774,N_765);
or U929 (N_929,N_606,N_603);
xnor U930 (N_930,N_651,N_646);
and U931 (N_931,N_609,N_797);
and U932 (N_932,N_786,N_633);
and U933 (N_933,N_612,N_770);
nor U934 (N_934,N_738,N_720);
or U935 (N_935,N_796,N_773);
and U936 (N_936,N_602,N_690);
nor U937 (N_937,N_765,N_664);
xor U938 (N_938,N_748,N_682);
nor U939 (N_939,N_708,N_674);
nor U940 (N_940,N_647,N_792);
and U941 (N_941,N_704,N_771);
nor U942 (N_942,N_736,N_643);
xnor U943 (N_943,N_670,N_664);
or U944 (N_944,N_703,N_609);
and U945 (N_945,N_722,N_736);
nand U946 (N_946,N_740,N_607);
nor U947 (N_947,N_795,N_772);
nand U948 (N_948,N_770,N_781);
nand U949 (N_949,N_675,N_673);
and U950 (N_950,N_786,N_626);
and U951 (N_951,N_667,N_774);
nor U952 (N_952,N_608,N_787);
or U953 (N_953,N_741,N_698);
nor U954 (N_954,N_688,N_691);
nor U955 (N_955,N_754,N_662);
nand U956 (N_956,N_731,N_655);
xnor U957 (N_957,N_697,N_623);
nor U958 (N_958,N_737,N_664);
nand U959 (N_959,N_640,N_631);
nand U960 (N_960,N_746,N_651);
nor U961 (N_961,N_770,N_737);
xor U962 (N_962,N_753,N_771);
nand U963 (N_963,N_638,N_768);
nor U964 (N_964,N_739,N_694);
or U965 (N_965,N_750,N_710);
and U966 (N_966,N_741,N_691);
nand U967 (N_967,N_782,N_758);
nor U968 (N_968,N_619,N_724);
and U969 (N_969,N_740,N_741);
and U970 (N_970,N_772,N_648);
xor U971 (N_971,N_765,N_696);
nand U972 (N_972,N_686,N_675);
xnor U973 (N_973,N_780,N_763);
nor U974 (N_974,N_625,N_747);
nand U975 (N_975,N_638,N_647);
nor U976 (N_976,N_723,N_728);
nand U977 (N_977,N_729,N_632);
or U978 (N_978,N_695,N_780);
xnor U979 (N_979,N_749,N_628);
or U980 (N_980,N_654,N_600);
nand U981 (N_981,N_603,N_751);
and U982 (N_982,N_608,N_601);
nand U983 (N_983,N_677,N_612);
nand U984 (N_984,N_624,N_752);
nand U985 (N_985,N_721,N_689);
or U986 (N_986,N_743,N_791);
or U987 (N_987,N_619,N_740);
nand U988 (N_988,N_724,N_720);
and U989 (N_989,N_641,N_788);
xor U990 (N_990,N_755,N_750);
or U991 (N_991,N_673,N_742);
or U992 (N_992,N_734,N_642);
and U993 (N_993,N_607,N_644);
or U994 (N_994,N_634,N_706);
nand U995 (N_995,N_635,N_628);
xnor U996 (N_996,N_666,N_766);
xor U997 (N_997,N_785,N_730);
xnor U998 (N_998,N_679,N_760);
nand U999 (N_999,N_764,N_695);
nor U1000 (N_1000,N_814,N_808);
nand U1001 (N_1001,N_820,N_837);
xnor U1002 (N_1002,N_932,N_922);
nand U1003 (N_1003,N_842,N_869);
and U1004 (N_1004,N_892,N_945);
and U1005 (N_1005,N_817,N_961);
nor U1006 (N_1006,N_880,N_877);
nor U1007 (N_1007,N_935,N_901);
nand U1008 (N_1008,N_900,N_946);
nor U1009 (N_1009,N_910,N_891);
nand U1010 (N_1010,N_850,N_840);
nand U1011 (N_1011,N_934,N_841);
nor U1012 (N_1012,N_896,N_940);
and U1013 (N_1013,N_983,N_870);
nand U1014 (N_1014,N_960,N_907);
nor U1015 (N_1015,N_815,N_970);
and U1016 (N_1016,N_927,N_936);
xor U1017 (N_1017,N_996,N_810);
nor U1018 (N_1018,N_822,N_944);
and U1019 (N_1019,N_802,N_987);
nand U1020 (N_1020,N_807,N_884);
nand U1021 (N_1021,N_911,N_821);
xor U1022 (N_1022,N_941,N_957);
xor U1023 (N_1023,N_918,N_975);
and U1024 (N_1024,N_967,N_885);
xor U1025 (N_1025,N_883,N_836);
or U1026 (N_1026,N_929,N_858);
nand U1027 (N_1027,N_978,N_893);
nand U1028 (N_1028,N_931,N_980);
nand U1029 (N_1029,N_966,N_865);
and U1030 (N_1030,N_873,N_976);
nor U1031 (N_1031,N_906,N_832);
nand U1032 (N_1032,N_871,N_991);
xor U1033 (N_1033,N_845,N_888);
and U1034 (N_1034,N_834,N_851);
or U1035 (N_1035,N_823,N_833);
and U1036 (N_1036,N_952,N_926);
or U1037 (N_1037,N_992,N_997);
and U1038 (N_1038,N_812,N_999);
xor U1039 (N_1039,N_835,N_848);
and U1040 (N_1040,N_855,N_872);
xnor U1041 (N_1041,N_829,N_874);
xor U1042 (N_1042,N_894,N_838);
nor U1043 (N_1043,N_990,N_824);
or U1044 (N_1044,N_857,N_861);
xnor U1045 (N_1045,N_909,N_816);
nor U1046 (N_1046,N_953,N_844);
or U1047 (N_1047,N_956,N_813);
nand U1048 (N_1048,N_819,N_879);
or U1049 (N_1049,N_947,N_801);
nand U1050 (N_1050,N_854,N_915);
nor U1051 (N_1051,N_925,N_859);
and U1052 (N_1052,N_917,N_866);
xnor U1053 (N_1053,N_959,N_809);
xor U1054 (N_1054,N_862,N_951);
nor U1055 (N_1055,N_914,N_899);
or U1056 (N_1056,N_890,N_895);
and U1057 (N_1057,N_867,N_981);
xor U1058 (N_1058,N_818,N_928);
and U1059 (N_1059,N_864,N_803);
and U1060 (N_1060,N_964,N_973);
or U1061 (N_1061,N_852,N_839);
or U1062 (N_1062,N_958,N_924);
and U1063 (N_1063,N_827,N_887);
and U1064 (N_1064,N_942,N_828);
nor U1065 (N_1065,N_830,N_876);
nand U1066 (N_1066,N_889,N_912);
nand U1067 (N_1067,N_902,N_982);
nor U1068 (N_1068,N_979,N_863);
nor U1069 (N_1069,N_943,N_804);
nor U1070 (N_1070,N_984,N_995);
xor U1071 (N_1071,N_955,N_939);
nor U1072 (N_1072,N_938,N_849);
or U1073 (N_1073,N_806,N_994);
nand U1074 (N_1074,N_969,N_847);
and U1075 (N_1075,N_988,N_962);
nand U1076 (N_1076,N_856,N_963);
or U1077 (N_1077,N_933,N_954);
xor U1078 (N_1078,N_968,N_974);
xor U1079 (N_1079,N_868,N_881);
nor U1080 (N_1080,N_905,N_937);
and U1081 (N_1081,N_972,N_825);
nor U1082 (N_1082,N_805,N_977);
nor U1083 (N_1083,N_921,N_886);
and U1084 (N_1084,N_882,N_989);
nand U1085 (N_1085,N_846,N_965);
xor U1086 (N_1086,N_949,N_913);
xor U1087 (N_1087,N_908,N_860);
xnor U1088 (N_1088,N_811,N_993);
nor U1089 (N_1089,N_875,N_897);
xor U1090 (N_1090,N_923,N_919);
or U1091 (N_1091,N_903,N_904);
xor U1092 (N_1092,N_986,N_920);
xnor U1093 (N_1093,N_930,N_898);
or U1094 (N_1094,N_878,N_843);
or U1095 (N_1095,N_826,N_800);
xor U1096 (N_1096,N_948,N_950);
or U1097 (N_1097,N_916,N_998);
and U1098 (N_1098,N_971,N_853);
and U1099 (N_1099,N_831,N_985);
nand U1100 (N_1100,N_819,N_826);
nor U1101 (N_1101,N_964,N_950);
or U1102 (N_1102,N_960,N_930);
or U1103 (N_1103,N_957,N_884);
nand U1104 (N_1104,N_928,N_961);
or U1105 (N_1105,N_977,N_951);
and U1106 (N_1106,N_874,N_980);
xnor U1107 (N_1107,N_953,N_842);
nor U1108 (N_1108,N_838,N_892);
xnor U1109 (N_1109,N_978,N_940);
or U1110 (N_1110,N_869,N_952);
xor U1111 (N_1111,N_903,N_873);
nor U1112 (N_1112,N_840,N_929);
or U1113 (N_1113,N_829,N_824);
xnor U1114 (N_1114,N_836,N_974);
or U1115 (N_1115,N_887,N_904);
or U1116 (N_1116,N_867,N_835);
or U1117 (N_1117,N_992,N_958);
and U1118 (N_1118,N_929,N_935);
xor U1119 (N_1119,N_987,N_959);
and U1120 (N_1120,N_945,N_987);
nand U1121 (N_1121,N_964,N_810);
or U1122 (N_1122,N_999,N_940);
and U1123 (N_1123,N_846,N_950);
nor U1124 (N_1124,N_953,N_841);
nor U1125 (N_1125,N_949,N_918);
nand U1126 (N_1126,N_929,N_842);
nand U1127 (N_1127,N_983,N_881);
nor U1128 (N_1128,N_872,N_823);
and U1129 (N_1129,N_885,N_890);
nor U1130 (N_1130,N_998,N_927);
or U1131 (N_1131,N_943,N_934);
and U1132 (N_1132,N_828,N_971);
and U1133 (N_1133,N_852,N_978);
nand U1134 (N_1134,N_900,N_926);
nor U1135 (N_1135,N_862,N_864);
xnor U1136 (N_1136,N_858,N_891);
nand U1137 (N_1137,N_999,N_903);
or U1138 (N_1138,N_806,N_856);
and U1139 (N_1139,N_898,N_988);
or U1140 (N_1140,N_869,N_991);
and U1141 (N_1141,N_802,N_901);
nor U1142 (N_1142,N_927,N_957);
nand U1143 (N_1143,N_954,N_979);
or U1144 (N_1144,N_803,N_800);
and U1145 (N_1145,N_957,N_839);
xor U1146 (N_1146,N_960,N_840);
and U1147 (N_1147,N_966,N_826);
xor U1148 (N_1148,N_937,N_900);
or U1149 (N_1149,N_892,N_815);
nand U1150 (N_1150,N_960,N_863);
or U1151 (N_1151,N_997,N_853);
or U1152 (N_1152,N_861,N_932);
nor U1153 (N_1153,N_943,N_885);
nor U1154 (N_1154,N_864,N_998);
nand U1155 (N_1155,N_872,N_926);
xnor U1156 (N_1156,N_872,N_937);
xor U1157 (N_1157,N_889,N_869);
or U1158 (N_1158,N_974,N_927);
nand U1159 (N_1159,N_934,N_951);
nand U1160 (N_1160,N_899,N_894);
or U1161 (N_1161,N_881,N_971);
nor U1162 (N_1162,N_909,N_936);
nor U1163 (N_1163,N_887,N_805);
nand U1164 (N_1164,N_973,N_872);
and U1165 (N_1165,N_953,N_826);
and U1166 (N_1166,N_917,N_931);
and U1167 (N_1167,N_903,N_933);
nor U1168 (N_1168,N_871,N_892);
and U1169 (N_1169,N_896,N_869);
nor U1170 (N_1170,N_823,N_828);
nor U1171 (N_1171,N_894,N_983);
nor U1172 (N_1172,N_803,N_858);
nand U1173 (N_1173,N_854,N_929);
xor U1174 (N_1174,N_838,N_923);
xnor U1175 (N_1175,N_821,N_813);
xor U1176 (N_1176,N_979,N_826);
and U1177 (N_1177,N_962,N_976);
or U1178 (N_1178,N_961,N_859);
xnor U1179 (N_1179,N_946,N_953);
or U1180 (N_1180,N_843,N_894);
nor U1181 (N_1181,N_973,N_889);
nor U1182 (N_1182,N_836,N_948);
nand U1183 (N_1183,N_939,N_941);
or U1184 (N_1184,N_991,N_823);
nor U1185 (N_1185,N_842,N_877);
or U1186 (N_1186,N_991,N_909);
or U1187 (N_1187,N_817,N_939);
xnor U1188 (N_1188,N_945,N_890);
xnor U1189 (N_1189,N_934,N_889);
nor U1190 (N_1190,N_972,N_878);
nor U1191 (N_1191,N_919,N_951);
nor U1192 (N_1192,N_957,N_890);
nand U1193 (N_1193,N_971,N_926);
or U1194 (N_1194,N_867,N_998);
xnor U1195 (N_1195,N_855,N_951);
or U1196 (N_1196,N_826,N_915);
nand U1197 (N_1197,N_996,N_813);
and U1198 (N_1198,N_939,N_834);
or U1199 (N_1199,N_924,N_938);
and U1200 (N_1200,N_1002,N_1145);
and U1201 (N_1201,N_1042,N_1184);
xnor U1202 (N_1202,N_1045,N_1072);
and U1203 (N_1203,N_1140,N_1120);
xnor U1204 (N_1204,N_1025,N_1096);
nor U1205 (N_1205,N_1044,N_1074);
and U1206 (N_1206,N_1185,N_1060);
or U1207 (N_1207,N_1170,N_1158);
nor U1208 (N_1208,N_1136,N_1021);
nor U1209 (N_1209,N_1063,N_1017);
nor U1210 (N_1210,N_1113,N_1093);
nor U1211 (N_1211,N_1097,N_1103);
nand U1212 (N_1212,N_1116,N_1159);
or U1213 (N_1213,N_1182,N_1121);
or U1214 (N_1214,N_1026,N_1034);
and U1215 (N_1215,N_1156,N_1066);
nor U1216 (N_1216,N_1019,N_1050);
and U1217 (N_1217,N_1027,N_1062);
or U1218 (N_1218,N_1181,N_1127);
and U1219 (N_1219,N_1149,N_1101);
xor U1220 (N_1220,N_1051,N_1055);
nor U1221 (N_1221,N_1117,N_1197);
or U1222 (N_1222,N_1082,N_1146);
nand U1223 (N_1223,N_1118,N_1067);
or U1224 (N_1224,N_1162,N_1171);
or U1225 (N_1225,N_1141,N_1137);
xor U1226 (N_1226,N_1052,N_1176);
nand U1227 (N_1227,N_1195,N_1194);
and U1228 (N_1228,N_1020,N_1180);
nor U1229 (N_1229,N_1188,N_1179);
nor U1230 (N_1230,N_1196,N_1166);
or U1231 (N_1231,N_1148,N_1164);
or U1232 (N_1232,N_1088,N_1129);
nor U1233 (N_1233,N_1030,N_1153);
nor U1234 (N_1234,N_1155,N_1135);
and U1235 (N_1235,N_1183,N_1057);
or U1236 (N_1236,N_1080,N_1091);
or U1237 (N_1237,N_1092,N_1190);
nor U1238 (N_1238,N_1102,N_1187);
or U1239 (N_1239,N_1154,N_1069);
or U1240 (N_1240,N_1112,N_1032);
nor U1241 (N_1241,N_1005,N_1024);
or U1242 (N_1242,N_1107,N_1157);
nor U1243 (N_1243,N_1108,N_1014);
and U1244 (N_1244,N_1161,N_1192);
xor U1245 (N_1245,N_1064,N_1177);
xor U1246 (N_1246,N_1083,N_1077);
and U1247 (N_1247,N_1075,N_1009);
nand U1248 (N_1248,N_1001,N_1084);
xnor U1249 (N_1249,N_1011,N_1022);
nand U1250 (N_1250,N_1076,N_1168);
nor U1251 (N_1251,N_1079,N_1047);
and U1252 (N_1252,N_1125,N_1008);
and U1253 (N_1253,N_1173,N_1100);
xnor U1254 (N_1254,N_1152,N_1099);
or U1255 (N_1255,N_1006,N_1175);
and U1256 (N_1256,N_1143,N_1128);
xnor U1257 (N_1257,N_1058,N_1018);
and U1258 (N_1258,N_1048,N_1172);
and U1259 (N_1259,N_1086,N_1081);
nor U1260 (N_1260,N_1169,N_1105);
and U1261 (N_1261,N_1111,N_1191);
nor U1262 (N_1262,N_1073,N_1189);
nand U1263 (N_1263,N_1036,N_1056);
nand U1264 (N_1264,N_1174,N_1033);
and U1265 (N_1265,N_1012,N_1028);
or U1266 (N_1266,N_1139,N_1038);
and U1267 (N_1267,N_1040,N_1198);
xor U1268 (N_1268,N_1115,N_1061);
nor U1269 (N_1269,N_1163,N_1110);
and U1270 (N_1270,N_1160,N_1165);
xor U1271 (N_1271,N_1031,N_1142);
nor U1272 (N_1272,N_1003,N_1059);
nor U1273 (N_1273,N_1151,N_1126);
or U1274 (N_1274,N_1114,N_1186);
nor U1275 (N_1275,N_1123,N_1106);
or U1276 (N_1276,N_1029,N_1013);
xnor U1277 (N_1277,N_1109,N_1007);
nor U1278 (N_1278,N_1131,N_1000);
or U1279 (N_1279,N_1094,N_1098);
nand U1280 (N_1280,N_1087,N_1133);
and U1281 (N_1281,N_1090,N_1134);
nand U1282 (N_1282,N_1095,N_1104);
nand U1283 (N_1283,N_1015,N_1041);
and U1284 (N_1284,N_1147,N_1071);
and U1285 (N_1285,N_1144,N_1124);
xnor U1286 (N_1286,N_1037,N_1130);
nand U1287 (N_1287,N_1065,N_1119);
or U1288 (N_1288,N_1178,N_1089);
nor U1289 (N_1289,N_1085,N_1167);
xor U1290 (N_1290,N_1132,N_1150);
nor U1291 (N_1291,N_1070,N_1043);
nand U1292 (N_1292,N_1068,N_1016);
nand U1293 (N_1293,N_1039,N_1199);
nand U1294 (N_1294,N_1010,N_1049);
xor U1295 (N_1295,N_1023,N_1035);
or U1296 (N_1296,N_1078,N_1122);
or U1297 (N_1297,N_1004,N_1054);
nor U1298 (N_1298,N_1193,N_1046);
xnor U1299 (N_1299,N_1138,N_1053);
xnor U1300 (N_1300,N_1048,N_1006);
nand U1301 (N_1301,N_1048,N_1003);
xor U1302 (N_1302,N_1177,N_1033);
nor U1303 (N_1303,N_1188,N_1120);
nor U1304 (N_1304,N_1086,N_1015);
nor U1305 (N_1305,N_1009,N_1155);
xor U1306 (N_1306,N_1024,N_1177);
or U1307 (N_1307,N_1033,N_1106);
or U1308 (N_1308,N_1082,N_1191);
or U1309 (N_1309,N_1075,N_1071);
or U1310 (N_1310,N_1135,N_1150);
nor U1311 (N_1311,N_1196,N_1155);
xor U1312 (N_1312,N_1138,N_1048);
nand U1313 (N_1313,N_1168,N_1112);
nand U1314 (N_1314,N_1141,N_1147);
nor U1315 (N_1315,N_1163,N_1044);
or U1316 (N_1316,N_1004,N_1161);
or U1317 (N_1317,N_1011,N_1021);
and U1318 (N_1318,N_1055,N_1139);
xnor U1319 (N_1319,N_1055,N_1166);
or U1320 (N_1320,N_1071,N_1049);
xor U1321 (N_1321,N_1184,N_1114);
nand U1322 (N_1322,N_1076,N_1192);
xor U1323 (N_1323,N_1111,N_1110);
or U1324 (N_1324,N_1137,N_1164);
and U1325 (N_1325,N_1141,N_1044);
nor U1326 (N_1326,N_1012,N_1107);
xor U1327 (N_1327,N_1049,N_1149);
nand U1328 (N_1328,N_1076,N_1198);
nand U1329 (N_1329,N_1099,N_1024);
xor U1330 (N_1330,N_1046,N_1119);
nand U1331 (N_1331,N_1010,N_1051);
xnor U1332 (N_1332,N_1053,N_1128);
nor U1333 (N_1333,N_1080,N_1074);
nor U1334 (N_1334,N_1088,N_1041);
xnor U1335 (N_1335,N_1146,N_1059);
nand U1336 (N_1336,N_1152,N_1104);
nand U1337 (N_1337,N_1155,N_1191);
nor U1338 (N_1338,N_1119,N_1146);
or U1339 (N_1339,N_1035,N_1055);
xor U1340 (N_1340,N_1093,N_1029);
xor U1341 (N_1341,N_1107,N_1005);
or U1342 (N_1342,N_1176,N_1097);
nor U1343 (N_1343,N_1126,N_1191);
nand U1344 (N_1344,N_1190,N_1057);
and U1345 (N_1345,N_1090,N_1084);
or U1346 (N_1346,N_1105,N_1194);
nor U1347 (N_1347,N_1042,N_1070);
xnor U1348 (N_1348,N_1167,N_1068);
xnor U1349 (N_1349,N_1055,N_1193);
or U1350 (N_1350,N_1075,N_1169);
xnor U1351 (N_1351,N_1006,N_1104);
xnor U1352 (N_1352,N_1097,N_1114);
xnor U1353 (N_1353,N_1199,N_1144);
nor U1354 (N_1354,N_1166,N_1056);
nor U1355 (N_1355,N_1034,N_1016);
or U1356 (N_1356,N_1104,N_1001);
nand U1357 (N_1357,N_1020,N_1135);
nand U1358 (N_1358,N_1143,N_1032);
and U1359 (N_1359,N_1089,N_1058);
nor U1360 (N_1360,N_1082,N_1076);
and U1361 (N_1361,N_1169,N_1046);
xor U1362 (N_1362,N_1073,N_1045);
or U1363 (N_1363,N_1083,N_1124);
nand U1364 (N_1364,N_1040,N_1159);
xor U1365 (N_1365,N_1087,N_1013);
and U1366 (N_1366,N_1088,N_1034);
or U1367 (N_1367,N_1075,N_1110);
nand U1368 (N_1368,N_1019,N_1053);
nand U1369 (N_1369,N_1118,N_1126);
xnor U1370 (N_1370,N_1084,N_1131);
nor U1371 (N_1371,N_1006,N_1090);
or U1372 (N_1372,N_1156,N_1061);
and U1373 (N_1373,N_1146,N_1083);
and U1374 (N_1374,N_1155,N_1000);
or U1375 (N_1375,N_1076,N_1171);
xor U1376 (N_1376,N_1154,N_1143);
and U1377 (N_1377,N_1177,N_1166);
or U1378 (N_1378,N_1158,N_1028);
xor U1379 (N_1379,N_1157,N_1187);
xnor U1380 (N_1380,N_1134,N_1006);
xnor U1381 (N_1381,N_1071,N_1081);
xnor U1382 (N_1382,N_1157,N_1170);
nor U1383 (N_1383,N_1096,N_1084);
nor U1384 (N_1384,N_1133,N_1050);
nor U1385 (N_1385,N_1132,N_1095);
xnor U1386 (N_1386,N_1001,N_1108);
xor U1387 (N_1387,N_1036,N_1183);
and U1388 (N_1388,N_1039,N_1151);
nor U1389 (N_1389,N_1021,N_1046);
and U1390 (N_1390,N_1059,N_1057);
and U1391 (N_1391,N_1074,N_1017);
or U1392 (N_1392,N_1119,N_1073);
xnor U1393 (N_1393,N_1094,N_1056);
and U1394 (N_1394,N_1110,N_1088);
nand U1395 (N_1395,N_1119,N_1177);
or U1396 (N_1396,N_1136,N_1186);
nor U1397 (N_1397,N_1049,N_1150);
nand U1398 (N_1398,N_1142,N_1182);
nor U1399 (N_1399,N_1123,N_1137);
xnor U1400 (N_1400,N_1278,N_1393);
nand U1401 (N_1401,N_1382,N_1265);
and U1402 (N_1402,N_1331,N_1343);
xnor U1403 (N_1403,N_1294,N_1310);
or U1404 (N_1404,N_1222,N_1376);
nor U1405 (N_1405,N_1326,N_1271);
nand U1406 (N_1406,N_1311,N_1314);
nor U1407 (N_1407,N_1321,N_1272);
xor U1408 (N_1408,N_1253,N_1322);
xnor U1409 (N_1409,N_1318,N_1361);
or U1410 (N_1410,N_1209,N_1229);
and U1411 (N_1411,N_1224,N_1342);
xor U1412 (N_1412,N_1360,N_1238);
nor U1413 (N_1413,N_1217,N_1218);
nand U1414 (N_1414,N_1341,N_1230);
nand U1415 (N_1415,N_1205,N_1358);
nand U1416 (N_1416,N_1355,N_1249);
xnor U1417 (N_1417,N_1384,N_1204);
xor U1418 (N_1418,N_1369,N_1232);
or U1419 (N_1419,N_1263,N_1200);
nor U1420 (N_1420,N_1383,N_1228);
nor U1421 (N_1421,N_1291,N_1211);
nor U1422 (N_1422,N_1388,N_1324);
or U1423 (N_1423,N_1337,N_1395);
nand U1424 (N_1424,N_1338,N_1208);
and U1425 (N_1425,N_1289,N_1368);
nor U1426 (N_1426,N_1389,N_1373);
xor U1427 (N_1427,N_1375,N_1240);
nor U1428 (N_1428,N_1365,N_1279);
nor U1429 (N_1429,N_1367,N_1267);
nor U1430 (N_1430,N_1379,N_1247);
nor U1431 (N_1431,N_1219,N_1359);
or U1432 (N_1432,N_1259,N_1241);
nor U1433 (N_1433,N_1213,N_1214);
and U1434 (N_1434,N_1244,N_1352);
nand U1435 (N_1435,N_1348,N_1206);
and U1436 (N_1436,N_1227,N_1254);
xnor U1437 (N_1437,N_1235,N_1297);
nand U1438 (N_1438,N_1397,N_1275);
xor U1439 (N_1439,N_1345,N_1286);
nand U1440 (N_1440,N_1323,N_1266);
nand U1441 (N_1441,N_1216,N_1307);
nor U1442 (N_1442,N_1242,N_1334);
or U1443 (N_1443,N_1335,N_1203);
xnor U1444 (N_1444,N_1258,N_1333);
xor U1445 (N_1445,N_1372,N_1317);
or U1446 (N_1446,N_1277,N_1304);
and U1447 (N_1447,N_1243,N_1387);
or U1448 (N_1448,N_1293,N_1329);
nand U1449 (N_1449,N_1396,N_1308);
or U1450 (N_1450,N_1221,N_1210);
nor U1451 (N_1451,N_1299,N_1276);
and U1452 (N_1452,N_1377,N_1262);
nand U1453 (N_1453,N_1261,N_1251);
and U1454 (N_1454,N_1285,N_1269);
or U1455 (N_1455,N_1225,N_1336);
xor U1456 (N_1456,N_1357,N_1234);
nand U1457 (N_1457,N_1270,N_1264);
nor U1458 (N_1458,N_1282,N_1394);
nor U1459 (N_1459,N_1256,N_1273);
and U1460 (N_1460,N_1370,N_1281);
nand U1461 (N_1461,N_1363,N_1246);
nand U1462 (N_1462,N_1245,N_1300);
nand U1463 (N_1463,N_1378,N_1305);
or U1464 (N_1464,N_1292,N_1351);
nor U1465 (N_1465,N_1380,N_1362);
nand U1466 (N_1466,N_1316,N_1215);
nand U1467 (N_1467,N_1353,N_1315);
and U1468 (N_1468,N_1231,N_1313);
nor U1469 (N_1469,N_1250,N_1381);
and U1470 (N_1470,N_1385,N_1309);
nor U1471 (N_1471,N_1386,N_1349);
nor U1472 (N_1472,N_1296,N_1356);
or U1473 (N_1473,N_1371,N_1354);
and U1474 (N_1474,N_1301,N_1298);
or U1475 (N_1475,N_1290,N_1302);
and U1476 (N_1476,N_1332,N_1330);
xnor U1477 (N_1477,N_1390,N_1220);
nor U1478 (N_1478,N_1306,N_1319);
nor U1479 (N_1479,N_1274,N_1257);
and U1480 (N_1480,N_1392,N_1248);
and U1481 (N_1481,N_1255,N_1347);
or U1482 (N_1482,N_1398,N_1295);
or U1483 (N_1483,N_1223,N_1327);
and U1484 (N_1484,N_1207,N_1325);
nor U1485 (N_1485,N_1350,N_1202);
or U1486 (N_1486,N_1239,N_1236);
xnor U1487 (N_1487,N_1252,N_1268);
or U1488 (N_1488,N_1212,N_1346);
xor U1489 (N_1489,N_1287,N_1328);
nor U1490 (N_1490,N_1340,N_1303);
or U1491 (N_1491,N_1320,N_1283);
nor U1492 (N_1492,N_1366,N_1233);
nor U1493 (N_1493,N_1226,N_1344);
nor U1494 (N_1494,N_1312,N_1339);
and U1495 (N_1495,N_1280,N_1364);
nor U1496 (N_1496,N_1284,N_1260);
nor U1497 (N_1497,N_1399,N_1288);
and U1498 (N_1498,N_1391,N_1201);
nor U1499 (N_1499,N_1237,N_1374);
xor U1500 (N_1500,N_1330,N_1348);
nand U1501 (N_1501,N_1315,N_1327);
xnor U1502 (N_1502,N_1386,N_1251);
nand U1503 (N_1503,N_1258,N_1276);
and U1504 (N_1504,N_1332,N_1241);
xor U1505 (N_1505,N_1276,N_1319);
and U1506 (N_1506,N_1349,N_1364);
or U1507 (N_1507,N_1252,N_1276);
or U1508 (N_1508,N_1301,N_1284);
and U1509 (N_1509,N_1277,N_1228);
or U1510 (N_1510,N_1246,N_1230);
and U1511 (N_1511,N_1264,N_1279);
and U1512 (N_1512,N_1265,N_1207);
xor U1513 (N_1513,N_1211,N_1313);
and U1514 (N_1514,N_1216,N_1201);
or U1515 (N_1515,N_1395,N_1270);
nor U1516 (N_1516,N_1251,N_1344);
or U1517 (N_1517,N_1332,N_1260);
or U1518 (N_1518,N_1272,N_1377);
and U1519 (N_1519,N_1299,N_1301);
xor U1520 (N_1520,N_1380,N_1332);
nand U1521 (N_1521,N_1240,N_1319);
or U1522 (N_1522,N_1280,N_1337);
or U1523 (N_1523,N_1392,N_1234);
nor U1524 (N_1524,N_1218,N_1293);
nand U1525 (N_1525,N_1363,N_1389);
or U1526 (N_1526,N_1366,N_1389);
and U1527 (N_1527,N_1280,N_1299);
or U1528 (N_1528,N_1384,N_1292);
nor U1529 (N_1529,N_1261,N_1348);
and U1530 (N_1530,N_1275,N_1281);
xnor U1531 (N_1531,N_1346,N_1313);
and U1532 (N_1532,N_1312,N_1257);
nor U1533 (N_1533,N_1290,N_1346);
xnor U1534 (N_1534,N_1351,N_1232);
xnor U1535 (N_1535,N_1368,N_1372);
xnor U1536 (N_1536,N_1207,N_1394);
xnor U1537 (N_1537,N_1202,N_1228);
nand U1538 (N_1538,N_1357,N_1219);
or U1539 (N_1539,N_1308,N_1255);
xnor U1540 (N_1540,N_1343,N_1314);
xor U1541 (N_1541,N_1368,N_1320);
or U1542 (N_1542,N_1268,N_1290);
and U1543 (N_1543,N_1322,N_1389);
nor U1544 (N_1544,N_1204,N_1284);
nand U1545 (N_1545,N_1210,N_1369);
or U1546 (N_1546,N_1306,N_1289);
nor U1547 (N_1547,N_1343,N_1370);
nand U1548 (N_1548,N_1365,N_1292);
xor U1549 (N_1549,N_1271,N_1381);
nand U1550 (N_1550,N_1257,N_1219);
xnor U1551 (N_1551,N_1219,N_1349);
nor U1552 (N_1552,N_1202,N_1229);
xnor U1553 (N_1553,N_1206,N_1282);
and U1554 (N_1554,N_1225,N_1239);
and U1555 (N_1555,N_1357,N_1284);
nand U1556 (N_1556,N_1332,N_1223);
or U1557 (N_1557,N_1203,N_1353);
xor U1558 (N_1558,N_1310,N_1212);
and U1559 (N_1559,N_1364,N_1353);
and U1560 (N_1560,N_1244,N_1229);
xor U1561 (N_1561,N_1330,N_1255);
xnor U1562 (N_1562,N_1215,N_1227);
or U1563 (N_1563,N_1262,N_1226);
nand U1564 (N_1564,N_1322,N_1321);
and U1565 (N_1565,N_1399,N_1368);
and U1566 (N_1566,N_1226,N_1307);
xnor U1567 (N_1567,N_1271,N_1293);
and U1568 (N_1568,N_1356,N_1243);
nand U1569 (N_1569,N_1355,N_1288);
nand U1570 (N_1570,N_1208,N_1390);
nand U1571 (N_1571,N_1313,N_1322);
nor U1572 (N_1572,N_1230,N_1285);
and U1573 (N_1573,N_1317,N_1380);
nand U1574 (N_1574,N_1276,N_1261);
or U1575 (N_1575,N_1238,N_1241);
nand U1576 (N_1576,N_1287,N_1365);
xor U1577 (N_1577,N_1273,N_1393);
nor U1578 (N_1578,N_1291,N_1379);
or U1579 (N_1579,N_1280,N_1277);
nand U1580 (N_1580,N_1266,N_1331);
and U1581 (N_1581,N_1293,N_1383);
xor U1582 (N_1582,N_1338,N_1318);
xnor U1583 (N_1583,N_1344,N_1319);
or U1584 (N_1584,N_1215,N_1209);
xor U1585 (N_1585,N_1285,N_1311);
nor U1586 (N_1586,N_1326,N_1313);
and U1587 (N_1587,N_1272,N_1218);
and U1588 (N_1588,N_1268,N_1312);
or U1589 (N_1589,N_1357,N_1342);
or U1590 (N_1590,N_1259,N_1220);
or U1591 (N_1591,N_1288,N_1341);
and U1592 (N_1592,N_1361,N_1337);
xor U1593 (N_1593,N_1282,N_1334);
nor U1594 (N_1594,N_1317,N_1373);
nand U1595 (N_1595,N_1345,N_1332);
or U1596 (N_1596,N_1308,N_1270);
and U1597 (N_1597,N_1265,N_1395);
nand U1598 (N_1598,N_1379,N_1270);
and U1599 (N_1599,N_1216,N_1392);
nand U1600 (N_1600,N_1595,N_1424);
nor U1601 (N_1601,N_1587,N_1526);
nand U1602 (N_1602,N_1479,N_1461);
nor U1603 (N_1603,N_1540,N_1534);
nand U1604 (N_1604,N_1482,N_1580);
xor U1605 (N_1605,N_1583,N_1435);
xnor U1606 (N_1606,N_1505,N_1554);
and U1607 (N_1607,N_1557,N_1467);
and U1608 (N_1608,N_1458,N_1579);
or U1609 (N_1609,N_1430,N_1547);
and U1610 (N_1610,N_1406,N_1511);
and U1611 (N_1611,N_1468,N_1420);
nor U1612 (N_1612,N_1528,N_1447);
xor U1613 (N_1613,N_1499,N_1509);
nor U1614 (N_1614,N_1582,N_1408);
nand U1615 (N_1615,N_1454,N_1456);
or U1616 (N_1616,N_1485,N_1490);
xor U1617 (N_1617,N_1560,N_1586);
nand U1618 (N_1618,N_1597,N_1568);
nor U1619 (N_1619,N_1500,N_1551);
xor U1620 (N_1620,N_1413,N_1448);
nor U1621 (N_1621,N_1496,N_1571);
and U1622 (N_1622,N_1416,N_1489);
xnor U1623 (N_1623,N_1581,N_1402);
or U1624 (N_1624,N_1460,N_1512);
and U1625 (N_1625,N_1589,N_1535);
nor U1626 (N_1626,N_1522,N_1415);
nor U1627 (N_1627,N_1463,N_1441);
or U1628 (N_1628,N_1515,N_1513);
nand U1629 (N_1629,N_1539,N_1529);
xor U1630 (N_1630,N_1429,N_1561);
nand U1631 (N_1631,N_1562,N_1527);
and U1632 (N_1632,N_1543,N_1478);
and U1633 (N_1633,N_1472,N_1466);
or U1634 (N_1634,N_1436,N_1572);
nor U1635 (N_1635,N_1531,N_1550);
xor U1636 (N_1636,N_1409,N_1578);
and U1637 (N_1637,N_1410,N_1504);
or U1638 (N_1638,N_1514,N_1428);
nand U1639 (N_1639,N_1450,N_1525);
or U1640 (N_1640,N_1417,N_1446);
xnor U1641 (N_1641,N_1414,N_1412);
xnor U1642 (N_1642,N_1594,N_1474);
nand U1643 (N_1643,N_1486,N_1403);
nor U1644 (N_1644,N_1510,N_1439);
nor U1645 (N_1645,N_1459,N_1464);
nand U1646 (N_1646,N_1565,N_1518);
nor U1647 (N_1647,N_1549,N_1457);
nor U1648 (N_1648,N_1419,N_1411);
nor U1649 (N_1649,N_1563,N_1431);
nand U1650 (N_1650,N_1552,N_1443);
nand U1651 (N_1651,N_1471,N_1537);
nand U1652 (N_1652,N_1544,N_1596);
or U1653 (N_1653,N_1584,N_1524);
xnor U1654 (N_1654,N_1497,N_1542);
nand U1655 (N_1655,N_1426,N_1545);
or U1656 (N_1656,N_1400,N_1455);
or U1657 (N_1657,N_1442,N_1407);
xnor U1658 (N_1658,N_1538,N_1506);
nand U1659 (N_1659,N_1599,N_1590);
nand U1660 (N_1660,N_1492,N_1591);
nand U1661 (N_1661,N_1502,N_1520);
and U1662 (N_1662,N_1495,N_1517);
or U1663 (N_1663,N_1555,N_1541);
and U1664 (N_1664,N_1546,N_1427);
nand U1665 (N_1665,N_1519,N_1445);
nor U1666 (N_1666,N_1452,N_1477);
xor U1667 (N_1667,N_1548,N_1574);
nand U1668 (N_1668,N_1449,N_1508);
and U1669 (N_1669,N_1444,N_1438);
and U1670 (N_1670,N_1483,N_1418);
xnor U1671 (N_1671,N_1573,N_1501);
nand U1672 (N_1672,N_1576,N_1465);
nor U1673 (N_1673,N_1598,N_1521);
and U1674 (N_1674,N_1473,N_1421);
xnor U1675 (N_1675,N_1476,N_1536);
nor U1676 (N_1676,N_1491,N_1556);
or U1677 (N_1677,N_1437,N_1494);
nor U1678 (N_1678,N_1567,N_1493);
or U1679 (N_1679,N_1425,N_1592);
nand U1680 (N_1680,N_1401,N_1575);
and U1681 (N_1681,N_1453,N_1588);
and U1682 (N_1682,N_1593,N_1475);
and U1683 (N_1683,N_1480,N_1558);
nand U1684 (N_1684,N_1533,N_1530);
nor U1685 (N_1685,N_1488,N_1553);
xnor U1686 (N_1686,N_1559,N_1566);
nor U1687 (N_1687,N_1422,N_1434);
and U1688 (N_1688,N_1470,N_1423);
and U1689 (N_1689,N_1469,N_1564);
xor U1690 (N_1690,N_1577,N_1585);
nor U1691 (N_1691,N_1532,N_1498);
nor U1692 (N_1692,N_1481,N_1484);
and U1693 (N_1693,N_1432,N_1487);
or U1694 (N_1694,N_1451,N_1507);
and U1695 (N_1695,N_1405,N_1523);
or U1696 (N_1696,N_1440,N_1404);
nor U1697 (N_1697,N_1462,N_1569);
nand U1698 (N_1698,N_1570,N_1516);
and U1699 (N_1699,N_1433,N_1503);
nor U1700 (N_1700,N_1422,N_1462);
nor U1701 (N_1701,N_1458,N_1567);
or U1702 (N_1702,N_1535,N_1506);
nor U1703 (N_1703,N_1484,N_1523);
nor U1704 (N_1704,N_1493,N_1599);
and U1705 (N_1705,N_1516,N_1598);
xor U1706 (N_1706,N_1438,N_1574);
nor U1707 (N_1707,N_1486,N_1574);
nor U1708 (N_1708,N_1502,N_1554);
nand U1709 (N_1709,N_1472,N_1507);
nand U1710 (N_1710,N_1552,N_1479);
nand U1711 (N_1711,N_1447,N_1502);
nand U1712 (N_1712,N_1541,N_1571);
xnor U1713 (N_1713,N_1434,N_1466);
and U1714 (N_1714,N_1558,N_1574);
nor U1715 (N_1715,N_1543,N_1528);
or U1716 (N_1716,N_1467,N_1512);
xnor U1717 (N_1717,N_1408,N_1576);
xor U1718 (N_1718,N_1402,N_1458);
nand U1719 (N_1719,N_1539,N_1521);
and U1720 (N_1720,N_1539,N_1575);
nor U1721 (N_1721,N_1413,N_1472);
nor U1722 (N_1722,N_1573,N_1553);
or U1723 (N_1723,N_1471,N_1508);
or U1724 (N_1724,N_1469,N_1421);
nand U1725 (N_1725,N_1527,N_1530);
nor U1726 (N_1726,N_1541,N_1509);
or U1727 (N_1727,N_1444,N_1414);
nor U1728 (N_1728,N_1515,N_1449);
or U1729 (N_1729,N_1595,N_1534);
and U1730 (N_1730,N_1514,N_1453);
nand U1731 (N_1731,N_1556,N_1590);
xor U1732 (N_1732,N_1413,N_1500);
nand U1733 (N_1733,N_1463,N_1525);
nand U1734 (N_1734,N_1509,N_1403);
and U1735 (N_1735,N_1491,N_1476);
xor U1736 (N_1736,N_1440,N_1473);
and U1737 (N_1737,N_1513,N_1541);
or U1738 (N_1738,N_1530,N_1499);
nor U1739 (N_1739,N_1453,N_1445);
or U1740 (N_1740,N_1441,N_1561);
or U1741 (N_1741,N_1420,N_1517);
nand U1742 (N_1742,N_1491,N_1449);
nand U1743 (N_1743,N_1438,N_1562);
nand U1744 (N_1744,N_1591,N_1527);
nor U1745 (N_1745,N_1526,N_1409);
xnor U1746 (N_1746,N_1518,N_1400);
and U1747 (N_1747,N_1551,N_1502);
or U1748 (N_1748,N_1503,N_1567);
xor U1749 (N_1749,N_1494,N_1483);
or U1750 (N_1750,N_1583,N_1516);
nand U1751 (N_1751,N_1447,N_1486);
nor U1752 (N_1752,N_1460,N_1472);
nand U1753 (N_1753,N_1484,N_1478);
and U1754 (N_1754,N_1464,N_1452);
nand U1755 (N_1755,N_1595,N_1495);
nor U1756 (N_1756,N_1489,N_1415);
nor U1757 (N_1757,N_1491,N_1575);
xnor U1758 (N_1758,N_1461,N_1523);
nor U1759 (N_1759,N_1457,N_1472);
or U1760 (N_1760,N_1548,N_1417);
nand U1761 (N_1761,N_1432,N_1430);
or U1762 (N_1762,N_1589,N_1576);
or U1763 (N_1763,N_1592,N_1469);
and U1764 (N_1764,N_1516,N_1544);
or U1765 (N_1765,N_1456,N_1512);
nor U1766 (N_1766,N_1493,N_1558);
nor U1767 (N_1767,N_1457,N_1511);
and U1768 (N_1768,N_1442,N_1504);
nand U1769 (N_1769,N_1440,N_1408);
nand U1770 (N_1770,N_1508,N_1522);
xor U1771 (N_1771,N_1472,N_1448);
or U1772 (N_1772,N_1497,N_1500);
or U1773 (N_1773,N_1517,N_1431);
nand U1774 (N_1774,N_1518,N_1461);
xnor U1775 (N_1775,N_1472,N_1578);
and U1776 (N_1776,N_1531,N_1435);
nor U1777 (N_1777,N_1480,N_1485);
or U1778 (N_1778,N_1523,N_1541);
nor U1779 (N_1779,N_1402,N_1591);
or U1780 (N_1780,N_1533,N_1550);
xnor U1781 (N_1781,N_1470,N_1543);
and U1782 (N_1782,N_1498,N_1576);
and U1783 (N_1783,N_1466,N_1462);
and U1784 (N_1784,N_1542,N_1447);
and U1785 (N_1785,N_1422,N_1469);
nand U1786 (N_1786,N_1592,N_1450);
xor U1787 (N_1787,N_1497,N_1593);
nor U1788 (N_1788,N_1487,N_1421);
nand U1789 (N_1789,N_1505,N_1518);
and U1790 (N_1790,N_1559,N_1447);
and U1791 (N_1791,N_1524,N_1522);
nand U1792 (N_1792,N_1442,N_1413);
nand U1793 (N_1793,N_1538,N_1556);
nor U1794 (N_1794,N_1584,N_1428);
or U1795 (N_1795,N_1564,N_1597);
or U1796 (N_1796,N_1433,N_1580);
nor U1797 (N_1797,N_1489,N_1573);
and U1798 (N_1798,N_1469,N_1580);
or U1799 (N_1799,N_1430,N_1551);
or U1800 (N_1800,N_1705,N_1645);
or U1801 (N_1801,N_1701,N_1695);
nand U1802 (N_1802,N_1756,N_1779);
and U1803 (N_1803,N_1769,N_1679);
nand U1804 (N_1804,N_1642,N_1650);
or U1805 (N_1805,N_1714,N_1665);
nand U1806 (N_1806,N_1629,N_1640);
nand U1807 (N_1807,N_1758,N_1621);
nand U1808 (N_1808,N_1785,N_1661);
nand U1809 (N_1809,N_1658,N_1773);
nand U1810 (N_1810,N_1619,N_1707);
nor U1811 (N_1811,N_1611,N_1664);
nor U1812 (N_1812,N_1638,N_1681);
nand U1813 (N_1813,N_1699,N_1790);
nand U1814 (N_1814,N_1670,N_1602);
nor U1815 (N_1815,N_1666,N_1639);
nor U1816 (N_1816,N_1722,N_1624);
nor U1817 (N_1817,N_1609,N_1771);
and U1818 (N_1818,N_1637,N_1726);
and U1819 (N_1819,N_1703,N_1742);
xnor U1820 (N_1820,N_1649,N_1603);
nand U1821 (N_1821,N_1733,N_1716);
xnor U1822 (N_1822,N_1646,N_1713);
xor U1823 (N_1823,N_1618,N_1607);
nand U1824 (N_1824,N_1720,N_1676);
nand U1825 (N_1825,N_1648,N_1775);
nor U1826 (N_1826,N_1614,N_1751);
or U1827 (N_1827,N_1605,N_1796);
nand U1828 (N_1828,N_1715,N_1780);
or U1829 (N_1829,N_1612,N_1793);
nor U1830 (N_1830,N_1651,N_1753);
nand U1831 (N_1831,N_1749,N_1630);
or U1832 (N_1832,N_1702,N_1772);
nand U1833 (N_1833,N_1615,N_1739);
xnor U1834 (N_1834,N_1724,N_1655);
or U1835 (N_1835,N_1710,N_1709);
xor U1836 (N_1836,N_1697,N_1752);
and U1837 (N_1837,N_1704,N_1678);
and U1838 (N_1838,N_1660,N_1795);
and U1839 (N_1839,N_1672,N_1652);
and U1840 (N_1840,N_1731,N_1770);
nand U1841 (N_1841,N_1798,N_1634);
nor U1842 (N_1842,N_1685,N_1736);
and U1843 (N_1843,N_1784,N_1643);
xor U1844 (N_1844,N_1625,N_1719);
nor U1845 (N_1845,N_1765,N_1654);
or U1846 (N_1846,N_1711,N_1776);
or U1847 (N_1847,N_1606,N_1647);
xnor U1848 (N_1848,N_1735,N_1799);
nor U1849 (N_1849,N_1653,N_1669);
nor U1850 (N_1850,N_1667,N_1778);
and U1851 (N_1851,N_1692,N_1789);
nand U1852 (N_1852,N_1797,N_1766);
or U1853 (N_1853,N_1673,N_1777);
or U1854 (N_1854,N_1675,N_1718);
xnor U1855 (N_1855,N_1706,N_1748);
nor U1856 (N_1856,N_1750,N_1620);
xnor U1857 (N_1857,N_1662,N_1738);
or U1858 (N_1858,N_1723,N_1604);
and U1859 (N_1859,N_1668,N_1745);
or U1860 (N_1860,N_1633,N_1686);
nor U1861 (N_1861,N_1644,N_1659);
nand U1862 (N_1862,N_1761,N_1786);
and U1863 (N_1863,N_1622,N_1782);
xnor U1864 (N_1864,N_1743,N_1762);
nand U1865 (N_1865,N_1628,N_1641);
nand U1866 (N_1866,N_1768,N_1759);
xnor U1867 (N_1867,N_1656,N_1721);
xor U1868 (N_1868,N_1601,N_1684);
or U1869 (N_1869,N_1690,N_1610);
xnor U1870 (N_1870,N_1687,N_1682);
nand U1871 (N_1871,N_1698,N_1737);
and U1872 (N_1872,N_1663,N_1694);
or U1873 (N_1873,N_1754,N_1732);
nand U1874 (N_1874,N_1788,N_1740);
nor U1875 (N_1875,N_1693,N_1632);
and U1876 (N_1876,N_1741,N_1717);
xnor U1877 (N_1877,N_1623,N_1671);
nor U1878 (N_1878,N_1763,N_1728);
nor U1879 (N_1879,N_1635,N_1688);
nand U1880 (N_1880,N_1730,N_1613);
nor U1881 (N_1881,N_1700,N_1791);
nor U1882 (N_1882,N_1627,N_1708);
nor U1883 (N_1883,N_1608,N_1680);
and U1884 (N_1884,N_1787,N_1760);
and U1885 (N_1885,N_1657,N_1696);
nor U1886 (N_1886,N_1781,N_1712);
nor U1887 (N_1887,N_1764,N_1729);
xor U1888 (N_1888,N_1792,N_1725);
nand U1889 (N_1889,N_1674,N_1747);
nand U1890 (N_1890,N_1755,N_1689);
nor U1891 (N_1891,N_1757,N_1774);
or U1892 (N_1892,N_1636,N_1626);
nor U1893 (N_1893,N_1767,N_1783);
and U1894 (N_1894,N_1677,N_1691);
xor U1895 (N_1895,N_1727,N_1746);
nand U1896 (N_1896,N_1744,N_1734);
nand U1897 (N_1897,N_1600,N_1617);
nor U1898 (N_1898,N_1794,N_1631);
or U1899 (N_1899,N_1683,N_1616);
xor U1900 (N_1900,N_1607,N_1649);
nor U1901 (N_1901,N_1783,N_1606);
xnor U1902 (N_1902,N_1630,N_1655);
nor U1903 (N_1903,N_1668,N_1742);
or U1904 (N_1904,N_1674,N_1646);
nor U1905 (N_1905,N_1628,N_1634);
xor U1906 (N_1906,N_1600,N_1766);
nor U1907 (N_1907,N_1698,N_1632);
xnor U1908 (N_1908,N_1689,N_1774);
xnor U1909 (N_1909,N_1670,N_1736);
and U1910 (N_1910,N_1724,N_1770);
and U1911 (N_1911,N_1628,N_1614);
xnor U1912 (N_1912,N_1624,N_1605);
or U1913 (N_1913,N_1696,N_1792);
xnor U1914 (N_1914,N_1750,N_1738);
and U1915 (N_1915,N_1630,N_1616);
xor U1916 (N_1916,N_1783,N_1748);
or U1917 (N_1917,N_1786,N_1748);
and U1918 (N_1918,N_1722,N_1631);
xnor U1919 (N_1919,N_1601,N_1774);
nand U1920 (N_1920,N_1787,N_1752);
or U1921 (N_1921,N_1654,N_1696);
or U1922 (N_1922,N_1795,N_1642);
and U1923 (N_1923,N_1794,N_1740);
xnor U1924 (N_1924,N_1781,N_1603);
nor U1925 (N_1925,N_1664,N_1726);
xnor U1926 (N_1926,N_1665,N_1777);
or U1927 (N_1927,N_1775,N_1633);
or U1928 (N_1928,N_1753,N_1623);
nand U1929 (N_1929,N_1717,N_1720);
or U1930 (N_1930,N_1762,N_1619);
or U1931 (N_1931,N_1719,N_1674);
and U1932 (N_1932,N_1602,N_1611);
and U1933 (N_1933,N_1690,N_1672);
nor U1934 (N_1934,N_1773,N_1714);
nor U1935 (N_1935,N_1774,N_1703);
nand U1936 (N_1936,N_1740,N_1779);
nand U1937 (N_1937,N_1639,N_1762);
or U1938 (N_1938,N_1612,N_1637);
nand U1939 (N_1939,N_1695,N_1633);
and U1940 (N_1940,N_1601,N_1663);
xnor U1941 (N_1941,N_1759,N_1651);
or U1942 (N_1942,N_1662,N_1620);
nand U1943 (N_1943,N_1785,N_1747);
nand U1944 (N_1944,N_1600,N_1727);
or U1945 (N_1945,N_1747,N_1791);
nand U1946 (N_1946,N_1737,N_1763);
nand U1947 (N_1947,N_1659,N_1779);
and U1948 (N_1948,N_1609,N_1776);
nor U1949 (N_1949,N_1605,N_1633);
nand U1950 (N_1950,N_1716,N_1772);
xnor U1951 (N_1951,N_1635,N_1751);
nor U1952 (N_1952,N_1616,N_1633);
or U1953 (N_1953,N_1704,N_1782);
and U1954 (N_1954,N_1680,N_1690);
xor U1955 (N_1955,N_1697,N_1751);
nor U1956 (N_1956,N_1706,N_1752);
xor U1957 (N_1957,N_1698,N_1734);
nor U1958 (N_1958,N_1757,N_1713);
nand U1959 (N_1959,N_1676,N_1640);
xor U1960 (N_1960,N_1754,N_1673);
nand U1961 (N_1961,N_1711,N_1661);
xnor U1962 (N_1962,N_1755,N_1786);
nand U1963 (N_1963,N_1727,N_1629);
nand U1964 (N_1964,N_1665,N_1763);
nand U1965 (N_1965,N_1779,N_1603);
or U1966 (N_1966,N_1771,N_1684);
xor U1967 (N_1967,N_1647,N_1616);
xor U1968 (N_1968,N_1741,N_1757);
xor U1969 (N_1969,N_1639,N_1721);
xnor U1970 (N_1970,N_1679,N_1785);
nand U1971 (N_1971,N_1618,N_1694);
or U1972 (N_1972,N_1689,N_1624);
or U1973 (N_1973,N_1659,N_1671);
or U1974 (N_1974,N_1744,N_1660);
nor U1975 (N_1975,N_1762,N_1651);
nor U1976 (N_1976,N_1796,N_1616);
xnor U1977 (N_1977,N_1746,N_1658);
xnor U1978 (N_1978,N_1763,N_1739);
xor U1979 (N_1979,N_1638,N_1730);
xnor U1980 (N_1980,N_1762,N_1687);
nor U1981 (N_1981,N_1756,N_1635);
nor U1982 (N_1982,N_1639,N_1799);
and U1983 (N_1983,N_1671,N_1626);
and U1984 (N_1984,N_1728,N_1654);
and U1985 (N_1985,N_1608,N_1692);
and U1986 (N_1986,N_1770,N_1766);
or U1987 (N_1987,N_1725,N_1756);
nand U1988 (N_1988,N_1736,N_1606);
or U1989 (N_1989,N_1684,N_1696);
nor U1990 (N_1990,N_1797,N_1753);
and U1991 (N_1991,N_1698,N_1718);
xor U1992 (N_1992,N_1668,N_1728);
nand U1993 (N_1993,N_1722,N_1755);
and U1994 (N_1994,N_1600,N_1774);
nand U1995 (N_1995,N_1717,N_1700);
xnor U1996 (N_1996,N_1671,N_1656);
or U1997 (N_1997,N_1658,N_1794);
nor U1998 (N_1998,N_1790,N_1773);
nand U1999 (N_1999,N_1637,N_1702);
nand U2000 (N_2000,N_1809,N_1834);
or U2001 (N_2001,N_1881,N_1845);
and U2002 (N_2002,N_1841,N_1914);
or U2003 (N_2003,N_1849,N_1944);
and U2004 (N_2004,N_1890,N_1983);
or U2005 (N_2005,N_1970,N_1802);
xnor U2006 (N_2006,N_1876,N_1989);
or U2007 (N_2007,N_1918,N_1901);
and U2008 (N_2008,N_1953,N_1853);
nand U2009 (N_2009,N_1871,N_1893);
xor U2010 (N_2010,N_1882,N_1930);
nand U2011 (N_2011,N_1857,N_1839);
nand U2012 (N_2012,N_1819,N_1803);
and U2013 (N_2013,N_1813,N_1860);
nor U2014 (N_2014,N_1820,N_1800);
or U2015 (N_2015,N_1848,N_1910);
xnor U2016 (N_2016,N_1931,N_1879);
nand U2017 (N_2017,N_1869,N_1958);
nor U2018 (N_2018,N_1816,N_1974);
xor U2019 (N_2019,N_1924,N_1948);
xor U2020 (N_2020,N_1863,N_1965);
nand U2021 (N_2021,N_1998,N_1859);
or U2022 (N_2022,N_1905,N_1818);
and U2023 (N_2023,N_1887,N_1843);
or U2024 (N_2024,N_1904,N_1821);
and U2025 (N_2025,N_1969,N_1908);
or U2026 (N_2026,N_1927,N_1851);
or U2027 (N_2027,N_1868,N_1870);
nand U2028 (N_2028,N_1804,N_1939);
xnor U2029 (N_2029,N_1858,N_1942);
nor U2030 (N_2030,N_1866,N_1872);
or U2031 (N_2031,N_1894,N_1976);
xor U2032 (N_2032,N_1856,N_1832);
nand U2033 (N_2033,N_1999,N_1846);
and U2034 (N_2034,N_1961,N_1949);
nor U2035 (N_2035,N_1897,N_1885);
and U2036 (N_2036,N_1956,N_1847);
nand U2037 (N_2037,N_1815,N_1950);
or U2038 (N_2038,N_1929,N_1874);
or U2039 (N_2039,N_1824,N_1891);
or U2040 (N_2040,N_1896,N_1954);
or U2041 (N_2041,N_1862,N_1920);
and U2042 (N_2042,N_1917,N_1811);
nor U2043 (N_2043,N_1827,N_1867);
nand U2044 (N_2044,N_1826,N_1850);
and U2045 (N_2045,N_1875,N_1873);
or U2046 (N_2046,N_1806,N_1919);
or U2047 (N_2047,N_1943,N_1838);
nand U2048 (N_2048,N_1938,N_1928);
nor U2049 (N_2049,N_1993,N_1936);
nor U2050 (N_2050,N_1971,N_1984);
nor U2051 (N_2051,N_1842,N_1966);
nor U2052 (N_2052,N_1895,N_1996);
and U2053 (N_2053,N_1883,N_1903);
and U2054 (N_2054,N_1980,N_1955);
nand U2055 (N_2055,N_1889,N_1988);
and U2056 (N_2056,N_1822,N_1810);
nor U2057 (N_2057,N_1967,N_1829);
xor U2058 (N_2058,N_1801,N_1833);
or U2059 (N_2059,N_1884,N_1814);
nor U2060 (N_2060,N_1912,N_1864);
nand U2061 (N_2061,N_1991,N_1861);
nor U2062 (N_2062,N_1877,N_1925);
nor U2063 (N_2063,N_1972,N_1831);
xor U2064 (N_2064,N_1907,N_1830);
nand U2065 (N_2065,N_1952,N_1975);
nand U2066 (N_2066,N_1977,N_1902);
nor U2067 (N_2067,N_1964,N_1807);
or U2068 (N_2068,N_1978,N_1933);
nand U2069 (N_2069,N_1911,N_1968);
nor U2070 (N_2070,N_1994,N_1940);
xor U2071 (N_2071,N_1906,N_1888);
xnor U2072 (N_2072,N_1837,N_1995);
xor U2073 (N_2073,N_1945,N_1812);
nor U2074 (N_2074,N_1825,N_1937);
xnor U2075 (N_2075,N_1979,N_1854);
nand U2076 (N_2076,N_1899,N_1886);
or U2077 (N_2077,N_1844,N_1878);
nor U2078 (N_2078,N_1823,N_1951);
nand U2079 (N_2079,N_1973,N_1923);
nor U2080 (N_2080,N_1898,N_1828);
or U2081 (N_2081,N_1990,N_1963);
nand U2082 (N_2082,N_1922,N_1981);
and U2083 (N_2083,N_1921,N_1855);
and U2084 (N_2084,N_1808,N_1836);
nor U2085 (N_2085,N_1915,N_1982);
xnor U2086 (N_2086,N_1926,N_1913);
or U2087 (N_2087,N_1932,N_1947);
nor U2088 (N_2088,N_1900,N_1805);
or U2089 (N_2089,N_1941,N_1865);
nor U2090 (N_2090,N_1985,N_1960);
xor U2091 (N_2091,N_1909,N_1946);
and U2092 (N_2092,N_1959,N_1992);
nor U2093 (N_2093,N_1934,N_1916);
nor U2094 (N_2094,N_1817,N_1935);
or U2095 (N_2095,N_1835,N_1852);
nor U2096 (N_2096,N_1986,N_1892);
xor U2097 (N_2097,N_1987,N_1962);
and U2098 (N_2098,N_1997,N_1880);
nand U2099 (N_2099,N_1957,N_1840);
or U2100 (N_2100,N_1916,N_1821);
nand U2101 (N_2101,N_1834,N_1876);
and U2102 (N_2102,N_1984,N_1954);
nand U2103 (N_2103,N_1901,N_1972);
and U2104 (N_2104,N_1971,N_1923);
nor U2105 (N_2105,N_1865,N_1805);
xnor U2106 (N_2106,N_1826,N_1835);
and U2107 (N_2107,N_1920,N_1896);
nor U2108 (N_2108,N_1932,N_1902);
xor U2109 (N_2109,N_1943,N_1812);
nor U2110 (N_2110,N_1905,N_1800);
nand U2111 (N_2111,N_1916,N_1946);
xor U2112 (N_2112,N_1828,N_1974);
and U2113 (N_2113,N_1863,N_1839);
nor U2114 (N_2114,N_1868,N_1897);
nand U2115 (N_2115,N_1974,N_1924);
or U2116 (N_2116,N_1950,N_1886);
nand U2117 (N_2117,N_1936,N_1987);
nor U2118 (N_2118,N_1978,N_1905);
nand U2119 (N_2119,N_1986,N_1969);
nor U2120 (N_2120,N_1860,N_1935);
nand U2121 (N_2121,N_1901,N_1844);
or U2122 (N_2122,N_1802,N_1990);
and U2123 (N_2123,N_1910,N_1900);
xor U2124 (N_2124,N_1802,N_1945);
and U2125 (N_2125,N_1934,N_1809);
nor U2126 (N_2126,N_1934,N_1914);
xor U2127 (N_2127,N_1948,N_1938);
nor U2128 (N_2128,N_1983,N_1966);
xor U2129 (N_2129,N_1836,N_1958);
xor U2130 (N_2130,N_1870,N_1832);
nor U2131 (N_2131,N_1891,N_1811);
or U2132 (N_2132,N_1932,N_1896);
or U2133 (N_2133,N_1903,N_1969);
xor U2134 (N_2134,N_1810,N_1974);
nand U2135 (N_2135,N_1807,N_1992);
xor U2136 (N_2136,N_1930,N_1956);
nor U2137 (N_2137,N_1941,N_1947);
or U2138 (N_2138,N_1874,N_1821);
nor U2139 (N_2139,N_1875,N_1814);
nor U2140 (N_2140,N_1913,N_1990);
or U2141 (N_2141,N_1941,N_1847);
and U2142 (N_2142,N_1869,N_1849);
and U2143 (N_2143,N_1937,N_1983);
and U2144 (N_2144,N_1921,N_1940);
nand U2145 (N_2145,N_1975,N_1883);
xor U2146 (N_2146,N_1837,N_1806);
nor U2147 (N_2147,N_1936,N_1932);
or U2148 (N_2148,N_1932,N_1980);
nand U2149 (N_2149,N_1820,N_1817);
nor U2150 (N_2150,N_1808,N_1879);
nor U2151 (N_2151,N_1831,N_1880);
nand U2152 (N_2152,N_1813,N_1856);
or U2153 (N_2153,N_1941,N_1851);
or U2154 (N_2154,N_1994,N_1811);
and U2155 (N_2155,N_1824,N_1857);
xnor U2156 (N_2156,N_1899,N_1904);
xnor U2157 (N_2157,N_1812,N_1909);
nand U2158 (N_2158,N_1890,N_1988);
nor U2159 (N_2159,N_1825,N_1944);
or U2160 (N_2160,N_1871,N_1941);
nor U2161 (N_2161,N_1883,N_1919);
and U2162 (N_2162,N_1941,N_1919);
nor U2163 (N_2163,N_1908,N_1946);
and U2164 (N_2164,N_1895,N_1970);
nor U2165 (N_2165,N_1940,N_1892);
or U2166 (N_2166,N_1932,N_1807);
xnor U2167 (N_2167,N_1826,N_1841);
nand U2168 (N_2168,N_1857,N_1883);
nor U2169 (N_2169,N_1957,N_1922);
or U2170 (N_2170,N_1864,N_1923);
and U2171 (N_2171,N_1829,N_1868);
or U2172 (N_2172,N_1855,N_1840);
xor U2173 (N_2173,N_1973,N_1876);
and U2174 (N_2174,N_1844,N_1906);
and U2175 (N_2175,N_1934,N_1879);
xor U2176 (N_2176,N_1894,N_1992);
and U2177 (N_2177,N_1986,N_1883);
or U2178 (N_2178,N_1812,N_1857);
and U2179 (N_2179,N_1974,N_1841);
nand U2180 (N_2180,N_1978,N_1812);
and U2181 (N_2181,N_1995,N_1875);
and U2182 (N_2182,N_1928,N_1816);
nor U2183 (N_2183,N_1896,N_1860);
xor U2184 (N_2184,N_1865,N_1924);
nand U2185 (N_2185,N_1897,N_1916);
and U2186 (N_2186,N_1845,N_1823);
or U2187 (N_2187,N_1984,N_1946);
or U2188 (N_2188,N_1954,N_1899);
or U2189 (N_2189,N_1892,N_1842);
nor U2190 (N_2190,N_1995,N_1935);
nand U2191 (N_2191,N_1955,N_1957);
and U2192 (N_2192,N_1986,N_1956);
nor U2193 (N_2193,N_1806,N_1853);
or U2194 (N_2194,N_1890,N_1828);
and U2195 (N_2195,N_1960,N_1984);
and U2196 (N_2196,N_1864,N_1859);
nand U2197 (N_2197,N_1974,N_1897);
nor U2198 (N_2198,N_1874,N_1915);
nand U2199 (N_2199,N_1911,N_1879);
nand U2200 (N_2200,N_2080,N_2024);
nor U2201 (N_2201,N_2131,N_2137);
nor U2202 (N_2202,N_2098,N_2108);
nor U2203 (N_2203,N_2013,N_2079);
nor U2204 (N_2204,N_2068,N_2180);
nand U2205 (N_2205,N_2146,N_2158);
xnor U2206 (N_2206,N_2077,N_2006);
and U2207 (N_2207,N_2078,N_2076);
nor U2208 (N_2208,N_2015,N_2115);
and U2209 (N_2209,N_2103,N_2133);
and U2210 (N_2210,N_2136,N_2122);
xnor U2211 (N_2211,N_2190,N_2134);
or U2212 (N_2212,N_2163,N_2193);
or U2213 (N_2213,N_2094,N_2199);
nor U2214 (N_2214,N_2139,N_2121);
xor U2215 (N_2215,N_2007,N_2135);
and U2216 (N_2216,N_2197,N_2039);
or U2217 (N_2217,N_2184,N_2155);
and U2218 (N_2218,N_2052,N_2099);
xor U2219 (N_2219,N_2125,N_2093);
or U2220 (N_2220,N_2128,N_2160);
or U2221 (N_2221,N_2109,N_2161);
or U2222 (N_2222,N_2042,N_2111);
nor U2223 (N_2223,N_2063,N_2124);
nand U2224 (N_2224,N_2171,N_2038);
xor U2225 (N_2225,N_2172,N_2016);
nand U2226 (N_2226,N_2054,N_2130);
nand U2227 (N_2227,N_2048,N_2084);
nand U2228 (N_2228,N_2011,N_2150);
or U2229 (N_2229,N_2018,N_2085);
or U2230 (N_2230,N_2174,N_2120);
nand U2231 (N_2231,N_2144,N_2075);
xor U2232 (N_2232,N_2065,N_2058);
nor U2233 (N_2233,N_2166,N_2088);
or U2234 (N_2234,N_2176,N_2072);
xor U2235 (N_2235,N_2126,N_2100);
xor U2236 (N_2236,N_2169,N_2031);
nor U2237 (N_2237,N_2053,N_2110);
or U2238 (N_2238,N_2044,N_2097);
and U2239 (N_2239,N_2112,N_2026);
or U2240 (N_2240,N_2086,N_2025);
and U2241 (N_2241,N_2071,N_2089);
xor U2242 (N_2242,N_2141,N_2057);
and U2243 (N_2243,N_2001,N_2104);
and U2244 (N_2244,N_2185,N_2145);
and U2245 (N_2245,N_2188,N_2073);
nand U2246 (N_2246,N_2191,N_2138);
nand U2247 (N_2247,N_2004,N_2041);
or U2248 (N_2248,N_2147,N_2061);
xnor U2249 (N_2249,N_2021,N_2168);
or U2250 (N_2250,N_2183,N_2027);
nand U2251 (N_2251,N_2127,N_2037);
nand U2252 (N_2252,N_2173,N_2119);
and U2253 (N_2253,N_2095,N_2033);
nand U2254 (N_2254,N_2043,N_2192);
nand U2255 (N_2255,N_2036,N_2177);
or U2256 (N_2256,N_2090,N_2123);
nand U2257 (N_2257,N_2074,N_2096);
or U2258 (N_2258,N_2187,N_2114);
nand U2259 (N_2259,N_2181,N_2142);
xnor U2260 (N_2260,N_2092,N_2029);
xor U2261 (N_2261,N_2189,N_2028);
and U2262 (N_2262,N_2148,N_2106);
xor U2263 (N_2263,N_2164,N_2129);
nor U2264 (N_2264,N_2165,N_2175);
nand U2265 (N_2265,N_2149,N_2059);
nand U2266 (N_2266,N_2022,N_2170);
and U2267 (N_2267,N_2102,N_2051);
or U2268 (N_2268,N_2113,N_2049);
nand U2269 (N_2269,N_2046,N_2194);
or U2270 (N_2270,N_2087,N_2000);
nand U2271 (N_2271,N_2014,N_2017);
xor U2272 (N_2272,N_2082,N_2010);
nor U2273 (N_2273,N_2101,N_2034);
xnor U2274 (N_2274,N_2159,N_2140);
or U2275 (N_2275,N_2045,N_2009);
nor U2276 (N_2276,N_2157,N_2091);
nor U2277 (N_2277,N_2047,N_2196);
or U2278 (N_2278,N_2156,N_2020);
nor U2279 (N_2279,N_2023,N_2083);
xnor U2280 (N_2280,N_2153,N_2005);
xor U2281 (N_2281,N_2060,N_2067);
xnor U2282 (N_2282,N_2002,N_2008);
nand U2283 (N_2283,N_2195,N_2132);
or U2284 (N_2284,N_2056,N_2062);
xor U2285 (N_2285,N_2066,N_2117);
nor U2286 (N_2286,N_2178,N_2167);
nor U2287 (N_2287,N_2032,N_2154);
nand U2288 (N_2288,N_2182,N_2019);
nand U2289 (N_2289,N_2003,N_2064);
xnor U2290 (N_2290,N_2105,N_2143);
and U2291 (N_2291,N_2070,N_2179);
nor U2292 (N_2292,N_2081,N_2012);
xor U2293 (N_2293,N_2055,N_2030);
xor U2294 (N_2294,N_2152,N_2186);
nor U2295 (N_2295,N_2162,N_2151);
nor U2296 (N_2296,N_2050,N_2107);
nand U2297 (N_2297,N_2118,N_2069);
and U2298 (N_2298,N_2035,N_2040);
or U2299 (N_2299,N_2116,N_2198);
and U2300 (N_2300,N_2166,N_2184);
and U2301 (N_2301,N_2105,N_2018);
and U2302 (N_2302,N_2054,N_2096);
or U2303 (N_2303,N_2012,N_2017);
xnor U2304 (N_2304,N_2053,N_2178);
nor U2305 (N_2305,N_2124,N_2176);
xnor U2306 (N_2306,N_2094,N_2191);
nand U2307 (N_2307,N_2083,N_2051);
or U2308 (N_2308,N_2028,N_2039);
nand U2309 (N_2309,N_2071,N_2115);
nor U2310 (N_2310,N_2170,N_2062);
and U2311 (N_2311,N_2069,N_2036);
nand U2312 (N_2312,N_2050,N_2095);
xor U2313 (N_2313,N_2187,N_2040);
nand U2314 (N_2314,N_2016,N_2176);
and U2315 (N_2315,N_2035,N_2120);
xnor U2316 (N_2316,N_2051,N_2141);
nand U2317 (N_2317,N_2126,N_2058);
nor U2318 (N_2318,N_2194,N_2022);
nand U2319 (N_2319,N_2047,N_2010);
or U2320 (N_2320,N_2163,N_2087);
or U2321 (N_2321,N_2032,N_2178);
nand U2322 (N_2322,N_2193,N_2003);
nor U2323 (N_2323,N_2151,N_2062);
xnor U2324 (N_2324,N_2177,N_2126);
nand U2325 (N_2325,N_2126,N_2154);
and U2326 (N_2326,N_2136,N_2073);
nand U2327 (N_2327,N_2184,N_2068);
nand U2328 (N_2328,N_2002,N_2125);
and U2329 (N_2329,N_2012,N_2085);
or U2330 (N_2330,N_2010,N_2022);
nor U2331 (N_2331,N_2076,N_2034);
and U2332 (N_2332,N_2116,N_2070);
xnor U2333 (N_2333,N_2131,N_2109);
nor U2334 (N_2334,N_2018,N_2054);
nand U2335 (N_2335,N_2177,N_2093);
nand U2336 (N_2336,N_2090,N_2051);
xnor U2337 (N_2337,N_2185,N_2077);
and U2338 (N_2338,N_2105,N_2180);
nand U2339 (N_2339,N_2193,N_2063);
nand U2340 (N_2340,N_2042,N_2188);
and U2341 (N_2341,N_2007,N_2138);
nor U2342 (N_2342,N_2087,N_2103);
or U2343 (N_2343,N_2116,N_2171);
nor U2344 (N_2344,N_2187,N_2029);
or U2345 (N_2345,N_2017,N_2049);
nand U2346 (N_2346,N_2171,N_2196);
nor U2347 (N_2347,N_2076,N_2090);
xor U2348 (N_2348,N_2072,N_2087);
xor U2349 (N_2349,N_2033,N_2189);
xor U2350 (N_2350,N_2195,N_2196);
nand U2351 (N_2351,N_2104,N_2164);
or U2352 (N_2352,N_2091,N_2183);
nand U2353 (N_2353,N_2196,N_2133);
or U2354 (N_2354,N_2125,N_2131);
nor U2355 (N_2355,N_2007,N_2069);
and U2356 (N_2356,N_2081,N_2138);
nor U2357 (N_2357,N_2068,N_2162);
nand U2358 (N_2358,N_2025,N_2045);
nand U2359 (N_2359,N_2009,N_2029);
xor U2360 (N_2360,N_2094,N_2088);
and U2361 (N_2361,N_2180,N_2109);
nand U2362 (N_2362,N_2009,N_2190);
nor U2363 (N_2363,N_2149,N_2150);
xnor U2364 (N_2364,N_2193,N_2100);
nor U2365 (N_2365,N_2163,N_2003);
nand U2366 (N_2366,N_2167,N_2090);
nand U2367 (N_2367,N_2102,N_2112);
or U2368 (N_2368,N_2081,N_2129);
nor U2369 (N_2369,N_2096,N_2122);
or U2370 (N_2370,N_2109,N_2018);
nor U2371 (N_2371,N_2157,N_2005);
or U2372 (N_2372,N_2056,N_2078);
and U2373 (N_2373,N_2100,N_2176);
and U2374 (N_2374,N_2133,N_2034);
nand U2375 (N_2375,N_2070,N_2098);
and U2376 (N_2376,N_2002,N_2100);
and U2377 (N_2377,N_2171,N_2076);
or U2378 (N_2378,N_2103,N_2040);
and U2379 (N_2379,N_2009,N_2140);
nor U2380 (N_2380,N_2069,N_2040);
nor U2381 (N_2381,N_2081,N_2114);
nor U2382 (N_2382,N_2119,N_2101);
and U2383 (N_2383,N_2003,N_2187);
nor U2384 (N_2384,N_2047,N_2186);
nand U2385 (N_2385,N_2020,N_2192);
or U2386 (N_2386,N_2068,N_2002);
and U2387 (N_2387,N_2154,N_2146);
nand U2388 (N_2388,N_2101,N_2170);
or U2389 (N_2389,N_2154,N_2088);
or U2390 (N_2390,N_2036,N_2099);
nand U2391 (N_2391,N_2046,N_2049);
and U2392 (N_2392,N_2195,N_2036);
xor U2393 (N_2393,N_2109,N_2148);
nor U2394 (N_2394,N_2137,N_2121);
xor U2395 (N_2395,N_2043,N_2194);
nand U2396 (N_2396,N_2120,N_2033);
xor U2397 (N_2397,N_2001,N_2184);
nor U2398 (N_2398,N_2013,N_2099);
nand U2399 (N_2399,N_2045,N_2161);
xor U2400 (N_2400,N_2331,N_2344);
nor U2401 (N_2401,N_2268,N_2320);
xor U2402 (N_2402,N_2307,N_2236);
nor U2403 (N_2403,N_2241,N_2222);
or U2404 (N_2404,N_2248,N_2308);
xor U2405 (N_2405,N_2330,N_2257);
or U2406 (N_2406,N_2359,N_2285);
xnor U2407 (N_2407,N_2319,N_2276);
xnor U2408 (N_2408,N_2382,N_2376);
or U2409 (N_2409,N_2314,N_2312);
nand U2410 (N_2410,N_2315,N_2295);
nor U2411 (N_2411,N_2203,N_2289);
nor U2412 (N_2412,N_2323,N_2290);
nand U2413 (N_2413,N_2372,N_2354);
nor U2414 (N_2414,N_2322,N_2357);
or U2415 (N_2415,N_2393,N_2262);
and U2416 (N_2416,N_2286,N_2238);
nand U2417 (N_2417,N_2346,N_2250);
and U2418 (N_2418,N_2387,N_2399);
nand U2419 (N_2419,N_2209,N_2227);
nor U2420 (N_2420,N_2326,N_2324);
or U2421 (N_2421,N_2310,N_2215);
nor U2422 (N_2422,N_2208,N_2242);
or U2423 (N_2423,N_2362,N_2366);
nand U2424 (N_2424,N_2282,N_2259);
nand U2425 (N_2425,N_2380,N_2240);
and U2426 (N_2426,N_2304,N_2321);
or U2427 (N_2427,N_2339,N_2228);
and U2428 (N_2428,N_2235,N_2297);
xnor U2429 (N_2429,N_2337,N_2234);
or U2430 (N_2430,N_2274,N_2288);
nand U2431 (N_2431,N_2340,N_2313);
or U2432 (N_2432,N_2309,N_2206);
nand U2433 (N_2433,N_2266,N_2394);
xnor U2434 (N_2434,N_2223,N_2389);
nand U2435 (N_2435,N_2244,N_2249);
nand U2436 (N_2436,N_2218,N_2378);
xnor U2437 (N_2437,N_2329,N_2260);
nor U2438 (N_2438,N_2349,N_2332);
xor U2439 (N_2439,N_2233,N_2284);
nor U2440 (N_2440,N_2371,N_2367);
or U2441 (N_2441,N_2316,N_2267);
nor U2442 (N_2442,N_2377,N_2336);
nand U2443 (N_2443,N_2296,N_2224);
nand U2444 (N_2444,N_2258,N_2201);
or U2445 (N_2445,N_2369,N_2395);
and U2446 (N_2446,N_2300,N_2255);
nand U2447 (N_2447,N_2353,N_2390);
or U2448 (N_2448,N_2303,N_2375);
or U2449 (N_2449,N_2271,N_2318);
nand U2450 (N_2450,N_2239,N_2202);
and U2451 (N_2451,N_2247,N_2213);
and U2452 (N_2452,N_2293,N_2343);
nand U2453 (N_2453,N_2216,N_2200);
and U2454 (N_2454,N_2335,N_2392);
xnor U2455 (N_2455,N_2269,N_2325);
nor U2456 (N_2456,N_2384,N_2230);
nand U2457 (N_2457,N_2370,N_2365);
or U2458 (N_2458,N_2270,N_2298);
xnor U2459 (N_2459,N_2381,N_2229);
nand U2460 (N_2460,N_2272,N_2342);
nor U2461 (N_2461,N_2283,N_2292);
nand U2462 (N_2462,N_2205,N_2275);
or U2463 (N_2463,N_2356,N_2306);
and U2464 (N_2464,N_2386,N_2221);
nor U2465 (N_2465,N_2214,N_2252);
xnor U2466 (N_2466,N_2251,N_2364);
nand U2467 (N_2467,N_2279,N_2226);
nor U2468 (N_2468,N_2207,N_2397);
and U2469 (N_2469,N_2338,N_2265);
xor U2470 (N_2470,N_2287,N_2305);
xnor U2471 (N_2471,N_2245,N_2273);
xnor U2472 (N_2472,N_2294,N_2263);
and U2473 (N_2473,N_2211,N_2280);
and U2474 (N_2474,N_2351,N_2256);
or U2475 (N_2475,N_2210,N_2352);
or U2476 (N_2476,N_2345,N_2361);
and U2477 (N_2477,N_2311,N_2281);
nand U2478 (N_2478,N_2301,N_2341);
nand U2479 (N_2479,N_2363,N_2374);
xnor U2480 (N_2480,N_2385,N_2254);
or U2481 (N_2481,N_2379,N_2264);
and U2482 (N_2482,N_2383,N_2398);
nor U2483 (N_2483,N_2348,N_2246);
and U2484 (N_2484,N_2277,N_2355);
nand U2485 (N_2485,N_2396,N_2278);
xnor U2486 (N_2486,N_2334,N_2333);
or U2487 (N_2487,N_2220,N_2391);
or U2488 (N_2488,N_2243,N_2373);
or U2489 (N_2489,N_2368,N_2231);
xor U2490 (N_2490,N_2317,N_2388);
xor U2491 (N_2491,N_2360,N_2253);
and U2492 (N_2492,N_2299,N_2232);
nand U2493 (N_2493,N_2350,N_2358);
xor U2494 (N_2494,N_2212,N_2327);
nor U2495 (N_2495,N_2261,N_2219);
nor U2496 (N_2496,N_2225,N_2204);
or U2497 (N_2497,N_2217,N_2291);
and U2498 (N_2498,N_2347,N_2302);
nand U2499 (N_2499,N_2328,N_2237);
nor U2500 (N_2500,N_2291,N_2327);
xor U2501 (N_2501,N_2390,N_2230);
nand U2502 (N_2502,N_2369,N_2363);
or U2503 (N_2503,N_2247,N_2288);
nor U2504 (N_2504,N_2255,N_2226);
nand U2505 (N_2505,N_2277,N_2339);
and U2506 (N_2506,N_2309,N_2379);
nor U2507 (N_2507,N_2257,N_2357);
nor U2508 (N_2508,N_2344,N_2286);
nand U2509 (N_2509,N_2292,N_2272);
and U2510 (N_2510,N_2201,N_2343);
and U2511 (N_2511,N_2258,N_2302);
nand U2512 (N_2512,N_2204,N_2223);
nor U2513 (N_2513,N_2313,N_2278);
nand U2514 (N_2514,N_2226,N_2336);
nand U2515 (N_2515,N_2337,N_2232);
xnor U2516 (N_2516,N_2314,N_2347);
nor U2517 (N_2517,N_2317,N_2289);
nand U2518 (N_2518,N_2264,N_2346);
and U2519 (N_2519,N_2375,N_2255);
nor U2520 (N_2520,N_2305,N_2247);
and U2521 (N_2521,N_2247,N_2328);
nor U2522 (N_2522,N_2269,N_2231);
or U2523 (N_2523,N_2251,N_2292);
or U2524 (N_2524,N_2349,N_2393);
or U2525 (N_2525,N_2363,N_2251);
or U2526 (N_2526,N_2327,N_2286);
nor U2527 (N_2527,N_2216,N_2236);
nand U2528 (N_2528,N_2234,N_2230);
and U2529 (N_2529,N_2315,N_2217);
nor U2530 (N_2530,N_2314,N_2244);
nor U2531 (N_2531,N_2300,N_2267);
or U2532 (N_2532,N_2250,N_2373);
nand U2533 (N_2533,N_2280,N_2345);
nand U2534 (N_2534,N_2334,N_2297);
xor U2535 (N_2535,N_2307,N_2262);
nor U2536 (N_2536,N_2269,N_2221);
nor U2537 (N_2537,N_2242,N_2327);
nand U2538 (N_2538,N_2333,N_2250);
xor U2539 (N_2539,N_2380,N_2271);
or U2540 (N_2540,N_2338,N_2253);
xor U2541 (N_2541,N_2246,N_2256);
or U2542 (N_2542,N_2325,N_2320);
and U2543 (N_2543,N_2395,N_2200);
xnor U2544 (N_2544,N_2270,N_2233);
or U2545 (N_2545,N_2227,N_2252);
and U2546 (N_2546,N_2355,N_2259);
nand U2547 (N_2547,N_2332,N_2253);
nand U2548 (N_2548,N_2314,N_2262);
xnor U2549 (N_2549,N_2315,N_2286);
nand U2550 (N_2550,N_2360,N_2340);
or U2551 (N_2551,N_2230,N_2241);
xnor U2552 (N_2552,N_2266,N_2338);
nand U2553 (N_2553,N_2362,N_2298);
nor U2554 (N_2554,N_2362,N_2247);
or U2555 (N_2555,N_2214,N_2211);
and U2556 (N_2556,N_2274,N_2258);
nor U2557 (N_2557,N_2344,N_2306);
nor U2558 (N_2558,N_2381,N_2297);
and U2559 (N_2559,N_2362,N_2233);
or U2560 (N_2560,N_2218,N_2303);
and U2561 (N_2561,N_2268,N_2271);
nand U2562 (N_2562,N_2322,N_2257);
nor U2563 (N_2563,N_2372,N_2389);
nor U2564 (N_2564,N_2376,N_2374);
nand U2565 (N_2565,N_2322,N_2260);
nor U2566 (N_2566,N_2237,N_2371);
or U2567 (N_2567,N_2336,N_2371);
nand U2568 (N_2568,N_2287,N_2240);
nor U2569 (N_2569,N_2209,N_2347);
xnor U2570 (N_2570,N_2331,N_2260);
xnor U2571 (N_2571,N_2346,N_2273);
or U2572 (N_2572,N_2233,N_2280);
nor U2573 (N_2573,N_2392,N_2233);
nor U2574 (N_2574,N_2396,N_2316);
and U2575 (N_2575,N_2205,N_2320);
xnor U2576 (N_2576,N_2235,N_2267);
nor U2577 (N_2577,N_2238,N_2200);
xor U2578 (N_2578,N_2207,N_2297);
and U2579 (N_2579,N_2360,N_2217);
nand U2580 (N_2580,N_2382,N_2337);
nand U2581 (N_2581,N_2222,N_2237);
and U2582 (N_2582,N_2323,N_2209);
and U2583 (N_2583,N_2293,N_2391);
and U2584 (N_2584,N_2293,N_2322);
xnor U2585 (N_2585,N_2329,N_2351);
and U2586 (N_2586,N_2254,N_2389);
nor U2587 (N_2587,N_2359,N_2236);
nand U2588 (N_2588,N_2338,N_2210);
or U2589 (N_2589,N_2314,N_2343);
nor U2590 (N_2590,N_2231,N_2356);
and U2591 (N_2591,N_2357,N_2261);
or U2592 (N_2592,N_2354,N_2336);
nand U2593 (N_2593,N_2265,N_2392);
nor U2594 (N_2594,N_2262,N_2322);
nand U2595 (N_2595,N_2378,N_2323);
and U2596 (N_2596,N_2379,N_2297);
nand U2597 (N_2597,N_2218,N_2288);
nand U2598 (N_2598,N_2399,N_2358);
and U2599 (N_2599,N_2239,N_2332);
and U2600 (N_2600,N_2596,N_2588);
nand U2601 (N_2601,N_2547,N_2589);
or U2602 (N_2602,N_2467,N_2514);
and U2603 (N_2603,N_2470,N_2541);
nor U2604 (N_2604,N_2409,N_2485);
and U2605 (N_2605,N_2402,N_2445);
and U2606 (N_2606,N_2460,N_2560);
nor U2607 (N_2607,N_2508,N_2568);
or U2608 (N_2608,N_2487,N_2517);
xnor U2609 (N_2609,N_2524,N_2439);
nand U2610 (N_2610,N_2537,N_2522);
xnor U2611 (N_2611,N_2571,N_2552);
or U2612 (N_2612,N_2546,N_2493);
nand U2613 (N_2613,N_2489,N_2488);
nand U2614 (N_2614,N_2490,N_2437);
nor U2615 (N_2615,N_2421,N_2406);
nor U2616 (N_2616,N_2598,N_2486);
xor U2617 (N_2617,N_2576,N_2431);
nor U2618 (N_2618,N_2449,N_2503);
and U2619 (N_2619,N_2566,N_2559);
or U2620 (N_2620,N_2574,N_2408);
or U2621 (N_2621,N_2511,N_2479);
xnor U2622 (N_2622,N_2443,N_2474);
or U2623 (N_2623,N_2450,N_2415);
nand U2624 (N_2624,N_2553,N_2498);
nand U2625 (N_2625,N_2533,N_2535);
and U2626 (N_2626,N_2412,N_2531);
xnor U2627 (N_2627,N_2575,N_2453);
nor U2628 (N_2628,N_2536,N_2454);
xor U2629 (N_2629,N_2513,N_2496);
xnor U2630 (N_2630,N_2400,N_2497);
or U2631 (N_2631,N_2519,N_2480);
or U2632 (N_2632,N_2591,N_2452);
or U2633 (N_2633,N_2581,N_2469);
nand U2634 (N_2634,N_2482,N_2595);
and U2635 (N_2635,N_2520,N_2464);
nor U2636 (N_2636,N_2407,N_2554);
nor U2637 (N_2637,N_2424,N_2426);
nor U2638 (N_2638,N_2599,N_2401);
or U2639 (N_2639,N_2572,N_2567);
xnor U2640 (N_2640,N_2446,N_2416);
nand U2641 (N_2641,N_2548,N_2465);
or U2642 (N_2642,N_2532,N_2459);
or U2643 (N_2643,N_2573,N_2504);
or U2644 (N_2644,N_2477,N_2577);
xor U2645 (N_2645,N_2475,N_2455);
xnor U2646 (N_2646,N_2563,N_2441);
nor U2647 (N_2647,N_2538,N_2448);
and U2648 (N_2648,N_2410,N_2413);
and U2649 (N_2649,N_2587,N_2580);
and U2650 (N_2650,N_2405,N_2420);
nor U2651 (N_2651,N_2428,N_2423);
xnor U2652 (N_2652,N_2510,N_2447);
or U2653 (N_2653,N_2462,N_2468);
xnor U2654 (N_2654,N_2505,N_2411);
nor U2655 (N_2655,N_2417,N_2433);
or U2656 (N_2656,N_2458,N_2509);
nor U2657 (N_2657,N_2463,N_2436);
nor U2658 (N_2658,N_2419,N_2570);
and U2659 (N_2659,N_2429,N_2515);
or U2660 (N_2660,N_2478,N_2471);
or U2661 (N_2661,N_2414,N_2530);
nand U2662 (N_2662,N_2523,N_2473);
nor U2663 (N_2663,N_2521,N_2582);
nor U2664 (N_2664,N_2444,N_2484);
xor U2665 (N_2665,N_2518,N_2438);
xor U2666 (N_2666,N_2425,N_2483);
nor U2667 (N_2667,N_2579,N_2555);
nor U2668 (N_2668,N_2481,N_2491);
nor U2669 (N_2669,N_2543,N_2435);
nand U2670 (N_2670,N_2528,N_2569);
or U2671 (N_2671,N_2525,N_2561);
nand U2672 (N_2672,N_2557,N_2526);
or U2673 (N_2673,N_2594,N_2451);
nor U2674 (N_2674,N_2418,N_2457);
or U2675 (N_2675,N_2590,N_2472);
or U2676 (N_2676,N_2494,N_2502);
nand U2677 (N_2677,N_2544,N_2404);
xor U2678 (N_2678,N_2597,N_2539);
nand U2679 (N_2679,N_2593,N_2461);
or U2680 (N_2680,N_2564,N_2527);
nor U2681 (N_2681,N_2427,N_2432);
or U2682 (N_2682,N_2456,N_2545);
xnor U2683 (N_2683,N_2540,N_2585);
or U2684 (N_2684,N_2550,N_2507);
xnor U2685 (N_2685,N_2549,N_2403);
or U2686 (N_2686,N_2434,N_2500);
nand U2687 (N_2687,N_2492,N_2440);
nor U2688 (N_2688,N_2495,N_2592);
nand U2689 (N_2689,N_2556,N_2558);
nor U2690 (N_2690,N_2501,N_2578);
xnor U2691 (N_2691,N_2534,N_2586);
nor U2692 (N_2692,N_2422,N_2430);
nor U2693 (N_2693,N_2442,N_2542);
and U2694 (N_2694,N_2583,N_2516);
nand U2695 (N_2695,N_2529,N_2476);
nor U2696 (N_2696,N_2466,N_2512);
nor U2697 (N_2697,N_2562,N_2565);
xnor U2698 (N_2698,N_2584,N_2499);
or U2699 (N_2699,N_2506,N_2551);
nor U2700 (N_2700,N_2413,N_2448);
and U2701 (N_2701,N_2476,N_2574);
and U2702 (N_2702,N_2467,N_2533);
or U2703 (N_2703,N_2548,N_2597);
nand U2704 (N_2704,N_2503,N_2406);
nand U2705 (N_2705,N_2579,N_2403);
and U2706 (N_2706,N_2534,N_2514);
xor U2707 (N_2707,N_2514,N_2578);
xnor U2708 (N_2708,N_2411,N_2497);
nor U2709 (N_2709,N_2460,N_2525);
xnor U2710 (N_2710,N_2405,N_2410);
xor U2711 (N_2711,N_2562,N_2493);
and U2712 (N_2712,N_2475,N_2576);
xor U2713 (N_2713,N_2577,N_2534);
or U2714 (N_2714,N_2458,N_2523);
nand U2715 (N_2715,N_2556,N_2497);
and U2716 (N_2716,N_2521,N_2416);
nand U2717 (N_2717,N_2442,N_2548);
xor U2718 (N_2718,N_2407,N_2506);
or U2719 (N_2719,N_2574,N_2471);
or U2720 (N_2720,N_2448,N_2444);
xor U2721 (N_2721,N_2405,N_2577);
nor U2722 (N_2722,N_2469,N_2572);
xnor U2723 (N_2723,N_2404,N_2474);
xnor U2724 (N_2724,N_2504,N_2531);
nand U2725 (N_2725,N_2461,N_2427);
and U2726 (N_2726,N_2571,N_2434);
xor U2727 (N_2727,N_2507,N_2471);
and U2728 (N_2728,N_2439,N_2536);
or U2729 (N_2729,N_2515,N_2446);
or U2730 (N_2730,N_2504,N_2412);
nand U2731 (N_2731,N_2518,N_2514);
or U2732 (N_2732,N_2544,N_2571);
nand U2733 (N_2733,N_2583,N_2500);
xnor U2734 (N_2734,N_2539,N_2406);
and U2735 (N_2735,N_2507,N_2454);
and U2736 (N_2736,N_2498,N_2597);
nor U2737 (N_2737,N_2520,N_2452);
nand U2738 (N_2738,N_2598,N_2470);
nor U2739 (N_2739,N_2452,N_2519);
nand U2740 (N_2740,N_2477,N_2540);
nor U2741 (N_2741,N_2513,N_2452);
nand U2742 (N_2742,N_2408,N_2465);
nand U2743 (N_2743,N_2546,N_2440);
and U2744 (N_2744,N_2456,N_2493);
or U2745 (N_2745,N_2452,N_2492);
or U2746 (N_2746,N_2584,N_2560);
or U2747 (N_2747,N_2447,N_2509);
nor U2748 (N_2748,N_2521,N_2586);
or U2749 (N_2749,N_2568,N_2448);
or U2750 (N_2750,N_2428,N_2417);
nor U2751 (N_2751,N_2528,N_2499);
nand U2752 (N_2752,N_2465,N_2490);
xor U2753 (N_2753,N_2479,N_2550);
or U2754 (N_2754,N_2560,N_2463);
nand U2755 (N_2755,N_2460,N_2567);
xnor U2756 (N_2756,N_2406,N_2548);
or U2757 (N_2757,N_2478,N_2579);
xor U2758 (N_2758,N_2418,N_2407);
and U2759 (N_2759,N_2569,N_2506);
or U2760 (N_2760,N_2540,N_2481);
and U2761 (N_2761,N_2519,N_2514);
nor U2762 (N_2762,N_2526,N_2408);
and U2763 (N_2763,N_2425,N_2599);
and U2764 (N_2764,N_2493,N_2474);
or U2765 (N_2765,N_2456,N_2597);
nor U2766 (N_2766,N_2523,N_2479);
and U2767 (N_2767,N_2483,N_2512);
xor U2768 (N_2768,N_2474,N_2544);
nand U2769 (N_2769,N_2524,N_2423);
nand U2770 (N_2770,N_2463,N_2561);
or U2771 (N_2771,N_2401,N_2558);
nand U2772 (N_2772,N_2468,N_2428);
xnor U2773 (N_2773,N_2438,N_2487);
or U2774 (N_2774,N_2407,N_2568);
nand U2775 (N_2775,N_2437,N_2529);
and U2776 (N_2776,N_2424,N_2589);
and U2777 (N_2777,N_2402,N_2536);
and U2778 (N_2778,N_2452,N_2540);
nor U2779 (N_2779,N_2491,N_2548);
and U2780 (N_2780,N_2590,N_2532);
and U2781 (N_2781,N_2525,N_2474);
and U2782 (N_2782,N_2544,N_2526);
or U2783 (N_2783,N_2432,N_2561);
and U2784 (N_2784,N_2461,N_2595);
nor U2785 (N_2785,N_2516,N_2571);
nand U2786 (N_2786,N_2422,N_2563);
and U2787 (N_2787,N_2545,N_2550);
and U2788 (N_2788,N_2596,N_2433);
or U2789 (N_2789,N_2518,N_2437);
nor U2790 (N_2790,N_2589,N_2445);
nor U2791 (N_2791,N_2548,N_2554);
and U2792 (N_2792,N_2458,N_2431);
xor U2793 (N_2793,N_2478,N_2453);
xor U2794 (N_2794,N_2437,N_2567);
or U2795 (N_2795,N_2576,N_2530);
nand U2796 (N_2796,N_2419,N_2451);
xor U2797 (N_2797,N_2431,N_2560);
and U2798 (N_2798,N_2513,N_2594);
nand U2799 (N_2799,N_2413,N_2506);
nor U2800 (N_2800,N_2766,N_2749);
nor U2801 (N_2801,N_2797,N_2673);
nand U2802 (N_2802,N_2646,N_2635);
or U2803 (N_2803,N_2779,N_2736);
or U2804 (N_2804,N_2791,N_2771);
and U2805 (N_2805,N_2618,N_2627);
xor U2806 (N_2806,N_2704,N_2742);
xor U2807 (N_2807,N_2665,N_2664);
nor U2808 (N_2808,N_2645,N_2757);
xnor U2809 (N_2809,N_2753,N_2686);
nor U2810 (N_2810,N_2726,N_2649);
and U2811 (N_2811,N_2734,N_2630);
xnor U2812 (N_2812,N_2624,N_2735);
and U2813 (N_2813,N_2617,N_2681);
or U2814 (N_2814,N_2751,N_2728);
or U2815 (N_2815,N_2731,N_2659);
or U2816 (N_2816,N_2651,N_2746);
nor U2817 (N_2817,N_2705,N_2614);
nand U2818 (N_2818,N_2677,N_2756);
nand U2819 (N_2819,N_2615,N_2729);
nor U2820 (N_2820,N_2698,N_2701);
nor U2821 (N_2821,N_2727,N_2653);
nor U2822 (N_2822,N_2755,N_2773);
nor U2823 (N_2823,N_2619,N_2752);
or U2824 (N_2824,N_2777,N_2616);
nor U2825 (N_2825,N_2785,N_2693);
xor U2826 (N_2826,N_2781,N_2603);
xnor U2827 (N_2827,N_2715,N_2765);
nand U2828 (N_2828,N_2798,N_2799);
and U2829 (N_2829,N_2625,N_2789);
nand U2830 (N_2830,N_2720,N_2759);
xnor U2831 (N_2831,N_2682,N_2638);
nor U2832 (N_2832,N_2769,N_2600);
nor U2833 (N_2833,N_2655,N_2606);
nand U2834 (N_2834,N_2629,N_2744);
nand U2835 (N_2835,N_2671,N_2633);
and U2836 (N_2836,N_2611,N_2763);
xor U2837 (N_2837,N_2709,N_2652);
and U2838 (N_2838,N_2634,N_2691);
xor U2839 (N_2839,N_2708,N_2672);
nand U2840 (N_2840,N_2641,N_2764);
nor U2841 (N_2841,N_2737,N_2724);
and U2842 (N_2842,N_2605,N_2702);
xor U2843 (N_2843,N_2761,N_2644);
nor U2844 (N_2844,N_2772,N_2620);
xor U2845 (N_2845,N_2741,N_2748);
nand U2846 (N_2846,N_2788,N_2666);
nand U2847 (N_2847,N_2722,N_2662);
nand U2848 (N_2848,N_2739,N_2784);
nor U2849 (N_2849,N_2783,N_2675);
nor U2850 (N_2850,N_2707,N_2657);
nand U2851 (N_2851,N_2695,N_2639);
nand U2852 (N_2852,N_2650,N_2713);
nor U2853 (N_2853,N_2740,N_2621);
nand U2854 (N_2854,N_2636,N_2745);
nor U2855 (N_2855,N_2714,N_2775);
nand U2856 (N_2856,N_2626,N_2623);
and U2857 (N_2857,N_2692,N_2793);
and U2858 (N_2858,N_2654,N_2703);
xnor U2859 (N_2859,N_2712,N_2706);
and U2860 (N_2860,N_2792,N_2632);
xor U2861 (N_2861,N_2684,N_2679);
xnor U2862 (N_2862,N_2747,N_2725);
xnor U2863 (N_2863,N_2774,N_2609);
and U2864 (N_2864,N_2710,N_2676);
nor U2865 (N_2865,N_2640,N_2648);
nor U2866 (N_2866,N_2670,N_2796);
nor U2867 (N_2867,N_2663,N_2719);
and U2868 (N_2868,N_2667,N_2711);
or U2869 (N_2869,N_2697,N_2656);
nand U2870 (N_2870,N_2754,N_2685);
and U2871 (N_2871,N_2612,N_2628);
nand U2872 (N_2872,N_2718,N_2699);
xor U2873 (N_2873,N_2782,N_2680);
or U2874 (N_2874,N_2601,N_2608);
xor U2875 (N_2875,N_2758,N_2700);
nor U2876 (N_2876,N_2658,N_2716);
nor U2877 (N_2877,N_2668,N_2794);
nand U2878 (N_2878,N_2787,N_2690);
nand U2879 (N_2879,N_2750,N_2694);
and U2880 (N_2880,N_2767,N_2732);
or U2881 (N_2881,N_2760,N_2669);
nand U2882 (N_2882,N_2613,N_2683);
nor U2883 (N_2883,N_2786,N_2642);
and U2884 (N_2884,N_2778,N_2643);
xor U2885 (N_2885,N_2660,N_2602);
and U2886 (N_2886,N_2743,N_2795);
or U2887 (N_2887,N_2790,N_2610);
nand U2888 (N_2888,N_2674,N_2762);
nand U2889 (N_2889,N_2717,N_2723);
and U2890 (N_2890,N_2780,N_2776);
nand U2891 (N_2891,N_2688,N_2733);
nand U2892 (N_2892,N_2622,N_2738);
nor U2893 (N_2893,N_2637,N_2604);
or U2894 (N_2894,N_2607,N_2647);
nand U2895 (N_2895,N_2730,N_2687);
nand U2896 (N_2896,N_2661,N_2631);
or U2897 (N_2897,N_2696,N_2689);
nand U2898 (N_2898,N_2768,N_2678);
or U2899 (N_2899,N_2721,N_2770);
or U2900 (N_2900,N_2755,N_2737);
and U2901 (N_2901,N_2702,N_2782);
nand U2902 (N_2902,N_2792,N_2718);
nor U2903 (N_2903,N_2758,N_2799);
and U2904 (N_2904,N_2719,N_2632);
and U2905 (N_2905,N_2678,N_2706);
nand U2906 (N_2906,N_2703,N_2781);
nor U2907 (N_2907,N_2773,N_2725);
xnor U2908 (N_2908,N_2775,N_2626);
and U2909 (N_2909,N_2669,N_2750);
nand U2910 (N_2910,N_2737,N_2680);
nand U2911 (N_2911,N_2615,N_2654);
nand U2912 (N_2912,N_2749,N_2600);
nor U2913 (N_2913,N_2777,N_2765);
nand U2914 (N_2914,N_2735,N_2661);
nand U2915 (N_2915,N_2767,N_2722);
nor U2916 (N_2916,N_2656,N_2670);
and U2917 (N_2917,N_2786,N_2757);
or U2918 (N_2918,N_2798,N_2667);
nand U2919 (N_2919,N_2703,N_2660);
nand U2920 (N_2920,N_2796,N_2766);
xor U2921 (N_2921,N_2719,N_2739);
and U2922 (N_2922,N_2617,N_2696);
nor U2923 (N_2923,N_2786,N_2713);
or U2924 (N_2924,N_2703,N_2796);
and U2925 (N_2925,N_2646,N_2626);
nor U2926 (N_2926,N_2690,N_2645);
or U2927 (N_2927,N_2668,N_2685);
or U2928 (N_2928,N_2686,N_2682);
nor U2929 (N_2929,N_2722,N_2695);
and U2930 (N_2930,N_2739,N_2658);
or U2931 (N_2931,N_2642,N_2608);
nand U2932 (N_2932,N_2656,N_2741);
or U2933 (N_2933,N_2612,N_2631);
xor U2934 (N_2934,N_2672,N_2707);
and U2935 (N_2935,N_2756,N_2769);
xnor U2936 (N_2936,N_2794,N_2709);
nor U2937 (N_2937,N_2671,N_2674);
xor U2938 (N_2938,N_2612,N_2604);
and U2939 (N_2939,N_2781,N_2629);
nand U2940 (N_2940,N_2729,N_2633);
xor U2941 (N_2941,N_2656,N_2639);
xor U2942 (N_2942,N_2604,N_2693);
nand U2943 (N_2943,N_2752,N_2710);
nand U2944 (N_2944,N_2766,N_2625);
or U2945 (N_2945,N_2633,N_2647);
nor U2946 (N_2946,N_2731,N_2624);
xor U2947 (N_2947,N_2658,N_2786);
nand U2948 (N_2948,N_2769,N_2665);
and U2949 (N_2949,N_2649,N_2749);
and U2950 (N_2950,N_2678,N_2742);
xor U2951 (N_2951,N_2648,N_2714);
and U2952 (N_2952,N_2692,N_2600);
and U2953 (N_2953,N_2645,N_2776);
or U2954 (N_2954,N_2772,N_2712);
nand U2955 (N_2955,N_2681,N_2735);
and U2956 (N_2956,N_2674,N_2664);
nor U2957 (N_2957,N_2721,N_2724);
and U2958 (N_2958,N_2717,N_2680);
xor U2959 (N_2959,N_2773,N_2697);
or U2960 (N_2960,N_2681,N_2623);
nand U2961 (N_2961,N_2689,N_2624);
xor U2962 (N_2962,N_2645,N_2743);
and U2963 (N_2963,N_2788,N_2642);
or U2964 (N_2964,N_2757,N_2703);
nor U2965 (N_2965,N_2647,N_2774);
nand U2966 (N_2966,N_2613,N_2620);
or U2967 (N_2967,N_2792,N_2647);
or U2968 (N_2968,N_2783,N_2617);
xnor U2969 (N_2969,N_2679,N_2628);
or U2970 (N_2970,N_2685,N_2745);
and U2971 (N_2971,N_2791,N_2796);
xnor U2972 (N_2972,N_2746,N_2686);
nand U2973 (N_2973,N_2785,N_2716);
and U2974 (N_2974,N_2783,N_2759);
and U2975 (N_2975,N_2684,N_2753);
xnor U2976 (N_2976,N_2636,N_2606);
nor U2977 (N_2977,N_2685,N_2733);
xor U2978 (N_2978,N_2746,N_2654);
and U2979 (N_2979,N_2607,N_2771);
nand U2980 (N_2980,N_2717,N_2652);
xnor U2981 (N_2981,N_2790,N_2611);
and U2982 (N_2982,N_2615,N_2777);
or U2983 (N_2983,N_2796,N_2684);
and U2984 (N_2984,N_2786,N_2769);
and U2985 (N_2985,N_2603,N_2762);
nor U2986 (N_2986,N_2698,N_2726);
and U2987 (N_2987,N_2748,N_2692);
nand U2988 (N_2988,N_2617,N_2688);
or U2989 (N_2989,N_2787,N_2696);
xnor U2990 (N_2990,N_2654,N_2680);
nor U2991 (N_2991,N_2734,N_2606);
and U2992 (N_2992,N_2756,N_2688);
nor U2993 (N_2993,N_2645,N_2763);
nor U2994 (N_2994,N_2628,N_2727);
and U2995 (N_2995,N_2769,N_2682);
or U2996 (N_2996,N_2763,N_2630);
nand U2997 (N_2997,N_2700,N_2733);
xor U2998 (N_2998,N_2623,N_2774);
and U2999 (N_2999,N_2654,N_2685);
and U3000 (N_3000,N_2967,N_2878);
nand U3001 (N_3001,N_2830,N_2884);
xor U3002 (N_3002,N_2882,N_2933);
xnor U3003 (N_3003,N_2950,N_2981);
xnor U3004 (N_3004,N_2879,N_2937);
nor U3005 (N_3005,N_2996,N_2863);
or U3006 (N_3006,N_2940,N_2908);
and U3007 (N_3007,N_2998,N_2883);
nor U3008 (N_3008,N_2976,N_2954);
or U3009 (N_3009,N_2892,N_2914);
nand U3010 (N_3010,N_2887,N_2855);
xnor U3011 (N_3011,N_2849,N_2868);
nor U3012 (N_3012,N_2875,N_2971);
xnor U3013 (N_3013,N_2949,N_2886);
xor U3014 (N_3014,N_2873,N_2861);
xor U3015 (N_3015,N_2943,N_2842);
nor U3016 (N_3016,N_2989,N_2839);
nor U3017 (N_3017,N_2904,N_2815);
and U3018 (N_3018,N_2806,N_2961);
and U3019 (N_3019,N_2856,N_2959);
nand U3020 (N_3020,N_2801,N_2936);
xnor U3021 (N_3021,N_2910,N_2828);
xor U3022 (N_3022,N_2820,N_2927);
and U3023 (N_3023,N_2888,N_2941);
and U3024 (N_3024,N_2953,N_2957);
and U3025 (N_3025,N_2893,N_2935);
and U3026 (N_3026,N_2903,N_2827);
xor U3027 (N_3027,N_2979,N_2938);
xor U3028 (N_3028,N_2926,N_2930);
xor U3029 (N_3029,N_2891,N_2984);
nor U3030 (N_3030,N_2869,N_2913);
and U3031 (N_3031,N_2925,N_2966);
and U3032 (N_3032,N_2948,N_2955);
nor U3033 (N_3033,N_2972,N_2974);
or U3034 (N_3034,N_2871,N_2980);
or U3035 (N_3035,N_2947,N_2915);
nor U3036 (N_3036,N_2911,N_2991);
xor U3037 (N_3037,N_2858,N_2983);
or U3038 (N_3038,N_2951,N_2982);
nor U3039 (N_3039,N_2896,N_2866);
nand U3040 (N_3040,N_2968,N_2837);
nor U3041 (N_3041,N_2859,N_2814);
xnor U3042 (N_3042,N_2821,N_2918);
or U3043 (N_3043,N_2958,N_2919);
nor U3044 (N_3044,N_2848,N_2800);
and U3045 (N_3045,N_2822,N_2894);
nand U3046 (N_3046,N_2898,N_2928);
and U3047 (N_3047,N_2988,N_2909);
xnor U3048 (N_3048,N_2995,N_2843);
nor U3049 (N_3049,N_2877,N_2934);
and U3050 (N_3050,N_2841,N_2862);
nor U3051 (N_3051,N_2803,N_2846);
or U3052 (N_3052,N_2923,N_2900);
nor U3053 (N_3053,N_2804,N_2899);
nand U3054 (N_3054,N_2946,N_2867);
nor U3055 (N_3055,N_2870,N_2817);
xnor U3056 (N_3056,N_2876,N_2956);
nor U3057 (N_3057,N_2962,N_2992);
xnor U3058 (N_3058,N_2874,N_2844);
and U3059 (N_3059,N_2978,N_2997);
or U3060 (N_3060,N_2897,N_2872);
and U3061 (N_3061,N_2836,N_2819);
nor U3062 (N_3062,N_2853,N_2921);
xnor U3063 (N_3063,N_2902,N_2880);
nor U3064 (N_3064,N_2810,N_2999);
or U3065 (N_3065,N_2890,N_2973);
xnor U3066 (N_3066,N_2885,N_2960);
nand U3067 (N_3067,N_2929,N_2970);
nor U3068 (N_3068,N_2813,N_2823);
xnor U3069 (N_3069,N_2826,N_2977);
and U3070 (N_3070,N_2889,N_2847);
nand U3071 (N_3071,N_2952,N_2924);
nand U3072 (N_3072,N_2833,N_2805);
nand U3073 (N_3073,N_2986,N_2920);
or U3074 (N_3074,N_2964,N_2993);
and U3075 (N_3075,N_2939,N_2857);
xnor U3076 (N_3076,N_2852,N_2965);
or U3077 (N_3077,N_2945,N_2831);
nor U3078 (N_3078,N_2807,N_2864);
xor U3079 (N_3079,N_2808,N_2942);
and U3080 (N_3080,N_2985,N_2881);
nand U3081 (N_3081,N_2854,N_2922);
nor U3082 (N_3082,N_2905,N_2840);
xnor U3083 (N_3083,N_2802,N_2917);
xnor U3084 (N_3084,N_2845,N_2835);
and U3085 (N_3085,N_2812,N_2824);
nor U3086 (N_3086,N_2932,N_2816);
nand U3087 (N_3087,N_2832,N_2916);
nor U3088 (N_3088,N_2906,N_2895);
or U3089 (N_3089,N_2907,N_2825);
and U3090 (N_3090,N_2990,N_2969);
or U3091 (N_3091,N_2811,N_2829);
nand U3092 (N_3092,N_2850,N_2818);
and U3093 (N_3093,N_2963,N_2865);
nor U3094 (N_3094,N_2975,N_2809);
and U3095 (N_3095,N_2838,N_2987);
nor U3096 (N_3096,N_2851,N_2944);
xor U3097 (N_3097,N_2931,N_2901);
xnor U3098 (N_3098,N_2994,N_2860);
or U3099 (N_3099,N_2912,N_2834);
xnor U3100 (N_3100,N_2970,N_2918);
nand U3101 (N_3101,N_2989,N_2812);
or U3102 (N_3102,N_2943,N_2856);
or U3103 (N_3103,N_2939,N_2866);
or U3104 (N_3104,N_2908,N_2990);
nand U3105 (N_3105,N_2946,N_2951);
xnor U3106 (N_3106,N_2866,N_2824);
nor U3107 (N_3107,N_2958,N_2938);
or U3108 (N_3108,N_2949,N_2857);
xor U3109 (N_3109,N_2894,N_2933);
nor U3110 (N_3110,N_2951,N_2901);
nand U3111 (N_3111,N_2955,N_2821);
and U3112 (N_3112,N_2891,N_2987);
nor U3113 (N_3113,N_2857,N_2906);
nand U3114 (N_3114,N_2881,N_2937);
xor U3115 (N_3115,N_2850,N_2989);
nand U3116 (N_3116,N_2955,N_2818);
nand U3117 (N_3117,N_2926,N_2810);
nand U3118 (N_3118,N_2967,N_2973);
nand U3119 (N_3119,N_2925,N_2913);
or U3120 (N_3120,N_2985,N_2826);
or U3121 (N_3121,N_2906,N_2868);
xor U3122 (N_3122,N_2864,N_2897);
xor U3123 (N_3123,N_2897,N_2939);
xnor U3124 (N_3124,N_2977,N_2983);
nor U3125 (N_3125,N_2824,N_2977);
and U3126 (N_3126,N_2897,N_2831);
and U3127 (N_3127,N_2829,N_2897);
or U3128 (N_3128,N_2809,N_2815);
nor U3129 (N_3129,N_2882,N_2950);
nor U3130 (N_3130,N_2955,N_2949);
and U3131 (N_3131,N_2920,N_2828);
and U3132 (N_3132,N_2830,N_2874);
or U3133 (N_3133,N_2984,N_2866);
nor U3134 (N_3134,N_2999,N_2886);
xor U3135 (N_3135,N_2818,N_2883);
or U3136 (N_3136,N_2987,N_2841);
nor U3137 (N_3137,N_2802,N_2963);
xnor U3138 (N_3138,N_2878,N_2903);
nand U3139 (N_3139,N_2917,N_2838);
nor U3140 (N_3140,N_2853,N_2930);
nand U3141 (N_3141,N_2830,N_2946);
or U3142 (N_3142,N_2822,N_2984);
nor U3143 (N_3143,N_2832,N_2972);
or U3144 (N_3144,N_2809,N_2864);
nand U3145 (N_3145,N_2988,N_2834);
or U3146 (N_3146,N_2904,N_2992);
or U3147 (N_3147,N_2935,N_2945);
or U3148 (N_3148,N_2874,N_2904);
xnor U3149 (N_3149,N_2805,N_2982);
nor U3150 (N_3150,N_2852,N_2999);
nand U3151 (N_3151,N_2921,N_2852);
xor U3152 (N_3152,N_2991,N_2910);
or U3153 (N_3153,N_2849,N_2978);
nor U3154 (N_3154,N_2952,N_2893);
and U3155 (N_3155,N_2804,N_2861);
nor U3156 (N_3156,N_2910,N_2915);
nor U3157 (N_3157,N_2845,N_2951);
or U3158 (N_3158,N_2985,N_2932);
xor U3159 (N_3159,N_2973,N_2871);
nand U3160 (N_3160,N_2976,N_2982);
nand U3161 (N_3161,N_2887,N_2894);
and U3162 (N_3162,N_2875,N_2906);
and U3163 (N_3163,N_2899,N_2859);
and U3164 (N_3164,N_2918,N_2980);
or U3165 (N_3165,N_2918,N_2829);
nand U3166 (N_3166,N_2930,N_2854);
xor U3167 (N_3167,N_2802,N_2886);
xnor U3168 (N_3168,N_2935,N_2952);
or U3169 (N_3169,N_2970,N_2874);
and U3170 (N_3170,N_2981,N_2853);
nor U3171 (N_3171,N_2980,N_2974);
xnor U3172 (N_3172,N_2952,N_2832);
nand U3173 (N_3173,N_2911,N_2863);
or U3174 (N_3174,N_2983,N_2984);
and U3175 (N_3175,N_2997,N_2922);
nand U3176 (N_3176,N_2981,N_2903);
xnor U3177 (N_3177,N_2878,N_2913);
and U3178 (N_3178,N_2947,N_2974);
nand U3179 (N_3179,N_2915,N_2997);
nand U3180 (N_3180,N_2898,N_2982);
nor U3181 (N_3181,N_2930,N_2857);
and U3182 (N_3182,N_2994,N_2911);
nor U3183 (N_3183,N_2802,N_2996);
xor U3184 (N_3184,N_2889,N_2860);
xor U3185 (N_3185,N_2849,N_2862);
and U3186 (N_3186,N_2942,N_2987);
xnor U3187 (N_3187,N_2846,N_2898);
xor U3188 (N_3188,N_2997,N_2927);
xor U3189 (N_3189,N_2902,N_2913);
or U3190 (N_3190,N_2811,N_2934);
nor U3191 (N_3191,N_2846,N_2880);
nor U3192 (N_3192,N_2926,N_2850);
xnor U3193 (N_3193,N_2972,N_2920);
and U3194 (N_3194,N_2973,N_2800);
xnor U3195 (N_3195,N_2938,N_2994);
nor U3196 (N_3196,N_2985,N_2821);
nor U3197 (N_3197,N_2981,N_2910);
or U3198 (N_3198,N_2904,N_2923);
nor U3199 (N_3199,N_2920,N_2968);
or U3200 (N_3200,N_3106,N_3169);
nand U3201 (N_3201,N_3146,N_3161);
nand U3202 (N_3202,N_3156,N_3090);
or U3203 (N_3203,N_3126,N_3071);
nand U3204 (N_3204,N_3187,N_3048);
or U3205 (N_3205,N_3148,N_3099);
nor U3206 (N_3206,N_3180,N_3149);
and U3207 (N_3207,N_3107,N_3085);
nor U3208 (N_3208,N_3007,N_3104);
xor U3209 (N_3209,N_3109,N_3134);
or U3210 (N_3210,N_3191,N_3153);
or U3211 (N_3211,N_3022,N_3097);
xor U3212 (N_3212,N_3178,N_3130);
nor U3213 (N_3213,N_3006,N_3133);
and U3214 (N_3214,N_3021,N_3036);
or U3215 (N_3215,N_3159,N_3184);
or U3216 (N_3216,N_3186,N_3074);
nor U3217 (N_3217,N_3035,N_3073);
xor U3218 (N_3218,N_3183,N_3162);
or U3219 (N_3219,N_3112,N_3100);
nor U3220 (N_3220,N_3078,N_3120);
or U3221 (N_3221,N_3033,N_3166);
nor U3222 (N_3222,N_3151,N_3194);
and U3223 (N_3223,N_3055,N_3069);
nor U3224 (N_3224,N_3119,N_3038);
nor U3225 (N_3225,N_3131,N_3094);
or U3226 (N_3226,N_3102,N_3014);
or U3227 (N_3227,N_3111,N_3056);
nor U3228 (N_3228,N_3072,N_3052);
or U3229 (N_3229,N_3011,N_3193);
xnor U3230 (N_3230,N_3020,N_3128);
or U3231 (N_3231,N_3057,N_3028);
nand U3232 (N_3232,N_3061,N_3173);
or U3233 (N_3233,N_3122,N_3096);
nor U3234 (N_3234,N_3049,N_3092);
or U3235 (N_3235,N_3076,N_3198);
xor U3236 (N_3236,N_3140,N_3155);
and U3237 (N_3237,N_3070,N_3065);
xor U3238 (N_3238,N_3045,N_3044);
nor U3239 (N_3239,N_3087,N_3172);
or U3240 (N_3240,N_3103,N_3095);
nand U3241 (N_3241,N_3182,N_3117);
nand U3242 (N_3242,N_3135,N_3143);
or U3243 (N_3243,N_3129,N_3026);
nor U3244 (N_3244,N_3137,N_3176);
and U3245 (N_3245,N_3029,N_3171);
or U3246 (N_3246,N_3115,N_3123);
and U3247 (N_3247,N_3093,N_3145);
and U3248 (N_3248,N_3042,N_3031);
and U3249 (N_3249,N_3152,N_3017);
xnor U3250 (N_3250,N_3110,N_3060);
and U3251 (N_3251,N_3077,N_3105);
nand U3252 (N_3252,N_3003,N_3098);
xor U3253 (N_3253,N_3116,N_3142);
or U3254 (N_3254,N_3064,N_3136);
and U3255 (N_3255,N_3027,N_3015);
nor U3256 (N_3256,N_3144,N_3068);
nand U3257 (N_3257,N_3139,N_3165);
nand U3258 (N_3258,N_3091,N_3185);
and U3259 (N_3259,N_3158,N_3010);
or U3260 (N_3260,N_3199,N_3192);
or U3261 (N_3261,N_3001,N_3088);
xor U3262 (N_3262,N_3179,N_3127);
xor U3263 (N_3263,N_3188,N_3177);
nor U3264 (N_3264,N_3062,N_3150);
xor U3265 (N_3265,N_3082,N_3004);
and U3266 (N_3266,N_3034,N_3118);
nor U3267 (N_3267,N_3018,N_3089);
and U3268 (N_3268,N_3157,N_3164);
xnor U3269 (N_3269,N_3000,N_3121);
or U3270 (N_3270,N_3113,N_3047);
or U3271 (N_3271,N_3012,N_3125);
xnor U3272 (N_3272,N_3174,N_3080);
and U3273 (N_3273,N_3075,N_3040);
and U3274 (N_3274,N_3163,N_3086);
and U3275 (N_3275,N_3050,N_3114);
and U3276 (N_3276,N_3170,N_3175);
nand U3277 (N_3277,N_3053,N_3016);
xnor U3278 (N_3278,N_3167,N_3009);
xor U3279 (N_3279,N_3066,N_3005);
xor U3280 (N_3280,N_3160,N_3124);
nand U3281 (N_3281,N_3030,N_3101);
or U3282 (N_3282,N_3002,N_3141);
xor U3283 (N_3283,N_3046,N_3197);
and U3284 (N_3284,N_3043,N_3168);
xnor U3285 (N_3285,N_3008,N_3132);
xor U3286 (N_3286,N_3037,N_3025);
and U3287 (N_3287,N_3189,N_3063);
nor U3288 (N_3288,N_3195,N_3023);
xnor U3289 (N_3289,N_3054,N_3181);
nor U3290 (N_3290,N_3013,N_3024);
nand U3291 (N_3291,N_3138,N_3083);
and U3292 (N_3292,N_3067,N_3019);
or U3293 (N_3293,N_3079,N_3041);
xor U3294 (N_3294,N_3039,N_3108);
nor U3295 (N_3295,N_3081,N_3154);
nor U3296 (N_3296,N_3032,N_3059);
or U3297 (N_3297,N_3084,N_3190);
xnor U3298 (N_3298,N_3147,N_3058);
nor U3299 (N_3299,N_3051,N_3196);
or U3300 (N_3300,N_3189,N_3115);
and U3301 (N_3301,N_3132,N_3022);
nand U3302 (N_3302,N_3041,N_3010);
nand U3303 (N_3303,N_3191,N_3164);
nand U3304 (N_3304,N_3003,N_3047);
nor U3305 (N_3305,N_3024,N_3125);
nor U3306 (N_3306,N_3118,N_3183);
or U3307 (N_3307,N_3197,N_3021);
and U3308 (N_3308,N_3193,N_3089);
or U3309 (N_3309,N_3102,N_3085);
or U3310 (N_3310,N_3096,N_3107);
nor U3311 (N_3311,N_3000,N_3196);
nor U3312 (N_3312,N_3131,N_3148);
nor U3313 (N_3313,N_3007,N_3161);
xnor U3314 (N_3314,N_3145,N_3097);
xnor U3315 (N_3315,N_3125,N_3089);
nor U3316 (N_3316,N_3151,N_3092);
nor U3317 (N_3317,N_3006,N_3114);
nor U3318 (N_3318,N_3071,N_3106);
xnor U3319 (N_3319,N_3055,N_3188);
and U3320 (N_3320,N_3175,N_3196);
or U3321 (N_3321,N_3195,N_3183);
nand U3322 (N_3322,N_3152,N_3032);
and U3323 (N_3323,N_3052,N_3178);
and U3324 (N_3324,N_3077,N_3053);
nor U3325 (N_3325,N_3048,N_3179);
and U3326 (N_3326,N_3122,N_3002);
or U3327 (N_3327,N_3137,N_3110);
xor U3328 (N_3328,N_3136,N_3129);
nand U3329 (N_3329,N_3047,N_3122);
nor U3330 (N_3330,N_3114,N_3055);
or U3331 (N_3331,N_3000,N_3166);
nor U3332 (N_3332,N_3135,N_3053);
xnor U3333 (N_3333,N_3141,N_3191);
xnor U3334 (N_3334,N_3002,N_3011);
nor U3335 (N_3335,N_3072,N_3004);
nand U3336 (N_3336,N_3002,N_3151);
xor U3337 (N_3337,N_3181,N_3155);
and U3338 (N_3338,N_3012,N_3048);
or U3339 (N_3339,N_3134,N_3164);
or U3340 (N_3340,N_3190,N_3046);
nor U3341 (N_3341,N_3081,N_3178);
and U3342 (N_3342,N_3176,N_3100);
nand U3343 (N_3343,N_3184,N_3074);
and U3344 (N_3344,N_3110,N_3015);
nand U3345 (N_3345,N_3191,N_3145);
nor U3346 (N_3346,N_3189,N_3199);
nor U3347 (N_3347,N_3039,N_3091);
nand U3348 (N_3348,N_3102,N_3023);
nand U3349 (N_3349,N_3095,N_3132);
xnor U3350 (N_3350,N_3141,N_3172);
and U3351 (N_3351,N_3128,N_3173);
xor U3352 (N_3352,N_3121,N_3137);
or U3353 (N_3353,N_3040,N_3131);
nor U3354 (N_3354,N_3007,N_3138);
xor U3355 (N_3355,N_3086,N_3159);
xor U3356 (N_3356,N_3017,N_3052);
or U3357 (N_3357,N_3068,N_3003);
nor U3358 (N_3358,N_3045,N_3016);
nand U3359 (N_3359,N_3153,N_3110);
nand U3360 (N_3360,N_3041,N_3103);
xnor U3361 (N_3361,N_3187,N_3154);
and U3362 (N_3362,N_3190,N_3138);
nand U3363 (N_3363,N_3156,N_3095);
nor U3364 (N_3364,N_3012,N_3101);
nand U3365 (N_3365,N_3001,N_3180);
and U3366 (N_3366,N_3034,N_3064);
or U3367 (N_3367,N_3190,N_3073);
and U3368 (N_3368,N_3062,N_3161);
nor U3369 (N_3369,N_3026,N_3102);
nand U3370 (N_3370,N_3053,N_3007);
nor U3371 (N_3371,N_3092,N_3026);
nand U3372 (N_3372,N_3168,N_3076);
xnor U3373 (N_3373,N_3025,N_3005);
and U3374 (N_3374,N_3117,N_3101);
nand U3375 (N_3375,N_3028,N_3092);
or U3376 (N_3376,N_3065,N_3108);
nand U3377 (N_3377,N_3007,N_3157);
xor U3378 (N_3378,N_3017,N_3080);
or U3379 (N_3379,N_3196,N_3018);
nand U3380 (N_3380,N_3137,N_3030);
nand U3381 (N_3381,N_3098,N_3087);
xor U3382 (N_3382,N_3034,N_3123);
nor U3383 (N_3383,N_3112,N_3056);
nand U3384 (N_3384,N_3016,N_3092);
or U3385 (N_3385,N_3189,N_3009);
or U3386 (N_3386,N_3048,N_3071);
nor U3387 (N_3387,N_3113,N_3064);
nand U3388 (N_3388,N_3145,N_3156);
nand U3389 (N_3389,N_3125,N_3128);
nor U3390 (N_3390,N_3065,N_3021);
xnor U3391 (N_3391,N_3157,N_3075);
or U3392 (N_3392,N_3037,N_3138);
xor U3393 (N_3393,N_3078,N_3067);
nor U3394 (N_3394,N_3119,N_3043);
nand U3395 (N_3395,N_3150,N_3186);
or U3396 (N_3396,N_3179,N_3117);
xnor U3397 (N_3397,N_3074,N_3183);
xnor U3398 (N_3398,N_3177,N_3127);
nand U3399 (N_3399,N_3187,N_3059);
nor U3400 (N_3400,N_3204,N_3317);
or U3401 (N_3401,N_3324,N_3339);
nand U3402 (N_3402,N_3252,N_3312);
xor U3403 (N_3403,N_3332,N_3266);
or U3404 (N_3404,N_3237,N_3265);
and U3405 (N_3405,N_3211,N_3370);
or U3406 (N_3406,N_3248,N_3257);
or U3407 (N_3407,N_3208,N_3256);
or U3408 (N_3408,N_3271,N_3285);
xor U3409 (N_3409,N_3336,N_3367);
nor U3410 (N_3410,N_3360,N_3251);
nand U3411 (N_3411,N_3361,N_3222);
nand U3412 (N_3412,N_3281,N_3386);
nand U3413 (N_3413,N_3287,N_3348);
nand U3414 (N_3414,N_3245,N_3286);
nor U3415 (N_3415,N_3225,N_3246);
nor U3416 (N_3416,N_3275,N_3309);
nand U3417 (N_3417,N_3331,N_3234);
nand U3418 (N_3418,N_3220,N_3314);
or U3419 (N_3419,N_3319,N_3368);
nor U3420 (N_3420,N_3231,N_3372);
or U3421 (N_3421,N_3349,N_3235);
and U3422 (N_3422,N_3294,N_3201);
nor U3423 (N_3423,N_3200,N_3350);
nor U3424 (N_3424,N_3293,N_3274);
nor U3425 (N_3425,N_3276,N_3303);
or U3426 (N_3426,N_3295,N_3392);
and U3427 (N_3427,N_3379,N_3329);
nand U3428 (N_3428,N_3226,N_3206);
and U3429 (N_3429,N_3270,N_3327);
or U3430 (N_3430,N_3255,N_3284);
and U3431 (N_3431,N_3279,N_3316);
nor U3432 (N_3432,N_3377,N_3202);
xor U3433 (N_3433,N_3346,N_3359);
nand U3434 (N_3434,N_3278,N_3291);
and U3435 (N_3435,N_3352,N_3355);
nand U3436 (N_3436,N_3306,N_3300);
xnor U3437 (N_3437,N_3304,N_3390);
nand U3438 (N_3438,N_3337,N_3388);
nand U3439 (N_3439,N_3260,N_3366);
xor U3440 (N_3440,N_3243,N_3362);
or U3441 (N_3441,N_3269,N_3325);
nand U3442 (N_3442,N_3399,N_3207);
and U3443 (N_3443,N_3383,N_3322);
nand U3444 (N_3444,N_3321,N_3380);
nand U3445 (N_3445,N_3356,N_3333);
nand U3446 (N_3446,N_3283,N_3272);
or U3447 (N_3447,N_3232,N_3262);
nand U3448 (N_3448,N_3323,N_3363);
or U3449 (N_3449,N_3229,N_3347);
nor U3450 (N_3450,N_3263,N_3254);
xnor U3451 (N_3451,N_3259,N_3341);
xnor U3452 (N_3452,N_3223,N_3230);
or U3453 (N_3453,N_3330,N_3240);
or U3454 (N_3454,N_3344,N_3369);
or U3455 (N_3455,N_3374,N_3311);
nor U3456 (N_3456,N_3389,N_3233);
nor U3457 (N_3457,N_3268,N_3296);
nor U3458 (N_3458,N_3395,N_3318);
or U3459 (N_3459,N_3241,N_3334);
nor U3460 (N_3460,N_3228,N_3313);
and U3461 (N_3461,N_3290,N_3375);
nand U3462 (N_3462,N_3282,N_3217);
or U3463 (N_3463,N_3289,N_3247);
and U3464 (N_3464,N_3381,N_3342);
nand U3465 (N_3465,N_3326,N_3373);
or U3466 (N_3466,N_3299,N_3242);
nor U3467 (N_3467,N_3354,N_3305);
nand U3468 (N_3468,N_3371,N_3219);
xor U3469 (N_3469,N_3273,N_3236);
xnor U3470 (N_3470,N_3357,N_3301);
nand U3471 (N_3471,N_3239,N_3343);
nand U3472 (N_3472,N_3218,N_3398);
or U3473 (N_3473,N_3213,N_3280);
and U3474 (N_3474,N_3210,N_3351);
or U3475 (N_3475,N_3244,N_3267);
or U3476 (N_3476,N_3203,N_3315);
nor U3477 (N_3477,N_3358,N_3387);
and U3478 (N_3478,N_3382,N_3353);
nand U3479 (N_3479,N_3288,N_3238);
xnor U3480 (N_3480,N_3209,N_3385);
xnor U3481 (N_3481,N_3297,N_3216);
xnor U3482 (N_3482,N_3397,N_3340);
or U3483 (N_3483,N_3298,N_3384);
nand U3484 (N_3484,N_3365,N_3264);
or U3485 (N_3485,N_3364,N_3215);
nand U3486 (N_3486,N_3224,N_3292);
or U3487 (N_3487,N_3376,N_3328);
xnor U3488 (N_3488,N_3258,N_3310);
xor U3489 (N_3489,N_3345,N_3302);
nor U3490 (N_3490,N_3335,N_3308);
nand U3491 (N_3491,N_3227,N_3396);
and U3492 (N_3492,N_3205,N_3250);
nor U3493 (N_3493,N_3277,N_3253);
nor U3494 (N_3494,N_3307,N_3320);
or U3495 (N_3495,N_3393,N_3214);
nand U3496 (N_3496,N_3391,N_3261);
or U3497 (N_3497,N_3394,N_3378);
or U3498 (N_3498,N_3249,N_3221);
and U3499 (N_3499,N_3212,N_3338);
nor U3500 (N_3500,N_3331,N_3279);
nand U3501 (N_3501,N_3206,N_3300);
xor U3502 (N_3502,N_3337,N_3294);
nand U3503 (N_3503,N_3290,N_3297);
nor U3504 (N_3504,N_3361,N_3329);
xor U3505 (N_3505,N_3358,N_3231);
or U3506 (N_3506,N_3279,N_3349);
nand U3507 (N_3507,N_3263,N_3265);
nor U3508 (N_3508,N_3280,N_3235);
nand U3509 (N_3509,N_3240,N_3349);
nand U3510 (N_3510,N_3249,N_3245);
or U3511 (N_3511,N_3201,N_3228);
nand U3512 (N_3512,N_3355,N_3311);
and U3513 (N_3513,N_3309,N_3386);
or U3514 (N_3514,N_3297,N_3302);
or U3515 (N_3515,N_3375,N_3263);
or U3516 (N_3516,N_3305,N_3346);
or U3517 (N_3517,N_3392,N_3245);
and U3518 (N_3518,N_3327,N_3355);
and U3519 (N_3519,N_3349,N_3357);
nand U3520 (N_3520,N_3348,N_3257);
nor U3521 (N_3521,N_3389,N_3378);
nor U3522 (N_3522,N_3251,N_3391);
nand U3523 (N_3523,N_3390,N_3236);
xor U3524 (N_3524,N_3344,N_3282);
or U3525 (N_3525,N_3360,N_3362);
xor U3526 (N_3526,N_3385,N_3371);
nand U3527 (N_3527,N_3230,N_3247);
or U3528 (N_3528,N_3290,N_3345);
nor U3529 (N_3529,N_3227,N_3261);
or U3530 (N_3530,N_3263,N_3270);
nor U3531 (N_3531,N_3324,N_3351);
xnor U3532 (N_3532,N_3368,N_3377);
nand U3533 (N_3533,N_3383,N_3395);
and U3534 (N_3534,N_3327,N_3235);
and U3535 (N_3535,N_3207,N_3223);
or U3536 (N_3536,N_3355,N_3211);
nand U3537 (N_3537,N_3212,N_3380);
nor U3538 (N_3538,N_3318,N_3250);
nand U3539 (N_3539,N_3315,N_3217);
nor U3540 (N_3540,N_3294,N_3310);
and U3541 (N_3541,N_3334,N_3337);
or U3542 (N_3542,N_3202,N_3222);
and U3543 (N_3543,N_3315,N_3366);
or U3544 (N_3544,N_3286,N_3335);
nand U3545 (N_3545,N_3247,N_3243);
and U3546 (N_3546,N_3211,N_3391);
and U3547 (N_3547,N_3251,N_3332);
nand U3548 (N_3548,N_3255,N_3360);
nand U3549 (N_3549,N_3234,N_3205);
nor U3550 (N_3550,N_3228,N_3231);
xor U3551 (N_3551,N_3372,N_3258);
nor U3552 (N_3552,N_3312,N_3352);
or U3553 (N_3553,N_3228,N_3272);
nand U3554 (N_3554,N_3211,N_3250);
nor U3555 (N_3555,N_3208,N_3395);
and U3556 (N_3556,N_3204,N_3276);
or U3557 (N_3557,N_3252,N_3311);
nor U3558 (N_3558,N_3209,N_3220);
nand U3559 (N_3559,N_3288,N_3337);
nand U3560 (N_3560,N_3330,N_3231);
and U3561 (N_3561,N_3373,N_3279);
nand U3562 (N_3562,N_3282,N_3379);
nor U3563 (N_3563,N_3323,N_3263);
nand U3564 (N_3564,N_3305,N_3392);
xnor U3565 (N_3565,N_3277,N_3216);
xnor U3566 (N_3566,N_3248,N_3297);
and U3567 (N_3567,N_3332,N_3364);
and U3568 (N_3568,N_3282,N_3210);
nand U3569 (N_3569,N_3218,N_3217);
and U3570 (N_3570,N_3323,N_3340);
nand U3571 (N_3571,N_3220,N_3207);
and U3572 (N_3572,N_3320,N_3239);
xor U3573 (N_3573,N_3212,N_3237);
xor U3574 (N_3574,N_3204,N_3369);
or U3575 (N_3575,N_3267,N_3217);
and U3576 (N_3576,N_3363,N_3230);
xor U3577 (N_3577,N_3313,N_3289);
xnor U3578 (N_3578,N_3231,N_3399);
nor U3579 (N_3579,N_3312,N_3357);
xnor U3580 (N_3580,N_3326,N_3334);
and U3581 (N_3581,N_3264,N_3278);
and U3582 (N_3582,N_3253,N_3293);
nor U3583 (N_3583,N_3391,N_3396);
nand U3584 (N_3584,N_3397,N_3241);
nand U3585 (N_3585,N_3240,N_3226);
nor U3586 (N_3586,N_3323,N_3288);
and U3587 (N_3587,N_3291,N_3334);
xnor U3588 (N_3588,N_3396,N_3220);
xor U3589 (N_3589,N_3394,N_3257);
and U3590 (N_3590,N_3360,N_3373);
or U3591 (N_3591,N_3398,N_3337);
xnor U3592 (N_3592,N_3216,N_3352);
and U3593 (N_3593,N_3309,N_3264);
or U3594 (N_3594,N_3260,N_3292);
or U3595 (N_3595,N_3290,N_3241);
and U3596 (N_3596,N_3341,N_3329);
nor U3597 (N_3597,N_3341,N_3305);
nand U3598 (N_3598,N_3323,N_3339);
xor U3599 (N_3599,N_3222,N_3342);
nor U3600 (N_3600,N_3411,N_3584);
xor U3601 (N_3601,N_3470,N_3593);
and U3602 (N_3602,N_3433,N_3421);
nor U3603 (N_3603,N_3521,N_3468);
nor U3604 (N_3604,N_3402,N_3588);
nand U3605 (N_3605,N_3479,N_3507);
xnor U3606 (N_3606,N_3571,N_3419);
nand U3607 (N_3607,N_3573,N_3474);
nand U3608 (N_3608,N_3489,N_3485);
xnor U3609 (N_3609,N_3455,N_3579);
or U3610 (N_3610,N_3541,N_3523);
and U3611 (N_3611,N_3502,N_3425);
nand U3612 (N_3612,N_3515,N_3565);
nor U3613 (N_3613,N_3572,N_3475);
nand U3614 (N_3614,N_3436,N_3553);
or U3615 (N_3615,N_3430,N_3492);
or U3616 (N_3616,N_3554,N_3415);
nand U3617 (N_3617,N_3536,N_3514);
xor U3618 (N_3618,N_3578,N_3528);
xnor U3619 (N_3619,N_3484,N_3451);
and U3620 (N_3620,N_3452,N_3459);
xor U3621 (N_3621,N_3444,N_3517);
nand U3622 (N_3622,N_3574,N_3581);
nand U3623 (N_3623,N_3405,N_3486);
and U3624 (N_3624,N_3499,N_3560);
xnor U3625 (N_3625,N_3465,N_3491);
and U3626 (N_3626,N_3568,N_3466);
or U3627 (N_3627,N_3490,N_3567);
nand U3628 (N_3628,N_3413,N_3500);
xnor U3629 (N_3629,N_3580,N_3535);
xnor U3630 (N_3630,N_3527,N_3570);
nor U3631 (N_3631,N_3562,N_3495);
or U3632 (N_3632,N_3542,N_3561);
nor U3633 (N_3633,N_3464,N_3414);
xnor U3634 (N_3634,N_3446,N_3529);
nand U3635 (N_3635,N_3587,N_3458);
and U3636 (N_3636,N_3505,N_3556);
nor U3637 (N_3637,N_3538,N_3540);
or U3638 (N_3638,N_3469,N_3438);
nand U3639 (N_3639,N_3467,N_3422);
or U3640 (N_3640,N_3482,N_3597);
xnor U3641 (N_3641,N_3497,N_3437);
nor U3642 (N_3642,N_3555,N_3478);
and U3643 (N_3643,N_3428,N_3552);
and U3644 (N_3644,N_3524,N_3439);
and U3645 (N_3645,N_3462,N_3404);
nor U3646 (N_3646,N_3582,N_3598);
xnor U3647 (N_3647,N_3412,N_3432);
nor U3648 (N_3648,N_3449,N_3551);
nand U3649 (N_3649,N_3576,N_3595);
and U3650 (N_3650,N_3481,N_3532);
xnor U3651 (N_3651,N_3501,N_3416);
nor U3652 (N_3652,N_3589,N_3418);
or U3653 (N_3653,N_3487,N_3518);
nor U3654 (N_3654,N_3577,N_3423);
xor U3655 (N_3655,N_3457,N_3509);
nor U3656 (N_3656,N_3592,N_3558);
or U3657 (N_3657,N_3520,N_3448);
nand U3658 (N_3658,N_3543,N_3410);
and U3659 (N_3659,N_3401,N_3559);
nor U3660 (N_3660,N_3454,N_3534);
nor U3661 (N_3661,N_3594,N_3566);
or U3662 (N_3662,N_3434,N_3511);
and U3663 (N_3663,N_3522,N_3488);
and U3664 (N_3664,N_3546,N_3563);
or U3665 (N_3665,N_3461,N_3493);
nor U3666 (N_3666,N_3525,N_3549);
or U3667 (N_3667,N_3503,N_3583);
xor U3668 (N_3668,N_3506,N_3564);
or U3669 (N_3669,N_3441,N_3427);
nor U3670 (N_3670,N_3477,N_3591);
and U3671 (N_3671,N_3408,N_3443);
or U3672 (N_3672,N_3400,N_3512);
or U3673 (N_3673,N_3429,N_3575);
or U3674 (N_3674,N_3460,N_3453);
nor U3675 (N_3675,N_3456,N_3406);
nor U3676 (N_3676,N_3557,N_3409);
nor U3677 (N_3677,N_3513,N_3537);
and U3678 (N_3678,N_3516,N_3585);
and U3679 (N_3679,N_3545,N_3407);
and U3680 (N_3680,N_3476,N_3420);
or U3681 (N_3681,N_3544,N_3445);
nor U3682 (N_3682,N_3526,N_3510);
and U3683 (N_3683,N_3508,N_3548);
xor U3684 (N_3684,N_3450,N_3440);
nor U3685 (N_3685,N_3473,N_3403);
nor U3686 (N_3686,N_3569,N_3463);
xnor U3687 (N_3687,N_3586,N_3426);
nor U3688 (N_3688,N_3539,N_3431);
nand U3689 (N_3689,N_3424,N_3531);
nand U3690 (N_3690,N_3504,N_3550);
xor U3691 (N_3691,N_3483,N_3494);
or U3692 (N_3692,N_3435,N_3442);
nand U3693 (N_3693,N_3417,N_3596);
or U3694 (N_3694,N_3599,N_3496);
nor U3695 (N_3695,N_3547,N_3533);
nor U3696 (N_3696,N_3471,N_3590);
and U3697 (N_3697,N_3498,N_3519);
xnor U3698 (N_3698,N_3447,N_3530);
nor U3699 (N_3699,N_3472,N_3480);
nor U3700 (N_3700,N_3580,N_3507);
xnor U3701 (N_3701,N_3462,N_3490);
or U3702 (N_3702,N_3411,N_3580);
xor U3703 (N_3703,N_3479,N_3509);
and U3704 (N_3704,N_3439,N_3508);
or U3705 (N_3705,N_3452,N_3422);
or U3706 (N_3706,N_3441,N_3434);
xor U3707 (N_3707,N_3443,N_3582);
or U3708 (N_3708,N_3437,N_3422);
nand U3709 (N_3709,N_3472,N_3556);
nand U3710 (N_3710,N_3555,N_3534);
nor U3711 (N_3711,N_3586,N_3427);
nor U3712 (N_3712,N_3583,N_3557);
and U3713 (N_3713,N_3507,N_3473);
and U3714 (N_3714,N_3585,N_3419);
nor U3715 (N_3715,N_3533,N_3474);
nor U3716 (N_3716,N_3592,N_3457);
xor U3717 (N_3717,N_3500,N_3431);
or U3718 (N_3718,N_3504,N_3412);
nand U3719 (N_3719,N_3414,N_3461);
nand U3720 (N_3720,N_3586,N_3550);
or U3721 (N_3721,N_3444,N_3414);
or U3722 (N_3722,N_3532,N_3592);
xor U3723 (N_3723,N_3402,N_3599);
or U3724 (N_3724,N_3550,N_3496);
nand U3725 (N_3725,N_3590,N_3576);
xor U3726 (N_3726,N_3426,N_3424);
nor U3727 (N_3727,N_3591,N_3470);
nand U3728 (N_3728,N_3401,N_3571);
or U3729 (N_3729,N_3571,N_3539);
or U3730 (N_3730,N_3400,N_3476);
or U3731 (N_3731,N_3508,N_3559);
and U3732 (N_3732,N_3513,N_3485);
and U3733 (N_3733,N_3584,N_3558);
or U3734 (N_3734,N_3414,N_3496);
nor U3735 (N_3735,N_3579,N_3417);
nor U3736 (N_3736,N_3511,N_3435);
nand U3737 (N_3737,N_3430,N_3417);
and U3738 (N_3738,N_3536,N_3590);
xnor U3739 (N_3739,N_3426,N_3541);
or U3740 (N_3740,N_3434,N_3472);
and U3741 (N_3741,N_3467,N_3401);
nor U3742 (N_3742,N_3429,N_3473);
nand U3743 (N_3743,N_3521,N_3564);
nor U3744 (N_3744,N_3454,N_3440);
or U3745 (N_3745,N_3538,N_3489);
nor U3746 (N_3746,N_3490,N_3483);
and U3747 (N_3747,N_3450,N_3457);
xor U3748 (N_3748,N_3460,N_3442);
or U3749 (N_3749,N_3574,N_3588);
xor U3750 (N_3750,N_3596,N_3539);
xnor U3751 (N_3751,N_3413,N_3406);
and U3752 (N_3752,N_3540,N_3407);
or U3753 (N_3753,N_3410,N_3582);
nand U3754 (N_3754,N_3583,N_3564);
xnor U3755 (N_3755,N_3455,N_3411);
and U3756 (N_3756,N_3577,N_3534);
and U3757 (N_3757,N_3409,N_3486);
xnor U3758 (N_3758,N_3504,N_3482);
or U3759 (N_3759,N_3589,N_3482);
nand U3760 (N_3760,N_3466,N_3516);
and U3761 (N_3761,N_3446,N_3405);
or U3762 (N_3762,N_3443,N_3484);
nor U3763 (N_3763,N_3599,N_3499);
and U3764 (N_3764,N_3506,N_3427);
or U3765 (N_3765,N_3429,N_3579);
and U3766 (N_3766,N_3460,N_3553);
xor U3767 (N_3767,N_3512,N_3547);
nand U3768 (N_3768,N_3527,N_3528);
and U3769 (N_3769,N_3586,N_3509);
nand U3770 (N_3770,N_3536,N_3418);
nor U3771 (N_3771,N_3540,N_3510);
nand U3772 (N_3772,N_3463,N_3449);
nor U3773 (N_3773,N_3505,N_3412);
or U3774 (N_3774,N_3575,N_3428);
or U3775 (N_3775,N_3422,N_3407);
and U3776 (N_3776,N_3475,N_3563);
or U3777 (N_3777,N_3538,N_3569);
nand U3778 (N_3778,N_3484,N_3429);
and U3779 (N_3779,N_3402,N_3519);
nand U3780 (N_3780,N_3417,N_3537);
nor U3781 (N_3781,N_3512,N_3595);
xnor U3782 (N_3782,N_3484,N_3454);
nor U3783 (N_3783,N_3509,N_3584);
nand U3784 (N_3784,N_3543,N_3405);
nor U3785 (N_3785,N_3472,N_3519);
xor U3786 (N_3786,N_3515,N_3519);
xor U3787 (N_3787,N_3568,N_3558);
nand U3788 (N_3788,N_3402,N_3410);
nor U3789 (N_3789,N_3442,N_3422);
and U3790 (N_3790,N_3588,N_3411);
nand U3791 (N_3791,N_3451,N_3472);
nor U3792 (N_3792,N_3522,N_3553);
nor U3793 (N_3793,N_3413,N_3508);
and U3794 (N_3794,N_3585,N_3495);
or U3795 (N_3795,N_3411,N_3454);
nor U3796 (N_3796,N_3490,N_3539);
nand U3797 (N_3797,N_3422,N_3469);
nand U3798 (N_3798,N_3486,N_3561);
and U3799 (N_3799,N_3435,N_3408);
or U3800 (N_3800,N_3752,N_3745);
and U3801 (N_3801,N_3685,N_3781);
nor U3802 (N_3802,N_3762,N_3607);
or U3803 (N_3803,N_3628,N_3718);
or U3804 (N_3804,N_3796,N_3707);
nor U3805 (N_3805,N_3701,N_3784);
nor U3806 (N_3806,N_3642,N_3743);
nor U3807 (N_3807,N_3790,N_3658);
xor U3808 (N_3808,N_3690,N_3791);
xnor U3809 (N_3809,N_3744,N_3664);
or U3810 (N_3810,N_3732,N_3671);
and U3811 (N_3811,N_3770,N_3632);
nand U3812 (N_3812,N_3742,N_3644);
and U3813 (N_3813,N_3794,N_3719);
or U3814 (N_3814,N_3786,N_3666);
and U3815 (N_3815,N_3720,N_3747);
or U3816 (N_3816,N_3624,N_3733);
or U3817 (N_3817,N_3736,N_3767);
xnor U3818 (N_3818,N_3660,N_3697);
nand U3819 (N_3819,N_3604,N_3649);
xnor U3820 (N_3820,N_3731,N_3764);
nand U3821 (N_3821,N_3645,N_3708);
nand U3822 (N_3822,N_3651,N_3616);
and U3823 (N_3823,N_3689,N_3799);
nand U3824 (N_3824,N_3655,N_3798);
nor U3825 (N_3825,N_3759,N_3676);
xor U3826 (N_3826,N_3713,N_3748);
nor U3827 (N_3827,N_3627,N_3758);
nor U3828 (N_3828,N_3686,N_3797);
nand U3829 (N_3829,N_3674,N_3605);
nor U3830 (N_3830,N_3638,N_3612);
xor U3831 (N_3831,N_3600,N_3668);
or U3832 (N_3832,N_3782,N_3654);
xnor U3833 (N_3833,N_3618,N_3679);
xor U3834 (N_3834,N_3661,N_3741);
or U3835 (N_3835,N_3740,N_3785);
and U3836 (N_3836,N_3634,N_3656);
or U3837 (N_3837,N_3776,N_3688);
and U3838 (N_3838,N_3646,N_3780);
nand U3839 (N_3839,N_3637,N_3702);
xnor U3840 (N_3840,N_3768,N_3691);
xor U3841 (N_3841,N_3619,N_3611);
and U3842 (N_3842,N_3777,N_3705);
nand U3843 (N_3843,N_3728,N_3709);
nand U3844 (N_3844,N_3641,N_3749);
and U3845 (N_3845,N_3723,N_3783);
nand U3846 (N_3846,N_3615,N_3631);
and U3847 (N_3847,N_3695,N_3734);
nor U3848 (N_3848,N_3602,N_3775);
and U3849 (N_3849,N_3699,N_3703);
nand U3850 (N_3850,N_3670,N_3769);
or U3851 (N_3851,N_3684,N_3773);
or U3852 (N_3852,N_3787,N_3636);
or U3853 (N_3853,N_3650,N_3601);
and U3854 (N_3854,N_3696,N_3724);
and U3855 (N_3855,N_3669,N_3738);
or U3856 (N_3856,N_3635,N_3725);
xor U3857 (N_3857,N_3606,N_3761);
and U3858 (N_3858,N_3662,N_3771);
or U3859 (N_3859,N_3754,N_3663);
xnor U3860 (N_3860,N_3756,N_3737);
xnor U3861 (N_3861,N_3665,N_3680);
xnor U3862 (N_3862,N_3630,N_3779);
nor U3863 (N_3863,N_3652,N_3735);
xnor U3864 (N_3864,N_3608,N_3710);
and U3865 (N_3865,N_3755,N_3712);
nand U3866 (N_3866,N_3792,N_3639);
and U3867 (N_3867,N_3778,N_3698);
xor U3868 (N_3868,N_3717,N_3677);
xor U3869 (N_3869,N_3706,N_3727);
nor U3870 (N_3870,N_3711,N_3739);
or U3871 (N_3871,N_3774,N_3772);
nor U3872 (N_3872,N_3620,N_3647);
xor U3873 (N_3873,N_3683,N_3673);
or U3874 (N_3874,N_3704,N_3757);
nand U3875 (N_3875,N_3760,N_3687);
xor U3876 (N_3876,N_3753,N_3726);
or U3877 (N_3877,N_3626,N_3623);
and U3878 (N_3878,N_3682,N_3617);
and U3879 (N_3879,N_3681,N_3672);
or U3880 (N_3880,N_3657,N_3692);
and U3881 (N_3881,N_3621,N_3633);
nand U3882 (N_3882,N_3700,N_3795);
xnor U3883 (N_3883,N_3716,N_3648);
or U3884 (N_3884,N_3750,N_3653);
xor U3885 (N_3885,N_3721,N_3722);
xor U3886 (N_3886,N_3614,N_3765);
nand U3887 (N_3887,N_3659,N_3694);
xor U3888 (N_3888,N_3751,N_3693);
or U3889 (N_3889,N_3609,N_3629);
and U3890 (N_3890,N_3667,N_3714);
nor U3891 (N_3891,N_3613,N_3730);
nand U3892 (N_3892,N_3603,N_3675);
nor U3893 (N_3893,N_3788,N_3715);
nor U3894 (N_3894,N_3622,N_3746);
nand U3895 (N_3895,N_3610,N_3789);
and U3896 (N_3896,N_3763,N_3678);
nand U3897 (N_3897,N_3643,N_3729);
nand U3898 (N_3898,N_3640,N_3793);
nor U3899 (N_3899,N_3625,N_3766);
nor U3900 (N_3900,N_3626,N_3693);
nor U3901 (N_3901,N_3675,N_3661);
xnor U3902 (N_3902,N_3629,N_3616);
nand U3903 (N_3903,N_3695,N_3610);
nor U3904 (N_3904,N_3630,N_3600);
or U3905 (N_3905,N_3669,N_3758);
nand U3906 (N_3906,N_3632,N_3640);
or U3907 (N_3907,N_3682,N_3692);
and U3908 (N_3908,N_3715,N_3739);
and U3909 (N_3909,N_3772,N_3702);
and U3910 (N_3910,N_3600,N_3695);
and U3911 (N_3911,N_3761,N_3756);
nor U3912 (N_3912,N_3711,N_3791);
nand U3913 (N_3913,N_3652,N_3635);
or U3914 (N_3914,N_3795,N_3642);
xor U3915 (N_3915,N_3798,N_3693);
nor U3916 (N_3916,N_3712,N_3781);
nand U3917 (N_3917,N_3710,N_3622);
xnor U3918 (N_3918,N_3639,N_3669);
or U3919 (N_3919,N_3757,N_3701);
xnor U3920 (N_3920,N_3753,N_3671);
or U3921 (N_3921,N_3662,N_3784);
nor U3922 (N_3922,N_3618,N_3691);
nand U3923 (N_3923,N_3757,N_3710);
nand U3924 (N_3924,N_3710,N_3787);
or U3925 (N_3925,N_3782,N_3645);
or U3926 (N_3926,N_3614,N_3756);
and U3927 (N_3927,N_3721,N_3760);
nand U3928 (N_3928,N_3791,N_3706);
nor U3929 (N_3929,N_3783,N_3754);
or U3930 (N_3930,N_3768,N_3769);
xor U3931 (N_3931,N_3754,N_3600);
and U3932 (N_3932,N_3621,N_3793);
or U3933 (N_3933,N_3762,N_3777);
and U3934 (N_3934,N_3626,N_3660);
nor U3935 (N_3935,N_3755,N_3717);
and U3936 (N_3936,N_3654,N_3761);
nor U3937 (N_3937,N_3618,N_3667);
or U3938 (N_3938,N_3633,N_3650);
nand U3939 (N_3939,N_3601,N_3638);
and U3940 (N_3940,N_3657,N_3682);
and U3941 (N_3941,N_3654,N_3789);
xor U3942 (N_3942,N_3684,N_3711);
nor U3943 (N_3943,N_3602,N_3696);
nand U3944 (N_3944,N_3703,N_3692);
nor U3945 (N_3945,N_3625,N_3624);
nand U3946 (N_3946,N_3712,N_3738);
and U3947 (N_3947,N_3757,N_3792);
xor U3948 (N_3948,N_3767,N_3772);
xor U3949 (N_3949,N_3727,N_3622);
and U3950 (N_3950,N_3683,N_3687);
and U3951 (N_3951,N_3627,N_3792);
or U3952 (N_3952,N_3748,N_3722);
nand U3953 (N_3953,N_3704,N_3721);
nor U3954 (N_3954,N_3657,N_3752);
xor U3955 (N_3955,N_3775,N_3736);
nor U3956 (N_3956,N_3732,N_3758);
and U3957 (N_3957,N_3682,N_3679);
nand U3958 (N_3958,N_3604,N_3720);
nand U3959 (N_3959,N_3771,N_3785);
nor U3960 (N_3960,N_3610,N_3767);
nor U3961 (N_3961,N_3786,N_3729);
nor U3962 (N_3962,N_3685,N_3604);
and U3963 (N_3963,N_3713,N_3680);
nand U3964 (N_3964,N_3678,N_3655);
nor U3965 (N_3965,N_3756,N_3637);
and U3966 (N_3966,N_3693,N_3642);
or U3967 (N_3967,N_3691,N_3755);
and U3968 (N_3968,N_3758,N_3794);
or U3969 (N_3969,N_3766,N_3684);
and U3970 (N_3970,N_3708,N_3631);
nor U3971 (N_3971,N_3717,N_3728);
and U3972 (N_3972,N_3602,N_3620);
nor U3973 (N_3973,N_3695,N_3669);
nand U3974 (N_3974,N_3644,N_3705);
and U3975 (N_3975,N_3771,N_3651);
nor U3976 (N_3976,N_3711,N_3700);
or U3977 (N_3977,N_3661,N_3654);
xnor U3978 (N_3978,N_3699,N_3740);
nand U3979 (N_3979,N_3739,N_3735);
nor U3980 (N_3980,N_3685,N_3646);
nor U3981 (N_3981,N_3777,N_3634);
or U3982 (N_3982,N_3767,N_3674);
nor U3983 (N_3983,N_3797,N_3629);
xnor U3984 (N_3984,N_3701,N_3746);
xor U3985 (N_3985,N_3601,N_3666);
and U3986 (N_3986,N_3622,N_3655);
nand U3987 (N_3987,N_3667,N_3699);
nand U3988 (N_3988,N_3715,N_3642);
and U3989 (N_3989,N_3632,N_3627);
nand U3990 (N_3990,N_3669,N_3716);
or U3991 (N_3991,N_3651,N_3733);
or U3992 (N_3992,N_3638,N_3740);
nand U3993 (N_3993,N_3644,N_3753);
or U3994 (N_3994,N_3752,N_3730);
or U3995 (N_3995,N_3673,N_3763);
and U3996 (N_3996,N_3630,N_3719);
and U3997 (N_3997,N_3690,N_3655);
or U3998 (N_3998,N_3719,N_3620);
xnor U3999 (N_3999,N_3654,N_3713);
nand U4000 (N_4000,N_3837,N_3830);
xor U4001 (N_4001,N_3850,N_3977);
nor U4002 (N_4002,N_3891,N_3807);
xor U4003 (N_4003,N_3862,N_3923);
and U4004 (N_4004,N_3967,N_3946);
or U4005 (N_4005,N_3903,N_3829);
nor U4006 (N_4006,N_3984,N_3904);
or U4007 (N_4007,N_3831,N_3918);
nand U4008 (N_4008,N_3908,N_3812);
or U4009 (N_4009,N_3851,N_3893);
xor U4010 (N_4010,N_3979,N_3939);
and U4011 (N_4011,N_3847,N_3856);
or U4012 (N_4012,N_3951,N_3991);
nand U4013 (N_4013,N_3915,N_3959);
xnor U4014 (N_4014,N_3810,N_3818);
and U4015 (N_4015,N_3888,N_3973);
and U4016 (N_4016,N_3974,N_3952);
xor U4017 (N_4017,N_3824,N_3986);
nor U4018 (N_4018,N_3826,N_3828);
nor U4019 (N_4019,N_3931,N_3942);
nand U4020 (N_4020,N_3976,N_3928);
or U4021 (N_4021,N_3917,N_3901);
and U4022 (N_4022,N_3880,N_3896);
nand U4023 (N_4023,N_3811,N_3982);
and U4024 (N_4024,N_3874,N_3940);
nand U4025 (N_4025,N_3846,N_3802);
nor U4026 (N_4026,N_3912,N_3869);
or U4027 (N_4027,N_3889,N_3963);
xnor U4028 (N_4028,N_3859,N_3965);
nand U4029 (N_4029,N_3884,N_3838);
nand U4030 (N_4030,N_3932,N_3962);
xor U4031 (N_4031,N_3845,N_3873);
nor U4032 (N_4032,N_3895,N_3985);
or U4033 (N_4033,N_3841,N_3815);
or U4034 (N_4034,N_3855,N_3953);
nor U4035 (N_4035,N_3950,N_3806);
or U4036 (N_4036,N_3836,N_3966);
xnor U4037 (N_4037,N_3968,N_3906);
xor U4038 (N_4038,N_3927,N_3972);
nand U4039 (N_4039,N_3910,N_3899);
nand U4040 (N_4040,N_3930,N_3929);
and U4041 (N_4041,N_3821,N_3844);
nor U4042 (N_4042,N_3877,N_3848);
and U4043 (N_4043,N_3994,N_3937);
xnor U4044 (N_4044,N_3870,N_3887);
nor U4045 (N_4045,N_3957,N_3805);
and U4046 (N_4046,N_3925,N_3817);
nand U4047 (N_4047,N_3970,N_3922);
nand U4048 (N_4048,N_3867,N_3894);
xor U4049 (N_4049,N_3854,N_3866);
nor U4050 (N_4050,N_3840,N_3964);
nand U4051 (N_4051,N_3809,N_3800);
or U4052 (N_4052,N_3993,N_3881);
nand U4053 (N_4053,N_3849,N_3947);
xnor U4054 (N_4054,N_3938,N_3820);
or U4055 (N_4055,N_3843,N_3833);
nand U4056 (N_4056,N_3956,N_3936);
or U4057 (N_4057,N_3934,N_3960);
nand U4058 (N_4058,N_3961,N_3913);
or U4059 (N_4059,N_3943,N_3808);
and U4060 (N_4060,N_3892,N_3998);
nand U4061 (N_4061,N_3905,N_3827);
nor U4062 (N_4062,N_3865,N_3933);
nand U4063 (N_4063,N_3911,N_3803);
xor U4064 (N_4064,N_3819,N_3839);
nor U4065 (N_4065,N_3935,N_3944);
xor U4066 (N_4066,N_3955,N_3909);
or U4067 (N_4067,N_3919,N_3898);
nor U4068 (N_4068,N_3988,N_3969);
xor U4069 (N_4069,N_3864,N_3814);
or U4070 (N_4070,N_3878,N_3825);
or U4071 (N_4071,N_3978,N_3975);
nor U4072 (N_4072,N_3948,N_3990);
xor U4073 (N_4073,N_3857,N_3900);
or U4074 (N_4074,N_3907,N_3858);
nand U4075 (N_4075,N_3914,N_3983);
or U4076 (N_4076,N_3822,N_3834);
nor U4077 (N_4077,N_3842,N_3868);
nor U4078 (N_4078,N_3997,N_3989);
xor U4079 (N_4079,N_3996,N_3816);
or U4080 (N_4080,N_3872,N_3995);
and U4081 (N_4081,N_3971,N_3863);
and U4082 (N_4082,N_3945,N_3897);
nand U4083 (N_4083,N_3921,N_3835);
nor U4084 (N_4084,N_3871,N_3853);
and U4085 (N_4085,N_3981,N_3804);
and U4086 (N_4086,N_3916,N_3926);
or U4087 (N_4087,N_3980,N_3876);
xor U4088 (N_4088,N_3920,N_3883);
nor U4089 (N_4089,N_3861,N_3813);
and U4090 (N_4090,N_3958,N_3886);
xor U4091 (N_4091,N_3992,N_3902);
xor U4092 (N_4092,N_3832,N_3882);
or U4093 (N_4093,N_3924,N_3885);
nand U4094 (N_4094,N_3875,N_3954);
xor U4095 (N_4095,N_3823,N_3941);
or U4096 (N_4096,N_3801,N_3879);
nand U4097 (N_4097,N_3999,N_3949);
nand U4098 (N_4098,N_3987,N_3860);
and U4099 (N_4099,N_3852,N_3890);
and U4100 (N_4100,N_3836,N_3887);
and U4101 (N_4101,N_3803,N_3909);
xnor U4102 (N_4102,N_3855,N_3826);
and U4103 (N_4103,N_3961,N_3846);
xor U4104 (N_4104,N_3955,N_3896);
xnor U4105 (N_4105,N_3807,N_3886);
or U4106 (N_4106,N_3976,N_3931);
and U4107 (N_4107,N_3919,N_3968);
xnor U4108 (N_4108,N_3834,N_3851);
nor U4109 (N_4109,N_3807,N_3943);
or U4110 (N_4110,N_3910,N_3882);
nor U4111 (N_4111,N_3998,N_3966);
nor U4112 (N_4112,N_3855,N_3845);
and U4113 (N_4113,N_3944,N_3822);
xor U4114 (N_4114,N_3860,N_3936);
or U4115 (N_4115,N_3888,N_3901);
xor U4116 (N_4116,N_3925,N_3950);
nor U4117 (N_4117,N_3810,N_3847);
nand U4118 (N_4118,N_3890,N_3888);
and U4119 (N_4119,N_3831,N_3883);
nor U4120 (N_4120,N_3873,N_3823);
xor U4121 (N_4121,N_3879,N_3800);
or U4122 (N_4122,N_3863,N_3889);
and U4123 (N_4123,N_3832,N_3871);
or U4124 (N_4124,N_3835,N_3977);
xnor U4125 (N_4125,N_3906,N_3904);
and U4126 (N_4126,N_3833,N_3886);
xor U4127 (N_4127,N_3847,N_3953);
xor U4128 (N_4128,N_3907,N_3863);
nor U4129 (N_4129,N_3950,N_3913);
xor U4130 (N_4130,N_3811,N_3963);
nor U4131 (N_4131,N_3808,N_3831);
and U4132 (N_4132,N_3996,N_3847);
xnor U4133 (N_4133,N_3932,N_3844);
xor U4134 (N_4134,N_3854,N_3983);
xor U4135 (N_4135,N_3891,N_3951);
or U4136 (N_4136,N_3842,N_3978);
nand U4137 (N_4137,N_3978,N_3812);
and U4138 (N_4138,N_3803,N_3838);
and U4139 (N_4139,N_3961,N_3929);
or U4140 (N_4140,N_3951,N_3867);
nand U4141 (N_4141,N_3891,N_3839);
nand U4142 (N_4142,N_3807,N_3870);
nand U4143 (N_4143,N_3968,N_3838);
nor U4144 (N_4144,N_3987,N_3844);
or U4145 (N_4145,N_3987,N_3806);
nor U4146 (N_4146,N_3934,N_3850);
or U4147 (N_4147,N_3854,N_3921);
or U4148 (N_4148,N_3906,N_3899);
xor U4149 (N_4149,N_3998,N_3987);
xnor U4150 (N_4150,N_3863,N_3990);
nand U4151 (N_4151,N_3875,N_3918);
nor U4152 (N_4152,N_3832,N_3897);
nor U4153 (N_4153,N_3907,N_3984);
or U4154 (N_4154,N_3917,N_3906);
xnor U4155 (N_4155,N_3935,N_3979);
nand U4156 (N_4156,N_3992,N_3904);
and U4157 (N_4157,N_3926,N_3864);
xnor U4158 (N_4158,N_3858,N_3929);
nor U4159 (N_4159,N_3918,N_3932);
xor U4160 (N_4160,N_3973,N_3852);
or U4161 (N_4161,N_3968,N_3939);
nor U4162 (N_4162,N_3813,N_3849);
nor U4163 (N_4163,N_3899,N_3870);
nor U4164 (N_4164,N_3883,N_3986);
and U4165 (N_4165,N_3862,N_3812);
xor U4166 (N_4166,N_3800,N_3911);
nor U4167 (N_4167,N_3857,N_3942);
or U4168 (N_4168,N_3981,N_3994);
or U4169 (N_4169,N_3938,N_3972);
nor U4170 (N_4170,N_3949,N_3878);
nor U4171 (N_4171,N_3976,N_3939);
nor U4172 (N_4172,N_3908,N_3871);
xor U4173 (N_4173,N_3999,N_3985);
or U4174 (N_4174,N_3999,N_3832);
nand U4175 (N_4175,N_3863,N_3862);
nand U4176 (N_4176,N_3947,N_3900);
nor U4177 (N_4177,N_3868,N_3962);
nor U4178 (N_4178,N_3819,N_3939);
nor U4179 (N_4179,N_3883,N_3919);
xor U4180 (N_4180,N_3921,N_3874);
and U4181 (N_4181,N_3864,N_3949);
xor U4182 (N_4182,N_3849,N_3942);
and U4183 (N_4183,N_3916,N_3801);
xnor U4184 (N_4184,N_3812,N_3824);
xnor U4185 (N_4185,N_3998,N_3822);
or U4186 (N_4186,N_3873,N_3809);
nor U4187 (N_4187,N_3859,N_3889);
xnor U4188 (N_4188,N_3894,N_3918);
and U4189 (N_4189,N_3829,N_3854);
and U4190 (N_4190,N_3898,N_3968);
or U4191 (N_4191,N_3971,N_3869);
or U4192 (N_4192,N_3960,N_3965);
xor U4193 (N_4193,N_3975,N_3850);
nor U4194 (N_4194,N_3947,N_3901);
nand U4195 (N_4195,N_3936,N_3933);
xnor U4196 (N_4196,N_3949,N_3819);
nor U4197 (N_4197,N_3948,N_3994);
nor U4198 (N_4198,N_3834,N_3867);
xor U4199 (N_4199,N_3950,N_3847);
and U4200 (N_4200,N_4026,N_4162);
nand U4201 (N_4201,N_4013,N_4030);
and U4202 (N_4202,N_4166,N_4146);
or U4203 (N_4203,N_4140,N_4045);
nor U4204 (N_4204,N_4059,N_4124);
nand U4205 (N_4205,N_4049,N_4056);
nor U4206 (N_4206,N_4084,N_4086);
nand U4207 (N_4207,N_4067,N_4085);
and U4208 (N_4208,N_4163,N_4088);
nand U4209 (N_4209,N_4091,N_4099);
xnor U4210 (N_4210,N_4193,N_4071);
and U4211 (N_4211,N_4157,N_4009);
and U4212 (N_4212,N_4178,N_4113);
and U4213 (N_4213,N_4001,N_4159);
nor U4214 (N_4214,N_4083,N_4130);
and U4215 (N_4215,N_4177,N_4106);
and U4216 (N_4216,N_4198,N_4016);
or U4217 (N_4217,N_4053,N_4047);
nand U4218 (N_4218,N_4002,N_4102);
and U4219 (N_4219,N_4080,N_4074);
or U4220 (N_4220,N_4090,N_4142);
xnor U4221 (N_4221,N_4191,N_4164);
xor U4222 (N_4222,N_4199,N_4019);
and U4223 (N_4223,N_4087,N_4182);
and U4224 (N_4224,N_4097,N_4003);
xor U4225 (N_4225,N_4109,N_4076);
nand U4226 (N_4226,N_4111,N_4044);
nand U4227 (N_4227,N_4025,N_4137);
nor U4228 (N_4228,N_4107,N_4195);
and U4229 (N_4229,N_4165,N_4141);
xor U4230 (N_4230,N_4148,N_4161);
or U4231 (N_4231,N_4125,N_4129);
nor U4232 (N_4232,N_4119,N_4062);
xor U4233 (N_4233,N_4179,N_4055);
and U4234 (N_4234,N_4024,N_4171);
or U4235 (N_4235,N_4063,N_4104);
nor U4236 (N_4236,N_4185,N_4188);
nand U4237 (N_4237,N_4022,N_4128);
xor U4238 (N_4238,N_4153,N_4154);
or U4239 (N_4239,N_4079,N_4040);
and U4240 (N_4240,N_4108,N_4028);
nor U4241 (N_4241,N_4064,N_4114);
and U4242 (N_4242,N_4082,N_4068);
xnor U4243 (N_4243,N_4050,N_4038);
and U4244 (N_4244,N_4190,N_4187);
nand U4245 (N_4245,N_4121,N_4158);
or U4246 (N_4246,N_4155,N_4115);
nor U4247 (N_4247,N_4034,N_4020);
xnor U4248 (N_4248,N_4035,N_4173);
or U4249 (N_4249,N_4183,N_4105);
nor U4250 (N_4250,N_4112,N_4041);
nand U4251 (N_4251,N_4000,N_4012);
nand U4252 (N_4252,N_4094,N_4120);
nand U4253 (N_4253,N_4150,N_4132);
or U4254 (N_4254,N_4169,N_4031);
nor U4255 (N_4255,N_4118,N_4135);
and U4256 (N_4256,N_4052,N_4189);
xnor U4257 (N_4257,N_4123,N_4110);
nor U4258 (N_4258,N_4138,N_4077);
or U4259 (N_4259,N_4096,N_4008);
or U4260 (N_4260,N_4027,N_4039);
nand U4261 (N_4261,N_4054,N_4015);
or U4262 (N_4262,N_4194,N_4131);
nor U4263 (N_4263,N_4078,N_4073);
nor U4264 (N_4264,N_4037,N_4010);
and U4265 (N_4265,N_4101,N_4042);
nand U4266 (N_4266,N_4032,N_4048);
xnor U4267 (N_4267,N_4151,N_4176);
or U4268 (N_4268,N_4100,N_4147);
nor U4269 (N_4269,N_4060,N_4181);
or U4270 (N_4270,N_4023,N_4018);
nor U4271 (N_4271,N_4057,N_4103);
nor U4272 (N_4272,N_4180,N_4144);
and U4273 (N_4273,N_4069,N_4136);
nand U4274 (N_4274,N_4098,N_4081);
or U4275 (N_4275,N_4046,N_4092);
and U4276 (N_4276,N_4072,N_4116);
nor U4277 (N_4277,N_4036,N_4058);
xor U4278 (N_4278,N_4061,N_4006);
nor U4279 (N_4279,N_4065,N_4051);
and U4280 (N_4280,N_4184,N_4174);
nand U4281 (N_4281,N_4029,N_4122);
and U4282 (N_4282,N_4133,N_4021);
nor U4283 (N_4283,N_4167,N_4089);
or U4284 (N_4284,N_4117,N_4134);
and U4285 (N_4285,N_4156,N_4011);
nor U4286 (N_4286,N_4043,N_4093);
xnor U4287 (N_4287,N_4175,N_4160);
xnor U4288 (N_4288,N_4170,N_4186);
and U4289 (N_4289,N_4149,N_4152);
and U4290 (N_4290,N_4172,N_4143);
and U4291 (N_4291,N_4007,N_4066);
or U4292 (N_4292,N_4075,N_4139);
nand U4293 (N_4293,N_4145,N_4004);
or U4294 (N_4294,N_4005,N_4197);
xnor U4295 (N_4295,N_4127,N_4126);
or U4296 (N_4296,N_4017,N_4033);
xnor U4297 (N_4297,N_4095,N_4168);
nand U4298 (N_4298,N_4192,N_4196);
nand U4299 (N_4299,N_4070,N_4014);
and U4300 (N_4300,N_4116,N_4141);
xor U4301 (N_4301,N_4008,N_4045);
or U4302 (N_4302,N_4173,N_4081);
nand U4303 (N_4303,N_4133,N_4037);
or U4304 (N_4304,N_4167,N_4170);
nand U4305 (N_4305,N_4156,N_4109);
and U4306 (N_4306,N_4089,N_4151);
nor U4307 (N_4307,N_4077,N_4169);
or U4308 (N_4308,N_4024,N_4033);
xnor U4309 (N_4309,N_4000,N_4062);
nor U4310 (N_4310,N_4187,N_4095);
xor U4311 (N_4311,N_4088,N_4098);
nor U4312 (N_4312,N_4161,N_4056);
and U4313 (N_4313,N_4139,N_4073);
xor U4314 (N_4314,N_4080,N_4114);
nor U4315 (N_4315,N_4085,N_4082);
nand U4316 (N_4316,N_4067,N_4108);
nor U4317 (N_4317,N_4034,N_4107);
and U4318 (N_4318,N_4178,N_4156);
and U4319 (N_4319,N_4069,N_4082);
nor U4320 (N_4320,N_4058,N_4080);
and U4321 (N_4321,N_4030,N_4127);
or U4322 (N_4322,N_4185,N_4148);
and U4323 (N_4323,N_4016,N_4194);
xnor U4324 (N_4324,N_4005,N_4185);
and U4325 (N_4325,N_4157,N_4197);
and U4326 (N_4326,N_4142,N_4064);
nor U4327 (N_4327,N_4078,N_4092);
nand U4328 (N_4328,N_4109,N_4106);
nand U4329 (N_4329,N_4095,N_4073);
nor U4330 (N_4330,N_4180,N_4028);
xnor U4331 (N_4331,N_4155,N_4102);
or U4332 (N_4332,N_4138,N_4086);
nor U4333 (N_4333,N_4151,N_4137);
and U4334 (N_4334,N_4113,N_4184);
and U4335 (N_4335,N_4143,N_4122);
and U4336 (N_4336,N_4098,N_4030);
nor U4337 (N_4337,N_4051,N_4011);
xor U4338 (N_4338,N_4118,N_4025);
and U4339 (N_4339,N_4127,N_4133);
nor U4340 (N_4340,N_4168,N_4146);
nand U4341 (N_4341,N_4083,N_4154);
or U4342 (N_4342,N_4146,N_4177);
nor U4343 (N_4343,N_4109,N_4175);
and U4344 (N_4344,N_4067,N_4154);
nand U4345 (N_4345,N_4159,N_4151);
and U4346 (N_4346,N_4069,N_4146);
and U4347 (N_4347,N_4048,N_4198);
xor U4348 (N_4348,N_4090,N_4165);
and U4349 (N_4349,N_4147,N_4040);
nor U4350 (N_4350,N_4196,N_4175);
or U4351 (N_4351,N_4070,N_4003);
or U4352 (N_4352,N_4115,N_4007);
and U4353 (N_4353,N_4164,N_4111);
xor U4354 (N_4354,N_4032,N_4034);
xor U4355 (N_4355,N_4040,N_4016);
nand U4356 (N_4356,N_4017,N_4123);
and U4357 (N_4357,N_4167,N_4100);
nand U4358 (N_4358,N_4105,N_4052);
or U4359 (N_4359,N_4074,N_4064);
or U4360 (N_4360,N_4033,N_4094);
xor U4361 (N_4361,N_4008,N_4198);
and U4362 (N_4362,N_4116,N_4019);
and U4363 (N_4363,N_4129,N_4016);
nand U4364 (N_4364,N_4121,N_4198);
xnor U4365 (N_4365,N_4056,N_4140);
nor U4366 (N_4366,N_4006,N_4065);
nand U4367 (N_4367,N_4036,N_4073);
or U4368 (N_4368,N_4008,N_4169);
nor U4369 (N_4369,N_4019,N_4132);
xor U4370 (N_4370,N_4105,N_4040);
xnor U4371 (N_4371,N_4107,N_4023);
or U4372 (N_4372,N_4091,N_4176);
xor U4373 (N_4373,N_4018,N_4102);
xor U4374 (N_4374,N_4133,N_4001);
nor U4375 (N_4375,N_4095,N_4107);
or U4376 (N_4376,N_4031,N_4186);
nand U4377 (N_4377,N_4146,N_4068);
nor U4378 (N_4378,N_4067,N_4134);
nor U4379 (N_4379,N_4172,N_4036);
xnor U4380 (N_4380,N_4153,N_4052);
or U4381 (N_4381,N_4126,N_4118);
and U4382 (N_4382,N_4032,N_4060);
nor U4383 (N_4383,N_4115,N_4100);
xor U4384 (N_4384,N_4051,N_4028);
xnor U4385 (N_4385,N_4123,N_4140);
or U4386 (N_4386,N_4140,N_4034);
and U4387 (N_4387,N_4063,N_4012);
xnor U4388 (N_4388,N_4140,N_4120);
and U4389 (N_4389,N_4037,N_4120);
xnor U4390 (N_4390,N_4186,N_4192);
or U4391 (N_4391,N_4166,N_4068);
and U4392 (N_4392,N_4061,N_4074);
nor U4393 (N_4393,N_4156,N_4135);
and U4394 (N_4394,N_4076,N_4053);
xor U4395 (N_4395,N_4058,N_4100);
nand U4396 (N_4396,N_4082,N_4105);
and U4397 (N_4397,N_4169,N_4027);
nand U4398 (N_4398,N_4165,N_4108);
or U4399 (N_4399,N_4023,N_4123);
xnor U4400 (N_4400,N_4252,N_4242);
xor U4401 (N_4401,N_4327,N_4292);
xor U4402 (N_4402,N_4270,N_4306);
and U4403 (N_4403,N_4365,N_4346);
nand U4404 (N_4404,N_4229,N_4384);
or U4405 (N_4405,N_4353,N_4288);
and U4406 (N_4406,N_4255,N_4393);
nand U4407 (N_4407,N_4345,N_4303);
nor U4408 (N_4408,N_4247,N_4271);
and U4409 (N_4409,N_4230,N_4222);
nor U4410 (N_4410,N_4387,N_4326);
nor U4411 (N_4411,N_4265,N_4262);
and U4412 (N_4412,N_4315,N_4269);
nor U4413 (N_4413,N_4227,N_4274);
nor U4414 (N_4414,N_4377,N_4366);
and U4415 (N_4415,N_4337,N_4237);
or U4416 (N_4416,N_4398,N_4300);
nand U4417 (N_4417,N_4301,N_4395);
nor U4418 (N_4418,N_4381,N_4243);
nand U4419 (N_4419,N_4212,N_4201);
and U4420 (N_4420,N_4207,N_4342);
or U4421 (N_4421,N_4200,N_4344);
nand U4422 (N_4422,N_4235,N_4329);
and U4423 (N_4423,N_4287,N_4215);
and U4424 (N_4424,N_4364,N_4399);
or U4425 (N_4425,N_4386,N_4253);
nand U4426 (N_4426,N_4378,N_4347);
nor U4427 (N_4427,N_4354,N_4338);
xnor U4428 (N_4428,N_4296,N_4249);
xnor U4429 (N_4429,N_4361,N_4362);
and U4430 (N_4430,N_4258,N_4310);
nand U4431 (N_4431,N_4285,N_4330);
nor U4432 (N_4432,N_4341,N_4375);
nor U4433 (N_4433,N_4283,N_4376);
or U4434 (N_4434,N_4221,N_4232);
nand U4435 (N_4435,N_4323,N_4313);
or U4436 (N_4436,N_4311,N_4290);
nor U4437 (N_4437,N_4322,N_4246);
xor U4438 (N_4438,N_4360,N_4309);
or U4439 (N_4439,N_4234,N_4307);
or U4440 (N_4440,N_4273,N_4276);
nand U4441 (N_4441,N_4336,N_4349);
xnor U4442 (N_4442,N_4213,N_4348);
nor U4443 (N_4443,N_4328,N_4363);
nand U4444 (N_4444,N_4299,N_4209);
xor U4445 (N_4445,N_4204,N_4340);
nand U4446 (N_4446,N_4351,N_4205);
nand U4447 (N_4447,N_4314,N_4263);
xor U4448 (N_4448,N_4220,N_4216);
and U4449 (N_4449,N_4282,N_4324);
nand U4450 (N_4450,N_4266,N_4251);
or U4451 (N_4451,N_4352,N_4367);
or U4452 (N_4452,N_4390,N_4278);
nor U4453 (N_4453,N_4259,N_4397);
nand U4454 (N_4454,N_4225,N_4239);
nor U4455 (N_4455,N_4359,N_4391);
and U4456 (N_4456,N_4343,N_4202);
xor U4457 (N_4457,N_4223,N_4389);
or U4458 (N_4458,N_4280,N_4248);
nand U4459 (N_4459,N_4332,N_4350);
nand U4460 (N_4460,N_4368,N_4286);
xor U4461 (N_4461,N_4335,N_4302);
xnor U4462 (N_4462,N_4379,N_4394);
or U4463 (N_4463,N_4305,N_4241);
xnor U4464 (N_4464,N_4317,N_4228);
xor U4465 (N_4465,N_4250,N_4275);
xnor U4466 (N_4466,N_4264,N_4268);
nor U4467 (N_4467,N_4226,N_4325);
nor U4468 (N_4468,N_4383,N_4293);
nand U4469 (N_4469,N_4331,N_4320);
nor U4470 (N_4470,N_4257,N_4304);
nand U4471 (N_4471,N_4333,N_4357);
nor U4472 (N_4472,N_4334,N_4203);
or U4473 (N_4473,N_4272,N_4318);
or U4474 (N_4474,N_4217,N_4289);
xor U4475 (N_4475,N_4214,N_4339);
xnor U4476 (N_4476,N_4369,N_4267);
and U4477 (N_4477,N_4294,N_4260);
nand U4478 (N_4478,N_4308,N_4210);
and U4479 (N_4479,N_4240,N_4231);
or U4480 (N_4480,N_4256,N_4233);
and U4481 (N_4481,N_4355,N_4372);
and U4482 (N_4482,N_4291,N_4380);
and U4483 (N_4483,N_4356,N_4245);
and U4484 (N_4484,N_4316,N_4319);
and U4485 (N_4485,N_4277,N_4396);
nand U4486 (N_4486,N_4211,N_4358);
or U4487 (N_4487,N_4218,N_4238);
xnor U4488 (N_4488,N_4281,N_4295);
nand U4489 (N_4489,N_4321,N_4206);
or U4490 (N_4490,N_4388,N_4297);
and U4491 (N_4491,N_4236,N_4219);
nor U4492 (N_4492,N_4370,N_4244);
and U4493 (N_4493,N_4279,N_4385);
and U4494 (N_4494,N_4254,N_4312);
or U4495 (N_4495,N_4373,N_4208);
or U4496 (N_4496,N_4224,N_4374);
or U4497 (N_4497,N_4261,N_4371);
nand U4498 (N_4498,N_4298,N_4392);
nand U4499 (N_4499,N_4284,N_4382);
nor U4500 (N_4500,N_4213,N_4288);
xnor U4501 (N_4501,N_4238,N_4393);
nand U4502 (N_4502,N_4228,N_4202);
nand U4503 (N_4503,N_4389,N_4244);
nand U4504 (N_4504,N_4367,N_4242);
and U4505 (N_4505,N_4228,N_4343);
and U4506 (N_4506,N_4329,N_4242);
and U4507 (N_4507,N_4319,N_4379);
nand U4508 (N_4508,N_4221,N_4310);
nand U4509 (N_4509,N_4312,N_4245);
nand U4510 (N_4510,N_4229,N_4246);
or U4511 (N_4511,N_4343,N_4252);
nand U4512 (N_4512,N_4391,N_4296);
nor U4513 (N_4513,N_4255,N_4322);
nand U4514 (N_4514,N_4261,N_4367);
and U4515 (N_4515,N_4362,N_4352);
or U4516 (N_4516,N_4260,N_4399);
xnor U4517 (N_4517,N_4344,N_4374);
nand U4518 (N_4518,N_4336,N_4335);
nand U4519 (N_4519,N_4387,N_4262);
or U4520 (N_4520,N_4333,N_4380);
nor U4521 (N_4521,N_4312,N_4205);
and U4522 (N_4522,N_4288,N_4233);
nor U4523 (N_4523,N_4308,N_4243);
nand U4524 (N_4524,N_4283,N_4284);
nand U4525 (N_4525,N_4243,N_4280);
xnor U4526 (N_4526,N_4388,N_4254);
nor U4527 (N_4527,N_4266,N_4329);
nor U4528 (N_4528,N_4386,N_4246);
nor U4529 (N_4529,N_4207,N_4237);
or U4530 (N_4530,N_4215,N_4241);
nand U4531 (N_4531,N_4256,N_4246);
and U4532 (N_4532,N_4282,N_4302);
and U4533 (N_4533,N_4223,N_4368);
nor U4534 (N_4534,N_4237,N_4288);
xnor U4535 (N_4535,N_4336,N_4345);
nand U4536 (N_4536,N_4299,N_4320);
xor U4537 (N_4537,N_4268,N_4258);
xnor U4538 (N_4538,N_4266,N_4272);
or U4539 (N_4539,N_4268,N_4348);
and U4540 (N_4540,N_4263,N_4244);
or U4541 (N_4541,N_4354,N_4225);
or U4542 (N_4542,N_4244,N_4289);
nand U4543 (N_4543,N_4318,N_4324);
and U4544 (N_4544,N_4386,N_4224);
xnor U4545 (N_4545,N_4280,N_4348);
xnor U4546 (N_4546,N_4361,N_4300);
nand U4547 (N_4547,N_4349,N_4219);
nor U4548 (N_4548,N_4248,N_4295);
nor U4549 (N_4549,N_4342,N_4388);
xnor U4550 (N_4550,N_4393,N_4336);
or U4551 (N_4551,N_4396,N_4302);
or U4552 (N_4552,N_4300,N_4239);
nor U4553 (N_4553,N_4284,N_4285);
and U4554 (N_4554,N_4321,N_4292);
nor U4555 (N_4555,N_4354,N_4245);
nor U4556 (N_4556,N_4311,N_4253);
nor U4557 (N_4557,N_4377,N_4264);
or U4558 (N_4558,N_4321,N_4312);
or U4559 (N_4559,N_4371,N_4369);
nor U4560 (N_4560,N_4301,N_4370);
nor U4561 (N_4561,N_4275,N_4216);
xor U4562 (N_4562,N_4315,N_4314);
xor U4563 (N_4563,N_4319,N_4243);
and U4564 (N_4564,N_4282,N_4326);
and U4565 (N_4565,N_4340,N_4382);
or U4566 (N_4566,N_4276,N_4385);
or U4567 (N_4567,N_4201,N_4267);
xnor U4568 (N_4568,N_4286,N_4312);
or U4569 (N_4569,N_4281,N_4320);
xnor U4570 (N_4570,N_4343,N_4325);
nor U4571 (N_4571,N_4268,N_4251);
xnor U4572 (N_4572,N_4321,N_4210);
and U4573 (N_4573,N_4369,N_4341);
and U4574 (N_4574,N_4351,N_4303);
or U4575 (N_4575,N_4240,N_4270);
nand U4576 (N_4576,N_4326,N_4310);
xnor U4577 (N_4577,N_4345,N_4368);
nand U4578 (N_4578,N_4327,N_4236);
and U4579 (N_4579,N_4262,N_4291);
nor U4580 (N_4580,N_4282,N_4321);
xor U4581 (N_4581,N_4355,N_4200);
nor U4582 (N_4582,N_4274,N_4243);
and U4583 (N_4583,N_4298,N_4256);
or U4584 (N_4584,N_4201,N_4293);
nand U4585 (N_4585,N_4203,N_4288);
nor U4586 (N_4586,N_4334,N_4255);
and U4587 (N_4587,N_4246,N_4397);
nand U4588 (N_4588,N_4320,N_4340);
xor U4589 (N_4589,N_4327,N_4254);
xnor U4590 (N_4590,N_4288,N_4335);
nand U4591 (N_4591,N_4278,N_4223);
or U4592 (N_4592,N_4320,N_4297);
nor U4593 (N_4593,N_4391,N_4348);
and U4594 (N_4594,N_4218,N_4354);
xor U4595 (N_4595,N_4330,N_4392);
and U4596 (N_4596,N_4260,N_4365);
or U4597 (N_4597,N_4391,N_4336);
nand U4598 (N_4598,N_4295,N_4344);
or U4599 (N_4599,N_4201,N_4351);
xnor U4600 (N_4600,N_4444,N_4495);
xor U4601 (N_4601,N_4471,N_4429);
or U4602 (N_4602,N_4527,N_4590);
and U4603 (N_4603,N_4447,N_4455);
and U4604 (N_4604,N_4426,N_4583);
xor U4605 (N_4605,N_4541,N_4441);
xnor U4606 (N_4606,N_4529,N_4420);
and U4607 (N_4607,N_4468,N_4438);
xnor U4608 (N_4608,N_4538,N_4599);
and U4609 (N_4609,N_4596,N_4557);
nor U4610 (N_4610,N_4479,N_4450);
nor U4611 (N_4611,N_4485,N_4416);
or U4612 (N_4612,N_4500,N_4404);
or U4613 (N_4613,N_4452,N_4475);
and U4614 (N_4614,N_4586,N_4491);
and U4615 (N_4615,N_4524,N_4577);
nor U4616 (N_4616,N_4554,N_4511);
and U4617 (N_4617,N_4476,N_4510);
xor U4618 (N_4618,N_4509,N_4503);
nor U4619 (N_4619,N_4517,N_4477);
xnor U4620 (N_4620,N_4564,N_4448);
or U4621 (N_4621,N_4446,N_4546);
and U4622 (N_4622,N_4421,N_4490);
or U4623 (N_4623,N_4506,N_4542);
nor U4624 (N_4624,N_4443,N_4515);
or U4625 (N_4625,N_4432,N_4526);
nor U4626 (N_4626,N_4464,N_4502);
and U4627 (N_4627,N_4530,N_4562);
nor U4628 (N_4628,N_4427,N_4551);
nand U4629 (N_4629,N_4466,N_4439);
xnor U4630 (N_4630,N_4496,N_4410);
nor U4631 (N_4631,N_4574,N_4474);
xor U4632 (N_4632,N_4433,N_4540);
nand U4633 (N_4633,N_4547,N_4480);
nor U4634 (N_4634,N_4431,N_4560);
nand U4635 (N_4635,N_4498,N_4435);
nor U4636 (N_4636,N_4593,N_4584);
nand U4637 (N_4637,N_4481,N_4520);
or U4638 (N_4638,N_4425,N_4545);
xnor U4639 (N_4639,N_4499,N_4482);
nor U4640 (N_4640,N_4413,N_4430);
nand U4641 (N_4641,N_4436,N_4456);
and U4642 (N_4642,N_4550,N_4451);
xnor U4643 (N_4643,N_4488,N_4406);
nand U4644 (N_4644,N_4423,N_4531);
xor U4645 (N_4645,N_4587,N_4408);
nand U4646 (N_4646,N_4414,N_4484);
or U4647 (N_4647,N_4454,N_4516);
nand U4648 (N_4648,N_4411,N_4457);
nand U4649 (N_4649,N_4553,N_4445);
or U4650 (N_4650,N_4533,N_4566);
xor U4651 (N_4651,N_4569,N_4534);
or U4652 (N_4652,N_4505,N_4563);
nand U4653 (N_4653,N_4597,N_4513);
and U4654 (N_4654,N_4543,N_4573);
nor U4655 (N_4655,N_4483,N_4489);
or U4656 (N_4656,N_4501,N_4522);
nand U4657 (N_4657,N_4582,N_4519);
nand U4658 (N_4658,N_4440,N_4472);
and U4659 (N_4659,N_4552,N_4585);
nand U4660 (N_4660,N_4419,N_4535);
or U4661 (N_4661,N_4403,N_4588);
xnor U4662 (N_4662,N_4571,N_4561);
nand U4663 (N_4663,N_4402,N_4467);
xnor U4664 (N_4664,N_4514,N_4463);
or U4665 (N_4665,N_4437,N_4598);
xor U4666 (N_4666,N_4508,N_4473);
xor U4667 (N_4667,N_4459,N_4528);
nand U4668 (N_4668,N_4544,N_4417);
or U4669 (N_4669,N_4572,N_4493);
xor U4670 (N_4670,N_4422,N_4409);
xnor U4671 (N_4671,N_4537,N_4525);
nor U4672 (N_4672,N_4497,N_4556);
xor U4673 (N_4673,N_4532,N_4549);
and U4674 (N_4674,N_4494,N_4559);
or U4675 (N_4675,N_4412,N_4453);
nand U4676 (N_4676,N_4536,N_4589);
and U4677 (N_4677,N_4405,N_4580);
or U4678 (N_4678,N_4478,N_4575);
nand U4679 (N_4679,N_4492,N_4592);
xor U4680 (N_4680,N_4460,N_4548);
nor U4681 (N_4681,N_4578,N_4424);
and U4682 (N_4682,N_4565,N_4461);
and U4683 (N_4683,N_4401,N_4407);
or U4684 (N_4684,N_4487,N_4567);
nand U4685 (N_4685,N_4594,N_4591);
or U4686 (N_4686,N_4428,N_4400);
nor U4687 (N_4687,N_4449,N_4415);
nor U4688 (N_4688,N_4442,N_4558);
or U4689 (N_4689,N_4418,N_4568);
nand U4690 (N_4690,N_4470,N_4523);
xor U4691 (N_4691,N_4469,N_4486);
and U4692 (N_4692,N_4595,N_4581);
nor U4693 (N_4693,N_4570,N_4576);
or U4694 (N_4694,N_4521,N_4518);
nor U4695 (N_4695,N_4507,N_4465);
or U4696 (N_4696,N_4504,N_4555);
and U4697 (N_4697,N_4462,N_4539);
xor U4698 (N_4698,N_4512,N_4579);
nor U4699 (N_4699,N_4458,N_4434);
nand U4700 (N_4700,N_4419,N_4503);
nand U4701 (N_4701,N_4473,N_4450);
xnor U4702 (N_4702,N_4561,N_4429);
nand U4703 (N_4703,N_4464,N_4536);
xor U4704 (N_4704,N_4495,N_4485);
xor U4705 (N_4705,N_4554,N_4495);
xnor U4706 (N_4706,N_4451,N_4562);
nand U4707 (N_4707,N_4570,N_4444);
xor U4708 (N_4708,N_4419,N_4422);
nand U4709 (N_4709,N_4529,N_4547);
nor U4710 (N_4710,N_4461,N_4473);
nor U4711 (N_4711,N_4531,N_4413);
xor U4712 (N_4712,N_4435,N_4523);
nand U4713 (N_4713,N_4472,N_4585);
nor U4714 (N_4714,N_4485,N_4421);
nor U4715 (N_4715,N_4500,N_4597);
or U4716 (N_4716,N_4591,N_4552);
or U4717 (N_4717,N_4433,N_4483);
nor U4718 (N_4718,N_4562,N_4581);
and U4719 (N_4719,N_4445,N_4454);
and U4720 (N_4720,N_4474,N_4411);
and U4721 (N_4721,N_4552,N_4402);
nor U4722 (N_4722,N_4462,N_4488);
nand U4723 (N_4723,N_4544,N_4561);
nand U4724 (N_4724,N_4571,N_4519);
xnor U4725 (N_4725,N_4417,N_4559);
nor U4726 (N_4726,N_4472,N_4485);
or U4727 (N_4727,N_4581,N_4493);
nor U4728 (N_4728,N_4408,N_4416);
nand U4729 (N_4729,N_4467,N_4418);
nand U4730 (N_4730,N_4561,N_4423);
nor U4731 (N_4731,N_4468,N_4555);
nand U4732 (N_4732,N_4582,N_4554);
nand U4733 (N_4733,N_4407,N_4487);
nor U4734 (N_4734,N_4520,N_4560);
nor U4735 (N_4735,N_4585,N_4425);
or U4736 (N_4736,N_4501,N_4490);
nand U4737 (N_4737,N_4514,N_4566);
nand U4738 (N_4738,N_4594,N_4533);
nor U4739 (N_4739,N_4436,N_4513);
or U4740 (N_4740,N_4516,N_4571);
or U4741 (N_4741,N_4431,N_4442);
nor U4742 (N_4742,N_4599,N_4573);
and U4743 (N_4743,N_4515,N_4574);
nor U4744 (N_4744,N_4599,N_4539);
nand U4745 (N_4745,N_4511,N_4587);
nor U4746 (N_4746,N_4543,N_4439);
xor U4747 (N_4747,N_4462,N_4598);
and U4748 (N_4748,N_4540,N_4503);
xnor U4749 (N_4749,N_4432,N_4554);
nor U4750 (N_4750,N_4416,N_4450);
nand U4751 (N_4751,N_4476,N_4447);
xor U4752 (N_4752,N_4497,N_4544);
and U4753 (N_4753,N_4466,N_4566);
nand U4754 (N_4754,N_4492,N_4530);
xnor U4755 (N_4755,N_4424,N_4496);
xor U4756 (N_4756,N_4584,N_4566);
nor U4757 (N_4757,N_4422,N_4447);
nand U4758 (N_4758,N_4531,N_4453);
or U4759 (N_4759,N_4524,N_4454);
or U4760 (N_4760,N_4409,N_4483);
nand U4761 (N_4761,N_4556,N_4583);
and U4762 (N_4762,N_4535,N_4575);
nand U4763 (N_4763,N_4560,N_4511);
or U4764 (N_4764,N_4529,N_4469);
and U4765 (N_4765,N_4407,N_4463);
and U4766 (N_4766,N_4416,N_4480);
nor U4767 (N_4767,N_4552,N_4460);
and U4768 (N_4768,N_4520,N_4556);
and U4769 (N_4769,N_4443,N_4596);
nand U4770 (N_4770,N_4551,N_4487);
xor U4771 (N_4771,N_4592,N_4477);
and U4772 (N_4772,N_4486,N_4508);
xor U4773 (N_4773,N_4545,N_4577);
nand U4774 (N_4774,N_4591,N_4489);
nor U4775 (N_4775,N_4496,N_4494);
nand U4776 (N_4776,N_4514,N_4509);
nor U4777 (N_4777,N_4566,N_4554);
nand U4778 (N_4778,N_4475,N_4522);
nand U4779 (N_4779,N_4502,N_4435);
xnor U4780 (N_4780,N_4574,N_4432);
or U4781 (N_4781,N_4436,N_4551);
and U4782 (N_4782,N_4438,N_4537);
and U4783 (N_4783,N_4583,N_4466);
xor U4784 (N_4784,N_4456,N_4415);
nand U4785 (N_4785,N_4588,N_4425);
nor U4786 (N_4786,N_4490,N_4474);
or U4787 (N_4787,N_4534,N_4519);
or U4788 (N_4788,N_4546,N_4464);
and U4789 (N_4789,N_4595,N_4493);
nand U4790 (N_4790,N_4548,N_4578);
nor U4791 (N_4791,N_4597,N_4569);
and U4792 (N_4792,N_4485,N_4555);
nand U4793 (N_4793,N_4428,N_4536);
nor U4794 (N_4794,N_4492,N_4523);
nand U4795 (N_4795,N_4554,N_4507);
and U4796 (N_4796,N_4547,N_4599);
and U4797 (N_4797,N_4599,N_4421);
xor U4798 (N_4798,N_4554,N_4480);
nor U4799 (N_4799,N_4546,N_4431);
nor U4800 (N_4800,N_4675,N_4705);
and U4801 (N_4801,N_4682,N_4715);
nor U4802 (N_4802,N_4681,N_4701);
xnor U4803 (N_4803,N_4753,N_4757);
and U4804 (N_4804,N_4781,N_4629);
nand U4805 (N_4805,N_4607,N_4673);
nand U4806 (N_4806,N_4685,N_4646);
xor U4807 (N_4807,N_4643,N_4718);
nand U4808 (N_4808,N_4683,N_4779);
nor U4809 (N_4809,N_4774,N_4672);
and U4810 (N_4810,N_4628,N_4704);
nor U4811 (N_4811,N_4692,N_4766);
xnor U4812 (N_4812,N_4676,N_4623);
and U4813 (N_4813,N_4617,N_4644);
nand U4814 (N_4814,N_4703,N_4729);
nand U4815 (N_4815,N_4669,N_4730);
and U4816 (N_4816,N_4654,N_4785);
nor U4817 (N_4817,N_4773,N_4776);
nand U4818 (N_4818,N_4625,N_4737);
nor U4819 (N_4819,N_4631,N_4618);
nand U4820 (N_4820,N_4719,N_4640);
nor U4821 (N_4821,N_4615,N_4602);
nor U4822 (N_4822,N_4797,N_4613);
xnor U4823 (N_4823,N_4700,N_4714);
and U4824 (N_4824,N_4661,N_4759);
or U4825 (N_4825,N_4659,N_4688);
and U4826 (N_4826,N_4667,N_4777);
and U4827 (N_4827,N_4755,N_4722);
nand U4828 (N_4828,N_4798,N_4707);
nor U4829 (N_4829,N_4680,N_4696);
nand U4830 (N_4830,N_4735,N_4780);
and U4831 (N_4831,N_4632,N_4764);
or U4832 (N_4832,N_4698,N_4726);
or U4833 (N_4833,N_4699,N_4686);
or U4834 (N_4834,N_4662,N_4712);
nand U4835 (N_4835,N_4711,N_4634);
nand U4836 (N_4836,N_4650,N_4621);
nand U4837 (N_4837,N_4684,N_4741);
and U4838 (N_4838,N_4736,N_4734);
nand U4839 (N_4839,N_4750,N_4791);
nand U4840 (N_4840,N_4651,N_4649);
nand U4841 (N_4841,N_4771,N_4619);
xor U4842 (N_4842,N_4616,N_4656);
nand U4843 (N_4843,N_4784,N_4727);
xnor U4844 (N_4844,N_4724,N_4691);
xor U4845 (N_4845,N_4763,N_4609);
nor U4846 (N_4846,N_4765,N_4678);
nand U4847 (N_4847,N_4733,N_4670);
nor U4848 (N_4848,N_4600,N_4713);
or U4849 (N_4849,N_4679,N_4639);
or U4850 (N_4850,N_4740,N_4767);
xnor U4851 (N_4851,N_4738,N_4725);
or U4852 (N_4852,N_4645,N_4663);
and U4853 (N_4853,N_4744,N_4743);
nor U4854 (N_4854,N_4604,N_4709);
or U4855 (N_4855,N_4605,N_4633);
nand U4856 (N_4856,N_4723,N_4695);
or U4857 (N_4857,N_4608,N_4665);
and U4858 (N_4858,N_4636,N_4756);
nand U4859 (N_4859,N_4638,N_4769);
nand U4860 (N_4860,N_4664,N_4620);
or U4861 (N_4861,N_4627,N_4768);
and U4862 (N_4862,N_4706,N_4742);
nor U4863 (N_4863,N_4748,N_4793);
and U4864 (N_4864,N_4697,N_4622);
and U4865 (N_4865,N_4610,N_4787);
xnor U4866 (N_4866,N_4652,N_4749);
nand U4867 (N_4867,N_4642,N_4612);
xor U4868 (N_4868,N_4790,N_4648);
nor U4869 (N_4869,N_4796,N_4666);
xor U4870 (N_4870,N_4671,N_4746);
and U4871 (N_4871,N_4624,N_4660);
nand U4872 (N_4872,N_4694,N_4782);
and U4873 (N_4873,N_4788,N_4693);
or U4874 (N_4874,N_4606,N_4770);
or U4875 (N_4875,N_4603,N_4687);
nor U4876 (N_4876,N_4637,N_4601);
nand U4877 (N_4877,N_4658,N_4655);
nor U4878 (N_4878,N_4728,N_4747);
and U4879 (N_4879,N_4775,N_4794);
and U4880 (N_4880,N_4795,N_4635);
nand U4881 (N_4881,N_4674,N_4641);
nand U4882 (N_4882,N_4745,N_4630);
nand U4883 (N_4883,N_4614,N_4721);
xor U4884 (N_4884,N_4732,N_4611);
xor U4885 (N_4885,N_4689,N_4786);
xor U4886 (N_4886,N_4783,N_4720);
nor U4887 (N_4887,N_4772,N_4702);
nor U4888 (N_4888,N_4690,N_4677);
nand U4889 (N_4889,N_4799,N_4647);
nor U4890 (N_4890,N_4657,N_4760);
or U4891 (N_4891,N_4792,N_4778);
and U4892 (N_4892,N_4716,N_4731);
and U4893 (N_4893,N_4762,N_4708);
xnor U4894 (N_4894,N_4752,N_4653);
and U4895 (N_4895,N_4710,N_4789);
or U4896 (N_4896,N_4668,N_4626);
xor U4897 (N_4897,N_4758,N_4717);
xnor U4898 (N_4898,N_4751,N_4754);
or U4899 (N_4899,N_4739,N_4761);
nor U4900 (N_4900,N_4733,N_4660);
nand U4901 (N_4901,N_4768,N_4619);
or U4902 (N_4902,N_4621,N_4609);
or U4903 (N_4903,N_4752,N_4758);
and U4904 (N_4904,N_4798,N_4686);
or U4905 (N_4905,N_4726,N_4774);
nand U4906 (N_4906,N_4680,N_4753);
nand U4907 (N_4907,N_4704,N_4629);
nor U4908 (N_4908,N_4741,N_4614);
nand U4909 (N_4909,N_4673,N_4704);
nor U4910 (N_4910,N_4754,N_4774);
and U4911 (N_4911,N_4640,N_4602);
or U4912 (N_4912,N_4668,N_4716);
nor U4913 (N_4913,N_4692,N_4760);
nor U4914 (N_4914,N_4720,N_4688);
or U4915 (N_4915,N_4650,N_4791);
or U4916 (N_4916,N_4730,N_4792);
nand U4917 (N_4917,N_4758,N_4704);
nor U4918 (N_4918,N_4762,N_4612);
and U4919 (N_4919,N_4653,N_4641);
or U4920 (N_4920,N_4644,N_4735);
and U4921 (N_4921,N_4649,N_4731);
and U4922 (N_4922,N_4650,N_4677);
or U4923 (N_4923,N_4778,N_4739);
nor U4924 (N_4924,N_4784,N_4750);
nand U4925 (N_4925,N_4668,N_4706);
and U4926 (N_4926,N_4630,N_4703);
xor U4927 (N_4927,N_4719,N_4768);
and U4928 (N_4928,N_4796,N_4691);
nor U4929 (N_4929,N_4656,N_4632);
xor U4930 (N_4930,N_4655,N_4712);
xnor U4931 (N_4931,N_4756,N_4652);
and U4932 (N_4932,N_4794,N_4605);
or U4933 (N_4933,N_4781,N_4603);
xor U4934 (N_4934,N_4677,N_4630);
or U4935 (N_4935,N_4678,N_4607);
xnor U4936 (N_4936,N_4710,N_4627);
xnor U4937 (N_4937,N_4669,N_4664);
xnor U4938 (N_4938,N_4784,N_4693);
nand U4939 (N_4939,N_4648,N_4720);
or U4940 (N_4940,N_4703,N_4695);
xnor U4941 (N_4941,N_4713,N_4719);
nand U4942 (N_4942,N_4748,N_4602);
nor U4943 (N_4943,N_4648,N_4782);
and U4944 (N_4944,N_4749,N_4684);
xnor U4945 (N_4945,N_4685,N_4607);
or U4946 (N_4946,N_4720,N_4759);
nand U4947 (N_4947,N_4741,N_4775);
or U4948 (N_4948,N_4680,N_4668);
xnor U4949 (N_4949,N_4608,N_4726);
or U4950 (N_4950,N_4707,N_4672);
nand U4951 (N_4951,N_4776,N_4639);
and U4952 (N_4952,N_4760,N_4711);
nand U4953 (N_4953,N_4662,N_4645);
nor U4954 (N_4954,N_4781,N_4651);
or U4955 (N_4955,N_4618,N_4683);
nand U4956 (N_4956,N_4703,N_4757);
and U4957 (N_4957,N_4641,N_4720);
nor U4958 (N_4958,N_4626,N_4685);
and U4959 (N_4959,N_4639,N_4668);
nand U4960 (N_4960,N_4659,N_4760);
nor U4961 (N_4961,N_4616,N_4701);
nand U4962 (N_4962,N_4638,N_4728);
nand U4963 (N_4963,N_4700,N_4786);
nor U4964 (N_4964,N_4731,N_4626);
or U4965 (N_4965,N_4686,N_4702);
and U4966 (N_4966,N_4668,N_4743);
and U4967 (N_4967,N_4703,N_4799);
nand U4968 (N_4968,N_4635,N_4725);
or U4969 (N_4969,N_4612,N_4670);
xnor U4970 (N_4970,N_4635,N_4739);
or U4971 (N_4971,N_4747,N_4696);
and U4972 (N_4972,N_4727,N_4743);
and U4973 (N_4973,N_4779,N_4636);
or U4974 (N_4974,N_4638,N_4757);
nor U4975 (N_4975,N_4755,N_4733);
and U4976 (N_4976,N_4734,N_4691);
xnor U4977 (N_4977,N_4661,N_4603);
or U4978 (N_4978,N_4760,N_4707);
or U4979 (N_4979,N_4636,N_4607);
nand U4980 (N_4980,N_4682,N_4799);
and U4981 (N_4981,N_4757,N_4740);
and U4982 (N_4982,N_4753,N_4701);
nor U4983 (N_4983,N_4733,N_4673);
nor U4984 (N_4984,N_4640,N_4765);
xor U4985 (N_4985,N_4757,N_4736);
nor U4986 (N_4986,N_4788,N_4701);
nand U4987 (N_4987,N_4729,N_4787);
xnor U4988 (N_4988,N_4649,N_4686);
xnor U4989 (N_4989,N_4621,N_4688);
or U4990 (N_4990,N_4669,N_4722);
and U4991 (N_4991,N_4673,N_4611);
nor U4992 (N_4992,N_4742,N_4653);
and U4993 (N_4993,N_4796,N_4633);
and U4994 (N_4994,N_4656,N_4701);
nor U4995 (N_4995,N_4780,N_4731);
nand U4996 (N_4996,N_4642,N_4684);
or U4997 (N_4997,N_4713,N_4768);
nand U4998 (N_4998,N_4703,N_4603);
or U4999 (N_4999,N_4644,N_4619);
xor UO_0 (O_0,N_4986,N_4848);
and UO_1 (O_1,N_4942,N_4852);
xnor UO_2 (O_2,N_4991,N_4907);
nor UO_3 (O_3,N_4875,N_4914);
or UO_4 (O_4,N_4882,N_4893);
nand UO_5 (O_5,N_4844,N_4885);
xnor UO_6 (O_6,N_4902,N_4845);
or UO_7 (O_7,N_4856,N_4934);
nand UO_8 (O_8,N_4825,N_4941);
xor UO_9 (O_9,N_4888,N_4952);
and UO_10 (O_10,N_4829,N_4842);
nor UO_11 (O_11,N_4815,N_4828);
nand UO_12 (O_12,N_4905,N_4827);
and UO_13 (O_13,N_4841,N_4992);
or UO_14 (O_14,N_4910,N_4811);
nand UO_15 (O_15,N_4831,N_4822);
or UO_16 (O_16,N_4994,N_4923);
nor UO_17 (O_17,N_4961,N_4887);
xor UO_18 (O_18,N_4931,N_4977);
nand UO_19 (O_19,N_4834,N_4929);
nand UO_20 (O_20,N_4908,N_4801);
xor UO_21 (O_21,N_4884,N_4832);
and UO_22 (O_22,N_4867,N_4853);
nand UO_23 (O_23,N_4843,N_4917);
xnor UO_24 (O_24,N_4974,N_4805);
or UO_25 (O_25,N_4895,N_4964);
and UO_26 (O_26,N_4944,N_4836);
xnor UO_27 (O_27,N_4879,N_4892);
nor UO_28 (O_28,N_4876,N_4904);
nor UO_29 (O_29,N_4847,N_4881);
nand UO_30 (O_30,N_4824,N_4948);
xor UO_31 (O_31,N_4858,N_4963);
or UO_32 (O_32,N_4913,N_4800);
and UO_33 (O_33,N_4803,N_4850);
xor UO_34 (O_34,N_4901,N_4922);
or UO_35 (O_35,N_4936,N_4990);
and UO_36 (O_36,N_4810,N_4973);
xnor UO_37 (O_37,N_4865,N_4826);
xnor UO_38 (O_38,N_4946,N_4863);
nand UO_39 (O_39,N_4804,N_4846);
nand UO_40 (O_40,N_4982,N_4959);
xnor UO_41 (O_41,N_4838,N_4993);
or UO_42 (O_42,N_4808,N_4956);
or UO_43 (O_43,N_4919,N_4864);
xnor UO_44 (O_44,N_4812,N_4969);
and UO_45 (O_45,N_4997,N_4830);
nor UO_46 (O_46,N_4880,N_4967);
nor UO_47 (O_47,N_4980,N_4872);
nor UO_48 (O_48,N_4840,N_4947);
xor UO_49 (O_49,N_4886,N_4983);
xnor UO_50 (O_50,N_4978,N_4814);
or UO_51 (O_51,N_4839,N_4817);
nand UO_52 (O_52,N_4945,N_4849);
or UO_53 (O_53,N_4894,N_4968);
nor UO_54 (O_54,N_4949,N_4932);
xnor UO_55 (O_55,N_4873,N_4860);
xor UO_56 (O_56,N_4897,N_4938);
or UO_57 (O_57,N_4970,N_4954);
or UO_58 (O_58,N_4871,N_4889);
and UO_59 (O_59,N_4813,N_4926);
xor UO_60 (O_60,N_4943,N_4918);
nand UO_61 (O_61,N_4953,N_4855);
and UO_62 (O_62,N_4976,N_4835);
xnor UO_63 (O_63,N_4806,N_4935);
nor UO_64 (O_64,N_4821,N_4870);
nand UO_65 (O_65,N_4999,N_4837);
and UO_66 (O_66,N_4874,N_4899);
and UO_67 (O_67,N_4869,N_4903);
or UO_68 (O_68,N_4998,N_4960);
nor UO_69 (O_69,N_4933,N_4802);
or UO_70 (O_70,N_4915,N_4818);
nor UO_71 (O_71,N_4951,N_4891);
nand UO_72 (O_72,N_4854,N_4920);
nor UO_73 (O_73,N_4912,N_4866);
nor UO_74 (O_74,N_4996,N_4950);
nor UO_75 (O_75,N_4809,N_4987);
and UO_76 (O_76,N_4966,N_4930);
or UO_77 (O_77,N_4816,N_4962);
nor UO_78 (O_78,N_4971,N_4958);
and UO_79 (O_79,N_4957,N_4911);
nand UO_80 (O_80,N_4972,N_4979);
or UO_81 (O_81,N_4906,N_4833);
or UO_82 (O_82,N_4900,N_4916);
xnor UO_83 (O_83,N_4862,N_4927);
nor UO_84 (O_84,N_4820,N_4878);
and UO_85 (O_85,N_4995,N_4859);
nor UO_86 (O_86,N_4861,N_4940);
nor UO_87 (O_87,N_4988,N_4890);
and UO_88 (O_88,N_4896,N_4985);
xnor UO_89 (O_89,N_4955,N_4989);
xor UO_90 (O_90,N_4883,N_4819);
or UO_91 (O_91,N_4937,N_4851);
nand UO_92 (O_92,N_4823,N_4924);
nor UO_93 (O_93,N_4877,N_4965);
xnor UO_94 (O_94,N_4928,N_4921);
xnor UO_95 (O_95,N_4925,N_4857);
nor UO_96 (O_96,N_4898,N_4939);
xnor UO_97 (O_97,N_4981,N_4868);
xor UO_98 (O_98,N_4984,N_4909);
xor UO_99 (O_99,N_4975,N_4807);
and UO_100 (O_100,N_4957,N_4837);
nor UO_101 (O_101,N_4906,N_4814);
nor UO_102 (O_102,N_4964,N_4801);
and UO_103 (O_103,N_4922,N_4951);
nand UO_104 (O_104,N_4999,N_4891);
xor UO_105 (O_105,N_4933,N_4864);
and UO_106 (O_106,N_4846,N_4993);
nor UO_107 (O_107,N_4827,N_4961);
nor UO_108 (O_108,N_4888,N_4911);
xnor UO_109 (O_109,N_4942,N_4827);
nor UO_110 (O_110,N_4856,N_4994);
or UO_111 (O_111,N_4888,N_4968);
xnor UO_112 (O_112,N_4917,N_4981);
and UO_113 (O_113,N_4974,N_4944);
nor UO_114 (O_114,N_4954,N_4880);
or UO_115 (O_115,N_4963,N_4929);
xnor UO_116 (O_116,N_4958,N_4816);
xnor UO_117 (O_117,N_4818,N_4874);
xnor UO_118 (O_118,N_4926,N_4916);
xor UO_119 (O_119,N_4826,N_4916);
nor UO_120 (O_120,N_4814,N_4857);
or UO_121 (O_121,N_4924,N_4876);
xor UO_122 (O_122,N_4893,N_4886);
and UO_123 (O_123,N_4883,N_4988);
xnor UO_124 (O_124,N_4975,N_4987);
xnor UO_125 (O_125,N_4912,N_4837);
nor UO_126 (O_126,N_4981,N_4950);
xor UO_127 (O_127,N_4940,N_4944);
nor UO_128 (O_128,N_4835,N_4910);
xor UO_129 (O_129,N_4946,N_4868);
or UO_130 (O_130,N_4855,N_4885);
and UO_131 (O_131,N_4997,N_4978);
nor UO_132 (O_132,N_4889,N_4822);
or UO_133 (O_133,N_4938,N_4872);
xnor UO_134 (O_134,N_4830,N_4932);
and UO_135 (O_135,N_4813,N_4929);
xor UO_136 (O_136,N_4938,N_4860);
nor UO_137 (O_137,N_4953,N_4822);
and UO_138 (O_138,N_4838,N_4823);
or UO_139 (O_139,N_4870,N_4800);
and UO_140 (O_140,N_4981,N_4997);
xor UO_141 (O_141,N_4861,N_4880);
or UO_142 (O_142,N_4886,N_4861);
nand UO_143 (O_143,N_4823,N_4907);
nand UO_144 (O_144,N_4984,N_4883);
and UO_145 (O_145,N_4822,N_4890);
nand UO_146 (O_146,N_4837,N_4908);
xor UO_147 (O_147,N_4830,N_4990);
nand UO_148 (O_148,N_4939,N_4967);
nor UO_149 (O_149,N_4822,N_4825);
nor UO_150 (O_150,N_4832,N_4833);
or UO_151 (O_151,N_4919,N_4913);
or UO_152 (O_152,N_4860,N_4939);
and UO_153 (O_153,N_4972,N_4826);
or UO_154 (O_154,N_4877,N_4810);
nand UO_155 (O_155,N_4858,N_4948);
and UO_156 (O_156,N_4905,N_4832);
nand UO_157 (O_157,N_4822,N_4981);
or UO_158 (O_158,N_4905,N_4952);
and UO_159 (O_159,N_4804,N_4996);
and UO_160 (O_160,N_4804,N_4904);
nand UO_161 (O_161,N_4855,N_4923);
and UO_162 (O_162,N_4961,N_4997);
and UO_163 (O_163,N_4863,N_4902);
xnor UO_164 (O_164,N_4805,N_4821);
nor UO_165 (O_165,N_4828,N_4804);
and UO_166 (O_166,N_4967,N_4831);
nand UO_167 (O_167,N_4819,N_4838);
nand UO_168 (O_168,N_4901,N_4852);
nand UO_169 (O_169,N_4892,N_4992);
nand UO_170 (O_170,N_4956,N_4879);
or UO_171 (O_171,N_4986,N_4909);
xor UO_172 (O_172,N_4887,N_4928);
nand UO_173 (O_173,N_4989,N_4883);
or UO_174 (O_174,N_4987,N_4981);
nand UO_175 (O_175,N_4866,N_4979);
nand UO_176 (O_176,N_4918,N_4953);
nand UO_177 (O_177,N_4835,N_4811);
or UO_178 (O_178,N_4975,N_4888);
or UO_179 (O_179,N_4838,N_4850);
or UO_180 (O_180,N_4905,N_4851);
nand UO_181 (O_181,N_4870,N_4888);
nand UO_182 (O_182,N_4810,N_4845);
or UO_183 (O_183,N_4827,N_4851);
xor UO_184 (O_184,N_4924,N_4884);
nand UO_185 (O_185,N_4949,N_4888);
or UO_186 (O_186,N_4874,N_4992);
nor UO_187 (O_187,N_4955,N_4851);
xnor UO_188 (O_188,N_4896,N_4815);
nor UO_189 (O_189,N_4880,N_4957);
or UO_190 (O_190,N_4878,N_4806);
and UO_191 (O_191,N_4959,N_4848);
and UO_192 (O_192,N_4878,N_4974);
xnor UO_193 (O_193,N_4863,N_4800);
nand UO_194 (O_194,N_4963,N_4924);
xor UO_195 (O_195,N_4864,N_4968);
xnor UO_196 (O_196,N_4840,N_4948);
nor UO_197 (O_197,N_4899,N_4960);
nor UO_198 (O_198,N_4957,N_4914);
nand UO_199 (O_199,N_4858,N_4968);
or UO_200 (O_200,N_4808,N_4868);
nand UO_201 (O_201,N_4854,N_4989);
nand UO_202 (O_202,N_4953,N_4930);
nor UO_203 (O_203,N_4847,N_4899);
xor UO_204 (O_204,N_4806,N_4856);
xnor UO_205 (O_205,N_4997,N_4982);
nor UO_206 (O_206,N_4808,N_4930);
xor UO_207 (O_207,N_4851,N_4954);
nor UO_208 (O_208,N_4866,N_4917);
or UO_209 (O_209,N_4976,N_4862);
or UO_210 (O_210,N_4905,N_4862);
nor UO_211 (O_211,N_4908,N_4988);
and UO_212 (O_212,N_4874,N_4844);
nor UO_213 (O_213,N_4872,N_4987);
xor UO_214 (O_214,N_4884,N_4803);
nand UO_215 (O_215,N_4845,N_4822);
or UO_216 (O_216,N_4821,N_4928);
and UO_217 (O_217,N_4862,N_4986);
xnor UO_218 (O_218,N_4926,N_4891);
nor UO_219 (O_219,N_4835,N_4966);
xor UO_220 (O_220,N_4910,N_4812);
xor UO_221 (O_221,N_4948,N_4958);
and UO_222 (O_222,N_4900,N_4801);
nor UO_223 (O_223,N_4974,N_4946);
or UO_224 (O_224,N_4825,N_4924);
and UO_225 (O_225,N_4905,N_4990);
nor UO_226 (O_226,N_4893,N_4861);
nand UO_227 (O_227,N_4987,N_4978);
nor UO_228 (O_228,N_4802,N_4961);
nand UO_229 (O_229,N_4806,N_4862);
xnor UO_230 (O_230,N_4981,N_4978);
xor UO_231 (O_231,N_4938,N_4944);
nand UO_232 (O_232,N_4937,N_4888);
or UO_233 (O_233,N_4933,N_4857);
nand UO_234 (O_234,N_4869,N_4964);
or UO_235 (O_235,N_4832,N_4893);
nor UO_236 (O_236,N_4910,N_4902);
nor UO_237 (O_237,N_4876,N_4933);
nand UO_238 (O_238,N_4947,N_4909);
nor UO_239 (O_239,N_4844,N_4806);
xnor UO_240 (O_240,N_4851,N_4847);
or UO_241 (O_241,N_4849,N_4979);
or UO_242 (O_242,N_4993,N_4820);
xnor UO_243 (O_243,N_4957,N_4947);
xnor UO_244 (O_244,N_4821,N_4862);
nand UO_245 (O_245,N_4908,N_4967);
nor UO_246 (O_246,N_4993,N_4832);
or UO_247 (O_247,N_4834,N_4920);
xnor UO_248 (O_248,N_4949,N_4934);
xnor UO_249 (O_249,N_4888,N_4981);
nand UO_250 (O_250,N_4817,N_4997);
nand UO_251 (O_251,N_4842,N_4964);
nor UO_252 (O_252,N_4825,N_4844);
or UO_253 (O_253,N_4835,N_4987);
xnor UO_254 (O_254,N_4991,N_4996);
or UO_255 (O_255,N_4898,N_4964);
and UO_256 (O_256,N_4828,N_4964);
or UO_257 (O_257,N_4823,N_4895);
and UO_258 (O_258,N_4842,N_4811);
and UO_259 (O_259,N_4915,N_4945);
or UO_260 (O_260,N_4933,N_4911);
or UO_261 (O_261,N_4935,N_4844);
xor UO_262 (O_262,N_4841,N_4845);
or UO_263 (O_263,N_4899,N_4817);
and UO_264 (O_264,N_4983,N_4823);
and UO_265 (O_265,N_4996,N_4833);
nor UO_266 (O_266,N_4896,N_4963);
xor UO_267 (O_267,N_4928,N_4929);
xnor UO_268 (O_268,N_4892,N_4956);
nor UO_269 (O_269,N_4822,N_4861);
and UO_270 (O_270,N_4889,N_4839);
xor UO_271 (O_271,N_4859,N_4993);
nand UO_272 (O_272,N_4800,N_4918);
nor UO_273 (O_273,N_4810,N_4908);
or UO_274 (O_274,N_4907,N_4934);
nor UO_275 (O_275,N_4816,N_4830);
nor UO_276 (O_276,N_4883,N_4923);
or UO_277 (O_277,N_4931,N_4823);
and UO_278 (O_278,N_4929,N_4974);
or UO_279 (O_279,N_4964,N_4825);
nor UO_280 (O_280,N_4871,N_4929);
nand UO_281 (O_281,N_4869,N_4974);
nand UO_282 (O_282,N_4948,N_4857);
xor UO_283 (O_283,N_4812,N_4811);
nand UO_284 (O_284,N_4837,N_4909);
nand UO_285 (O_285,N_4860,N_4931);
xnor UO_286 (O_286,N_4845,N_4961);
nand UO_287 (O_287,N_4944,N_4922);
or UO_288 (O_288,N_4922,N_4948);
nand UO_289 (O_289,N_4854,N_4897);
xnor UO_290 (O_290,N_4924,N_4836);
xnor UO_291 (O_291,N_4864,N_4830);
and UO_292 (O_292,N_4874,N_4993);
nor UO_293 (O_293,N_4963,N_4944);
and UO_294 (O_294,N_4881,N_4978);
or UO_295 (O_295,N_4820,N_4903);
and UO_296 (O_296,N_4939,N_4829);
nand UO_297 (O_297,N_4921,N_4916);
and UO_298 (O_298,N_4912,N_4819);
xnor UO_299 (O_299,N_4935,N_4829);
nor UO_300 (O_300,N_4997,N_4966);
and UO_301 (O_301,N_4999,N_4822);
nand UO_302 (O_302,N_4955,N_4862);
or UO_303 (O_303,N_4842,N_4900);
nand UO_304 (O_304,N_4858,N_4885);
xnor UO_305 (O_305,N_4988,N_4893);
xor UO_306 (O_306,N_4895,N_4829);
xor UO_307 (O_307,N_4987,N_4924);
and UO_308 (O_308,N_4852,N_4974);
and UO_309 (O_309,N_4993,N_4929);
xor UO_310 (O_310,N_4962,N_4911);
and UO_311 (O_311,N_4990,N_4821);
nor UO_312 (O_312,N_4994,N_4876);
or UO_313 (O_313,N_4897,N_4807);
nor UO_314 (O_314,N_4979,N_4896);
and UO_315 (O_315,N_4949,N_4913);
nor UO_316 (O_316,N_4997,N_4962);
nand UO_317 (O_317,N_4898,N_4977);
xor UO_318 (O_318,N_4817,N_4964);
nand UO_319 (O_319,N_4891,N_4873);
xnor UO_320 (O_320,N_4910,N_4973);
and UO_321 (O_321,N_4886,N_4991);
or UO_322 (O_322,N_4874,N_4894);
and UO_323 (O_323,N_4878,N_4857);
nor UO_324 (O_324,N_4859,N_4954);
or UO_325 (O_325,N_4817,N_4963);
nor UO_326 (O_326,N_4902,N_4911);
nand UO_327 (O_327,N_4830,N_4894);
nor UO_328 (O_328,N_4832,N_4859);
and UO_329 (O_329,N_4997,N_4827);
nor UO_330 (O_330,N_4854,N_4803);
or UO_331 (O_331,N_4876,N_4886);
or UO_332 (O_332,N_4999,N_4874);
and UO_333 (O_333,N_4964,N_4805);
nand UO_334 (O_334,N_4965,N_4827);
nor UO_335 (O_335,N_4891,N_4833);
and UO_336 (O_336,N_4838,N_4841);
xnor UO_337 (O_337,N_4866,N_4901);
and UO_338 (O_338,N_4830,N_4821);
or UO_339 (O_339,N_4860,N_4868);
nor UO_340 (O_340,N_4949,N_4931);
nor UO_341 (O_341,N_4987,N_4832);
nand UO_342 (O_342,N_4837,N_4818);
and UO_343 (O_343,N_4935,N_4889);
xor UO_344 (O_344,N_4991,N_4880);
nand UO_345 (O_345,N_4957,N_4996);
nand UO_346 (O_346,N_4833,N_4912);
nor UO_347 (O_347,N_4945,N_4909);
nand UO_348 (O_348,N_4964,N_4823);
and UO_349 (O_349,N_4933,N_4807);
and UO_350 (O_350,N_4980,N_4910);
and UO_351 (O_351,N_4918,N_4841);
or UO_352 (O_352,N_4991,N_4941);
nand UO_353 (O_353,N_4813,N_4821);
or UO_354 (O_354,N_4895,N_4903);
or UO_355 (O_355,N_4877,N_4804);
nand UO_356 (O_356,N_4904,N_4906);
or UO_357 (O_357,N_4818,N_4867);
and UO_358 (O_358,N_4858,N_4834);
or UO_359 (O_359,N_4845,N_4994);
or UO_360 (O_360,N_4904,N_4998);
and UO_361 (O_361,N_4828,N_4931);
and UO_362 (O_362,N_4898,N_4931);
and UO_363 (O_363,N_4964,N_4972);
nand UO_364 (O_364,N_4898,N_4829);
and UO_365 (O_365,N_4914,N_4864);
and UO_366 (O_366,N_4863,N_4856);
nor UO_367 (O_367,N_4835,N_4864);
nand UO_368 (O_368,N_4807,N_4991);
nand UO_369 (O_369,N_4988,N_4830);
or UO_370 (O_370,N_4801,N_4830);
or UO_371 (O_371,N_4865,N_4959);
nor UO_372 (O_372,N_4867,N_4850);
or UO_373 (O_373,N_4876,N_4856);
and UO_374 (O_374,N_4933,N_4805);
and UO_375 (O_375,N_4824,N_4977);
and UO_376 (O_376,N_4973,N_4996);
nor UO_377 (O_377,N_4996,N_4933);
nand UO_378 (O_378,N_4919,N_4946);
nand UO_379 (O_379,N_4983,N_4975);
or UO_380 (O_380,N_4852,N_4964);
nor UO_381 (O_381,N_4917,N_4803);
or UO_382 (O_382,N_4852,N_4809);
nor UO_383 (O_383,N_4936,N_4814);
or UO_384 (O_384,N_4893,N_4985);
nand UO_385 (O_385,N_4902,N_4893);
nor UO_386 (O_386,N_4875,N_4902);
nand UO_387 (O_387,N_4976,N_4879);
xor UO_388 (O_388,N_4939,N_4938);
xnor UO_389 (O_389,N_4861,N_4885);
xnor UO_390 (O_390,N_4844,N_4882);
and UO_391 (O_391,N_4919,N_4966);
or UO_392 (O_392,N_4929,N_4828);
nor UO_393 (O_393,N_4807,N_4839);
nor UO_394 (O_394,N_4805,N_4865);
or UO_395 (O_395,N_4883,N_4964);
nor UO_396 (O_396,N_4972,N_4977);
xnor UO_397 (O_397,N_4987,N_4914);
and UO_398 (O_398,N_4951,N_4903);
and UO_399 (O_399,N_4846,N_4888);
nor UO_400 (O_400,N_4913,N_4971);
and UO_401 (O_401,N_4886,N_4951);
and UO_402 (O_402,N_4997,N_4977);
nand UO_403 (O_403,N_4855,N_4859);
or UO_404 (O_404,N_4972,N_4858);
xnor UO_405 (O_405,N_4937,N_4906);
or UO_406 (O_406,N_4983,N_4824);
nor UO_407 (O_407,N_4926,N_4940);
or UO_408 (O_408,N_4885,N_4847);
xnor UO_409 (O_409,N_4885,N_4955);
or UO_410 (O_410,N_4837,N_4921);
nand UO_411 (O_411,N_4837,N_4905);
nor UO_412 (O_412,N_4902,N_4825);
and UO_413 (O_413,N_4837,N_4858);
or UO_414 (O_414,N_4962,N_4852);
nand UO_415 (O_415,N_4805,N_4948);
and UO_416 (O_416,N_4943,N_4833);
and UO_417 (O_417,N_4857,N_4843);
xor UO_418 (O_418,N_4916,N_4966);
nand UO_419 (O_419,N_4837,N_4982);
nand UO_420 (O_420,N_4802,N_4921);
or UO_421 (O_421,N_4895,N_4979);
or UO_422 (O_422,N_4828,N_4984);
nand UO_423 (O_423,N_4801,N_4945);
and UO_424 (O_424,N_4951,N_4906);
nor UO_425 (O_425,N_4902,N_4888);
and UO_426 (O_426,N_4867,N_4843);
nand UO_427 (O_427,N_4823,N_4985);
nand UO_428 (O_428,N_4897,N_4931);
or UO_429 (O_429,N_4880,N_4859);
xor UO_430 (O_430,N_4818,N_4888);
nor UO_431 (O_431,N_4822,N_4812);
xnor UO_432 (O_432,N_4942,N_4945);
nor UO_433 (O_433,N_4957,N_4828);
and UO_434 (O_434,N_4905,N_4870);
nand UO_435 (O_435,N_4841,N_4835);
xor UO_436 (O_436,N_4958,N_4966);
and UO_437 (O_437,N_4993,N_4814);
xor UO_438 (O_438,N_4957,N_4928);
or UO_439 (O_439,N_4822,N_4884);
or UO_440 (O_440,N_4839,N_4856);
xor UO_441 (O_441,N_4973,N_4987);
xor UO_442 (O_442,N_4950,N_4908);
xor UO_443 (O_443,N_4834,N_4962);
and UO_444 (O_444,N_4850,N_4907);
xor UO_445 (O_445,N_4810,N_4966);
or UO_446 (O_446,N_4806,N_4803);
xor UO_447 (O_447,N_4967,N_4882);
and UO_448 (O_448,N_4929,N_4896);
nor UO_449 (O_449,N_4839,N_4914);
xnor UO_450 (O_450,N_4951,N_4809);
and UO_451 (O_451,N_4909,N_4899);
nand UO_452 (O_452,N_4879,N_4904);
nor UO_453 (O_453,N_4877,N_4989);
nor UO_454 (O_454,N_4927,N_4994);
nand UO_455 (O_455,N_4993,N_4987);
xor UO_456 (O_456,N_4966,N_4909);
nand UO_457 (O_457,N_4970,N_4852);
or UO_458 (O_458,N_4820,N_4836);
or UO_459 (O_459,N_4832,N_4872);
nor UO_460 (O_460,N_4848,N_4842);
nor UO_461 (O_461,N_4976,N_4907);
nor UO_462 (O_462,N_4970,N_4995);
and UO_463 (O_463,N_4885,N_4970);
or UO_464 (O_464,N_4895,N_4890);
and UO_465 (O_465,N_4984,N_4840);
nand UO_466 (O_466,N_4951,N_4812);
nor UO_467 (O_467,N_4938,N_4937);
nand UO_468 (O_468,N_4999,N_4952);
and UO_469 (O_469,N_4950,N_4859);
xor UO_470 (O_470,N_4839,N_4873);
and UO_471 (O_471,N_4909,N_4940);
or UO_472 (O_472,N_4929,N_4899);
xnor UO_473 (O_473,N_4961,N_4826);
xor UO_474 (O_474,N_4979,N_4904);
nand UO_475 (O_475,N_4830,N_4950);
or UO_476 (O_476,N_4809,N_4988);
nand UO_477 (O_477,N_4994,N_4989);
nand UO_478 (O_478,N_4981,N_4957);
and UO_479 (O_479,N_4908,N_4982);
and UO_480 (O_480,N_4967,N_4957);
and UO_481 (O_481,N_4869,N_4917);
nor UO_482 (O_482,N_4937,N_4915);
or UO_483 (O_483,N_4945,N_4861);
xnor UO_484 (O_484,N_4920,N_4939);
nor UO_485 (O_485,N_4894,N_4984);
nand UO_486 (O_486,N_4811,N_4956);
xor UO_487 (O_487,N_4916,N_4863);
nand UO_488 (O_488,N_4943,N_4914);
nor UO_489 (O_489,N_4998,N_4978);
nand UO_490 (O_490,N_4845,N_4914);
xor UO_491 (O_491,N_4830,N_4882);
or UO_492 (O_492,N_4812,N_4943);
nor UO_493 (O_493,N_4941,N_4838);
nand UO_494 (O_494,N_4959,N_4859);
and UO_495 (O_495,N_4970,N_4860);
nand UO_496 (O_496,N_4919,N_4997);
or UO_497 (O_497,N_4865,N_4896);
and UO_498 (O_498,N_4906,N_4929);
and UO_499 (O_499,N_4855,N_4899);
or UO_500 (O_500,N_4967,N_4803);
xor UO_501 (O_501,N_4844,N_4991);
or UO_502 (O_502,N_4916,N_4913);
xor UO_503 (O_503,N_4853,N_4910);
nor UO_504 (O_504,N_4943,N_4857);
and UO_505 (O_505,N_4878,N_4860);
nor UO_506 (O_506,N_4928,N_4807);
nor UO_507 (O_507,N_4813,N_4875);
or UO_508 (O_508,N_4958,N_4830);
nand UO_509 (O_509,N_4943,N_4810);
nand UO_510 (O_510,N_4916,N_4825);
xnor UO_511 (O_511,N_4972,N_4867);
xnor UO_512 (O_512,N_4878,N_4922);
nand UO_513 (O_513,N_4958,N_4979);
nor UO_514 (O_514,N_4843,N_4929);
or UO_515 (O_515,N_4853,N_4851);
xnor UO_516 (O_516,N_4872,N_4809);
nor UO_517 (O_517,N_4850,N_4886);
nor UO_518 (O_518,N_4888,N_4880);
or UO_519 (O_519,N_4928,N_4920);
and UO_520 (O_520,N_4963,N_4987);
and UO_521 (O_521,N_4872,N_4921);
nor UO_522 (O_522,N_4966,N_4894);
and UO_523 (O_523,N_4802,N_4807);
xor UO_524 (O_524,N_4813,N_4842);
and UO_525 (O_525,N_4842,N_4927);
and UO_526 (O_526,N_4946,N_4826);
nor UO_527 (O_527,N_4948,N_4834);
and UO_528 (O_528,N_4922,N_4847);
nand UO_529 (O_529,N_4946,N_4925);
nor UO_530 (O_530,N_4872,N_4970);
xnor UO_531 (O_531,N_4837,N_4855);
nand UO_532 (O_532,N_4914,N_4962);
nand UO_533 (O_533,N_4868,N_4991);
nor UO_534 (O_534,N_4869,N_4884);
and UO_535 (O_535,N_4891,N_4915);
and UO_536 (O_536,N_4817,N_4824);
and UO_537 (O_537,N_4855,N_4988);
xnor UO_538 (O_538,N_4815,N_4950);
and UO_539 (O_539,N_4829,N_4967);
nand UO_540 (O_540,N_4879,N_4893);
nand UO_541 (O_541,N_4927,N_4931);
nand UO_542 (O_542,N_4859,N_4915);
xnor UO_543 (O_543,N_4934,N_4841);
nor UO_544 (O_544,N_4831,N_4931);
nor UO_545 (O_545,N_4866,N_4882);
nand UO_546 (O_546,N_4932,N_4982);
and UO_547 (O_547,N_4885,N_4866);
xor UO_548 (O_548,N_4816,N_4942);
nor UO_549 (O_549,N_4821,N_4940);
xnor UO_550 (O_550,N_4836,N_4863);
nand UO_551 (O_551,N_4881,N_4874);
or UO_552 (O_552,N_4870,N_4893);
nor UO_553 (O_553,N_4985,N_4845);
nor UO_554 (O_554,N_4814,N_4967);
xor UO_555 (O_555,N_4848,N_4871);
and UO_556 (O_556,N_4987,N_4820);
nand UO_557 (O_557,N_4960,N_4802);
xnor UO_558 (O_558,N_4812,N_4813);
or UO_559 (O_559,N_4965,N_4914);
nor UO_560 (O_560,N_4874,N_4997);
nand UO_561 (O_561,N_4870,N_4933);
or UO_562 (O_562,N_4863,N_4992);
or UO_563 (O_563,N_4963,N_4980);
nor UO_564 (O_564,N_4860,N_4827);
nor UO_565 (O_565,N_4815,N_4985);
xnor UO_566 (O_566,N_4873,N_4946);
nor UO_567 (O_567,N_4912,N_4812);
and UO_568 (O_568,N_4840,N_4942);
and UO_569 (O_569,N_4852,N_4872);
xnor UO_570 (O_570,N_4961,N_4890);
or UO_571 (O_571,N_4918,N_4803);
and UO_572 (O_572,N_4995,N_4918);
xnor UO_573 (O_573,N_4913,N_4948);
and UO_574 (O_574,N_4805,N_4811);
nand UO_575 (O_575,N_4812,N_4939);
xor UO_576 (O_576,N_4856,N_4975);
or UO_577 (O_577,N_4831,N_4827);
and UO_578 (O_578,N_4983,N_4856);
or UO_579 (O_579,N_4874,N_4902);
or UO_580 (O_580,N_4980,N_4971);
nand UO_581 (O_581,N_4968,N_4990);
or UO_582 (O_582,N_4906,N_4848);
nand UO_583 (O_583,N_4855,N_4935);
and UO_584 (O_584,N_4961,N_4859);
nor UO_585 (O_585,N_4865,N_4848);
xor UO_586 (O_586,N_4923,N_4891);
and UO_587 (O_587,N_4848,N_4876);
xor UO_588 (O_588,N_4872,N_4946);
or UO_589 (O_589,N_4808,N_4994);
xnor UO_590 (O_590,N_4938,N_4934);
nand UO_591 (O_591,N_4976,N_4893);
or UO_592 (O_592,N_4828,N_4993);
xnor UO_593 (O_593,N_4950,N_4888);
xnor UO_594 (O_594,N_4814,N_4917);
and UO_595 (O_595,N_4997,N_4931);
and UO_596 (O_596,N_4873,N_4927);
nor UO_597 (O_597,N_4945,N_4885);
and UO_598 (O_598,N_4991,N_4937);
or UO_599 (O_599,N_4869,N_4910);
and UO_600 (O_600,N_4846,N_4840);
nand UO_601 (O_601,N_4825,N_4866);
and UO_602 (O_602,N_4841,N_4929);
nand UO_603 (O_603,N_4964,N_4879);
and UO_604 (O_604,N_4881,N_4971);
and UO_605 (O_605,N_4904,N_4938);
or UO_606 (O_606,N_4948,N_4823);
xnor UO_607 (O_607,N_4952,N_4894);
or UO_608 (O_608,N_4996,N_4825);
or UO_609 (O_609,N_4859,N_4823);
xor UO_610 (O_610,N_4958,N_4959);
nand UO_611 (O_611,N_4985,N_4824);
and UO_612 (O_612,N_4950,N_4898);
nand UO_613 (O_613,N_4837,N_4913);
or UO_614 (O_614,N_4807,N_4987);
xnor UO_615 (O_615,N_4977,N_4991);
xnor UO_616 (O_616,N_4992,N_4846);
or UO_617 (O_617,N_4899,N_4934);
and UO_618 (O_618,N_4914,N_4933);
or UO_619 (O_619,N_4877,N_4913);
or UO_620 (O_620,N_4803,N_4821);
nand UO_621 (O_621,N_4928,N_4911);
nor UO_622 (O_622,N_4835,N_4963);
or UO_623 (O_623,N_4919,N_4961);
or UO_624 (O_624,N_4906,N_4889);
or UO_625 (O_625,N_4988,N_4840);
and UO_626 (O_626,N_4803,N_4979);
nand UO_627 (O_627,N_4880,N_4817);
xnor UO_628 (O_628,N_4829,N_4824);
nor UO_629 (O_629,N_4901,N_4960);
or UO_630 (O_630,N_4851,N_4830);
xor UO_631 (O_631,N_4925,N_4871);
or UO_632 (O_632,N_4841,N_4836);
and UO_633 (O_633,N_4953,N_4846);
and UO_634 (O_634,N_4920,N_4911);
xnor UO_635 (O_635,N_4882,N_4991);
and UO_636 (O_636,N_4941,N_4923);
nor UO_637 (O_637,N_4881,N_4990);
and UO_638 (O_638,N_4831,N_4987);
nand UO_639 (O_639,N_4820,N_4846);
and UO_640 (O_640,N_4929,N_4867);
xnor UO_641 (O_641,N_4883,N_4805);
nor UO_642 (O_642,N_4873,N_4884);
and UO_643 (O_643,N_4951,N_4934);
or UO_644 (O_644,N_4836,N_4855);
nand UO_645 (O_645,N_4816,N_4921);
and UO_646 (O_646,N_4842,N_4905);
and UO_647 (O_647,N_4830,N_4860);
xor UO_648 (O_648,N_4943,N_4930);
or UO_649 (O_649,N_4824,N_4952);
nor UO_650 (O_650,N_4865,N_4869);
and UO_651 (O_651,N_4936,N_4865);
or UO_652 (O_652,N_4883,N_4910);
and UO_653 (O_653,N_4860,N_4940);
nor UO_654 (O_654,N_4869,N_4914);
and UO_655 (O_655,N_4817,N_4966);
nand UO_656 (O_656,N_4891,N_4912);
xnor UO_657 (O_657,N_4985,N_4869);
and UO_658 (O_658,N_4952,N_4802);
and UO_659 (O_659,N_4963,N_4844);
xor UO_660 (O_660,N_4888,N_4807);
nor UO_661 (O_661,N_4841,N_4982);
nand UO_662 (O_662,N_4954,N_4931);
xor UO_663 (O_663,N_4875,N_4968);
nor UO_664 (O_664,N_4952,N_4815);
or UO_665 (O_665,N_4886,N_4914);
nand UO_666 (O_666,N_4816,N_4843);
xor UO_667 (O_667,N_4970,N_4881);
nand UO_668 (O_668,N_4887,N_4951);
xnor UO_669 (O_669,N_4980,N_4916);
nor UO_670 (O_670,N_4880,N_4846);
and UO_671 (O_671,N_4818,N_4894);
and UO_672 (O_672,N_4870,N_4921);
and UO_673 (O_673,N_4914,N_4991);
and UO_674 (O_674,N_4905,N_4882);
or UO_675 (O_675,N_4986,N_4838);
xnor UO_676 (O_676,N_4953,N_4980);
xor UO_677 (O_677,N_4955,N_4816);
nand UO_678 (O_678,N_4956,N_4832);
nand UO_679 (O_679,N_4865,N_4850);
or UO_680 (O_680,N_4845,N_4996);
or UO_681 (O_681,N_4940,N_4827);
or UO_682 (O_682,N_4951,N_4950);
xor UO_683 (O_683,N_4881,N_4878);
or UO_684 (O_684,N_4979,N_4875);
nand UO_685 (O_685,N_4903,N_4962);
or UO_686 (O_686,N_4890,N_4891);
nand UO_687 (O_687,N_4893,N_4977);
or UO_688 (O_688,N_4866,N_4950);
nand UO_689 (O_689,N_4837,N_4956);
or UO_690 (O_690,N_4991,N_4864);
or UO_691 (O_691,N_4990,N_4975);
or UO_692 (O_692,N_4952,N_4848);
xor UO_693 (O_693,N_4897,N_4907);
nor UO_694 (O_694,N_4985,N_4836);
nand UO_695 (O_695,N_4856,N_4958);
nor UO_696 (O_696,N_4908,N_4871);
nor UO_697 (O_697,N_4938,N_4804);
xor UO_698 (O_698,N_4804,N_4832);
nand UO_699 (O_699,N_4945,N_4857);
nand UO_700 (O_700,N_4998,N_4913);
nand UO_701 (O_701,N_4814,N_4853);
and UO_702 (O_702,N_4899,N_4806);
and UO_703 (O_703,N_4839,N_4991);
nand UO_704 (O_704,N_4865,N_4957);
and UO_705 (O_705,N_4880,N_4981);
nand UO_706 (O_706,N_4960,N_4971);
and UO_707 (O_707,N_4807,N_4924);
nand UO_708 (O_708,N_4982,N_4995);
nor UO_709 (O_709,N_4851,N_4907);
xnor UO_710 (O_710,N_4918,N_4849);
nand UO_711 (O_711,N_4813,N_4800);
nand UO_712 (O_712,N_4854,N_4917);
and UO_713 (O_713,N_4820,N_4853);
xor UO_714 (O_714,N_4960,N_4804);
or UO_715 (O_715,N_4958,N_4986);
nand UO_716 (O_716,N_4978,N_4824);
xnor UO_717 (O_717,N_4937,N_4993);
or UO_718 (O_718,N_4910,N_4970);
and UO_719 (O_719,N_4939,N_4893);
xor UO_720 (O_720,N_4837,N_4943);
nor UO_721 (O_721,N_4979,N_4974);
nand UO_722 (O_722,N_4888,N_4820);
or UO_723 (O_723,N_4834,N_4906);
or UO_724 (O_724,N_4873,N_4983);
and UO_725 (O_725,N_4840,N_4861);
or UO_726 (O_726,N_4968,N_4887);
or UO_727 (O_727,N_4839,N_4879);
xnor UO_728 (O_728,N_4886,N_4800);
and UO_729 (O_729,N_4849,N_4924);
and UO_730 (O_730,N_4934,N_4883);
nand UO_731 (O_731,N_4946,N_4857);
xnor UO_732 (O_732,N_4903,N_4875);
nor UO_733 (O_733,N_4855,N_4866);
xnor UO_734 (O_734,N_4920,N_4865);
and UO_735 (O_735,N_4919,N_4877);
or UO_736 (O_736,N_4892,N_4903);
xnor UO_737 (O_737,N_4856,N_4973);
nor UO_738 (O_738,N_4902,N_4940);
or UO_739 (O_739,N_4837,N_4915);
xnor UO_740 (O_740,N_4825,N_4840);
nor UO_741 (O_741,N_4837,N_4845);
nor UO_742 (O_742,N_4902,N_4958);
or UO_743 (O_743,N_4872,N_4904);
and UO_744 (O_744,N_4993,N_4844);
or UO_745 (O_745,N_4817,N_4832);
nor UO_746 (O_746,N_4896,N_4923);
and UO_747 (O_747,N_4943,N_4800);
xor UO_748 (O_748,N_4923,N_4986);
nor UO_749 (O_749,N_4854,N_4991);
and UO_750 (O_750,N_4987,N_4898);
and UO_751 (O_751,N_4803,N_4843);
nand UO_752 (O_752,N_4815,N_4850);
nor UO_753 (O_753,N_4840,N_4821);
and UO_754 (O_754,N_4891,N_4835);
xnor UO_755 (O_755,N_4939,N_4964);
nor UO_756 (O_756,N_4996,N_4931);
nor UO_757 (O_757,N_4907,N_4915);
and UO_758 (O_758,N_4902,N_4838);
nor UO_759 (O_759,N_4894,N_4941);
xor UO_760 (O_760,N_4852,N_4814);
and UO_761 (O_761,N_4883,N_4832);
nor UO_762 (O_762,N_4935,N_4905);
and UO_763 (O_763,N_4821,N_4933);
or UO_764 (O_764,N_4944,N_4952);
nor UO_765 (O_765,N_4829,N_4984);
and UO_766 (O_766,N_4912,N_4934);
and UO_767 (O_767,N_4934,N_4825);
nor UO_768 (O_768,N_4888,N_4924);
nor UO_769 (O_769,N_4853,N_4838);
nor UO_770 (O_770,N_4881,N_4997);
nor UO_771 (O_771,N_4970,N_4832);
and UO_772 (O_772,N_4983,N_4979);
xnor UO_773 (O_773,N_4991,N_4918);
nor UO_774 (O_774,N_4960,N_4886);
nand UO_775 (O_775,N_4836,N_4947);
nor UO_776 (O_776,N_4895,N_4801);
nor UO_777 (O_777,N_4905,N_4841);
xnor UO_778 (O_778,N_4908,N_4869);
nand UO_779 (O_779,N_4806,N_4852);
nand UO_780 (O_780,N_4999,N_4856);
nand UO_781 (O_781,N_4917,N_4897);
and UO_782 (O_782,N_4924,N_4886);
xnor UO_783 (O_783,N_4883,N_4882);
xnor UO_784 (O_784,N_4874,N_4915);
nor UO_785 (O_785,N_4960,N_4893);
or UO_786 (O_786,N_4810,N_4956);
and UO_787 (O_787,N_4845,N_4935);
or UO_788 (O_788,N_4842,N_4928);
nand UO_789 (O_789,N_4919,N_4977);
or UO_790 (O_790,N_4927,N_4996);
or UO_791 (O_791,N_4836,N_4962);
nor UO_792 (O_792,N_4871,N_4820);
or UO_793 (O_793,N_4832,N_4984);
xor UO_794 (O_794,N_4915,N_4807);
xor UO_795 (O_795,N_4958,N_4822);
nand UO_796 (O_796,N_4855,N_4984);
or UO_797 (O_797,N_4851,N_4837);
nor UO_798 (O_798,N_4958,N_4812);
xor UO_799 (O_799,N_4886,N_4870);
nor UO_800 (O_800,N_4925,N_4802);
and UO_801 (O_801,N_4870,N_4938);
xnor UO_802 (O_802,N_4998,N_4874);
or UO_803 (O_803,N_4881,N_4943);
nor UO_804 (O_804,N_4807,N_4881);
nand UO_805 (O_805,N_4928,N_4940);
nand UO_806 (O_806,N_4842,N_4812);
nand UO_807 (O_807,N_4941,N_4852);
or UO_808 (O_808,N_4804,N_4822);
and UO_809 (O_809,N_4832,N_4854);
nor UO_810 (O_810,N_4829,N_4840);
xnor UO_811 (O_811,N_4814,N_4921);
nor UO_812 (O_812,N_4847,N_4908);
nor UO_813 (O_813,N_4839,N_4910);
or UO_814 (O_814,N_4920,N_4914);
nor UO_815 (O_815,N_4917,N_4922);
xnor UO_816 (O_816,N_4875,N_4825);
and UO_817 (O_817,N_4992,N_4839);
nand UO_818 (O_818,N_4942,N_4995);
and UO_819 (O_819,N_4947,N_4964);
or UO_820 (O_820,N_4925,N_4851);
nor UO_821 (O_821,N_4972,N_4939);
xnor UO_822 (O_822,N_4822,N_4820);
or UO_823 (O_823,N_4884,N_4912);
xnor UO_824 (O_824,N_4854,N_4850);
and UO_825 (O_825,N_4869,N_4982);
nor UO_826 (O_826,N_4865,N_4997);
xnor UO_827 (O_827,N_4983,N_4948);
xor UO_828 (O_828,N_4817,N_4876);
xnor UO_829 (O_829,N_4860,N_4988);
nor UO_830 (O_830,N_4865,N_4886);
nand UO_831 (O_831,N_4955,N_4850);
or UO_832 (O_832,N_4874,N_4848);
or UO_833 (O_833,N_4832,N_4814);
or UO_834 (O_834,N_4939,N_4921);
nand UO_835 (O_835,N_4929,N_4979);
and UO_836 (O_836,N_4904,N_4916);
or UO_837 (O_837,N_4890,N_4864);
or UO_838 (O_838,N_4817,N_4866);
nor UO_839 (O_839,N_4956,N_4965);
nor UO_840 (O_840,N_4994,N_4993);
nor UO_841 (O_841,N_4991,N_4848);
nand UO_842 (O_842,N_4849,N_4892);
and UO_843 (O_843,N_4841,N_4890);
nor UO_844 (O_844,N_4992,N_4953);
or UO_845 (O_845,N_4838,N_4835);
nand UO_846 (O_846,N_4834,N_4848);
or UO_847 (O_847,N_4801,N_4983);
or UO_848 (O_848,N_4955,N_4911);
nor UO_849 (O_849,N_4986,N_4830);
xor UO_850 (O_850,N_4880,N_4895);
and UO_851 (O_851,N_4850,N_4942);
nor UO_852 (O_852,N_4988,N_4805);
xor UO_853 (O_853,N_4960,N_4831);
and UO_854 (O_854,N_4909,N_4876);
nand UO_855 (O_855,N_4973,N_4907);
xor UO_856 (O_856,N_4885,N_4846);
nand UO_857 (O_857,N_4937,N_4988);
xnor UO_858 (O_858,N_4912,N_4937);
and UO_859 (O_859,N_4897,N_4851);
nand UO_860 (O_860,N_4867,N_4963);
or UO_861 (O_861,N_4900,N_4949);
or UO_862 (O_862,N_4964,N_4938);
and UO_863 (O_863,N_4867,N_4863);
nand UO_864 (O_864,N_4872,N_4803);
xor UO_865 (O_865,N_4810,N_4971);
nand UO_866 (O_866,N_4973,N_4864);
nand UO_867 (O_867,N_4855,N_4871);
or UO_868 (O_868,N_4891,N_4906);
nor UO_869 (O_869,N_4966,N_4818);
or UO_870 (O_870,N_4880,N_4807);
and UO_871 (O_871,N_4875,N_4909);
xor UO_872 (O_872,N_4848,N_4826);
xnor UO_873 (O_873,N_4804,N_4851);
nand UO_874 (O_874,N_4887,N_4918);
xnor UO_875 (O_875,N_4935,N_4881);
xnor UO_876 (O_876,N_4871,N_4894);
nand UO_877 (O_877,N_4949,N_4833);
or UO_878 (O_878,N_4813,N_4844);
or UO_879 (O_879,N_4812,N_4980);
nor UO_880 (O_880,N_4910,N_4941);
nor UO_881 (O_881,N_4843,N_4955);
xnor UO_882 (O_882,N_4961,N_4969);
xor UO_883 (O_883,N_4996,N_4911);
xor UO_884 (O_884,N_4925,N_4924);
or UO_885 (O_885,N_4965,N_4992);
and UO_886 (O_886,N_4942,N_4962);
nor UO_887 (O_887,N_4842,N_4893);
xor UO_888 (O_888,N_4947,N_4887);
nand UO_889 (O_889,N_4858,N_4882);
and UO_890 (O_890,N_4914,N_4992);
or UO_891 (O_891,N_4827,N_4878);
xor UO_892 (O_892,N_4986,N_4881);
nor UO_893 (O_893,N_4916,N_4816);
and UO_894 (O_894,N_4927,N_4848);
nor UO_895 (O_895,N_4911,N_4815);
or UO_896 (O_896,N_4936,N_4892);
nor UO_897 (O_897,N_4814,N_4915);
nand UO_898 (O_898,N_4901,N_4918);
nand UO_899 (O_899,N_4923,N_4989);
or UO_900 (O_900,N_4856,N_4939);
and UO_901 (O_901,N_4833,N_4903);
or UO_902 (O_902,N_4911,N_4967);
and UO_903 (O_903,N_4826,N_4881);
nor UO_904 (O_904,N_4866,N_4897);
xor UO_905 (O_905,N_4972,N_4922);
and UO_906 (O_906,N_4845,N_4904);
or UO_907 (O_907,N_4988,N_4917);
nand UO_908 (O_908,N_4976,N_4874);
and UO_909 (O_909,N_4820,N_4960);
xnor UO_910 (O_910,N_4840,N_4875);
xor UO_911 (O_911,N_4914,N_4821);
or UO_912 (O_912,N_4829,N_4878);
nor UO_913 (O_913,N_4832,N_4925);
xor UO_914 (O_914,N_4952,N_4906);
xor UO_915 (O_915,N_4914,N_4942);
xnor UO_916 (O_916,N_4853,N_4909);
xnor UO_917 (O_917,N_4850,N_4839);
nor UO_918 (O_918,N_4905,N_4911);
xor UO_919 (O_919,N_4847,N_4807);
nand UO_920 (O_920,N_4862,N_4861);
and UO_921 (O_921,N_4905,N_4961);
xor UO_922 (O_922,N_4800,N_4887);
and UO_923 (O_923,N_4947,N_4928);
nor UO_924 (O_924,N_4991,N_4931);
nand UO_925 (O_925,N_4975,N_4806);
nand UO_926 (O_926,N_4832,N_4966);
and UO_927 (O_927,N_4968,N_4825);
and UO_928 (O_928,N_4813,N_4879);
xnor UO_929 (O_929,N_4827,N_4838);
nand UO_930 (O_930,N_4866,N_4816);
xnor UO_931 (O_931,N_4851,N_4874);
nand UO_932 (O_932,N_4902,N_4964);
or UO_933 (O_933,N_4898,N_4899);
and UO_934 (O_934,N_4925,N_4860);
or UO_935 (O_935,N_4983,N_4829);
nand UO_936 (O_936,N_4976,N_4981);
and UO_937 (O_937,N_4955,N_4809);
xnor UO_938 (O_938,N_4994,N_4844);
xor UO_939 (O_939,N_4881,N_4963);
nor UO_940 (O_940,N_4838,N_4894);
or UO_941 (O_941,N_4855,N_4928);
xnor UO_942 (O_942,N_4831,N_4948);
xnor UO_943 (O_943,N_4977,N_4857);
nor UO_944 (O_944,N_4947,N_4927);
nor UO_945 (O_945,N_4934,N_4990);
or UO_946 (O_946,N_4903,N_4984);
nor UO_947 (O_947,N_4991,N_4988);
nor UO_948 (O_948,N_4825,N_4857);
xnor UO_949 (O_949,N_4877,N_4844);
nor UO_950 (O_950,N_4882,N_4879);
xor UO_951 (O_951,N_4889,N_4957);
nor UO_952 (O_952,N_4838,N_4932);
or UO_953 (O_953,N_4951,N_4874);
xor UO_954 (O_954,N_4931,N_4854);
nand UO_955 (O_955,N_4984,N_4987);
nor UO_956 (O_956,N_4971,N_4979);
nand UO_957 (O_957,N_4928,N_4808);
or UO_958 (O_958,N_4888,N_4851);
or UO_959 (O_959,N_4896,N_4913);
and UO_960 (O_960,N_4800,N_4853);
nor UO_961 (O_961,N_4885,N_4919);
or UO_962 (O_962,N_4825,N_4905);
xor UO_963 (O_963,N_4945,N_4887);
and UO_964 (O_964,N_4899,N_4904);
nor UO_965 (O_965,N_4860,N_4915);
or UO_966 (O_966,N_4846,N_4931);
xor UO_967 (O_967,N_4845,N_4954);
xnor UO_968 (O_968,N_4828,N_4897);
or UO_969 (O_969,N_4989,N_4818);
nand UO_970 (O_970,N_4938,N_4854);
nand UO_971 (O_971,N_4937,N_4878);
nand UO_972 (O_972,N_4825,N_4969);
and UO_973 (O_973,N_4831,N_4848);
or UO_974 (O_974,N_4807,N_4994);
nand UO_975 (O_975,N_4873,N_4847);
nand UO_976 (O_976,N_4973,N_4812);
nand UO_977 (O_977,N_4852,N_4876);
and UO_978 (O_978,N_4938,N_4920);
and UO_979 (O_979,N_4923,N_4962);
xor UO_980 (O_980,N_4934,N_4835);
nor UO_981 (O_981,N_4954,N_4972);
nand UO_982 (O_982,N_4887,N_4919);
or UO_983 (O_983,N_4981,N_4988);
or UO_984 (O_984,N_4905,N_4926);
xnor UO_985 (O_985,N_4885,N_4954);
or UO_986 (O_986,N_4910,N_4838);
nand UO_987 (O_987,N_4957,N_4999);
or UO_988 (O_988,N_4804,N_4912);
nand UO_989 (O_989,N_4918,N_4972);
or UO_990 (O_990,N_4877,N_4821);
or UO_991 (O_991,N_4871,N_4953);
xnor UO_992 (O_992,N_4958,N_4933);
and UO_993 (O_993,N_4903,N_4857);
or UO_994 (O_994,N_4863,N_4855);
xor UO_995 (O_995,N_4960,N_4837);
xor UO_996 (O_996,N_4817,N_4881);
and UO_997 (O_997,N_4977,N_4820);
or UO_998 (O_998,N_4843,N_4858);
nor UO_999 (O_999,N_4919,N_4963);
endmodule