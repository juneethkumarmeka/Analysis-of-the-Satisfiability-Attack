module basic_750_5000_1000_10_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_281,In_261);
nand U1 (N_1,In_99,In_688);
nand U2 (N_2,In_483,In_622);
xor U3 (N_3,In_153,In_141);
or U4 (N_4,In_524,In_647);
nand U5 (N_5,In_119,In_683);
nand U6 (N_6,In_232,In_749);
nand U7 (N_7,In_746,In_5);
nand U8 (N_8,In_385,In_418);
or U9 (N_9,In_446,In_510);
or U10 (N_10,In_492,In_550);
nand U11 (N_11,In_325,In_745);
nor U12 (N_12,In_727,In_528);
or U13 (N_13,In_149,In_620);
nand U14 (N_14,In_731,In_630);
nor U15 (N_15,In_270,In_225);
nor U16 (N_16,In_458,In_531);
or U17 (N_17,In_125,In_632);
nand U18 (N_18,In_147,In_359);
nand U19 (N_19,In_461,In_354);
and U20 (N_20,In_652,In_552);
nor U21 (N_21,In_157,In_182);
or U22 (N_22,In_172,In_181);
nand U23 (N_23,In_422,In_431);
or U24 (N_24,In_693,In_491);
nor U25 (N_25,In_176,In_519);
or U26 (N_26,In_660,In_584);
or U27 (N_27,In_409,In_52);
or U28 (N_28,In_703,In_668);
or U29 (N_29,In_735,In_152);
nor U30 (N_30,In_242,In_583);
and U31 (N_31,In_407,In_14);
and U32 (N_32,In_223,In_503);
nand U33 (N_33,In_593,In_601);
nand U34 (N_34,In_180,In_608);
nand U35 (N_35,In_406,In_717);
nand U36 (N_36,In_611,In_439);
or U37 (N_37,In_233,In_687);
and U38 (N_38,In_8,In_419);
or U39 (N_39,In_525,In_317);
nor U40 (N_40,In_344,In_291);
and U41 (N_41,In_222,In_135);
nor U42 (N_42,In_37,In_244);
nor U43 (N_43,In_564,In_357);
nand U44 (N_44,In_399,In_424);
nor U45 (N_45,In_81,In_251);
and U46 (N_46,In_643,In_451);
and U47 (N_47,In_22,In_23);
or U48 (N_48,In_656,In_297);
and U49 (N_49,In_477,In_113);
nor U50 (N_50,In_128,In_436);
and U51 (N_51,In_209,In_86);
nor U52 (N_52,In_38,In_274);
nand U53 (N_53,In_576,In_379);
and U54 (N_54,In_537,In_644);
and U55 (N_55,In_376,In_586);
xnor U56 (N_56,In_708,In_732);
and U57 (N_57,In_437,In_423);
or U58 (N_58,In_504,In_741);
or U59 (N_59,In_684,In_729);
nand U60 (N_60,In_674,In_450);
nand U61 (N_61,In_306,In_129);
nor U62 (N_62,In_341,In_547);
nand U63 (N_63,In_410,In_162);
or U64 (N_64,In_736,In_467);
nand U65 (N_65,In_592,In_338);
and U66 (N_66,In_452,In_267);
nor U67 (N_67,In_453,In_594);
nand U68 (N_68,In_441,In_621);
nand U69 (N_69,In_571,In_68);
nand U70 (N_70,In_440,In_569);
or U71 (N_71,In_337,In_105);
and U72 (N_72,In_435,In_529);
nand U73 (N_73,In_645,In_282);
nand U74 (N_74,In_459,In_575);
nor U75 (N_75,In_743,In_744);
or U76 (N_76,In_390,In_533);
nand U77 (N_77,In_397,In_80);
or U78 (N_78,In_130,In_285);
nor U79 (N_79,In_739,In_293);
or U80 (N_80,In_605,In_53);
and U81 (N_81,In_2,In_55);
and U82 (N_82,In_187,In_123);
or U83 (N_83,In_432,In_664);
xor U84 (N_84,In_195,In_208);
nor U85 (N_85,In_616,In_470);
nor U86 (N_86,In_495,In_484);
and U87 (N_87,In_574,In_188);
and U88 (N_88,In_733,In_73);
nand U89 (N_89,In_34,In_370);
and U90 (N_90,In_175,In_50);
nand U91 (N_91,In_694,In_196);
nand U92 (N_92,In_543,In_610);
nand U93 (N_93,In_114,In_500);
xor U94 (N_94,In_604,In_277);
nor U95 (N_95,In_79,In_567);
nand U96 (N_96,In_40,In_725);
nor U97 (N_97,In_460,In_184);
nor U98 (N_98,In_480,In_515);
nor U99 (N_99,In_343,In_220);
nor U100 (N_100,In_454,In_665);
and U101 (N_101,In_348,In_561);
and U102 (N_102,In_512,In_151);
or U103 (N_103,In_597,In_201);
nor U104 (N_104,In_599,In_136);
nor U105 (N_105,In_589,In_32);
nor U106 (N_106,In_497,In_280);
nand U107 (N_107,In_18,In_655);
nor U108 (N_108,In_568,In_143);
or U109 (N_109,In_661,In_144);
or U110 (N_110,In_69,In_26);
nor U111 (N_111,In_702,In_150);
nand U112 (N_112,In_250,In_488);
and U113 (N_113,In_697,In_408);
and U114 (N_114,In_494,In_260);
and U115 (N_115,In_246,In_49);
nand U116 (N_116,In_174,In_64);
or U117 (N_117,In_563,In_737);
and U118 (N_118,In_265,In_95);
nor U119 (N_119,In_168,In_164);
or U120 (N_120,In_65,In_462);
xor U121 (N_121,In_132,In_425);
nor U122 (N_122,In_205,In_216);
or U123 (N_123,In_284,In_332);
nor U124 (N_124,In_724,In_628);
xnor U125 (N_125,In_185,In_46);
nand U126 (N_126,In_641,In_165);
nor U127 (N_127,In_417,In_75);
nand U128 (N_128,In_301,In_485);
and U129 (N_129,In_191,In_318);
and U130 (N_130,In_349,In_221);
nor U131 (N_131,In_612,In_456);
nand U132 (N_132,In_302,In_228);
nand U133 (N_133,In_76,In_699);
nor U134 (N_134,In_25,In_62);
and U135 (N_135,In_723,In_206);
nand U136 (N_136,In_189,In_623);
and U137 (N_137,In_548,In_701);
and U138 (N_138,In_66,In_673);
nand U139 (N_139,In_322,In_468);
and U140 (N_140,In_298,In_371);
or U141 (N_141,In_421,In_101);
nand U142 (N_142,In_3,In_420);
and U143 (N_143,In_229,In_243);
or U144 (N_144,In_326,In_642);
nand U145 (N_145,In_39,In_566);
nor U146 (N_146,In_296,In_190);
or U147 (N_147,In_544,In_77);
nand U148 (N_148,In_139,In_94);
nand U149 (N_149,In_449,In_438);
nor U150 (N_150,In_287,In_514);
or U151 (N_151,In_295,In_20);
and U152 (N_152,In_355,In_670);
and U153 (N_153,In_200,In_249);
and U154 (N_154,In_539,In_672);
or U155 (N_155,In_169,In_442);
or U156 (N_156,In_33,In_678);
nor U157 (N_157,In_648,In_254);
or U158 (N_158,In_177,In_212);
and U159 (N_159,In_559,In_108);
nand U160 (N_160,In_607,In_726);
nand U161 (N_161,In_234,In_6);
nor U162 (N_162,In_689,In_330);
or U163 (N_163,In_363,In_507);
nor U164 (N_164,In_629,In_405);
nand U165 (N_165,In_695,In_478);
xnor U166 (N_166,In_581,In_546);
and U167 (N_167,In_489,In_373);
or U168 (N_168,In_331,In_538);
and U169 (N_169,In_535,In_577);
nor U170 (N_170,In_381,In_82);
nor U171 (N_171,In_17,In_626);
or U172 (N_172,In_372,In_320);
nand U173 (N_173,In_473,In_704);
or U174 (N_174,In_156,In_676);
nand U175 (N_175,In_264,In_327);
or U176 (N_176,In_636,In_598);
or U177 (N_177,In_316,In_553);
and U178 (N_178,In_304,In_572);
and U179 (N_179,In_426,In_4);
nor U180 (N_180,In_573,In_602);
nand U181 (N_181,In_93,In_443);
and U182 (N_182,In_257,In_738);
or U183 (N_183,In_268,In_96);
or U184 (N_184,In_193,In_748);
or U185 (N_185,In_198,In_718);
nor U186 (N_186,In_118,In_12);
xnor U187 (N_187,In_197,In_402);
and U188 (N_188,In_98,In_110);
and U189 (N_189,In_475,In_361);
and U190 (N_190,In_312,In_134);
nor U191 (N_191,In_161,In_633);
nor U192 (N_192,In_562,In_479);
nand U193 (N_193,In_279,In_170);
or U194 (N_194,In_339,In_218);
nand U195 (N_195,In_523,In_269);
or U196 (N_196,In_83,In_166);
nor U197 (N_197,In_625,In_447);
nor U198 (N_198,In_305,In_502);
or U199 (N_199,In_517,In_142);
nor U200 (N_200,In_518,In_207);
and U201 (N_201,In_380,In_398);
or U202 (N_202,In_681,In_72);
nand U203 (N_203,In_155,In_84);
or U204 (N_204,In_482,In_35);
nand U205 (N_205,In_131,In_606);
nor U206 (N_206,In_377,In_682);
or U207 (N_207,In_658,In_530);
nand U208 (N_208,In_685,In_591);
and U209 (N_209,In_618,In_71);
nand U210 (N_210,In_653,In_145);
and U211 (N_211,In_639,In_691);
nand U212 (N_212,In_505,In_255);
and U213 (N_213,In_613,In_627);
nand U214 (N_214,In_651,In_362);
nand U215 (N_215,In_27,In_721);
and U216 (N_216,In_536,In_579);
nand U217 (N_217,In_444,In_711);
and U218 (N_218,In_400,In_13);
nand U219 (N_219,In_412,In_635);
or U220 (N_220,In_382,In_707);
and U221 (N_221,In_252,In_179);
and U222 (N_222,In_516,In_545);
and U223 (N_223,In_464,In_353);
nor U224 (N_224,In_367,In_266);
and U225 (N_225,In_289,In_308);
nand U226 (N_226,In_107,In_522);
and U227 (N_227,In_414,In_219);
or U228 (N_228,In_121,In_556);
and U229 (N_229,In_97,In_47);
or U230 (N_230,In_137,In_677);
nor U231 (N_231,In_342,In_10);
nand U232 (N_232,In_91,In_669);
or U233 (N_233,In_716,In_271);
nand U234 (N_234,In_106,In_347);
nor U235 (N_235,In_712,In_465);
nor U236 (N_236,In_294,In_403);
or U237 (N_237,In_375,In_742);
nor U238 (N_238,In_474,In_650);
nor U239 (N_239,In_321,In_247);
nor U240 (N_240,In_89,In_680);
and U241 (N_241,In_235,In_619);
nor U242 (N_242,In_313,In_56);
nor U243 (N_243,In_74,In_173);
nor U244 (N_244,In_323,In_24);
nor U245 (N_245,In_272,In_15);
nand U246 (N_246,In_63,In_213);
and U247 (N_247,In_138,In_389);
or U248 (N_248,In_51,In_163);
nor U249 (N_249,In_466,In_640);
or U250 (N_250,In_78,In_383);
nand U251 (N_251,In_508,In_541);
or U252 (N_252,In_7,In_44);
and U253 (N_253,In_603,In_19);
nand U254 (N_254,In_273,In_366);
or U255 (N_255,In_369,In_48);
nor U256 (N_256,In_521,In_290);
nor U257 (N_257,In_705,In_117);
and U258 (N_258,In_671,In_226);
nand U259 (N_259,In_388,In_148);
nor U260 (N_260,In_102,In_9);
nor U261 (N_261,In_329,In_551);
or U262 (N_262,In_126,In_360);
nand U263 (N_263,In_248,In_358);
and U264 (N_264,In_600,In_124);
and U265 (N_265,In_31,In_540);
nand U266 (N_266,In_520,In_57);
nor U267 (N_267,In_224,In_311);
and U268 (N_268,In_657,In_85);
or U269 (N_269,In_542,In_340);
and U270 (N_270,In_159,In_580);
or U271 (N_271,In_245,In_30);
or U272 (N_272,In_416,In_328);
and U273 (N_273,In_513,In_236);
nand U274 (N_274,In_570,In_481);
or U275 (N_275,In_713,In_146);
or U276 (N_276,In_710,In_374);
xor U277 (N_277,In_309,In_127);
or U278 (N_278,In_386,In_430);
and U279 (N_279,In_307,In_624);
nand U280 (N_280,In_43,In_217);
and U281 (N_281,In_231,In_549);
or U282 (N_282,In_204,In_214);
nand U283 (N_283,In_532,In_582);
nand U284 (N_284,In_637,In_210);
nand U285 (N_285,In_496,In_486);
nor U286 (N_286,In_300,In_649);
nor U287 (N_287,In_706,In_429);
nand U288 (N_288,In_103,In_122);
and U289 (N_289,In_734,In_45);
nand U290 (N_290,In_472,In_554);
nand U291 (N_291,In_526,In_476);
or U292 (N_292,In_666,In_211);
xor U293 (N_293,In_28,In_654);
and U294 (N_294,In_490,In_116);
nand U295 (N_295,In_275,In_698);
and U296 (N_296,In_587,In_167);
and U297 (N_297,In_42,In_509);
nand U298 (N_298,In_463,In_120);
nor U299 (N_299,In_238,In_368);
or U300 (N_300,In_351,In_747);
and U301 (N_301,In_160,In_378);
or U302 (N_302,In_457,In_720);
and U303 (N_303,In_384,In_511);
nand U304 (N_304,In_183,In_675);
or U305 (N_305,In_719,In_740);
and U306 (N_306,In_667,In_395);
nand U307 (N_307,In_499,In_241);
nor U308 (N_308,In_560,In_614);
and U309 (N_309,In_392,In_227);
and U310 (N_310,In_140,In_286);
nand U311 (N_311,In_192,In_21);
and U312 (N_312,In_61,In_240);
nand U313 (N_313,In_615,In_88);
or U314 (N_314,In_411,In_345);
or U315 (N_315,In_364,In_336);
nor U316 (N_316,In_310,In_262);
nand U317 (N_317,In_324,In_239);
nand U318 (N_318,In_588,In_36);
nor U319 (N_319,In_394,In_534);
nand U320 (N_320,In_29,In_283);
xor U321 (N_321,In_0,In_288);
or U322 (N_322,In_186,In_112);
nand U323 (N_323,In_203,In_413);
or U324 (N_324,In_646,In_595);
or U325 (N_325,In_314,In_11);
xor U326 (N_326,In_278,In_199);
or U327 (N_327,In_299,In_578);
or U328 (N_328,In_178,In_90);
and U329 (N_329,In_100,In_335);
nor U330 (N_330,In_194,In_631);
or U331 (N_331,In_709,In_634);
nand U332 (N_332,In_334,In_433);
or U333 (N_333,In_487,In_202);
or U334 (N_334,In_471,In_714);
nand U335 (N_335,In_154,In_104);
nand U336 (N_336,In_730,In_396);
and U337 (N_337,In_276,In_356);
xnor U338 (N_338,In_158,In_59);
or U339 (N_339,In_230,In_527);
or U340 (N_340,In_319,In_41);
or U341 (N_341,In_253,In_434);
nor U342 (N_342,In_92,In_60);
or U343 (N_343,In_87,In_555);
nand U344 (N_344,In_303,In_346);
xnor U345 (N_345,In_498,In_133);
or U346 (N_346,In_292,In_215);
or U347 (N_347,In_415,In_696);
or U348 (N_348,In_686,In_662);
nand U349 (N_349,In_258,In_111);
and U350 (N_350,In_722,In_67);
nand U351 (N_351,In_263,In_448);
xnor U352 (N_352,In_427,In_333);
nor U353 (N_353,In_506,In_256);
nor U354 (N_354,In_315,In_16);
and U355 (N_355,In_58,In_455);
or U356 (N_356,In_393,In_590);
nand U357 (N_357,In_109,In_609);
and U358 (N_358,In_352,In_585);
nor U359 (N_359,In_171,In_596);
and U360 (N_360,In_679,In_350);
nor U361 (N_361,In_259,In_659);
or U362 (N_362,In_70,In_493);
nor U363 (N_363,In_700,In_663);
nor U364 (N_364,In_715,In_365);
nand U365 (N_365,In_558,In_428);
or U366 (N_366,In_469,In_115);
nor U367 (N_367,In_391,In_728);
and U368 (N_368,In_237,In_404);
or U369 (N_369,In_445,In_565);
and U370 (N_370,In_617,In_1);
nor U371 (N_371,In_638,In_692);
and U372 (N_372,In_690,In_501);
or U373 (N_373,In_54,In_557);
and U374 (N_374,In_387,In_401);
and U375 (N_375,In_746,In_398);
nand U376 (N_376,In_646,In_368);
xnor U377 (N_377,In_684,In_33);
and U378 (N_378,In_387,In_169);
or U379 (N_379,In_15,In_247);
or U380 (N_380,In_609,In_649);
nor U381 (N_381,In_69,In_257);
or U382 (N_382,In_58,In_404);
nand U383 (N_383,In_242,In_251);
nand U384 (N_384,In_128,In_568);
or U385 (N_385,In_128,In_497);
nor U386 (N_386,In_95,In_35);
nor U387 (N_387,In_414,In_746);
nand U388 (N_388,In_228,In_87);
nand U389 (N_389,In_16,In_583);
or U390 (N_390,In_402,In_214);
nor U391 (N_391,In_660,In_140);
or U392 (N_392,In_213,In_233);
and U393 (N_393,In_315,In_40);
and U394 (N_394,In_452,In_265);
nand U395 (N_395,In_249,In_8);
nor U396 (N_396,In_724,In_610);
or U397 (N_397,In_260,In_450);
nand U398 (N_398,In_585,In_47);
and U399 (N_399,In_139,In_165);
nor U400 (N_400,In_91,In_382);
nor U401 (N_401,In_529,In_286);
and U402 (N_402,In_741,In_8);
or U403 (N_403,In_369,In_733);
and U404 (N_404,In_484,In_3);
nor U405 (N_405,In_260,In_82);
nor U406 (N_406,In_206,In_582);
nand U407 (N_407,In_93,In_411);
xnor U408 (N_408,In_523,In_612);
or U409 (N_409,In_193,In_675);
nand U410 (N_410,In_318,In_526);
nor U411 (N_411,In_73,In_116);
nand U412 (N_412,In_513,In_619);
nand U413 (N_413,In_434,In_575);
or U414 (N_414,In_256,In_118);
and U415 (N_415,In_307,In_146);
nand U416 (N_416,In_65,In_471);
nand U417 (N_417,In_503,In_412);
and U418 (N_418,In_49,In_575);
and U419 (N_419,In_411,In_117);
nand U420 (N_420,In_312,In_266);
and U421 (N_421,In_369,In_98);
and U422 (N_422,In_671,In_28);
nand U423 (N_423,In_536,In_480);
nand U424 (N_424,In_670,In_43);
nand U425 (N_425,In_383,In_739);
nor U426 (N_426,In_745,In_266);
nor U427 (N_427,In_221,In_655);
and U428 (N_428,In_463,In_337);
or U429 (N_429,In_645,In_96);
or U430 (N_430,In_44,In_251);
nor U431 (N_431,In_68,In_467);
nor U432 (N_432,In_506,In_387);
nor U433 (N_433,In_301,In_339);
or U434 (N_434,In_279,In_336);
and U435 (N_435,In_745,In_326);
nand U436 (N_436,In_17,In_527);
nand U437 (N_437,In_138,In_524);
or U438 (N_438,In_443,In_364);
nor U439 (N_439,In_517,In_92);
or U440 (N_440,In_719,In_438);
nand U441 (N_441,In_592,In_735);
or U442 (N_442,In_81,In_749);
nor U443 (N_443,In_85,In_124);
and U444 (N_444,In_354,In_675);
nor U445 (N_445,In_108,In_667);
nor U446 (N_446,In_67,In_404);
or U447 (N_447,In_225,In_66);
nand U448 (N_448,In_227,In_22);
nor U449 (N_449,In_381,In_294);
and U450 (N_450,In_79,In_638);
nand U451 (N_451,In_90,In_240);
nand U452 (N_452,In_75,In_392);
and U453 (N_453,In_450,In_105);
nor U454 (N_454,In_78,In_734);
and U455 (N_455,In_469,In_256);
or U456 (N_456,In_643,In_262);
nand U457 (N_457,In_570,In_20);
xnor U458 (N_458,In_555,In_574);
or U459 (N_459,In_166,In_84);
xnor U460 (N_460,In_685,In_157);
and U461 (N_461,In_25,In_222);
and U462 (N_462,In_462,In_464);
or U463 (N_463,In_711,In_5);
or U464 (N_464,In_652,In_554);
or U465 (N_465,In_335,In_478);
nor U466 (N_466,In_235,In_617);
or U467 (N_467,In_726,In_579);
nor U468 (N_468,In_456,In_455);
nand U469 (N_469,In_119,In_607);
nor U470 (N_470,In_389,In_517);
nand U471 (N_471,In_708,In_724);
nand U472 (N_472,In_168,In_292);
nor U473 (N_473,In_611,In_190);
and U474 (N_474,In_120,In_344);
nand U475 (N_475,In_709,In_378);
and U476 (N_476,In_409,In_72);
nand U477 (N_477,In_122,In_578);
nand U478 (N_478,In_250,In_326);
and U479 (N_479,In_725,In_473);
or U480 (N_480,In_62,In_453);
and U481 (N_481,In_501,In_521);
xnor U482 (N_482,In_423,In_639);
nand U483 (N_483,In_531,In_346);
nor U484 (N_484,In_246,In_569);
nor U485 (N_485,In_114,In_74);
nand U486 (N_486,In_3,In_113);
nand U487 (N_487,In_457,In_327);
nand U488 (N_488,In_424,In_14);
and U489 (N_489,In_313,In_398);
nand U490 (N_490,In_692,In_701);
and U491 (N_491,In_234,In_193);
xnor U492 (N_492,In_127,In_558);
nand U493 (N_493,In_264,In_61);
nand U494 (N_494,In_109,In_540);
nor U495 (N_495,In_582,In_142);
and U496 (N_496,In_614,In_237);
nand U497 (N_497,In_740,In_315);
or U498 (N_498,In_2,In_500);
nor U499 (N_499,In_705,In_405);
and U500 (N_500,N_469,N_402);
or U501 (N_501,N_446,N_426);
and U502 (N_502,N_292,N_104);
nor U503 (N_503,N_182,N_202);
nand U504 (N_504,N_78,N_266);
nand U505 (N_505,N_221,N_203);
nor U506 (N_506,N_264,N_488);
or U507 (N_507,N_44,N_484);
and U508 (N_508,N_366,N_495);
or U509 (N_509,N_369,N_85);
and U510 (N_510,N_279,N_443);
or U511 (N_511,N_176,N_476);
or U512 (N_512,N_316,N_435);
nor U513 (N_513,N_454,N_135);
nand U514 (N_514,N_374,N_438);
and U515 (N_515,N_333,N_155);
nor U516 (N_516,N_33,N_385);
or U517 (N_517,N_56,N_413);
nor U518 (N_518,N_7,N_204);
nor U519 (N_519,N_347,N_38);
or U520 (N_520,N_238,N_68);
nand U521 (N_521,N_280,N_231);
nand U522 (N_522,N_340,N_48);
nor U523 (N_523,N_113,N_335);
and U524 (N_524,N_299,N_424);
and U525 (N_525,N_425,N_167);
and U526 (N_526,N_31,N_98);
or U527 (N_527,N_130,N_437);
nor U528 (N_528,N_383,N_143);
nand U529 (N_529,N_122,N_213);
or U530 (N_530,N_233,N_74);
nand U531 (N_531,N_323,N_372);
nand U532 (N_532,N_51,N_99);
nand U533 (N_533,N_62,N_186);
and U534 (N_534,N_380,N_195);
and U535 (N_535,N_132,N_447);
nor U536 (N_536,N_28,N_448);
nand U537 (N_537,N_368,N_246);
nor U538 (N_538,N_36,N_81);
nand U539 (N_539,N_154,N_171);
and U540 (N_540,N_392,N_27);
or U541 (N_541,N_322,N_489);
nor U542 (N_542,N_14,N_309);
or U543 (N_543,N_285,N_190);
or U544 (N_544,N_270,N_459);
or U545 (N_545,N_4,N_326);
nand U546 (N_546,N_139,N_406);
and U547 (N_547,N_445,N_441);
nor U548 (N_548,N_52,N_70);
nor U549 (N_549,N_242,N_403);
nor U550 (N_550,N_145,N_364);
xnor U551 (N_551,N_283,N_228);
nand U552 (N_552,N_183,N_397);
nor U553 (N_553,N_90,N_318);
nand U554 (N_554,N_290,N_388);
xnor U555 (N_555,N_331,N_46);
or U556 (N_556,N_152,N_61);
and U557 (N_557,N_229,N_207);
nor U558 (N_558,N_365,N_158);
or U559 (N_559,N_162,N_470);
and U560 (N_560,N_259,N_352);
and U561 (N_561,N_140,N_430);
and U562 (N_562,N_381,N_219);
nand U563 (N_563,N_327,N_80);
xnor U564 (N_564,N_253,N_197);
or U565 (N_565,N_467,N_357);
xor U566 (N_566,N_465,N_288);
nand U567 (N_567,N_26,N_261);
nand U568 (N_568,N_217,N_421);
nor U569 (N_569,N_225,N_324);
nand U570 (N_570,N_419,N_105);
nand U571 (N_571,N_268,N_308);
and U572 (N_572,N_198,N_54);
and U573 (N_573,N_344,N_147);
nor U574 (N_574,N_449,N_82);
nand U575 (N_575,N_311,N_291);
or U576 (N_576,N_250,N_144);
nor U577 (N_577,N_422,N_452);
nand U578 (N_578,N_245,N_483);
or U579 (N_579,N_84,N_88);
nand U580 (N_580,N_274,N_209);
nor U581 (N_581,N_87,N_96);
nand U582 (N_582,N_386,N_42);
or U583 (N_583,N_119,N_396);
or U584 (N_584,N_110,N_149);
nand U585 (N_585,N_95,N_282);
and U586 (N_586,N_407,N_360);
and U587 (N_587,N_211,N_133);
nor U588 (N_588,N_464,N_196);
xnor U589 (N_589,N_214,N_482);
and U590 (N_590,N_296,N_350);
or U591 (N_591,N_227,N_434);
and U592 (N_592,N_312,N_93);
or U593 (N_593,N_194,N_164);
and U594 (N_594,N_475,N_159);
and U595 (N_595,N_57,N_22);
and U596 (N_596,N_20,N_479);
or U597 (N_597,N_260,N_247);
nor U598 (N_598,N_398,N_305);
or U599 (N_599,N_287,N_16);
and U600 (N_600,N_379,N_265);
nor U601 (N_601,N_237,N_193);
or U602 (N_602,N_497,N_359);
nor U603 (N_603,N_462,N_378);
xor U604 (N_604,N_65,N_492);
or U605 (N_605,N_432,N_375);
nor U606 (N_606,N_477,N_343);
xnor U607 (N_607,N_19,N_86);
nor U608 (N_608,N_83,N_67);
nand U609 (N_609,N_451,N_306);
nor U610 (N_610,N_339,N_478);
nor U611 (N_611,N_123,N_243);
and U612 (N_612,N_136,N_236);
and U613 (N_613,N_49,N_298);
nand U614 (N_614,N_433,N_138);
nand U615 (N_615,N_348,N_240);
or U616 (N_616,N_410,N_373);
or U617 (N_617,N_457,N_116);
xnor U618 (N_618,N_252,N_399);
or U619 (N_619,N_181,N_263);
or U620 (N_620,N_226,N_187);
nand U621 (N_621,N_393,N_401);
or U622 (N_622,N_220,N_415);
or U623 (N_623,N_269,N_480);
and U624 (N_624,N_349,N_455);
or U625 (N_625,N_436,N_428);
and U626 (N_626,N_66,N_112);
and U627 (N_627,N_420,N_1);
and U628 (N_628,N_239,N_60);
nand U629 (N_629,N_45,N_188);
nor U630 (N_630,N_29,N_142);
nand U631 (N_631,N_278,N_168);
or U632 (N_632,N_184,N_126);
or U633 (N_633,N_150,N_458);
xor U634 (N_634,N_101,N_146);
nand U635 (N_635,N_493,N_321);
or U636 (N_636,N_103,N_320);
or U637 (N_637,N_39,N_315);
nor U638 (N_638,N_64,N_248);
or U639 (N_639,N_400,N_10);
and U640 (N_640,N_9,N_92);
nor U641 (N_641,N_473,N_313);
nor U642 (N_642,N_474,N_418);
nand U643 (N_643,N_295,N_409);
or U644 (N_644,N_76,N_153);
nor U645 (N_645,N_199,N_341);
nand U646 (N_646,N_129,N_241);
nor U647 (N_647,N_404,N_351);
and U648 (N_648,N_18,N_300);
or U649 (N_649,N_370,N_25);
nand U650 (N_650,N_463,N_405);
or U651 (N_651,N_390,N_91);
and U652 (N_652,N_151,N_254);
or U653 (N_653,N_262,N_163);
or U654 (N_654,N_487,N_201);
nor U655 (N_655,N_58,N_75);
nand U656 (N_656,N_0,N_102);
or U657 (N_657,N_346,N_40);
nor U658 (N_658,N_354,N_11);
or U659 (N_659,N_361,N_412);
or U660 (N_660,N_485,N_107);
or U661 (N_661,N_89,N_3);
or U662 (N_662,N_496,N_170);
nor U663 (N_663,N_255,N_72);
nand U664 (N_664,N_121,N_2);
nand U665 (N_665,N_294,N_376);
and U666 (N_666,N_442,N_275);
and U667 (N_667,N_134,N_117);
nor U668 (N_668,N_106,N_389);
nor U669 (N_669,N_192,N_115);
nand U670 (N_670,N_391,N_114);
and U671 (N_671,N_328,N_206);
nor U672 (N_672,N_423,N_148);
or U673 (N_673,N_55,N_35);
and U674 (N_674,N_69,N_286);
or U675 (N_675,N_257,N_230);
or U676 (N_676,N_178,N_200);
or U677 (N_677,N_137,N_281);
and U678 (N_678,N_127,N_330);
nor U679 (N_679,N_120,N_32);
and U680 (N_680,N_411,N_125);
and U681 (N_681,N_439,N_358);
nand U682 (N_682,N_314,N_94);
and U683 (N_683,N_332,N_108);
nand U684 (N_684,N_124,N_453);
nand U685 (N_685,N_486,N_218);
nand U686 (N_686,N_244,N_345);
nor U687 (N_687,N_50,N_267);
and U688 (N_688,N_79,N_222);
and U689 (N_689,N_355,N_128);
or U690 (N_690,N_293,N_276);
nor U691 (N_691,N_490,N_481);
and U692 (N_692,N_191,N_173);
nor U693 (N_693,N_249,N_160);
or U694 (N_694,N_161,N_97);
nand U695 (N_695,N_30,N_336);
or U696 (N_696,N_24,N_47);
and U697 (N_697,N_456,N_367);
nor U698 (N_698,N_304,N_356);
or U699 (N_699,N_177,N_258);
nand U700 (N_700,N_429,N_284);
nor U701 (N_701,N_337,N_297);
or U702 (N_702,N_212,N_37);
or U703 (N_703,N_111,N_256);
and U704 (N_704,N_41,N_303);
and U705 (N_705,N_6,N_444);
and U706 (N_706,N_118,N_431);
xnor U707 (N_707,N_17,N_414);
nor U708 (N_708,N_141,N_23);
or U709 (N_709,N_189,N_223);
or U710 (N_710,N_251,N_185);
and U711 (N_711,N_21,N_175);
nand U712 (N_712,N_169,N_174);
xnor U713 (N_713,N_384,N_363);
or U714 (N_714,N_210,N_73);
and U715 (N_715,N_15,N_450);
nand U716 (N_716,N_395,N_59);
nand U717 (N_717,N_13,N_468);
or U718 (N_718,N_382,N_12);
nor U719 (N_719,N_377,N_63);
nand U720 (N_720,N_234,N_338);
nor U721 (N_721,N_71,N_289);
nor U722 (N_722,N_215,N_466);
or U723 (N_723,N_208,N_53);
and U724 (N_724,N_224,N_34);
nand U725 (N_725,N_100,N_491);
and U726 (N_726,N_471,N_408);
and U727 (N_727,N_77,N_394);
or U728 (N_728,N_109,N_371);
nor U729 (N_729,N_277,N_494);
and U730 (N_730,N_272,N_271);
or U731 (N_731,N_319,N_179);
or U732 (N_732,N_131,N_310);
or U733 (N_733,N_180,N_166);
and U734 (N_734,N_325,N_232);
nor U735 (N_735,N_235,N_461);
or U736 (N_736,N_440,N_334);
or U737 (N_737,N_417,N_43);
nor U738 (N_738,N_362,N_156);
nor U739 (N_739,N_472,N_342);
and U740 (N_740,N_353,N_307);
nor U741 (N_741,N_329,N_427);
nand U742 (N_742,N_273,N_157);
nand U743 (N_743,N_205,N_216);
nand U744 (N_744,N_387,N_302);
and U745 (N_745,N_8,N_499);
nand U746 (N_746,N_498,N_460);
or U747 (N_747,N_317,N_5);
nor U748 (N_748,N_165,N_301);
nor U749 (N_749,N_416,N_172);
and U750 (N_750,N_157,N_453);
and U751 (N_751,N_68,N_390);
nor U752 (N_752,N_141,N_10);
nor U753 (N_753,N_96,N_130);
and U754 (N_754,N_246,N_285);
or U755 (N_755,N_275,N_108);
nand U756 (N_756,N_261,N_497);
nor U757 (N_757,N_427,N_203);
nand U758 (N_758,N_314,N_148);
xor U759 (N_759,N_404,N_298);
and U760 (N_760,N_275,N_206);
or U761 (N_761,N_193,N_366);
and U762 (N_762,N_16,N_294);
and U763 (N_763,N_340,N_85);
xnor U764 (N_764,N_357,N_455);
or U765 (N_765,N_343,N_475);
and U766 (N_766,N_119,N_231);
and U767 (N_767,N_185,N_117);
or U768 (N_768,N_408,N_260);
nor U769 (N_769,N_323,N_441);
nor U770 (N_770,N_344,N_341);
and U771 (N_771,N_158,N_458);
nand U772 (N_772,N_276,N_75);
or U773 (N_773,N_499,N_396);
nand U774 (N_774,N_218,N_149);
and U775 (N_775,N_477,N_459);
xnor U776 (N_776,N_6,N_48);
and U777 (N_777,N_130,N_137);
and U778 (N_778,N_111,N_372);
nand U779 (N_779,N_475,N_135);
and U780 (N_780,N_465,N_376);
or U781 (N_781,N_17,N_144);
nand U782 (N_782,N_313,N_9);
nor U783 (N_783,N_471,N_201);
or U784 (N_784,N_104,N_433);
nor U785 (N_785,N_26,N_297);
nand U786 (N_786,N_425,N_461);
nor U787 (N_787,N_139,N_200);
or U788 (N_788,N_25,N_116);
and U789 (N_789,N_268,N_278);
nor U790 (N_790,N_465,N_413);
nor U791 (N_791,N_226,N_181);
nand U792 (N_792,N_499,N_212);
nand U793 (N_793,N_198,N_263);
nor U794 (N_794,N_319,N_439);
nor U795 (N_795,N_92,N_56);
or U796 (N_796,N_40,N_295);
or U797 (N_797,N_52,N_395);
nor U798 (N_798,N_47,N_368);
nand U799 (N_799,N_418,N_288);
or U800 (N_800,N_238,N_83);
or U801 (N_801,N_60,N_261);
nand U802 (N_802,N_76,N_203);
nor U803 (N_803,N_446,N_307);
nor U804 (N_804,N_90,N_180);
or U805 (N_805,N_400,N_80);
or U806 (N_806,N_110,N_131);
nor U807 (N_807,N_226,N_447);
and U808 (N_808,N_180,N_74);
or U809 (N_809,N_352,N_35);
and U810 (N_810,N_154,N_152);
and U811 (N_811,N_30,N_142);
nor U812 (N_812,N_190,N_34);
or U813 (N_813,N_360,N_325);
nand U814 (N_814,N_8,N_70);
and U815 (N_815,N_102,N_147);
or U816 (N_816,N_274,N_394);
and U817 (N_817,N_67,N_227);
or U818 (N_818,N_463,N_496);
nor U819 (N_819,N_138,N_460);
and U820 (N_820,N_32,N_411);
nand U821 (N_821,N_104,N_94);
or U822 (N_822,N_474,N_57);
nand U823 (N_823,N_133,N_273);
nor U824 (N_824,N_290,N_154);
nand U825 (N_825,N_418,N_491);
xnor U826 (N_826,N_308,N_396);
nor U827 (N_827,N_344,N_362);
nand U828 (N_828,N_345,N_469);
nor U829 (N_829,N_359,N_84);
or U830 (N_830,N_110,N_12);
nand U831 (N_831,N_106,N_26);
nor U832 (N_832,N_275,N_427);
and U833 (N_833,N_387,N_425);
and U834 (N_834,N_343,N_322);
or U835 (N_835,N_240,N_2);
or U836 (N_836,N_338,N_284);
and U837 (N_837,N_403,N_205);
nand U838 (N_838,N_485,N_315);
and U839 (N_839,N_237,N_280);
or U840 (N_840,N_307,N_238);
nor U841 (N_841,N_68,N_418);
or U842 (N_842,N_439,N_406);
nand U843 (N_843,N_473,N_327);
nor U844 (N_844,N_224,N_287);
nor U845 (N_845,N_197,N_95);
or U846 (N_846,N_417,N_289);
and U847 (N_847,N_53,N_64);
nor U848 (N_848,N_299,N_276);
or U849 (N_849,N_66,N_474);
and U850 (N_850,N_49,N_492);
nor U851 (N_851,N_238,N_268);
and U852 (N_852,N_175,N_221);
and U853 (N_853,N_34,N_309);
or U854 (N_854,N_313,N_95);
or U855 (N_855,N_178,N_167);
and U856 (N_856,N_129,N_382);
and U857 (N_857,N_271,N_92);
nand U858 (N_858,N_458,N_148);
and U859 (N_859,N_458,N_489);
nor U860 (N_860,N_358,N_476);
nand U861 (N_861,N_223,N_472);
nand U862 (N_862,N_251,N_219);
and U863 (N_863,N_443,N_456);
and U864 (N_864,N_475,N_383);
nor U865 (N_865,N_185,N_190);
nand U866 (N_866,N_420,N_293);
nor U867 (N_867,N_70,N_68);
or U868 (N_868,N_352,N_23);
nor U869 (N_869,N_409,N_276);
nor U870 (N_870,N_219,N_326);
and U871 (N_871,N_270,N_259);
and U872 (N_872,N_220,N_50);
nor U873 (N_873,N_491,N_302);
nand U874 (N_874,N_155,N_4);
nand U875 (N_875,N_405,N_441);
nand U876 (N_876,N_250,N_162);
nor U877 (N_877,N_215,N_312);
and U878 (N_878,N_250,N_108);
or U879 (N_879,N_332,N_232);
and U880 (N_880,N_401,N_151);
and U881 (N_881,N_426,N_44);
nor U882 (N_882,N_59,N_276);
nor U883 (N_883,N_356,N_78);
or U884 (N_884,N_375,N_111);
and U885 (N_885,N_71,N_0);
and U886 (N_886,N_328,N_497);
nor U887 (N_887,N_86,N_347);
and U888 (N_888,N_214,N_292);
nor U889 (N_889,N_282,N_216);
or U890 (N_890,N_49,N_53);
nand U891 (N_891,N_236,N_221);
or U892 (N_892,N_356,N_391);
and U893 (N_893,N_395,N_175);
nand U894 (N_894,N_244,N_231);
nand U895 (N_895,N_474,N_457);
nor U896 (N_896,N_105,N_60);
and U897 (N_897,N_401,N_244);
or U898 (N_898,N_250,N_85);
nand U899 (N_899,N_83,N_369);
and U900 (N_900,N_22,N_9);
or U901 (N_901,N_92,N_337);
and U902 (N_902,N_365,N_346);
nor U903 (N_903,N_326,N_116);
or U904 (N_904,N_309,N_416);
or U905 (N_905,N_300,N_3);
nand U906 (N_906,N_404,N_213);
nor U907 (N_907,N_315,N_351);
nand U908 (N_908,N_117,N_441);
nand U909 (N_909,N_391,N_326);
nor U910 (N_910,N_308,N_191);
nand U911 (N_911,N_196,N_427);
nor U912 (N_912,N_386,N_311);
or U913 (N_913,N_236,N_322);
nor U914 (N_914,N_445,N_166);
nor U915 (N_915,N_18,N_22);
nor U916 (N_916,N_292,N_256);
nand U917 (N_917,N_353,N_410);
xnor U918 (N_918,N_286,N_218);
or U919 (N_919,N_19,N_395);
nand U920 (N_920,N_486,N_232);
or U921 (N_921,N_428,N_447);
or U922 (N_922,N_192,N_50);
nor U923 (N_923,N_225,N_421);
nand U924 (N_924,N_436,N_270);
nor U925 (N_925,N_252,N_142);
nor U926 (N_926,N_499,N_68);
and U927 (N_927,N_137,N_314);
nand U928 (N_928,N_477,N_150);
nor U929 (N_929,N_289,N_32);
and U930 (N_930,N_34,N_11);
xnor U931 (N_931,N_401,N_73);
or U932 (N_932,N_204,N_229);
nand U933 (N_933,N_26,N_241);
nor U934 (N_934,N_483,N_449);
nand U935 (N_935,N_220,N_84);
xnor U936 (N_936,N_372,N_175);
nand U937 (N_937,N_264,N_21);
and U938 (N_938,N_236,N_478);
and U939 (N_939,N_156,N_22);
or U940 (N_940,N_226,N_150);
nor U941 (N_941,N_0,N_61);
nand U942 (N_942,N_346,N_340);
nor U943 (N_943,N_394,N_28);
nand U944 (N_944,N_236,N_474);
nand U945 (N_945,N_452,N_495);
and U946 (N_946,N_72,N_379);
and U947 (N_947,N_153,N_438);
or U948 (N_948,N_337,N_415);
and U949 (N_949,N_404,N_427);
or U950 (N_950,N_1,N_364);
nor U951 (N_951,N_292,N_217);
or U952 (N_952,N_134,N_41);
or U953 (N_953,N_127,N_278);
and U954 (N_954,N_355,N_118);
nand U955 (N_955,N_36,N_485);
and U956 (N_956,N_80,N_191);
nor U957 (N_957,N_252,N_32);
nand U958 (N_958,N_208,N_256);
nand U959 (N_959,N_258,N_243);
and U960 (N_960,N_256,N_439);
and U961 (N_961,N_57,N_174);
nand U962 (N_962,N_5,N_489);
nor U963 (N_963,N_275,N_77);
nand U964 (N_964,N_125,N_33);
or U965 (N_965,N_360,N_168);
and U966 (N_966,N_1,N_226);
and U967 (N_967,N_472,N_44);
and U968 (N_968,N_184,N_104);
and U969 (N_969,N_234,N_57);
and U970 (N_970,N_180,N_193);
nand U971 (N_971,N_319,N_117);
or U972 (N_972,N_7,N_437);
nand U973 (N_973,N_323,N_459);
nand U974 (N_974,N_95,N_356);
nand U975 (N_975,N_499,N_11);
nor U976 (N_976,N_345,N_462);
or U977 (N_977,N_277,N_86);
nor U978 (N_978,N_478,N_435);
or U979 (N_979,N_497,N_229);
nor U980 (N_980,N_282,N_293);
nand U981 (N_981,N_451,N_113);
and U982 (N_982,N_146,N_6);
nand U983 (N_983,N_399,N_331);
nand U984 (N_984,N_113,N_61);
and U985 (N_985,N_256,N_164);
and U986 (N_986,N_412,N_98);
nor U987 (N_987,N_274,N_228);
nor U988 (N_988,N_92,N_357);
nand U989 (N_989,N_186,N_64);
nand U990 (N_990,N_436,N_237);
and U991 (N_991,N_71,N_81);
xor U992 (N_992,N_424,N_243);
nand U993 (N_993,N_154,N_18);
nor U994 (N_994,N_462,N_323);
nand U995 (N_995,N_479,N_9);
or U996 (N_996,N_15,N_288);
nand U997 (N_997,N_186,N_480);
or U998 (N_998,N_331,N_332);
or U999 (N_999,N_33,N_251);
nand U1000 (N_1000,N_675,N_864);
or U1001 (N_1001,N_503,N_670);
nor U1002 (N_1002,N_919,N_827);
or U1003 (N_1003,N_790,N_854);
or U1004 (N_1004,N_597,N_927);
or U1005 (N_1005,N_542,N_617);
and U1006 (N_1006,N_502,N_903);
nor U1007 (N_1007,N_628,N_632);
or U1008 (N_1008,N_876,N_633);
or U1009 (N_1009,N_582,N_557);
nand U1010 (N_1010,N_920,N_507);
or U1011 (N_1011,N_626,N_546);
and U1012 (N_1012,N_567,N_933);
and U1013 (N_1013,N_992,N_783);
and U1014 (N_1014,N_866,N_614);
and U1015 (N_1015,N_640,N_731);
nand U1016 (N_1016,N_777,N_859);
nand U1017 (N_1017,N_797,N_742);
or U1018 (N_1018,N_713,N_774);
and U1019 (N_1019,N_826,N_666);
nor U1020 (N_1020,N_725,N_645);
and U1021 (N_1021,N_709,N_631);
nand U1022 (N_1022,N_805,N_894);
and U1023 (N_1023,N_836,N_701);
or U1024 (N_1024,N_697,N_811);
or U1025 (N_1025,N_668,N_586);
nand U1026 (N_1026,N_729,N_880);
or U1027 (N_1027,N_667,N_948);
and U1028 (N_1028,N_504,N_543);
nand U1029 (N_1029,N_759,N_551);
xnor U1030 (N_1030,N_739,N_559);
xnor U1031 (N_1031,N_893,N_821);
nor U1032 (N_1032,N_657,N_702);
xor U1033 (N_1033,N_999,N_665);
nor U1034 (N_1034,N_878,N_890);
nor U1035 (N_1035,N_850,N_772);
and U1036 (N_1036,N_793,N_712);
or U1037 (N_1037,N_803,N_984);
nor U1038 (N_1038,N_521,N_598);
or U1039 (N_1039,N_509,N_838);
nand U1040 (N_1040,N_929,N_969);
or U1041 (N_1041,N_527,N_804);
nor U1042 (N_1042,N_817,N_660);
nand U1043 (N_1043,N_610,N_724);
nand U1044 (N_1044,N_837,N_500);
nand U1045 (N_1045,N_942,N_681);
nor U1046 (N_1046,N_553,N_647);
and U1047 (N_1047,N_511,N_792);
nand U1048 (N_1048,N_718,N_923);
nor U1049 (N_1049,N_990,N_569);
and U1050 (N_1050,N_965,N_961);
nor U1051 (N_1051,N_762,N_775);
or U1052 (N_1052,N_515,N_734);
nand U1053 (N_1053,N_911,N_771);
nor U1054 (N_1054,N_900,N_525);
nand U1055 (N_1055,N_678,N_841);
nand U1056 (N_1056,N_530,N_889);
and U1057 (N_1057,N_596,N_987);
nor U1058 (N_1058,N_698,N_625);
nand U1059 (N_1059,N_711,N_552);
nand U1060 (N_1060,N_799,N_536);
and U1061 (N_1061,N_523,N_656);
nand U1062 (N_1062,N_595,N_940);
and U1063 (N_1063,N_908,N_727);
xor U1064 (N_1064,N_563,N_917);
or U1065 (N_1065,N_513,N_851);
xor U1066 (N_1066,N_839,N_620);
nand U1067 (N_1067,N_891,N_937);
or U1068 (N_1068,N_907,N_550);
and U1069 (N_1069,N_798,N_829);
or U1070 (N_1070,N_538,N_534);
nand U1071 (N_1071,N_578,N_566);
or U1072 (N_1072,N_636,N_548);
nand U1073 (N_1073,N_561,N_974);
and U1074 (N_1074,N_671,N_868);
or U1075 (N_1075,N_820,N_533);
and U1076 (N_1076,N_761,N_673);
and U1077 (N_1077,N_930,N_787);
nor U1078 (N_1078,N_767,N_539);
or U1079 (N_1079,N_510,N_949);
nor U1080 (N_1080,N_606,N_652);
nand U1081 (N_1081,N_683,N_902);
or U1082 (N_1082,N_649,N_540);
nor U1083 (N_1083,N_863,N_743);
and U1084 (N_1084,N_862,N_782);
and U1085 (N_1085,N_684,N_594);
or U1086 (N_1086,N_730,N_770);
nand U1087 (N_1087,N_603,N_897);
and U1088 (N_1088,N_717,N_815);
nor U1089 (N_1089,N_705,N_519);
xor U1090 (N_1090,N_831,N_576);
and U1091 (N_1091,N_952,N_882);
nor U1092 (N_1092,N_544,N_785);
nor U1093 (N_1093,N_605,N_745);
or U1094 (N_1094,N_840,N_505);
or U1095 (N_1095,N_524,N_806);
or U1096 (N_1096,N_870,N_922);
nand U1097 (N_1097,N_788,N_621);
or U1098 (N_1098,N_537,N_776);
or U1099 (N_1099,N_736,N_912);
or U1100 (N_1100,N_593,N_579);
and U1101 (N_1101,N_791,N_802);
or U1102 (N_1102,N_693,N_562);
nand U1103 (N_1103,N_520,N_737);
nor U1104 (N_1104,N_874,N_583);
nand U1105 (N_1105,N_951,N_813);
or U1106 (N_1106,N_720,N_514);
or U1107 (N_1107,N_612,N_872);
or U1108 (N_1108,N_924,N_662);
nor U1109 (N_1109,N_565,N_516);
nor U1110 (N_1110,N_637,N_950);
nor U1111 (N_1111,N_795,N_573);
or U1112 (N_1112,N_858,N_852);
nor U1113 (N_1113,N_918,N_800);
nand U1114 (N_1114,N_973,N_898);
nor U1115 (N_1115,N_710,N_769);
and U1116 (N_1116,N_825,N_983);
and U1117 (N_1117,N_570,N_564);
xor U1118 (N_1118,N_968,N_856);
nor U1119 (N_1119,N_699,N_959);
nand U1120 (N_1120,N_692,N_602);
nand U1121 (N_1121,N_735,N_715);
or U1122 (N_1122,N_664,N_832);
and U1123 (N_1123,N_744,N_871);
and U1124 (N_1124,N_558,N_843);
and U1125 (N_1125,N_855,N_953);
and U1126 (N_1126,N_574,N_756);
nor U1127 (N_1127,N_997,N_716);
and U1128 (N_1128,N_816,N_584);
and U1129 (N_1129,N_629,N_809);
and U1130 (N_1130,N_758,N_604);
or U1131 (N_1131,N_810,N_989);
nand U1132 (N_1132,N_853,N_752);
and U1133 (N_1133,N_846,N_634);
and U1134 (N_1134,N_661,N_726);
or U1135 (N_1135,N_757,N_676);
nor U1136 (N_1136,N_979,N_695);
nor U1137 (N_1137,N_823,N_580);
and U1138 (N_1138,N_877,N_857);
and U1139 (N_1139,N_687,N_635);
or U1140 (N_1140,N_738,N_679);
or U1141 (N_1141,N_904,N_995);
and U1142 (N_1142,N_963,N_532);
nand U1143 (N_1143,N_977,N_925);
and U1144 (N_1144,N_556,N_590);
and U1145 (N_1145,N_945,N_914);
and U1146 (N_1146,N_936,N_690);
nand U1147 (N_1147,N_910,N_887);
nand U1148 (N_1148,N_921,N_913);
and U1149 (N_1149,N_905,N_512);
and U1150 (N_1150,N_916,N_972);
nor U1151 (N_1151,N_658,N_834);
nand U1152 (N_1152,N_719,N_659);
nand U1153 (N_1153,N_672,N_547);
nand U1154 (N_1154,N_619,N_824);
nand U1155 (N_1155,N_786,N_873);
nand U1156 (N_1156,N_939,N_518);
nand U1157 (N_1157,N_796,N_694);
or U1158 (N_1158,N_967,N_609);
and U1159 (N_1159,N_822,N_935);
or U1160 (N_1160,N_808,N_707);
and U1161 (N_1161,N_998,N_909);
and U1162 (N_1162,N_674,N_528);
nand U1163 (N_1163,N_773,N_971);
nor U1164 (N_1164,N_982,N_646);
and U1165 (N_1165,N_780,N_861);
nor U1166 (N_1166,N_981,N_644);
nor U1167 (N_1167,N_886,N_895);
nand U1168 (N_1168,N_932,N_991);
nand U1169 (N_1169,N_860,N_686);
nor U1170 (N_1170,N_819,N_941);
and U1171 (N_1171,N_615,N_696);
nand U1172 (N_1172,N_733,N_884);
nand U1173 (N_1173,N_529,N_976);
nand U1174 (N_1174,N_571,N_749);
or U1175 (N_1175,N_753,N_526);
or U1176 (N_1176,N_611,N_833);
or U1177 (N_1177,N_766,N_956);
nor U1178 (N_1178,N_642,N_608);
nand U1179 (N_1179,N_944,N_549);
or U1180 (N_1180,N_869,N_708);
and U1181 (N_1181,N_655,N_748);
or U1182 (N_1182,N_568,N_993);
and U1183 (N_1183,N_622,N_835);
nand U1184 (N_1184,N_653,N_560);
or U1185 (N_1185,N_955,N_741);
or U1186 (N_1186,N_740,N_581);
or U1187 (N_1187,N_946,N_669);
and U1188 (N_1188,N_896,N_592);
or U1189 (N_1189,N_732,N_728);
and U1190 (N_1190,N_688,N_865);
or U1191 (N_1191,N_781,N_650);
nor U1192 (N_1192,N_630,N_607);
or U1193 (N_1193,N_814,N_828);
nor U1194 (N_1194,N_721,N_848);
or U1195 (N_1195,N_763,N_881);
or U1196 (N_1196,N_691,N_892);
nand U1197 (N_1197,N_591,N_706);
or U1198 (N_1198,N_750,N_875);
and U1199 (N_1199,N_535,N_879);
nor U1200 (N_1200,N_765,N_980);
or U1201 (N_1201,N_830,N_970);
xor U1202 (N_1202,N_888,N_589);
and U1203 (N_1203,N_682,N_641);
nor U1204 (N_1204,N_943,N_975);
or U1205 (N_1205,N_928,N_760);
nand U1206 (N_1206,N_784,N_677);
and U1207 (N_1207,N_689,N_754);
and U1208 (N_1208,N_957,N_883);
and U1209 (N_1209,N_714,N_747);
or U1210 (N_1210,N_812,N_985);
or U1211 (N_1211,N_585,N_958);
nor U1212 (N_1212,N_599,N_847);
xnor U1213 (N_1213,N_842,N_704);
nor U1214 (N_1214,N_915,N_849);
nand U1215 (N_1215,N_960,N_723);
or U1216 (N_1216,N_555,N_867);
or U1217 (N_1217,N_947,N_700);
or U1218 (N_1218,N_966,N_901);
and U1219 (N_1219,N_541,N_964);
and U1220 (N_1220,N_554,N_994);
nand U1221 (N_1221,N_755,N_601);
and U1222 (N_1222,N_685,N_988);
nor U1223 (N_1223,N_954,N_807);
nand U1224 (N_1224,N_794,N_768);
nand U1225 (N_1225,N_643,N_844);
and U1226 (N_1226,N_764,N_722);
or U1227 (N_1227,N_663,N_986);
nand U1228 (N_1228,N_996,N_680);
and U1229 (N_1229,N_506,N_517);
nand U1230 (N_1230,N_931,N_638);
or U1231 (N_1231,N_651,N_934);
nor U1232 (N_1232,N_613,N_587);
nand U1233 (N_1233,N_845,N_746);
nand U1234 (N_1234,N_926,N_588);
or U1235 (N_1235,N_938,N_623);
nand U1236 (N_1236,N_818,N_899);
nor U1237 (N_1237,N_648,N_789);
and U1238 (N_1238,N_624,N_618);
and U1239 (N_1239,N_531,N_522);
nor U1240 (N_1240,N_703,N_577);
nor U1241 (N_1241,N_906,N_654);
or U1242 (N_1242,N_639,N_545);
nand U1243 (N_1243,N_501,N_508);
nand U1244 (N_1244,N_600,N_575);
and U1245 (N_1245,N_751,N_801);
and U1246 (N_1246,N_778,N_962);
nor U1247 (N_1247,N_779,N_572);
nand U1248 (N_1248,N_978,N_627);
nor U1249 (N_1249,N_616,N_885);
xor U1250 (N_1250,N_823,N_777);
nor U1251 (N_1251,N_580,N_630);
and U1252 (N_1252,N_869,N_526);
or U1253 (N_1253,N_880,N_757);
and U1254 (N_1254,N_712,N_796);
and U1255 (N_1255,N_687,N_571);
or U1256 (N_1256,N_916,N_963);
and U1257 (N_1257,N_687,N_827);
nand U1258 (N_1258,N_736,N_583);
or U1259 (N_1259,N_668,N_530);
nand U1260 (N_1260,N_572,N_909);
and U1261 (N_1261,N_917,N_733);
or U1262 (N_1262,N_760,N_809);
and U1263 (N_1263,N_700,N_801);
and U1264 (N_1264,N_943,N_736);
nand U1265 (N_1265,N_533,N_852);
or U1266 (N_1266,N_936,N_733);
and U1267 (N_1267,N_807,N_699);
and U1268 (N_1268,N_742,N_910);
nor U1269 (N_1269,N_764,N_587);
nand U1270 (N_1270,N_648,N_534);
nor U1271 (N_1271,N_668,N_504);
or U1272 (N_1272,N_728,N_733);
xor U1273 (N_1273,N_562,N_586);
or U1274 (N_1274,N_916,N_781);
and U1275 (N_1275,N_838,N_835);
nand U1276 (N_1276,N_624,N_974);
and U1277 (N_1277,N_740,N_630);
nor U1278 (N_1278,N_785,N_840);
or U1279 (N_1279,N_540,N_520);
nor U1280 (N_1280,N_921,N_974);
or U1281 (N_1281,N_628,N_848);
or U1282 (N_1282,N_728,N_533);
nand U1283 (N_1283,N_925,N_741);
nor U1284 (N_1284,N_579,N_588);
and U1285 (N_1285,N_860,N_583);
and U1286 (N_1286,N_947,N_935);
nand U1287 (N_1287,N_659,N_744);
or U1288 (N_1288,N_955,N_866);
nor U1289 (N_1289,N_845,N_543);
and U1290 (N_1290,N_842,N_629);
or U1291 (N_1291,N_916,N_629);
and U1292 (N_1292,N_879,N_537);
nand U1293 (N_1293,N_951,N_663);
nor U1294 (N_1294,N_549,N_648);
nand U1295 (N_1295,N_781,N_677);
nor U1296 (N_1296,N_988,N_935);
nand U1297 (N_1297,N_642,N_662);
and U1298 (N_1298,N_932,N_874);
nand U1299 (N_1299,N_849,N_889);
and U1300 (N_1300,N_688,N_976);
nand U1301 (N_1301,N_726,N_636);
and U1302 (N_1302,N_872,N_847);
nor U1303 (N_1303,N_882,N_924);
nor U1304 (N_1304,N_934,N_863);
nor U1305 (N_1305,N_629,N_565);
and U1306 (N_1306,N_507,N_575);
nor U1307 (N_1307,N_916,N_637);
or U1308 (N_1308,N_638,N_819);
nand U1309 (N_1309,N_771,N_770);
nor U1310 (N_1310,N_687,N_850);
and U1311 (N_1311,N_696,N_598);
and U1312 (N_1312,N_898,N_855);
xor U1313 (N_1313,N_993,N_583);
nor U1314 (N_1314,N_787,N_947);
and U1315 (N_1315,N_651,N_621);
or U1316 (N_1316,N_816,N_614);
nor U1317 (N_1317,N_817,N_912);
and U1318 (N_1318,N_825,N_720);
nor U1319 (N_1319,N_932,N_516);
or U1320 (N_1320,N_765,N_775);
or U1321 (N_1321,N_833,N_906);
nand U1322 (N_1322,N_910,N_939);
and U1323 (N_1323,N_584,N_969);
or U1324 (N_1324,N_512,N_943);
nor U1325 (N_1325,N_626,N_828);
nand U1326 (N_1326,N_926,N_881);
and U1327 (N_1327,N_545,N_641);
nor U1328 (N_1328,N_892,N_687);
or U1329 (N_1329,N_966,N_894);
nand U1330 (N_1330,N_976,N_709);
and U1331 (N_1331,N_578,N_762);
nand U1332 (N_1332,N_527,N_740);
nor U1333 (N_1333,N_543,N_836);
and U1334 (N_1334,N_729,N_924);
or U1335 (N_1335,N_885,N_647);
nand U1336 (N_1336,N_546,N_694);
or U1337 (N_1337,N_755,N_992);
nand U1338 (N_1338,N_569,N_571);
nor U1339 (N_1339,N_714,N_992);
nand U1340 (N_1340,N_679,N_554);
or U1341 (N_1341,N_837,N_640);
and U1342 (N_1342,N_856,N_764);
and U1343 (N_1343,N_983,N_997);
nand U1344 (N_1344,N_941,N_725);
or U1345 (N_1345,N_701,N_609);
or U1346 (N_1346,N_509,N_553);
nor U1347 (N_1347,N_537,N_733);
nor U1348 (N_1348,N_668,N_523);
and U1349 (N_1349,N_545,N_853);
and U1350 (N_1350,N_616,N_973);
nor U1351 (N_1351,N_946,N_893);
nor U1352 (N_1352,N_720,N_538);
and U1353 (N_1353,N_904,N_770);
nor U1354 (N_1354,N_995,N_600);
or U1355 (N_1355,N_771,N_938);
nand U1356 (N_1356,N_601,N_777);
nor U1357 (N_1357,N_592,N_821);
nand U1358 (N_1358,N_827,N_686);
and U1359 (N_1359,N_521,N_908);
or U1360 (N_1360,N_736,N_825);
nand U1361 (N_1361,N_525,N_606);
nand U1362 (N_1362,N_662,N_775);
and U1363 (N_1363,N_582,N_844);
or U1364 (N_1364,N_533,N_667);
xnor U1365 (N_1365,N_560,N_887);
nand U1366 (N_1366,N_705,N_512);
or U1367 (N_1367,N_674,N_831);
nor U1368 (N_1368,N_999,N_821);
and U1369 (N_1369,N_738,N_616);
nor U1370 (N_1370,N_525,N_732);
or U1371 (N_1371,N_585,N_502);
or U1372 (N_1372,N_953,N_678);
or U1373 (N_1373,N_786,N_813);
or U1374 (N_1374,N_800,N_731);
nor U1375 (N_1375,N_957,N_655);
nand U1376 (N_1376,N_742,N_887);
or U1377 (N_1377,N_662,N_966);
and U1378 (N_1378,N_770,N_607);
nand U1379 (N_1379,N_746,N_747);
or U1380 (N_1380,N_967,N_548);
or U1381 (N_1381,N_921,N_772);
nand U1382 (N_1382,N_891,N_788);
nand U1383 (N_1383,N_842,N_764);
nand U1384 (N_1384,N_560,N_835);
and U1385 (N_1385,N_769,N_978);
and U1386 (N_1386,N_651,N_898);
and U1387 (N_1387,N_544,N_600);
nor U1388 (N_1388,N_772,N_929);
and U1389 (N_1389,N_617,N_870);
and U1390 (N_1390,N_764,N_936);
or U1391 (N_1391,N_845,N_505);
or U1392 (N_1392,N_552,N_940);
or U1393 (N_1393,N_848,N_599);
nor U1394 (N_1394,N_695,N_939);
nor U1395 (N_1395,N_632,N_508);
nand U1396 (N_1396,N_531,N_943);
nand U1397 (N_1397,N_689,N_570);
nand U1398 (N_1398,N_521,N_633);
or U1399 (N_1399,N_791,N_522);
nor U1400 (N_1400,N_952,N_710);
nand U1401 (N_1401,N_926,N_700);
nor U1402 (N_1402,N_647,N_592);
and U1403 (N_1403,N_506,N_855);
and U1404 (N_1404,N_788,N_652);
and U1405 (N_1405,N_813,N_849);
and U1406 (N_1406,N_656,N_920);
nor U1407 (N_1407,N_728,N_843);
or U1408 (N_1408,N_927,N_556);
or U1409 (N_1409,N_834,N_522);
nand U1410 (N_1410,N_702,N_762);
or U1411 (N_1411,N_699,N_792);
nand U1412 (N_1412,N_521,N_935);
and U1413 (N_1413,N_521,N_951);
nor U1414 (N_1414,N_736,N_740);
nor U1415 (N_1415,N_637,N_515);
nand U1416 (N_1416,N_864,N_861);
and U1417 (N_1417,N_709,N_728);
nor U1418 (N_1418,N_775,N_973);
nand U1419 (N_1419,N_616,N_965);
nor U1420 (N_1420,N_899,N_676);
and U1421 (N_1421,N_511,N_851);
or U1422 (N_1422,N_910,N_593);
or U1423 (N_1423,N_503,N_755);
nand U1424 (N_1424,N_694,N_810);
xnor U1425 (N_1425,N_707,N_502);
or U1426 (N_1426,N_757,N_681);
and U1427 (N_1427,N_689,N_852);
and U1428 (N_1428,N_906,N_776);
nor U1429 (N_1429,N_831,N_565);
nand U1430 (N_1430,N_543,N_512);
and U1431 (N_1431,N_914,N_813);
or U1432 (N_1432,N_599,N_653);
and U1433 (N_1433,N_760,N_530);
nand U1434 (N_1434,N_728,N_581);
or U1435 (N_1435,N_609,N_643);
nor U1436 (N_1436,N_580,N_670);
and U1437 (N_1437,N_873,N_664);
nor U1438 (N_1438,N_708,N_770);
or U1439 (N_1439,N_519,N_901);
nand U1440 (N_1440,N_585,N_552);
and U1441 (N_1441,N_508,N_791);
or U1442 (N_1442,N_984,N_741);
nand U1443 (N_1443,N_789,N_807);
nand U1444 (N_1444,N_697,N_976);
and U1445 (N_1445,N_868,N_586);
or U1446 (N_1446,N_672,N_912);
or U1447 (N_1447,N_911,N_604);
nor U1448 (N_1448,N_900,N_519);
or U1449 (N_1449,N_522,N_991);
or U1450 (N_1450,N_982,N_651);
or U1451 (N_1451,N_751,N_507);
nor U1452 (N_1452,N_614,N_780);
nand U1453 (N_1453,N_803,N_733);
and U1454 (N_1454,N_665,N_731);
nand U1455 (N_1455,N_556,N_570);
and U1456 (N_1456,N_979,N_997);
or U1457 (N_1457,N_594,N_839);
or U1458 (N_1458,N_694,N_524);
or U1459 (N_1459,N_928,N_856);
nor U1460 (N_1460,N_630,N_964);
nand U1461 (N_1461,N_893,N_517);
nor U1462 (N_1462,N_670,N_892);
nand U1463 (N_1463,N_956,N_810);
and U1464 (N_1464,N_995,N_735);
and U1465 (N_1465,N_960,N_586);
nor U1466 (N_1466,N_762,N_946);
nor U1467 (N_1467,N_502,N_605);
nand U1468 (N_1468,N_850,N_829);
nand U1469 (N_1469,N_895,N_648);
nand U1470 (N_1470,N_605,N_927);
and U1471 (N_1471,N_933,N_825);
nor U1472 (N_1472,N_993,N_955);
nor U1473 (N_1473,N_706,N_639);
nor U1474 (N_1474,N_827,N_584);
nand U1475 (N_1475,N_742,N_705);
nor U1476 (N_1476,N_700,N_925);
nor U1477 (N_1477,N_627,N_618);
and U1478 (N_1478,N_730,N_851);
and U1479 (N_1479,N_705,N_699);
xor U1480 (N_1480,N_959,N_557);
or U1481 (N_1481,N_787,N_911);
nor U1482 (N_1482,N_707,N_842);
or U1483 (N_1483,N_757,N_532);
or U1484 (N_1484,N_981,N_663);
or U1485 (N_1485,N_843,N_877);
nor U1486 (N_1486,N_975,N_571);
xor U1487 (N_1487,N_658,N_962);
nor U1488 (N_1488,N_958,N_688);
or U1489 (N_1489,N_861,N_815);
nand U1490 (N_1490,N_828,N_915);
and U1491 (N_1491,N_538,N_661);
or U1492 (N_1492,N_825,N_583);
xor U1493 (N_1493,N_725,N_724);
or U1494 (N_1494,N_728,N_965);
nor U1495 (N_1495,N_507,N_543);
or U1496 (N_1496,N_707,N_871);
nand U1497 (N_1497,N_794,N_511);
nand U1498 (N_1498,N_662,N_997);
nor U1499 (N_1499,N_546,N_811);
and U1500 (N_1500,N_1456,N_1187);
nand U1501 (N_1501,N_1258,N_1133);
nor U1502 (N_1502,N_1252,N_1440);
nor U1503 (N_1503,N_1293,N_1011);
nor U1504 (N_1504,N_1354,N_1194);
nand U1505 (N_1505,N_1027,N_1334);
nand U1506 (N_1506,N_1193,N_1461);
nand U1507 (N_1507,N_1409,N_1043);
or U1508 (N_1508,N_1405,N_1146);
and U1509 (N_1509,N_1127,N_1363);
and U1510 (N_1510,N_1198,N_1131);
and U1511 (N_1511,N_1230,N_1094);
or U1512 (N_1512,N_1115,N_1176);
nor U1513 (N_1513,N_1054,N_1220);
nor U1514 (N_1514,N_1271,N_1186);
or U1515 (N_1515,N_1457,N_1147);
nand U1516 (N_1516,N_1154,N_1423);
nand U1517 (N_1517,N_1077,N_1372);
nor U1518 (N_1518,N_1101,N_1025);
nor U1519 (N_1519,N_1199,N_1447);
or U1520 (N_1520,N_1095,N_1426);
and U1521 (N_1521,N_1494,N_1343);
nor U1522 (N_1522,N_1174,N_1404);
nand U1523 (N_1523,N_1317,N_1138);
and U1524 (N_1524,N_1202,N_1316);
nor U1525 (N_1525,N_1029,N_1016);
nor U1526 (N_1526,N_1493,N_1166);
nor U1527 (N_1527,N_1270,N_1120);
or U1528 (N_1528,N_1212,N_1454);
nand U1529 (N_1529,N_1318,N_1192);
nand U1530 (N_1530,N_1032,N_1465);
nor U1531 (N_1531,N_1374,N_1434);
or U1532 (N_1532,N_1282,N_1313);
or U1533 (N_1533,N_1495,N_1468);
nand U1534 (N_1534,N_1414,N_1288);
and U1535 (N_1535,N_1472,N_1099);
nor U1536 (N_1536,N_1368,N_1393);
nand U1537 (N_1537,N_1344,N_1180);
or U1538 (N_1538,N_1328,N_1375);
nor U1539 (N_1539,N_1227,N_1417);
or U1540 (N_1540,N_1234,N_1010);
nor U1541 (N_1541,N_1265,N_1163);
nor U1542 (N_1542,N_1428,N_1200);
nand U1543 (N_1543,N_1251,N_1411);
or U1544 (N_1544,N_1069,N_1416);
and U1545 (N_1545,N_1490,N_1051);
and U1546 (N_1546,N_1152,N_1459);
nand U1547 (N_1547,N_1040,N_1118);
or U1548 (N_1548,N_1184,N_1349);
nand U1549 (N_1549,N_1398,N_1063);
and U1550 (N_1550,N_1320,N_1145);
nand U1551 (N_1551,N_1243,N_1073);
and U1552 (N_1552,N_1306,N_1074);
and U1553 (N_1553,N_1470,N_1276);
nor U1554 (N_1554,N_1137,N_1022);
or U1555 (N_1555,N_1275,N_1272);
nor U1556 (N_1556,N_1453,N_1460);
or U1557 (N_1557,N_1155,N_1356);
nand U1558 (N_1558,N_1290,N_1448);
and U1559 (N_1559,N_1058,N_1250);
nand U1560 (N_1560,N_1452,N_1443);
and U1561 (N_1561,N_1325,N_1371);
or U1562 (N_1562,N_1439,N_1274);
nand U1563 (N_1563,N_1132,N_1231);
or U1564 (N_1564,N_1483,N_1103);
or U1565 (N_1565,N_1098,N_1229);
nor U1566 (N_1566,N_1491,N_1214);
and U1567 (N_1567,N_1064,N_1013);
and U1568 (N_1568,N_1024,N_1340);
or U1569 (N_1569,N_1382,N_1033);
and U1570 (N_1570,N_1464,N_1072);
nand U1571 (N_1571,N_1116,N_1053);
or U1572 (N_1572,N_1246,N_1066);
and U1573 (N_1573,N_1402,N_1266);
and U1574 (N_1574,N_1226,N_1475);
or U1575 (N_1575,N_1353,N_1224);
nor U1576 (N_1576,N_1441,N_1242);
nor U1577 (N_1577,N_1210,N_1042);
nor U1578 (N_1578,N_1397,N_1394);
and U1579 (N_1579,N_1299,N_1237);
xnor U1580 (N_1580,N_1091,N_1020);
nor U1581 (N_1581,N_1062,N_1195);
and U1582 (N_1582,N_1004,N_1373);
nand U1583 (N_1583,N_1264,N_1474);
and U1584 (N_1584,N_1135,N_1143);
nand U1585 (N_1585,N_1451,N_1466);
xnor U1586 (N_1586,N_1435,N_1076);
or U1587 (N_1587,N_1232,N_1188);
nor U1588 (N_1588,N_1412,N_1122);
and U1589 (N_1589,N_1005,N_1018);
or U1590 (N_1590,N_1012,N_1241);
or U1591 (N_1591,N_1129,N_1379);
and U1592 (N_1592,N_1216,N_1097);
and U1593 (N_1593,N_1168,N_1159);
or U1594 (N_1594,N_1158,N_1425);
nor U1595 (N_1595,N_1370,N_1323);
nor U1596 (N_1596,N_1326,N_1236);
nand U1597 (N_1597,N_1486,N_1253);
and U1598 (N_1598,N_1102,N_1294);
nor U1599 (N_1599,N_1481,N_1124);
nor U1600 (N_1600,N_1204,N_1395);
nand U1601 (N_1601,N_1014,N_1437);
nor U1602 (N_1602,N_1151,N_1009);
and U1603 (N_1603,N_1113,N_1307);
and U1604 (N_1604,N_1125,N_1136);
nand U1605 (N_1605,N_1311,N_1107);
xor U1606 (N_1606,N_1348,N_1057);
or U1607 (N_1607,N_1287,N_1477);
and U1608 (N_1608,N_1396,N_1269);
nor U1609 (N_1609,N_1002,N_1105);
nand U1610 (N_1610,N_1182,N_1341);
and U1611 (N_1611,N_1355,N_1028);
or U1612 (N_1612,N_1429,N_1114);
nand U1613 (N_1613,N_1314,N_1181);
and U1614 (N_1614,N_1256,N_1003);
and U1615 (N_1615,N_1338,N_1207);
nand U1616 (N_1616,N_1419,N_1172);
and U1617 (N_1617,N_1342,N_1084);
nand U1618 (N_1618,N_1436,N_1399);
or U1619 (N_1619,N_1498,N_1302);
nor U1620 (N_1620,N_1044,N_1046);
nand U1621 (N_1621,N_1104,N_1281);
or U1622 (N_1622,N_1444,N_1111);
and U1623 (N_1623,N_1403,N_1364);
or U1624 (N_1624,N_1208,N_1268);
nand U1625 (N_1625,N_1427,N_1038);
nor U1626 (N_1626,N_1380,N_1424);
nor U1627 (N_1627,N_1039,N_1119);
nor U1628 (N_1628,N_1463,N_1392);
nor U1629 (N_1629,N_1479,N_1164);
nand U1630 (N_1630,N_1065,N_1415);
nand U1631 (N_1631,N_1171,N_1142);
nor U1632 (N_1632,N_1139,N_1362);
and U1633 (N_1633,N_1408,N_1123);
or U1634 (N_1634,N_1322,N_1418);
nand U1635 (N_1635,N_1450,N_1165);
nand U1636 (N_1636,N_1089,N_1153);
or U1637 (N_1637,N_1496,N_1406);
nand U1638 (N_1638,N_1090,N_1446);
and U1639 (N_1639,N_1420,N_1050);
nor U1640 (N_1640,N_1190,N_1467);
or U1641 (N_1641,N_1140,N_1488);
or U1642 (N_1642,N_1161,N_1036);
and U1643 (N_1643,N_1023,N_1128);
xor U1644 (N_1644,N_1278,N_1352);
xnor U1645 (N_1645,N_1361,N_1345);
nand U1646 (N_1646,N_1480,N_1068);
nor U1647 (N_1647,N_1263,N_1078);
nor U1648 (N_1648,N_1000,N_1254);
and U1649 (N_1649,N_1223,N_1007);
or U1650 (N_1650,N_1286,N_1169);
nand U1651 (N_1651,N_1489,N_1017);
nand U1652 (N_1652,N_1047,N_1482);
nand U1653 (N_1653,N_1346,N_1308);
xnor U1654 (N_1654,N_1121,N_1445);
nor U1655 (N_1655,N_1096,N_1499);
or U1656 (N_1656,N_1359,N_1369);
nand U1657 (N_1657,N_1144,N_1217);
and U1658 (N_1658,N_1331,N_1401);
or U1659 (N_1659,N_1350,N_1430);
nor U1660 (N_1660,N_1283,N_1432);
nand U1661 (N_1661,N_1367,N_1067);
nand U1662 (N_1662,N_1484,N_1366);
nand U1663 (N_1663,N_1389,N_1126);
nand U1664 (N_1664,N_1462,N_1141);
or U1665 (N_1665,N_1244,N_1109);
nor U1666 (N_1666,N_1209,N_1421);
nor U1667 (N_1667,N_1309,N_1431);
nand U1668 (N_1668,N_1222,N_1471);
and U1669 (N_1669,N_1173,N_1228);
and U1670 (N_1670,N_1259,N_1400);
nand U1671 (N_1671,N_1442,N_1075);
nand U1672 (N_1672,N_1458,N_1031);
nor U1673 (N_1673,N_1298,N_1289);
nor U1674 (N_1674,N_1257,N_1061);
and U1675 (N_1675,N_1255,N_1130);
nand U1676 (N_1676,N_1260,N_1150);
nor U1677 (N_1677,N_1279,N_1175);
nand U1678 (N_1678,N_1183,N_1292);
or U1679 (N_1679,N_1413,N_1205);
or U1680 (N_1680,N_1189,N_1178);
nor U1681 (N_1681,N_1315,N_1335);
and U1682 (N_1682,N_1487,N_1324);
nand U1683 (N_1683,N_1052,N_1332);
and U1684 (N_1684,N_1384,N_1358);
nor U1685 (N_1685,N_1034,N_1301);
and U1686 (N_1686,N_1081,N_1006);
xnor U1687 (N_1687,N_1303,N_1245);
nor U1688 (N_1688,N_1455,N_1304);
or U1689 (N_1689,N_1296,N_1378);
and U1690 (N_1690,N_1284,N_1386);
nor U1691 (N_1691,N_1319,N_1196);
or U1692 (N_1692,N_1037,N_1015);
nor U1693 (N_1693,N_1387,N_1410);
and U1694 (N_1694,N_1422,N_1206);
or U1695 (N_1695,N_1170,N_1085);
or U1696 (N_1696,N_1079,N_1238);
or U1697 (N_1697,N_1247,N_1219);
and U1698 (N_1698,N_1218,N_1071);
nor U1699 (N_1699,N_1280,N_1157);
or U1700 (N_1700,N_1221,N_1240);
or U1701 (N_1701,N_1148,N_1385);
or U1702 (N_1702,N_1160,N_1327);
and U1703 (N_1703,N_1473,N_1235);
nand U1704 (N_1704,N_1357,N_1360);
or U1705 (N_1705,N_1197,N_1026);
and U1706 (N_1706,N_1049,N_1381);
and U1707 (N_1707,N_1112,N_1008);
or U1708 (N_1708,N_1351,N_1365);
nand U1709 (N_1709,N_1106,N_1433);
and U1710 (N_1710,N_1225,N_1476);
nand U1711 (N_1711,N_1100,N_1239);
or U1712 (N_1712,N_1438,N_1055);
nand U1713 (N_1713,N_1108,N_1086);
or U1714 (N_1714,N_1201,N_1295);
and U1715 (N_1715,N_1185,N_1117);
or U1716 (N_1716,N_1347,N_1110);
nand U1717 (N_1717,N_1001,N_1300);
nand U1718 (N_1718,N_1449,N_1262);
nor U1719 (N_1719,N_1261,N_1203);
nor U1720 (N_1720,N_1082,N_1291);
or U1721 (N_1721,N_1485,N_1329);
nand U1722 (N_1722,N_1215,N_1233);
or U1723 (N_1723,N_1030,N_1248);
xnor U1724 (N_1724,N_1478,N_1285);
and U1725 (N_1725,N_1407,N_1267);
nand U1726 (N_1726,N_1339,N_1177);
xnor U1727 (N_1727,N_1045,N_1497);
and U1728 (N_1728,N_1162,N_1191);
or U1729 (N_1729,N_1156,N_1333);
or U1730 (N_1730,N_1388,N_1087);
and U1731 (N_1731,N_1019,N_1093);
nand U1732 (N_1732,N_1391,N_1070);
nor U1733 (N_1733,N_1060,N_1083);
or U1734 (N_1734,N_1297,N_1048);
xnor U1735 (N_1735,N_1249,N_1273);
nand U1736 (N_1736,N_1492,N_1337);
nand U1737 (N_1737,N_1310,N_1383);
nand U1738 (N_1738,N_1021,N_1167);
nor U1739 (N_1739,N_1035,N_1088);
and U1740 (N_1740,N_1390,N_1312);
nor U1741 (N_1741,N_1056,N_1134);
or U1742 (N_1742,N_1149,N_1336);
or U1743 (N_1743,N_1376,N_1469);
nand U1744 (N_1744,N_1179,N_1041);
nor U1745 (N_1745,N_1277,N_1377);
and U1746 (N_1746,N_1080,N_1092);
nor U1747 (N_1747,N_1059,N_1211);
xnor U1748 (N_1748,N_1213,N_1305);
nand U1749 (N_1749,N_1321,N_1330);
nand U1750 (N_1750,N_1003,N_1321);
or U1751 (N_1751,N_1456,N_1034);
nor U1752 (N_1752,N_1368,N_1017);
nand U1753 (N_1753,N_1353,N_1436);
nor U1754 (N_1754,N_1355,N_1046);
nand U1755 (N_1755,N_1104,N_1199);
and U1756 (N_1756,N_1004,N_1249);
nand U1757 (N_1757,N_1189,N_1070);
nand U1758 (N_1758,N_1075,N_1088);
xor U1759 (N_1759,N_1061,N_1248);
and U1760 (N_1760,N_1028,N_1044);
or U1761 (N_1761,N_1398,N_1403);
nand U1762 (N_1762,N_1140,N_1253);
nor U1763 (N_1763,N_1333,N_1417);
nand U1764 (N_1764,N_1361,N_1378);
nor U1765 (N_1765,N_1119,N_1252);
xnor U1766 (N_1766,N_1288,N_1194);
or U1767 (N_1767,N_1073,N_1301);
or U1768 (N_1768,N_1178,N_1352);
nor U1769 (N_1769,N_1244,N_1218);
and U1770 (N_1770,N_1309,N_1491);
nor U1771 (N_1771,N_1312,N_1166);
nand U1772 (N_1772,N_1246,N_1195);
xor U1773 (N_1773,N_1016,N_1076);
and U1774 (N_1774,N_1166,N_1395);
and U1775 (N_1775,N_1486,N_1219);
and U1776 (N_1776,N_1271,N_1301);
nand U1777 (N_1777,N_1443,N_1354);
and U1778 (N_1778,N_1353,N_1143);
xnor U1779 (N_1779,N_1072,N_1085);
nand U1780 (N_1780,N_1318,N_1426);
nand U1781 (N_1781,N_1214,N_1035);
nand U1782 (N_1782,N_1231,N_1244);
nor U1783 (N_1783,N_1434,N_1112);
and U1784 (N_1784,N_1466,N_1046);
nand U1785 (N_1785,N_1369,N_1479);
nand U1786 (N_1786,N_1058,N_1343);
nor U1787 (N_1787,N_1476,N_1430);
nand U1788 (N_1788,N_1320,N_1316);
nand U1789 (N_1789,N_1420,N_1483);
nand U1790 (N_1790,N_1007,N_1480);
nor U1791 (N_1791,N_1152,N_1467);
or U1792 (N_1792,N_1178,N_1232);
or U1793 (N_1793,N_1490,N_1377);
or U1794 (N_1794,N_1235,N_1428);
or U1795 (N_1795,N_1218,N_1073);
or U1796 (N_1796,N_1002,N_1209);
or U1797 (N_1797,N_1436,N_1313);
and U1798 (N_1798,N_1405,N_1206);
or U1799 (N_1799,N_1420,N_1041);
nand U1800 (N_1800,N_1387,N_1103);
nor U1801 (N_1801,N_1394,N_1439);
nor U1802 (N_1802,N_1033,N_1371);
and U1803 (N_1803,N_1280,N_1391);
nand U1804 (N_1804,N_1147,N_1320);
nor U1805 (N_1805,N_1003,N_1199);
nor U1806 (N_1806,N_1050,N_1129);
or U1807 (N_1807,N_1223,N_1178);
nand U1808 (N_1808,N_1265,N_1218);
nand U1809 (N_1809,N_1211,N_1217);
and U1810 (N_1810,N_1249,N_1195);
nand U1811 (N_1811,N_1131,N_1448);
nor U1812 (N_1812,N_1368,N_1135);
nand U1813 (N_1813,N_1217,N_1133);
and U1814 (N_1814,N_1413,N_1153);
xor U1815 (N_1815,N_1380,N_1344);
nand U1816 (N_1816,N_1270,N_1474);
and U1817 (N_1817,N_1089,N_1022);
or U1818 (N_1818,N_1308,N_1123);
and U1819 (N_1819,N_1430,N_1066);
nand U1820 (N_1820,N_1036,N_1438);
nor U1821 (N_1821,N_1317,N_1498);
or U1822 (N_1822,N_1064,N_1150);
nand U1823 (N_1823,N_1332,N_1160);
or U1824 (N_1824,N_1499,N_1139);
and U1825 (N_1825,N_1319,N_1073);
nor U1826 (N_1826,N_1359,N_1402);
nor U1827 (N_1827,N_1103,N_1407);
nand U1828 (N_1828,N_1032,N_1249);
or U1829 (N_1829,N_1332,N_1293);
nand U1830 (N_1830,N_1144,N_1405);
and U1831 (N_1831,N_1043,N_1001);
nor U1832 (N_1832,N_1327,N_1139);
xnor U1833 (N_1833,N_1023,N_1399);
and U1834 (N_1834,N_1078,N_1020);
nor U1835 (N_1835,N_1241,N_1152);
nand U1836 (N_1836,N_1163,N_1236);
and U1837 (N_1837,N_1162,N_1073);
or U1838 (N_1838,N_1306,N_1294);
xnor U1839 (N_1839,N_1386,N_1485);
nand U1840 (N_1840,N_1355,N_1200);
nor U1841 (N_1841,N_1247,N_1493);
or U1842 (N_1842,N_1096,N_1373);
or U1843 (N_1843,N_1065,N_1439);
and U1844 (N_1844,N_1261,N_1157);
nor U1845 (N_1845,N_1091,N_1171);
or U1846 (N_1846,N_1295,N_1241);
and U1847 (N_1847,N_1020,N_1416);
nor U1848 (N_1848,N_1434,N_1336);
and U1849 (N_1849,N_1267,N_1170);
and U1850 (N_1850,N_1062,N_1258);
and U1851 (N_1851,N_1099,N_1058);
or U1852 (N_1852,N_1191,N_1021);
xnor U1853 (N_1853,N_1395,N_1340);
and U1854 (N_1854,N_1394,N_1427);
and U1855 (N_1855,N_1117,N_1308);
nor U1856 (N_1856,N_1322,N_1111);
nand U1857 (N_1857,N_1367,N_1397);
or U1858 (N_1858,N_1222,N_1147);
or U1859 (N_1859,N_1262,N_1276);
or U1860 (N_1860,N_1044,N_1397);
nor U1861 (N_1861,N_1376,N_1458);
and U1862 (N_1862,N_1344,N_1017);
nor U1863 (N_1863,N_1224,N_1384);
nand U1864 (N_1864,N_1327,N_1080);
nor U1865 (N_1865,N_1127,N_1364);
or U1866 (N_1866,N_1447,N_1354);
and U1867 (N_1867,N_1010,N_1442);
and U1868 (N_1868,N_1003,N_1276);
nand U1869 (N_1869,N_1455,N_1309);
xor U1870 (N_1870,N_1258,N_1332);
and U1871 (N_1871,N_1180,N_1061);
or U1872 (N_1872,N_1421,N_1148);
and U1873 (N_1873,N_1461,N_1013);
nand U1874 (N_1874,N_1256,N_1355);
nor U1875 (N_1875,N_1444,N_1038);
and U1876 (N_1876,N_1057,N_1231);
and U1877 (N_1877,N_1072,N_1336);
and U1878 (N_1878,N_1391,N_1264);
and U1879 (N_1879,N_1231,N_1160);
nand U1880 (N_1880,N_1286,N_1439);
nor U1881 (N_1881,N_1121,N_1441);
and U1882 (N_1882,N_1474,N_1317);
and U1883 (N_1883,N_1482,N_1271);
and U1884 (N_1884,N_1250,N_1005);
or U1885 (N_1885,N_1077,N_1067);
nand U1886 (N_1886,N_1345,N_1044);
nor U1887 (N_1887,N_1193,N_1104);
nand U1888 (N_1888,N_1373,N_1119);
and U1889 (N_1889,N_1152,N_1402);
nor U1890 (N_1890,N_1105,N_1417);
nand U1891 (N_1891,N_1421,N_1486);
nor U1892 (N_1892,N_1218,N_1275);
and U1893 (N_1893,N_1135,N_1284);
nor U1894 (N_1894,N_1061,N_1050);
nand U1895 (N_1895,N_1177,N_1401);
or U1896 (N_1896,N_1380,N_1270);
nor U1897 (N_1897,N_1196,N_1132);
nand U1898 (N_1898,N_1307,N_1425);
nor U1899 (N_1899,N_1102,N_1486);
or U1900 (N_1900,N_1398,N_1108);
nand U1901 (N_1901,N_1276,N_1180);
nor U1902 (N_1902,N_1090,N_1417);
nor U1903 (N_1903,N_1055,N_1064);
and U1904 (N_1904,N_1365,N_1023);
and U1905 (N_1905,N_1290,N_1263);
xnor U1906 (N_1906,N_1279,N_1075);
nor U1907 (N_1907,N_1280,N_1308);
nand U1908 (N_1908,N_1072,N_1251);
and U1909 (N_1909,N_1359,N_1049);
nand U1910 (N_1910,N_1171,N_1081);
nor U1911 (N_1911,N_1187,N_1005);
nand U1912 (N_1912,N_1220,N_1092);
nor U1913 (N_1913,N_1371,N_1147);
or U1914 (N_1914,N_1210,N_1192);
and U1915 (N_1915,N_1314,N_1116);
xor U1916 (N_1916,N_1455,N_1066);
or U1917 (N_1917,N_1427,N_1365);
or U1918 (N_1918,N_1404,N_1047);
nor U1919 (N_1919,N_1067,N_1153);
or U1920 (N_1920,N_1228,N_1389);
nand U1921 (N_1921,N_1014,N_1204);
nor U1922 (N_1922,N_1179,N_1482);
nor U1923 (N_1923,N_1165,N_1389);
or U1924 (N_1924,N_1393,N_1067);
nand U1925 (N_1925,N_1423,N_1022);
and U1926 (N_1926,N_1050,N_1261);
nand U1927 (N_1927,N_1125,N_1352);
nor U1928 (N_1928,N_1085,N_1122);
nor U1929 (N_1929,N_1414,N_1216);
nor U1930 (N_1930,N_1372,N_1054);
nor U1931 (N_1931,N_1451,N_1065);
or U1932 (N_1932,N_1427,N_1422);
nand U1933 (N_1933,N_1323,N_1132);
and U1934 (N_1934,N_1086,N_1389);
and U1935 (N_1935,N_1322,N_1225);
nor U1936 (N_1936,N_1219,N_1330);
and U1937 (N_1937,N_1008,N_1071);
or U1938 (N_1938,N_1178,N_1032);
or U1939 (N_1939,N_1242,N_1363);
or U1940 (N_1940,N_1067,N_1144);
or U1941 (N_1941,N_1114,N_1402);
and U1942 (N_1942,N_1228,N_1443);
nor U1943 (N_1943,N_1402,N_1471);
or U1944 (N_1944,N_1343,N_1172);
xnor U1945 (N_1945,N_1145,N_1384);
nor U1946 (N_1946,N_1065,N_1318);
xor U1947 (N_1947,N_1128,N_1119);
nor U1948 (N_1948,N_1210,N_1492);
and U1949 (N_1949,N_1414,N_1376);
nand U1950 (N_1950,N_1045,N_1414);
xnor U1951 (N_1951,N_1250,N_1453);
and U1952 (N_1952,N_1311,N_1350);
nor U1953 (N_1953,N_1286,N_1174);
nand U1954 (N_1954,N_1389,N_1444);
or U1955 (N_1955,N_1275,N_1214);
nand U1956 (N_1956,N_1323,N_1180);
and U1957 (N_1957,N_1363,N_1123);
nand U1958 (N_1958,N_1020,N_1113);
nand U1959 (N_1959,N_1158,N_1166);
nor U1960 (N_1960,N_1331,N_1141);
nor U1961 (N_1961,N_1170,N_1496);
or U1962 (N_1962,N_1285,N_1453);
nor U1963 (N_1963,N_1148,N_1302);
nand U1964 (N_1964,N_1148,N_1231);
or U1965 (N_1965,N_1366,N_1066);
nand U1966 (N_1966,N_1137,N_1402);
or U1967 (N_1967,N_1152,N_1047);
and U1968 (N_1968,N_1232,N_1339);
and U1969 (N_1969,N_1019,N_1256);
and U1970 (N_1970,N_1472,N_1093);
and U1971 (N_1971,N_1165,N_1122);
or U1972 (N_1972,N_1238,N_1229);
nor U1973 (N_1973,N_1228,N_1321);
or U1974 (N_1974,N_1316,N_1356);
and U1975 (N_1975,N_1096,N_1252);
nor U1976 (N_1976,N_1211,N_1175);
nand U1977 (N_1977,N_1010,N_1232);
or U1978 (N_1978,N_1073,N_1354);
and U1979 (N_1979,N_1319,N_1356);
nor U1980 (N_1980,N_1490,N_1075);
nor U1981 (N_1981,N_1285,N_1455);
nor U1982 (N_1982,N_1161,N_1244);
and U1983 (N_1983,N_1258,N_1220);
nand U1984 (N_1984,N_1322,N_1059);
nand U1985 (N_1985,N_1352,N_1270);
nand U1986 (N_1986,N_1206,N_1125);
or U1987 (N_1987,N_1434,N_1169);
nor U1988 (N_1988,N_1455,N_1259);
and U1989 (N_1989,N_1317,N_1238);
and U1990 (N_1990,N_1010,N_1132);
nand U1991 (N_1991,N_1228,N_1101);
nor U1992 (N_1992,N_1020,N_1460);
or U1993 (N_1993,N_1418,N_1389);
nor U1994 (N_1994,N_1435,N_1075);
nor U1995 (N_1995,N_1369,N_1457);
nand U1996 (N_1996,N_1373,N_1333);
or U1997 (N_1997,N_1426,N_1328);
and U1998 (N_1998,N_1369,N_1449);
nand U1999 (N_1999,N_1191,N_1370);
and U2000 (N_2000,N_1792,N_1642);
and U2001 (N_2001,N_1538,N_1713);
and U2002 (N_2002,N_1520,N_1552);
nand U2003 (N_2003,N_1803,N_1758);
and U2004 (N_2004,N_1968,N_1998);
nand U2005 (N_2005,N_1536,N_1540);
and U2006 (N_2006,N_1711,N_1869);
or U2007 (N_2007,N_1645,N_1911);
nand U2008 (N_2008,N_1929,N_1509);
nor U2009 (N_2009,N_1507,N_1866);
nand U2010 (N_2010,N_1996,N_1700);
or U2011 (N_2011,N_1639,N_1916);
or U2012 (N_2012,N_1926,N_1731);
or U2013 (N_2013,N_1886,N_1952);
nand U2014 (N_2014,N_1810,N_1832);
and U2015 (N_2015,N_1707,N_1859);
nand U2016 (N_2016,N_1769,N_1892);
nor U2017 (N_2017,N_1880,N_1638);
or U2018 (N_2018,N_1740,N_1785);
and U2019 (N_2019,N_1864,N_1807);
or U2020 (N_2020,N_1871,N_1992);
nor U2021 (N_2021,N_1741,N_1837);
and U2022 (N_2022,N_1826,N_1838);
and U2023 (N_2023,N_1857,N_1574);
nor U2024 (N_2024,N_1526,N_1767);
and U2025 (N_2025,N_1945,N_1979);
or U2026 (N_2026,N_1861,N_1908);
xor U2027 (N_2027,N_1681,N_1891);
nand U2028 (N_2028,N_1894,N_1919);
nor U2029 (N_2029,N_1946,N_1999);
nor U2030 (N_2030,N_1889,N_1882);
or U2031 (N_2031,N_1963,N_1783);
nor U2032 (N_2032,N_1896,N_1967);
or U2033 (N_2033,N_1955,N_1565);
or U2034 (N_2034,N_1531,N_1523);
or U2035 (N_2035,N_1879,N_1953);
nand U2036 (N_2036,N_1609,N_1544);
nor U2037 (N_2037,N_1974,N_1885);
and U2038 (N_2038,N_1678,N_1559);
nand U2039 (N_2039,N_1931,N_1875);
nor U2040 (N_2040,N_1688,N_1725);
or U2041 (N_2041,N_1641,N_1628);
nor U2042 (N_2042,N_1934,N_1671);
nor U2043 (N_2043,N_1790,N_1691);
and U2044 (N_2044,N_1787,N_1561);
nor U2045 (N_2045,N_1611,N_1663);
or U2046 (N_2046,N_1510,N_1951);
and U2047 (N_2047,N_1578,N_1789);
nand U2048 (N_2048,N_1560,N_1813);
nand U2049 (N_2049,N_1853,N_1768);
or U2050 (N_2050,N_1545,N_1847);
and U2051 (N_2051,N_1918,N_1577);
nand U2052 (N_2052,N_1772,N_1774);
nand U2053 (N_2053,N_1851,N_1806);
nor U2054 (N_2054,N_1930,N_1612);
or U2055 (N_2055,N_1957,N_1596);
or U2056 (N_2056,N_1654,N_1925);
nor U2057 (N_2057,N_1562,N_1670);
or U2058 (N_2058,N_1901,N_1786);
nor U2059 (N_2059,N_1634,N_1595);
nor U2060 (N_2060,N_1710,N_1695);
or U2061 (N_2061,N_1883,N_1662);
nand U2062 (N_2062,N_1555,N_1960);
nand U2063 (N_2063,N_1550,N_1677);
nand U2064 (N_2064,N_1912,N_1680);
nor U2065 (N_2065,N_1948,N_1718);
or U2066 (N_2066,N_1805,N_1760);
and U2067 (N_2067,N_1753,N_1557);
nand U2068 (N_2068,N_1860,N_1547);
and U2069 (N_2069,N_1701,N_1682);
and U2070 (N_2070,N_1702,N_1633);
nor U2071 (N_2071,N_1610,N_1933);
nor U2072 (N_2072,N_1714,N_1534);
nand U2073 (N_2073,N_1679,N_1971);
nor U2074 (N_2074,N_1759,N_1924);
nor U2075 (N_2075,N_1820,N_1516);
and U2076 (N_2076,N_1721,N_1719);
and U2077 (N_2077,N_1533,N_1747);
nand U2078 (N_2078,N_1553,N_1615);
nor U2079 (N_2079,N_1877,N_1692);
nor U2080 (N_2080,N_1737,N_1618);
and U2081 (N_2081,N_1500,N_1842);
or U2082 (N_2082,N_1804,N_1524);
and U2083 (N_2083,N_1909,N_1907);
nor U2084 (N_2084,N_1636,N_1729);
nand U2085 (N_2085,N_1821,N_1938);
or U2086 (N_2086,N_1809,N_1897);
or U2087 (N_2087,N_1850,N_1503);
nor U2088 (N_2088,N_1839,N_1674);
and U2089 (N_2089,N_1863,N_1716);
nor U2090 (N_2090,N_1608,N_1522);
and U2091 (N_2091,N_1604,N_1870);
nand U2092 (N_2092,N_1512,N_1818);
or U2093 (N_2093,N_1727,N_1514);
nor U2094 (N_2094,N_1601,N_1862);
and U2095 (N_2095,N_1980,N_1582);
nor U2096 (N_2096,N_1749,N_1685);
or U2097 (N_2097,N_1872,N_1920);
and U2098 (N_2098,N_1653,N_1505);
or U2099 (N_2099,N_1732,N_1613);
nor U2100 (N_2100,N_1959,N_1981);
nor U2101 (N_2101,N_1917,N_1566);
or U2102 (N_2102,N_1928,N_1841);
or U2103 (N_2103,N_1969,N_1833);
nand U2104 (N_2104,N_1942,N_1583);
and U2105 (N_2105,N_1873,N_1508);
and U2106 (N_2106,N_1814,N_1984);
and U2107 (N_2107,N_1705,N_1935);
nor U2108 (N_2108,N_1812,N_1905);
and U2109 (N_2109,N_1698,N_1899);
nor U2110 (N_2110,N_1811,N_1782);
nor U2111 (N_2111,N_1976,N_1659);
or U2112 (N_2112,N_1651,N_1644);
nand U2113 (N_2113,N_1586,N_1537);
xor U2114 (N_2114,N_1655,N_1669);
and U2115 (N_2115,N_1964,N_1827);
and U2116 (N_2116,N_1699,N_1855);
and U2117 (N_2117,N_1858,N_1735);
or U2118 (N_2118,N_1745,N_1791);
and U2119 (N_2119,N_1902,N_1535);
or U2120 (N_2120,N_1530,N_1637);
and U2121 (N_2121,N_1541,N_1779);
nand U2122 (N_2122,N_1888,N_1546);
nand U2123 (N_2123,N_1597,N_1756);
or U2124 (N_2124,N_1708,N_1567);
nor U2125 (N_2125,N_1693,N_1965);
or U2126 (N_2126,N_1724,N_1937);
or U2127 (N_2127,N_1843,N_1835);
nor U2128 (N_2128,N_1656,N_1985);
or U2129 (N_2129,N_1978,N_1944);
nor U2130 (N_2130,N_1631,N_1650);
or U2131 (N_2131,N_1730,N_1706);
or U2132 (N_2132,N_1624,N_1598);
or U2133 (N_2133,N_1778,N_1748);
nor U2134 (N_2134,N_1599,N_1584);
and U2135 (N_2135,N_1617,N_1525);
nand U2136 (N_2136,N_1548,N_1606);
nor U2137 (N_2137,N_1982,N_1966);
or U2138 (N_2138,N_1846,N_1519);
nand U2139 (N_2139,N_1836,N_1751);
and U2140 (N_2140,N_1961,N_1777);
and U2141 (N_2141,N_1607,N_1922);
or U2142 (N_2142,N_1672,N_1904);
or U2143 (N_2143,N_1580,N_1781);
nor U2144 (N_2144,N_1709,N_1585);
and U2145 (N_2145,N_1986,N_1893);
nand U2146 (N_2146,N_1549,N_1646);
nor U2147 (N_2147,N_1775,N_1589);
nor U2148 (N_2148,N_1627,N_1848);
nor U2149 (N_2149,N_1868,N_1773);
nand U2150 (N_2150,N_1600,N_1554);
nor U2151 (N_2151,N_1587,N_1958);
nand U2152 (N_2152,N_1903,N_1849);
nand U2153 (N_2153,N_1954,N_1649);
nor U2154 (N_2154,N_1532,N_1990);
nand U2155 (N_2155,N_1906,N_1518);
or U2156 (N_2156,N_1703,N_1665);
and U2157 (N_2157,N_1771,N_1723);
and U2158 (N_2158,N_1630,N_1932);
or U2159 (N_2159,N_1995,N_1801);
and U2160 (N_2160,N_1570,N_1579);
nand U2161 (N_2161,N_1590,N_1823);
or U2162 (N_2162,N_1513,N_1874);
nand U2163 (N_2163,N_1983,N_1854);
or U2164 (N_2164,N_1720,N_1742);
nand U2165 (N_2165,N_1593,N_1660);
and U2166 (N_2166,N_1923,N_1991);
or U2167 (N_2167,N_1939,N_1506);
nor U2168 (N_2168,N_1666,N_1687);
nor U2169 (N_2169,N_1797,N_1798);
nor U2170 (N_2170,N_1591,N_1844);
nor U2171 (N_2171,N_1558,N_1616);
nand U2172 (N_2172,N_1770,N_1800);
nand U2173 (N_2173,N_1876,N_1936);
and U2174 (N_2174,N_1815,N_1543);
and U2175 (N_2175,N_1704,N_1575);
or U2176 (N_2176,N_1764,N_1648);
nor U2177 (N_2177,N_1563,N_1970);
nand U2178 (N_2178,N_1673,N_1890);
and U2179 (N_2179,N_1867,N_1539);
nor U2180 (N_2180,N_1752,N_1840);
nand U2181 (N_2181,N_1750,N_1602);
nand U2182 (N_2182,N_1620,N_1761);
or U2183 (N_2183,N_1675,N_1822);
or U2184 (N_2184,N_1527,N_1757);
nand U2185 (N_2185,N_1972,N_1776);
or U2186 (N_2186,N_1551,N_1845);
nand U2187 (N_2187,N_1898,N_1728);
and U2188 (N_2188,N_1502,N_1973);
xor U2189 (N_2189,N_1943,N_1743);
and U2190 (N_2190,N_1799,N_1564);
nor U2191 (N_2191,N_1795,N_1796);
nor U2192 (N_2192,N_1556,N_1825);
or U2193 (N_2193,N_1994,N_1542);
and U2194 (N_2194,N_1856,N_1528);
nor U2195 (N_2195,N_1573,N_1975);
nor U2196 (N_2196,N_1622,N_1726);
nor U2197 (N_2197,N_1588,N_1915);
nand U2198 (N_2198,N_1689,N_1658);
nand U2199 (N_2199,N_1824,N_1632);
nand U2200 (N_2200,N_1712,N_1619);
nor U2201 (N_2201,N_1571,N_1722);
or U2202 (N_2202,N_1921,N_1834);
nor U2203 (N_2203,N_1738,N_1762);
or U2204 (N_2204,N_1829,N_1950);
and U2205 (N_2205,N_1988,N_1676);
nand U2206 (N_2206,N_1683,N_1736);
nand U2207 (N_2207,N_1664,N_1746);
nor U2208 (N_2208,N_1569,N_1755);
or U2209 (N_2209,N_1517,N_1865);
nor U2210 (N_2210,N_1754,N_1733);
nand U2211 (N_2211,N_1734,N_1852);
and U2212 (N_2212,N_1657,N_1793);
or U2213 (N_2213,N_1993,N_1572);
nand U2214 (N_2214,N_1521,N_1763);
nor U2215 (N_2215,N_1884,N_1940);
nand U2216 (N_2216,N_1977,N_1887);
nor U2217 (N_2217,N_1511,N_1690);
or U2218 (N_2218,N_1949,N_1501);
nand U2219 (N_2219,N_1684,N_1717);
or U2220 (N_2220,N_1962,N_1640);
or U2221 (N_2221,N_1997,N_1614);
or U2222 (N_2222,N_1794,N_1603);
nand U2223 (N_2223,N_1581,N_1780);
nand U2224 (N_2224,N_1643,N_1529);
nand U2225 (N_2225,N_1788,N_1895);
nand U2226 (N_2226,N_1819,N_1697);
nand U2227 (N_2227,N_1830,N_1576);
nand U2228 (N_2228,N_1802,N_1647);
nor U2229 (N_2229,N_1621,N_1784);
or U2230 (N_2230,N_1765,N_1766);
nor U2231 (N_2231,N_1625,N_1817);
nand U2232 (N_2232,N_1605,N_1914);
and U2233 (N_2233,N_1947,N_1900);
nor U2234 (N_2234,N_1989,N_1927);
nand U2235 (N_2235,N_1635,N_1878);
nor U2236 (N_2236,N_1696,N_1831);
and U2237 (N_2237,N_1594,N_1661);
and U2238 (N_2238,N_1808,N_1629);
nand U2239 (N_2239,N_1515,N_1816);
and U2240 (N_2240,N_1686,N_1739);
and U2241 (N_2241,N_1881,N_1623);
nand U2242 (N_2242,N_1694,N_1956);
nand U2243 (N_2243,N_1913,N_1592);
or U2244 (N_2244,N_1568,N_1828);
or U2245 (N_2245,N_1504,N_1715);
nand U2246 (N_2246,N_1910,N_1652);
nor U2247 (N_2247,N_1987,N_1668);
or U2248 (N_2248,N_1626,N_1667);
nor U2249 (N_2249,N_1744,N_1941);
nor U2250 (N_2250,N_1965,N_1614);
and U2251 (N_2251,N_1917,N_1637);
or U2252 (N_2252,N_1605,N_1961);
or U2253 (N_2253,N_1551,N_1682);
nand U2254 (N_2254,N_1641,N_1599);
nand U2255 (N_2255,N_1647,N_1991);
nor U2256 (N_2256,N_1582,N_1763);
or U2257 (N_2257,N_1944,N_1911);
or U2258 (N_2258,N_1839,N_1961);
or U2259 (N_2259,N_1683,N_1598);
nand U2260 (N_2260,N_1909,N_1634);
and U2261 (N_2261,N_1914,N_1643);
or U2262 (N_2262,N_1910,N_1965);
nand U2263 (N_2263,N_1716,N_1814);
nand U2264 (N_2264,N_1744,N_1806);
nand U2265 (N_2265,N_1768,N_1744);
nor U2266 (N_2266,N_1827,N_1916);
or U2267 (N_2267,N_1634,N_1626);
nor U2268 (N_2268,N_1730,N_1865);
and U2269 (N_2269,N_1636,N_1611);
nand U2270 (N_2270,N_1579,N_1506);
and U2271 (N_2271,N_1554,N_1969);
and U2272 (N_2272,N_1786,N_1920);
or U2273 (N_2273,N_1673,N_1814);
or U2274 (N_2274,N_1822,N_1986);
nor U2275 (N_2275,N_1989,N_1979);
and U2276 (N_2276,N_1768,N_1696);
nor U2277 (N_2277,N_1714,N_1987);
nor U2278 (N_2278,N_1542,N_1673);
xnor U2279 (N_2279,N_1876,N_1787);
nand U2280 (N_2280,N_1723,N_1517);
nand U2281 (N_2281,N_1614,N_1546);
nor U2282 (N_2282,N_1609,N_1718);
or U2283 (N_2283,N_1889,N_1537);
nand U2284 (N_2284,N_1630,N_1652);
nand U2285 (N_2285,N_1507,N_1712);
nand U2286 (N_2286,N_1669,N_1757);
or U2287 (N_2287,N_1925,N_1960);
or U2288 (N_2288,N_1685,N_1934);
or U2289 (N_2289,N_1761,N_1615);
and U2290 (N_2290,N_1988,N_1531);
and U2291 (N_2291,N_1949,N_1672);
nand U2292 (N_2292,N_1783,N_1641);
nand U2293 (N_2293,N_1639,N_1881);
and U2294 (N_2294,N_1677,N_1552);
nor U2295 (N_2295,N_1565,N_1847);
or U2296 (N_2296,N_1642,N_1851);
or U2297 (N_2297,N_1736,N_1535);
or U2298 (N_2298,N_1761,N_1924);
nor U2299 (N_2299,N_1771,N_1796);
nand U2300 (N_2300,N_1551,N_1958);
nand U2301 (N_2301,N_1805,N_1546);
or U2302 (N_2302,N_1780,N_1754);
or U2303 (N_2303,N_1887,N_1622);
or U2304 (N_2304,N_1770,N_1844);
and U2305 (N_2305,N_1943,N_1907);
nor U2306 (N_2306,N_1955,N_1835);
nand U2307 (N_2307,N_1759,N_1846);
and U2308 (N_2308,N_1878,N_1859);
nand U2309 (N_2309,N_1655,N_1590);
nor U2310 (N_2310,N_1508,N_1847);
and U2311 (N_2311,N_1663,N_1694);
nor U2312 (N_2312,N_1922,N_1621);
or U2313 (N_2313,N_1583,N_1789);
nand U2314 (N_2314,N_1776,N_1714);
nor U2315 (N_2315,N_1611,N_1648);
nor U2316 (N_2316,N_1602,N_1696);
nand U2317 (N_2317,N_1719,N_1532);
nand U2318 (N_2318,N_1510,N_1965);
or U2319 (N_2319,N_1573,N_1645);
and U2320 (N_2320,N_1897,N_1668);
or U2321 (N_2321,N_1610,N_1576);
nand U2322 (N_2322,N_1799,N_1751);
or U2323 (N_2323,N_1899,N_1951);
nor U2324 (N_2324,N_1967,N_1924);
or U2325 (N_2325,N_1507,N_1501);
or U2326 (N_2326,N_1890,N_1629);
nand U2327 (N_2327,N_1790,N_1905);
or U2328 (N_2328,N_1810,N_1557);
nor U2329 (N_2329,N_1781,N_1656);
nand U2330 (N_2330,N_1754,N_1658);
or U2331 (N_2331,N_1655,N_1707);
or U2332 (N_2332,N_1565,N_1547);
nand U2333 (N_2333,N_1998,N_1881);
and U2334 (N_2334,N_1918,N_1743);
nand U2335 (N_2335,N_1938,N_1901);
xor U2336 (N_2336,N_1880,N_1965);
and U2337 (N_2337,N_1916,N_1655);
and U2338 (N_2338,N_1835,N_1750);
nor U2339 (N_2339,N_1704,N_1634);
and U2340 (N_2340,N_1529,N_1577);
nor U2341 (N_2341,N_1648,N_1838);
and U2342 (N_2342,N_1630,N_1612);
and U2343 (N_2343,N_1938,N_1971);
nor U2344 (N_2344,N_1839,N_1702);
nand U2345 (N_2345,N_1626,N_1961);
nand U2346 (N_2346,N_1794,N_1890);
nand U2347 (N_2347,N_1738,N_1966);
and U2348 (N_2348,N_1910,N_1781);
and U2349 (N_2349,N_1812,N_1680);
nor U2350 (N_2350,N_1669,N_1699);
nand U2351 (N_2351,N_1960,N_1613);
nor U2352 (N_2352,N_1657,N_1953);
or U2353 (N_2353,N_1815,N_1552);
and U2354 (N_2354,N_1682,N_1877);
nand U2355 (N_2355,N_1814,N_1701);
nand U2356 (N_2356,N_1920,N_1772);
or U2357 (N_2357,N_1614,N_1754);
and U2358 (N_2358,N_1545,N_1778);
and U2359 (N_2359,N_1665,N_1910);
nor U2360 (N_2360,N_1836,N_1728);
or U2361 (N_2361,N_1705,N_1511);
or U2362 (N_2362,N_1626,N_1594);
or U2363 (N_2363,N_1681,N_1865);
nand U2364 (N_2364,N_1535,N_1817);
or U2365 (N_2365,N_1572,N_1939);
nor U2366 (N_2366,N_1527,N_1979);
nand U2367 (N_2367,N_1936,N_1698);
nor U2368 (N_2368,N_1677,N_1544);
nor U2369 (N_2369,N_1667,N_1649);
xnor U2370 (N_2370,N_1976,N_1536);
nand U2371 (N_2371,N_1835,N_1805);
nand U2372 (N_2372,N_1988,N_1579);
and U2373 (N_2373,N_1537,N_1553);
nand U2374 (N_2374,N_1737,N_1543);
nand U2375 (N_2375,N_1777,N_1584);
or U2376 (N_2376,N_1947,N_1697);
nor U2377 (N_2377,N_1828,N_1508);
xor U2378 (N_2378,N_1671,N_1931);
nand U2379 (N_2379,N_1618,N_1690);
and U2380 (N_2380,N_1834,N_1604);
or U2381 (N_2381,N_1744,N_1903);
nor U2382 (N_2382,N_1912,N_1896);
nand U2383 (N_2383,N_1634,N_1682);
nor U2384 (N_2384,N_1708,N_1718);
xnor U2385 (N_2385,N_1594,N_1513);
or U2386 (N_2386,N_1662,N_1824);
nor U2387 (N_2387,N_1597,N_1718);
or U2388 (N_2388,N_1699,N_1574);
or U2389 (N_2389,N_1992,N_1557);
and U2390 (N_2390,N_1674,N_1847);
nand U2391 (N_2391,N_1857,N_1598);
nand U2392 (N_2392,N_1994,N_1736);
xnor U2393 (N_2393,N_1849,N_1652);
nor U2394 (N_2394,N_1634,N_1644);
and U2395 (N_2395,N_1666,N_1522);
or U2396 (N_2396,N_1943,N_1991);
or U2397 (N_2397,N_1509,N_1578);
xnor U2398 (N_2398,N_1603,N_1720);
xor U2399 (N_2399,N_1741,N_1830);
or U2400 (N_2400,N_1653,N_1557);
nand U2401 (N_2401,N_1892,N_1832);
nand U2402 (N_2402,N_1863,N_1859);
and U2403 (N_2403,N_1723,N_1694);
and U2404 (N_2404,N_1937,N_1595);
nand U2405 (N_2405,N_1865,N_1530);
nand U2406 (N_2406,N_1817,N_1770);
xor U2407 (N_2407,N_1939,N_1916);
nand U2408 (N_2408,N_1693,N_1782);
nor U2409 (N_2409,N_1979,N_1774);
or U2410 (N_2410,N_1817,N_1772);
or U2411 (N_2411,N_1894,N_1946);
or U2412 (N_2412,N_1626,N_1951);
nor U2413 (N_2413,N_1631,N_1694);
nand U2414 (N_2414,N_1504,N_1626);
and U2415 (N_2415,N_1671,N_1707);
nand U2416 (N_2416,N_1798,N_1917);
nand U2417 (N_2417,N_1680,N_1975);
and U2418 (N_2418,N_1872,N_1806);
and U2419 (N_2419,N_1504,N_1851);
or U2420 (N_2420,N_1794,N_1951);
or U2421 (N_2421,N_1710,N_1886);
and U2422 (N_2422,N_1636,N_1634);
nand U2423 (N_2423,N_1807,N_1776);
nand U2424 (N_2424,N_1592,N_1898);
or U2425 (N_2425,N_1973,N_1869);
nor U2426 (N_2426,N_1863,N_1700);
nand U2427 (N_2427,N_1871,N_1851);
xor U2428 (N_2428,N_1752,N_1722);
nor U2429 (N_2429,N_1782,N_1643);
nor U2430 (N_2430,N_1935,N_1647);
nor U2431 (N_2431,N_1597,N_1986);
nor U2432 (N_2432,N_1888,N_1835);
or U2433 (N_2433,N_1551,N_1967);
and U2434 (N_2434,N_1647,N_1849);
nor U2435 (N_2435,N_1643,N_1693);
and U2436 (N_2436,N_1793,N_1911);
nand U2437 (N_2437,N_1698,N_1990);
and U2438 (N_2438,N_1591,N_1598);
and U2439 (N_2439,N_1942,N_1608);
and U2440 (N_2440,N_1873,N_1559);
and U2441 (N_2441,N_1639,N_1594);
or U2442 (N_2442,N_1664,N_1572);
and U2443 (N_2443,N_1591,N_1641);
nand U2444 (N_2444,N_1857,N_1702);
nor U2445 (N_2445,N_1729,N_1960);
nor U2446 (N_2446,N_1731,N_1639);
or U2447 (N_2447,N_1536,N_1966);
and U2448 (N_2448,N_1651,N_1964);
and U2449 (N_2449,N_1845,N_1633);
nand U2450 (N_2450,N_1508,N_1833);
nand U2451 (N_2451,N_1927,N_1646);
or U2452 (N_2452,N_1653,N_1713);
nand U2453 (N_2453,N_1984,N_1883);
xor U2454 (N_2454,N_1582,N_1991);
nor U2455 (N_2455,N_1663,N_1615);
nand U2456 (N_2456,N_1614,N_1989);
and U2457 (N_2457,N_1768,N_1949);
or U2458 (N_2458,N_1588,N_1534);
or U2459 (N_2459,N_1502,N_1983);
nand U2460 (N_2460,N_1562,N_1922);
or U2461 (N_2461,N_1598,N_1512);
or U2462 (N_2462,N_1692,N_1850);
and U2463 (N_2463,N_1613,N_1746);
nand U2464 (N_2464,N_1917,N_1893);
and U2465 (N_2465,N_1679,N_1835);
nand U2466 (N_2466,N_1696,N_1684);
and U2467 (N_2467,N_1506,N_1652);
xnor U2468 (N_2468,N_1782,N_1559);
nor U2469 (N_2469,N_1752,N_1897);
nand U2470 (N_2470,N_1858,N_1812);
or U2471 (N_2471,N_1660,N_1554);
xnor U2472 (N_2472,N_1880,N_1675);
nor U2473 (N_2473,N_1674,N_1859);
and U2474 (N_2474,N_1955,N_1539);
nand U2475 (N_2475,N_1664,N_1961);
and U2476 (N_2476,N_1958,N_1784);
and U2477 (N_2477,N_1894,N_1802);
and U2478 (N_2478,N_1763,N_1766);
and U2479 (N_2479,N_1926,N_1796);
nand U2480 (N_2480,N_1616,N_1614);
or U2481 (N_2481,N_1978,N_1574);
or U2482 (N_2482,N_1991,N_1998);
nand U2483 (N_2483,N_1555,N_1579);
or U2484 (N_2484,N_1522,N_1638);
or U2485 (N_2485,N_1607,N_1806);
and U2486 (N_2486,N_1521,N_1535);
and U2487 (N_2487,N_1863,N_1914);
nor U2488 (N_2488,N_1683,N_1891);
and U2489 (N_2489,N_1784,N_1505);
nor U2490 (N_2490,N_1891,N_1919);
and U2491 (N_2491,N_1590,N_1799);
nand U2492 (N_2492,N_1899,N_1831);
nand U2493 (N_2493,N_1778,N_1608);
and U2494 (N_2494,N_1657,N_1858);
nand U2495 (N_2495,N_1757,N_1783);
or U2496 (N_2496,N_1938,N_1939);
nor U2497 (N_2497,N_1928,N_1788);
and U2498 (N_2498,N_1571,N_1995);
or U2499 (N_2499,N_1699,N_1907);
and U2500 (N_2500,N_2073,N_2284);
or U2501 (N_2501,N_2424,N_2233);
or U2502 (N_2502,N_2287,N_2382);
and U2503 (N_2503,N_2057,N_2412);
nor U2504 (N_2504,N_2294,N_2102);
nand U2505 (N_2505,N_2147,N_2394);
or U2506 (N_2506,N_2099,N_2471);
and U2507 (N_2507,N_2276,N_2184);
or U2508 (N_2508,N_2070,N_2144);
nand U2509 (N_2509,N_2337,N_2479);
nand U2510 (N_2510,N_2186,N_2122);
xor U2511 (N_2511,N_2422,N_2464);
or U2512 (N_2512,N_2261,N_2039);
or U2513 (N_2513,N_2248,N_2267);
or U2514 (N_2514,N_2333,N_2413);
and U2515 (N_2515,N_2243,N_2487);
and U2516 (N_2516,N_2035,N_2086);
and U2517 (N_2517,N_2262,N_2058);
nor U2518 (N_2518,N_2236,N_2133);
nand U2519 (N_2519,N_2385,N_2069);
and U2520 (N_2520,N_2112,N_2223);
or U2521 (N_2521,N_2062,N_2209);
nand U2522 (N_2522,N_2389,N_2029);
xnor U2523 (N_2523,N_2085,N_2254);
nand U2524 (N_2524,N_2020,N_2410);
nor U2525 (N_2525,N_2059,N_2375);
or U2526 (N_2526,N_2170,N_2264);
or U2527 (N_2527,N_2492,N_2229);
nor U2528 (N_2528,N_2338,N_2392);
nand U2529 (N_2529,N_2381,N_2414);
nand U2530 (N_2530,N_2190,N_2369);
nor U2531 (N_2531,N_2352,N_2119);
or U2532 (N_2532,N_2089,N_2242);
nor U2533 (N_2533,N_2280,N_2279);
and U2534 (N_2534,N_2449,N_2241);
or U2535 (N_2535,N_2444,N_2151);
or U2536 (N_2536,N_2308,N_2169);
nand U2537 (N_2537,N_2268,N_2436);
and U2538 (N_2538,N_2297,N_2218);
nand U2539 (N_2539,N_2149,N_2051);
and U2540 (N_2540,N_2012,N_2165);
or U2541 (N_2541,N_2457,N_2499);
or U2542 (N_2542,N_2328,N_2216);
and U2543 (N_2543,N_2494,N_2025);
or U2544 (N_2544,N_2423,N_2010);
or U2545 (N_2545,N_2143,N_2238);
or U2546 (N_2546,N_2040,N_2088);
and U2547 (N_2547,N_2019,N_2235);
nor U2548 (N_2548,N_2068,N_2199);
nor U2549 (N_2549,N_2317,N_2015);
or U2550 (N_2550,N_2038,N_2082);
nor U2551 (N_2551,N_2446,N_2314);
or U2552 (N_2552,N_2318,N_2316);
or U2553 (N_2553,N_2064,N_2275);
nor U2554 (N_2554,N_2255,N_2386);
nand U2555 (N_2555,N_2176,N_2211);
nor U2556 (N_2556,N_2077,N_2008);
nor U2557 (N_2557,N_2072,N_2116);
and U2558 (N_2558,N_2101,N_2154);
or U2559 (N_2559,N_2166,N_2074);
nor U2560 (N_2560,N_2439,N_2152);
xor U2561 (N_2561,N_2331,N_2044);
or U2562 (N_2562,N_2431,N_2196);
nor U2563 (N_2563,N_2193,N_2053);
and U2564 (N_2564,N_2172,N_2142);
xor U2565 (N_2565,N_2079,N_2266);
nor U2566 (N_2566,N_2213,N_2183);
xnor U2567 (N_2567,N_2167,N_2452);
and U2568 (N_2568,N_2356,N_2031);
and U2569 (N_2569,N_2360,N_2127);
nand U2570 (N_2570,N_2011,N_2107);
or U2571 (N_2571,N_2054,N_2226);
nor U2572 (N_2572,N_2168,N_2370);
or U2573 (N_2573,N_2322,N_2249);
xor U2574 (N_2574,N_2456,N_2002);
nand U2575 (N_2575,N_2361,N_2036);
and U2576 (N_2576,N_2140,N_2081);
nor U2577 (N_2577,N_2224,N_2001);
nor U2578 (N_2578,N_2174,N_2427);
or U2579 (N_2579,N_2451,N_2357);
nand U2580 (N_2580,N_2365,N_2293);
or U2581 (N_2581,N_2027,N_2030);
nor U2582 (N_2582,N_2239,N_2497);
or U2583 (N_2583,N_2372,N_2325);
or U2584 (N_2584,N_2055,N_2219);
or U2585 (N_2585,N_2378,N_2335);
and U2586 (N_2586,N_2201,N_2390);
xor U2587 (N_2587,N_2334,N_2164);
nor U2588 (N_2588,N_2117,N_2398);
or U2589 (N_2589,N_2206,N_2135);
nand U2590 (N_2590,N_2221,N_2013);
nor U2591 (N_2591,N_2491,N_2026);
nor U2592 (N_2592,N_2336,N_2046);
and U2593 (N_2593,N_2182,N_2292);
or U2594 (N_2594,N_2300,N_2438);
or U2595 (N_2595,N_2291,N_2084);
nand U2596 (N_2596,N_2366,N_2047);
and U2597 (N_2597,N_2227,N_2091);
and U2598 (N_2598,N_2415,N_2230);
or U2599 (N_2599,N_2159,N_2490);
nand U2600 (N_2600,N_2472,N_2130);
nand U2601 (N_2601,N_2194,N_2080);
nor U2602 (N_2602,N_2161,N_2245);
xor U2603 (N_2603,N_2450,N_2309);
nand U2604 (N_2604,N_2098,N_2087);
nand U2605 (N_2605,N_2049,N_2045);
or U2606 (N_2606,N_2301,N_2124);
nor U2607 (N_2607,N_2401,N_2028);
nand U2608 (N_2608,N_2063,N_2484);
nand U2609 (N_2609,N_2203,N_2353);
nor U2610 (N_2610,N_2374,N_2037);
nor U2611 (N_2611,N_2195,N_2106);
nor U2612 (N_2612,N_2368,N_2111);
or U2613 (N_2613,N_2437,N_2380);
or U2614 (N_2614,N_2488,N_2339);
nand U2615 (N_2615,N_2480,N_2260);
or U2616 (N_2616,N_2426,N_2313);
and U2617 (N_2617,N_2458,N_2495);
nand U2618 (N_2618,N_2420,N_2327);
nand U2619 (N_2619,N_2061,N_2018);
nand U2620 (N_2620,N_2258,N_2311);
nor U2621 (N_2621,N_2312,N_2232);
and U2622 (N_2622,N_2060,N_2470);
nand U2623 (N_2623,N_2179,N_2278);
nor U2624 (N_2624,N_2461,N_2024);
nand U2625 (N_2625,N_2173,N_2104);
nand U2626 (N_2626,N_2341,N_2425);
nor U2627 (N_2627,N_2421,N_2139);
nand U2628 (N_2628,N_2187,N_2363);
nand U2629 (N_2629,N_2468,N_2498);
and U2630 (N_2630,N_2185,N_2113);
and U2631 (N_2631,N_2406,N_2244);
xor U2632 (N_2632,N_2282,N_2343);
nand U2633 (N_2633,N_2296,N_2396);
and U2634 (N_2634,N_2136,N_2197);
and U2635 (N_2635,N_2347,N_2283);
and U2636 (N_2636,N_2092,N_2453);
nand U2637 (N_2637,N_2114,N_2340);
nor U2638 (N_2638,N_2065,N_2475);
or U2639 (N_2639,N_2447,N_2489);
nor U2640 (N_2640,N_2274,N_2295);
nor U2641 (N_2641,N_2402,N_2319);
and U2642 (N_2642,N_2251,N_2052);
or U2643 (N_2643,N_2463,N_2007);
or U2644 (N_2644,N_2466,N_2324);
nor U2645 (N_2645,N_2332,N_2156);
nor U2646 (N_2646,N_2289,N_2455);
nor U2647 (N_2647,N_2393,N_2105);
and U2648 (N_2648,N_2126,N_2141);
and U2649 (N_2649,N_2477,N_2454);
nor U2650 (N_2650,N_2417,N_2004);
nand U2651 (N_2651,N_2407,N_2342);
nand U2652 (N_2652,N_2399,N_2348);
nand U2653 (N_2653,N_2305,N_2178);
and U2654 (N_2654,N_2066,N_2288);
and U2655 (N_2655,N_2000,N_2355);
nor U2656 (N_2656,N_2465,N_2388);
nor U2657 (N_2657,N_2003,N_2162);
nand U2658 (N_2658,N_2071,N_2033);
nand U2659 (N_2659,N_2397,N_2171);
or U2660 (N_2660,N_2391,N_2448);
xnor U2661 (N_2661,N_2434,N_2217);
nor U2662 (N_2662,N_2009,N_2097);
nor U2663 (N_2663,N_2210,N_2181);
and U2664 (N_2664,N_2253,N_2250);
or U2665 (N_2665,N_2202,N_2485);
and U2666 (N_2666,N_2138,N_2272);
nor U2667 (N_2667,N_2376,N_2359);
and U2668 (N_2668,N_2377,N_2271);
nand U2669 (N_2669,N_2125,N_2215);
nand U2670 (N_2670,N_2323,N_2214);
or U2671 (N_2671,N_2281,N_2017);
nor U2672 (N_2672,N_2474,N_2299);
or U2673 (N_2673,N_2100,N_2428);
or U2674 (N_2674,N_2307,N_2345);
nor U2675 (N_2675,N_2373,N_2022);
and U2676 (N_2676,N_2096,N_2445);
and U2677 (N_2677,N_2131,N_2443);
nand U2678 (N_2678,N_2351,N_2483);
or U2679 (N_2679,N_2408,N_2432);
nand U2680 (N_2680,N_2270,N_2304);
or U2681 (N_2681,N_2042,N_2109);
or U2682 (N_2682,N_2234,N_2459);
nand U2683 (N_2683,N_2405,N_2371);
and U2684 (N_2684,N_2212,N_2076);
and U2685 (N_2685,N_2032,N_2358);
nor U2686 (N_2686,N_2330,N_2277);
nand U2687 (N_2687,N_2155,N_2403);
nand U2688 (N_2688,N_2418,N_2259);
nand U2689 (N_2689,N_2476,N_2481);
or U2690 (N_2690,N_2191,N_2128);
or U2691 (N_2691,N_2257,N_2429);
or U2692 (N_2692,N_2469,N_2188);
and U2693 (N_2693,N_2349,N_2246);
nand U2694 (N_2694,N_2048,N_2460);
nand U2695 (N_2695,N_2326,N_2200);
nor U2696 (N_2696,N_2228,N_2329);
and U2697 (N_2697,N_2362,N_2043);
nor U2698 (N_2698,N_2321,N_2050);
nor U2699 (N_2699,N_2384,N_2198);
nand U2700 (N_2700,N_2462,N_2220);
nor U2701 (N_2701,N_2237,N_2387);
and U2702 (N_2702,N_2482,N_2120);
and U2703 (N_2703,N_2067,N_2473);
nor U2704 (N_2704,N_2395,N_2041);
and U2705 (N_2705,N_2177,N_2416);
or U2706 (N_2706,N_2435,N_2346);
nor U2707 (N_2707,N_2145,N_2252);
or U2708 (N_2708,N_2129,N_2146);
nor U2709 (N_2709,N_2240,N_2180);
and U2710 (N_2710,N_2354,N_2192);
and U2711 (N_2711,N_2021,N_2285);
and U2712 (N_2712,N_2083,N_2404);
nor U2713 (N_2713,N_2400,N_2350);
or U2714 (N_2714,N_2023,N_2110);
or U2715 (N_2715,N_2442,N_2430);
or U2716 (N_2716,N_2419,N_2189);
and U2717 (N_2717,N_2411,N_2263);
nand U2718 (N_2718,N_2163,N_2302);
nor U2719 (N_2719,N_2409,N_2175);
nand U2720 (N_2720,N_2364,N_2379);
and U2721 (N_2721,N_2005,N_2231);
and U2722 (N_2722,N_2290,N_2134);
and U2723 (N_2723,N_2310,N_2440);
or U2724 (N_2724,N_2467,N_2075);
or U2725 (N_2725,N_2123,N_2132);
nor U2726 (N_2726,N_2486,N_2222);
and U2727 (N_2727,N_2496,N_2150);
nor U2728 (N_2728,N_2014,N_2121);
or U2729 (N_2729,N_2208,N_2108);
and U2730 (N_2730,N_2148,N_2090);
nand U2731 (N_2731,N_2247,N_2094);
or U2732 (N_2732,N_2383,N_2153);
nand U2733 (N_2733,N_2315,N_2256);
or U2734 (N_2734,N_2303,N_2367);
or U2735 (N_2735,N_2137,N_2158);
nand U2736 (N_2736,N_2306,N_2093);
and U2737 (N_2737,N_2034,N_2016);
or U2738 (N_2738,N_2103,N_2118);
and U2739 (N_2739,N_2441,N_2269);
and U2740 (N_2740,N_2433,N_2207);
xor U2741 (N_2741,N_2204,N_2115);
nand U2742 (N_2742,N_2265,N_2205);
nand U2743 (N_2743,N_2320,N_2078);
or U2744 (N_2744,N_2478,N_2006);
or U2745 (N_2745,N_2286,N_2273);
or U2746 (N_2746,N_2298,N_2157);
or U2747 (N_2747,N_2056,N_2225);
or U2748 (N_2748,N_2344,N_2160);
nor U2749 (N_2749,N_2493,N_2095);
or U2750 (N_2750,N_2397,N_2027);
nand U2751 (N_2751,N_2487,N_2286);
nand U2752 (N_2752,N_2471,N_2127);
or U2753 (N_2753,N_2290,N_2076);
nor U2754 (N_2754,N_2141,N_2379);
or U2755 (N_2755,N_2105,N_2427);
nand U2756 (N_2756,N_2053,N_2211);
and U2757 (N_2757,N_2258,N_2029);
nand U2758 (N_2758,N_2008,N_2090);
nor U2759 (N_2759,N_2478,N_2288);
nor U2760 (N_2760,N_2412,N_2153);
and U2761 (N_2761,N_2328,N_2055);
nor U2762 (N_2762,N_2470,N_2378);
or U2763 (N_2763,N_2210,N_2279);
and U2764 (N_2764,N_2279,N_2251);
nand U2765 (N_2765,N_2188,N_2291);
and U2766 (N_2766,N_2477,N_2357);
nand U2767 (N_2767,N_2106,N_2077);
or U2768 (N_2768,N_2130,N_2383);
nor U2769 (N_2769,N_2386,N_2232);
and U2770 (N_2770,N_2262,N_2258);
and U2771 (N_2771,N_2247,N_2076);
nand U2772 (N_2772,N_2188,N_2384);
nor U2773 (N_2773,N_2144,N_2427);
or U2774 (N_2774,N_2027,N_2174);
and U2775 (N_2775,N_2232,N_2293);
nand U2776 (N_2776,N_2325,N_2046);
nor U2777 (N_2777,N_2198,N_2490);
and U2778 (N_2778,N_2217,N_2435);
and U2779 (N_2779,N_2457,N_2317);
and U2780 (N_2780,N_2260,N_2359);
or U2781 (N_2781,N_2065,N_2271);
nor U2782 (N_2782,N_2488,N_2074);
nor U2783 (N_2783,N_2422,N_2258);
or U2784 (N_2784,N_2257,N_2075);
or U2785 (N_2785,N_2135,N_2047);
and U2786 (N_2786,N_2315,N_2247);
or U2787 (N_2787,N_2171,N_2174);
or U2788 (N_2788,N_2342,N_2065);
or U2789 (N_2789,N_2400,N_2007);
or U2790 (N_2790,N_2257,N_2471);
nand U2791 (N_2791,N_2294,N_2430);
or U2792 (N_2792,N_2204,N_2022);
nand U2793 (N_2793,N_2275,N_2305);
nand U2794 (N_2794,N_2245,N_2270);
nor U2795 (N_2795,N_2321,N_2092);
nand U2796 (N_2796,N_2024,N_2447);
and U2797 (N_2797,N_2339,N_2121);
nor U2798 (N_2798,N_2307,N_2406);
nor U2799 (N_2799,N_2183,N_2032);
xor U2800 (N_2800,N_2384,N_2336);
nand U2801 (N_2801,N_2015,N_2269);
nor U2802 (N_2802,N_2362,N_2405);
or U2803 (N_2803,N_2363,N_2380);
nand U2804 (N_2804,N_2210,N_2390);
or U2805 (N_2805,N_2287,N_2017);
or U2806 (N_2806,N_2208,N_2082);
and U2807 (N_2807,N_2180,N_2297);
or U2808 (N_2808,N_2016,N_2423);
or U2809 (N_2809,N_2485,N_2419);
or U2810 (N_2810,N_2258,N_2451);
xnor U2811 (N_2811,N_2075,N_2099);
nand U2812 (N_2812,N_2088,N_2248);
and U2813 (N_2813,N_2179,N_2011);
and U2814 (N_2814,N_2056,N_2374);
nand U2815 (N_2815,N_2255,N_2491);
nor U2816 (N_2816,N_2466,N_2221);
or U2817 (N_2817,N_2217,N_2208);
nand U2818 (N_2818,N_2037,N_2174);
and U2819 (N_2819,N_2358,N_2224);
nor U2820 (N_2820,N_2143,N_2178);
and U2821 (N_2821,N_2423,N_2349);
nand U2822 (N_2822,N_2144,N_2187);
or U2823 (N_2823,N_2486,N_2213);
xor U2824 (N_2824,N_2263,N_2259);
nand U2825 (N_2825,N_2191,N_2059);
and U2826 (N_2826,N_2079,N_2480);
and U2827 (N_2827,N_2499,N_2243);
and U2828 (N_2828,N_2432,N_2193);
and U2829 (N_2829,N_2101,N_2057);
and U2830 (N_2830,N_2069,N_2362);
and U2831 (N_2831,N_2366,N_2485);
or U2832 (N_2832,N_2295,N_2479);
or U2833 (N_2833,N_2307,N_2125);
or U2834 (N_2834,N_2497,N_2124);
and U2835 (N_2835,N_2344,N_2304);
and U2836 (N_2836,N_2388,N_2222);
or U2837 (N_2837,N_2456,N_2373);
or U2838 (N_2838,N_2078,N_2278);
or U2839 (N_2839,N_2132,N_2220);
or U2840 (N_2840,N_2138,N_2415);
or U2841 (N_2841,N_2065,N_2399);
and U2842 (N_2842,N_2254,N_2224);
nor U2843 (N_2843,N_2191,N_2196);
nand U2844 (N_2844,N_2198,N_2113);
nor U2845 (N_2845,N_2121,N_2056);
nand U2846 (N_2846,N_2147,N_2287);
xnor U2847 (N_2847,N_2015,N_2421);
and U2848 (N_2848,N_2148,N_2154);
and U2849 (N_2849,N_2386,N_2213);
or U2850 (N_2850,N_2081,N_2153);
nand U2851 (N_2851,N_2082,N_2014);
xor U2852 (N_2852,N_2479,N_2332);
and U2853 (N_2853,N_2389,N_2417);
or U2854 (N_2854,N_2315,N_2171);
or U2855 (N_2855,N_2465,N_2053);
nand U2856 (N_2856,N_2311,N_2145);
nor U2857 (N_2857,N_2470,N_2077);
and U2858 (N_2858,N_2104,N_2150);
nor U2859 (N_2859,N_2067,N_2376);
nor U2860 (N_2860,N_2304,N_2024);
or U2861 (N_2861,N_2272,N_2346);
or U2862 (N_2862,N_2496,N_2292);
or U2863 (N_2863,N_2250,N_2418);
and U2864 (N_2864,N_2331,N_2023);
nand U2865 (N_2865,N_2384,N_2279);
or U2866 (N_2866,N_2335,N_2422);
or U2867 (N_2867,N_2219,N_2359);
nor U2868 (N_2868,N_2384,N_2429);
nand U2869 (N_2869,N_2290,N_2082);
nor U2870 (N_2870,N_2220,N_2192);
or U2871 (N_2871,N_2249,N_2052);
nand U2872 (N_2872,N_2119,N_2422);
and U2873 (N_2873,N_2398,N_2153);
or U2874 (N_2874,N_2372,N_2312);
nor U2875 (N_2875,N_2060,N_2153);
nand U2876 (N_2876,N_2349,N_2468);
or U2877 (N_2877,N_2226,N_2393);
or U2878 (N_2878,N_2057,N_2493);
or U2879 (N_2879,N_2197,N_2206);
or U2880 (N_2880,N_2495,N_2005);
and U2881 (N_2881,N_2212,N_2186);
or U2882 (N_2882,N_2383,N_2176);
or U2883 (N_2883,N_2189,N_2090);
nand U2884 (N_2884,N_2203,N_2335);
and U2885 (N_2885,N_2312,N_2049);
nor U2886 (N_2886,N_2051,N_2054);
nor U2887 (N_2887,N_2393,N_2308);
and U2888 (N_2888,N_2419,N_2147);
or U2889 (N_2889,N_2491,N_2186);
or U2890 (N_2890,N_2144,N_2432);
and U2891 (N_2891,N_2217,N_2029);
nor U2892 (N_2892,N_2113,N_2422);
and U2893 (N_2893,N_2196,N_2041);
nor U2894 (N_2894,N_2370,N_2492);
and U2895 (N_2895,N_2328,N_2035);
nand U2896 (N_2896,N_2413,N_2320);
or U2897 (N_2897,N_2120,N_2021);
or U2898 (N_2898,N_2445,N_2195);
or U2899 (N_2899,N_2423,N_2252);
nor U2900 (N_2900,N_2080,N_2326);
or U2901 (N_2901,N_2355,N_2223);
xnor U2902 (N_2902,N_2116,N_2388);
and U2903 (N_2903,N_2317,N_2158);
nor U2904 (N_2904,N_2077,N_2420);
or U2905 (N_2905,N_2477,N_2191);
or U2906 (N_2906,N_2056,N_2360);
or U2907 (N_2907,N_2107,N_2341);
and U2908 (N_2908,N_2087,N_2078);
nand U2909 (N_2909,N_2336,N_2035);
and U2910 (N_2910,N_2317,N_2315);
nand U2911 (N_2911,N_2061,N_2387);
nand U2912 (N_2912,N_2115,N_2195);
xor U2913 (N_2913,N_2108,N_2177);
nor U2914 (N_2914,N_2087,N_2287);
and U2915 (N_2915,N_2044,N_2201);
nor U2916 (N_2916,N_2357,N_2150);
nand U2917 (N_2917,N_2412,N_2229);
xor U2918 (N_2918,N_2064,N_2300);
or U2919 (N_2919,N_2029,N_2174);
and U2920 (N_2920,N_2153,N_2418);
nand U2921 (N_2921,N_2064,N_2216);
and U2922 (N_2922,N_2459,N_2456);
nor U2923 (N_2923,N_2331,N_2370);
nor U2924 (N_2924,N_2458,N_2196);
or U2925 (N_2925,N_2443,N_2207);
xnor U2926 (N_2926,N_2007,N_2464);
or U2927 (N_2927,N_2499,N_2486);
or U2928 (N_2928,N_2139,N_2131);
nand U2929 (N_2929,N_2335,N_2051);
or U2930 (N_2930,N_2108,N_2169);
or U2931 (N_2931,N_2414,N_2403);
nand U2932 (N_2932,N_2071,N_2294);
or U2933 (N_2933,N_2039,N_2487);
or U2934 (N_2934,N_2098,N_2121);
nand U2935 (N_2935,N_2047,N_2329);
nand U2936 (N_2936,N_2009,N_2450);
or U2937 (N_2937,N_2351,N_2441);
or U2938 (N_2938,N_2172,N_2127);
and U2939 (N_2939,N_2271,N_2349);
or U2940 (N_2940,N_2260,N_2381);
and U2941 (N_2941,N_2296,N_2458);
or U2942 (N_2942,N_2021,N_2084);
nor U2943 (N_2943,N_2354,N_2347);
or U2944 (N_2944,N_2400,N_2153);
nor U2945 (N_2945,N_2083,N_2081);
and U2946 (N_2946,N_2048,N_2205);
or U2947 (N_2947,N_2288,N_2309);
or U2948 (N_2948,N_2123,N_2040);
nor U2949 (N_2949,N_2195,N_2496);
nor U2950 (N_2950,N_2313,N_2035);
and U2951 (N_2951,N_2013,N_2010);
and U2952 (N_2952,N_2074,N_2202);
or U2953 (N_2953,N_2132,N_2331);
nor U2954 (N_2954,N_2012,N_2497);
nor U2955 (N_2955,N_2213,N_2207);
nor U2956 (N_2956,N_2076,N_2285);
nor U2957 (N_2957,N_2385,N_2001);
or U2958 (N_2958,N_2187,N_2474);
or U2959 (N_2959,N_2177,N_2245);
nor U2960 (N_2960,N_2271,N_2228);
nand U2961 (N_2961,N_2196,N_2042);
and U2962 (N_2962,N_2399,N_2146);
or U2963 (N_2963,N_2499,N_2049);
and U2964 (N_2964,N_2178,N_2229);
nor U2965 (N_2965,N_2331,N_2115);
nor U2966 (N_2966,N_2385,N_2479);
nand U2967 (N_2967,N_2180,N_2446);
nand U2968 (N_2968,N_2406,N_2462);
nand U2969 (N_2969,N_2410,N_2266);
or U2970 (N_2970,N_2081,N_2222);
nand U2971 (N_2971,N_2125,N_2145);
nor U2972 (N_2972,N_2359,N_2477);
or U2973 (N_2973,N_2231,N_2125);
and U2974 (N_2974,N_2136,N_2369);
nand U2975 (N_2975,N_2118,N_2077);
xor U2976 (N_2976,N_2227,N_2271);
and U2977 (N_2977,N_2019,N_2303);
nor U2978 (N_2978,N_2254,N_2291);
or U2979 (N_2979,N_2216,N_2407);
and U2980 (N_2980,N_2406,N_2204);
and U2981 (N_2981,N_2360,N_2028);
xor U2982 (N_2982,N_2338,N_2239);
and U2983 (N_2983,N_2148,N_2475);
or U2984 (N_2984,N_2056,N_2291);
and U2985 (N_2985,N_2135,N_2025);
and U2986 (N_2986,N_2411,N_2426);
nand U2987 (N_2987,N_2303,N_2033);
nor U2988 (N_2988,N_2347,N_2005);
nand U2989 (N_2989,N_2463,N_2054);
or U2990 (N_2990,N_2303,N_2161);
or U2991 (N_2991,N_2411,N_2015);
nor U2992 (N_2992,N_2474,N_2152);
nand U2993 (N_2993,N_2183,N_2253);
nor U2994 (N_2994,N_2194,N_2103);
nor U2995 (N_2995,N_2336,N_2252);
nor U2996 (N_2996,N_2255,N_2021);
and U2997 (N_2997,N_2448,N_2230);
and U2998 (N_2998,N_2072,N_2274);
xnor U2999 (N_2999,N_2044,N_2245);
or U3000 (N_3000,N_2765,N_2700);
nand U3001 (N_3001,N_2792,N_2626);
or U3002 (N_3002,N_2972,N_2523);
nor U3003 (N_3003,N_2546,N_2576);
nand U3004 (N_3004,N_2808,N_2959);
or U3005 (N_3005,N_2529,N_2885);
or U3006 (N_3006,N_2917,N_2839);
nor U3007 (N_3007,N_2579,N_2571);
nand U3008 (N_3008,N_2535,N_2977);
nand U3009 (N_3009,N_2658,N_2630);
nand U3010 (N_3010,N_2807,N_2887);
nand U3011 (N_3011,N_2766,N_2914);
and U3012 (N_3012,N_2545,N_2679);
nor U3013 (N_3013,N_2804,N_2548);
or U3014 (N_3014,N_2783,N_2607);
and U3015 (N_3015,N_2553,N_2821);
nand U3016 (N_3016,N_2517,N_2729);
or U3017 (N_3017,N_2528,N_2895);
and U3018 (N_3018,N_2526,N_2787);
and U3019 (N_3019,N_2997,N_2777);
nand U3020 (N_3020,N_2978,N_2536);
and U3021 (N_3021,N_2996,N_2583);
or U3022 (N_3022,N_2936,N_2738);
or U3023 (N_3023,N_2613,N_2882);
nor U3024 (N_3024,N_2843,N_2877);
nor U3025 (N_3025,N_2805,N_2721);
and U3026 (N_3026,N_2860,N_2519);
or U3027 (N_3027,N_2920,N_2648);
nand U3028 (N_3028,N_2965,N_2889);
and U3029 (N_3029,N_2952,N_2511);
and U3030 (N_3030,N_2706,N_2503);
or U3031 (N_3031,N_2638,N_2662);
nand U3032 (N_3032,N_2934,N_2761);
and U3033 (N_3033,N_2675,N_2866);
nor U3034 (N_3034,N_2861,N_2764);
or U3035 (N_3035,N_2768,N_2999);
or U3036 (N_3036,N_2680,N_2522);
or U3037 (N_3037,N_2849,N_2689);
nand U3038 (N_3038,N_2995,N_2868);
and U3039 (N_3039,N_2784,N_2803);
nor U3040 (N_3040,N_2651,N_2994);
or U3041 (N_3041,N_2544,N_2875);
nand U3042 (N_3042,N_2916,N_2527);
and U3043 (N_3043,N_2743,N_2773);
nor U3044 (N_3044,N_2525,N_2670);
nor U3045 (N_3045,N_2964,N_2970);
nand U3046 (N_3046,N_2541,N_2898);
or U3047 (N_3047,N_2586,N_2534);
nor U3048 (N_3048,N_2793,N_2949);
and U3049 (N_3049,N_2930,N_2785);
xor U3050 (N_3050,N_2570,N_2696);
or U3051 (N_3051,N_2874,N_2833);
or U3052 (N_3052,N_2557,N_2590);
nor U3053 (N_3053,N_2826,N_2581);
nor U3054 (N_3054,N_2911,N_2718);
nor U3055 (N_3055,N_2666,N_2663);
and U3056 (N_3056,N_2615,N_2708);
or U3057 (N_3057,N_2817,N_2824);
nor U3058 (N_3058,N_2575,N_2789);
nand U3059 (N_3059,N_2669,N_2870);
or U3060 (N_3060,N_2744,N_2776);
or U3061 (N_3061,N_2888,N_2852);
nor U3062 (N_3062,N_2886,N_2775);
or U3063 (N_3063,N_2715,N_2802);
nor U3064 (N_3064,N_2984,N_2954);
and U3065 (N_3065,N_2893,N_2846);
and U3066 (N_3066,N_2509,N_2726);
nor U3067 (N_3067,N_2906,N_2565);
and U3068 (N_3068,N_2688,N_2909);
nand U3069 (N_3069,N_2656,N_2739);
nor U3070 (N_3070,N_2871,N_2512);
and U3071 (N_3071,N_2944,N_2747);
nand U3072 (N_3072,N_2629,N_2958);
or U3073 (N_3073,N_2791,N_2790);
nand U3074 (N_3074,N_2500,N_2732);
nand U3075 (N_3075,N_2676,N_2842);
and U3076 (N_3076,N_2634,N_2514);
nor U3077 (N_3077,N_2554,N_2502);
nor U3078 (N_3078,N_2928,N_2705);
nor U3079 (N_3079,N_2587,N_2598);
and U3080 (N_3080,N_2608,N_2844);
nand U3081 (N_3081,N_2961,N_2851);
and U3082 (N_3082,N_2814,N_2660);
and U3083 (N_3083,N_2505,N_2707);
or U3084 (N_3084,N_2655,N_2904);
nand U3085 (N_3085,N_2756,N_2683);
or U3086 (N_3086,N_2753,N_2653);
nand U3087 (N_3087,N_2899,N_2919);
nor U3088 (N_3088,N_2876,N_2574);
and U3089 (N_3089,N_2872,N_2672);
nor U3090 (N_3090,N_2588,N_2604);
nor U3091 (N_3091,N_2504,N_2837);
or U3092 (N_3092,N_2690,N_2645);
nand U3093 (N_3093,N_2813,N_2838);
or U3094 (N_3094,N_2563,N_2730);
or U3095 (N_3095,N_2508,N_2968);
nor U3096 (N_3096,N_2810,N_2760);
nor U3097 (N_3097,N_2682,N_2749);
nand U3098 (N_3098,N_2720,N_2903);
or U3099 (N_3099,N_2945,N_2606);
or U3100 (N_3100,N_2892,N_2782);
and U3101 (N_3101,N_2735,N_2521);
or U3102 (N_3102,N_2603,N_2797);
nor U3103 (N_3103,N_2585,N_2712);
or U3104 (N_3104,N_2767,N_2755);
and U3105 (N_3105,N_2639,N_2896);
or U3106 (N_3106,N_2533,N_2642);
and U3107 (N_3107,N_2991,N_2596);
xor U3108 (N_3108,N_2982,N_2652);
nand U3109 (N_3109,N_2897,N_2507);
nand U3110 (N_3110,N_2649,N_2723);
nand U3111 (N_3111,N_2741,N_2962);
and U3112 (N_3112,N_2880,N_2562);
nor U3113 (N_3113,N_2635,N_2901);
nor U3114 (N_3114,N_2524,N_2931);
nor U3115 (N_3115,N_2677,N_2580);
nor U3116 (N_3116,N_2569,N_2539);
and U3117 (N_3117,N_2647,N_2664);
or U3118 (N_3118,N_2905,N_2734);
nand U3119 (N_3119,N_2857,N_2678);
nor U3120 (N_3120,N_2573,N_2907);
nor U3121 (N_3121,N_2845,N_2622);
and U3122 (N_3122,N_2686,N_2543);
xnor U3123 (N_3123,N_2924,N_2819);
nand U3124 (N_3124,N_2549,N_2832);
and U3125 (N_3125,N_2616,N_2908);
and U3126 (N_3126,N_2912,N_2956);
and U3127 (N_3127,N_2589,N_2890);
nor U3128 (N_3128,N_2619,N_2520);
or U3129 (N_3129,N_2532,N_2811);
nand U3130 (N_3130,N_2746,N_2988);
nand U3131 (N_3131,N_2927,N_2702);
and U3132 (N_3132,N_2980,N_2929);
nor U3133 (N_3133,N_2542,N_2795);
nor U3134 (N_3134,N_2611,N_2750);
nand U3135 (N_3135,N_2836,N_2657);
or U3136 (N_3136,N_2973,N_2993);
or U3137 (N_3137,N_2618,N_2620);
and U3138 (N_3138,N_2617,N_2601);
nand U3139 (N_3139,N_2834,N_2591);
or U3140 (N_3140,N_2752,N_2640);
or U3141 (N_3141,N_2659,N_2922);
and U3142 (N_3142,N_2673,N_2740);
nor U3143 (N_3143,N_2825,N_2925);
nor U3144 (N_3144,N_2665,N_2711);
nor U3145 (N_3145,N_2884,N_2850);
and U3146 (N_3146,N_2989,N_2695);
xnor U3147 (N_3147,N_2883,N_2998);
nor U3148 (N_3148,N_2710,N_2551);
or U3149 (N_3149,N_2625,N_2831);
nor U3150 (N_3150,N_2698,N_2862);
or U3151 (N_3151,N_2537,N_2939);
and U3152 (N_3152,N_2841,N_2736);
nand U3153 (N_3153,N_2704,N_2778);
nand U3154 (N_3154,N_2624,N_2560);
or U3155 (N_3155,N_2891,N_2694);
and U3156 (N_3156,N_2812,N_2697);
nand U3157 (N_3157,N_2902,N_2572);
and U3158 (N_3158,N_2963,N_2742);
and U3159 (N_3159,N_2725,N_2801);
nand U3160 (N_3160,N_2681,N_2650);
and U3161 (N_3161,N_2967,N_2758);
nor U3162 (N_3162,N_2853,N_2828);
or U3163 (N_3163,N_2796,N_2863);
and U3164 (N_3164,N_2538,N_2960);
and U3165 (N_3165,N_2559,N_2722);
nand U3166 (N_3166,N_2724,N_2654);
nor U3167 (N_3167,N_2786,N_2564);
nor U3168 (N_3168,N_2913,N_2530);
or U3169 (N_3169,N_2516,N_2727);
or U3170 (N_3170,N_2667,N_2864);
nand U3171 (N_3171,N_2701,N_2771);
nand U3172 (N_3172,N_2582,N_2687);
nor U3173 (N_3173,N_2781,N_2774);
nor U3174 (N_3174,N_2602,N_2858);
nor U3175 (N_3175,N_2806,N_2894);
or U3176 (N_3176,N_2628,N_2829);
or U3177 (N_3177,N_2879,N_2501);
and U3178 (N_3178,N_2643,N_2685);
or U3179 (N_3179,N_2878,N_2609);
or U3180 (N_3180,N_2873,N_2915);
and U3181 (N_3181,N_2748,N_2910);
or U3182 (N_3182,N_2926,N_2728);
nor U3183 (N_3183,N_2780,N_2992);
nand U3184 (N_3184,N_2976,N_2631);
nand U3185 (N_3185,N_2568,N_2614);
nand U3186 (N_3186,N_2633,N_2578);
nor U3187 (N_3187,N_2921,N_2577);
nor U3188 (N_3188,N_2555,N_2900);
nor U3189 (N_3189,N_2599,N_2693);
nor U3190 (N_3190,N_2800,N_2757);
or U3191 (N_3191,N_2584,N_2558);
nor U3192 (N_3192,N_2933,N_2646);
or U3193 (N_3193,N_2869,N_2809);
nand U3194 (N_3194,N_2938,N_2798);
nor U3195 (N_3195,N_2847,N_2816);
nor U3196 (N_3196,N_2840,N_2594);
nor U3197 (N_3197,N_2547,N_2918);
nor U3198 (N_3198,N_2595,N_2957);
nand U3199 (N_3199,N_2703,N_2865);
nor U3200 (N_3200,N_2600,N_2567);
nor U3201 (N_3201,N_2762,N_2955);
nor U3202 (N_3202,N_2923,N_2621);
and U3203 (N_3203,N_2822,N_2610);
or U3204 (N_3204,N_2940,N_2943);
nand U3205 (N_3205,N_2947,N_2515);
xnor U3206 (N_3206,N_2605,N_2592);
nor U3207 (N_3207,N_2820,N_2942);
nor U3208 (N_3208,N_2794,N_2745);
nand U3209 (N_3209,N_2935,N_2531);
or U3210 (N_3210,N_2779,N_2751);
or U3211 (N_3211,N_2692,N_2510);
or U3212 (N_3212,N_2987,N_2856);
nor U3213 (N_3213,N_2716,N_2661);
nor U3214 (N_3214,N_2540,N_2731);
or U3215 (N_3215,N_2932,N_2763);
xor U3216 (N_3216,N_2859,N_2627);
or U3217 (N_3217,N_2772,N_2979);
or U3218 (N_3218,N_2881,N_2799);
or U3219 (N_3219,N_2975,N_2941);
and U3220 (N_3220,N_2953,N_2937);
and U3221 (N_3221,N_2855,N_2966);
nand U3222 (N_3222,N_2714,N_2983);
xor U3223 (N_3223,N_2719,N_2717);
or U3224 (N_3224,N_2674,N_2699);
and U3225 (N_3225,N_2830,N_2566);
and U3226 (N_3226,N_2969,N_2737);
nand U3227 (N_3227,N_2684,N_2691);
and U3228 (N_3228,N_2671,N_2815);
and U3229 (N_3229,N_2770,N_2644);
nor U3230 (N_3230,N_2593,N_2848);
or U3231 (N_3231,N_2835,N_2974);
nor U3232 (N_3232,N_2597,N_2769);
or U3233 (N_3233,N_2668,N_2552);
xnor U3234 (N_3234,N_2632,N_2641);
xor U3235 (N_3235,N_2854,N_2636);
nand U3236 (N_3236,N_2754,N_2950);
nor U3237 (N_3237,N_2951,N_2713);
or U3238 (N_3238,N_2709,N_2733);
or U3239 (N_3239,N_2948,N_2867);
or U3240 (N_3240,N_2946,N_2818);
nor U3241 (N_3241,N_2612,N_2637);
or U3242 (N_3242,N_2827,N_2788);
nor U3243 (N_3243,N_2623,N_2518);
or U3244 (N_3244,N_2759,N_2550);
xor U3245 (N_3245,N_2986,N_2556);
and U3246 (N_3246,N_2823,N_2990);
nor U3247 (N_3247,N_2561,N_2971);
and U3248 (N_3248,N_2985,N_2513);
nor U3249 (N_3249,N_2981,N_2506);
nand U3250 (N_3250,N_2711,N_2910);
or U3251 (N_3251,N_2647,N_2977);
nand U3252 (N_3252,N_2735,N_2656);
nand U3253 (N_3253,N_2986,N_2701);
nand U3254 (N_3254,N_2612,N_2713);
nand U3255 (N_3255,N_2581,N_2709);
or U3256 (N_3256,N_2765,N_2653);
nor U3257 (N_3257,N_2589,N_2770);
nand U3258 (N_3258,N_2571,N_2874);
nor U3259 (N_3259,N_2678,N_2769);
nor U3260 (N_3260,N_2943,N_2968);
and U3261 (N_3261,N_2993,N_2793);
or U3262 (N_3262,N_2956,N_2741);
or U3263 (N_3263,N_2946,N_2903);
and U3264 (N_3264,N_2853,N_2925);
and U3265 (N_3265,N_2987,N_2826);
nand U3266 (N_3266,N_2612,N_2663);
or U3267 (N_3267,N_2892,N_2713);
nor U3268 (N_3268,N_2692,N_2767);
nand U3269 (N_3269,N_2678,N_2980);
and U3270 (N_3270,N_2787,N_2574);
or U3271 (N_3271,N_2734,N_2504);
nand U3272 (N_3272,N_2912,N_2991);
nor U3273 (N_3273,N_2665,N_2542);
nor U3274 (N_3274,N_2531,N_2740);
and U3275 (N_3275,N_2824,N_2729);
nor U3276 (N_3276,N_2957,N_2607);
and U3277 (N_3277,N_2502,N_2508);
or U3278 (N_3278,N_2615,N_2796);
or U3279 (N_3279,N_2712,N_2686);
or U3280 (N_3280,N_2959,N_2831);
nand U3281 (N_3281,N_2649,N_2843);
or U3282 (N_3282,N_2825,N_2564);
and U3283 (N_3283,N_2896,N_2935);
nor U3284 (N_3284,N_2558,N_2748);
or U3285 (N_3285,N_2582,N_2605);
or U3286 (N_3286,N_2979,N_2816);
or U3287 (N_3287,N_2532,N_2819);
nor U3288 (N_3288,N_2971,N_2598);
or U3289 (N_3289,N_2947,N_2766);
nand U3290 (N_3290,N_2595,N_2867);
nand U3291 (N_3291,N_2972,N_2500);
nand U3292 (N_3292,N_2577,N_2847);
and U3293 (N_3293,N_2728,N_2592);
or U3294 (N_3294,N_2934,N_2683);
nand U3295 (N_3295,N_2969,N_2897);
or U3296 (N_3296,N_2546,N_2941);
or U3297 (N_3297,N_2677,N_2841);
nand U3298 (N_3298,N_2691,N_2952);
nor U3299 (N_3299,N_2565,N_2746);
or U3300 (N_3300,N_2816,N_2845);
nand U3301 (N_3301,N_2765,N_2611);
nand U3302 (N_3302,N_2982,N_2883);
nor U3303 (N_3303,N_2757,N_2735);
or U3304 (N_3304,N_2524,N_2753);
nor U3305 (N_3305,N_2665,N_2596);
and U3306 (N_3306,N_2750,N_2682);
or U3307 (N_3307,N_2852,N_2909);
nor U3308 (N_3308,N_2836,N_2611);
nor U3309 (N_3309,N_2759,N_2656);
nor U3310 (N_3310,N_2695,N_2978);
xor U3311 (N_3311,N_2839,N_2988);
or U3312 (N_3312,N_2996,N_2586);
and U3313 (N_3313,N_2552,N_2993);
and U3314 (N_3314,N_2718,N_2531);
nor U3315 (N_3315,N_2822,N_2826);
xnor U3316 (N_3316,N_2566,N_2508);
and U3317 (N_3317,N_2692,N_2965);
or U3318 (N_3318,N_2730,N_2785);
nand U3319 (N_3319,N_2520,N_2526);
nor U3320 (N_3320,N_2782,N_2809);
nor U3321 (N_3321,N_2907,N_2992);
nor U3322 (N_3322,N_2786,N_2751);
or U3323 (N_3323,N_2835,N_2949);
nor U3324 (N_3324,N_2519,N_2796);
or U3325 (N_3325,N_2677,N_2995);
and U3326 (N_3326,N_2771,N_2994);
or U3327 (N_3327,N_2733,N_2887);
xnor U3328 (N_3328,N_2860,N_2710);
xnor U3329 (N_3329,N_2842,N_2575);
and U3330 (N_3330,N_2726,N_2917);
or U3331 (N_3331,N_2890,N_2938);
xnor U3332 (N_3332,N_2561,N_2573);
nor U3333 (N_3333,N_2521,N_2853);
or U3334 (N_3334,N_2582,N_2739);
and U3335 (N_3335,N_2680,N_2717);
or U3336 (N_3336,N_2762,N_2791);
or U3337 (N_3337,N_2670,N_2774);
and U3338 (N_3338,N_2925,N_2796);
xnor U3339 (N_3339,N_2506,N_2906);
or U3340 (N_3340,N_2517,N_2579);
or U3341 (N_3341,N_2949,N_2909);
nand U3342 (N_3342,N_2779,N_2690);
nor U3343 (N_3343,N_2806,N_2678);
nand U3344 (N_3344,N_2654,N_2812);
or U3345 (N_3345,N_2854,N_2672);
nand U3346 (N_3346,N_2661,N_2837);
or U3347 (N_3347,N_2868,N_2828);
nor U3348 (N_3348,N_2539,N_2590);
nor U3349 (N_3349,N_2865,N_2578);
nor U3350 (N_3350,N_2789,N_2837);
and U3351 (N_3351,N_2671,N_2672);
xnor U3352 (N_3352,N_2673,N_2763);
or U3353 (N_3353,N_2865,N_2898);
nand U3354 (N_3354,N_2886,N_2677);
nor U3355 (N_3355,N_2524,N_2584);
xor U3356 (N_3356,N_2637,N_2684);
and U3357 (N_3357,N_2838,N_2584);
nand U3358 (N_3358,N_2625,N_2566);
and U3359 (N_3359,N_2719,N_2662);
nor U3360 (N_3360,N_2965,N_2922);
nand U3361 (N_3361,N_2505,N_2801);
nand U3362 (N_3362,N_2804,N_2598);
or U3363 (N_3363,N_2650,N_2829);
or U3364 (N_3364,N_2626,N_2945);
nor U3365 (N_3365,N_2778,N_2601);
nor U3366 (N_3366,N_2816,N_2654);
and U3367 (N_3367,N_2986,N_2856);
nor U3368 (N_3368,N_2587,N_2554);
nand U3369 (N_3369,N_2826,N_2972);
nand U3370 (N_3370,N_2663,N_2534);
nor U3371 (N_3371,N_2773,N_2882);
nand U3372 (N_3372,N_2794,N_2530);
nand U3373 (N_3373,N_2761,N_2820);
nand U3374 (N_3374,N_2637,N_2799);
and U3375 (N_3375,N_2666,N_2737);
nor U3376 (N_3376,N_2815,N_2989);
and U3377 (N_3377,N_2521,N_2799);
or U3378 (N_3378,N_2655,N_2979);
nand U3379 (N_3379,N_2777,N_2511);
nand U3380 (N_3380,N_2823,N_2586);
or U3381 (N_3381,N_2642,N_2743);
nand U3382 (N_3382,N_2954,N_2857);
and U3383 (N_3383,N_2639,N_2589);
or U3384 (N_3384,N_2731,N_2582);
and U3385 (N_3385,N_2595,N_2994);
nand U3386 (N_3386,N_2522,N_2974);
and U3387 (N_3387,N_2895,N_2978);
nand U3388 (N_3388,N_2978,N_2580);
nor U3389 (N_3389,N_2646,N_2742);
and U3390 (N_3390,N_2523,N_2880);
nor U3391 (N_3391,N_2786,N_2796);
xor U3392 (N_3392,N_2710,N_2545);
and U3393 (N_3393,N_2797,N_2864);
nand U3394 (N_3394,N_2913,N_2893);
or U3395 (N_3395,N_2716,N_2504);
and U3396 (N_3396,N_2825,N_2689);
or U3397 (N_3397,N_2898,N_2560);
nor U3398 (N_3398,N_2745,N_2718);
and U3399 (N_3399,N_2944,N_2756);
nand U3400 (N_3400,N_2697,N_2886);
nand U3401 (N_3401,N_2817,N_2532);
nand U3402 (N_3402,N_2712,N_2615);
or U3403 (N_3403,N_2913,N_2653);
nor U3404 (N_3404,N_2697,N_2575);
and U3405 (N_3405,N_2729,N_2536);
and U3406 (N_3406,N_2519,N_2721);
or U3407 (N_3407,N_2613,N_2832);
nand U3408 (N_3408,N_2895,N_2558);
or U3409 (N_3409,N_2796,N_2634);
nor U3410 (N_3410,N_2726,N_2806);
nand U3411 (N_3411,N_2729,N_2507);
nand U3412 (N_3412,N_2766,N_2739);
nor U3413 (N_3413,N_2616,N_2831);
nand U3414 (N_3414,N_2985,N_2502);
or U3415 (N_3415,N_2792,N_2599);
or U3416 (N_3416,N_2745,N_2608);
and U3417 (N_3417,N_2618,N_2672);
nor U3418 (N_3418,N_2540,N_2905);
nor U3419 (N_3419,N_2783,N_2714);
and U3420 (N_3420,N_2537,N_2575);
nor U3421 (N_3421,N_2678,N_2991);
or U3422 (N_3422,N_2903,N_2664);
nor U3423 (N_3423,N_2672,N_2576);
nor U3424 (N_3424,N_2532,N_2716);
nor U3425 (N_3425,N_2508,N_2585);
or U3426 (N_3426,N_2954,N_2867);
and U3427 (N_3427,N_2941,N_2960);
nor U3428 (N_3428,N_2789,N_2925);
and U3429 (N_3429,N_2715,N_2720);
nor U3430 (N_3430,N_2952,N_2807);
nand U3431 (N_3431,N_2561,N_2751);
and U3432 (N_3432,N_2729,N_2721);
or U3433 (N_3433,N_2534,N_2601);
and U3434 (N_3434,N_2552,N_2903);
and U3435 (N_3435,N_2532,N_2796);
and U3436 (N_3436,N_2534,N_2599);
and U3437 (N_3437,N_2845,N_2611);
and U3438 (N_3438,N_2560,N_2947);
or U3439 (N_3439,N_2738,N_2646);
and U3440 (N_3440,N_2942,N_2593);
and U3441 (N_3441,N_2925,N_2628);
nand U3442 (N_3442,N_2572,N_2735);
and U3443 (N_3443,N_2733,N_2706);
nand U3444 (N_3444,N_2640,N_2803);
or U3445 (N_3445,N_2935,N_2556);
or U3446 (N_3446,N_2508,N_2945);
or U3447 (N_3447,N_2726,N_2876);
nor U3448 (N_3448,N_2726,N_2900);
nand U3449 (N_3449,N_2890,N_2548);
nor U3450 (N_3450,N_2868,N_2920);
nor U3451 (N_3451,N_2779,N_2935);
and U3452 (N_3452,N_2550,N_2766);
nand U3453 (N_3453,N_2740,N_2626);
nor U3454 (N_3454,N_2760,N_2898);
and U3455 (N_3455,N_2971,N_2923);
nand U3456 (N_3456,N_2836,N_2723);
and U3457 (N_3457,N_2684,N_2527);
or U3458 (N_3458,N_2591,N_2819);
or U3459 (N_3459,N_2921,N_2611);
nor U3460 (N_3460,N_2632,N_2585);
or U3461 (N_3461,N_2961,N_2786);
and U3462 (N_3462,N_2727,N_2896);
nor U3463 (N_3463,N_2953,N_2853);
nand U3464 (N_3464,N_2562,N_2787);
nor U3465 (N_3465,N_2665,N_2950);
nand U3466 (N_3466,N_2955,N_2584);
or U3467 (N_3467,N_2819,N_2790);
nand U3468 (N_3468,N_2835,N_2792);
and U3469 (N_3469,N_2879,N_2730);
nor U3470 (N_3470,N_2900,N_2891);
nor U3471 (N_3471,N_2768,N_2967);
or U3472 (N_3472,N_2908,N_2965);
or U3473 (N_3473,N_2669,N_2628);
and U3474 (N_3474,N_2685,N_2589);
and U3475 (N_3475,N_2865,N_2938);
nor U3476 (N_3476,N_2862,N_2877);
nand U3477 (N_3477,N_2931,N_2862);
nand U3478 (N_3478,N_2502,N_2780);
nand U3479 (N_3479,N_2612,N_2613);
and U3480 (N_3480,N_2709,N_2861);
nand U3481 (N_3481,N_2854,N_2828);
nor U3482 (N_3482,N_2736,N_2519);
and U3483 (N_3483,N_2723,N_2964);
nand U3484 (N_3484,N_2680,N_2534);
or U3485 (N_3485,N_2705,N_2956);
nand U3486 (N_3486,N_2645,N_2601);
and U3487 (N_3487,N_2609,N_2522);
or U3488 (N_3488,N_2624,N_2603);
or U3489 (N_3489,N_2652,N_2833);
nand U3490 (N_3490,N_2536,N_2753);
and U3491 (N_3491,N_2604,N_2744);
xor U3492 (N_3492,N_2574,N_2887);
nand U3493 (N_3493,N_2542,N_2562);
or U3494 (N_3494,N_2714,N_2857);
and U3495 (N_3495,N_2726,N_2748);
nand U3496 (N_3496,N_2524,N_2935);
or U3497 (N_3497,N_2876,N_2674);
nand U3498 (N_3498,N_2770,N_2844);
and U3499 (N_3499,N_2810,N_2914);
nor U3500 (N_3500,N_3436,N_3154);
nand U3501 (N_3501,N_3437,N_3474);
nand U3502 (N_3502,N_3152,N_3447);
or U3503 (N_3503,N_3172,N_3469);
nand U3504 (N_3504,N_3106,N_3260);
and U3505 (N_3505,N_3457,N_3214);
nand U3506 (N_3506,N_3382,N_3180);
and U3507 (N_3507,N_3285,N_3332);
or U3508 (N_3508,N_3085,N_3265);
nor U3509 (N_3509,N_3092,N_3031);
and U3510 (N_3510,N_3270,N_3372);
nand U3511 (N_3511,N_3212,N_3290);
nor U3512 (N_3512,N_3241,N_3479);
and U3513 (N_3513,N_3462,N_3383);
or U3514 (N_3514,N_3103,N_3206);
nand U3515 (N_3515,N_3304,N_3319);
xnor U3516 (N_3516,N_3105,N_3418);
nor U3517 (N_3517,N_3042,N_3393);
nor U3518 (N_3518,N_3317,N_3416);
nor U3519 (N_3519,N_3312,N_3450);
nand U3520 (N_3520,N_3200,N_3489);
and U3521 (N_3521,N_3174,N_3033);
nand U3522 (N_3522,N_3122,N_3355);
or U3523 (N_3523,N_3003,N_3146);
nand U3524 (N_3524,N_3282,N_3448);
nand U3525 (N_3525,N_3252,N_3297);
nor U3526 (N_3526,N_3009,N_3158);
and U3527 (N_3527,N_3113,N_3077);
nor U3528 (N_3528,N_3468,N_3432);
xnor U3529 (N_3529,N_3164,N_3371);
or U3530 (N_3530,N_3150,N_3050);
and U3531 (N_3531,N_3037,N_3365);
xnor U3532 (N_3532,N_3095,N_3108);
or U3533 (N_3533,N_3300,N_3098);
nand U3534 (N_3534,N_3151,N_3499);
nor U3535 (N_3535,N_3153,N_3359);
and U3536 (N_3536,N_3331,N_3109);
and U3537 (N_3537,N_3013,N_3441);
or U3538 (N_3538,N_3134,N_3074);
or U3539 (N_3539,N_3305,N_3081);
nand U3540 (N_3540,N_3268,N_3217);
or U3541 (N_3541,N_3339,N_3406);
nand U3542 (N_3542,N_3353,N_3376);
nand U3543 (N_3543,N_3186,N_3222);
xor U3544 (N_3544,N_3254,N_3140);
and U3545 (N_3545,N_3478,N_3229);
nand U3546 (N_3546,N_3123,N_3367);
nor U3547 (N_3547,N_3024,N_3221);
nand U3548 (N_3548,N_3277,N_3173);
and U3549 (N_3549,N_3192,N_3067);
and U3550 (N_3550,N_3089,N_3093);
and U3551 (N_3551,N_3384,N_3345);
nor U3552 (N_3552,N_3328,N_3420);
and U3553 (N_3553,N_3047,N_3476);
xor U3554 (N_3554,N_3494,N_3149);
and U3555 (N_3555,N_3127,N_3073);
nand U3556 (N_3556,N_3043,N_3480);
nor U3557 (N_3557,N_3482,N_3204);
or U3558 (N_3558,N_3336,N_3057);
xnor U3559 (N_3559,N_3492,N_3280);
nor U3560 (N_3560,N_3400,N_3101);
and U3561 (N_3561,N_3491,N_3190);
and U3562 (N_3562,N_3213,N_3148);
or U3563 (N_3563,N_3230,N_3368);
xnor U3564 (N_3564,N_3251,N_3256);
nand U3565 (N_3565,N_3231,N_3329);
nand U3566 (N_3566,N_3263,N_3308);
or U3567 (N_3567,N_3198,N_3284);
and U3568 (N_3568,N_3159,N_3433);
nand U3569 (N_3569,N_3326,N_3264);
nand U3570 (N_3570,N_3205,N_3320);
nand U3571 (N_3571,N_3118,N_3288);
nor U3572 (N_3572,N_3028,N_3286);
and U3573 (N_3573,N_3082,N_3323);
nor U3574 (N_3574,N_3129,N_3216);
and U3575 (N_3575,N_3170,N_3340);
and U3576 (N_3576,N_3177,N_3207);
or U3577 (N_3577,N_3396,N_3071);
and U3578 (N_3578,N_3182,N_3488);
nor U3579 (N_3579,N_3338,N_3357);
nor U3580 (N_3580,N_3236,N_3049);
or U3581 (N_3581,N_3453,N_3160);
nor U3582 (N_3582,N_3327,N_3090);
nand U3583 (N_3583,N_3412,N_3379);
nor U3584 (N_3584,N_3070,N_3135);
and U3585 (N_3585,N_3211,N_3132);
nand U3586 (N_3586,N_3116,N_3165);
nand U3587 (N_3587,N_3008,N_3218);
and U3588 (N_3588,N_3343,N_3208);
nor U3589 (N_3589,N_3258,N_3004);
nor U3590 (N_3590,N_3012,N_3010);
and U3591 (N_3591,N_3321,N_3374);
and U3592 (N_3592,N_3193,N_3334);
and U3593 (N_3593,N_3295,N_3341);
or U3594 (N_3594,N_3189,N_3246);
or U3595 (N_3595,N_3114,N_3021);
nand U3596 (N_3596,N_3375,N_3157);
or U3597 (N_3597,N_3238,N_3446);
nand U3598 (N_3598,N_3032,N_3361);
or U3599 (N_3599,N_3459,N_3240);
and U3600 (N_3600,N_3405,N_3058);
nor U3601 (N_3601,N_3407,N_3387);
nor U3602 (N_3602,N_3318,N_3209);
nor U3603 (N_3603,N_3112,N_3066);
or U3604 (N_3604,N_3099,N_3171);
or U3605 (N_3605,N_3431,N_3039);
nor U3606 (N_3606,N_3451,N_3188);
or U3607 (N_3607,N_3430,N_3166);
nor U3608 (N_3608,N_3124,N_3036);
and U3609 (N_3609,N_3181,N_3274);
or U3610 (N_3610,N_3235,N_3460);
nand U3611 (N_3611,N_3377,N_3397);
and U3612 (N_3612,N_3056,N_3197);
xnor U3613 (N_3613,N_3360,N_3344);
nor U3614 (N_3614,N_3015,N_3248);
nand U3615 (N_3615,N_3237,N_3139);
and U3616 (N_3616,N_3141,N_3117);
nand U3617 (N_3617,N_3404,N_3311);
nand U3618 (N_3618,N_3330,N_3034);
and U3619 (N_3619,N_3120,N_3219);
and U3620 (N_3620,N_3275,N_3273);
or U3621 (N_3621,N_3322,N_3096);
or U3622 (N_3622,N_3363,N_3445);
and U3623 (N_3623,N_3429,N_3027);
nor U3624 (N_3624,N_3391,N_3084);
nand U3625 (N_3625,N_3271,N_3495);
and U3626 (N_3626,N_3194,N_3335);
or U3627 (N_3627,N_3267,N_3228);
and U3628 (N_3628,N_3247,N_3086);
and U3629 (N_3629,N_3473,N_3041);
and U3630 (N_3630,N_3060,N_3061);
or U3631 (N_3631,N_3310,N_3006);
nand U3632 (N_3632,N_3234,N_3301);
or U3633 (N_3633,N_3419,N_3244);
and U3634 (N_3634,N_3409,N_3121);
and U3635 (N_3635,N_3399,N_3401);
nor U3636 (N_3636,N_3131,N_3055);
nor U3637 (N_3637,N_3220,N_3291);
and U3638 (N_3638,N_3102,N_3294);
or U3639 (N_3639,N_3210,N_3444);
nor U3640 (N_3640,N_3163,N_3455);
nand U3641 (N_3641,N_3485,N_3381);
and U3642 (N_3642,N_3350,N_3201);
and U3643 (N_3643,N_3296,N_3410);
and U3644 (N_3644,N_3496,N_3063);
nor U3645 (N_3645,N_3463,N_3023);
nor U3646 (N_3646,N_3126,N_3225);
nor U3647 (N_3647,N_3438,N_3155);
nor U3648 (N_3648,N_3348,N_3456);
nand U3649 (N_3649,N_3133,N_3100);
xor U3650 (N_3650,N_3486,N_3064);
nand U3651 (N_3651,N_3094,N_3333);
nor U3652 (N_3652,N_3239,N_3424);
nand U3653 (N_3653,N_3342,N_3029);
nor U3654 (N_3654,N_3187,N_3325);
and U3655 (N_3655,N_3156,N_3421);
nor U3656 (N_3656,N_3232,N_3428);
or U3657 (N_3657,N_3179,N_3402);
nand U3658 (N_3658,N_3293,N_3005);
and U3659 (N_3659,N_3035,N_3169);
nor U3660 (N_3660,N_3000,N_3195);
and U3661 (N_3661,N_3119,N_3045);
and U3662 (N_3662,N_3366,N_3162);
and U3663 (N_3663,N_3227,N_3481);
and U3664 (N_3664,N_3255,N_3378);
nor U3665 (N_3665,N_3075,N_3143);
nor U3666 (N_3666,N_3097,N_3398);
nor U3667 (N_3667,N_3142,N_3083);
nand U3668 (N_3668,N_3422,N_3088);
nand U3669 (N_3669,N_3471,N_3349);
or U3670 (N_3670,N_3007,N_3487);
nor U3671 (N_3671,N_3245,N_3337);
or U3672 (N_3672,N_3373,N_3369);
and U3673 (N_3673,N_3426,N_3269);
and U3674 (N_3674,N_3253,N_3191);
and U3675 (N_3675,N_3415,N_3266);
and U3676 (N_3676,N_3395,N_3356);
or U3677 (N_3677,N_3014,N_3307);
nand U3678 (N_3678,N_3283,N_3130);
or U3679 (N_3679,N_3002,N_3168);
nand U3680 (N_3680,N_3138,N_3137);
and U3681 (N_3681,N_3440,N_3467);
nor U3682 (N_3682,N_3287,N_3223);
or U3683 (N_3683,N_3423,N_3046);
and U3684 (N_3684,N_3324,N_3026);
nand U3685 (N_3685,N_3392,N_3203);
nand U3686 (N_3686,N_3178,N_3370);
and U3687 (N_3687,N_3249,N_3261);
or U3688 (N_3688,N_3449,N_3040);
nor U3689 (N_3689,N_3389,N_3115);
or U3690 (N_3690,N_3062,N_3452);
or U3691 (N_3691,N_3016,N_3425);
and U3692 (N_3692,N_3025,N_3477);
nand U3693 (N_3693,N_3072,N_3443);
or U3694 (N_3694,N_3313,N_3069);
nand U3695 (N_3695,N_3362,N_3125);
and U3696 (N_3696,N_3272,N_3048);
nand U3697 (N_3697,N_3483,N_3161);
nand U3698 (N_3698,N_3059,N_3175);
or U3699 (N_3699,N_3314,N_3001);
nor U3700 (N_3700,N_3196,N_3454);
nor U3701 (N_3701,N_3281,N_3202);
nor U3702 (N_3702,N_3242,N_3104);
nand U3703 (N_3703,N_3298,N_3472);
and U3704 (N_3704,N_3018,N_3380);
nor U3705 (N_3705,N_3386,N_3167);
nand U3706 (N_3706,N_3465,N_3226);
and U3707 (N_3707,N_3078,N_3484);
nand U3708 (N_3708,N_3408,N_3352);
or U3709 (N_3709,N_3411,N_3414);
nor U3710 (N_3710,N_3019,N_3107);
nor U3711 (N_3711,N_3427,N_3315);
or U3712 (N_3712,N_3302,N_3136);
or U3713 (N_3713,N_3358,N_3091);
nand U3714 (N_3714,N_3289,N_3347);
nand U3715 (N_3715,N_3184,N_3493);
or U3716 (N_3716,N_3306,N_3199);
nor U3717 (N_3717,N_3038,N_3257);
nor U3718 (N_3718,N_3215,N_3299);
nor U3719 (N_3719,N_3128,N_3185);
nand U3720 (N_3720,N_3110,N_3434);
nand U3721 (N_3721,N_3458,N_3316);
and U3722 (N_3722,N_3262,N_3076);
and U3723 (N_3723,N_3011,N_3054);
nor U3724 (N_3724,N_3183,N_3346);
nor U3725 (N_3725,N_3497,N_3030);
or U3726 (N_3726,N_3292,N_3144);
nand U3727 (N_3727,N_3388,N_3243);
and U3728 (N_3728,N_3464,N_3435);
or U3729 (N_3729,N_3020,N_3080);
nand U3730 (N_3730,N_3475,N_3390);
and U3731 (N_3731,N_3490,N_3354);
or U3732 (N_3732,N_3224,N_3051);
or U3733 (N_3733,N_3276,N_3279);
or U3734 (N_3734,N_3022,N_3309);
nor U3735 (N_3735,N_3233,N_3394);
nand U3736 (N_3736,N_3498,N_3147);
nor U3737 (N_3737,N_3087,N_3461);
nand U3738 (N_3738,N_3466,N_3145);
xnor U3739 (N_3739,N_3470,N_3259);
nand U3740 (N_3740,N_3017,N_3278);
and U3741 (N_3741,N_3079,N_3403);
and U3742 (N_3742,N_3044,N_3111);
nor U3743 (N_3743,N_3439,N_3417);
nand U3744 (N_3744,N_3351,N_3385);
and U3745 (N_3745,N_3364,N_3053);
or U3746 (N_3746,N_3052,N_3413);
nor U3747 (N_3747,N_3176,N_3442);
nor U3748 (N_3748,N_3068,N_3303);
and U3749 (N_3749,N_3250,N_3065);
or U3750 (N_3750,N_3075,N_3436);
nor U3751 (N_3751,N_3245,N_3138);
or U3752 (N_3752,N_3155,N_3444);
nor U3753 (N_3753,N_3026,N_3101);
nand U3754 (N_3754,N_3354,N_3274);
nand U3755 (N_3755,N_3411,N_3484);
nor U3756 (N_3756,N_3401,N_3475);
nor U3757 (N_3757,N_3120,N_3172);
nand U3758 (N_3758,N_3363,N_3364);
xor U3759 (N_3759,N_3409,N_3274);
and U3760 (N_3760,N_3256,N_3257);
nand U3761 (N_3761,N_3455,N_3377);
nor U3762 (N_3762,N_3453,N_3454);
or U3763 (N_3763,N_3163,N_3231);
or U3764 (N_3764,N_3044,N_3446);
xor U3765 (N_3765,N_3082,N_3261);
nand U3766 (N_3766,N_3471,N_3497);
nor U3767 (N_3767,N_3131,N_3265);
nand U3768 (N_3768,N_3486,N_3302);
nor U3769 (N_3769,N_3093,N_3134);
and U3770 (N_3770,N_3424,N_3049);
nor U3771 (N_3771,N_3128,N_3447);
and U3772 (N_3772,N_3435,N_3044);
nor U3773 (N_3773,N_3143,N_3097);
nand U3774 (N_3774,N_3457,N_3199);
nand U3775 (N_3775,N_3039,N_3151);
and U3776 (N_3776,N_3153,N_3364);
nand U3777 (N_3777,N_3450,N_3091);
nor U3778 (N_3778,N_3342,N_3192);
nor U3779 (N_3779,N_3020,N_3180);
and U3780 (N_3780,N_3426,N_3265);
nor U3781 (N_3781,N_3293,N_3200);
or U3782 (N_3782,N_3209,N_3230);
nand U3783 (N_3783,N_3486,N_3250);
and U3784 (N_3784,N_3492,N_3482);
or U3785 (N_3785,N_3160,N_3052);
nor U3786 (N_3786,N_3224,N_3072);
and U3787 (N_3787,N_3128,N_3270);
nand U3788 (N_3788,N_3095,N_3060);
xnor U3789 (N_3789,N_3253,N_3025);
nor U3790 (N_3790,N_3070,N_3288);
and U3791 (N_3791,N_3361,N_3179);
xor U3792 (N_3792,N_3203,N_3193);
or U3793 (N_3793,N_3130,N_3002);
nor U3794 (N_3794,N_3441,N_3070);
and U3795 (N_3795,N_3092,N_3450);
xor U3796 (N_3796,N_3381,N_3356);
or U3797 (N_3797,N_3077,N_3116);
nand U3798 (N_3798,N_3191,N_3126);
nand U3799 (N_3799,N_3406,N_3156);
nand U3800 (N_3800,N_3380,N_3270);
nor U3801 (N_3801,N_3119,N_3219);
and U3802 (N_3802,N_3313,N_3039);
or U3803 (N_3803,N_3127,N_3453);
and U3804 (N_3804,N_3269,N_3028);
or U3805 (N_3805,N_3031,N_3491);
and U3806 (N_3806,N_3487,N_3405);
nand U3807 (N_3807,N_3309,N_3429);
nand U3808 (N_3808,N_3330,N_3060);
nand U3809 (N_3809,N_3125,N_3215);
or U3810 (N_3810,N_3297,N_3092);
nor U3811 (N_3811,N_3022,N_3051);
and U3812 (N_3812,N_3379,N_3328);
nor U3813 (N_3813,N_3178,N_3332);
and U3814 (N_3814,N_3368,N_3201);
and U3815 (N_3815,N_3406,N_3400);
and U3816 (N_3816,N_3478,N_3256);
nor U3817 (N_3817,N_3462,N_3339);
or U3818 (N_3818,N_3047,N_3442);
nor U3819 (N_3819,N_3448,N_3105);
or U3820 (N_3820,N_3465,N_3388);
or U3821 (N_3821,N_3368,N_3496);
or U3822 (N_3822,N_3143,N_3273);
nand U3823 (N_3823,N_3041,N_3403);
and U3824 (N_3824,N_3383,N_3107);
and U3825 (N_3825,N_3444,N_3465);
nor U3826 (N_3826,N_3007,N_3080);
nor U3827 (N_3827,N_3070,N_3008);
nor U3828 (N_3828,N_3033,N_3220);
or U3829 (N_3829,N_3075,N_3015);
nor U3830 (N_3830,N_3017,N_3387);
nor U3831 (N_3831,N_3111,N_3016);
nor U3832 (N_3832,N_3413,N_3261);
nor U3833 (N_3833,N_3010,N_3472);
or U3834 (N_3834,N_3216,N_3371);
and U3835 (N_3835,N_3392,N_3181);
and U3836 (N_3836,N_3448,N_3075);
and U3837 (N_3837,N_3010,N_3118);
or U3838 (N_3838,N_3202,N_3079);
and U3839 (N_3839,N_3107,N_3126);
nand U3840 (N_3840,N_3254,N_3117);
and U3841 (N_3841,N_3066,N_3424);
nor U3842 (N_3842,N_3482,N_3047);
or U3843 (N_3843,N_3287,N_3005);
or U3844 (N_3844,N_3273,N_3073);
or U3845 (N_3845,N_3186,N_3266);
or U3846 (N_3846,N_3326,N_3187);
or U3847 (N_3847,N_3239,N_3479);
or U3848 (N_3848,N_3181,N_3371);
and U3849 (N_3849,N_3341,N_3063);
and U3850 (N_3850,N_3027,N_3209);
or U3851 (N_3851,N_3015,N_3056);
nand U3852 (N_3852,N_3187,N_3110);
nor U3853 (N_3853,N_3222,N_3285);
or U3854 (N_3854,N_3362,N_3325);
xor U3855 (N_3855,N_3084,N_3260);
nor U3856 (N_3856,N_3089,N_3121);
nand U3857 (N_3857,N_3090,N_3056);
nand U3858 (N_3858,N_3311,N_3476);
nor U3859 (N_3859,N_3392,N_3257);
and U3860 (N_3860,N_3325,N_3277);
or U3861 (N_3861,N_3102,N_3496);
or U3862 (N_3862,N_3374,N_3422);
nand U3863 (N_3863,N_3157,N_3069);
nand U3864 (N_3864,N_3035,N_3045);
and U3865 (N_3865,N_3346,N_3229);
or U3866 (N_3866,N_3030,N_3150);
nand U3867 (N_3867,N_3139,N_3172);
and U3868 (N_3868,N_3055,N_3491);
nor U3869 (N_3869,N_3009,N_3148);
nand U3870 (N_3870,N_3345,N_3482);
and U3871 (N_3871,N_3193,N_3305);
nand U3872 (N_3872,N_3151,N_3215);
or U3873 (N_3873,N_3067,N_3108);
or U3874 (N_3874,N_3431,N_3093);
or U3875 (N_3875,N_3179,N_3078);
nand U3876 (N_3876,N_3360,N_3260);
nand U3877 (N_3877,N_3390,N_3417);
and U3878 (N_3878,N_3360,N_3409);
nand U3879 (N_3879,N_3467,N_3035);
nor U3880 (N_3880,N_3167,N_3311);
nor U3881 (N_3881,N_3284,N_3227);
and U3882 (N_3882,N_3324,N_3074);
or U3883 (N_3883,N_3089,N_3373);
nor U3884 (N_3884,N_3243,N_3197);
nor U3885 (N_3885,N_3249,N_3089);
and U3886 (N_3886,N_3128,N_3024);
and U3887 (N_3887,N_3481,N_3499);
or U3888 (N_3888,N_3261,N_3490);
or U3889 (N_3889,N_3310,N_3288);
nor U3890 (N_3890,N_3261,N_3246);
xnor U3891 (N_3891,N_3171,N_3054);
or U3892 (N_3892,N_3099,N_3424);
nand U3893 (N_3893,N_3354,N_3223);
and U3894 (N_3894,N_3145,N_3237);
or U3895 (N_3895,N_3173,N_3391);
nor U3896 (N_3896,N_3265,N_3277);
or U3897 (N_3897,N_3195,N_3149);
or U3898 (N_3898,N_3256,N_3249);
and U3899 (N_3899,N_3145,N_3320);
or U3900 (N_3900,N_3192,N_3372);
nand U3901 (N_3901,N_3199,N_3114);
or U3902 (N_3902,N_3004,N_3227);
or U3903 (N_3903,N_3121,N_3247);
or U3904 (N_3904,N_3179,N_3339);
nor U3905 (N_3905,N_3023,N_3085);
nand U3906 (N_3906,N_3182,N_3268);
and U3907 (N_3907,N_3043,N_3004);
or U3908 (N_3908,N_3288,N_3028);
xor U3909 (N_3909,N_3392,N_3401);
or U3910 (N_3910,N_3397,N_3290);
and U3911 (N_3911,N_3478,N_3195);
or U3912 (N_3912,N_3403,N_3277);
and U3913 (N_3913,N_3457,N_3207);
nor U3914 (N_3914,N_3415,N_3465);
nand U3915 (N_3915,N_3277,N_3012);
nand U3916 (N_3916,N_3329,N_3215);
or U3917 (N_3917,N_3115,N_3099);
nand U3918 (N_3918,N_3198,N_3032);
and U3919 (N_3919,N_3012,N_3137);
xnor U3920 (N_3920,N_3477,N_3092);
nor U3921 (N_3921,N_3258,N_3401);
and U3922 (N_3922,N_3452,N_3229);
and U3923 (N_3923,N_3096,N_3249);
nand U3924 (N_3924,N_3054,N_3063);
and U3925 (N_3925,N_3292,N_3197);
nand U3926 (N_3926,N_3486,N_3301);
nand U3927 (N_3927,N_3001,N_3145);
nand U3928 (N_3928,N_3037,N_3021);
or U3929 (N_3929,N_3410,N_3454);
nor U3930 (N_3930,N_3467,N_3442);
nor U3931 (N_3931,N_3441,N_3113);
and U3932 (N_3932,N_3112,N_3274);
or U3933 (N_3933,N_3094,N_3209);
nand U3934 (N_3934,N_3348,N_3008);
and U3935 (N_3935,N_3204,N_3237);
or U3936 (N_3936,N_3313,N_3212);
and U3937 (N_3937,N_3094,N_3044);
or U3938 (N_3938,N_3179,N_3026);
xnor U3939 (N_3939,N_3055,N_3310);
and U3940 (N_3940,N_3045,N_3396);
or U3941 (N_3941,N_3194,N_3174);
xor U3942 (N_3942,N_3190,N_3005);
or U3943 (N_3943,N_3487,N_3213);
and U3944 (N_3944,N_3111,N_3440);
nor U3945 (N_3945,N_3387,N_3226);
and U3946 (N_3946,N_3084,N_3329);
or U3947 (N_3947,N_3455,N_3493);
or U3948 (N_3948,N_3040,N_3212);
or U3949 (N_3949,N_3342,N_3363);
nand U3950 (N_3950,N_3335,N_3128);
nand U3951 (N_3951,N_3069,N_3307);
nor U3952 (N_3952,N_3383,N_3016);
nor U3953 (N_3953,N_3411,N_3095);
nor U3954 (N_3954,N_3043,N_3089);
nor U3955 (N_3955,N_3009,N_3359);
nand U3956 (N_3956,N_3320,N_3296);
nand U3957 (N_3957,N_3382,N_3191);
nand U3958 (N_3958,N_3390,N_3362);
or U3959 (N_3959,N_3116,N_3287);
or U3960 (N_3960,N_3106,N_3155);
nor U3961 (N_3961,N_3351,N_3250);
or U3962 (N_3962,N_3359,N_3417);
or U3963 (N_3963,N_3420,N_3238);
and U3964 (N_3964,N_3475,N_3441);
nand U3965 (N_3965,N_3481,N_3138);
or U3966 (N_3966,N_3473,N_3470);
nand U3967 (N_3967,N_3170,N_3254);
xnor U3968 (N_3968,N_3484,N_3280);
nor U3969 (N_3969,N_3325,N_3215);
or U3970 (N_3970,N_3364,N_3211);
or U3971 (N_3971,N_3008,N_3369);
nand U3972 (N_3972,N_3463,N_3069);
and U3973 (N_3973,N_3242,N_3434);
or U3974 (N_3974,N_3482,N_3453);
nor U3975 (N_3975,N_3164,N_3030);
nand U3976 (N_3976,N_3474,N_3073);
or U3977 (N_3977,N_3312,N_3224);
nand U3978 (N_3978,N_3499,N_3452);
nand U3979 (N_3979,N_3265,N_3159);
or U3980 (N_3980,N_3464,N_3465);
nand U3981 (N_3981,N_3255,N_3345);
nand U3982 (N_3982,N_3235,N_3360);
xor U3983 (N_3983,N_3344,N_3347);
and U3984 (N_3984,N_3280,N_3069);
and U3985 (N_3985,N_3385,N_3228);
and U3986 (N_3986,N_3333,N_3415);
or U3987 (N_3987,N_3391,N_3177);
nand U3988 (N_3988,N_3016,N_3480);
nand U3989 (N_3989,N_3048,N_3367);
nor U3990 (N_3990,N_3352,N_3349);
nor U3991 (N_3991,N_3137,N_3472);
and U3992 (N_3992,N_3273,N_3217);
nor U3993 (N_3993,N_3208,N_3255);
or U3994 (N_3994,N_3325,N_3145);
nor U3995 (N_3995,N_3204,N_3008);
nand U3996 (N_3996,N_3048,N_3267);
and U3997 (N_3997,N_3235,N_3191);
nor U3998 (N_3998,N_3301,N_3448);
and U3999 (N_3999,N_3164,N_3429);
or U4000 (N_4000,N_3743,N_3593);
and U4001 (N_4001,N_3956,N_3837);
or U4002 (N_4002,N_3876,N_3615);
nand U4003 (N_4003,N_3985,N_3852);
or U4004 (N_4004,N_3941,N_3963);
or U4005 (N_4005,N_3730,N_3927);
nand U4006 (N_4006,N_3920,N_3755);
xor U4007 (N_4007,N_3713,N_3564);
xnor U4008 (N_4008,N_3895,N_3514);
or U4009 (N_4009,N_3558,N_3717);
and U4010 (N_4010,N_3687,N_3982);
nand U4011 (N_4011,N_3664,N_3708);
nor U4012 (N_4012,N_3691,N_3747);
and U4013 (N_4013,N_3732,N_3809);
nor U4014 (N_4014,N_3516,N_3770);
nor U4015 (N_4015,N_3517,N_3889);
nand U4016 (N_4016,N_3991,N_3614);
and U4017 (N_4017,N_3644,N_3653);
or U4018 (N_4018,N_3539,N_3825);
nor U4019 (N_4019,N_3741,N_3734);
or U4020 (N_4020,N_3648,N_3938);
and U4021 (N_4021,N_3573,N_3853);
or U4022 (N_4022,N_3598,N_3638);
or U4023 (N_4023,N_3948,N_3595);
and U4024 (N_4024,N_3946,N_3739);
or U4025 (N_4025,N_3822,N_3665);
and U4026 (N_4026,N_3900,N_3726);
nand U4027 (N_4027,N_3906,N_3523);
nor U4028 (N_4028,N_3542,N_3931);
nand U4029 (N_4029,N_3894,N_3570);
nand U4030 (N_4030,N_3702,N_3681);
nor U4031 (N_4031,N_3908,N_3675);
and U4032 (N_4032,N_3830,N_3792);
nor U4033 (N_4033,N_3879,N_3515);
or U4034 (N_4034,N_3567,N_3707);
nor U4035 (N_4035,N_3628,N_3987);
nor U4036 (N_4036,N_3738,N_3596);
nand U4037 (N_4037,N_3674,N_3538);
nand U4038 (N_4038,N_3947,N_3700);
nand U4039 (N_4039,N_3817,N_3580);
nand U4040 (N_4040,N_3623,N_3880);
nor U4041 (N_4041,N_3694,N_3582);
nor U4042 (N_4042,N_3972,N_3912);
and U4043 (N_4043,N_3609,N_3957);
and U4044 (N_4044,N_3836,N_3682);
or U4045 (N_4045,N_3866,N_3629);
and U4046 (N_4046,N_3923,N_3530);
and U4047 (N_4047,N_3806,N_3521);
or U4048 (N_4048,N_3658,N_3905);
and U4049 (N_4049,N_3603,N_3684);
and U4050 (N_4050,N_3773,N_3627);
nor U4051 (N_4051,N_3696,N_3834);
or U4052 (N_4052,N_3916,N_3630);
nor U4053 (N_4053,N_3502,N_3725);
and U4054 (N_4054,N_3529,N_3958);
nand U4055 (N_4055,N_3531,N_3996);
and U4056 (N_4056,N_3798,N_3998);
nor U4057 (N_4057,N_3796,N_3507);
and U4058 (N_4058,N_3731,N_3533);
nand U4059 (N_4059,N_3504,N_3509);
nand U4060 (N_4060,N_3970,N_3710);
or U4061 (N_4061,N_3581,N_3683);
or U4062 (N_4062,N_3760,N_3654);
and U4063 (N_4063,N_3723,N_3679);
nor U4064 (N_4064,N_3791,N_3922);
and U4065 (N_4065,N_3522,N_3569);
nor U4066 (N_4066,N_3728,N_3503);
nor U4067 (N_4067,N_3859,N_3960);
nand U4068 (N_4068,N_3804,N_3518);
and U4069 (N_4069,N_3951,N_3869);
nand U4070 (N_4070,N_3622,N_3612);
nand U4071 (N_4071,N_3877,N_3984);
or U4072 (N_4072,N_3961,N_3552);
and U4073 (N_4073,N_3608,N_3505);
nor U4074 (N_4074,N_3903,N_3875);
nand U4075 (N_4075,N_3902,N_3882);
or U4076 (N_4076,N_3867,N_3733);
nand U4077 (N_4077,N_3952,N_3950);
or U4078 (N_4078,N_3785,N_3508);
nor U4079 (N_4079,N_3568,N_3661);
nor U4080 (N_4080,N_3547,N_3692);
nand U4081 (N_4081,N_3907,N_3759);
and U4082 (N_4082,N_3635,N_3742);
or U4083 (N_4083,N_3892,N_3745);
nor U4084 (N_4084,N_3693,N_3645);
and U4085 (N_4085,N_3765,N_3964);
nor U4086 (N_4086,N_3788,N_3617);
nor U4087 (N_4087,N_3714,N_3563);
or U4088 (N_4088,N_3973,N_3962);
nand U4089 (N_4089,N_3857,N_3783);
and U4090 (N_4090,N_3851,N_3697);
and U4091 (N_4091,N_3878,N_3613);
and U4092 (N_4092,N_3959,N_3729);
nor U4093 (N_4093,N_3967,N_3914);
nand U4094 (N_4094,N_3935,N_3643);
xnor U4095 (N_4095,N_3856,N_3977);
nor U4096 (N_4096,N_3835,N_3579);
and U4097 (N_4097,N_3861,N_3858);
nand U4098 (N_4098,N_3698,N_3727);
and U4099 (N_4099,N_3764,N_3936);
nand U4100 (N_4100,N_3855,N_3775);
xor U4101 (N_4101,N_3527,N_3666);
nor U4102 (N_4102,N_3887,N_3561);
and U4103 (N_4103,N_3863,N_3715);
nand U4104 (N_4104,N_3939,N_3735);
or U4105 (N_4105,N_3757,N_3601);
and U4106 (N_4106,N_3901,N_3676);
or U4107 (N_4107,N_3979,N_3896);
or U4108 (N_4108,N_3893,N_3562);
nor U4109 (N_4109,N_3592,N_3924);
nand U4110 (N_4110,N_3736,N_3805);
nor U4111 (N_4111,N_3616,N_3821);
and U4112 (N_4112,N_3546,N_3565);
nand U4113 (N_4113,N_3662,N_3719);
and U4114 (N_4114,N_3704,N_3797);
and U4115 (N_4115,N_3810,N_3624);
or U4116 (N_4116,N_3640,N_3955);
or U4117 (N_4117,N_3911,N_3993);
nor U4118 (N_4118,N_3621,N_3776);
xnor U4119 (N_4119,N_3602,N_3583);
and U4120 (N_4120,N_3537,N_3655);
xnor U4121 (N_4121,N_3651,N_3641);
and U4122 (N_4122,N_3917,N_3652);
nand U4123 (N_4123,N_3656,N_3749);
nor U4124 (N_4124,N_3589,N_3827);
or U4125 (N_4125,N_3845,N_3812);
nand U4126 (N_4126,N_3718,N_3519);
nand U4127 (N_4127,N_3535,N_3590);
nor U4128 (N_4128,N_3820,N_3949);
nor U4129 (N_4129,N_3868,N_3918);
and U4130 (N_4130,N_3932,N_3862);
nor U4131 (N_4131,N_3545,N_3781);
or U4132 (N_4132,N_3826,N_3588);
or U4133 (N_4133,N_3680,N_3705);
or U4134 (N_4134,N_3926,N_3659);
nor U4135 (N_4135,N_3510,N_3767);
and U4136 (N_4136,N_3766,N_3511);
nor U4137 (N_4137,N_3607,N_3611);
nor U4138 (N_4138,N_3541,N_3871);
nor U4139 (N_4139,N_3793,N_3824);
nor U4140 (N_4140,N_3829,N_3799);
or U4141 (N_4141,N_3965,N_3966);
or U4142 (N_4142,N_3591,N_3904);
or U4143 (N_4143,N_3536,N_3716);
or U4144 (N_4144,N_3997,N_3572);
or U4145 (N_4145,N_3975,N_3832);
or U4146 (N_4146,N_3620,N_3689);
or U4147 (N_4147,N_3649,N_3777);
and U4148 (N_4148,N_3795,N_3823);
nand U4149 (N_4149,N_3919,N_3971);
nand U4150 (N_4150,N_3703,N_3842);
and U4151 (N_4151,N_3988,N_3873);
or U4152 (N_4152,N_3548,N_3642);
and U4153 (N_4153,N_3721,N_3699);
or U4154 (N_4154,N_3524,N_3647);
nand U4155 (N_4155,N_3898,N_3534);
xnor U4156 (N_4156,N_3610,N_3780);
or U4157 (N_4157,N_3688,N_3833);
nand U4158 (N_4158,N_3578,N_3915);
and U4159 (N_4159,N_3969,N_3650);
and U4160 (N_4160,N_3671,N_3512);
nor U4161 (N_4161,N_3670,N_3831);
nor U4162 (N_4162,N_3543,N_3800);
and U4163 (N_4163,N_3597,N_3577);
nor U4164 (N_4164,N_3992,N_3841);
nor U4165 (N_4165,N_3818,N_3778);
nor U4166 (N_4166,N_3910,N_3819);
and U4167 (N_4167,N_3594,N_3974);
xor U4168 (N_4168,N_3500,N_3934);
or U4169 (N_4169,N_3940,N_3790);
nor U4170 (N_4170,N_3928,N_3808);
or U4171 (N_4171,N_3762,N_3575);
and U4172 (N_4172,N_3706,N_3802);
nand U4173 (N_4173,N_3763,N_3753);
and U4174 (N_4174,N_3549,N_3989);
and U4175 (N_4175,N_3870,N_3978);
nor U4176 (N_4176,N_3525,N_3968);
or U4177 (N_4177,N_3712,N_3625);
and U4178 (N_4178,N_3909,N_3983);
xnor U4179 (N_4179,N_3786,N_3600);
or U4180 (N_4180,N_3605,N_3551);
nand U4181 (N_4181,N_3571,N_3618);
or U4182 (N_4182,N_3872,N_3606);
nand U4183 (N_4183,N_3854,N_3891);
nand U4184 (N_4184,N_3913,N_3690);
nand U4185 (N_4185,N_3849,N_3874);
nand U4186 (N_4186,N_3724,N_3844);
nand U4187 (N_4187,N_3555,N_3746);
nor U4188 (N_4188,N_3520,N_3540);
and U4189 (N_4189,N_3994,N_3584);
nor U4190 (N_4190,N_3669,N_3814);
nor U4191 (N_4191,N_3864,N_3758);
nand U4192 (N_4192,N_3815,N_3550);
nor U4193 (N_4193,N_3646,N_3976);
nor U4194 (N_4194,N_3890,N_3794);
nor U4195 (N_4195,N_3557,N_3981);
or U4196 (N_4196,N_3774,N_3737);
nor U4197 (N_4197,N_3803,N_3888);
nor U4198 (N_4198,N_3945,N_3772);
or U4199 (N_4199,N_3633,N_3953);
nor U4200 (N_4200,N_3840,N_3816);
nor U4201 (N_4201,N_3846,N_3779);
nand U4202 (N_4202,N_3769,N_3701);
or U4203 (N_4203,N_3672,N_3828);
nand U4204 (N_4204,N_3711,N_3513);
nor U4205 (N_4205,N_3604,N_3942);
nand U4206 (N_4206,N_3673,N_3771);
nor U4207 (N_4207,N_3752,N_3883);
nor U4208 (N_4208,N_3768,N_3990);
nand U4209 (N_4209,N_3850,N_3528);
nor U4210 (N_4210,N_3929,N_3933);
or U4211 (N_4211,N_3686,N_3709);
and U4212 (N_4212,N_3678,N_3943);
or U4213 (N_4213,N_3544,N_3986);
or U4214 (N_4214,N_3881,N_3663);
nand U4215 (N_4215,N_3576,N_3838);
nand U4216 (N_4216,N_3668,N_3637);
nor U4217 (N_4217,N_3761,N_3750);
nand U4218 (N_4218,N_3667,N_3695);
nand U4219 (N_4219,N_3501,N_3839);
xnor U4220 (N_4220,N_3574,N_3848);
and U4221 (N_4221,N_3722,N_3789);
nand U4222 (N_4222,N_3925,N_3754);
nor U4223 (N_4223,N_3657,N_3744);
nand U4224 (N_4224,N_3532,N_3865);
or U4225 (N_4225,N_3599,N_3677);
nor U4226 (N_4226,N_3885,N_3619);
nand U4227 (N_4227,N_3811,N_3566);
nand U4228 (N_4228,N_3553,N_3585);
nor U4229 (N_4229,N_3751,N_3782);
nor U4230 (N_4230,N_3807,N_3899);
and U4231 (N_4231,N_3632,N_3886);
nand U4232 (N_4232,N_3685,N_3884);
nor U4233 (N_4233,N_3980,N_3860);
nor U4234 (N_4234,N_3660,N_3847);
xor U4235 (N_4235,N_3526,N_3801);
nand U4236 (N_4236,N_3999,N_3897);
or U4237 (N_4237,N_3756,N_3740);
nand U4238 (N_4238,N_3636,N_3944);
and U4239 (N_4239,N_3843,N_3626);
nand U4240 (N_4240,N_3586,N_3559);
and U4241 (N_4241,N_3937,N_3634);
nor U4242 (N_4242,N_3930,N_3639);
nor U4243 (N_4243,N_3921,N_3787);
nor U4244 (N_4244,N_3720,N_3995);
nor U4245 (N_4245,N_3560,N_3587);
nor U4246 (N_4246,N_3556,N_3748);
or U4247 (N_4247,N_3554,N_3954);
xor U4248 (N_4248,N_3631,N_3813);
nor U4249 (N_4249,N_3506,N_3784);
nand U4250 (N_4250,N_3877,N_3644);
or U4251 (N_4251,N_3616,N_3594);
or U4252 (N_4252,N_3599,N_3925);
nor U4253 (N_4253,N_3822,N_3599);
nor U4254 (N_4254,N_3911,N_3856);
nor U4255 (N_4255,N_3738,N_3750);
nor U4256 (N_4256,N_3823,N_3507);
nand U4257 (N_4257,N_3762,N_3885);
and U4258 (N_4258,N_3865,N_3933);
nand U4259 (N_4259,N_3628,N_3860);
or U4260 (N_4260,N_3831,N_3609);
or U4261 (N_4261,N_3550,N_3899);
and U4262 (N_4262,N_3727,N_3922);
nand U4263 (N_4263,N_3503,N_3552);
nand U4264 (N_4264,N_3892,N_3754);
and U4265 (N_4265,N_3614,N_3746);
or U4266 (N_4266,N_3572,N_3924);
and U4267 (N_4267,N_3846,N_3823);
and U4268 (N_4268,N_3657,N_3950);
or U4269 (N_4269,N_3697,N_3616);
nor U4270 (N_4270,N_3539,N_3817);
and U4271 (N_4271,N_3833,N_3776);
nand U4272 (N_4272,N_3540,N_3808);
nand U4273 (N_4273,N_3985,N_3695);
nor U4274 (N_4274,N_3530,N_3960);
and U4275 (N_4275,N_3917,N_3763);
and U4276 (N_4276,N_3981,N_3545);
nand U4277 (N_4277,N_3648,N_3937);
nor U4278 (N_4278,N_3984,N_3789);
and U4279 (N_4279,N_3506,N_3642);
or U4280 (N_4280,N_3645,N_3701);
nor U4281 (N_4281,N_3628,N_3767);
and U4282 (N_4282,N_3768,N_3506);
nor U4283 (N_4283,N_3916,N_3872);
nor U4284 (N_4284,N_3998,N_3841);
nor U4285 (N_4285,N_3943,N_3702);
nor U4286 (N_4286,N_3515,N_3961);
and U4287 (N_4287,N_3788,N_3860);
nor U4288 (N_4288,N_3889,N_3808);
and U4289 (N_4289,N_3733,N_3790);
and U4290 (N_4290,N_3660,N_3938);
nand U4291 (N_4291,N_3666,N_3975);
nor U4292 (N_4292,N_3757,N_3934);
nand U4293 (N_4293,N_3552,N_3625);
nor U4294 (N_4294,N_3538,N_3648);
nor U4295 (N_4295,N_3550,N_3628);
nand U4296 (N_4296,N_3741,N_3645);
nand U4297 (N_4297,N_3771,N_3763);
and U4298 (N_4298,N_3753,N_3711);
and U4299 (N_4299,N_3952,N_3589);
nor U4300 (N_4300,N_3629,N_3662);
or U4301 (N_4301,N_3538,N_3726);
nor U4302 (N_4302,N_3976,N_3877);
or U4303 (N_4303,N_3825,N_3637);
nor U4304 (N_4304,N_3841,N_3931);
or U4305 (N_4305,N_3585,N_3719);
nor U4306 (N_4306,N_3587,N_3992);
nor U4307 (N_4307,N_3637,N_3994);
nand U4308 (N_4308,N_3857,N_3547);
and U4309 (N_4309,N_3923,N_3793);
and U4310 (N_4310,N_3723,N_3952);
or U4311 (N_4311,N_3636,N_3727);
and U4312 (N_4312,N_3702,N_3507);
xor U4313 (N_4313,N_3743,N_3779);
nor U4314 (N_4314,N_3618,N_3964);
nand U4315 (N_4315,N_3567,N_3506);
nand U4316 (N_4316,N_3858,N_3916);
nor U4317 (N_4317,N_3970,N_3671);
nor U4318 (N_4318,N_3941,N_3922);
nand U4319 (N_4319,N_3586,N_3642);
or U4320 (N_4320,N_3715,N_3644);
and U4321 (N_4321,N_3520,N_3654);
or U4322 (N_4322,N_3739,N_3738);
or U4323 (N_4323,N_3972,N_3854);
nor U4324 (N_4324,N_3770,N_3793);
or U4325 (N_4325,N_3914,N_3854);
or U4326 (N_4326,N_3533,N_3931);
nor U4327 (N_4327,N_3739,N_3956);
and U4328 (N_4328,N_3590,N_3827);
or U4329 (N_4329,N_3836,N_3878);
or U4330 (N_4330,N_3903,N_3823);
and U4331 (N_4331,N_3938,N_3711);
nand U4332 (N_4332,N_3863,N_3735);
nor U4333 (N_4333,N_3562,N_3517);
or U4334 (N_4334,N_3744,N_3980);
and U4335 (N_4335,N_3933,N_3512);
or U4336 (N_4336,N_3963,N_3720);
and U4337 (N_4337,N_3718,N_3924);
nand U4338 (N_4338,N_3809,N_3850);
nor U4339 (N_4339,N_3729,N_3539);
and U4340 (N_4340,N_3636,N_3873);
or U4341 (N_4341,N_3898,N_3859);
nand U4342 (N_4342,N_3667,N_3739);
and U4343 (N_4343,N_3794,N_3587);
or U4344 (N_4344,N_3889,N_3750);
or U4345 (N_4345,N_3951,N_3618);
nand U4346 (N_4346,N_3869,N_3571);
xor U4347 (N_4347,N_3544,N_3614);
or U4348 (N_4348,N_3942,N_3874);
nor U4349 (N_4349,N_3677,N_3766);
nand U4350 (N_4350,N_3667,N_3559);
nand U4351 (N_4351,N_3843,N_3914);
nand U4352 (N_4352,N_3907,N_3851);
or U4353 (N_4353,N_3924,N_3983);
xor U4354 (N_4354,N_3760,N_3848);
or U4355 (N_4355,N_3648,N_3819);
and U4356 (N_4356,N_3544,N_3824);
or U4357 (N_4357,N_3802,N_3784);
nand U4358 (N_4358,N_3893,N_3681);
and U4359 (N_4359,N_3818,N_3954);
nand U4360 (N_4360,N_3890,N_3651);
nor U4361 (N_4361,N_3880,N_3837);
nor U4362 (N_4362,N_3947,N_3626);
or U4363 (N_4363,N_3967,N_3582);
or U4364 (N_4364,N_3987,N_3876);
nor U4365 (N_4365,N_3600,N_3673);
or U4366 (N_4366,N_3743,N_3777);
nand U4367 (N_4367,N_3590,N_3751);
nand U4368 (N_4368,N_3677,N_3737);
nor U4369 (N_4369,N_3814,N_3722);
and U4370 (N_4370,N_3500,N_3840);
nor U4371 (N_4371,N_3680,N_3520);
nor U4372 (N_4372,N_3517,N_3882);
or U4373 (N_4373,N_3705,N_3992);
and U4374 (N_4374,N_3589,N_3804);
nand U4375 (N_4375,N_3977,N_3708);
or U4376 (N_4376,N_3855,N_3917);
nor U4377 (N_4377,N_3703,N_3695);
or U4378 (N_4378,N_3591,N_3905);
nor U4379 (N_4379,N_3843,N_3644);
or U4380 (N_4380,N_3591,N_3722);
or U4381 (N_4381,N_3575,N_3615);
nand U4382 (N_4382,N_3740,N_3609);
and U4383 (N_4383,N_3814,N_3510);
xnor U4384 (N_4384,N_3778,N_3982);
or U4385 (N_4385,N_3683,N_3585);
nand U4386 (N_4386,N_3995,N_3606);
nand U4387 (N_4387,N_3932,N_3504);
xnor U4388 (N_4388,N_3997,N_3779);
and U4389 (N_4389,N_3717,N_3972);
nor U4390 (N_4390,N_3841,N_3684);
and U4391 (N_4391,N_3853,N_3640);
xnor U4392 (N_4392,N_3715,N_3948);
nor U4393 (N_4393,N_3646,N_3675);
and U4394 (N_4394,N_3672,N_3912);
nand U4395 (N_4395,N_3714,N_3851);
and U4396 (N_4396,N_3740,N_3554);
and U4397 (N_4397,N_3567,N_3730);
nor U4398 (N_4398,N_3739,N_3553);
nand U4399 (N_4399,N_3897,N_3961);
or U4400 (N_4400,N_3639,N_3594);
nor U4401 (N_4401,N_3954,N_3627);
nor U4402 (N_4402,N_3965,N_3723);
or U4403 (N_4403,N_3678,N_3757);
nor U4404 (N_4404,N_3627,N_3572);
or U4405 (N_4405,N_3816,N_3753);
nand U4406 (N_4406,N_3502,N_3547);
or U4407 (N_4407,N_3867,N_3741);
nand U4408 (N_4408,N_3840,N_3720);
nand U4409 (N_4409,N_3732,N_3682);
and U4410 (N_4410,N_3583,N_3741);
nor U4411 (N_4411,N_3663,N_3500);
nor U4412 (N_4412,N_3603,N_3549);
xor U4413 (N_4413,N_3512,N_3996);
nand U4414 (N_4414,N_3921,N_3915);
and U4415 (N_4415,N_3587,N_3509);
and U4416 (N_4416,N_3622,N_3693);
nand U4417 (N_4417,N_3921,N_3686);
nand U4418 (N_4418,N_3850,N_3636);
and U4419 (N_4419,N_3679,N_3813);
and U4420 (N_4420,N_3531,N_3940);
or U4421 (N_4421,N_3988,N_3700);
nand U4422 (N_4422,N_3558,N_3534);
and U4423 (N_4423,N_3591,N_3600);
and U4424 (N_4424,N_3858,N_3897);
nand U4425 (N_4425,N_3648,N_3850);
nor U4426 (N_4426,N_3534,N_3796);
nor U4427 (N_4427,N_3865,N_3837);
xnor U4428 (N_4428,N_3510,N_3764);
or U4429 (N_4429,N_3965,N_3809);
nor U4430 (N_4430,N_3769,N_3866);
and U4431 (N_4431,N_3832,N_3851);
or U4432 (N_4432,N_3750,N_3634);
nor U4433 (N_4433,N_3645,N_3941);
nand U4434 (N_4434,N_3726,N_3717);
or U4435 (N_4435,N_3826,N_3512);
nand U4436 (N_4436,N_3761,N_3648);
or U4437 (N_4437,N_3989,N_3935);
and U4438 (N_4438,N_3626,N_3751);
and U4439 (N_4439,N_3719,N_3760);
nand U4440 (N_4440,N_3835,N_3635);
and U4441 (N_4441,N_3552,N_3576);
or U4442 (N_4442,N_3527,N_3960);
or U4443 (N_4443,N_3521,N_3972);
and U4444 (N_4444,N_3714,N_3757);
nand U4445 (N_4445,N_3562,N_3707);
or U4446 (N_4446,N_3796,N_3814);
xnor U4447 (N_4447,N_3943,N_3608);
and U4448 (N_4448,N_3547,N_3881);
and U4449 (N_4449,N_3578,N_3862);
nand U4450 (N_4450,N_3994,N_3806);
or U4451 (N_4451,N_3833,N_3790);
nor U4452 (N_4452,N_3654,N_3688);
or U4453 (N_4453,N_3592,N_3931);
nor U4454 (N_4454,N_3863,N_3818);
nor U4455 (N_4455,N_3671,N_3966);
nor U4456 (N_4456,N_3972,N_3631);
or U4457 (N_4457,N_3989,N_3878);
and U4458 (N_4458,N_3769,N_3958);
nand U4459 (N_4459,N_3546,N_3830);
nor U4460 (N_4460,N_3795,N_3553);
nor U4461 (N_4461,N_3781,N_3778);
xnor U4462 (N_4462,N_3679,N_3838);
nand U4463 (N_4463,N_3548,N_3679);
nand U4464 (N_4464,N_3598,N_3829);
xor U4465 (N_4465,N_3700,N_3981);
or U4466 (N_4466,N_3649,N_3783);
nand U4467 (N_4467,N_3760,N_3944);
or U4468 (N_4468,N_3906,N_3943);
nor U4469 (N_4469,N_3642,N_3747);
and U4470 (N_4470,N_3696,N_3706);
xnor U4471 (N_4471,N_3887,N_3648);
or U4472 (N_4472,N_3686,N_3717);
nand U4473 (N_4473,N_3532,N_3955);
nand U4474 (N_4474,N_3968,N_3959);
or U4475 (N_4475,N_3633,N_3619);
and U4476 (N_4476,N_3637,N_3787);
nand U4477 (N_4477,N_3951,N_3579);
nor U4478 (N_4478,N_3533,N_3729);
nor U4479 (N_4479,N_3842,N_3883);
or U4480 (N_4480,N_3864,N_3730);
and U4481 (N_4481,N_3833,N_3585);
nand U4482 (N_4482,N_3657,N_3689);
xor U4483 (N_4483,N_3568,N_3556);
or U4484 (N_4484,N_3908,N_3709);
nand U4485 (N_4485,N_3649,N_3712);
or U4486 (N_4486,N_3750,N_3739);
nor U4487 (N_4487,N_3543,N_3901);
nor U4488 (N_4488,N_3797,N_3546);
nor U4489 (N_4489,N_3797,N_3979);
or U4490 (N_4490,N_3980,N_3624);
nand U4491 (N_4491,N_3692,N_3651);
nor U4492 (N_4492,N_3939,N_3973);
and U4493 (N_4493,N_3938,N_3996);
or U4494 (N_4494,N_3566,N_3591);
nand U4495 (N_4495,N_3833,N_3574);
nand U4496 (N_4496,N_3648,N_3514);
nor U4497 (N_4497,N_3882,N_3996);
nand U4498 (N_4498,N_3945,N_3563);
nor U4499 (N_4499,N_3862,N_3518);
or U4500 (N_4500,N_4427,N_4261);
and U4501 (N_4501,N_4316,N_4010);
or U4502 (N_4502,N_4410,N_4407);
or U4503 (N_4503,N_4092,N_4201);
nand U4504 (N_4504,N_4298,N_4174);
and U4505 (N_4505,N_4441,N_4205);
or U4506 (N_4506,N_4465,N_4428);
and U4507 (N_4507,N_4045,N_4227);
and U4508 (N_4508,N_4021,N_4145);
or U4509 (N_4509,N_4479,N_4161);
and U4510 (N_4510,N_4393,N_4443);
nand U4511 (N_4511,N_4209,N_4102);
and U4512 (N_4512,N_4058,N_4402);
xnor U4513 (N_4513,N_4116,N_4474);
xor U4514 (N_4514,N_4398,N_4198);
or U4515 (N_4515,N_4421,N_4213);
or U4516 (N_4516,N_4403,N_4275);
nor U4517 (N_4517,N_4446,N_4311);
nand U4518 (N_4518,N_4222,N_4260);
nand U4519 (N_4519,N_4018,N_4169);
and U4520 (N_4520,N_4130,N_4050);
nor U4521 (N_4521,N_4158,N_4162);
nor U4522 (N_4522,N_4252,N_4131);
nor U4523 (N_4523,N_4194,N_4476);
or U4524 (N_4524,N_4293,N_4345);
nor U4525 (N_4525,N_4376,N_4342);
or U4526 (N_4526,N_4433,N_4333);
nor U4527 (N_4527,N_4085,N_4070);
nand U4528 (N_4528,N_4218,N_4394);
nand U4529 (N_4529,N_4464,N_4000);
nand U4530 (N_4530,N_4312,N_4334);
or U4531 (N_4531,N_4250,N_4041);
and U4532 (N_4532,N_4240,N_4196);
xor U4533 (N_4533,N_4432,N_4297);
xor U4534 (N_4534,N_4079,N_4255);
and U4535 (N_4535,N_4365,N_4165);
nor U4536 (N_4536,N_4272,N_4224);
or U4537 (N_4537,N_4253,N_4192);
or U4538 (N_4538,N_4239,N_4026);
nand U4539 (N_4539,N_4061,N_4400);
and U4540 (N_4540,N_4324,N_4491);
nand U4541 (N_4541,N_4246,N_4495);
nand U4542 (N_4542,N_4121,N_4448);
nand U4543 (N_4543,N_4177,N_4258);
and U4544 (N_4544,N_4069,N_4451);
and U4545 (N_4545,N_4294,N_4105);
or U4546 (N_4546,N_4313,N_4133);
and U4547 (N_4547,N_4020,N_4355);
nor U4548 (N_4548,N_4319,N_4278);
or U4549 (N_4549,N_4389,N_4339);
or U4550 (N_4550,N_4125,N_4004);
nor U4551 (N_4551,N_4099,N_4093);
and U4552 (N_4552,N_4435,N_4126);
and U4553 (N_4553,N_4309,N_4470);
and U4554 (N_4554,N_4195,N_4122);
nand U4555 (N_4555,N_4152,N_4219);
and U4556 (N_4556,N_4191,N_4181);
nand U4557 (N_4557,N_4331,N_4039);
and U4558 (N_4558,N_4285,N_4097);
nor U4559 (N_4559,N_4327,N_4426);
nor U4560 (N_4560,N_4414,N_4193);
nor U4561 (N_4561,N_4247,N_4006);
or U4562 (N_4562,N_4024,N_4053);
and U4563 (N_4563,N_4211,N_4153);
nor U4564 (N_4564,N_4361,N_4086);
nand U4565 (N_4565,N_4498,N_4462);
nor U4566 (N_4566,N_4387,N_4112);
nor U4567 (N_4567,N_4235,N_4134);
nor U4568 (N_4568,N_4080,N_4359);
nand U4569 (N_4569,N_4005,N_4371);
nand U4570 (N_4570,N_4489,N_4088);
or U4571 (N_4571,N_4439,N_4372);
nand U4572 (N_4572,N_4042,N_4067);
and U4573 (N_4573,N_4274,N_4008);
nand U4574 (N_4574,N_4496,N_4185);
nor U4575 (N_4575,N_4416,N_4481);
nor U4576 (N_4576,N_4472,N_4335);
and U4577 (N_4577,N_4332,N_4019);
and U4578 (N_4578,N_4111,N_4109);
nand U4579 (N_4579,N_4082,N_4175);
and U4580 (N_4580,N_4392,N_4492);
or U4581 (N_4581,N_4485,N_4017);
nor U4582 (N_4582,N_4031,N_4113);
and U4583 (N_4583,N_4475,N_4138);
or U4584 (N_4584,N_4388,N_4100);
and U4585 (N_4585,N_4302,N_4156);
and U4586 (N_4586,N_4373,N_4210);
nand U4587 (N_4587,N_4101,N_4207);
nand U4588 (N_4588,N_4199,N_4282);
nor U4589 (N_4589,N_4450,N_4442);
nand U4590 (N_4590,N_4150,N_4089);
or U4591 (N_4591,N_4187,N_4007);
nor U4592 (N_4592,N_4379,N_4328);
or U4593 (N_4593,N_4159,N_4283);
nor U4594 (N_4594,N_4351,N_4396);
nor U4595 (N_4595,N_4065,N_4486);
or U4596 (N_4596,N_4103,N_4415);
nand U4597 (N_4597,N_4461,N_4182);
nand U4598 (N_4598,N_4487,N_4043);
and U4599 (N_4599,N_4230,N_4363);
nand U4600 (N_4600,N_4269,N_4466);
nor U4601 (N_4601,N_4108,N_4300);
nand U4602 (N_4602,N_4076,N_4027);
nor U4603 (N_4603,N_4323,N_4494);
nand U4604 (N_4604,N_4074,N_4425);
or U4605 (N_4605,N_4368,N_4289);
nor U4606 (N_4606,N_4242,N_4378);
and U4607 (N_4607,N_4263,N_4136);
nand U4608 (N_4608,N_4090,N_4436);
and U4609 (N_4609,N_4059,N_4304);
nor U4610 (N_4610,N_4038,N_4216);
nor U4611 (N_4611,N_4401,N_4110);
or U4612 (N_4612,N_4455,N_4452);
nand U4613 (N_4613,N_4095,N_4214);
nor U4614 (N_4614,N_4064,N_4276);
nor U4615 (N_4615,N_4154,N_4062);
nor U4616 (N_4616,N_4399,N_4155);
nand U4617 (N_4617,N_4279,N_4003);
and U4618 (N_4618,N_4030,N_4139);
or U4619 (N_4619,N_4423,N_4029);
or U4620 (N_4620,N_4066,N_4167);
nand U4621 (N_4621,N_4237,N_4320);
nand U4622 (N_4622,N_4340,N_4457);
and U4623 (N_4623,N_4262,N_4128);
nor U4624 (N_4624,N_4002,N_4215);
and U4625 (N_4625,N_4160,N_4186);
nor U4626 (N_4626,N_4197,N_4084);
or U4627 (N_4627,N_4094,N_4437);
nor U4628 (N_4628,N_4073,N_4206);
nor U4629 (N_4629,N_4225,N_4056);
and U4630 (N_4630,N_4106,N_4364);
and U4631 (N_4631,N_4404,N_4083);
nor U4632 (N_4632,N_4163,N_4183);
nand U4633 (N_4633,N_4232,N_4135);
nor U4634 (N_4634,N_4411,N_4001);
nor U4635 (N_4635,N_4200,N_4395);
nor U4636 (N_4636,N_4129,N_4023);
xnor U4637 (N_4637,N_4418,N_4347);
nand U4638 (N_4638,N_4249,N_4308);
nor U4639 (N_4639,N_4238,N_4391);
and U4640 (N_4640,N_4422,N_4490);
or U4641 (N_4641,N_4132,N_4348);
or U4642 (N_4642,N_4384,N_4497);
nand U4643 (N_4643,N_4463,N_4322);
and U4644 (N_4644,N_4284,N_4413);
and U4645 (N_4645,N_4321,N_4499);
and U4646 (N_4646,N_4028,N_4458);
and U4647 (N_4647,N_4137,N_4176);
nor U4648 (N_4648,N_4016,N_4068);
or U4649 (N_4649,N_4075,N_4114);
and U4650 (N_4650,N_4374,N_4014);
or U4651 (N_4651,N_4420,N_4078);
or U4652 (N_4652,N_4296,N_4180);
nand U4653 (N_4653,N_4119,N_4344);
nand U4654 (N_4654,N_4254,N_4234);
nand U4655 (N_4655,N_4170,N_4318);
and U4656 (N_4656,N_4358,N_4115);
and U4657 (N_4657,N_4350,N_4049);
nand U4658 (N_4658,N_4330,N_4229);
and U4659 (N_4659,N_4051,N_4190);
nor U4660 (N_4660,N_4143,N_4098);
or U4661 (N_4661,N_4173,N_4168);
or U4662 (N_4662,N_4142,N_4375);
or U4663 (N_4663,N_4047,N_4248);
nor U4664 (N_4664,N_4469,N_4268);
and U4665 (N_4665,N_4157,N_4251);
nand U4666 (N_4666,N_4013,N_4104);
nand U4667 (N_4667,N_4273,N_4397);
nand U4668 (N_4668,N_4341,N_4048);
or U4669 (N_4669,N_4301,N_4203);
nand U4670 (N_4670,N_4337,N_4406);
or U4671 (N_4671,N_4315,N_4245);
nand U4672 (N_4672,N_4453,N_4354);
nor U4673 (N_4673,N_4149,N_4267);
xnor U4674 (N_4674,N_4178,N_4317);
nor U4675 (N_4675,N_4025,N_4015);
and U4676 (N_4676,N_4424,N_4447);
or U4677 (N_4677,N_4270,N_4360);
or U4678 (N_4678,N_4381,N_4459);
and U4679 (N_4679,N_4338,N_4184);
or U4680 (N_4680,N_4471,N_4383);
or U4681 (N_4681,N_4012,N_4046);
nor U4682 (N_4682,N_4265,N_4390);
nor U4683 (N_4683,N_4357,N_4478);
nand U4684 (N_4684,N_4223,N_4292);
nor U4685 (N_4685,N_4366,N_4009);
nand U4686 (N_4686,N_4440,N_4037);
nor U4687 (N_4687,N_4431,N_4445);
or U4688 (N_4688,N_4438,N_4473);
nand U4689 (N_4689,N_4204,N_4164);
or U4690 (N_4690,N_4266,N_4054);
nor U4691 (N_4691,N_4052,N_4057);
nand U4692 (N_4692,N_4419,N_4456);
nand U4693 (N_4693,N_4291,N_4022);
or U4694 (N_4694,N_4483,N_4107);
nor U4695 (N_4695,N_4236,N_4343);
nor U4696 (N_4696,N_4124,N_4148);
nand U4697 (N_4697,N_4179,N_4352);
nand U4698 (N_4698,N_4325,N_4349);
or U4699 (N_4699,N_4123,N_4264);
and U4700 (N_4700,N_4417,N_4329);
nor U4701 (N_4701,N_4141,N_4172);
or U4702 (N_4702,N_4228,N_4202);
and U4703 (N_4703,N_4280,N_4147);
nor U4704 (N_4704,N_4468,N_4217);
nand U4705 (N_4705,N_4233,N_4467);
nor U4706 (N_4706,N_4336,N_4299);
nand U4707 (N_4707,N_4036,N_4034);
xor U4708 (N_4708,N_4306,N_4412);
and U4709 (N_4709,N_4288,N_4171);
nor U4710 (N_4710,N_4303,N_4281);
or U4711 (N_4711,N_4310,N_4208);
nand U4712 (N_4712,N_4409,N_4188);
or U4713 (N_4713,N_4295,N_4243);
and U4714 (N_4714,N_4408,N_4346);
nand U4715 (N_4715,N_4060,N_4480);
nor U4716 (N_4716,N_4353,N_4033);
and U4717 (N_4717,N_4449,N_4221);
nor U4718 (N_4718,N_4032,N_4189);
nand U4719 (N_4719,N_4120,N_4460);
nand U4720 (N_4720,N_4362,N_4063);
and U4721 (N_4721,N_4484,N_4151);
and U4722 (N_4722,N_4385,N_4166);
nand U4723 (N_4723,N_4146,N_4386);
and U4724 (N_4724,N_4326,N_4434);
and U4725 (N_4725,N_4244,N_4055);
nand U4726 (N_4726,N_4040,N_4127);
nor U4727 (N_4727,N_4277,N_4430);
nor U4728 (N_4728,N_4356,N_4444);
or U4729 (N_4729,N_4256,N_4096);
nor U4730 (N_4730,N_4144,N_4477);
nor U4731 (N_4731,N_4231,N_4286);
nor U4732 (N_4732,N_4482,N_4077);
xor U4733 (N_4733,N_4044,N_4377);
xnor U4734 (N_4734,N_4035,N_4380);
nor U4735 (N_4735,N_4220,N_4493);
or U4736 (N_4736,N_4117,N_4287);
nand U4737 (N_4737,N_4369,N_4305);
nand U4738 (N_4738,N_4091,N_4072);
nand U4739 (N_4739,N_4118,N_4307);
nand U4740 (N_4740,N_4454,N_4314);
nor U4741 (N_4741,N_4370,N_4087);
nor U4742 (N_4742,N_4071,N_4259);
or U4743 (N_4743,N_4382,N_4257);
and U4744 (N_4744,N_4290,N_4140);
nand U4745 (N_4745,N_4271,N_4367);
and U4746 (N_4746,N_4011,N_4241);
and U4747 (N_4747,N_4212,N_4488);
xnor U4748 (N_4748,N_4226,N_4405);
xor U4749 (N_4749,N_4081,N_4429);
nor U4750 (N_4750,N_4106,N_4400);
nand U4751 (N_4751,N_4227,N_4465);
nor U4752 (N_4752,N_4205,N_4129);
or U4753 (N_4753,N_4447,N_4076);
nor U4754 (N_4754,N_4481,N_4436);
nand U4755 (N_4755,N_4245,N_4228);
nand U4756 (N_4756,N_4155,N_4287);
nand U4757 (N_4757,N_4482,N_4214);
nand U4758 (N_4758,N_4106,N_4383);
and U4759 (N_4759,N_4192,N_4188);
and U4760 (N_4760,N_4165,N_4408);
and U4761 (N_4761,N_4100,N_4192);
and U4762 (N_4762,N_4041,N_4195);
nand U4763 (N_4763,N_4217,N_4381);
and U4764 (N_4764,N_4253,N_4310);
and U4765 (N_4765,N_4055,N_4203);
nor U4766 (N_4766,N_4290,N_4214);
nor U4767 (N_4767,N_4162,N_4251);
or U4768 (N_4768,N_4304,N_4465);
and U4769 (N_4769,N_4197,N_4105);
and U4770 (N_4770,N_4465,N_4111);
or U4771 (N_4771,N_4491,N_4023);
or U4772 (N_4772,N_4245,N_4131);
or U4773 (N_4773,N_4172,N_4437);
nor U4774 (N_4774,N_4391,N_4063);
nand U4775 (N_4775,N_4355,N_4059);
and U4776 (N_4776,N_4063,N_4361);
nand U4777 (N_4777,N_4174,N_4362);
xor U4778 (N_4778,N_4477,N_4302);
and U4779 (N_4779,N_4422,N_4355);
nand U4780 (N_4780,N_4033,N_4485);
and U4781 (N_4781,N_4215,N_4444);
nor U4782 (N_4782,N_4213,N_4135);
or U4783 (N_4783,N_4156,N_4385);
or U4784 (N_4784,N_4262,N_4047);
nor U4785 (N_4785,N_4486,N_4058);
nor U4786 (N_4786,N_4357,N_4385);
or U4787 (N_4787,N_4411,N_4068);
nor U4788 (N_4788,N_4411,N_4404);
and U4789 (N_4789,N_4449,N_4290);
nand U4790 (N_4790,N_4258,N_4221);
or U4791 (N_4791,N_4404,N_4309);
and U4792 (N_4792,N_4349,N_4418);
or U4793 (N_4793,N_4476,N_4218);
and U4794 (N_4794,N_4211,N_4366);
nand U4795 (N_4795,N_4461,N_4083);
or U4796 (N_4796,N_4185,N_4291);
and U4797 (N_4797,N_4238,N_4360);
nand U4798 (N_4798,N_4244,N_4417);
and U4799 (N_4799,N_4013,N_4371);
nand U4800 (N_4800,N_4277,N_4438);
nor U4801 (N_4801,N_4337,N_4249);
nand U4802 (N_4802,N_4042,N_4315);
or U4803 (N_4803,N_4010,N_4188);
or U4804 (N_4804,N_4344,N_4387);
nor U4805 (N_4805,N_4427,N_4011);
nand U4806 (N_4806,N_4297,N_4468);
nor U4807 (N_4807,N_4023,N_4204);
nand U4808 (N_4808,N_4083,N_4074);
nand U4809 (N_4809,N_4019,N_4070);
and U4810 (N_4810,N_4121,N_4140);
nor U4811 (N_4811,N_4391,N_4095);
nor U4812 (N_4812,N_4486,N_4070);
nand U4813 (N_4813,N_4468,N_4048);
and U4814 (N_4814,N_4081,N_4495);
or U4815 (N_4815,N_4181,N_4227);
and U4816 (N_4816,N_4271,N_4221);
nand U4817 (N_4817,N_4409,N_4272);
nor U4818 (N_4818,N_4349,N_4403);
nand U4819 (N_4819,N_4270,N_4493);
and U4820 (N_4820,N_4020,N_4407);
nor U4821 (N_4821,N_4384,N_4354);
nand U4822 (N_4822,N_4364,N_4121);
nor U4823 (N_4823,N_4169,N_4285);
or U4824 (N_4824,N_4406,N_4007);
nand U4825 (N_4825,N_4444,N_4121);
nand U4826 (N_4826,N_4217,N_4377);
or U4827 (N_4827,N_4439,N_4434);
nor U4828 (N_4828,N_4064,N_4446);
or U4829 (N_4829,N_4003,N_4061);
xor U4830 (N_4830,N_4168,N_4049);
nand U4831 (N_4831,N_4129,N_4329);
or U4832 (N_4832,N_4386,N_4462);
nor U4833 (N_4833,N_4289,N_4212);
nand U4834 (N_4834,N_4236,N_4100);
nor U4835 (N_4835,N_4473,N_4257);
and U4836 (N_4836,N_4228,N_4026);
nor U4837 (N_4837,N_4089,N_4313);
or U4838 (N_4838,N_4227,N_4078);
or U4839 (N_4839,N_4254,N_4329);
or U4840 (N_4840,N_4478,N_4259);
or U4841 (N_4841,N_4149,N_4261);
and U4842 (N_4842,N_4401,N_4349);
xnor U4843 (N_4843,N_4399,N_4367);
nand U4844 (N_4844,N_4015,N_4068);
nand U4845 (N_4845,N_4074,N_4298);
nor U4846 (N_4846,N_4483,N_4296);
nand U4847 (N_4847,N_4124,N_4257);
and U4848 (N_4848,N_4320,N_4367);
nor U4849 (N_4849,N_4069,N_4194);
nand U4850 (N_4850,N_4242,N_4339);
nor U4851 (N_4851,N_4365,N_4382);
nand U4852 (N_4852,N_4029,N_4470);
nand U4853 (N_4853,N_4484,N_4104);
nand U4854 (N_4854,N_4494,N_4284);
nand U4855 (N_4855,N_4144,N_4451);
and U4856 (N_4856,N_4309,N_4455);
nand U4857 (N_4857,N_4370,N_4271);
or U4858 (N_4858,N_4098,N_4418);
or U4859 (N_4859,N_4040,N_4165);
nor U4860 (N_4860,N_4314,N_4205);
nor U4861 (N_4861,N_4478,N_4309);
or U4862 (N_4862,N_4089,N_4296);
or U4863 (N_4863,N_4376,N_4248);
and U4864 (N_4864,N_4310,N_4141);
nand U4865 (N_4865,N_4008,N_4004);
or U4866 (N_4866,N_4019,N_4091);
nand U4867 (N_4867,N_4217,N_4129);
or U4868 (N_4868,N_4325,N_4331);
and U4869 (N_4869,N_4078,N_4213);
nand U4870 (N_4870,N_4043,N_4071);
or U4871 (N_4871,N_4026,N_4065);
nand U4872 (N_4872,N_4364,N_4191);
nor U4873 (N_4873,N_4017,N_4109);
or U4874 (N_4874,N_4297,N_4062);
or U4875 (N_4875,N_4090,N_4373);
or U4876 (N_4876,N_4294,N_4393);
and U4877 (N_4877,N_4173,N_4077);
nand U4878 (N_4878,N_4338,N_4226);
or U4879 (N_4879,N_4143,N_4322);
and U4880 (N_4880,N_4192,N_4327);
and U4881 (N_4881,N_4487,N_4351);
xor U4882 (N_4882,N_4078,N_4143);
and U4883 (N_4883,N_4305,N_4292);
nor U4884 (N_4884,N_4375,N_4360);
nor U4885 (N_4885,N_4394,N_4358);
nand U4886 (N_4886,N_4461,N_4271);
and U4887 (N_4887,N_4131,N_4099);
nor U4888 (N_4888,N_4423,N_4074);
nand U4889 (N_4889,N_4259,N_4201);
and U4890 (N_4890,N_4340,N_4345);
and U4891 (N_4891,N_4006,N_4099);
or U4892 (N_4892,N_4073,N_4466);
or U4893 (N_4893,N_4097,N_4329);
nand U4894 (N_4894,N_4048,N_4030);
and U4895 (N_4895,N_4152,N_4088);
nor U4896 (N_4896,N_4236,N_4323);
nor U4897 (N_4897,N_4361,N_4029);
nand U4898 (N_4898,N_4019,N_4184);
nor U4899 (N_4899,N_4324,N_4280);
nand U4900 (N_4900,N_4056,N_4091);
or U4901 (N_4901,N_4414,N_4371);
and U4902 (N_4902,N_4476,N_4478);
and U4903 (N_4903,N_4023,N_4498);
or U4904 (N_4904,N_4186,N_4118);
xor U4905 (N_4905,N_4323,N_4130);
and U4906 (N_4906,N_4306,N_4197);
or U4907 (N_4907,N_4133,N_4457);
and U4908 (N_4908,N_4324,N_4273);
nor U4909 (N_4909,N_4048,N_4180);
and U4910 (N_4910,N_4422,N_4230);
nand U4911 (N_4911,N_4168,N_4368);
nor U4912 (N_4912,N_4458,N_4130);
or U4913 (N_4913,N_4361,N_4058);
nand U4914 (N_4914,N_4426,N_4414);
nand U4915 (N_4915,N_4436,N_4357);
or U4916 (N_4916,N_4308,N_4476);
or U4917 (N_4917,N_4312,N_4210);
or U4918 (N_4918,N_4220,N_4031);
nor U4919 (N_4919,N_4082,N_4443);
and U4920 (N_4920,N_4288,N_4398);
or U4921 (N_4921,N_4340,N_4281);
or U4922 (N_4922,N_4215,N_4246);
and U4923 (N_4923,N_4284,N_4393);
nor U4924 (N_4924,N_4283,N_4305);
nor U4925 (N_4925,N_4007,N_4464);
xnor U4926 (N_4926,N_4248,N_4405);
xnor U4927 (N_4927,N_4415,N_4255);
nor U4928 (N_4928,N_4242,N_4094);
nor U4929 (N_4929,N_4047,N_4169);
nor U4930 (N_4930,N_4139,N_4244);
xnor U4931 (N_4931,N_4391,N_4493);
and U4932 (N_4932,N_4300,N_4255);
and U4933 (N_4933,N_4046,N_4065);
or U4934 (N_4934,N_4220,N_4302);
or U4935 (N_4935,N_4496,N_4435);
nand U4936 (N_4936,N_4428,N_4396);
and U4937 (N_4937,N_4202,N_4261);
nand U4938 (N_4938,N_4455,N_4194);
nor U4939 (N_4939,N_4159,N_4338);
and U4940 (N_4940,N_4065,N_4430);
nor U4941 (N_4941,N_4083,N_4208);
nor U4942 (N_4942,N_4486,N_4484);
or U4943 (N_4943,N_4426,N_4488);
or U4944 (N_4944,N_4187,N_4276);
xor U4945 (N_4945,N_4033,N_4341);
or U4946 (N_4946,N_4433,N_4485);
or U4947 (N_4947,N_4441,N_4075);
and U4948 (N_4948,N_4321,N_4391);
nand U4949 (N_4949,N_4489,N_4106);
nor U4950 (N_4950,N_4465,N_4456);
or U4951 (N_4951,N_4449,N_4329);
nor U4952 (N_4952,N_4101,N_4469);
and U4953 (N_4953,N_4436,N_4291);
nand U4954 (N_4954,N_4076,N_4185);
or U4955 (N_4955,N_4237,N_4406);
and U4956 (N_4956,N_4165,N_4268);
nor U4957 (N_4957,N_4488,N_4190);
nor U4958 (N_4958,N_4305,N_4255);
and U4959 (N_4959,N_4281,N_4218);
nand U4960 (N_4960,N_4487,N_4175);
nand U4961 (N_4961,N_4385,N_4339);
and U4962 (N_4962,N_4312,N_4223);
nor U4963 (N_4963,N_4004,N_4422);
and U4964 (N_4964,N_4050,N_4146);
or U4965 (N_4965,N_4170,N_4358);
and U4966 (N_4966,N_4222,N_4333);
and U4967 (N_4967,N_4134,N_4249);
and U4968 (N_4968,N_4499,N_4039);
or U4969 (N_4969,N_4200,N_4485);
nand U4970 (N_4970,N_4389,N_4379);
nand U4971 (N_4971,N_4299,N_4002);
xor U4972 (N_4972,N_4317,N_4016);
or U4973 (N_4973,N_4205,N_4159);
nor U4974 (N_4974,N_4495,N_4079);
xor U4975 (N_4975,N_4009,N_4160);
nand U4976 (N_4976,N_4331,N_4086);
and U4977 (N_4977,N_4287,N_4040);
nand U4978 (N_4978,N_4170,N_4103);
nand U4979 (N_4979,N_4421,N_4447);
nand U4980 (N_4980,N_4459,N_4360);
nor U4981 (N_4981,N_4013,N_4077);
and U4982 (N_4982,N_4092,N_4436);
nor U4983 (N_4983,N_4388,N_4308);
xor U4984 (N_4984,N_4000,N_4447);
or U4985 (N_4985,N_4298,N_4348);
and U4986 (N_4986,N_4107,N_4182);
nand U4987 (N_4987,N_4302,N_4329);
and U4988 (N_4988,N_4481,N_4313);
xor U4989 (N_4989,N_4143,N_4184);
or U4990 (N_4990,N_4298,N_4270);
nand U4991 (N_4991,N_4490,N_4083);
nand U4992 (N_4992,N_4254,N_4027);
or U4993 (N_4993,N_4453,N_4062);
or U4994 (N_4994,N_4006,N_4213);
nand U4995 (N_4995,N_4438,N_4087);
nand U4996 (N_4996,N_4313,N_4016);
or U4997 (N_4997,N_4147,N_4051);
nand U4998 (N_4998,N_4382,N_4236);
nand U4999 (N_4999,N_4015,N_4221);
nor UO_0 (O_0,N_4986,N_4768);
nor UO_1 (O_1,N_4784,N_4687);
nand UO_2 (O_2,N_4971,N_4609);
nor UO_3 (O_3,N_4705,N_4693);
and UO_4 (O_4,N_4782,N_4887);
nor UO_5 (O_5,N_4763,N_4973);
or UO_6 (O_6,N_4822,N_4544);
and UO_7 (O_7,N_4649,N_4723);
and UO_8 (O_8,N_4837,N_4740);
nor UO_9 (O_9,N_4663,N_4951);
nor UO_10 (O_10,N_4580,N_4512);
nand UO_11 (O_11,N_4500,N_4890);
and UO_12 (O_12,N_4787,N_4721);
nand UO_13 (O_13,N_4853,N_4588);
nor UO_14 (O_14,N_4574,N_4965);
nor UO_15 (O_15,N_4848,N_4682);
and UO_16 (O_16,N_4896,N_4621);
nor UO_17 (O_17,N_4550,N_4689);
nand UO_18 (O_18,N_4828,N_4913);
or UO_19 (O_19,N_4888,N_4651);
nor UO_20 (O_20,N_4850,N_4586);
nor UO_21 (O_21,N_4697,N_4805);
nor UO_22 (O_22,N_4751,N_4849);
and UO_23 (O_23,N_4694,N_4708);
nand UO_24 (O_24,N_4819,N_4940);
nand UO_25 (O_25,N_4519,N_4843);
or UO_26 (O_26,N_4540,N_4629);
nor UO_27 (O_27,N_4615,N_4900);
or UO_28 (O_28,N_4801,N_4939);
nand UO_29 (O_29,N_4741,N_4765);
or UO_30 (O_30,N_4812,N_4963);
or UO_31 (O_31,N_4683,N_4882);
and UO_32 (O_32,N_4509,N_4815);
and UO_33 (O_33,N_4794,N_4792);
and UO_34 (O_34,N_4561,N_4551);
nand UO_35 (O_35,N_4781,N_4933);
nand UO_36 (O_36,N_4902,N_4710);
nand UO_37 (O_37,N_4823,N_4713);
nor UO_38 (O_38,N_4987,N_4817);
xor UO_39 (O_39,N_4614,N_4881);
nor UO_40 (O_40,N_4730,N_4516);
and UO_41 (O_41,N_4799,N_4545);
nor UO_42 (O_42,N_4922,N_4575);
nor UO_43 (O_43,N_4686,N_4994);
or UO_44 (O_44,N_4982,N_4591);
or UO_45 (O_45,N_4780,N_4759);
and UO_46 (O_46,N_4742,N_4958);
and UO_47 (O_47,N_4997,N_4993);
or UO_48 (O_48,N_4593,N_4706);
nand UO_49 (O_49,N_4852,N_4569);
nand UO_50 (O_50,N_4789,N_4797);
nand UO_51 (O_51,N_4531,N_4524);
and UO_52 (O_52,N_4967,N_4511);
or UO_53 (O_53,N_4895,N_4626);
and UO_54 (O_54,N_4908,N_4957);
and UO_55 (O_55,N_4602,N_4937);
nand UO_56 (O_56,N_4685,N_4684);
nand UO_57 (O_57,N_4860,N_4873);
nor UO_58 (O_58,N_4909,N_4899);
nand UO_59 (O_59,N_4962,N_4582);
nor UO_60 (O_60,N_4827,N_4749);
and UO_61 (O_61,N_4798,N_4875);
nor UO_62 (O_62,N_4716,N_4952);
nor UO_63 (O_63,N_4522,N_4866);
and UO_64 (O_64,N_4983,N_4622);
or UO_65 (O_65,N_4595,N_4560);
or UO_66 (O_66,N_4661,N_4979);
and UO_67 (O_67,N_4897,N_4835);
and UO_68 (O_68,N_4660,N_4729);
and UO_69 (O_69,N_4670,N_4665);
and UO_70 (O_70,N_4513,N_4655);
or UO_71 (O_71,N_4923,N_4688);
xor UO_72 (O_72,N_4767,N_4924);
and UO_73 (O_73,N_4755,N_4772);
nor UO_74 (O_74,N_4563,N_4526);
nand UO_75 (O_75,N_4558,N_4840);
or UO_76 (O_76,N_4856,N_4793);
nand UO_77 (O_77,N_4508,N_4754);
nor UO_78 (O_78,N_4985,N_4573);
nand UO_79 (O_79,N_4715,N_4521);
or UO_80 (O_80,N_4528,N_4669);
or UO_81 (O_81,N_4946,N_4631);
nand UO_82 (O_82,N_4568,N_4590);
and UO_83 (O_83,N_4931,N_4611);
nand UO_84 (O_84,N_4510,N_4692);
nor UO_85 (O_85,N_4935,N_4681);
nor UO_86 (O_86,N_4562,N_4879);
and UO_87 (O_87,N_4889,N_4776);
nor UO_88 (O_88,N_4567,N_4546);
nor UO_89 (O_89,N_4932,N_4704);
or UO_90 (O_90,N_4928,N_4737);
or UO_91 (O_91,N_4543,N_4829);
nor UO_92 (O_92,N_4620,N_4757);
and UO_93 (O_93,N_4731,N_4641);
nor UO_94 (O_94,N_4904,N_4834);
or UO_95 (O_95,N_4943,N_4844);
nand UO_96 (O_96,N_4745,N_4734);
nand UO_97 (O_97,N_4846,N_4648);
xor UO_98 (O_98,N_4527,N_4691);
nor UO_99 (O_99,N_4938,N_4653);
or UO_100 (O_100,N_4936,N_4668);
nand UO_101 (O_101,N_4953,N_4585);
xor UO_102 (O_102,N_4501,N_4947);
or UO_103 (O_103,N_4724,N_4867);
nand UO_104 (O_104,N_4604,N_4566);
or UO_105 (O_105,N_4581,N_4981);
and UO_106 (O_106,N_4825,N_4547);
nor UO_107 (O_107,N_4824,N_4820);
nor UO_108 (O_108,N_4530,N_4814);
nor UO_109 (O_109,N_4821,N_4725);
nand UO_110 (O_110,N_4605,N_4969);
nor UO_111 (O_111,N_4603,N_4906);
and UO_112 (O_112,N_4659,N_4714);
nor UO_113 (O_113,N_4656,N_4750);
nand UO_114 (O_114,N_4639,N_4743);
nor UO_115 (O_115,N_4771,N_4720);
or UO_116 (O_116,N_4752,N_4638);
and UO_117 (O_117,N_4869,N_4892);
or UO_118 (O_118,N_4919,N_4642);
and UO_119 (O_119,N_4676,N_4803);
nand UO_120 (O_120,N_4934,N_4650);
and UO_121 (O_121,N_4636,N_4859);
nand UO_122 (O_122,N_4597,N_4758);
nor UO_123 (O_123,N_4523,N_4628);
nor UO_124 (O_124,N_4921,N_4532);
xnor UO_125 (O_125,N_4589,N_4832);
nand UO_126 (O_126,N_4826,N_4916);
nand UO_127 (O_127,N_4839,N_4808);
and UO_128 (O_128,N_4645,N_4876);
nor UO_129 (O_129,N_4858,N_4942);
and UO_130 (O_130,N_4893,N_4635);
nor UO_131 (O_131,N_4961,N_4845);
nand UO_132 (O_132,N_4520,N_4525);
nand UO_133 (O_133,N_4555,N_4583);
nor UO_134 (O_134,N_4594,N_4788);
nor UO_135 (O_135,N_4579,N_4806);
or UO_136 (O_136,N_4877,N_4700);
nand UO_137 (O_137,N_4637,N_4914);
nor UO_138 (O_138,N_4918,N_4672);
and UO_139 (O_139,N_4619,N_4795);
nor UO_140 (O_140,N_4964,N_4503);
or UO_141 (O_141,N_4880,N_4662);
and UO_142 (O_142,N_4874,N_4842);
nor UO_143 (O_143,N_4862,N_4847);
nand UO_144 (O_144,N_4800,N_4907);
and UO_145 (O_145,N_4701,N_4679);
nand UO_146 (O_146,N_4977,N_4564);
nor UO_147 (O_147,N_4868,N_4779);
nand UO_148 (O_148,N_4671,N_4640);
nand UO_149 (O_149,N_4930,N_4732);
nand UO_150 (O_150,N_4954,N_4865);
nand UO_151 (O_151,N_4984,N_4735);
nor UO_152 (O_152,N_4813,N_4598);
and UO_153 (O_153,N_4905,N_4883);
nand UO_154 (O_154,N_4871,N_4811);
and UO_155 (O_155,N_4855,N_4926);
nor UO_156 (O_156,N_4587,N_4506);
nand UO_157 (O_157,N_4998,N_4851);
nor UO_158 (O_158,N_4553,N_4557);
nand UO_159 (O_159,N_4744,N_4816);
nor UO_160 (O_160,N_4539,N_4515);
nor UO_161 (O_161,N_4556,N_4802);
and UO_162 (O_162,N_4753,N_4927);
or UO_163 (O_163,N_4891,N_4728);
or UO_164 (O_164,N_4790,N_4770);
or UO_165 (O_165,N_4576,N_4929);
nor UO_166 (O_166,N_4831,N_4643);
nor UO_167 (O_167,N_4956,N_4578);
and UO_168 (O_168,N_4719,N_4854);
or UO_169 (O_169,N_4657,N_4596);
or UO_170 (O_170,N_4677,N_4777);
nand UO_171 (O_171,N_4709,N_4747);
xor UO_172 (O_172,N_4975,N_4833);
or UO_173 (O_173,N_4535,N_4970);
and UO_174 (O_174,N_4948,N_4507);
and UO_175 (O_175,N_4712,N_4992);
nand UO_176 (O_176,N_4807,N_4733);
or UO_177 (O_177,N_4861,N_4915);
and UO_178 (O_178,N_4617,N_4756);
or UO_179 (O_179,N_4974,N_4945);
nor UO_180 (O_180,N_4864,N_4610);
nand UO_181 (O_181,N_4972,N_4976);
and UO_182 (O_182,N_4796,N_4678);
nand UO_183 (O_183,N_4529,N_4870);
or UO_184 (O_184,N_4996,N_4785);
or UO_185 (O_185,N_4592,N_4748);
or UO_186 (O_186,N_4572,N_4804);
nand UO_187 (O_187,N_4791,N_4894);
nand UO_188 (O_188,N_4775,N_4608);
nand UO_189 (O_189,N_4702,N_4612);
and UO_190 (O_190,N_4537,N_4517);
xnor UO_191 (O_191,N_4886,N_4577);
and UO_192 (O_192,N_4634,N_4674);
and UO_193 (O_193,N_4601,N_4627);
nor UO_194 (O_194,N_4783,N_4722);
nand UO_195 (O_195,N_4917,N_4901);
and UO_196 (O_196,N_4978,N_4616);
nor UO_197 (O_197,N_4607,N_4717);
and UO_198 (O_198,N_4559,N_4623);
nand UO_199 (O_199,N_4959,N_4552);
nand UO_200 (O_200,N_4618,N_4726);
or UO_201 (O_201,N_4565,N_4647);
nor UO_202 (O_202,N_4673,N_4654);
and UO_203 (O_203,N_4695,N_4966);
nand UO_204 (O_204,N_4990,N_4644);
nor UO_205 (O_205,N_4911,N_4761);
nor UO_206 (O_206,N_4533,N_4898);
and UO_207 (O_207,N_4941,N_4711);
or UO_208 (O_208,N_4884,N_4857);
nand UO_209 (O_209,N_4863,N_4736);
nand UO_210 (O_210,N_4955,N_4727);
nor UO_211 (O_211,N_4989,N_4949);
or UO_212 (O_212,N_4738,N_4538);
nor UO_213 (O_213,N_4810,N_4584);
nor UO_214 (O_214,N_4666,N_4624);
nor UO_215 (O_215,N_4571,N_4836);
nand UO_216 (O_216,N_4652,N_4554);
and UO_217 (O_217,N_4841,N_4991);
nand UO_218 (O_218,N_4746,N_4690);
or UO_219 (O_219,N_4698,N_4613);
nand UO_220 (O_220,N_4534,N_4699);
xnor UO_221 (O_221,N_4995,N_4630);
nor UO_222 (O_222,N_4760,N_4518);
nand UO_223 (O_223,N_4664,N_4707);
nand UO_224 (O_224,N_4980,N_4830);
and UO_225 (O_225,N_4548,N_4878);
nand UO_226 (O_226,N_4675,N_4988);
or UO_227 (O_227,N_4838,N_4549);
nand UO_228 (O_228,N_4625,N_4885);
nand UO_229 (O_229,N_4809,N_4570);
nor UO_230 (O_230,N_4632,N_4950);
nor UO_231 (O_231,N_4773,N_4667);
nand UO_232 (O_232,N_4541,N_4762);
or UO_233 (O_233,N_4504,N_4960);
and UO_234 (O_234,N_4536,N_4872);
and UO_235 (O_235,N_4769,N_4912);
nand UO_236 (O_236,N_4786,N_4766);
xor UO_237 (O_237,N_4542,N_4680);
or UO_238 (O_238,N_4718,N_4502);
or UO_239 (O_239,N_4920,N_4633);
and UO_240 (O_240,N_4505,N_4658);
nand UO_241 (O_241,N_4703,N_4774);
and UO_242 (O_242,N_4999,N_4925);
and UO_243 (O_243,N_4944,N_4606);
nand UO_244 (O_244,N_4778,N_4599);
nand UO_245 (O_245,N_4696,N_4646);
and UO_246 (O_246,N_4514,N_4739);
nor UO_247 (O_247,N_4600,N_4968);
and UO_248 (O_248,N_4903,N_4818);
and UO_249 (O_249,N_4764,N_4910);
nand UO_250 (O_250,N_4946,N_4890);
nand UO_251 (O_251,N_4590,N_4577);
and UO_252 (O_252,N_4993,N_4564);
nor UO_253 (O_253,N_4585,N_4529);
or UO_254 (O_254,N_4973,N_4890);
and UO_255 (O_255,N_4943,N_4710);
and UO_256 (O_256,N_4682,N_4881);
or UO_257 (O_257,N_4834,N_4748);
and UO_258 (O_258,N_4828,N_4757);
xnor UO_259 (O_259,N_4558,N_4745);
or UO_260 (O_260,N_4620,N_4810);
nor UO_261 (O_261,N_4980,N_4856);
or UO_262 (O_262,N_4935,N_4561);
nor UO_263 (O_263,N_4545,N_4701);
nor UO_264 (O_264,N_4846,N_4752);
or UO_265 (O_265,N_4844,N_4680);
and UO_266 (O_266,N_4581,N_4836);
and UO_267 (O_267,N_4836,N_4659);
and UO_268 (O_268,N_4847,N_4792);
nand UO_269 (O_269,N_4774,N_4967);
nor UO_270 (O_270,N_4935,N_4680);
or UO_271 (O_271,N_4764,N_4902);
or UO_272 (O_272,N_4728,N_4505);
nor UO_273 (O_273,N_4527,N_4957);
nor UO_274 (O_274,N_4542,N_4892);
or UO_275 (O_275,N_4580,N_4926);
and UO_276 (O_276,N_4973,N_4978);
nand UO_277 (O_277,N_4790,N_4967);
xnor UO_278 (O_278,N_4548,N_4520);
or UO_279 (O_279,N_4861,N_4564);
or UO_280 (O_280,N_4540,N_4688);
nor UO_281 (O_281,N_4972,N_4831);
nand UO_282 (O_282,N_4754,N_4566);
or UO_283 (O_283,N_4719,N_4984);
and UO_284 (O_284,N_4516,N_4711);
and UO_285 (O_285,N_4560,N_4694);
nor UO_286 (O_286,N_4956,N_4779);
and UO_287 (O_287,N_4579,N_4893);
xnor UO_288 (O_288,N_4555,N_4566);
and UO_289 (O_289,N_4714,N_4670);
nand UO_290 (O_290,N_4773,N_4604);
nor UO_291 (O_291,N_4617,N_4508);
and UO_292 (O_292,N_4674,N_4667);
and UO_293 (O_293,N_4706,N_4588);
nor UO_294 (O_294,N_4981,N_4625);
and UO_295 (O_295,N_4735,N_4563);
nand UO_296 (O_296,N_4611,N_4672);
nor UO_297 (O_297,N_4675,N_4902);
nand UO_298 (O_298,N_4651,N_4561);
and UO_299 (O_299,N_4792,N_4781);
nor UO_300 (O_300,N_4771,N_4869);
or UO_301 (O_301,N_4537,N_4918);
nand UO_302 (O_302,N_4852,N_4600);
nand UO_303 (O_303,N_4627,N_4774);
nor UO_304 (O_304,N_4975,N_4910);
nor UO_305 (O_305,N_4568,N_4582);
nor UO_306 (O_306,N_4790,N_4883);
nand UO_307 (O_307,N_4752,N_4935);
or UO_308 (O_308,N_4674,N_4874);
nand UO_309 (O_309,N_4941,N_4990);
or UO_310 (O_310,N_4727,N_4548);
or UO_311 (O_311,N_4500,N_4749);
and UO_312 (O_312,N_4827,N_4870);
and UO_313 (O_313,N_4949,N_4751);
nor UO_314 (O_314,N_4873,N_4892);
nor UO_315 (O_315,N_4573,N_4586);
and UO_316 (O_316,N_4859,N_4771);
nand UO_317 (O_317,N_4896,N_4659);
or UO_318 (O_318,N_4864,N_4624);
or UO_319 (O_319,N_4843,N_4882);
or UO_320 (O_320,N_4958,N_4510);
nor UO_321 (O_321,N_4982,N_4625);
and UO_322 (O_322,N_4925,N_4741);
and UO_323 (O_323,N_4940,N_4880);
nand UO_324 (O_324,N_4913,N_4539);
or UO_325 (O_325,N_4617,N_4941);
and UO_326 (O_326,N_4534,N_4897);
and UO_327 (O_327,N_4707,N_4962);
nand UO_328 (O_328,N_4627,N_4959);
or UO_329 (O_329,N_4740,N_4660);
nor UO_330 (O_330,N_4634,N_4624);
nor UO_331 (O_331,N_4673,N_4801);
nand UO_332 (O_332,N_4747,N_4625);
nor UO_333 (O_333,N_4919,N_4587);
and UO_334 (O_334,N_4766,N_4899);
nor UO_335 (O_335,N_4925,N_4699);
or UO_336 (O_336,N_4877,N_4733);
nor UO_337 (O_337,N_4547,N_4855);
or UO_338 (O_338,N_4673,N_4670);
nand UO_339 (O_339,N_4710,N_4727);
nor UO_340 (O_340,N_4776,N_4600);
or UO_341 (O_341,N_4917,N_4785);
nand UO_342 (O_342,N_4951,N_4532);
nand UO_343 (O_343,N_4772,N_4941);
or UO_344 (O_344,N_4606,N_4996);
nand UO_345 (O_345,N_4624,N_4738);
nand UO_346 (O_346,N_4522,N_4552);
and UO_347 (O_347,N_4541,N_4604);
and UO_348 (O_348,N_4849,N_4708);
nand UO_349 (O_349,N_4522,N_4735);
nand UO_350 (O_350,N_4794,N_4700);
nand UO_351 (O_351,N_4966,N_4696);
nor UO_352 (O_352,N_4872,N_4772);
nand UO_353 (O_353,N_4734,N_4655);
nor UO_354 (O_354,N_4749,N_4676);
and UO_355 (O_355,N_4741,N_4772);
nand UO_356 (O_356,N_4792,N_4643);
or UO_357 (O_357,N_4583,N_4948);
and UO_358 (O_358,N_4685,N_4873);
nand UO_359 (O_359,N_4571,N_4826);
and UO_360 (O_360,N_4580,N_4996);
or UO_361 (O_361,N_4504,N_4992);
nand UO_362 (O_362,N_4604,N_4950);
or UO_363 (O_363,N_4675,N_4926);
nor UO_364 (O_364,N_4549,N_4583);
and UO_365 (O_365,N_4598,N_4841);
or UO_366 (O_366,N_4859,N_4581);
nor UO_367 (O_367,N_4607,N_4734);
nor UO_368 (O_368,N_4851,N_4546);
nand UO_369 (O_369,N_4753,N_4847);
or UO_370 (O_370,N_4604,N_4998);
and UO_371 (O_371,N_4795,N_4598);
nand UO_372 (O_372,N_4561,N_4809);
or UO_373 (O_373,N_4574,N_4964);
or UO_374 (O_374,N_4617,N_4521);
nor UO_375 (O_375,N_4996,N_4906);
nor UO_376 (O_376,N_4793,N_4778);
nor UO_377 (O_377,N_4880,N_4952);
and UO_378 (O_378,N_4604,N_4772);
or UO_379 (O_379,N_4645,N_4572);
nor UO_380 (O_380,N_4718,N_4972);
nor UO_381 (O_381,N_4563,N_4610);
nand UO_382 (O_382,N_4682,N_4970);
nand UO_383 (O_383,N_4560,N_4922);
nand UO_384 (O_384,N_4822,N_4741);
and UO_385 (O_385,N_4759,N_4675);
nand UO_386 (O_386,N_4676,N_4841);
or UO_387 (O_387,N_4614,N_4649);
nor UO_388 (O_388,N_4759,N_4916);
and UO_389 (O_389,N_4640,N_4594);
nor UO_390 (O_390,N_4886,N_4858);
and UO_391 (O_391,N_4580,N_4741);
nor UO_392 (O_392,N_4519,N_4528);
and UO_393 (O_393,N_4979,N_4950);
nand UO_394 (O_394,N_4607,N_4919);
or UO_395 (O_395,N_4922,N_4533);
and UO_396 (O_396,N_4903,N_4786);
or UO_397 (O_397,N_4887,N_4876);
nand UO_398 (O_398,N_4885,N_4955);
nand UO_399 (O_399,N_4558,N_4794);
and UO_400 (O_400,N_4976,N_4716);
or UO_401 (O_401,N_4865,N_4837);
nor UO_402 (O_402,N_4929,N_4817);
and UO_403 (O_403,N_4760,N_4844);
nor UO_404 (O_404,N_4716,N_4506);
and UO_405 (O_405,N_4953,N_4507);
and UO_406 (O_406,N_4518,N_4693);
nor UO_407 (O_407,N_4789,N_4782);
or UO_408 (O_408,N_4874,N_4828);
xnor UO_409 (O_409,N_4923,N_4638);
and UO_410 (O_410,N_4555,N_4973);
nor UO_411 (O_411,N_4598,N_4668);
nand UO_412 (O_412,N_4710,N_4718);
nor UO_413 (O_413,N_4744,N_4740);
nand UO_414 (O_414,N_4603,N_4549);
or UO_415 (O_415,N_4958,N_4599);
and UO_416 (O_416,N_4981,N_4847);
or UO_417 (O_417,N_4603,N_4970);
nand UO_418 (O_418,N_4550,N_4876);
nor UO_419 (O_419,N_4517,N_4701);
or UO_420 (O_420,N_4819,N_4842);
nand UO_421 (O_421,N_4784,N_4695);
and UO_422 (O_422,N_4837,N_4702);
nor UO_423 (O_423,N_4713,N_4663);
nor UO_424 (O_424,N_4782,N_4505);
nand UO_425 (O_425,N_4803,N_4547);
nor UO_426 (O_426,N_4791,N_4705);
xor UO_427 (O_427,N_4623,N_4691);
nand UO_428 (O_428,N_4577,N_4724);
or UO_429 (O_429,N_4941,N_4704);
or UO_430 (O_430,N_4720,N_4606);
nand UO_431 (O_431,N_4781,N_4712);
nor UO_432 (O_432,N_4554,N_4740);
or UO_433 (O_433,N_4630,N_4907);
or UO_434 (O_434,N_4574,N_4989);
nand UO_435 (O_435,N_4807,N_4563);
xnor UO_436 (O_436,N_4775,N_4809);
or UO_437 (O_437,N_4680,N_4573);
nor UO_438 (O_438,N_4802,N_4710);
nand UO_439 (O_439,N_4537,N_4688);
nand UO_440 (O_440,N_4813,N_4696);
nor UO_441 (O_441,N_4729,N_4511);
nor UO_442 (O_442,N_4937,N_4963);
nand UO_443 (O_443,N_4542,N_4558);
and UO_444 (O_444,N_4845,N_4518);
or UO_445 (O_445,N_4574,N_4757);
and UO_446 (O_446,N_4915,N_4519);
or UO_447 (O_447,N_4509,N_4886);
or UO_448 (O_448,N_4895,N_4947);
or UO_449 (O_449,N_4500,N_4695);
or UO_450 (O_450,N_4607,N_4956);
nor UO_451 (O_451,N_4967,N_4806);
nand UO_452 (O_452,N_4871,N_4929);
or UO_453 (O_453,N_4670,N_4861);
nand UO_454 (O_454,N_4799,N_4696);
nor UO_455 (O_455,N_4549,N_4716);
nor UO_456 (O_456,N_4842,N_4886);
nor UO_457 (O_457,N_4828,N_4510);
nand UO_458 (O_458,N_4756,N_4736);
nand UO_459 (O_459,N_4869,N_4894);
or UO_460 (O_460,N_4723,N_4718);
and UO_461 (O_461,N_4666,N_4694);
nand UO_462 (O_462,N_4935,N_4933);
nand UO_463 (O_463,N_4852,N_4867);
nand UO_464 (O_464,N_4788,N_4938);
or UO_465 (O_465,N_4670,N_4951);
nand UO_466 (O_466,N_4735,N_4921);
or UO_467 (O_467,N_4664,N_4840);
nand UO_468 (O_468,N_4754,N_4619);
nor UO_469 (O_469,N_4703,N_4598);
or UO_470 (O_470,N_4517,N_4987);
nand UO_471 (O_471,N_4866,N_4521);
or UO_472 (O_472,N_4652,N_4829);
and UO_473 (O_473,N_4814,N_4968);
and UO_474 (O_474,N_4976,N_4916);
or UO_475 (O_475,N_4784,N_4787);
or UO_476 (O_476,N_4868,N_4689);
nand UO_477 (O_477,N_4609,N_4562);
nand UO_478 (O_478,N_4698,N_4762);
nor UO_479 (O_479,N_4609,N_4925);
and UO_480 (O_480,N_4867,N_4502);
and UO_481 (O_481,N_4858,N_4965);
and UO_482 (O_482,N_4546,N_4758);
and UO_483 (O_483,N_4566,N_4936);
xor UO_484 (O_484,N_4666,N_4589);
and UO_485 (O_485,N_4787,N_4562);
and UO_486 (O_486,N_4723,N_4923);
and UO_487 (O_487,N_4761,N_4606);
or UO_488 (O_488,N_4695,N_4838);
or UO_489 (O_489,N_4935,N_4633);
nand UO_490 (O_490,N_4552,N_4628);
nand UO_491 (O_491,N_4692,N_4992);
and UO_492 (O_492,N_4904,N_4798);
nor UO_493 (O_493,N_4557,N_4667);
or UO_494 (O_494,N_4659,N_4844);
xnor UO_495 (O_495,N_4936,N_4725);
nand UO_496 (O_496,N_4697,N_4723);
or UO_497 (O_497,N_4823,N_4628);
and UO_498 (O_498,N_4542,N_4869);
or UO_499 (O_499,N_4884,N_4553);
nor UO_500 (O_500,N_4525,N_4870);
and UO_501 (O_501,N_4888,N_4647);
or UO_502 (O_502,N_4705,N_4812);
or UO_503 (O_503,N_4626,N_4593);
nor UO_504 (O_504,N_4720,N_4562);
and UO_505 (O_505,N_4792,N_4686);
nand UO_506 (O_506,N_4977,N_4639);
and UO_507 (O_507,N_4762,N_4688);
nor UO_508 (O_508,N_4577,N_4579);
and UO_509 (O_509,N_4900,N_4777);
or UO_510 (O_510,N_4834,N_4560);
nor UO_511 (O_511,N_4888,N_4829);
or UO_512 (O_512,N_4985,N_4925);
or UO_513 (O_513,N_4557,N_4538);
and UO_514 (O_514,N_4630,N_4761);
or UO_515 (O_515,N_4616,N_4618);
and UO_516 (O_516,N_4831,N_4574);
or UO_517 (O_517,N_4537,N_4658);
or UO_518 (O_518,N_4756,N_4722);
and UO_519 (O_519,N_4861,N_4651);
and UO_520 (O_520,N_4934,N_4541);
nand UO_521 (O_521,N_4723,N_4845);
or UO_522 (O_522,N_4613,N_4655);
or UO_523 (O_523,N_4593,N_4532);
nand UO_524 (O_524,N_4545,N_4840);
and UO_525 (O_525,N_4946,N_4923);
and UO_526 (O_526,N_4717,N_4596);
nand UO_527 (O_527,N_4547,N_4656);
xor UO_528 (O_528,N_4723,N_4748);
or UO_529 (O_529,N_4828,N_4537);
nor UO_530 (O_530,N_4890,N_4940);
and UO_531 (O_531,N_4823,N_4877);
or UO_532 (O_532,N_4972,N_4720);
nor UO_533 (O_533,N_4791,N_4606);
or UO_534 (O_534,N_4724,N_4738);
nor UO_535 (O_535,N_4658,N_4962);
nor UO_536 (O_536,N_4834,N_4865);
and UO_537 (O_537,N_4541,N_4565);
nand UO_538 (O_538,N_4600,N_4640);
nand UO_539 (O_539,N_4854,N_4858);
nor UO_540 (O_540,N_4709,N_4882);
or UO_541 (O_541,N_4838,N_4979);
and UO_542 (O_542,N_4782,N_4859);
nor UO_543 (O_543,N_4725,N_4509);
or UO_544 (O_544,N_4867,N_4680);
nand UO_545 (O_545,N_4838,N_4689);
and UO_546 (O_546,N_4589,N_4771);
and UO_547 (O_547,N_4904,N_4885);
or UO_548 (O_548,N_4857,N_4615);
or UO_549 (O_549,N_4651,N_4611);
and UO_550 (O_550,N_4531,N_4865);
nand UO_551 (O_551,N_4514,N_4906);
and UO_552 (O_552,N_4561,N_4560);
and UO_553 (O_553,N_4755,N_4976);
nand UO_554 (O_554,N_4622,N_4993);
and UO_555 (O_555,N_4900,N_4600);
nor UO_556 (O_556,N_4985,N_4928);
and UO_557 (O_557,N_4532,N_4726);
nor UO_558 (O_558,N_4510,N_4753);
and UO_559 (O_559,N_4652,N_4787);
nor UO_560 (O_560,N_4990,N_4709);
xnor UO_561 (O_561,N_4572,N_4888);
nand UO_562 (O_562,N_4697,N_4794);
nand UO_563 (O_563,N_4926,N_4979);
and UO_564 (O_564,N_4637,N_4688);
nand UO_565 (O_565,N_4542,N_4668);
or UO_566 (O_566,N_4849,N_4914);
and UO_567 (O_567,N_4766,N_4811);
or UO_568 (O_568,N_4583,N_4771);
nand UO_569 (O_569,N_4652,N_4977);
nor UO_570 (O_570,N_4827,N_4911);
or UO_571 (O_571,N_4985,N_4829);
or UO_572 (O_572,N_4785,N_4808);
nor UO_573 (O_573,N_4605,N_4757);
nand UO_574 (O_574,N_4547,N_4596);
and UO_575 (O_575,N_4861,N_4558);
nand UO_576 (O_576,N_4690,N_4626);
nor UO_577 (O_577,N_4578,N_4686);
and UO_578 (O_578,N_4756,N_4972);
or UO_579 (O_579,N_4975,N_4524);
and UO_580 (O_580,N_4639,N_4566);
and UO_581 (O_581,N_4914,N_4783);
or UO_582 (O_582,N_4953,N_4921);
nor UO_583 (O_583,N_4573,N_4670);
nand UO_584 (O_584,N_4782,N_4847);
nand UO_585 (O_585,N_4641,N_4684);
or UO_586 (O_586,N_4696,N_4840);
nor UO_587 (O_587,N_4934,N_4968);
and UO_588 (O_588,N_4855,N_4753);
nand UO_589 (O_589,N_4848,N_4753);
nand UO_590 (O_590,N_4629,N_4891);
or UO_591 (O_591,N_4579,N_4715);
nand UO_592 (O_592,N_4872,N_4859);
nand UO_593 (O_593,N_4959,N_4684);
nor UO_594 (O_594,N_4717,N_4604);
nand UO_595 (O_595,N_4541,N_4669);
nor UO_596 (O_596,N_4521,N_4668);
or UO_597 (O_597,N_4550,N_4599);
nand UO_598 (O_598,N_4791,N_4697);
nand UO_599 (O_599,N_4789,N_4868);
and UO_600 (O_600,N_4519,N_4880);
or UO_601 (O_601,N_4565,N_4582);
and UO_602 (O_602,N_4748,N_4778);
and UO_603 (O_603,N_4911,N_4633);
nand UO_604 (O_604,N_4511,N_4778);
nor UO_605 (O_605,N_4959,N_4925);
nor UO_606 (O_606,N_4729,N_4744);
nor UO_607 (O_607,N_4917,N_4963);
nor UO_608 (O_608,N_4862,N_4733);
nand UO_609 (O_609,N_4948,N_4962);
or UO_610 (O_610,N_4858,N_4865);
nand UO_611 (O_611,N_4506,N_4947);
or UO_612 (O_612,N_4828,N_4992);
and UO_613 (O_613,N_4523,N_4736);
nor UO_614 (O_614,N_4777,N_4686);
nand UO_615 (O_615,N_4987,N_4510);
and UO_616 (O_616,N_4605,N_4963);
nor UO_617 (O_617,N_4856,N_4622);
and UO_618 (O_618,N_4774,N_4655);
nand UO_619 (O_619,N_4568,N_4882);
or UO_620 (O_620,N_4708,N_4515);
and UO_621 (O_621,N_4991,N_4572);
and UO_622 (O_622,N_4574,N_4579);
or UO_623 (O_623,N_4548,N_4717);
nor UO_624 (O_624,N_4711,N_4782);
xor UO_625 (O_625,N_4653,N_4872);
nor UO_626 (O_626,N_4958,N_4826);
nand UO_627 (O_627,N_4809,N_4565);
nor UO_628 (O_628,N_4685,N_4688);
or UO_629 (O_629,N_4723,N_4506);
nor UO_630 (O_630,N_4610,N_4769);
nor UO_631 (O_631,N_4549,N_4826);
nor UO_632 (O_632,N_4905,N_4744);
nor UO_633 (O_633,N_4677,N_4866);
or UO_634 (O_634,N_4510,N_4884);
nand UO_635 (O_635,N_4706,N_4826);
nor UO_636 (O_636,N_4788,N_4889);
or UO_637 (O_637,N_4556,N_4794);
nor UO_638 (O_638,N_4930,N_4845);
and UO_639 (O_639,N_4878,N_4792);
and UO_640 (O_640,N_4646,N_4504);
or UO_641 (O_641,N_4612,N_4853);
nor UO_642 (O_642,N_4826,N_4961);
nand UO_643 (O_643,N_4508,N_4986);
nor UO_644 (O_644,N_4830,N_4535);
or UO_645 (O_645,N_4999,N_4932);
or UO_646 (O_646,N_4791,N_4661);
nand UO_647 (O_647,N_4866,N_4969);
nand UO_648 (O_648,N_4824,N_4819);
and UO_649 (O_649,N_4511,N_4996);
xnor UO_650 (O_650,N_4625,N_4657);
nor UO_651 (O_651,N_4887,N_4786);
and UO_652 (O_652,N_4503,N_4720);
nor UO_653 (O_653,N_4859,N_4816);
xor UO_654 (O_654,N_4900,N_4606);
nand UO_655 (O_655,N_4892,N_4956);
or UO_656 (O_656,N_4906,N_4691);
xor UO_657 (O_657,N_4929,N_4870);
nor UO_658 (O_658,N_4914,N_4678);
and UO_659 (O_659,N_4973,N_4970);
or UO_660 (O_660,N_4995,N_4640);
and UO_661 (O_661,N_4767,N_4890);
or UO_662 (O_662,N_4627,N_4645);
or UO_663 (O_663,N_4781,N_4794);
nand UO_664 (O_664,N_4528,N_4719);
and UO_665 (O_665,N_4912,N_4946);
and UO_666 (O_666,N_4662,N_4668);
or UO_667 (O_667,N_4922,N_4765);
or UO_668 (O_668,N_4572,N_4984);
nand UO_669 (O_669,N_4684,N_4688);
nand UO_670 (O_670,N_4873,N_4538);
nor UO_671 (O_671,N_4706,N_4688);
and UO_672 (O_672,N_4784,N_4581);
nand UO_673 (O_673,N_4791,N_4882);
and UO_674 (O_674,N_4501,N_4520);
nand UO_675 (O_675,N_4597,N_4667);
and UO_676 (O_676,N_4825,N_4779);
and UO_677 (O_677,N_4895,N_4639);
nor UO_678 (O_678,N_4556,N_4725);
xnor UO_679 (O_679,N_4811,N_4733);
or UO_680 (O_680,N_4626,N_4958);
or UO_681 (O_681,N_4584,N_4648);
nor UO_682 (O_682,N_4744,N_4520);
or UO_683 (O_683,N_4546,N_4693);
nor UO_684 (O_684,N_4891,N_4765);
nor UO_685 (O_685,N_4724,N_4507);
or UO_686 (O_686,N_4886,N_4695);
nand UO_687 (O_687,N_4547,N_4571);
and UO_688 (O_688,N_4744,N_4800);
nor UO_689 (O_689,N_4992,N_4975);
xor UO_690 (O_690,N_4758,N_4690);
or UO_691 (O_691,N_4812,N_4909);
and UO_692 (O_692,N_4834,N_4601);
and UO_693 (O_693,N_4794,N_4831);
nand UO_694 (O_694,N_4687,N_4604);
and UO_695 (O_695,N_4567,N_4982);
nor UO_696 (O_696,N_4790,N_4651);
or UO_697 (O_697,N_4677,N_4846);
and UO_698 (O_698,N_4733,N_4998);
or UO_699 (O_699,N_4500,N_4901);
or UO_700 (O_700,N_4843,N_4883);
and UO_701 (O_701,N_4876,N_4800);
and UO_702 (O_702,N_4865,N_4512);
and UO_703 (O_703,N_4798,N_4751);
or UO_704 (O_704,N_4653,N_4760);
nor UO_705 (O_705,N_4504,N_4903);
or UO_706 (O_706,N_4563,N_4947);
nor UO_707 (O_707,N_4646,N_4902);
nand UO_708 (O_708,N_4710,N_4515);
or UO_709 (O_709,N_4962,N_4673);
nand UO_710 (O_710,N_4678,N_4953);
nor UO_711 (O_711,N_4531,N_4821);
nand UO_712 (O_712,N_4953,N_4754);
and UO_713 (O_713,N_4919,N_4957);
or UO_714 (O_714,N_4913,N_4753);
and UO_715 (O_715,N_4795,N_4864);
nor UO_716 (O_716,N_4511,N_4695);
or UO_717 (O_717,N_4743,N_4688);
nand UO_718 (O_718,N_4546,N_4706);
or UO_719 (O_719,N_4963,N_4753);
nor UO_720 (O_720,N_4935,N_4526);
and UO_721 (O_721,N_4597,N_4911);
xnor UO_722 (O_722,N_4712,N_4919);
nand UO_723 (O_723,N_4819,N_4726);
xnor UO_724 (O_724,N_4945,N_4827);
and UO_725 (O_725,N_4907,N_4986);
or UO_726 (O_726,N_4959,N_4553);
nor UO_727 (O_727,N_4990,N_4596);
or UO_728 (O_728,N_4966,N_4987);
or UO_729 (O_729,N_4856,N_4683);
and UO_730 (O_730,N_4926,N_4716);
nand UO_731 (O_731,N_4744,N_4637);
nand UO_732 (O_732,N_4988,N_4807);
and UO_733 (O_733,N_4566,N_4869);
nor UO_734 (O_734,N_4731,N_4883);
or UO_735 (O_735,N_4687,N_4615);
nor UO_736 (O_736,N_4712,N_4658);
nor UO_737 (O_737,N_4889,N_4710);
nor UO_738 (O_738,N_4715,N_4898);
nand UO_739 (O_739,N_4751,N_4830);
or UO_740 (O_740,N_4542,N_4860);
nand UO_741 (O_741,N_4673,N_4835);
or UO_742 (O_742,N_4531,N_4975);
nor UO_743 (O_743,N_4626,N_4604);
or UO_744 (O_744,N_4805,N_4618);
or UO_745 (O_745,N_4836,N_4750);
xnor UO_746 (O_746,N_4778,N_4732);
or UO_747 (O_747,N_4907,N_4905);
and UO_748 (O_748,N_4519,N_4772);
nand UO_749 (O_749,N_4564,N_4650);
or UO_750 (O_750,N_4981,N_4537);
or UO_751 (O_751,N_4653,N_4934);
nand UO_752 (O_752,N_4924,N_4528);
xnor UO_753 (O_753,N_4789,N_4607);
and UO_754 (O_754,N_4517,N_4654);
or UO_755 (O_755,N_4632,N_4735);
or UO_756 (O_756,N_4619,N_4564);
nand UO_757 (O_757,N_4925,N_4587);
and UO_758 (O_758,N_4838,N_4641);
and UO_759 (O_759,N_4565,N_4500);
nand UO_760 (O_760,N_4600,N_4975);
nand UO_761 (O_761,N_4908,N_4711);
nand UO_762 (O_762,N_4802,N_4581);
nand UO_763 (O_763,N_4772,N_4994);
nand UO_764 (O_764,N_4731,N_4577);
nand UO_765 (O_765,N_4510,N_4931);
xnor UO_766 (O_766,N_4739,N_4669);
and UO_767 (O_767,N_4924,N_4806);
or UO_768 (O_768,N_4549,N_4789);
and UO_769 (O_769,N_4988,N_4937);
or UO_770 (O_770,N_4821,N_4670);
nor UO_771 (O_771,N_4713,N_4707);
or UO_772 (O_772,N_4995,N_4796);
and UO_773 (O_773,N_4653,N_4975);
nand UO_774 (O_774,N_4549,N_4651);
nor UO_775 (O_775,N_4932,N_4697);
nor UO_776 (O_776,N_4803,N_4519);
and UO_777 (O_777,N_4687,N_4523);
and UO_778 (O_778,N_4985,N_4831);
or UO_779 (O_779,N_4751,N_4596);
nand UO_780 (O_780,N_4661,N_4688);
or UO_781 (O_781,N_4573,N_4904);
or UO_782 (O_782,N_4654,N_4677);
or UO_783 (O_783,N_4985,N_4994);
and UO_784 (O_784,N_4736,N_4821);
nor UO_785 (O_785,N_4829,N_4986);
or UO_786 (O_786,N_4764,N_4632);
and UO_787 (O_787,N_4520,N_4685);
or UO_788 (O_788,N_4950,N_4573);
nand UO_789 (O_789,N_4849,N_4613);
nor UO_790 (O_790,N_4578,N_4563);
nand UO_791 (O_791,N_4642,N_4713);
and UO_792 (O_792,N_4892,N_4760);
nor UO_793 (O_793,N_4662,N_4787);
and UO_794 (O_794,N_4947,N_4601);
and UO_795 (O_795,N_4567,N_4917);
nor UO_796 (O_796,N_4919,N_4992);
and UO_797 (O_797,N_4839,N_4669);
nor UO_798 (O_798,N_4626,N_4715);
nor UO_799 (O_799,N_4824,N_4891);
nand UO_800 (O_800,N_4831,N_4777);
and UO_801 (O_801,N_4613,N_4910);
nand UO_802 (O_802,N_4521,N_4503);
nor UO_803 (O_803,N_4696,N_4906);
or UO_804 (O_804,N_4775,N_4814);
nor UO_805 (O_805,N_4838,N_4806);
nand UO_806 (O_806,N_4755,N_4873);
nor UO_807 (O_807,N_4903,N_4797);
and UO_808 (O_808,N_4924,N_4955);
nor UO_809 (O_809,N_4934,N_4665);
or UO_810 (O_810,N_4776,N_4883);
or UO_811 (O_811,N_4578,N_4570);
or UO_812 (O_812,N_4762,N_4500);
or UO_813 (O_813,N_4988,N_4571);
or UO_814 (O_814,N_4972,N_4770);
nand UO_815 (O_815,N_4948,N_4533);
nor UO_816 (O_816,N_4554,N_4600);
nand UO_817 (O_817,N_4525,N_4726);
and UO_818 (O_818,N_4878,N_4701);
and UO_819 (O_819,N_4760,N_4539);
and UO_820 (O_820,N_4931,N_4552);
nand UO_821 (O_821,N_4723,N_4523);
nand UO_822 (O_822,N_4924,N_4660);
and UO_823 (O_823,N_4853,N_4593);
nand UO_824 (O_824,N_4834,N_4910);
or UO_825 (O_825,N_4700,N_4995);
nand UO_826 (O_826,N_4720,N_4605);
xnor UO_827 (O_827,N_4678,N_4512);
or UO_828 (O_828,N_4759,N_4989);
nand UO_829 (O_829,N_4626,N_4713);
or UO_830 (O_830,N_4767,N_4542);
nor UO_831 (O_831,N_4887,N_4800);
nand UO_832 (O_832,N_4643,N_4758);
and UO_833 (O_833,N_4908,N_4890);
nor UO_834 (O_834,N_4845,N_4954);
nor UO_835 (O_835,N_4775,N_4877);
nand UO_836 (O_836,N_4507,N_4519);
nand UO_837 (O_837,N_4813,N_4990);
nand UO_838 (O_838,N_4875,N_4880);
and UO_839 (O_839,N_4649,N_4987);
nor UO_840 (O_840,N_4970,N_4654);
nor UO_841 (O_841,N_4869,N_4956);
nand UO_842 (O_842,N_4535,N_4945);
nor UO_843 (O_843,N_4675,N_4952);
nand UO_844 (O_844,N_4767,N_4668);
and UO_845 (O_845,N_4562,N_4958);
and UO_846 (O_846,N_4819,N_4665);
or UO_847 (O_847,N_4513,N_4697);
nand UO_848 (O_848,N_4515,N_4651);
nand UO_849 (O_849,N_4526,N_4648);
and UO_850 (O_850,N_4628,N_4942);
or UO_851 (O_851,N_4699,N_4815);
nor UO_852 (O_852,N_4789,N_4927);
and UO_853 (O_853,N_4982,N_4622);
or UO_854 (O_854,N_4678,N_4849);
nor UO_855 (O_855,N_4810,N_4782);
or UO_856 (O_856,N_4943,N_4633);
nand UO_857 (O_857,N_4600,N_4676);
nand UO_858 (O_858,N_4636,N_4674);
nor UO_859 (O_859,N_4801,N_4808);
nor UO_860 (O_860,N_4870,N_4749);
nand UO_861 (O_861,N_4558,N_4777);
and UO_862 (O_862,N_4687,N_4911);
nor UO_863 (O_863,N_4863,N_4874);
nand UO_864 (O_864,N_4874,N_4593);
or UO_865 (O_865,N_4704,N_4540);
nor UO_866 (O_866,N_4958,N_4653);
xnor UO_867 (O_867,N_4897,N_4668);
and UO_868 (O_868,N_4901,N_4918);
and UO_869 (O_869,N_4681,N_4871);
nor UO_870 (O_870,N_4675,N_4812);
nand UO_871 (O_871,N_4879,N_4639);
and UO_872 (O_872,N_4998,N_4841);
nor UO_873 (O_873,N_4848,N_4939);
or UO_874 (O_874,N_4957,N_4988);
xnor UO_875 (O_875,N_4581,N_4694);
or UO_876 (O_876,N_4946,N_4507);
or UO_877 (O_877,N_4542,N_4938);
nand UO_878 (O_878,N_4571,N_4533);
nand UO_879 (O_879,N_4575,N_4646);
or UO_880 (O_880,N_4672,N_4588);
nand UO_881 (O_881,N_4858,N_4971);
and UO_882 (O_882,N_4555,N_4877);
xnor UO_883 (O_883,N_4554,N_4641);
nor UO_884 (O_884,N_4923,N_4772);
nand UO_885 (O_885,N_4830,N_4701);
and UO_886 (O_886,N_4716,N_4749);
or UO_887 (O_887,N_4663,N_4996);
nand UO_888 (O_888,N_4621,N_4577);
and UO_889 (O_889,N_4533,N_4573);
nor UO_890 (O_890,N_4581,N_4689);
and UO_891 (O_891,N_4935,N_4528);
or UO_892 (O_892,N_4942,N_4999);
nand UO_893 (O_893,N_4647,N_4963);
xor UO_894 (O_894,N_4780,N_4566);
xor UO_895 (O_895,N_4755,N_4955);
nand UO_896 (O_896,N_4672,N_4906);
nand UO_897 (O_897,N_4693,N_4759);
or UO_898 (O_898,N_4641,N_4559);
nor UO_899 (O_899,N_4580,N_4750);
or UO_900 (O_900,N_4815,N_4941);
nand UO_901 (O_901,N_4593,N_4558);
or UO_902 (O_902,N_4791,N_4716);
nor UO_903 (O_903,N_4931,N_4667);
nand UO_904 (O_904,N_4711,N_4618);
xnor UO_905 (O_905,N_4921,N_4567);
or UO_906 (O_906,N_4833,N_4552);
and UO_907 (O_907,N_4564,N_4582);
nand UO_908 (O_908,N_4974,N_4843);
or UO_909 (O_909,N_4773,N_4797);
and UO_910 (O_910,N_4857,N_4837);
or UO_911 (O_911,N_4762,N_4863);
nor UO_912 (O_912,N_4879,N_4921);
or UO_913 (O_913,N_4520,N_4555);
nand UO_914 (O_914,N_4719,N_4619);
and UO_915 (O_915,N_4725,N_4580);
and UO_916 (O_916,N_4607,N_4592);
or UO_917 (O_917,N_4862,N_4566);
nor UO_918 (O_918,N_4976,N_4820);
and UO_919 (O_919,N_4720,N_4561);
and UO_920 (O_920,N_4781,N_4847);
and UO_921 (O_921,N_4554,N_4500);
nor UO_922 (O_922,N_4559,N_4714);
xor UO_923 (O_923,N_4876,N_4595);
or UO_924 (O_924,N_4949,N_4642);
nor UO_925 (O_925,N_4534,N_4575);
and UO_926 (O_926,N_4757,N_4551);
or UO_927 (O_927,N_4970,N_4756);
nor UO_928 (O_928,N_4514,N_4625);
or UO_929 (O_929,N_4534,N_4500);
nor UO_930 (O_930,N_4906,N_4774);
nor UO_931 (O_931,N_4759,N_4601);
or UO_932 (O_932,N_4847,N_4581);
and UO_933 (O_933,N_4766,N_4874);
nor UO_934 (O_934,N_4727,N_4783);
and UO_935 (O_935,N_4537,N_4948);
nor UO_936 (O_936,N_4691,N_4685);
nand UO_937 (O_937,N_4660,N_4668);
or UO_938 (O_938,N_4789,N_4745);
and UO_939 (O_939,N_4680,N_4546);
nand UO_940 (O_940,N_4887,N_4789);
xor UO_941 (O_941,N_4956,N_4858);
and UO_942 (O_942,N_4726,N_4820);
nand UO_943 (O_943,N_4564,N_4567);
or UO_944 (O_944,N_4807,N_4942);
and UO_945 (O_945,N_4845,N_4645);
nor UO_946 (O_946,N_4862,N_4634);
or UO_947 (O_947,N_4704,N_4559);
nor UO_948 (O_948,N_4941,N_4829);
or UO_949 (O_949,N_4573,N_4833);
nor UO_950 (O_950,N_4737,N_4542);
nand UO_951 (O_951,N_4984,N_4788);
nand UO_952 (O_952,N_4591,N_4767);
nand UO_953 (O_953,N_4793,N_4846);
nor UO_954 (O_954,N_4920,N_4611);
or UO_955 (O_955,N_4900,N_4764);
nand UO_956 (O_956,N_4604,N_4721);
nand UO_957 (O_957,N_4503,N_4678);
or UO_958 (O_958,N_4947,N_4731);
nand UO_959 (O_959,N_4743,N_4593);
and UO_960 (O_960,N_4666,N_4918);
nand UO_961 (O_961,N_4981,N_4922);
or UO_962 (O_962,N_4733,N_4963);
xor UO_963 (O_963,N_4630,N_4504);
nand UO_964 (O_964,N_4990,N_4628);
nor UO_965 (O_965,N_4708,N_4793);
and UO_966 (O_966,N_4823,N_4558);
and UO_967 (O_967,N_4737,N_4697);
nor UO_968 (O_968,N_4712,N_4523);
nor UO_969 (O_969,N_4644,N_4695);
or UO_970 (O_970,N_4869,N_4526);
nor UO_971 (O_971,N_4987,N_4643);
nand UO_972 (O_972,N_4504,N_4838);
and UO_973 (O_973,N_4710,N_4986);
nand UO_974 (O_974,N_4869,N_4880);
nor UO_975 (O_975,N_4554,N_4941);
and UO_976 (O_976,N_4787,N_4755);
nand UO_977 (O_977,N_4515,N_4864);
nor UO_978 (O_978,N_4594,N_4936);
nor UO_979 (O_979,N_4856,N_4598);
and UO_980 (O_980,N_4526,N_4918);
or UO_981 (O_981,N_4671,N_4692);
and UO_982 (O_982,N_4975,N_4744);
or UO_983 (O_983,N_4928,N_4671);
or UO_984 (O_984,N_4986,N_4570);
nand UO_985 (O_985,N_4994,N_4510);
or UO_986 (O_986,N_4886,N_4769);
nand UO_987 (O_987,N_4835,N_4714);
nand UO_988 (O_988,N_4681,N_4673);
or UO_989 (O_989,N_4545,N_4539);
or UO_990 (O_990,N_4563,N_4707);
xor UO_991 (O_991,N_4525,N_4581);
nand UO_992 (O_992,N_4717,N_4662);
nor UO_993 (O_993,N_4628,N_4932);
and UO_994 (O_994,N_4869,N_4944);
nand UO_995 (O_995,N_4603,N_4729);
nor UO_996 (O_996,N_4588,N_4573);
and UO_997 (O_997,N_4542,N_4970);
and UO_998 (O_998,N_4724,N_4510);
nand UO_999 (O_999,N_4932,N_4740);
endmodule