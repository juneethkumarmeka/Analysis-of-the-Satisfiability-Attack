module basic_500_3000_500_40_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_478,In_201);
or U1 (N_1,In_282,In_317);
xnor U2 (N_2,In_474,In_196);
xor U3 (N_3,In_98,In_384);
nor U4 (N_4,In_371,In_159);
nand U5 (N_5,In_482,In_252);
and U6 (N_6,In_111,In_467);
and U7 (N_7,In_119,In_276);
and U8 (N_8,In_149,In_355);
nor U9 (N_9,In_162,In_296);
and U10 (N_10,In_367,In_151);
xor U11 (N_11,In_448,In_408);
nand U12 (N_12,In_433,In_332);
or U13 (N_13,In_163,In_386);
xor U14 (N_14,In_186,In_22);
xor U15 (N_15,In_397,In_146);
or U16 (N_16,In_30,In_182);
and U17 (N_17,In_39,In_280);
nor U18 (N_18,In_166,In_364);
and U19 (N_19,In_285,In_243);
nand U20 (N_20,In_83,In_277);
nor U21 (N_21,In_41,In_54);
nor U22 (N_22,In_379,In_348);
nand U23 (N_23,In_233,In_323);
nor U24 (N_24,In_72,In_164);
nor U25 (N_25,In_158,In_192);
and U26 (N_26,In_475,In_132);
nand U27 (N_27,In_218,In_255);
xor U28 (N_28,In_157,In_87);
xor U29 (N_29,In_264,In_19);
or U30 (N_30,In_291,In_137);
nand U31 (N_31,In_2,In_199);
or U32 (N_32,In_238,In_213);
and U33 (N_33,In_9,In_324);
or U34 (N_34,In_465,In_321);
nor U35 (N_35,In_202,In_357);
or U36 (N_36,In_131,In_183);
or U37 (N_37,In_414,In_17);
or U38 (N_38,In_427,In_155);
nor U39 (N_39,In_256,In_331);
nand U40 (N_40,In_411,In_179);
nor U41 (N_41,In_451,In_14);
nand U42 (N_42,In_13,In_31);
nand U43 (N_43,In_148,In_156);
nor U44 (N_44,In_109,In_405);
xor U45 (N_45,In_229,In_319);
xor U46 (N_46,In_409,In_336);
nand U47 (N_47,In_366,In_191);
and U48 (N_48,In_267,In_140);
and U49 (N_49,In_34,In_128);
and U50 (N_50,In_308,In_175);
and U51 (N_51,In_26,In_413);
and U52 (N_52,In_82,In_426);
nand U53 (N_53,In_365,In_226);
and U54 (N_54,In_292,In_73);
xnor U55 (N_55,In_334,In_37);
or U56 (N_56,In_304,In_310);
and U57 (N_57,In_473,In_124);
nor U58 (N_58,In_372,In_272);
nor U59 (N_59,In_65,In_116);
and U60 (N_60,In_165,In_398);
or U61 (N_61,In_295,In_16);
xor U62 (N_62,In_176,In_198);
xnor U63 (N_63,In_85,In_471);
nor U64 (N_64,In_299,In_376);
nand U65 (N_65,In_139,In_143);
nand U66 (N_66,In_421,In_235);
nand U67 (N_67,In_268,In_358);
and U68 (N_68,In_245,In_187);
nor U69 (N_69,In_265,In_382);
nor U70 (N_70,In_4,In_499);
and U71 (N_71,In_195,In_3);
and U72 (N_72,In_377,In_214);
nand U73 (N_73,In_347,In_300);
nor U74 (N_74,In_350,In_305);
nand U75 (N_75,In_275,In_495);
nor U76 (N_76,In_95,In_286);
nand U77 (N_77,In_106,In_69);
nand U78 (N_78,N_69,In_232);
nand U79 (N_79,N_66,N_25);
nand U80 (N_80,In_101,In_374);
nand U81 (N_81,In_210,In_447);
nand U82 (N_82,In_62,In_328);
and U83 (N_83,In_395,In_211);
and U84 (N_84,In_215,In_28);
and U85 (N_85,In_320,N_54);
or U86 (N_86,In_351,In_112);
and U87 (N_87,N_47,In_220);
nor U88 (N_88,N_23,In_294);
xnor U89 (N_89,In_74,In_240);
nand U90 (N_90,In_25,In_154);
nand U91 (N_91,In_75,In_237);
or U92 (N_92,In_170,In_18);
or U93 (N_93,In_438,In_108);
nand U94 (N_94,In_345,In_407);
nand U95 (N_95,In_78,In_61);
nand U96 (N_96,In_446,In_416);
and U97 (N_97,In_423,In_242);
nand U98 (N_98,In_261,N_52);
nor U99 (N_99,In_488,In_47);
or U100 (N_100,In_429,In_144);
and U101 (N_101,In_129,In_417);
nor U102 (N_102,In_302,In_444);
nand U103 (N_103,In_193,In_346);
nor U104 (N_104,N_36,In_359);
or U105 (N_105,N_18,In_40);
nor U106 (N_106,In_127,In_27);
nor U107 (N_107,In_169,In_53);
nor U108 (N_108,N_32,In_160);
nor U109 (N_109,In_177,In_490);
nand U110 (N_110,N_73,In_466);
nor U111 (N_111,In_392,N_11);
nand U112 (N_112,In_410,In_307);
and U113 (N_113,In_469,In_254);
nor U114 (N_114,In_11,In_388);
nor U115 (N_115,In_221,In_103);
or U116 (N_116,In_477,In_102);
nor U117 (N_117,N_40,N_4);
nor U118 (N_118,In_32,In_418);
nor U119 (N_119,N_5,N_42);
nor U120 (N_120,In_114,In_396);
nand U121 (N_121,In_461,In_262);
nand U122 (N_122,In_208,In_306);
nand U123 (N_123,N_21,N_68);
nand U124 (N_124,In_76,In_441);
nor U125 (N_125,In_203,In_59);
or U126 (N_126,In_455,In_335);
nor U127 (N_127,In_412,In_253);
nand U128 (N_128,In_318,N_26);
nor U129 (N_129,In_0,In_489);
xnor U130 (N_130,In_459,N_65);
or U131 (N_131,In_123,In_250);
or U132 (N_132,In_227,In_216);
or U133 (N_133,In_207,In_230);
nor U134 (N_134,In_244,In_370);
nor U135 (N_135,In_117,In_493);
nor U136 (N_136,In_420,In_204);
nor U137 (N_137,In_309,In_437);
nor U138 (N_138,In_439,In_313);
or U139 (N_139,In_375,In_219);
nand U140 (N_140,In_188,In_273);
nand U141 (N_141,In_147,In_171);
or U142 (N_142,In_452,In_258);
nand U143 (N_143,N_74,N_20);
or U144 (N_144,In_178,In_298);
or U145 (N_145,In_24,In_274);
xnor U146 (N_146,In_209,In_481);
or U147 (N_147,In_297,In_314);
or U148 (N_148,In_15,In_51);
nor U149 (N_149,In_428,In_440);
and U150 (N_150,N_8,In_341);
and U151 (N_151,In_443,In_361);
and U152 (N_152,N_107,In_340);
nor U153 (N_153,N_132,In_20);
and U154 (N_154,In_45,In_404);
nand U155 (N_155,In_1,In_194);
and U156 (N_156,N_81,In_223);
nor U157 (N_157,In_138,In_491);
nand U158 (N_158,In_97,In_168);
xor U159 (N_159,In_432,In_425);
and U160 (N_160,N_115,In_480);
nand U161 (N_161,In_269,In_333);
or U162 (N_162,N_1,In_303);
nor U163 (N_163,In_52,In_167);
or U164 (N_164,N_27,In_94);
xnor U165 (N_165,In_206,N_143);
nand U166 (N_166,N_38,In_81);
nor U167 (N_167,In_121,N_44);
nand U168 (N_168,In_217,N_30);
and U169 (N_169,N_0,In_470);
nand U170 (N_170,In_145,In_284);
nand U171 (N_171,In_435,In_326);
nor U172 (N_172,N_109,N_14);
nor U173 (N_173,In_454,In_249);
xnor U174 (N_174,N_147,In_56);
nand U175 (N_175,In_399,N_106);
or U176 (N_176,In_312,In_290);
nor U177 (N_177,In_184,In_363);
xor U178 (N_178,In_498,In_107);
nor U179 (N_179,N_130,In_100);
nor U180 (N_180,N_97,N_128);
and U181 (N_181,N_80,N_76);
nand U182 (N_182,In_174,In_402);
nor U183 (N_183,In_36,N_95);
and U184 (N_184,N_116,N_135);
nor U185 (N_185,In_7,In_115);
or U186 (N_186,In_360,N_134);
or U187 (N_187,In_301,N_108);
xnor U188 (N_188,N_140,N_55);
nand U189 (N_189,In_63,N_61);
or U190 (N_190,In_181,In_90);
or U191 (N_191,In_391,In_401);
nand U192 (N_192,In_77,In_152);
or U193 (N_193,In_281,In_259);
nand U194 (N_194,In_278,In_60);
and U195 (N_195,In_67,In_105);
and U196 (N_196,In_70,In_125);
nand U197 (N_197,In_368,N_99);
and U198 (N_198,In_86,In_458);
nand U199 (N_199,N_110,In_118);
nand U200 (N_200,In_449,In_38);
xnor U201 (N_201,N_92,In_311);
and U202 (N_202,N_119,In_80);
nand U203 (N_203,In_436,In_173);
and U204 (N_204,N_75,N_88);
nor U205 (N_205,N_22,N_145);
nor U206 (N_206,N_60,In_89);
or U207 (N_207,N_58,N_139);
or U208 (N_208,N_136,In_486);
nand U209 (N_209,In_234,In_492);
and U210 (N_210,In_251,N_120);
nor U211 (N_211,In_29,In_231);
and U212 (N_212,In_380,In_456);
nand U213 (N_213,N_117,N_28);
nor U214 (N_214,In_247,N_43);
or U215 (N_215,In_485,N_91);
and U216 (N_216,In_212,In_394);
and U217 (N_217,N_137,In_450);
and U218 (N_218,In_430,In_354);
xor U219 (N_219,In_96,N_102);
nor U220 (N_220,N_10,N_37);
xor U221 (N_221,N_90,In_316);
and U222 (N_222,N_141,In_150);
or U223 (N_223,N_149,N_84);
xor U224 (N_224,In_55,N_13);
and U225 (N_225,In_43,N_113);
nor U226 (N_226,In_373,In_415);
nand U227 (N_227,N_103,N_39);
nor U228 (N_228,N_183,N_31);
or U229 (N_229,In_49,In_161);
nor U230 (N_230,In_442,In_322);
nor U231 (N_231,N_12,In_189);
or U232 (N_232,N_2,In_241);
nor U233 (N_233,N_87,In_141);
nand U234 (N_234,N_181,N_133);
nor U235 (N_235,N_129,N_173);
and U236 (N_236,N_78,In_271);
nor U237 (N_237,In_21,In_113);
nand U238 (N_238,N_112,In_224);
or U239 (N_239,In_288,N_178);
nand U240 (N_240,In_494,N_212);
and U241 (N_241,N_192,N_89);
and U242 (N_242,In_330,In_44);
nor U243 (N_243,In_344,N_163);
nand U244 (N_244,N_124,N_138);
nor U245 (N_245,N_53,In_134);
xor U246 (N_246,N_172,N_101);
or U247 (N_247,In_228,In_135);
or U248 (N_248,In_66,N_156);
or U249 (N_249,N_203,N_41);
nor U250 (N_250,N_50,In_205);
nand U251 (N_251,In_246,In_389);
nand U252 (N_252,N_59,N_209);
or U253 (N_253,N_49,N_67);
nor U254 (N_254,In_431,N_114);
nand U255 (N_255,N_123,N_16);
nor U256 (N_256,N_190,N_144);
xnor U257 (N_257,N_3,In_383);
xnor U258 (N_258,N_56,In_479);
nor U259 (N_259,In_185,In_369);
nor U260 (N_260,N_177,In_239);
or U261 (N_261,In_325,In_287);
and U262 (N_262,In_356,In_487);
and U263 (N_263,N_207,In_362);
or U264 (N_264,In_248,In_79);
or U265 (N_265,In_279,N_19);
nand U266 (N_266,N_154,N_94);
nor U267 (N_267,N_180,N_62);
xnor U268 (N_268,N_83,N_48);
nor U269 (N_269,N_17,In_353);
or U270 (N_270,N_175,In_422);
nand U271 (N_271,N_57,In_483);
and U272 (N_272,N_213,N_222);
nor U273 (N_273,In_257,In_484);
nor U274 (N_274,N_195,N_142);
and U275 (N_275,N_34,In_476);
nor U276 (N_276,N_202,N_77);
nand U277 (N_277,N_169,In_381);
nand U278 (N_278,In_120,N_111);
or U279 (N_279,N_205,In_91);
and U280 (N_280,N_131,N_9);
nor U281 (N_281,N_200,N_185);
or U282 (N_282,In_349,In_153);
nand U283 (N_283,In_197,In_460);
or U284 (N_284,N_161,N_118);
nor U285 (N_285,In_68,N_164);
nor U286 (N_286,In_46,In_462);
and U287 (N_287,In_6,N_179);
nor U288 (N_288,N_86,N_197);
nand U289 (N_289,In_180,N_170);
nand U290 (N_290,N_220,In_64);
nand U291 (N_291,In_126,N_33);
nor U292 (N_292,N_150,N_127);
nor U293 (N_293,N_171,N_165);
nand U294 (N_294,N_218,N_166);
nor U295 (N_295,In_23,In_50);
and U296 (N_296,N_122,N_79);
nor U297 (N_297,In_387,In_58);
nand U298 (N_298,N_121,In_342);
nor U299 (N_299,N_146,N_187);
or U300 (N_300,N_196,In_385);
nor U301 (N_301,N_250,In_339);
nand U302 (N_302,In_110,N_290);
nand U303 (N_303,N_215,N_208);
and U304 (N_304,In_8,N_206);
nand U305 (N_305,In_406,N_63);
xor U306 (N_306,N_6,In_457);
nor U307 (N_307,N_184,In_10);
or U308 (N_308,N_125,In_266);
nand U309 (N_309,N_275,In_445);
xor U310 (N_310,N_280,In_130);
and U311 (N_311,In_92,N_232);
nand U312 (N_312,N_189,N_228);
nor U313 (N_313,N_153,N_285);
nand U314 (N_314,N_298,N_223);
nand U315 (N_315,N_289,N_274);
and U316 (N_316,N_260,N_263);
or U317 (N_317,In_434,N_45);
and U318 (N_318,N_231,In_289);
nand U319 (N_319,N_72,N_188);
and U320 (N_320,In_293,In_263);
nand U321 (N_321,N_265,N_241);
nand U322 (N_322,N_258,N_227);
nand U323 (N_323,N_162,N_35);
and U324 (N_324,In_327,In_104);
nor U325 (N_325,In_142,N_29);
nand U326 (N_326,N_254,N_225);
or U327 (N_327,In_352,N_229);
or U328 (N_328,In_393,N_226);
and U329 (N_329,In_35,N_148);
nor U330 (N_330,N_159,N_221);
nand U331 (N_331,N_191,N_291);
nor U332 (N_332,N_247,N_255);
nand U333 (N_333,N_251,In_270);
nand U334 (N_334,N_211,N_268);
xor U335 (N_335,In_464,N_186);
xor U336 (N_336,N_279,In_84);
or U337 (N_337,N_64,N_270);
or U338 (N_338,In_343,N_176);
and U339 (N_339,In_338,N_267);
nand U340 (N_340,N_104,N_204);
or U341 (N_341,N_256,In_463);
nand U342 (N_342,In_33,N_157);
and U343 (N_343,In_225,N_82);
nor U344 (N_344,N_214,N_71);
xnor U345 (N_345,N_234,N_168);
or U346 (N_346,N_239,In_48);
and U347 (N_347,N_277,N_46);
nand U348 (N_348,N_160,N_155);
nor U349 (N_349,N_278,N_242);
nand U350 (N_350,In_400,N_51);
nand U351 (N_351,In_496,In_172);
nor U352 (N_352,N_299,N_243);
or U353 (N_353,In_88,N_24);
xor U354 (N_354,In_136,N_288);
and U355 (N_355,N_266,N_284);
nand U356 (N_356,In_283,N_262);
and U357 (N_357,N_235,N_272);
nor U358 (N_358,N_273,N_193);
and U359 (N_359,N_219,In_378);
nor U360 (N_360,N_167,In_42);
nor U361 (N_361,N_253,In_329);
nor U362 (N_362,N_98,N_93);
and U363 (N_363,N_216,N_264);
and U364 (N_364,N_126,In_260);
or U365 (N_365,In_5,N_100);
nor U366 (N_366,N_257,N_158);
or U367 (N_367,In_497,In_93);
nand U368 (N_368,N_182,N_233);
nor U369 (N_369,In_472,N_230);
nor U370 (N_370,N_246,N_85);
xnor U371 (N_371,In_57,N_194);
or U372 (N_372,N_281,In_12);
nor U373 (N_373,N_15,N_217);
or U374 (N_374,N_7,N_295);
nand U375 (N_375,N_312,N_244);
nor U376 (N_376,N_319,N_302);
and U377 (N_377,N_96,N_340);
nand U378 (N_378,N_338,N_346);
xor U379 (N_379,N_337,In_222);
nor U380 (N_380,In_390,N_306);
nor U381 (N_381,N_366,In_315);
nor U382 (N_382,N_283,In_200);
nor U383 (N_383,N_318,N_323);
or U384 (N_384,N_339,N_343);
and U385 (N_385,N_301,N_345);
xnor U386 (N_386,N_348,N_259);
nor U387 (N_387,In_236,N_330);
and U388 (N_388,N_350,N_252);
nor U389 (N_389,N_365,N_307);
or U390 (N_390,N_333,N_363);
nand U391 (N_391,N_370,N_336);
nor U392 (N_392,N_362,N_334);
and U393 (N_393,N_357,N_356);
and U394 (N_394,N_311,N_271);
nor U395 (N_395,N_198,N_248);
or U396 (N_396,N_368,N_369);
and U397 (N_397,N_351,N_315);
or U398 (N_398,N_210,N_358);
nand U399 (N_399,N_317,N_261);
or U400 (N_400,N_374,N_371);
xnor U401 (N_401,N_372,N_294);
nand U402 (N_402,N_364,N_314);
nor U403 (N_403,N_325,N_322);
or U404 (N_404,N_324,N_249);
and U405 (N_405,N_297,N_70);
and U406 (N_406,N_310,N_329);
or U407 (N_407,N_353,N_326);
nor U408 (N_408,N_335,In_453);
nand U409 (N_409,N_305,N_240);
or U410 (N_410,N_300,N_308);
or U411 (N_411,N_359,N_332);
xor U412 (N_412,In_71,N_352);
nor U413 (N_413,N_344,N_349);
xnor U414 (N_414,N_152,N_292);
and U415 (N_415,N_296,N_328);
nand U416 (N_416,In_99,N_287);
nor U417 (N_417,N_237,N_327);
xor U418 (N_418,N_151,N_342);
and U419 (N_419,In_190,N_293);
nand U420 (N_420,N_321,N_341);
and U421 (N_421,N_224,In_424);
nand U422 (N_422,N_354,N_304);
or U423 (N_423,N_316,N_303);
nand U424 (N_424,N_201,In_403);
or U425 (N_425,N_199,N_320);
or U426 (N_426,N_269,N_174);
xnor U427 (N_427,N_282,In_419);
nor U428 (N_428,N_360,In_133);
nand U429 (N_429,N_355,In_468);
or U430 (N_430,N_373,N_238);
nor U431 (N_431,N_347,In_337);
xnor U432 (N_432,N_367,N_309);
or U433 (N_433,N_313,N_276);
nand U434 (N_434,N_361,N_236);
and U435 (N_435,N_331,N_286);
nor U436 (N_436,In_122,N_245);
nor U437 (N_437,N_105,N_306);
nor U438 (N_438,N_320,In_453);
nor U439 (N_439,N_354,N_320);
or U440 (N_440,N_238,N_342);
and U441 (N_441,N_151,N_313);
nor U442 (N_442,In_419,N_323);
and U443 (N_443,N_335,N_201);
or U444 (N_444,N_321,N_339);
nand U445 (N_445,N_301,N_297);
xnor U446 (N_446,N_301,N_372);
and U447 (N_447,In_390,N_374);
nand U448 (N_448,In_236,N_276);
or U449 (N_449,In_222,N_152);
or U450 (N_450,N_389,N_381);
nand U451 (N_451,N_445,N_429);
nand U452 (N_452,N_405,N_416);
nor U453 (N_453,N_414,N_427);
nand U454 (N_454,N_379,N_431);
and U455 (N_455,N_421,N_396);
or U456 (N_456,N_391,N_438);
xnor U457 (N_457,N_384,N_388);
and U458 (N_458,N_444,N_432);
nor U459 (N_459,N_404,N_440);
or U460 (N_460,N_376,N_428);
xor U461 (N_461,N_383,N_378);
and U462 (N_462,N_401,N_375);
and U463 (N_463,N_393,N_382);
nand U464 (N_464,N_402,N_386);
and U465 (N_465,N_422,N_394);
nand U466 (N_466,N_392,N_434);
nor U467 (N_467,N_433,N_439);
or U468 (N_468,N_447,N_413);
nor U469 (N_469,N_448,N_412);
xor U470 (N_470,N_406,N_436);
nand U471 (N_471,N_403,N_387);
or U472 (N_472,N_442,N_420);
nand U473 (N_473,N_400,N_417);
nor U474 (N_474,N_377,N_449);
or U475 (N_475,N_426,N_415);
nand U476 (N_476,N_409,N_441);
nor U477 (N_477,N_380,N_423);
nand U478 (N_478,N_395,N_425);
or U479 (N_479,N_398,N_410);
xnor U480 (N_480,N_437,N_419);
and U481 (N_481,N_408,N_399);
nand U482 (N_482,N_424,N_430);
nor U483 (N_483,N_390,N_407);
or U484 (N_484,N_385,N_446);
or U485 (N_485,N_418,N_411);
nand U486 (N_486,N_443,N_435);
nor U487 (N_487,N_397,N_422);
nand U488 (N_488,N_404,N_434);
or U489 (N_489,N_430,N_415);
nand U490 (N_490,N_380,N_378);
or U491 (N_491,N_436,N_418);
and U492 (N_492,N_439,N_443);
nand U493 (N_493,N_413,N_384);
nor U494 (N_494,N_439,N_386);
or U495 (N_495,N_406,N_396);
nand U496 (N_496,N_416,N_430);
nor U497 (N_497,N_400,N_389);
nand U498 (N_498,N_429,N_415);
or U499 (N_499,N_409,N_417);
nand U500 (N_500,N_391,N_381);
xor U501 (N_501,N_425,N_408);
nor U502 (N_502,N_437,N_415);
nand U503 (N_503,N_400,N_406);
or U504 (N_504,N_415,N_402);
nor U505 (N_505,N_439,N_407);
nand U506 (N_506,N_442,N_419);
xnor U507 (N_507,N_448,N_424);
or U508 (N_508,N_438,N_418);
and U509 (N_509,N_410,N_412);
or U510 (N_510,N_406,N_383);
nand U511 (N_511,N_389,N_402);
nand U512 (N_512,N_417,N_437);
nor U513 (N_513,N_428,N_382);
xor U514 (N_514,N_436,N_447);
nand U515 (N_515,N_377,N_398);
and U516 (N_516,N_407,N_399);
nand U517 (N_517,N_398,N_434);
or U518 (N_518,N_448,N_391);
and U519 (N_519,N_419,N_449);
nor U520 (N_520,N_423,N_441);
or U521 (N_521,N_415,N_431);
and U522 (N_522,N_421,N_432);
nand U523 (N_523,N_423,N_419);
nor U524 (N_524,N_394,N_431);
or U525 (N_525,N_504,N_460);
or U526 (N_526,N_463,N_523);
and U527 (N_527,N_479,N_485);
or U528 (N_528,N_467,N_509);
or U529 (N_529,N_499,N_517);
nor U530 (N_530,N_472,N_494);
and U531 (N_531,N_461,N_511);
nor U532 (N_532,N_512,N_491);
nor U533 (N_533,N_468,N_458);
or U534 (N_534,N_508,N_484);
or U535 (N_535,N_462,N_521);
and U536 (N_536,N_505,N_454);
xnor U537 (N_537,N_497,N_510);
and U538 (N_538,N_486,N_475);
or U539 (N_539,N_520,N_513);
and U540 (N_540,N_492,N_481);
xor U541 (N_541,N_466,N_518);
nor U542 (N_542,N_498,N_465);
or U543 (N_543,N_487,N_483);
or U544 (N_544,N_515,N_471);
nor U545 (N_545,N_476,N_477);
nor U546 (N_546,N_503,N_524);
or U547 (N_547,N_522,N_516);
or U548 (N_548,N_459,N_456);
nand U549 (N_549,N_474,N_489);
xor U550 (N_550,N_500,N_464);
nor U551 (N_551,N_452,N_478);
nand U552 (N_552,N_490,N_470);
and U553 (N_553,N_514,N_507);
or U554 (N_554,N_455,N_451);
or U555 (N_555,N_480,N_469);
and U556 (N_556,N_473,N_501);
xnor U557 (N_557,N_482,N_496);
or U558 (N_558,N_519,N_495);
nand U559 (N_559,N_457,N_502);
and U560 (N_560,N_488,N_453);
xnor U561 (N_561,N_450,N_493);
nor U562 (N_562,N_506,N_463);
or U563 (N_563,N_470,N_511);
and U564 (N_564,N_506,N_473);
or U565 (N_565,N_457,N_511);
nand U566 (N_566,N_459,N_453);
or U567 (N_567,N_488,N_469);
nor U568 (N_568,N_507,N_478);
xnor U569 (N_569,N_512,N_470);
or U570 (N_570,N_508,N_520);
nand U571 (N_571,N_475,N_465);
nand U572 (N_572,N_494,N_514);
and U573 (N_573,N_470,N_505);
nor U574 (N_574,N_455,N_499);
or U575 (N_575,N_498,N_462);
nand U576 (N_576,N_459,N_457);
nand U577 (N_577,N_474,N_523);
and U578 (N_578,N_501,N_455);
xor U579 (N_579,N_508,N_516);
and U580 (N_580,N_471,N_495);
and U581 (N_581,N_521,N_457);
xnor U582 (N_582,N_459,N_512);
nand U583 (N_583,N_516,N_523);
xor U584 (N_584,N_483,N_471);
or U585 (N_585,N_505,N_497);
nand U586 (N_586,N_490,N_524);
nor U587 (N_587,N_478,N_454);
nand U588 (N_588,N_519,N_491);
nand U589 (N_589,N_522,N_484);
nor U590 (N_590,N_473,N_491);
nor U591 (N_591,N_487,N_481);
nor U592 (N_592,N_483,N_478);
xnor U593 (N_593,N_515,N_522);
and U594 (N_594,N_459,N_483);
nor U595 (N_595,N_477,N_491);
nor U596 (N_596,N_502,N_516);
xor U597 (N_597,N_523,N_511);
nor U598 (N_598,N_461,N_459);
nand U599 (N_599,N_459,N_510);
nand U600 (N_600,N_541,N_593);
nor U601 (N_601,N_545,N_531);
xor U602 (N_602,N_590,N_583);
nand U603 (N_603,N_571,N_586);
nand U604 (N_604,N_562,N_559);
and U605 (N_605,N_560,N_575);
and U606 (N_606,N_556,N_538);
or U607 (N_607,N_550,N_546);
xor U608 (N_608,N_529,N_533);
and U609 (N_609,N_567,N_554);
nor U610 (N_610,N_569,N_558);
nor U611 (N_611,N_535,N_599);
and U612 (N_612,N_580,N_551);
nand U613 (N_613,N_592,N_579);
or U614 (N_614,N_542,N_528);
nand U615 (N_615,N_587,N_594);
and U616 (N_616,N_591,N_588);
nor U617 (N_617,N_534,N_539);
and U618 (N_618,N_584,N_530);
and U619 (N_619,N_540,N_564);
or U620 (N_620,N_598,N_574);
nor U621 (N_621,N_537,N_536);
nor U622 (N_622,N_548,N_585);
nand U623 (N_623,N_570,N_572);
nand U624 (N_624,N_589,N_596);
nor U625 (N_625,N_555,N_595);
nor U626 (N_626,N_566,N_557);
nor U627 (N_627,N_581,N_578);
nor U628 (N_628,N_552,N_544);
nand U629 (N_629,N_553,N_526);
nor U630 (N_630,N_543,N_582);
or U631 (N_631,N_573,N_568);
or U632 (N_632,N_597,N_527);
nand U633 (N_633,N_561,N_525);
and U634 (N_634,N_549,N_565);
or U635 (N_635,N_547,N_577);
or U636 (N_636,N_576,N_532);
nand U637 (N_637,N_563,N_561);
nand U638 (N_638,N_583,N_572);
or U639 (N_639,N_594,N_583);
nand U640 (N_640,N_525,N_576);
nor U641 (N_641,N_568,N_553);
nand U642 (N_642,N_526,N_585);
and U643 (N_643,N_543,N_583);
nand U644 (N_644,N_596,N_541);
nand U645 (N_645,N_581,N_540);
nand U646 (N_646,N_567,N_540);
and U647 (N_647,N_592,N_599);
nor U648 (N_648,N_574,N_581);
and U649 (N_649,N_592,N_526);
nor U650 (N_650,N_598,N_536);
nor U651 (N_651,N_551,N_525);
or U652 (N_652,N_561,N_577);
nand U653 (N_653,N_594,N_569);
nand U654 (N_654,N_598,N_554);
nor U655 (N_655,N_540,N_580);
nand U656 (N_656,N_539,N_560);
or U657 (N_657,N_595,N_575);
and U658 (N_658,N_527,N_578);
or U659 (N_659,N_574,N_552);
nor U660 (N_660,N_535,N_543);
nand U661 (N_661,N_531,N_566);
xor U662 (N_662,N_599,N_528);
nor U663 (N_663,N_568,N_577);
or U664 (N_664,N_598,N_560);
xnor U665 (N_665,N_581,N_529);
or U666 (N_666,N_586,N_548);
xor U667 (N_667,N_593,N_571);
nand U668 (N_668,N_552,N_577);
nand U669 (N_669,N_546,N_530);
or U670 (N_670,N_525,N_527);
nor U671 (N_671,N_590,N_539);
xnor U672 (N_672,N_580,N_565);
and U673 (N_673,N_571,N_543);
or U674 (N_674,N_529,N_587);
nand U675 (N_675,N_635,N_605);
nor U676 (N_676,N_613,N_626);
or U677 (N_677,N_659,N_620);
nor U678 (N_678,N_623,N_636);
and U679 (N_679,N_640,N_603);
nor U680 (N_680,N_602,N_662);
nor U681 (N_681,N_665,N_646);
and U682 (N_682,N_604,N_651);
nor U683 (N_683,N_628,N_617);
and U684 (N_684,N_648,N_601);
nand U685 (N_685,N_647,N_629);
and U686 (N_686,N_667,N_672);
nor U687 (N_687,N_664,N_632);
nor U688 (N_688,N_666,N_600);
and U689 (N_689,N_649,N_621);
nand U690 (N_690,N_650,N_614);
nand U691 (N_691,N_637,N_643);
or U692 (N_692,N_634,N_656);
or U693 (N_693,N_616,N_663);
nand U694 (N_694,N_627,N_660);
nor U695 (N_695,N_609,N_624);
and U696 (N_696,N_652,N_608);
nand U697 (N_697,N_661,N_668);
or U698 (N_698,N_655,N_618);
nor U699 (N_699,N_639,N_630);
xor U700 (N_700,N_669,N_670);
nand U701 (N_701,N_645,N_611);
and U702 (N_702,N_644,N_631);
or U703 (N_703,N_657,N_610);
nand U704 (N_704,N_674,N_612);
nand U705 (N_705,N_615,N_671);
and U706 (N_706,N_653,N_625);
nand U707 (N_707,N_622,N_633);
or U708 (N_708,N_641,N_658);
nor U709 (N_709,N_606,N_673);
nand U710 (N_710,N_619,N_607);
and U711 (N_711,N_638,N_654);
or U712 (N_712,N_642,N_646);
or U713 (N_713,N_627,N_666);
nand U714 (N_714,N_666,N_642);
nor U715 (N_715,N_661,N_615);
and U716 (N_716,N_638,N_652);
nor U717 (N_717,N_601,N_632);
nand U718 (N_718,N_673,N_612);
and U719 (N_719,N_617,N_647);
nand U720 (N_720,N_604,N_606);
and U721 (N_721,N_645,N_651);
nor U722 (N_722,N_644,N_672);
and U723 (N_723,N_606,N_633);
xor U724 (N_724,N_669,N_658);
and U725 (N_725,N_640,N_643);
and U726 (N_726,N_610,N_666);
or U727 (N_727,N_641,N_627);
nand U728 (N_728,N_652,N_618);
and U729 (N_729,N_609,N_623);
and U730 (N_730,N_643,N_659);
or U731 (N_731,N_627,N_639);
and U732 (N_732,N_643,N_657);
nand U733 (N_733,N_657,N_617);
nor U734 (N_734,N_643,N_639);
nor U735 (N_735,N_648,N_625);
and U736 (N_736,N_666,N_645);
nor U737 (N_737,N_624,N_662);
and U738 (N_738,N_639,N_607);
or U739 (N_739,N_649,N_607);
nand U740 (N_740,N_628,N_661);
or U741 (N_741,N_672,N_654);
and U742 (N_742,N_645,N_621);
or U743 (N_743,N_617,N_608);
nand U744 (N_744,N_602,N_600);
and U745 (N_745,N_622,N_658);
and U746 (N_746,N_650,N_670);
nand U747 (N_747,N_647,N_638);
and U748 (N_748,N_647,N_643);
nand U749 (N_749,N_646,N_620);
or U750 (N_750,N_749,N_677);
and U751 (N_751,N_708,N_685);
and U752 (N_752,N_713,N_683);
nand U753 (N_753,N_746,N_701);
nor U754 (N_754,N_707,N_734);
nand U755 (N_755,N_699,N_735);
or U756 (N_756,N_748,N_730);
nand U757 (N_757,N_698,N_747);
and U758 (N_758,N_676,N_709);
nand U759 (N_759,N_724,N_678);
or U760 (N_760,N_681,N_731);
and U761 (N_761,N_736,N_738);
xnor U762 (N_762,N_718,N_702);
nand U763 (N_763,N_722,N_726);
or U764 (N_764,N_723,N_728);
xor U765 (N_765,N_680,N_682);
and U766 (N_766,N_740,N_689);
nand U767 (N_767,N_732,N_706);
and U768 (N_768,N_696,N_727);
nand U769 (N_769,N_743,N_692);
or U770 (N_770,N_687,N_714);
nor U771 (N_771,N_711,N_729);
and U772 (N_772,N_691,N_716);
and U773 (N_773,N_705,N_717);
or U774 (N_774,N_712,N_675);
nand U775 (N_775,N_737,N_688);
nor U776 (N_776,N_684,N_725);
nor U777 (N_777,N_690,N_686);
or U778 (N_778,N_694,N_744);
xnor U779 (N_779,N_695,N_720);
nand U780 (N_780,N_719,N_745);
xnor U781 (N_781,N_715,N_697);
and U782 (N_782,N_739,N_703);
or U783 (N_783,N_679,N_704);
nand U784 (N_784,N_700,N_710);
nand U785 (N_785,N_742,N_741);
nor U786 (N_786,N_721,N_693);
nand U787 (N_787,N_733,N_702);
nor U788 (N_788,N_733,N_684);
or U789 (N_789,N_747,N_717);
nand U790 (N_790,N_680,N_712);
or U791 (N_791,N_690,N_719);
and U792 (N_792,N_747,N_731);
xor U793 (N_793,N_701,N_691);
or U794 (N_794,N_709,N_691);
and U795 (N_795,N_728,N_678);
nor U796 (N_796,N_709,N_690);
xor U797 (N_797,N_702,N_706);
nand U798 (N_798,N_687,N_730);
nand U799 (N_799,N_743,N_688);
or U800 (N_800,N_680,N_733);
or U801 (N_801,N_718,N_694);
nor U802 (N_802,N_698,N_735);
nand U803 (N_803,N_702,N_741);
and U804 (N_804,N_704,N_718);
and U805 (N_805,N_746,N_738);
or U806 (N_806,N_681,N_704);
and U807 (N_807,N_691,N_736);
or U808 (N_808,N_711,N_726);
nand U809 (N_809,N_749,N_742);
and U810 (N_810,N_715,N_737);
xor U811 (N_811,N_737,N_697);
nor U812 (N_812,N_685,N_717);
nor U813 (N_813,N_730,N_707);
or U814 (N_814,N_724,N_702);
and U815 (N_815,N_676,N_696);
nor U816 (N_816,N_677,N_715);
and U817 (N_817,N_722,N_689);
xnor U818 (N_818,N_701,N_709);
nand U819 (N_819,N_697,N_729);
nand U820 (N_820,N_716,N_676);
and U821 (N_821,N_738,N_717);
and U822 (N_822,N_719,N_744);
and U823 (N_823,N_698,N_738);
nor U824 (N_824,N_718,N_697);
or U825 (N_825,N_808,N_762);
nand U826 (N_826,N_780,N_760);
or U827 (N_827,N_788,N_761);
xnor U828 (N_828,N_815,N_805);
nor U829 (N_829,N_811,N_810);
nor U830 (N_830,N_809,N_754);
nand U831 (N_831,N_786,N_803);
and U832 (N_832,N_814,N_763);
or U833 (N_833,N_776,N_751);
nor U834 (N_834,N_822,N_784);
or U835 (N_835,N_792,N_812);
nor U836 (N_836,N_806,N_782);
nor U837 (N_837,N_774,N_773);
or U838 (N_838,N_801,N_756);
nor U839 (N_839,N_785,N_793);
nor U840 (N_840,N_771,N_796);
xor U841 (N_841,N_781,N_816);
nor U842 (N_842,N_753,N_787);
xnor U843 (N_843,N_807,N_798);
nor U844 (N_844,N_772,N_821);
or U845 (N_845,N_804,N_797);
xnor U846 (N_846,N_818,N_824);
nand U847 (N_847,N_777,N_783);
and U848 (N_848,N_752,N_779);
xnor U849 (N_849,N_757,N_769);
nand U850 (N_850,N_800,N_759);
and U851 (N_851,N_770,N_819);
xnor U852 (N_852,N_758,N_791);
and U853 (N_853,N_802,N_750);
xor U854 (N_854,N_820,N_765);
and U855 (N_855,N_768,N_794);
nand U856 (N_856,N_775,N_799);
or U857 (N_857,N_755,N_790);
nor U858 (N_858,N_778,N_817);
nor U859 (N_859,N_823,N_789);
or U860 (N_860,N_813,N_767);
nand U861 (N_861,N_795,N_766);
nor U862 (N_862,N_764,N_823);
and U863 (N_863,N_797,N_758);
or U864 (N_864,N_767,N_784);
nor U865 (N_865,N_756,N_808);
nor U866 (N_866,N_793,N_808);
and U867 (N_867,N_800,N_779);
and U868 (N_868,N_760,N_809);
or U869 (N_869,N_799,N_800);
xnor U870 (N_870,N_818,N_758);
nand U871 (N_871,N_784,N_763);
xnor U872 (N_872,N_804,N_759);
and U873 (N_873,N_820,N_811);
nor U874 (N_874,N_815,N_763);
and U875 (N_875,N_761,N_775);
or U876 (N_876,N_751,N_818);
nor U877 (N_877,N_768,N_767);
nor U878 (N_878,N_771,N_770);
and U879 (N_879,N_772,N_799);
xor U880 (N_880,N_777,N_776);
nand U881 (N_881,N_816,N_797);
or U882 (N_882,N_811,N_769);
nor U883 (N_883,N_789,N_816);
nor U884 (N_884,N_794,N_783);
nand U885 (N_885,N_823,N_779);
nor U886 (N_886,N_792,N_791);
or U887 (N_887,N_800,N_803);
or U888 (N_888,N_775,N_801);
and U889 (N_889,N_782,N_800);
or U890 (N_890,N_816,N_756);
nand U891 (N_891,N_802,N_766);
nor U892 (N_892,N_818,N_814);
and U893 (N_893,N_757,N_810);
or U894 (N_894,N_752,N_766);
nor U895 (N_895,N_810,N_781);
nor U896 (N_896,N_782,N_808);
nor U897 (N_897,N_758,N_768);
and U898 (N_898,N_752,N_758);
and U899 (N_899,N_810,N_775);
or U900 (N_900,N_892,N_893);
and U901 (N_901,N_847,N_837);
nand U902 (N_902,N_859,N_876);
nor U903 (N_903,N_848,N_860);
and U904 (N_904,N_866,N_826);
and U905 (N_905,N_889,N_865);
nor U906 (N_906,N_838,N_899);
or U907 (N_907,N_835,N_861);
and U908 (N_908,N_845,N_862);
and U909 (N_909,N_831,N_842);
or U910 (N_910,N_884,N_843);
nor U911 (N_911,N_825,N_897);
or U912 (N_912,N_834,N_871);
nor U913 (N_913,N_858,N_857);
nor U914 (N_914,N_878,N_891);
or U915 (N_915,N_853,N_832);
nor U916 (N_916,N_856,N_875);
xnor U917 (N_917,N_887,N_827);
nand U918 (N_918,N_886,N_872);
or U919 (N_919,N_868,N_880);
nor U920 (N_920,N_894,N_883);
nand U921 (N_921,N_885,N_881);
or U922 (N_922,N_895,N_864);
nand U923 (N_923,N_888,N_890);
nor U924 (N_924,N_849,N_898);
or U925 (N_925,N_877,N_844);
or U926 (N_926,N_851,N_850);
nor U927 (N_927,N_833,N_869);
or U928 (N_928,N_846,N_829);
and U929 (N_929,N_896,N_836);
and U930 (N_930,N_828,N_873);
and U931 (N_931,N_839,N_852);
nor U932 (N_932,N_867,N_879);
nor U933 (N_933,N_874,N_840);
nand U934 (N_934,N_855,N_830);
nand U935 (N_935,N_854,N_882);
or U936 (N_936,N_863,N_841);
nor U937 (N_937,N_870,N_887);
and U938 (N_938,N_831,N_856);
xnor U939 (N_939,N_874,N_853);
nand U940 (N_940,N_825,N_878);
nor U941 (N_941,N_843,N_845);
or U942 (N_942,N_892,N_845);
xor U943 (N_943,N_834,N_864);
and U944 (N_944,N_843,N_827);
xnor U945 (N_945,N_844,N_842);
nor U946 (N_946,N_831,N_845);
xnor U947 (N_947,N_848,N_831);
nor U948 (N_948,N_839,N_863);
or U949 (N_949,N_874,N_865);
nor U950 (N_950,N_868,N_858);
nor U951 (N_951,N_881,N_889);
or U952 (N_952,N_838,N_847);
xor U953 (N_953,N_841,N_877);
nor U954 (N_954,N_882,N_893);
or U955 (N_955,N_842,N_882);
xor U956 (N_956,N_859,N_847);
nor U957 (N_957,N_879,N_891);
and U958 (N_958,N_827,N_842);
and U959 (N_959,N_828,N_857);
and U960 (N_960,N_880,N_886);
xnor U961 (N_961,N_893,N_826);
or U962 (N_962,N_870,N_895);
nor U963 (N_963,N_830,N_834);
or U964 (N_964,N_860,N_847);
xor U965 (N_965,N_861,N_863);
and U966 (N_966,N_890,N_837);
and U967 (N_967,N_841,N_888);
nor U968 (N_968,N_863,N_832);
nand U969 (N_969,N_853,N_847);
nand U970 (N_970,N_860,N_864);
nand U971 (N_971,N_838,N_869);
nor U972 (N_972,N_888,N_835);
or U973 (N_973,N_884,N_858);
nor U974 (N_974,N_836,N_883);
nand U975 (N_975,N_942,N_956);
and U976 (N_976,N_968,N_917);
or U977 (N_977,N_902,N_931);
nor U978 (N_978,N_904,N_954);
or U979 (N_979,N_903,N_906);
nor U980 (N_980,N_939,N_913);
and U981 (N_981,N_914,N_929);
nor U982 (N_982,N_951,N_947);
and U983 (N_983,N_952,N_948);
nand U984 (N_984,N_972,N_927);
and U985 (N_985,N_959,N_950);
or U986 (N_986,N_966,N_928);
or U987 (N_987,N_930,N_964);
xnor U988 (N_988,N_953,N_961);
xor U989 (N_989,N_936,N_923);
or U990 (N_990,N_900,N_940);
or U991 (N_991,N_958,N_925);
and U992 (N_992,N_949,N_965);
nand U993 (N_993,N_916,N_967);
nand U994 (N_994,N_907,N_970);
and U995 (N_995,N_901,N_915);
or U996 (N_996,N_919,N_973);
and U997 (N_997,N_908,N_920);
and U998 (N_998,N_905,N_938);
xor U999 (N_999,N_943,N_941);
nand U1000 (N_1000,N_924,N_918);
nand U1001 (N_1001,N_911,N_969);
or U1002 (N_1002,N_937,N_910);
and U1003 (N_1003,N_921,N_932);
nand U1004 (N_1004,N_971,N_935);
and U1005 (N_1005,N_946,N_974);
xor U1006 (N_1006,N_960,N_922);
and U1007 (N_1007,N_934,N_912);
and U1008 (N_1008,N_963,N_933);
nor U1009 (N_1009,N_955,N_962);
and U1010 (N_1010,N_945,N_957);
xnor U1011 (N_1011,N_909,N_926);
nor U1012 (N_1012,N_944,N_968);
nand U1013 (N_1013,N_913,N_917);
nor U1014 (N_1014,N_958,N_905);
nand U1015 (N_1015,N_912,N_944);
nor U1016 (N_1016,N_934,N_939);
nor U1017 (N_1017,N_920,N_973);
or U1018 (N_1018,N_940,N_906);
or U1019 (N_1019,N_924,N_973);
nand U1020 (N_1020,N_934,N_913);
or U1021 (N_1021,N_901,N_918);
nand U1022 (N_1022,N_955,N_973);
and U1023 (N_1023,N_974,N_907);
or U1024 (N_1024,N_969,N_964);
or U1025 (N_1025,N_950,N_903);
and U1026 (N_1026,N_908,N_933);
nor U1027 (N_1027,N_928,N_947);
nand U1028 (N_1028,N_947,N_931);
and U1029 (N_1029,N_921,N_945);
nand U1030 (N_1030,N_925,N_956);
and U1031 (N_1031,N_900,N_928);
or U1032 (N_1032,N_939,N_938);
nand U1033 (N_1033,N_902,N_932);
nand U1034 (N_1034,N_901,N_919);
nand U1035 (N_1035,N_930,N_927);
or U1036 (N_1036,N_930,N_952);
nor U1037 (N_1037,N_934,N_963);
nand U1038 (N_1038,N_901,N_920);
nor U1039 (N_1039,N_927,N_960);
and U1040 (N_1040,N_963,N_943);
and U1041 (N_1041,N_927,N_901);
nand U1042 (N_1042,N_958,N_912);
nor U1043 (N_1043,N_944,N_929);
and U1044 (N_1044,N_930,N_948);
and U1045 (N_1045,N_945,N_931);
xor U1046 (N_1046,N_925,N_937);
or U1047 (N_1047,N_957,N_933);
and U1048 (N_1048,N_972,N_931);
nor U1049 (N_1049,N_913,N_943);
nor U1050 (N_1050,N_1017,N_1023);
nor U1051 (N_1051,N_1013,N_1047);
nand U1052 (N_1052,N_998,N_1005);
nor U1053 (N_1053,N_992,N_991);
and U1054 (N_1054,N_996,N_1043);
xnor U1055 (N_1055,N_1008,N_988);
nor U1056 (N_1056,N_1015,N_1039);
nand U1057 (N_1057,N_1012,N_1027);
nor U1058 (N_1058,N_1024,N_1003);
nand U1059 (N_1059,N_1021,N_976);
nand U1060 (N_1060,N_981,N_994);
and U1061 (N_1061,N_1038,N_1025);
nor U1062 (N_1062,N_1009,N_1030);
nand U1063 (N_1063,N_990,N_985);
nand U1064 (N_1064,N_975,N_1018);
nand U1065 (N_1065,N_1034,N_983);
nand U1066 (N_1066,N_977,N_987);
nand U1067 (N_1067,N_1049,N_1033);
and U1068 (N_1068,N_993,N_989);
or U1069 (N_1069,N_1035,N_1045);
or U1070 (N_1070,N_1022,N_1036);
nor U1071 (N_1071,N_999,N_1002);
xor U1072 (N_1072,N_1001,N_1010);
nor U1073 (N_1073,N_1048,N_1044);
or U1074 (N_1074,N_1004,N_984);
nand U1075 (N_1075,N_1007,N_1026);
and U1076 (N_1076,N_1046,N_986);
nor U1077 (N_1077,N_1020,N_978);
and U1078 (N_1078,N_997,N_995);
nor U1079 (N_1079,N_1019,N_1011);
or U1080 (N_1080,N_1037,N_1031);
xnor U1081 (N_1081,N_1016,N_982);
nand U1082 (N_1082,N_1041,N_1032);
xnor U1083 (N_1083,N_1006,N_1042);
xor U1084 (N_1084,N_1029,N_1028);
nor U1085 (N_1085,N_1014,N_980);
xnor U1086 (N_1086,N_1000,N_979);
nor U1087 (N_1087,N_1040,N_1033);
nand U1088 (N_1088,N_1035,N_975);
and U1089 (N_1089,N_975,N_1009);
or U1090 (N_1090,N_1036,N_1000);
and U1091 (N_1091,N_992,N_1006);
nand U1092 (N_1092,N_1001,N_1021);
or U1093 (N_1093,N_1002,N_995);
nand U1094 (N_1094,N_979,N_1025);
and U1095 (N_1095,N_1046,N_1020);
and U1096 (N_1096,N_994,N_1033);
nor U1097 (N_1097,N_983,N_996);
or U1098 (N_1098,N_1034,N_1012);
and U1099 (N_1099,N_1027,N_1046);
and U1100 (N_1100,N_985,N_989);
nor U1101 (N_1101,N_1019,N_1035);
nand U1102 (N_1102,N_1006,N_995);
nor U1103 (N_1103,N_1028,N_1044);
nor U1104 (N_1104,N_985,N_1023);
and U1105 (N_1105,N_984,N_992);
or U1106 (N_1106,N_1039,N_1047);
and U1107 (N_1107,N_1041,N_1029);
nand U1108 (N_1108,N_1005,N_980);
or U1109 (N_1109,N_1008,N_1033);
nor U1110 (N_1110,N_977,N_989);
or U1111 (N_1111,N_1036,N_982);
xnor U1112 (N_1112,N_1014,N_1018);
or U1113 (N_1113,N_1024,N_1048);
or U1114 (N_1114,N_985,N_1037);
xor U1115 (N_1115,N_1007,N_1013);
nor U1116 (N_1116,N_991,N_1005);
or U1117 (N_1117,N_985,N_1009);
or U1118 (N_1118,N_992,N_1028);
or U1119 (N_1119,N_985,N_1043);
nand U1120 (N_1120,N_987,N_1027);
nand U1121 (N_1121,N_995,N_1008);
or U1122 (N_1122,N_993,N_998);
nand U1123 (N_1123,N_985,N_987);
nor U1124 (N_1124,N_1019,N_1022);
and U1125 (N_1125,N_1109,N_1120);
or U1126 (N_1126,N_1070,N_1051);
and U1127 (N_1127,N_1050,N_1122);
nor U1128 (N_1128,N_1092,N_1067);
nand U1129 (N_1129,N_1085,N_1076);
or U1130 (N_1130,N_1112,N_1077);
nor U1131 (N_1131,N_1061,N_1065);
and U1132 (N_1132,N_1091,N_1058);
or U1133 (N_1133,N_1062,N_1093);
nand U1134 (N_1134,N_1059,N_1089);
or U1135 (N_1135,N_1118,N_1094);
and U1136 (N_1136,N_1121,N_1055);
nand U1137 (N_1137,N_1066,N_1119);
and U1138 (N_1138,N_1056,N_1073);
or U1139 (N_1139,N_1105,N_1117);
and U1140 (N_1140,N_1079,N_1064);
nand U1141 (N_1141,N_1114,N_1069);
nor U1142 (N_1142,N_1088,N_1057);
nand U1143 (N_1143,N_1078,N_1095);
and U1144 (N_1144,N_1103,N_1074);
nor U1145 (N_1145,N_1100,N_1111);
or U1146 (N_1146,N_1107,N_1110);
or U1147 (N_1147,N_1099,N_1113);
and U1148 (N_1148,N_1084,N_1072);
xnor U1149 (N_1149,N_1086,N_1075);
nand U1150 (N_1150,N_1082,N_1081);
nand U1151 (N_1151,N_1087,N_1096);
nor U1152 (N_1152,N_1090,N_1063);
xnor U1153 (N_1153,N_1071,N_1054);
nor U1154 (N_1154,N_1108,N_1053);
or U1155 (N_1155,N_1098,N_1123);
nand U1156 (N_1156,N_1097,N_1052);
or U1157 (N_1157,N_1116,N_1083);
or U1158 (N_1158,N_1080,N_1101);
or U1159 (N_1159,N_1068,N_1115);
nor U1160 (N_1160,N_1060,N_1104);
nor U1161 (N_1161,N_1102,N_1106);
nand U1162 (N_1162,N_1124,N_1071);
or U1163 (N_1163,N_1058,N_1094);
and U1164 (N_1164,N_1110,N_1115);
xor U1165 (N_1165,N_1089,N_1102);
nand U1166 (N_1166,N_1061,N_1078);
nor U1167 (N_1167,N_1073,N_1103);
nor U1168 (N_1168,N_1075,N_1095);
nor U1169 (N_1169,N_1075,N_1104);
nand U1170 (N_1170,N_1071,N_1056);
nand U1171 (N_1171,N_1105,N_1087);
nand U1172 (N_1172,N_1056,N_1101);
or U1173 (N_1173,N_1085,N_1073);
and U1174 (N_1174,N_1057,N_1052);
and U1175 (N_1175,N_1109,N_1088);
nand U1176 (N_1176,N_1091,N_1082);
or U1177 (N_1177,N_1094,N_1060);
nor U1178 (N_1178,N_1109,N_1089);
or U1179 (N_1179,N_1050,N_1089);
nand U1180 (N_1180,N_1054,N_1050);
xnor U1181 (N_1181,N_1112,N_1080);
nand U1182 (N_1182,N_1115,N_1052);
and U1183 (N_1183,N_1118,N_1110);
or U1184 (N_1184,N_1060,N_1068);
xor U1185 (N_1185,N_1112,N_1108);
or U1186 (N_1186,N_1050,N_1109);
nand U1187 (N_1187,N_1068,N_1067);
nor U1188 (N_1188,N_1099,N_1064);
or U1189 (N_1189,N_1101,N_1066);
xnor U1190 (N_1190,N_1109,N_1090);
and U1191 (N_1191,N_1122,N_1124);
xnor U1192 (N_1192,N_1100,N_1116);
or U1193 (N_1193,N_1123,N_1054);
and U1194 (N_1194,N_1120,N_1074);
xnor U1195 (N_1195,N_1121,N_1095);
nand U1196 (N_1196,N_1113,N_1106);
or U1197 (N_1197,N_1108,N_1062);
or U1198 (N_1198,N_1069,N_1094);
nor U1199 (N_1199,N_1115,N_1095);
and U1200 (N_1200,N_1148,N_1131);
nor U1201 (N_1201,N_1195,N_1159);
xnor U1202 (N_1202,N_1156,N_1142);
or U1203 (N_1203,N_1145,N_1171);
nor U1204 (N_1204,N_1198,N_1187);
nand U1205 (N_1205,N_1193,N_1160);
and U1206 (N_1206,N_1194,N_1162);
or U1207 (N_1207,N_1140,N_1177);
nand U1208 (N_1208,N_1188,N_1185);
nand U1209 (N_1209,N_1146,N_1172);
or U1210 (N_1210,N_1143,N_1168);
nand U1211 (N_1211,N_1190,N_1178);
nand U1212 (N_1212,N_1191,N_1134);
nand U1213 (N_1213,N_1184,N_1157);
nand U1214 (N_1214,N_1136,N_1127);
and U1215 (N_1215,N_1129,N_1132);
or U1216 (N_1216,N_1135,N_1183);
and U1217 (N_1217,N_1169,N_1147);
and U1218 (N_1218,N_1176,N_1197);
nand U1219 (N_1219,N_1149,N_1181);
and U1220 (N_1220,N_1189,N_1166);
and U1221 (N_1221,N_1126,N_1161);
and U1222 (N_1222,N_1128,N_1180);
nor U1223 (N_1223,N_1155,N_1174);
nand U1224 (N_1224,N_1165,N_1125);
and U1225 (N_1225,N_1150,N_1179);
or U1226 (N_1226,N_1175,N_1152);
or U1227 (N_1227,N_1186,N_1167);
nand U1228 (N_1228,N_1138,N_1139);
and U1229 (N_1229,N_1170,N_1173);
nor U1230 (N_1230,N_1163,N_1158);
or U1231 (N_1231,N_1182,N_1154);
xnor U1232 (N_1232,N_1141,N_1199);
or U1233 (N_1233,N_1192,N_1151);
nand U1234 (N_1234,N_1133,N_1130);
nor U1235 (N_1235,N_1144,N_1153);
and U1236 (N_1236,N_1164,N_1196);
and U1237 (N_1237,N_1137,N_1179);
or U1238 (N_1238,N_1142,N_1189);
or U1239 (N_1239,N_1169,N_1166);
and U1240 (N_1240,N_1180,N_1181);
or U1241 (N_1241,N_1151,N_1148);
or U1242 (N_1242,N_1192,N_1141);
nor U1243 (N_1243,N_1198,N_1160);
and U1244 (N_1244,N_1191,N_1132);
nor U1245 (N_1245,N_1185,N_1193);
or U1246 (N_1246,N_1126,N_1160);
or U1247 (N_1247,N_1173,N_1133);
nor U1248 (N_1248,N_1171,N_1148);
or U1249 (N_1249,N_1178,N_1176);
or U1250 (N_1250,N_1171,N_1187);
or U1251 (N_1251,N_1152,N_1173);
nor U1252 (N_1252,N_1125,N_1127);
or U1253 (N_1253,N_1174,N_1156);
or U1254 (N_1254,N_1158,N_1184);
and U1255 (N_1255,N_1141,N_1193);
xor U1256 (N_1256,N_1199,N_1140);
nand U1257 (N_1257,N_1197,N_1137);
and U1258 (N_1258,N_1157,N_1194);
or U1259 (N_1259,N_1128,N_1157);
nand U1260 (N_1260,N_1182,N_1141);
nand U1261 (N_1261,N_1127,N_1197);
and U1262 (N_1262,N_1177,N_1178);
nor U1263 (N_1263,N_1142,N_1195);
nand U1264 (N_1264,N_1136,N_1129);
and U1265 (N_1265,N_1148,N_1167);
and U1266 (N_1266,N_1135,N_1130);
nor U1267 (N_1267,N_1151,N_1185);
and U1268 (N_1268,N_1194,N_1166);
nor U1269 (N_1269,N_1139,N_1135);
nand U1270 (N_1270,N_1150,N_1189);
nor U1271 (N_1271,N_1131,N_1147);
or U1272 (N_1272,N_1128,N_1199);
nand U1273 (N_1273,N_1146,N_1165);
and U1274 (N_1274,N_1153,N_1187);
nand U1275 (N_1275,N_1270,N_1210);
nand U1276 (N_1276,N_1215,N_1265);
or U1277 (N_1277,N_1220,N_1228);
or U1278 (N_1278,N_1233,N_1203);
and U1279 (N_1279,N_1227,N_1222);
and U1280 (N_1280,N_1245,N_1264);
and U1281 (N_1281,N_1256,N_1209);
nor U1282 (N_1282,N_1202,N_1218);
or U1283 (N_1283,N_1206,N_1208);
nand U1284 (N_1284,N_1235,N_1205);
and U1285 (N_1285,N_1259,N_1242);
nor U1286 (N_1286,N_1261,N_1244);
nand U1287 (N_1287,N_1201,N_1274);
or U1288 (N_1288,N_1239,N_1234);
or U1289 (N_1289,N_1250,N_1240);
nor U1290 (N_1290,N_1266,N_1272);
or U1291 (N_1291,N_1238,N_1251);
nand U1292 (N_1292,N_1212,N_1211);
and U1293 (N_1293,N_1207,N_1258);
nor U1294 (N_1294,N_1226,N_1260);
and U1295 (N_1295,N_1236,N_1204);
nand U1296 (N_1296,N_1217,N_1213);
nand U1297 (N_1297,N_1243,N_1248);
or U1298 (N_1298,N_1267,N_1219);
or U1299 (N_1299,N_1221,N_1225);
nand U1300 (N_1300,N_1214,N_1252);
nor U1301 (N_1301,N_1223,N_1247);
nand U1302 (N_1302,N_1232,N_1268);
and U1303 (N_1303,N_1246,N_1263);
or U1304 (N_1304,N_1254,N_1231);
and U1305 (N_1305,N_1216,N_1237);
and U1306 (N_1306,N_1229,N_1269);
and U1307 (N_1307,N_1200,N_1241);
nand U1308 (N_1308,N_1253,N_1257);
nand U1309 (N_1309,N_1249,N_1224);
and U1310 (N_1310,N_1262,N_1271);
or U1311 (N_1311,N_1255,N_1230);
xor U1312 (N_1312,N_1273,N_1221);
nor U1313 (N_1313,N_1226,N_1232);
and U1314 (N_1314,N_1224,N_1250);
or U1315 (N_1315,N_1208,N_1259);
xnor U1316 (N_1316,N_1260,N_1272);
or U1317 (N_1317,N_1257,N_1217);
nand U1318 (N_1318,N_1228,N_1230);
nand U1319 (N_1319,N_1223,N_1239);
xor U1320 (N_1320,N_1214,N_1218);
nand U1321 (N_1321,N_1263,N_1271);
and U1322 (N_1322,N_1205,N_1237);
or U1323 (N_1323,N_1244,N_1246);
and U1324 (N_1324,N_1254,N_1217);
or U1325 (N_1325,N_1239,N_1266);
nor U1326 (N_1326,N_1264,N_1218);
nand U1327 (N_1327,N_1228,N_1265);
nor U1328 (N_1328,N_1234,N_1220);
nor U1329 (N_1329,N_1262,N_1221);
nor U1330 (N_1330,N_1262,N_1243);
nor U1331 (N_1331,N_1200,N_1239);
and U1332 (N_1332,N_1268,N_1225);
xnor U1333 (N_1333,N_1244,N_1227);
nor U1334 (N_1334,N_1250,N_1201);
xor U1335 (N_1335,N_1245,N_1221);
and U1336 (N_1336,N_1204,N_1220);
and U1337 (N_1337,N_1253,N_1227);
and U1338 (N_1338,N_1235,N_1230);
nand U1339 (N_1339,N_1242,N_1215);
nor U1340 (N_1340,N_1256,N_1262);
or U1341 (N_1341,N_1263,N_1233);
nor U1342 (N_1342,N_1202,N_1247);
or U1343 (N_1343,N_1210,N_1265);
and U1344 (N_1344,N_1272,N_1257);
and U1345 (N_1345,N_1259,N_1238);
or U1346 (N_1346,N_1268,N_1257);
nand U1347 (N_1347,N_1262,N_1211);
and U1348 (N_1348,N_1257,N_1258);
nor U1349 (N_1349,N_1233,N_1231);
and U1350 (N_1350,N_1277,N_1309);
xnor U1351 (N_1351,N_1341,N_1283);
or U1352 (N_1352,N_1295,N_1275);
or U1353 (N_1353,N_1328,N_1312);
nor U1354 (N_1354,N_1299,N_1332);
or U1355 (N_1355,N_1282,N_1335);
or U1356 (N_1356,N_1294,N_1322);
and U1357 (N_1357,N_1305,N_1276);
or U1358 (N_1358,N_1344,N_1280);
or U1359 (N_1359,N_1318,N_1301);
nand U1360 (N_1360,N_1348,N_1325);
or U1361 (N_1361,N_1324,N_1346);
nand U1362 (N_1362,N_1284,N_1279);
nor U1363 (N_1363,N_1329,N_1298);
and U1364 (N_1364,N_1339,N_1278);
and U1365 (N_1365,N_1291,N_1314);
nand U1366 (N_1366,N_1297,N_1311);
or U1367 (N_1367,N_1327,N_1323);
or U1368 (N_1368,N_1289,N_1345);
and U1369 (N_1369,N_1286,N_1287);
xnor U1370 (N_1370,N_1296,N_1338);
nor U1371 (N_1371,N_1293,N_1308);
nor U1372 (N_1372,N_1288,N_1336);
nand U1373 (N_1373,N_1310,N_1321);
xor U1374 (N_1374,N_1333,N_1330);
nand U1375 (N_1375,N_1320,N_1315);
and U1376 (N_1376,N_1340,N_1292);
xnor U1377 (N_1377,N_1304,N_1281);
or U1378 (N_1378,N_1349,N_1307);
xor U1379 (N_1379,N_1337,N_1290);
nor U1380 (N_1380,N_1347,N_1317);
and U1381 (N_1381,N_1303,N_1313);
and U1382 (N_1382,N_1334,N_1342);
nand U1383 (N_1383,N_1302,N_1300);
and U1384 (N_1384,N_1343,N_1319);
nor U1385 (N_1385,N_1316,N_1326);
nor U1386 (N_1386,N_1306,N_1285);
and U1387 (N_1387,N_1331,N_1335);
and U1388 (N_1388,N_1316,N_1322);
or U1389 (N_1389,N_1347,N_1287);
or U1390 (N_1390,N_1305,N_1318);
nor U1391 (N_1391,N_1324,N_1318);
nor U1392 (N_1392,N_1310,N_1302);
nand U1393 (N_1393,N_1328,N_1338);
nand U1394 (N_1394,N_1279,N_1291);
and U1395 (N_1395,N_1313,N_1292);
and U1396 (N_1396,N_1304,N_1332);
nand U1397 (N_1397,N_1276,N_1299);
nand U1398 (N_1398,N_1309,N_1326);
nor U1399 (N_1399,N_1334,N_1325);
and U1400 (N_1400,N_1296,N_1294);
nor U1401 (N_1401,N_1319,N_1302);
and U1402 (N_1402,N_1300,N_1335);
xnor U1403 (N_1403,N_1315,N_1331);
nand U1404 (N_1404,N_1346,N_1287);
and U1405 (N_1405,N_1331,N_1329);
xor U1406 (N_1406,N_1347,N_1299);
xor U1407 (N_1407,N_1340,N_1286);
nor U1408 (N_1408,N_1288,N_1287);
and U1409 (N_1409,N_1305,N_1345);
xnor U1410 (N_1410,N_1286,N_1320);
and U1411 (N_1411,N_1279,N_1299);
nand U1412 (N_1412,N_1310,N_1299);
or U1413 (N_1413,N_1295,N_1346);
nor U1414 (N_1414,N_1302,N_1328);
nand U1415 (N_1415,N_1302,N_1299);
nor U1416 (N_1416,N_1301,N_1286);
and U1417 (N_1417,N_1295,N_1313);
or U1418 (N_1418,N_1277,N_1336);
nand U1419 (N_1419,N_1337,N_1294);
and U1420 (N_1420,N_1291,N_1339);
or U1421 (N_1421,N_1298,N_1293);
xor U1422 (N_1422,N_1341,N_1329);
and U1423 (N_1423,N_1288,N_1277);
and U1424 (N_1424,N_1276,N_1291);
and U1425 (N_1425,N_1376,N_1410);
nand U1426 (N_1426,N_1364,N_1391);
nor U1427 (N_1427,N_1396,N_1408);
nor U1428 (N_1428,N_1394,N_1407);
xor U1429 (N_1429,N_1399,N_1405);
and U1430 (N_1430,N_1397,N_1412);
or U1431 (N_1431,N_1402,N_1352);
nor U1432 (N_1432,N_1395,N_1423);
or U1433 (N_1433,N_1374,N_1388);
nor U1434 (N_1434,N_1356,N_1418);
nor U1435 (N_1435,N_1368,N_1379);
nand U1436 (N_1436,N_1361,N_1350);
nor U1437 (N_1437,N_1367,N_1351);
nor U1438 (N_1438,N_1387,N_1369);
and U1439 (N_1439,N_1421,N_1354);
or U1440 (N_1440,N_1363,N_1413);
xor U1441 (N_1441,N_1393,N_1381);
nor U1442 (N_1442,N_1416,N_1372);
and U1443 (N_1443,N_1414,N_1392);
nor U1444 (N_1444,N_1406,N_1404);
or U1445 (N_1445,N_1358,N_1362);
and U1446 (N_1446,N_1409,N_1357);
and U1447 (N_1447,N_1415,N_1389);
or U1448 (N_1448,N_1353,N_1373);
or U1449 (N_1449,N_1390,N_1417);
nand U1450 (N_1450,N_1386,N_1384);
and U1451 (N_1451,N_1411,N_1382);
and U1452 (N_1452,N_1385,N_1378);
and U1453 (N_1453,N_1424,N_1377);
xor U1454 (N_1454,N_1398,N_1383);
xnor U1455 (N_1455,N_1359,N_1401);
nor U1456 (N_1456,N_1366,N_1375);
nor U1457 (N_1457,N_1360,N_1355);
and U1458 (N_1458,N_1419,N_1400);
and U1459 (N_1459,N_1380,N_1370);
or U1460 (N_1460,N_1371,N_1420);
or U1461 (N_1461,N_1422,N_1403);
nand U1462 (N_1462,N_1365,N_1367);
and U1463 (N_1463,N_1399,N_1392);
or U1464 (N_1464,N_1358,N_1417);
and U1465 (N_1465,N_1395,N_1402);
and U1466 (N_1466,N_1406,N_1351);
nor U1467 (N_1467,N_1351,N_1424);
nand U1468 (N_1468,N_1420,N_1359);
and U1469 (N_1469,N_1367,N_1353);
or U1470 (N_1470,N_1382,N_1364);
or U1471 (N_1471,N_1419,N_1402);
or U1472 (N_1472,N_1368,N_1393);
nor U1473 (N_1473,N_1352,N_1413);
and U1474 (N_1474,N_1367,N_1414);
and U1475 (N_1475,N_1354,N_1378);
nand U1476 (N_1476,N_1414,N_1408);
or U1477 (N_1477,N_1372,N_1373);
nor U1478 (N_1478,N_1387,N_1374);
xnor U1479 (N_1479,N_1419,N_1417);
nor U1480 (N_1480,N_1351,N_1365);
and U1481 (N_1481,N_1359,N_1399);
and U1482 (N_1482,N_1393,N_1367);
nor U1483 (N_1483,N_1403,N_1381);
nand U1484 (N_1484,N_1377,N_1396);
and U1485 (N_1485,N_1373,N_1393);
nor U1486 (N_1486,N_1354,N_1398);
and U1487 (N_1487,N_1388,N_1371);
xnor U1488 (N_1488,N_1360,N_1413);
xnor U1489 (N_1489,N_1408,N_1387);
nand U1490 (N_1490,N_1357,N_1362);
and U1491 (N_1491,N_1403,N_1374);
nand U1492 (N_1492,N_1372,N_1375);
xor U1493 (N_1493,N_1422,N_1413);
and U1494 (N_1494,N_1382,N_1359);
nor U1495 (N_1495,N_1359,N_1405);
nor U1496 (N_1496,N_1410,N_1408);
xnor U1497 (N_1497,N_1362,N_1367);
nor U1498 (N_1498,N_1365,N_1371);
and U1499 (N_1499,N_1360,N_1378);
or U1500 (N_1500,N_1471,N_1478);
nand U1501 (N_1501,N_1441,N_1444);
and U1502 (N_1502,N_1480,N_1461);
or U1503 (N_1503,N_1470,N_1465);
xnor U1504 (N_1504,N_1492,N_1493);
xor U1505 (N_1505,N_1433,N_1435);
nand U1506 (N_1506,N_1484,N_1449);
and U1507 (N_1507,N_1432,N_1467);
and U1508 (N_1508,N_1482,N_1483);
nor U1509 (N_1509,N_1456,N_1489);
or U1510 (N_1510,N_1469,N_1496);
and U1511 (N_1511,N_1464,N_1430);
and U1512 (N_1512,N_1450,N_1499);
nor U1513 (N_1513,N_1447,N_1457);
and U1514 (N_1514,N_1440,N_1498);
nor U1515 (N_1515,N_1437,N_1425);
or U1516 (N_1516,N_1431,N_1486);
nor U1517 (N_1517,N_1477,N_1442);
and U1518 (N_1518,N_1448,N_1446);
and U1519 (N_1519,N_1439,N_1445);
nand U1520 (N_1520,N_1459,N_1474);
nand U1521 (N_1521,N_1479,N_1475);
or U1522 (N_1522,N_1451,N_1491);
and U1523 (N_1523,N_1494,N_1460);
nand U1524 (N_1524,N_1453,N_1490);
nor U1525 (N_1525,N_1438,N_1427);
and U1526 (N_1526,N_1426,N_1476);
and U1527 (N_1527,N_1454,N_1472);
nor U1528 (N_1528,N_1458,N_1488);
nor U1529 (N_1529,N_1463,N_1468);
xor U1530 (N_1530,N_1436,N_1452);
or U1531 (N_1531,N_1434,N_1455);
or U1532 (N_1532,N_1466,N_1473);
nor U1533 (N_1533,N_1462,N_1487);
nand U1534 (N_1534,N_1429,N_1481);
or U1535 (N_1535,N_1495,N_1497);
and U1536 (N_1536,N_1485,N_1443);
or U1537 (N_1537,N_1428,N_1440);
or U1538 (N_1538,N_1475,N_1456);
or U1539 (N_1539,N_1478,N_1499);
and U1540 (N_1540,N_1448,N_1480);
nand U1541 (N_1541,N_1473,N_1452);
and U1542 (N_1542,N_1477,N_1447);
and U1543 (N_1543,N_1437,N_1435);
or U1544 (N_1544,N_1488,N_1453);
nand U1545 (N_1545,N_1499,N_1445);
and U1546 (N_1546,N_1486,N_1430);
and U1547 (N_1547,N_1491,N_1473);
nor U1548 (N_1548,N_1439,N_1462);
or U1549 (N_1549,N_1434,N_1482);
and U1550 (N_1550,N_1437,N_1444);
and U1551 (N_1551,N_1455,N_1431);
or U1552 (N_1552,N_1435,N_1499);
nor U1553 (N_1553,N_1485,N_1426);
nand U1554 (N_1554,N_1494,N_1450);
nand U1555 (N_1555,N_1458,N_1477);
or U1556 (N_1556,N_1486,N_1472);
and U1557 (N_1557,N_1486,N_1497);
and U1558 (N_1558,N_1453,N_1427);
nand U1559 (N_1559,N_1482,N_1444);
xor U1560 (N_1560,N_1458,N_1444);
or U1561 (N_1561,N_1480,N_1430);
and U1562 (N_1562,N_1476,N_1468);
or U1563 (N_1563,N_1479,N_1466);
and U1564 (N_1564,N_1468,N_1450);
nand U1565 (N_1565,N_1485,N_1448);
nor U1566 (N_1566,N_1469,N_1494);
and U1567 (N_1567,N_1486,N_1492);
nor U1568 (N_1568,N_1489,N_1491);
nand U1569 (N_1569,N_1486,N_1477);
nor U1570 (N_1570,N_1460,N_1447);
nand U1571 (N_1571,N_1433,N_1489);
and U1572 (N_1572,N_1467,N_1452);
or U1573 (N_1573,N_1440,N_1481);
nand U1574 (N_1574,N_1454,N_1466);
or U1575 (N_1575,N_1511,N_1547);
and U1576 (N_1576,N_1522,N_1510);
or U1577 (N_1577,N_1562,N_1544);
and U1578 (N_1578,N_1503,N_1502);
nand U1579 (N_1579,N_1541,N_1500);
and U1580 (N_1580,N_1513,N_1564);
nand U1581 (N_1581,N_1516,N_1507);
xnor U1582 (N_1582,N_1529,N_1561);
and U1583 (N_1583,N_1543,N_1537);
or U1584 (N_1584,N_1518,N_1534);
nand U1585 (N_1585,N_1554,N_1538);
nand U1586 (N_1586,N_1521,N_1540);
nand U1587 (N_1587,N_1501,N_1536);
or U1588 (N_1588,N_1553,N_1509);
nand U1589 (N_1589,N_1569,N_1528);
nor U1590 (N_1590,N_1556,N_1568);
nand U1591 (N_1591,N_1505,N_1560);
or U1592 (N_1592,N_1546,N_1526);
and U1593 (N_1593,N_1525,N_1552);
and U1594 (N_1594,N_1550,N_1548);
nor U1595 (N_1595,N_1520,N_1527);
nand U1596 (N_1596,N_1542,N_1559);
and U1597 (N_1597,N_1557,N_1514);
nand U1598 (N_1598,N_1519,N_1532);
nand U1599 (N_1599,N_1555,N_1572);
nand U1600 (N_1600,N_1531,N_1549);
nor U1601 (N_1601,N_1515,N_1574);
nand U1602 (N_1602,N_1566,N_1506);
xor U1603 (N_1603,N_1570,N_1533);
nor U1604 (N_1604,N_1573,N_1517);
nand U1605 (N_1605,N_1535,N_1523);
or U1606 (N_1606,N_1565,N_1512);
nor U1607 (N_1607,N_1571,N_1530);
or U1608 (N_1608,N_1524,N_1563);
nor U1609 (N_1609,N_1508,N_1551);
nor U1610 (N_1610,N_1558,N_1539);
and U1611 (N_1611,N_1545,N_1504);
nor U1612 (N_1612,N_1567,N_1557);
or U1613 (N_1613,N_1570,N_1514);
or U1614 (N_1614,N_1545,N_1571);
nor U1615 (N_1615,N_1541,N_1545);
and U1616 (N_1616,N_1507,N_1523);
and U1617 (N_1617,N_1547,N_1538);
and U1618 (N_1618,N_1513,N_1551);
or U1619 (N_1619,N_1507,N_1529);
xor U1620 (N_1620,N_1521,N_1500);
or U1621 (N_1621,N_1546,N_1549);
nor U1622 (N_1622,N_1505,N_1541);
nor U1623 (N_1623,N_1523,N_1529);
nor U1624 (N_1624,N_1527,N_1526);
or U1625 (N_1625,N_1532,N_1554);
nand U1626 (N_1626,N_1536,N_1561);
nand U1627 (N_1627,N_1530,N_1561);
and U1628 (N_1628,N_1500,N_1556);
nor U1629 (N_1629,N_1557,N_1513);
or U1630 (N_1630,N_1550,N_1532);
and U1631 (N_1631,N_1535,N_1567);
and U1632 (N_1632,N_1542,N_1511);
or U1633 (N_1633,N_1561,N_1528);
and U1634 (N_1634,N_1530,N_1542);
nor U1635 (N_1635,N_1542,N_1539);
and U1636 (N_1636,N_1548,N_1551);
nor U1637 (N_1637,N_1528,N_1542);
nand U1638 (N_1638,N_1537,N_1514);
and U1639 (N_1639,N_1555,N_1525);
and U1640 (N_1640,N_1513,N_1523);
nor U1641 (N_1641,N_1504,N_1532);
and U1642 (N_1642,N_1558,N_1533);
or U1643 (N_1643,N_1541,N_1526);
nor U1644 (N_1644,N_1512,N_1566);
nand U1645 (N_1645,N_1515,N_1521);
xor U1646 (N_1646,N_1532,N_1548);
nor U1647 (N_1647,N_1561,N_1522);
nor U1648 (N_1648,N_1546,N_1522);
and U1649 (N_1649,N_1564,N_1565);
nor U1650 (N_1650,N_1638,N_1635);
nand U1651 (N_1651,N_1582,N_1623);
nor U1652 (N_1652,N_1606,N_1631);
and U1653 (N_1653,N_1637,N_1603);
and U1654 (N_1654,N_1611,N_1575);
nor U1655 (N_1655,N_1642,N_1579);
nor U1656 (N_1656,N_1593,N_1595);
or U1657 (N_1657,N_1604,N_1605);
and U1658 (N_1658,N_1597,N_1587);
and U1659 (N_1659,N_1577,N_1609);
nand U1660 (N_1660,N_1594,N_1646);
and U1661 (N_1661,N_1612,N_1602);
nor U1662 (N_1662,N_1592,N_1578);
nor U1663 (N_1663,N_1617,N_1636);
nand U1664 (N_1664,N_1616,N_1640);
nor U1665 (N_1665,N_1645,N_1580);
and U1666 (N_1666,N_1647,N_1625);
and U1667 (N_1667,N_1589,N_1614);
nand U1668 (N_1668,N_1586,N_1581);
and U1669 (N_1669,N_1622,N_1641);
nor U1670 (N_1670,N_1633,N_1607);
nand U1671 (N_1671,N_1600,N_1649);
or U1672 (N_1672,N_1624,N_1599);
xnor U1673 (N_1673,N_1615,N_1590);
nand U1674 (N_1674,N_1632,N_1584);
nand U1675 (N_1675,N_1585,N_1619);
and U1676 (N_1676,N_1644,N_1627);
nand U1677 (N_1677,N_1608,N_1601);
or U1678 (N_1678,N_1643,N_1576);
and U1679 (N_1679,N_1596,N_1588);
nor U1680 (N_1680,N_1630,N_1613);
nand U1681 (N_1681,N_1629,N_1626);
nand U1682 (N_1682,N_1618,N_1639);
nor U1683 (N_1683,N_1620,N_1591);
and U1684 (N_1684,N_1583,N_1610);
and U1685 (N_1685,N_1598,N_1621);
nand U1686 (N_1686,N_1634,N_1648);
xor U1687 (N_1687,N_1628,N_1606);
nor U1688 (N_1688,N_1585,N_1609);
xnor U1689 (N_1689,N_1609,N_1593);
nor U1690 (N_1690,N_1638,N_1640);
and U1691 (N_1691,N_1588,N_1627);
and U1692 (N_1692,N_1629,N_1634);
nand U1693 (N_1693,N_1642,N_1633);
nor U1694 (N_1694,N_1646,N_1622);
and U1695 (N_1695,N_1582,N_1587);
and U1696 (N_1696,N_1609,N_1626);
and U1697 (N_1697,N_1645,N_1583);
or U1698 (N_1698,N_1582,N_1586);
nor U1699 (N_1699,N_1608,N_1589);
xnor U1700 (N_1700,N_1621,N_1624);
nor U1701 (N_1701,N_1605,N_1592);
nand U1702 (N_1702,N_1622,N_1616);
nor U1703 (N_1703,N_1617,N_1648);
and U1704 (N_1704,N_1614,N_1579);
nand U1705 (N_1705,N_1590,N_1575);
xnor U1706 (N_1706,N_1598,N_1629);
xor U1707 (N_1707,N_1630,N_1611);
or U1708 (N_1708,N_1644,N_1615);
nor U1709 (N_1709,N_1613,N_1593);
nand U1710 (N_1710,N_1588,N_1603);
nand U1711 (N_1711,N_1619,N_1623);
and U1712 (N_1712,N_1631,N_1576);
nand U1713 (N_1713,N_1584,N_1596);
nor U1714 (N_1714,N_1576,N_1584);
or U1715 (N_1715,N_1605,N_1581);
nor U1716 (N_1716,N_1645,N_1579);
and U1717 (N_1717,N_1616,N_1620);
nand U1718 (N_1718,N_1619,N_1584);
and U1719 (N_1719,N_1637,N_1596);
and U1720 (N_1720,N_1639,N_1617);
nor U1721 (N_1721,N_1599,N_1620);
xnor U1722 (N_1722,N_1585,N_1633);
and U1723 (N_1723,N_1648,N_1591);
and U1724 (N_1724,N_1610,N_1636);
nor U1725 (N_1725,N_1668,N_1675);
and U1726 (N_1726,N_1687,N_1700);
nor U1727 (N_1727,N_1704,N_1692);
and U1728 (N_1728,N_1667,N_1683);
nor U1729 (N_1729,N_1682,N_1661);
xor U1730 (N_1730,N_1664,N_1694);
nor U1731 (N_1731,N_1669,N_1660);
nand U1732 (N_1732,N_1715,N_1685);
or U1733 (N_1733,N_1653,N_1714);
nand U1734 (N_1734,N_1674,N_1693);
nor U1735 (N_1735,N_1701,N_1721);
and U1736 (N_1736,N_1705,N_1658);
and U1737 (N_1737,N_1720,N_1695);
nor U1738 (N_1738,N_1670,N_1699);
or U1739 (N_1739,N_1652,N_1698);
nand U1740 (N_1740,N_1672,N_1688);
nor U1741 (N_1741,N_1723,N_1696);
and U1742 (N_1742,N_1656,N_1666);
nor U1743 (N_1743,N_1678,N_1718);
and U1744 (N_1744,N_1719,N_1717);
or U1745 (N_1745,N_1722,N_1679);
or U1746 (N_1746,N_1702,N_1716);
nand U1747 (N_1747,N_1663,N_1680);
nor U1748 (N_1748,N_1654,N_1651);
and U1749 (N_1749,N_1684,N_1662);
and U1750 (N_1750,N_1676,N_1657);
nand U1751 (N_1751,N_1713,N_1703);
nand U1752 (N_1752,N_1707,N_1665);
nor U1753 (N_1753,N_1673,N_1690);
nor U1754 (N_1754,N_1709,N_1708);
nor U1755 (N_1755,N_1671,N_1689);
or U1756 (N_1756,N_1697,N_1691);
and U1757 (N_1757,N_1659,N_1712);
or U1758 (N_1758,N_1724,N_1677);
nor U1759 (N_1759,N_1650,N_1686);
and U1760 (N_1760,N_1711,N_1655);
and U1761 (N_1761,N_1681,N_1706);
or U1762 (N_1762,N_1710,N_1692);
or U1763 (N_1763,N_1691,N_1678);
nand U1764 (N_1764,N_1700,N_1657);
nand U1765 (N_1765,N_1721,N_1690);
nor U1766 (N_1766,N_1721,N_1719);
nand U1767 (N_1767,N_1686,N_1688);
nor U1768 (N_1768,N_1692,N_1680);
nor U1769 (N_1769,N_1682,N_1681);
nand U1770 (N_1770,N_1659,N_1721);
and U1771 (N_1771,N_1710,N_1720);
and U1772 (N_1772,N_1694,N_1707);
nor U1773 (N_1773,N_1694,N_1658);
or U1774 (N_1774,N_1655,N_1707);
and U1775 (N_1775,N_1694,N_1650);
nand U1776 (N_1776,N_1663,N_1691);
nand U1777 (N_1777,N_1681,N_1667);
nand U1778 (N_1778,N_1682,N_1708);
nand U1779 (N_1779,N_1684,N_1687);
or U1780 (N_1780,N_1697,N_1690);
nand U1781 (N_1781,N_1699,N_1654);
nand U1782 (N_1782,N_1710,N_1664);
or U1783 (N_1783,N_1691,N_1690);
nand U1784 (N_1784,N_1652,N_1715);
nor U1785 (N_1785,N_1705,N_1706);
nand U1786 (N_1786,N_1717,N_1724);
nor U1787 (N_1787,N_1666,N_1673);
or U1788 (N_1788,N_1671,N_1723);
or U1789 (N_1789,N_1718,N_1713);
nand U1790 (N_1790,N_1656,N_1673);
nand U1791 (N_1791,N_1677,N_1703);
nor U1792 (N_1792,N_1709,N_1711);
nand U1793 (N_1793,N_1699,N_1661);
xnor U1794 (N_1794,N_1656,N_1689);
and U1795 (N_1795,N_1661,N_1701);
and U1796 (N_1796,N_1701,N_1666);
or U1797 (N_1797,N_1675,N_1678);
and U1798 (N_1798,N_1679,N_1672);
and U1799 (N_1799,N_1662,N_1707);
nand U1800 (N_1800,N_1733,N_1756);
nor U1801 (N_1801,N_1797,N_1774);
or U1802 (N_1802,N_1732,N_1785);
xor U1803 (N_1803,N_1752,N_1735);
and U1804 (N_1804,N_1795,N_1736);
nor U1805 (N_1805,N_1761,N_1777);
xor U1806 (N_1806,N_1757,N_1737);
nand U1807 (N_1807,N_1744,N_1741);
nor U1808 (N_1808,N_1755,N_1768);
nor U1809 (N_1809,N_1762,N_1759);
nand U1810 (N_1810,N_1798,N_1794);
nor U1811 (N_1811,N_1753,N_1725);
nand U1812 (N_1812,N_1751,N_1784);
xnor U1813 (N_1813,N_1779,N_1734);
and U1814 (N_1814,N_1739,N_1788);
or U1815 (N_1815,N_1748,N_1745);
or U1816 (N_1816,N_1787,N_1749);
and U1817 (N_1817,N_1758,N_1780);
or U1818 (N_1818,N_1767,N_1783);
nand U1819 (N_1819,N_1727,N_1782);
or U1820 (N_1820,N_1799,N_1731);
nor U1821 (N_1821,N_1791,N_1729);
nor U1822 (N_1822,N_1771,N_1746);
and U1823 (N_1823,N_1792,N_1743);
or U1824 (N_1824,N_1781,N_1760);
or U1825 (N_1825,N_1772,N_1793);
and U1826 (N_1826,N_1766,N_1754);
xor U1827 (N_1827,N_1728,N_1770);
nand U1828 (N_1828,N_1764,N_1765);
or U1829 (N_1829,N_1773,N_1796);
or U1830 (N_1830,N_1726,N_1769);
and U1831 (N_1831,N_1778,N_1786);
nor U1832 (N_1832,N_1750,N_1789);
and U1833 (N_1833,N_1742,N_1747);
xor U1834 (N_1834,N_1730,N_1775);
nor U1835 (N_1835,N_1776,N_1740);
and U1836 (N_1836,N_1738,N_1763);
and U1837 (N_1837,N_1790,N_1760);
nand U1838 (N_1838,N_1793,N_1748);
nor U1839 (N_1839,N_1798,N_1756);
or U1840 (N_1840,N_1796,N_1790);
or U1841 (N_1841,N_1792,N_1756);
nor U1842 (N_1842,N_1746,N_1792);
nand U1843 (N_1843,N_1742,N_1754);
and U1844 (N_1844,N_1748,N_1788);
and U1845 (N_1845,N_1760,N_1743);
nor U1846 (N_1846,N_1745,N_1789);
and U1847 (N_1847,N_1760,N_1746);
or U1848 (N_1848,N_1771,N_1797);
or U1849 (N_1849,N_1794,N_1770);
nor U1850 (N_1850,N_1740,N_1796);
nor U1851 (N_1851,N_1757,N_1792);
or U1852 (N_1852,N_1750,N_1757);
nor U1853 (N_1853,N_1788,N_1780);
nand U1854 (N_1854,N_1730,N_1759);
nor U1855 (N_1855,N_1735,N_1798);
or U1856 (N_1856,N_1750,N_1756);
nand U1857 (N_1857,N_1786,N_1744);
xnor U1858 (N_1858,N_1729,N_1762);
and U1859 (N_1859,N_1780,N_1797);
or U1860 (N_1860,N_1755,N_1756);
nand U1861 (N_1861,N_1766,N_1794);
or U1862 (N_1862,N_1730,N_1782);
or U1863 (N_1863,N_1741,N_1778);
and U1864 (N_1864,N_1774,N_1725);
nor U1865 (N_1865,N_1788,N_1781);
or U1866 (N_1866,N_1798,N_1777);
and U1867 (N_1867,N_1747,N_1728);
nor U1868 (N_1868,N_1746,N_1730);
nor U1869 (N_1869,N_1760,N_1729);
nand U1870 (N_1870,N_1747,N_1756);
nand U1871 (N_1871,N_1725,N_1758);
nand U1872 (N_1872,N_1773,N_1745);
nor U1873 (N_1873,N_1786,N_1740);
and U1874 (N_1874,N_1753,N_1793);
nand U1875 (N_1875,N_1807,N_1870);
or U1876 (N_1876,N_1828,N_1822);
nor U1877 (N_1877,N_1842,N_1848);
nand U1878 (N_1878,N_1839,N_1840);
nor U1879 (N_1879,N_1804,N_1872);
and U1880 (N_1880,N_1835,N_1868);
or U1881 (N_1881,N_1865,N_1847);
or U1882 (N_1882,N_1864,N_1866);
nand U1883 (N_1883,N_1831,N_1819);
or U1884 (N_1884,N_1873,N_1829);
or U1885 (N_1885,N_1874,N_1860);
nor U1886 (N_1886,N_1867,N_1817);
nor U1887 (N_1887,N_1802,N_1811);
nand U1888 (N_1888,N_1833,N_1845);
or U1889 (N_1889,N_1856,N_1869);
nor U1890 (N_1890,N_1812,N_1832);
and U1891 (N_1891,N_1814,N_1836);
and U1892 (N_1892,N_1827,N_1858);
nand U1893 (N_1893,N_1846,N_1859);
nor U1894 (N_1894,N_1809,N_1871);
or U1895 (N_1895,N_1826,N_1806);
nand U1896 (N_1896,N_1861,N_1815);
nor U1897 (N_1897,N_1821,N_1830);
or U1898 (N_1898,N_1844,N_1803);
nor U1899 (N_1899,N_1862,N_1805);
nand U1900 (N_1900,N_1853,N_1834);
nand U1901 (N_1901,N_1863,N_1838);
nand U1902 (N_1902,N_1810,N_1824);
and U1903 (N_1903,N_1857,N_1818);
and U1904 (N_1904,N_1813,N_1816);
and U1905 (N_1905,N_1808,N_1855);
nor U1906 (N_1906,N_1820,N_1841);
nand U1907 (N_1907,N_1849,N_1801);
nand U1908 (N_1908,N_1852,N_1837);
nor U1909 (N_1909,N_1851,N_1823);
or U1910 (N_1910,N_1854,N_1850);
or U1911 (N_1911,N_1800,N_1843);
and U1912 (N_1912,N_1825,N_1860);
nand U1913 (N_1913,N_1802,N_1867);
and U1914 (N_1914,N_1869,N_1852);
nor U1915 (N_1915,N_1840,N_1835);
or U1916 (N_1916,N_1858,N_1842);
xor U1917 (N_1917,N_1833,N_1822);
nor U1918 (N_1918,N_1868,N_1825);
or U1919 (N_1919,N_1820,N_1823);
and U1920 (N_1920,N_1839,N_1818);
and U1921 (N_1921,N_1855,N_1810);
nand U1922 (N_1922,N_1874,N_1810);
xor U1923 (N_1923,N_1850,N_1829);
xnor U1924 (N_1924,N_1812,N_1836);
or U1925 (N_1925,N_1865,N_1867);
nor U1926 (N_1926,N_1821,N_1868);
nor U1927 (N_1927,N_1826,N_1850);
or U1928 (N_1928,N_1869,N_1830);
and U1929 (N_1929,N_1822,N_1838);
nor U1930 (N_1930,N_1841,N_1827);
xor U1931 (N_1931,N_1830,N_1810);
and U1932 (N_1932,N_1804,N_1821);
nor U1933 (N_1933,N_1823,N_1847);
and U1934 (N_1934,N_1805,N_1866);
nor U1935 (N_1935,N_1827,N_1846);
and U1936 (N_1936,N_1845,N_1849);
xor U1937 (N_1937,N_1841,N_1874);
and U1938 (N_1938,N_1808,N_1807);
and U1939 (N_1939,N_1831,N_1818);
or U1940 (N_1940,N_1873,N_1804);
and U1941 (N_1941,N_1858,N_1818);
nor U1942 (N_1942,N_1849,N_1813);
or U1943 (N_1943,N_1842,N_1873);
or U1944 (N_1944,N_1837,N_1805);
nor U1945 (N_1945,N_1839,N_1856);
nand U1946 (N_1946,N_1854,N_1814);
and U1947 (N_1947,N_1852,N_1853);
nand U1948 (N_1948,N_1854,N_1831);
and U1949 (N_1949,N_1803,N_1804);
nand U1950 (N_1950,N_1887,N_1919);
nor U1951 (N_1951,N_1894,N_1876);
and U1952 (N_1952,N_1914,N_1881);
or U1953 (N_1953,N_1939,N_1913);
and U1954 (N_1954,N_1899,N_1908);
or U1955 (N_1955,N_1882,N_1893);
and U1956 (N_1956,N_1875,N_1909);
nand U1957 (N_1957,N_1884,N_1883);
and U1958 (N_1958,N_1912,N_1904);
or U1959 (N_1959,N_1937,N_1935);
nand U1960 (N_1960,N_1924,N_1885);
nand U1961 (N_1961,N_1945,N_1901);
and U1962 (N_1962,N_1920,N_1896);
nor U1963 (N_1963,N_1928,N_1949);
and U1964 (N_1964,N_1900,N_1891);
and U1965 (N_1965,N_1932,N_1898);
nor U1966 (N_1966,N_1948,N_1907);
xor U1967 (N_1967,N_1897,N_1933);
or U1968 (N_1968,N_1906,N_1890);
nand U1969 (N_1969,N_1944,N_1895);
xor U1970 (N_1970,N_1910,N_1930);
nand U1971 (N_1971,N_1936,N_1917);
or U1972 (N_1972,N_1931,N_1929);
xnor U1973 (N_1973,N_1892,N_1922);
and U1974 (N_1974,N_1886,N_1921);
and U1975 (N_1975,N_1905,N_1889);
and U1976 (N_1976,N_1878,N_1934);
nand U1977 (N_1977,N_1879,N_1915);
and U1978 (N_1978,N_1916,N_1902);
or U1979 (N_1979,N_1877,N_1946);
or U1980 (N_1980,N_1943,N_1911);
or U1981 (N_1981,N_1941,N_1923);
nor U1982 (N_1982,N_1938,N_1925);
or U1983 (N_1983,N_1942,N_1927);
and U1984 (N_1984,N_1947,N_1918);
nor U1985 (N_1985,N_1926,N_1940);
nor U1986 (N_1986,N_1888,N_1903);
nand U1987 (N_1987,N_1880,N_1894);
nand U1988 (N_1988,N_1904,N_1884);
nand U1989 (N_1989,N_1923,N_1916);
and U1990 (N_1990,N_1887,N_1941);
xnor U1991 (N_1991,N_1885,N_1929);
nand U1992 (N_1992,N_1886,N_1929);
or U1993 (N_1993,N_1907,N_1928);
and U1994 (N_1994,N_1943,N_1934);
and U1995 (N_1995,N_1875,N_1905);
nand U1996 (N_1996,N_1930,N_1933);
nor U1997 (N_1997,N_1945,N_1885);
and U1998 (N_1998,N_1902,N_1933);
and U1999 (N_1999,N_1890,N_1882);
or U2000 (N_2000,N_1878,N_1947);
nor U2001 (N_2001,N_1907,N_1919);
and U2002 (N_2002,N_1911,N_1885);
xor U2003 (N_2003,N_1927,N_1901);
or U2004 (N_2004,N_1935,N_1879);
nand U2005 (N_2005,N_1887,N_1942);
and U2006 (N_2006,N_1919,N_1915);
nand U2007 (N_2007,N_1925,N_1941);
nand U2008 (N_2008,N_1934,N_1923);
nor U2009 (N_2009,N_1949,N_1903);
or U2010 (N_2010,N_1905,N_1937);
nand U2011 (N_2011,N_1884,N_1917);
nand U2012 (N_2012,N_1889,N_1886);
nand U2013 (N_2013,N_1927,N_1932);
or U2014 (N_2014,N_1929,N_1936);
and U2015 (N_2015,N_1883,N_1903);
and U2016 (N_2016,N_1894,N_1897);
and U2017 (N_2017,N_1911,N_1923);
nor U2018 (N_2018,N_1902,N_1907);
nand U2019 (N_2019,N_1908,N_1893);
nand U2020 (N_2020,N_1883,N_1887);
nor U2021 (N_2021,N_1910,N_1886);
and U2022 (N_2022,N_1944,N_1906);
nand U2023 (N_2023,N_1881,N_1904);
nor U2024 (N_2024,N_1900,N_1932);
xnor U2025 (N_2025,N_1999,N_1952);
nand U2026 (N_2026,N_1978,N_1971);
or U2027 (N_2027,N_2020,N_2009);
nor U2028 (N_2028,N_2015,N_1968);
nor U2029 (N_2029,N_1959,N_1954);
nand U2030 (N_2030,N_2010,N_2014);
xor U2031 (N_2031,N_1996,N_1982);
and U2032 (N_2032,N_1989,N_1994);
xnor U2033 (N_2033,N_1970,N_2000);
and U2034 (N_2034,N_1960,N_1976);
and U2035 (N_2035,N_2018,N_1993);
or U2036 (N_2036,N_2004,N_1972);
xor U2037 (N_2037,N_2005,N_1969);
or U2038 (N_2038,N_1987,N_2003);
nand U2039 (N_2039,N_2017,N_2006);
and U2040 (N_2040,N_1951,N_1992);
nand U2041 (N_2041,N_1979,N_2024);
nand U2042 (N_2042,N_1958,N_1990);
xnor U2043 (N_2043,N_1974,N_1975);
or U2044 (N_2044,N_2011,N_1991);
or U2045 (N_2045,N_1984,N_1980);
nand U2046 (N_2046,N_1988,N_1985);
nand U2047 (N_2047,N_1986,N_1997);
nor U2048 (N_2048,N_2008,N_1956);
and U2049 (N_2049,N_1967,N_1998);
nand U2050 (N_2050,N_2016,N_1973);
nand U2051 (N_2051,N_1961,N_2012);
or U2052 (N_2052,N_1953,N_2013);
nor U2053 (N_2053,N_1983,N_1962);
nand U2054 (N_2054,N_2022,N_2007);
nor U2055 (N_2055,N_2002,N_2023);
or U2056 (N_2056,N_1981,N_1955);
and U2057 (N_2057,N_1965,N_1950);
or U2058 (N_2058,N_1977,N_1995);
nand U2059 (N_2059,N_2019,N_1963);
nand U2060 (N_2060,N_1964,N_1957);
or U2061 (N_2061,N_2021,N_1966);
nand U2062 (N_2062,N_2001,N_2000);
xnor U2063 (N_2063,N_2016,N_2001);
nand U2064 (N_2064,N_1962,N_1974);
and U2065 (N_2065,N_1950,N_2002);
or U2066 (N_2066,N_1980,N_1991);
or U2067 (N_2067,N_1956,N_1989);
and U2068 (N_2068,N_2006,N_1951);
and U2069 (N_2069,N_1975,N_1998);
nor U2070 (N_2070,N_1971,N_1997);
nand U2071 (N_2071,N_1979,N_2005);
nor U2072 (N_2072,N_2005,N_1993);
nand U2073 (N_2073,N_1968,N_2005);
nor U2074 (N_2074,N_1973,N_1998);
and U2075 (N_2075,N_1992,N_1994);
or U2076 (N_2076,N_1955,N_1953);
nor U2077 (N_2077,N_1985,N_1973);
or U2078 (N_2078,N_1979,N_1990);
or U2079 (N_2079,N_1995,N_1996);
nor U2080 (N_2080,N_1970,N_2013);
and U2081 (N_2081,N_2015,N_1974);
nor U2082 (N_2082,N_1991,N_1993);
nand U2083 (N_2083,N_2020,N_2023);
or U2084 (N_2084,N_1960,N_2012);
and U2085 (N_2085,N_1999,N_1967);
nor U2086 (N_2086,N_2004,N_2022);
xnor U2087 (N_2087,N_1994,N_1962);
and U2088 (N_2088,N_1959,N_1973);
or U2089 (N_2089,N_2014,N_1998);
nor U2090 (N_2090,N_1954,N_1990);
nand U2091 (N_2091,N_1967,N_1960);
or U2092 (N_2092,N_1954,N_2008);
or U2093 (N_2093,N_2014,N_1956);
nand U2094 (N_2094,N_1993,N_1979);
nand U2095 (N_2095,N_2008,N_1987);
nor U2096 (N_2096,N_1979,N_1992);
nand U2097 (N_2097,N_1951,N_2024);
and U2098 (N_2098,N_2014,N_2008);
and U2099 (N_2099,N_1960,N_2021);
nand U2100 (N_2100,N_2075,N_2064);
and U2101 (N_2101,N_2070,N_2078);
and U2102 (N_2102,N_2035,N_2028);
nand U2103 (N_2103,N_2030,N_2056);
nor U2104 (N_2104,N_2092,N_2032);
and U2105 (N_2105,N_2087,N_2036);
and U2106 (N_2106,N_2026,N_2029);
and U2107 (N_2107,N_2038,N_2068);
or U2108 (N_2108,N_2052,N_2096);
and U2109 (N_2109,N_2031,N_2053);
nor U2110 (N_2110,N_2054,N_2045);
and U2111 (N_2111,N_2097,N_2059);
xnor U2112 (N_2112,N_2050,N_2085);
nand U2113 (N_2113,N_2027,N_2037);
nor U2114 (N_2114,N_2025,N_2098);
xnor U2115 (N_2115,N_2079,N_2048);
or U2116 (N_2116,N_2071,N_2047);
and U2117 (N_2117,N_2088,N_2069);
or U2118 (N_2118,N_2034,N_2072);
nand U2119 (N_2119,N_2093,N_2043);
nand U2120 (N_2120,N_2080,N_2086);
and U2121 (N_2121,N_2099,N_2076);
nand U2122 (N_2122,N_2046,N_2065);
nand U2123 (N_2123,N_2074,N_2091);
or U2124 (N_2124,N_2095,N_2057);
nand U2125 (N_2125,N_2082,N_2084);
nand U2126 (N_2126,N_2042,N_2089);
nand U2127 (N_2127,N_2060,N_2077);
and U2128 (N_2128,N_2033,N_2062);
nor U2129 (N_2129,N_2041,N_2058);
and U2130 (N_2130,N_2055,N_2073);
and U2131 (N_2131,N_2090,N_2049);
nor U2132 (N_2132,N_2051,N_2081);
nor U2133 (N_2133,N_2044,N_2094);
and U2134 (N_2134,N_2067,N_2039);
or U2135 (N_2135,N_2083,N_2066);
or U2136 (N_2136,N_2040,N_2061);
nand U2137 (N_2137,N_2063,N_2050);
and U2138 (N_2138,N_2054,N_2026);
or U2139 (N_2139,N_2062,N_2098);
nor U2140 (N_2140,N_2091,N_2030);
xor U2141 (N_2141,N_2077,N_2069);
and U2142 (N_2142,N_2097,N_2068);
nor U2143 (N_2143,N_2098,N_2077);
nor U2144 (N_2144,N_2098,N_2068);
xor U2145 (N_2145,N_2079,N_2073);
and U2146 (N_2146,N_2044,N_2099);
and U2147 (N_2147,N_2093,N_2065);
or U2148 (N_2148,N_2060,N_2094);
and U2149 (N_2149,N_2077,N_2044);
nor U2150 (N_2150,N_2036,N_2078);
nand U2151 (N_2151,N_2037,N_2061);
nand U2152 (N_2152,N_2082,N_2041);
or U2153 (N_2153,N_2079,N_2040);
or U2154 (N_2154,N_2097,N_2073);
nor U2155 (N_2155,N_2080,N_2039);
nor U2156 (N_2156,N_2062,N_2063);
and U2157 (N_2157,N_2066,N_2095);
xor U2158 (N_2158,N_2099,N_2075);
and U2159 (N_2159,N_2084,N_2055);
nand U2160 (N_2160,N_2096,N_2067);
nand U2161 (N_2161,N_2094,N_2090);
nor U2162 (N_2162,N_2098,N_2087);
xor U2163 (N_2163,N_2074,N_2092);
nand U2164 (N_2164,N_2051,N_2068);
and U2165 (N_2165,N_2083,N_2074);
and U2166 (N_2166,N_2067,N_2045);
nand U2167 (N_2167,N_2061,N_2032);
nor U2168 (N_2168,N_2094,N_2065);
and U2169 (N_2169,N_2078,N_2069);
or U2170 (N_2170,N_2087,N_2031);
or U2171 (N_2171,N_2058,N_2046);
nor U2172 (N_2172,N_2098,N_2066);
and U2173 (N_2173,N_2064,N_2033);
and U2174 (N_2174,N_2054,N_2080);
nand U2175 (N_2175,N_2114,N_2146);
nor U2176 (N_2176,N_2168,N_2126);
nand U2177 (N_2177,N_2138,N_2117);
and U2178 (N_2178,N_2162,N_2110);
and U2179 (N_2179,N_2123,N_2103);
or U2180 (N_2180,N_2130,N_2129);
nor U2181 (N_2181,N_2165,N_2104);
nand U2182 (N_2182,N_2102,N_2158);
or U2183 (N_2183,N_2109,N_2159);
and U2184 (N_2184,N_2133,N_2160);
nor U2185 (N_2185,N_2100,N_2147);
and U2186 (N_2186,N_2134,N_2107);
nor U2187 (N_2187,N_2136,N_2173);
or U2188 (N_2188,N_2112,N_2145);
nor U2189 (N_2189,N_2151,N_2141);
or U2190 (N_2190,N_2161,N_2155);
nand U2191 (N_2191,N_2152,N_2144);
nand U2192 (N_2192,N_2101,N_2111);
or U2193 (N_2193,N_2148,N_2105);
nand U2194 (N_2194,N_2132,N_2113);
nand U2195 (N_2195,N_2116,N_2163);
and U2196 (N_2196,N_2122,N_2131);
nand U2197 (N_2197,N_2127,N_2139);
nand U2198 (N_2198,N_2174,N_2118);
and U2199 (N_2199,N_2135,N_2125);
nor U2200 (N_2200,N_2153,N_2167);
and U2201 (N_2201,N_2115,N_2143);
nand U2202 (N_2202,N_2137,N_2106);
nor U2203 (N_2203,N_2156,N_2172);
or U2204 (N_2204,N_2128,N_2108);
nand U2205 (N_2205,N_2124,N_2157);
nand U2206 (N_2206,N_2150,N_2121);
nor U2207 (N_2207,N_2119,N_2164);
or U2208 (N_2208,N_2149,N_2154);
nand U2209 (N_2209,N_2142,N_2170);
nor U2210 (N_2210,N_2166,N_2120);
nand U2211 (N_2211,N_2171,N_2140);
or U2212 (N_2212,N_2169,N_2112);
and U2213 (N_2213,N_2135,N_2110);
and U2214 (N_2214,N_2116,N_2114);
xor U2215 (N_2215,N_2120,N_2149);
nor U2216 (N_2216,N_2115,N_2102);
nand U2217 (N_2217,N_2169,N_2129);
and U2218 (N_2218,N_2155,N_2139);
or U2219 (N_2219,N_2154,N_2121);
nand U2220 (N_2220,N_2171,N_2125);
nor U2221 (N_2221,N_2127,N_2130);
nand U2222 (N_2222,N_2172,N_2138);
nor U2223 (N_2223,N_2112,N_2137);
and U2224 (N_2224,N_2105,N_2140);
nor U2225 (N_2225,N_2137,N_2136);
and U2226 (N_2226,N_2166,N_2167);
and U2227 (N_2227,N_2148,N_2126);
nand U2228 (N_2228,N_2164,N_2169);
or U2229 (N_2229,N_2161,N_2173);
nor U2230 (N_2230,N_2113,N_2142);
and U2231 (N_2231,N_2128,N_2105);
or U2232 (N_2232,N_2139,N_2124);
or U2233 (N_2233,N_2110,N_2126);
nand U2234 (N_2234,N_2117,N_2148);
nand U2235 (N_2235,N_2113,N_2107);
nand U2236 (N_2236,N_2122,N_2108);
or U2237 (N_2237,N_2140,N_2119);
nor U2238 (N_2238,N_2174,N_2163);
nor U2239 (N_2239,N_2111,N_2100);
and U2240 (N_2240,N_2154,N_2133);
or U2241 (N_2241,N_2121,N_2130);
nand U2242 (N_2242,N_2105,N_2110);
nor U2243 (N_2243,N_2172,N_2147);
nand U2244 (N_2244,N_2170,N_2162);
and U2245 (N_2245,N_2118,N_2144);
and U2246 (N_2246,N_2157,N_2143);
nand U2247 (N_2247,N_2121,N_2167);
and U2248 (N_2248,N_2146,N_2168);
or U2249 (N_2249,N_2105,N_2113);
or U2250 (N_2250,N_2208,N_2245);
or U2251 (N_2251,N_2209,N_2242);
nand U2252 (N_2252,N_2178,N_2221);
or U2253 (N_2253,N_2226,N_2193);
nor U2254 (N_2254,N_2187,N_2195);
nand U2255 (N_2255,N_2202,N_2216);
or U2256 (N_2256,N_2224,N_2211);
and U2257 (N_2257,N_2176,N_2228);
or U2258 (N_2258,N_2233,N_2212);
or U2259 (N_2259,N_2192,N_2239);
xnor U2260 (N_2260,N_2181,N_2227);
or U2261 (N_2261,N_2205,N_2213);
and U2262 (N_2262,N_2194,N_2215);
xnor U2263 (N_2263,N_2214,N_2219);
nand U2264 (N_2264,N_2236,N_2190);
nor U2265 (N_2265,N_2210,N_2198);
nand U2266 (N_2266,N_2201,N_2247);
and U2267 (N_2267,N_2238,N_2184);
nand U2268 (N_2268,N_2180,N_2177);
nor U2269 (N_2269,N_2243,N_2183);
and U2270 (N_2270,N_2218,N_2240);
or U2271 (N_2271,N_2234,N_2199);
nor U2272 (N_2272,N_2237,N_2222);
nand U2273 (N_2273,N_2189,N_2249);
nor U2274 (N_2274,N_2232,N_2207);
nand U2275 (N_2275,N_2200,N_2191);
nor U2276 (N_2276,N_2225,N_2223);
xnor U2277 (N_2277,N_2179,N_2197);
or U2278 (N_2278,N_2188,N_2220);
nand U2279 (N_2279,N_2182,N_2229);
nor U2280 (N_2280,N_2203,N_2204);
nand U2281 (N_2281,N_2175,N_2235);
nand U2282 (N_2282,N_2230,N_2246);
nand U2283 (N_2283,N_2244,N_2231);
nand U2284 (N_2284,N_2217,N_2241);
and U2285 (N_2285,N_2248,N_2196);
and U2286 (N_2286,N_2185,N_2206);
or U2287 (N_2287,N_2186,N_2198);
and U2288 (N_2288,N_2245,N_2195);
xor U2289 (N_2289,N_2215,N_2189);
nor U2290 (N_2290,N_2238,N_2249);
or U2291 (N_2291,N_2176,N_2213);
and U2292 (N_2292,N_2231,N_2241);
xnor U2293 (N_2293,N_2177,N_2176);
xor U2294 (N_2294,N_2202,N_2228);
and U2295 (N_2295,N_2192,N_2222);
xor U2296 (N_2296,N_2209,N_2192);
and U2297 (N_2297,N_2201,N_2175);
and U2298 (N_2298,N_2229,N_2196);
xnor U2299 (N_2299,N_2199,N_2217);
nor U2300 (N_2300,N_2244,N_2242);
and U2301 (N_2301,N_2194,N_2187);
or U2302 (N_2302,N_2209,N_2220);
and U2303 (N_2303,N_2196,N_2232);
and U2304 (N_2304,N_2248,N_2186);
nor U2305 (N_2305,N_2244,N_2177);
nand U2306 (N_2306,N_2229,N_2195);
nor U2307 (N_2307,N_2178,N_2224);
xor U2308 (N_2308,N_2236,N_2219);
and U2309 (N_2309,N_2248,N_2208);
or U2310 (N_2310,N_2207,N_2195);
nand U2311 (N_2311,N_2203,N_2178);
xor U2312 (N_2312,N_2213,N_2187);
nor U2313 (N_2313,N_2194,N_2221);
or U2314 (N_2314,N_2196,N_2184);
or U2315 (N_2315,N_2231,N_2195);
and U2316 (N_2316,N_2204,N_2192);
nor U2317 (N_2317,N_2176,N_2212);
nor U2318 (N_2318,N_2247,N_2211);
and U2319 (N_2319,N_2202,N_2237);
or U2320 (N_2320,N_2237,N_2208);
nand U2321 (N_2321,N_2227,N_2234);
or U2322 (N_2322,N_2207,N_2231);
and U2323 (N_2323,N_2206,N_2247);
nor U2324 (N_2324,N_2217,N_2184);
nand U2325 (N_2325,N_2253,N_2269);
nor U2326 (N_2326,N_2322,N_2289);
and U2327 (N_2327,N_2320,N_2297);
nand U2328 (N_2328,N_2318,N_2310);
nor U2329 (N_2329,N_2317,N_2279);
nor U2330 (N_2330,N_2324,N_2314);
nor U2331 (N_2331,N_2309,N_2255);
or U2332 (N_2332,N_2274,N_2272);
and U2333 (N_2333,N_2281,N_2256);
nor U2334 (N_2334,N_2296,N_2293);
nor U2335 (N_2335,N_2316,N_2267);
or U2336 (N_2336,N_2304,N_2263);
nand U2337 (N_2337,N_2271,N_2257);
xor U2338 (N_2338,N_2268,N_2291);
or U2339 (N_2339,N_2259,N_2299);
nand U2340 (N_2340,N_2292,N_2302);
nor U2341 (N_2341,N_2319,N_2276);
nor U2342 (N_2342,N_2311,N_2273);
or U2343 (N_2343,N_2258,N_2284);
or U2344 (N_2344,N_2303,N_2287);
or U2345 (N_2345,N_2278,N_2251);
or U2346 (N_2346,N_2321,N_2262);
and U2347 (N_2347,N_2254,N_2308);
nand U2348 (N_2348,N_2260,N_2275);
and U2349 (N_2349,N_2306,N_2286);
nor U2350 (N_2350,N_2250,N_2301);
nand U2351 (N_2351,N_2294,N_2277);
nand U2352 (N_2352,N_2312,N_2264);
or U2353 (N_2353,N_2270,N_2285);
and U2354 (N_2354,N_2283,N_2288);
or U2355 (N_2355,N_2290,N_2261);
nand U2356 (N_2356,N_2252,N_2313);
or U2357 (N_2357,N_2295,N_2298);
nand U2358 (N_2358,N_2280,N_2300);
and U2359 (N_2359,N_2315,N_2265);
nand U2360 (N_2360,N_2305,N_2266);
or U2361 (N_2361,N_2307,N_2282);
nand U2362 (N_2362,N_2323,N_2267);
or U2363 (N_2363,N_2321,N_2251);
or U2364 (N_2364,N_2281,N_2280);
and U2365 (N_2365,N_2251,N_2275);
nor U2366 (N_2366,N_2284,N_2286);
nand U2367 (N_2367,N_2257,N_2319);
and U2368 (N_2368,N_2262,N_2313);
or U2369 (N_2369,N_2280,N_2282);
nand U2370 (N_2370,N_2296,N_2270);
or U2371 (N_2371,N_2286,N_2323);
nor U2372 (N_2372,N_2251,N_2284);
nand U2373 (N_2373,N_2312,N_2258);
or U2374 (N_2374,N_2323,N_2319);
xnor U2375 (N_2375,N_2324,N_2285);
nor U2376 (N_2376,N_2254,N_2315);
and U2377 (N_2377,N_2265,N_2259);
nor U2378 (N_2378,N_2284,N_2292);
nor U2379 (N_2379,N_2291,N_2288);
nand U2380 (N_2380,N_2308,N_2294);
nand U2381 (N_2381,N_2317,N_2302);
nand U2382 (N_2382,N_2286,N_2313);
nor U2383 (N_2383,N_2290,N_2320);
and U2384 (N_2384,N_2295,N_2306);
and U2385 (N_2385,N_2262,N_2276);
xor U2386 (N_2386,N_2298,N_2251);
nand U2387 (N_2387,N_2293,N_2301);
nor U2388 (N_2388,N_2284,N_2296);
nor U2389 (N_2389,N_2303,N_2267);
and U2390 (N_2390,N_2277,N_2284);
xor U2391 (N_2391,N_2282,N_2264);
or U2392 (N_2392,N_2316,N_2252);
or U2393 (N_2393,N_2310,N_2282);
nand U2394 (N_2394,N_2322,N_2257);
nor U2395 (N_2395,N_2294,N_2316);
and U2396 (N_2396,N_2321,N_2319);
and U2397 (N_2397,N_2275,N_2257);
and U2398 (N_2398,N_2283,N_2255);
nor U2399 (N_2399,N_2263,N_2322);
nor U2400 (N_2400,N_2393,N_2370);
and U2401 (N_2401,N_2388,N_2377);
nor U2402 (N_2402,N_2334,N_2328);
nor U2403 (N_2403,N_2330,N_2378);
or U2404 (N_2404,N_2342,N_2349);
nand U2405 (N_2405,N_2351,N_2394);
nand U2406 (N_2406,N_2333,N_2327);
nor U2407 (N_2407,N_2354,N_2379);
nor U2408 (N_2408,N_2398,N_2364);
or U2409 (N_2409,N_2362,N_2332);
nand U2410 (N_2410,N_2343,N_2385);
or U2411 (N_2411,N_2365,N_2355);
xnor U2412 (N_2412,N_2360,N_2369);
nand U2413 (N_2413,N_2397,N_2372);
or U2414 (N_2414,N_2371,N_2346);
and U2415 (N_2415,N_2325,N_2340);
or U2416 (N_2416,N_2383,N_2341);
or U2417 (N_2417,N_2348,N_2344);
or U2418 (N_2418,N_2396,N_2338);
xor U2419 (N_2419,N_2337,N_2335);
and U2420 (N_2420,N_2392,N_2367);
and U2421 (N_2421,N_2381,N_2375);
nand U2422 (N_2422,N_2358,N_2384);
nand U2423 (N_2423,N_2363,N_2326);
nor U2424 (N_2424,N_2389,N_2376);
nand U2425 (N_2425,N_2359,N_2391);
nand U2426 (N_2426,N_2361,N_2352);
nor U2427 (N_2427,N_2357,N_2390);
xor U2428 (N_2428,N_2356,N_2373);
and U2429 (N_2429,N_2368,N_2374);
xnor U2430 (N_2430,N_2336,N_2382);
or U2431 (N_2431,N_2339,N_2345);
nand U2432 (N_2432,N_2380,N_2395);
xnor U2433 (N_2433,N_2331,N_2329);
xnor U2434 (N_2434,N_2399,N_2387);
nor U2435 (N_2435,N_2350,N_2386);
nor U2436 (N_2436,N_2353,N_2366);
or U2437 (N_2437,N_2347,N_2368);
or U2438 (N_2438,N_2393,N_2375);
nor U2439 (N_2439,N_2386,N_2381);
nor U2440 (N_2440,N_2385,N_2345);
or U2441 (N_2441,N_2325,N_2387);
and U2442 (N_2442,N_2398,N_2372);
nand U2443 (N_2443,N_2352,N_2334);
nand U2444 (N_2444,N_2328,N_2369);
and U2445 (N_2445,N_2365,N_2374);
nor U2446 (N_2446,N_2350,N_2371);
xnor U2447 (N_2447,N_2325,N_2336);
xnor U2448 (N_2448,N_2359,N_2326);
or U2449 (N_2449,N_2331,N_2333);
nand U2450 (N_2450,N_2355,N_2378);
and U2451 (N_2451,N_2372,N_2379);
and U2452 (N_2452,N_2354,N_2333);
nand U2453 (N_2453,N_2379,N_2378);
xor U2454 (N_2454,N_2384,N_2385);
nor U2455 (N_2455,N_2341,N_2375);
or U2456 (N_2456,N_2364,N_2346);
nand U2457 (N_2457,N_2332,N_2378);
nand U2458 (N_2458,N_2397,N_2366);
or U2459 (N_2459,N_2386,N_2382);
nand U2460 (N_2460,N_2375,N_2344);
nand U2461 (N_2461,N_2394,N_2340);
nor U2462 (N_2462,N_2343,N_2344);
nand U2463 (N_2463,N_2374,N_2370);
nand U2464 (N_2464,N_2386,N_2329);
or U2465 (N_2465,N_2336,N_2381);
nor U2466 (N_2466,N_2335,N_2344);
nand U2467 (N_2467,N_2359,N_2342);
nor U2468 (N_2468,N_2388,N_2380);
nand U2469 (N_2469,N_2365,N_2331);
or U2470 (N_2470,N_2383,N_2384);
nor U2471 (N_2471,N_2389,N_2333);
and U2472 (N_2472,N_2357,N_2399);
nand U2473 (N_2473,N_2360,N_2342);
or U2474 (N_2474,N_2398,N_2374);
nor U2475 (N_2475,N_2459,N_2417);
and U2476 (N_2476,N_2473,N_2448);
or U2477 (N_2477,N_2441,N_2444);
and U2478 (N_2478,N_2427,N_2465);
and U2479 (N_2479,N_2410,N_2467);
and U2480 (N_2480,N_2423,N_2453);
or U2481 (N_2481,N_2446,N_2419);
nor U2482 (N_2482,N_2440,N_2443);
or U2483 (N_2483,N_2470,N_2466);
nand U2484 (N_2484,N_2413,N_2455);
and U2485 (N_2485,N_2421,N_2412);
nand U2486 (N_2486,N_2432,N_2457);
or U2487 (N_2487,N_2431,N_2438);
and U2488 (N_2488,N_2452,N_2463);
nand U2489 (N_2489,N_2430,N_2451);
and U2490 (N_2490,N_2454,N_2418);
xnor U2491 (N_2491,N_2428,N_2469);
xor U2492 (N_2492,N_2400,N_2445);
and U2493 (N_2493,N_2411,N_2436);
or U2494 (N_2494,N_2456,N_2425);
or U2495 (N_2495,N_2442,N_2462);
xnor U2496 (N_2496,N_2404,N_2458);
nand U2497 (N_2497,N_2434,N_2415);
and U2498 (N_2498,N_2461,N_2402);
and U2499 (N_2499,N_2439,N_2409);
and U2500 (N_2500,N_2422,N_2471);
nand U2501 (N_2501,N_2437,N_2426);
nor U2502 (N_2502,N_2408,N_2460);
nand U2503 (N_2503,N_2447,N_2464);
or U2504 (N_2504,N_2450,N_2416);
and U2505 (N_2505,N_2468,N_2472);
and U2506 (N_2506,N_2420,N_2449);
or U2507 (N_2507,N_2424,N_2407);
nor U2508 (N_2508,N_2403,N_2433);
and U2509 (N_2509,N_2435,N_2429);
nand U2510 (N_2510,N_2401,N_2414);
or U2511 (N_2511,N_2406,N_2405);
and U2512 (N_2512,N_2474,N_2457);
xor U2513 (N_2513,N_2443,N_2408);
and U2514 (N_2514,N_2411,N_2426);
nor U2515 (N_2515,N_2412,N_2442);
and U2516 (N_2516,N_2454,N_2410);
and U2517 (N_2517,N_2420,N_2407);
or U2518 (N_2518,N_2413,N_2407);
nor U2519 (N_2519,N_2429,N_2400);
nor U2520 (N_2520,N_2461,N_2429);
nor U2521 (N_2521,N_2413,N_2402);
xnor U2522 (N_2522,N_2448,N_2471);
or U2523 (N_2523,N_2452,N_2442);
and U2524 (N_2524,N_2469,N_2405);
nand U2525 (N_2525,N_2406,N_2452);
nor U2526 (N_2526,N_2457,N_2433);
or U2527 (N_2527,N_2418,N_2436);
or U2528 (N_2528,N_2466,N_2469);
and U2529 (N_2529,N_2415,N_2401);
nor U2530 (N_2530,N_2461,N_2419);
or U2531 (N_2531,N_2466,N_2410);
or U2532 (N_2532,N_2428,N_2410);
nor U2533 (N_2533,N_2445,N_2446);
xnor U2534 (N_2534,N_2419,N_2411);
nor U2535 (N_2535,N_2420,N_2417);
nor U2536 (N_2536,N_2451,N_2435);
and U2537 (N_2537,N_2456,N_2401);
nand U2538 (N_2538,N_2417,N_2469);
xor U2539 (N_2539,N_2438,N_2442);
nor U2540 (N_2540,N_2402,N_2436);
nor U2541 (N_2541,N_2460,N_2467);
and U2542 (N_2542,N_2432,N_2426);
and U2543 (N_2543,N_2435,N_2443);
and U2544 (N_2544,N_2405,N_2441);
nor U2545 (N_2545,N_2433,N_2463);
xor U2546 (N_2546,N_2412,N_2455);
and U2547 (N_2547,N_2402,N_2435);
and U2548 (N_2548,N_2410,N_2421);
xor U2549 (N_2549,N_2442,N_2408);
nor U2550 (N_2550,N_2483,N_2517);
and U2551 (N_2551,N_2490,N_2504);
and U2552 (N_2552,N_2502,N_2496);
and U2553 (N_2553,N_2509,N_2511);
and U2554 (N_2554,N_2545,N_2503);
or U2555 (N_2555,N_2508,N_2528);
and U2556 (N_2556,N_2484,N_2497);
nand U2557 (N_2557,N_2537,N_2531);
or U2558 (N_2558,N_2533,N_2512);
nand U2559 (N_2559,N_2532,N_2506);
nor U2560 (N_2560,N_2507,N_2546);
xnor U2561 (N_2561,N_2485,N_2515);
nor U2562 (N_2562,N_2541,N_2486);
nand U2563 (N_2563,N_2495,N_2478);
and U2564 (N_2564,N_2518,N_2526);
xnor U2565 (N_2565,N_2501,N_2540);
nor U2566 (N_2566,N_2494,N_2534);
nor U2567 (N_2567,N_2480,N_2549);
and U2568 (N_2568,N_2539,N_2498);
nand U2569 (N_2569,N_2547,N_2513);
and U2570 (N_2570,N_2529,N_2482);
and U2571 (N_2571,N_2499,N_2535);
or U2572 (N_2572,N_2505,N_2530);
nand U2573 (N_2573,N_2514,N_2487);
or U2574 (N_2574,N_2476,N_2500);
or U2575 (N_2575,N_2542,N_2519);
and U2576 (N_2576,N_2523,N_2481);
nor U2577 (N_2577,N_2510,N_2522);
nand U2578 (N_2578,N_2548,N_2524);
nor U2579 (N_2579,N_2525,N_2520);
and U2580 (N_2580,N_2475,N_2516);
and U2581 (N_2581,N_2536,N_2493);
and U2582 (N_2582,N_2521,N_2488);
and U2583 (N_2583,N_2492,N_2477);
nand U2584 (N_2584,N_2544,N_2527);
or U2585 (N_2585,N_2479,N_2489);
nor U2586 (N_2586,N_2538,N_2491);
nand U2587 (N_2587,N_2543,N_2483);
xor U2588 (N_2588,N_2513,N_2523);
and U2589 (N_2589,N_2529,N_2500);
xnor U2590 (N_2590,N_2496,N_2481);
and U2591 (N_2591,N_2497,N_2527);
or U2592 (N_2592,N_2512,N_2539);
xor U2593 (N_2593,N_2488,N_2530);
nor U2594 (N_2594,N_2519,N_2521);
nor U2595 (N_2595,N_2478,N_2526);
nor U2596 (N_2596,N_2527,N_2548);
nand U2597 (N_2597,N_2481,N_2510);
nor U2598 (N_2598,N_2502,N_2513);
and U2599 (N_2599,N_2535,N_2497);
or U2600 (N_2600,N_2486,N_2548);
xor U2601 (N_2601,N_2523,N_2508);
and U2602 (N_2602,N_2526,N_2502);
and U2603 (N_2603,N_2546,N_2549);
and U2604 (N_2604,N_2476,N_2485);
and U2605 (N_2605,N_2485,N_2532);
nor U2606 (N_2606,N_2501,N_2547);
or U2607 (N_2607,N_2514,N_2496);
and U2608 (N_2608,N_2487,N_2530);
or U2609 (N_2609,N_2507,N_2534);
nand U2610 (N_2610,N_2534,N_2476);
xnor U2611 (N_2611,N_2501,N_2516);
and U2612 (N_2612,N_2546,N_2542);
and U2613 (N_2613,N_2515,N_2541);
nand U2614 (N_2614,N_2484,N_2510);
nand U2615 (N_2615,N_2541,N_2549);
nor U2616 (N_2616,N_2482,N_2547);
or U2617 (N_2617,N_2532,N_2482);
and U2618 (N_2618,N_2503,N_2476);
nor U2619 (N_2619,N_2505,N_2537);
xnor U2620 (N_2620,N_2516,N_2520);
xor U2621 (N_2621,N_2548,N_2518);
nand U2622 (N_2622,N_2476,N_2492);
nand U2623 (N_2623,N_2532,N_2486);
and U2624 (N_2624,N_2542,N_2540);
and U2625 (N_2625,N_2605,N_2590);
nand U2626 (N_2626,N_2559,N_2561);
and U2627 (N_2627,N_2602,N_2563);
or U2628 (N_2628,N_2610,N_2612);
or U2629 (N_2629,N_2623,N_2587);
or U2630 (N_2630,N_2586,N_2578);
nand U2631 (N_2631,N_2609,N_2614);
nand U2632 (N_2632,N_2568,N_2622);
nor U2633 (N_2633,N_2584,N_2617);
nand U2634 (N_2634,N_2571,N_2572);
xor U2635 (N_2635,N_2582,N_2577);
xnor U2636 (N_2636,N_2593,N_2599);
and U2637 (N_2637,N_2567,N_2594);
or U2638 (N_2638,N_2552,N_2611);
xor U2639 (N_2639,N_2575,N_2619);
nand U2640 (N_2640,N_2580,N_2585);
and U2641 (N_2641,N_2583,N_2558);
and U2642 (N_2642,N_2620,N_2615);
nand U2643 (N_2643,N_2595,N_2591);
xnor U2644 (N_2644,N_2574,N_2607);
nand U2645 (N_2645,N_2606,N_2581);
and U2646 (N_2646,N_2550,N_2600);
nand U2647 (N_2647,N_2624,N_2551);
and U2648 (N_2648,N_2621,N_2603);
xnor U2649 (N_2649,N_2589,N_2553);
and U2650 (N_2650,N_2570,N_2569);
nand U2651 (N_2651,N_2554,N_2597);
nand U2652 (N_2652,N_2573,N_2618);
or U2653 (N_2653,N_2555,N_2557);
and U2654 (N_2654,N_2562,N_2604);
nor U2655 (N_2655,N_2579,N_2556);
or U2656 (N_2656,N_2566,N_2576);
and U2657 (N_2657,N_2592,N_2601);
or U2658 (N_2658,N_2588,N_2596);
and U2659 (N_2659,N_2616,N_2564);
nor U2660 (N_2660,N_2598,N_2613);
and U2661 (N_2661,N_2565,N_2560);
nor U2662 (N_2662,N_2608,N_2585);
and U2663 (N_2663,N_2598,N_2618);
and U2664 (N_2664,N_2559,N_2551);
and U2665 (N_2665,N_2552,N_2580);
nand U2666 (N_2666,N_2582,N_2606);
nand U2667 (N_2667,N_2598,N_2553);
nor U2668 (N_2668,N_2589,N_2619);
or U2669 (N_2669,N_2577,N_2604);
xor U2670 (N_2670,N_2578,N_2603);
and U2671 (N_2671,N_2587,N_2624);
or U2672 (N_2672,N_2615,N_2566);
and U2673 (N_2673,N_2612,N_2614);
nor U2674 (N_2674,N_2552,N_2571);
and U2675 (N_2675,N_2605,N_2554);
nor U2676 (N_2676,N_2603,N_2596);
and U2677 (N_2677,N_2575,N_2590);
or U2678 (N_2678,N_2567,N_2572);
or U2679 (N_2679,N_2550,N_2576);
or U2680 (N_2680,N_2553,N_2613);
or U2681 (N_2681,N_2580,N_2587);
xor U2682 (N_2682,N_2578,N_2570);
nand U2683 (N_2683,N_2616,N_2552);
nor U2684 (N_2684,N_2550,N_2574);
or U2685 (N_2685,N_2563,N_2574);
nand U2686 (N_2686,N_2598,N_2620);
nand U2687 (N_2687,N_2557,N_2615);
nor U2688 (N_2688,N_2621,N_2551);
or U2689 (N_2689,N_2555,N_2554);
xnor U2690 (N_2690,N_2612,N_2623);
nor U2691 (N_2691,N_2574,N_2613);
xnor U2692 (N_2692,N_2562,N_2559);
nor U2693 (N_2693,N_2617,N_2569);
nand U2694 (N_2694,N_2591,N_2606);
xnor U2695 (N_2695,N_2552,N_2620);
and U2696 (N_2696,N_2594,N_2595);
nor U2697 (N_2697,N_2579,N_2575);
or U2698 (N_2698,N_2583,N_2611);
and U2699 (N_2699,N_2604,N_2598);
and U2700 (N_2700,N_2697,N_2664);
nand U2701 (N_2701,N_2642,N_2636);
nand U2702 (N_2702,N_2640,N_2692);
or U2703 (N_2703,N_2628,N_2644);
or U2704 (N_2704,N_2655,N_2646);
nand U2705 (N_2705,N_2651,N_2693);
nor U2706 (N_2706,N_2656,N_2659);
nand U2707 (N_2707,N_2665,N_2688);
and U2708 (N_2708,N_2698,N_2677);
nor U2709 (N_2709,N_2630,N_2694);
and U2710 (N_2710,N_2678,N_2627);
nor U2711 (N_2711,N_2639,N_2668);
nor U2712 (N_2712,N_2674,N_2666);
and U2713 (N_2713,N_2629,N_2658);
nor U2714 (N_2714,N_2626,N_2669);
or U2715 (N_2715,N_2683,N_2641);
xor U2716 (N_2716,N_2648,N_2653);
nor U2717 (N_2717,N_2673,N_2681);
nor U2718 (N_2718,N_2661,N_2637);
and U2719 (N_2719,N_2671,N_2643);
nand U2720 (N_2720,N_2679,N_2625);
nand U2721 (N_2721,N_2657,N_2696);
nor U2722 (N_2722,N_2685,N_2631);
nand U2723 (N_2723,N_2650,N_2645);
nor U2724 (N_2724,N_2676,N_2654);
and U2725 (N_2725,N_2633,N_2690);
xor U2726 (N_2726,N_2634,N_2672);
xor U2727 (N_2727,N_2647,N_2682);
xor U2728 (N_2728,N_2660,N_2662);
or U2729 (N_2729,N_2632,N_2663);
nand U2730 (N_2730,N_2680,N_2686);
nand U2731 (N_2731,N_2687,N_2652);
nor U2732 (N_2732,N_2695,N_2691);
and U2733 (N_2733,N_2684,N_2689);
nor U2734 (N_2734,N_2638,N_2675);
xor U2735 (N_2735,N_2649,N_2670);
nor U2736 (N_2736,N_2699,N_2667);
nand U2737 (N_2737,N_2635,N_2655);
nand U2738 (N_2738,N_2687,N_2672);
nand U2739 (N_2739,N_2630,N_2660);
and U2740 (N_2740,N_2631,N_2661);
and U2741 (N_2741,N_2661,N_2645);
and U2742 (N_2742,N_2696,N_2671);
or U2743 (N_2743,N_2698,N_2669);
xor U2744 (N_2744,N_2627,N_2688);
or U2745 (N_2745,N_2643,N_2672);
nand U2746 (N_2746,N_2627,N_2655);
or U2747 (N_2747,N_2642,N_2646);
nor U2748 (N_2748,N_2648,N_2652);
and U2749 (N_2749,N_2634,N_2650);
nand U2750 (N_2750,N_2636,N_2690);
nand U2751 (N_2751,N_2665,N_2662);
nand U2752 (N_2752,N_2648,N_2672);
nor U2753 (N_2753,N_2656,N_2682);
and U2754 (N_2754,N_2681,N_2648);
or U2755 (N_2755,N_2674,N_2656);
nand U2756 (N_2756,N_2682,N_2668);
and U2757 (N_2757,N_2682,N_2666);
xor U2758 (N_2758,N_2629,N_2681);
and U2759 (N_2759,N_2687,N_2640);
or U2760 (N_2760,N_2646,N_2666);
nor U2761 (N_2761,N_2693,N_2632);
or U2762 (N_2762,N_2649,N_2625);
xnor U2763 (N_2763,N_2667,N_2639);
nor U2764 (N_2764,N_2636,N_2689);
or U2765 (N_2765,N_2668,N_2686);
and U2766 (N_2766,N_2633,N_2682);
nand U2767 (N_2767,N_2641,N_2659);
or U2768 (N_2768,N_2682,N_2670);
or U2769 (N_2769,N_2695,N_2659);
nor U2770 (N_2770,N_2646,N_2664);
and U2771 (N_2771,N_2679,N_2629);
nand U2772 (N_2772,N_2641,N_2682);
nand U2773 (N_2773,N_2639,N_2674);
and U2774 (N_2774,N_2640,N_2656);
or U2775 (N_2775,N_2771,N_2737);
and U2776 (N_2776,N_2706,N_2769);
nand U2777 (N_2777,N_2700,N_2728);
or U2778 (N_2778,N_2765,N_2704);
nand U2779 (N_2779,N_2753,N_2736);
or U2780 (N_2780,N_2767,N_2768);
nand U2781 (N_2781,N_2755,N_2759);
xor U2782 (N_2782,N_2766,N_2761);
nand U2783 (N_2783,N_2701,N_2749);
xnor U2784 (N_2784,N_2734,N_2703);
nor U2785 (N_2785,N_2732,N_2727);
nand U2786 (N_2786,N_2739,N_2744);
and U2787 (N_2787,N_2717,N_2757);
nor U2788 (N_2788,N_2702,N_2731);
and U2789 (N_2789,N_2742,N_2733);
nor U2790 (N_2790,N_2735,N_2773);
or U2791 (N_2791,N_2705,N_2743);
and U2792 (N_2792,N_2756,N_2718);
and U2793 (N_2793,N_2762,N_2730);
nor U2794 (N_2794,N_2751,N_2747);
nor U2795 (N_2795,N_2758,N_2764);
or U2796 (N_2796,N_2774,N_2714);
xnor U2797 (N_2797,N_2772,N_2745);
and U2798 (N_2798,N_2738,N_2711);
or U2799 (N_2799,N_2712,N_2708);
and U2800 (N_2800,N_2707,N_2754);
nand U2801 (N_2801,N_2723,N_2725);
or U2802 (N_2802,N_2740,N_2722);
or U2803 (N_2803,N_2729,N_2716);
nand U2804 (N_2804,N_2750,N_2709);
nand U2805 (N_2805,N_2741,N_2726);
and U2806 (N_2806,N_2746,N_2770);
nand U2807 (N_2807,N_2720,N_2748);
nor U2808 (N_2808,N_2724,N_2710);
or U2809 (N_2809,N_2760,N_2715);
or U2810 (N_2810,N_2721,N_2752);
nor U2811 (N_2811,N_2719,N_2713);
and U2812 (N_2812,N_2763,N_2758);
nand U2813 (N_2813,N_2717,N_2751);
nor U2814 (N_2814,N_2755,N_2742);
nor U2815 (N_2815,N_2725,N_2740);
or U2816 (N_2816,N_2766,N_2728);
nand U2817 (N_2817,N_2722,N_2768);
xor U2818 (N_2818,N_2701,N_2726);
and U2819 (N_2819,N_2766,N_2713);
xor U2820 (N_2820,N_2740,N_2710);
or U2821 (N_2821,N_2744,N_2773);
and U2822 (N_2822,N_2700,N_2711);
nand U2823 (N_2823,N_2767,N_2750);
nand U2824 (N_2824,N_2770,N_2705);
or U2825 (N_2825,N_2763,N_2709);
nand U2826 (N_2826,N_2722,N_2763);
xor U2827 (N_2827,N_2735,N_2771);
nand U2828 (N_2828,N_2729,N_2730);
nor U2829 (N_2829,N_2773,N_2704);
or U2830 (N_2830,N_2733,N_2711);
nor U2831 (N_2831,N_2716,N_2708);
or U2832 (N_2832,N_2764,N_2771);
nor U2833 (N_2833,N_2773,N_2736);
nand U2834 (N_2834,N_2719,N_2764);
nor U2835 (N_2835,N_2746,N_2759);
nor U2836 (N_2836,N_2762,N_2772);
nor U2837 (N_2837,N_2732,N_2721);
nand U2838 (N_2838,N_2748,N_2719);
or U2839 (N_2839,N_2758,N_2754);
or U2840 (N_2840,N_2703,N_2707);
or U2841 (N_2841,N_2715,N_2742);
and U2842 (N_2842,N_2768,N_2741);
or U2843 (N_2843,N_2772,N_2740);
xnor U2844 (N_2844,N_2727,N_2742);
and U2845 (N_2845,N_2707,N_2736);
nor U2846 (N_2846,N_2749,N_2761);
and U2847 (N_2847,N_2742,N_2751);
and U2848 (N_2848,N_2745,N_2728);
and U2849 (N_2849,N_2758,N_2716);
and U2850 (N_2850,N_2842,N_2829);
nand U2851 (N_2851,N_2801,N_2784);
or U2852 (N_2852,N_2789,N_2810);
or U2853 (N_2853,N_2827,N_2797);
and U2854 (N_2854,N_2823,N_2786);
or U2855 (N_2855,N_2809,N_2839);
and U2856 (N_2856,N_2790,N_2830);
nor U2857 (N_2857,N_2845,N_2796);
nor U2858 (N_2858,N_2828,N_2781);
and U2859 (N_2859,N_2791,N_2779);
xor U2860 (N_2860,N_2782,N_2819);
xnor U2861 (N_2861,N_2844,N_2847);
xnor U2862 (N_2862,N_2778,N_2826);
or U2863 (N_2863,N_2846,N_2822);
and U2864 (N_2864,N_2804,N_2788);
nor U2865 (N_2865,N_2808,N_2793);
xnor U2866 (N_2866,N_2848,N_2785);
or U2867 (N_2867,N_2783,N_2814);
and U2868 (N_2868,N_2831,N_2825);
nor U2869 (N_2869,N_2818,N_2805);
nand U2870 (N_2870,N_2833,N_2775);
nand U2871 (N_2871,N_2815,N_2776);
or U2872 (N_2872,N_2806,N_2780);
nor U2873 (N_2873,N_2841,N_2820);
nor U2874 (N_2874,N_2800,N_2799);
and U2875 (N_2875,N_2843,N_2835);
and U2876 (N_2876,N_2838,N_2824);
or U2877 (N_2877,N_2794,N_2837);
or U2878 (N_2878,N_2777,N_2849);
xnor U2879 (N_2879,N_2802,N_2812);
or U2880 (N_2880,N_2817,N_2807);
nand U2881 (N_2881,N_2834,N_2798);
nor U2882 (N_2882,N_2821,N_2840);
nand U2883 (N_2883,N_2795,N_2816);
xor U2884 (N_2884,N_2792,N_2836);
xor U2885 (N_2885,N_2803,N_2787);
nand U2886 (N_2886,N_2832,N_2813);
or U2887 (N_2887,N_2811,N_2796);
nor U2888 (N_2888,N_2817,N_2839);
nor U2889 (N_2889,N_2779,N_2776);
nand U2890 (N_2890,N_2786,N_2820);
nand U2891 (N_2891,N_2821,N_2819);
nand U2892 (N_2892,N_2844,N_2816);
or U2893 (N_2893,N_2784,N_2815);
nor U2894 (N_2894,N_2816,N_2785);
nand U2895 (N_2895,N_2785,N_2837);
nor U2896 (N_2896,N_2786,N_2839);
xor U2897 (N_2897,N_2787,N_2835);
nor U2898 (N_2898,N_2783,N_2820);
xor U2899 (N_2899,N_2844,N_2843);
nor U2900 (N_2900,N_2839,N_2806);
nor U2901 (N_2901,N_2824,N_2827);
and U2902 (N_2902,N_2795,N_2787);
or U2903 (N_2903,N_2821,N_2801);
nand U2904 (N_2904,N_2823,N_2829);
and U2905 (N_2905,N_2849,N_2785);
nor U2906 (N_2906,N_2801,N_2810);
nand U2907 (N_2907,N_2799,N_2778);
or U2908 (N_2908,N_2845,N_2826);
or U2909 (N_2909,N_2829,N_2834);
nor U2910 (N_2910,N_2826,N_2808);
nor U2911 (N_2911,N_2785,N_2835);
xnor U2912 (N_2912,N_2841,N_2788);
or U2913 (N_2913,N_2828,N_2819);
or U2914 (N_2914,N_2834,N_2848);
nor U2915 (N_2915,N_2791,N_2792);
and U2916 (N_2916,N_2836,N_2779);
or U2917 (N_2917,N_2804,N_2815);
or U2918 (N_2918,N_2823,N_2808);
xor U2919 (N_2919,N_2801,N_2790);
or U2920 (N_2920,N_2846,N_2836);
xnor U2921 (N_2921,N_2831,N_2778);
or U2922 (N_2922,N_2806,N_2800);
or U2923 (N_2923,N_2832,N_2801);
nor U2924 (N_2924,N_2780,N_2784);
or U2925 (N_2925,N_2920,N_2901);
nand U2926 (N_2926,N_2900,N_2910);
nor U2927 (N_2927,N_2899,N_2879);
and U2928 (N_2928,N_2907,N_2876);
and U2929 (N_2929,N_2885,N_2856);
xor U2930 (N_2930,N_2863,N_2884);
and U2931 (N_2931,N_2857,N_2904);
nor U2932 (N_2932,N_2875,N_2883);
nand U2933 (N_2933,N_2867,N_2894);
nor U2934 (N_2934,N_2898,N_2871);
nor U2935 (N_2935,N_2914,N_2858);
and U2936 (N_2936,N_2874,N_2872);
nor U2937 (N_2937,N_2919,N_2915);
and U2938 (N_2938,N_2877,N_2896);
xor U2939 (N_2939,N_2866,N_2861);
or U2940 (N_2940,N_2889,N_2859);
nor U2941 (N_2941,N_2860,N_2913);
nand U2942 (N_2942,N_2868,N_2881);
or U2943 (N_2943,N_2923,N_2888);
nor U2944 (N_2944,N_2855,N_2912);
or U2945 (N_2945,N_2902,N_2851);
or U2946 (N_2946,N_2878,N_2869);
nor U2947 (N_2947,N_2882,N_2870);
or U2948 (N_2948,N_2890,N_2908);
or U2949 (N_2949,N_2924,N_2886);
or U2950 (N_2950,N_2905,N_2891);
and U2951 (N_2951,N_2852,N_2864);
xnor U2952 (N_2952,N_2892,N_2850);
xnor U2953 (N_2953,N_2897,N_2862);
nand U2954 (N_2954,N_2895,N_2865);
nand U2955 (N_2955,N_2922,N_2911);
and U2956 (N_2956,N_2918,N_2917);
nor U2957 (N_2957,N_2854,N_2893);
and U2958 (N_2958,N_2873,N_2916);
nor U2959 (N_2959,N_2909,N_2903);
or U2960 (N_2960,N_2880,N_2906);
and U2961 (N_2961,N_2887,N_2853);
and U2962 (N_2962,N_2921,N_2852);
and U2963 (N_2963,N_2917,N_2861);
or U2964 (N_2964,N_2892,N_2862);
nor U2965 (N_2965,N_2862,N_2921);
or U2966 (N_2966,N_2922,N_2915);
xor U2967 (N_2967,N_2862,N_2906);
nor U2968 (N_2968,N_2886,N_2916);
nor U2969 (N_2969,N_2909,N_2899);
nor U2970 (N_2970,N_2881,N_2860);
xor U2971 (N_2971,N_2875,N_2901);
and U2972 (N_2972,N_2911,N_2894);
or U2973 (N_2973,N_2850,N_2890);
or U2974 (N_2974,N_2851,N_2852);
xnor U2975 (N_2975,N_2909,N_2894);
nand U2976 (N_2976,N_2891,N_2877);
and U2977 (N_2977,N_2890,N_2916);
nand U2978 (N_2978,N_2895,N_2852);
nor U2979 (N_2979,N_2854,N_2911);
nand U2980 (N_2980,N_2891,N_2907);
nor U2981 (N_2981,N_2855,N_2905);
nand U2982 (N_2982,N_2924,N_2905);
nor U2983 (N_2983,N_2852,N_2854);
or U2984 (N_2984,N_2913,N_2884);
xor U2985 (N_2985,N_2918,N_2871);
nand U2986 (N_2986,N_2862,N_2852);
and U2987 (N_2987,N_2879,N_2922);
nor U2988 (N_2988,N_2904,N_2883);
and U2989 (N_2989,N_2860,N_2853);
or U2990 (N_2990,N_2858,N_2855);
xnor U2991 (N_2991,N_2882,N_2877);
and U2992 (N_2992,N_2903,N_2873);
xnor U2993 (N_2993,N_2880,N_2854);
or U2994 (N_2994,N_2879,N_2924);
and U2995 (N_2995,N_2871,N_2907);
nor U2996 (N_2996,N_2858,N_2903);
nand U2997 (N_2997,N_2918,N_2921);
nor U2998 (N_2998,N_2915,N_2912);
nor U2999 (N_2999,N_2918,N_2876);
nor UO_0 (O_0,N_2987,N_2979);
nor UO_1 (O_1,N_2939,N_2926);
or UO_2 (O_2,N_2929,N_2976);
and UO_3 (O_3,N_2942,N_2952);
xor UO_4 (O_4,N_2964,N_2949);
nor UO_5 (O_5,N_2948,N_2980);
and UO_6 (O_6,N_2984,N_2941);
nand UO_7 (O_7,N_2967,N_2955);
or UO_8 (O_8,N_2971,N_2994);
or UO_9 (O_9,N_2970,N_2988);
or UO_10 (O_10,N_2961,N_2936);
or UO_11 (O_11,N_2940,N_2953);
and UO_12 (O_12,N_2943,N_2990);
nor UO_13 (O_13,N_2934,N_2935);
nand UO_14 (O_14,N_2944,N_2928);
nand UO_15 (O_15,N_2974,N_2989);
nand UO_16 (O_16,N_2927,N_2946);
xnor UO_17 (O_17,N_2937,N_2975);
xnor UO_18 (O_18,N_2951,N_2983);
or UO_19 (O_19,N_2958,N_2993);
xnor UO_20 (O_20,N_2957,N_2991);
and UO_21 (O_21,N_2959,N_2985);
nand UO_22 (O_22,N_2930,N_2977);
and UO_23 (O_23,N_2947,N_2956);
xor UO_24 (O_24,N_2982,N_2981);
and UO_25 (O_25,N_2986,N_2965);
nand UO_26 (O_26,N_2966,N_2925);
and UO_27 (O_27,N_2973,N_2933);
and UO_28 (O_28,N_2931,N_2945);
nor UO_29 (O_29,N_2960,N_2962);
and UO_30 (O_30,N_2950,N_2997);
or UO_31 (O_31,N_2968,N_2969);
and UO_32 (O_32,N_2998,N_2978);
or UO_33 (O_33,N_2995,N_2932);
xnor UO_34 (O_34,N_2963,N_2992);
or UO_35 (O_35,N_2954,N_2996);
or UO_36 (O_36,N_2999,N_2972);
nor UO_37 (O_37,N_2938,N_2976);
or UO_38 (O_38,N_2943,N_2999);
xor UO_39 (O_39,N_2949,N_2979);
nand UO_40 (O_40,N_2926,N_2949);
nor UO_41 (O_41,N_2941,N_2964);
or UO_42 (O_42,N_2960,N_2983);
xnor UO_43 (O_43,N_2926,N_2966);
nand UO_44 (O_44,N_2956,N_2945);
and UO_45 (O_45,N_2940,N_2963);
nand UO_46 (O_46,N_2984,N_2949);
and UO_47 (O_47,N_2953,N_2998);
nor UO_48 (O_48,N_2929,N_2986);
nor UO_49 (O_49,N_2959,N_2934);
and UO_50 (O_50,N_2959,N_2983);
or UO_51 (O_51,N_2928,N_2947);
nor UO_52 (O_52,N_2981,N_2960);
and UO_53 (O_53,N_2985,N_2929);
nor UO_54 (O_54,N_2995,N_2980);
nor UO_55 (O_55,N_2928,N_2946);
xnor UO_56 (O_56,N_2937,N_2927);
nand UO_57 (O_57,N_2998,N_2973);
xnor UO_58 (O_58,N_2973,N_2949);
nor UO_59 (O_59,N_2940,N_2997);
and UO_60 (O_60,N_2954,N_2967);
nor UO_61 (O_61,N_2929,N_2959);
and UO_62 (O_62,N_2944,N_2929);
or UO_63 (O_63,N_2952,N_2939);
nand UO_64 (O_64,N_2938,N_2952);
xnor UO_65 (O_65,N_2926,N_2936);
xnor UO_66 (O_66,N_2940,N_2958);
and UO_67 (O_67,N_2979,N_2971);
nor UO_68 (O_68,N_2938,N_2940);
or UO_69 (O_69,N_2987,N_2967);
and UO_70 (O_70,N_2964,N_2927);
or UO_71 (O_71,N_2963,N_2953);
nor UO_72 (O_72,N_2969,N_2979);
and UO_73 (O_73,N_2941,N_2986);
nand UO_74 (O_74,N_2945,N_2991);
and UO_75 (O_75,N_2999,N_2934);
nor UO_76 (O_76,N_2942,N_2984);
nand UO_77 (O_77,N_2955,N_2928);
or UO_78 (O_78,N_2955,N_2985);
nand UO_79 (O_79,N_2984,N_2931);
xor UO_80 (O_80,N_2940,N_2990);
nand UO_81 (O_81,N_2961,N_2979);
and UO_82 (O_82,N_2997,N_2936);
and UO_83 (O_83,N_2950,N_2973);
nand UO_84 (O_84,N_2951,N_2949);
and UO_85 (O_85,N_2946,N_2997);
nand UO_86 (O_86,N_2939,N_2951);
or UO_87 (O_87,N_2935,N_2949);
nand UO_88 (O_88,N_2954,N_2997);
nand UO_89 (O_89,N_2975,N_2999);
or UO_90 (O_90,N_2932,N_2956);
or UO_91 (O_91,N_2967,N_2997);
nand UO_92 (O_92,N_2993,N_2950);
nand UO_93 (O_93,N_2936,N_2928);
nand UO_94 (O_94,N_2985,N_2946);
and UO_95 (O_95,N_2980,N_2946);
and UO_96 (O_96,N_2954,N_2973);
and UO_97 (O_97,N_2961,N_2984);
nand UO_98 (O_98,N_2968,N_2986);
nor UO_99 (O_99,N_2972,N_2981);
nor UO_100 (O_100,N_2976,N_2996);
or UO_101 (O_101,N_2943,N_2935);
nor UO_102 (O_102,N_2964,N_2935);
nor UO_103 (O_103,N_2937,N_2968);
nand UO_104 (O_104,N_2957,N_2980);
xnor UO_105 (O_105,N_2929,N_2925);
xor UO_106 (O_106,N_2973,N_2988);
or UO_107 (O_107,N_2999,N_2983);
nand UO_108 (O_108,N_2996,N_2942);
nand UO_109 (O_109,N_2995,N_2948);
xor UO_110 (O_110,N_2948,N_2989);
and UO_111 (O_111,N_2934,N_2958);
or UO_112 (O_112,N_2953,N_2947);
and UO_113 (O_113,N_2948,N_2986);
xnor UO_114 (O_114,N_2981,N_2955);
nand UO_115 (O_115,N_2998,N_2943);
nand UO_116 (O_116,N_2993,N_2937);
and UO_117 (O_117,N_2930,N_2979);
nand UO_118 (O_118,N_2990,N_2978);
and UO_119 (O_119,N_2950,N_2952);
xnor UO_120 (O_120,N_2994,N_2966);
nand UO_121 (O_121,N_2988,N_2946);
xor UO_122 (O_122,N_2930,N_2946);
xor UO_123 (O_123,N_2931,N_2941);
nor UO_124 (O_124,N_2963,N_2984);
and UO_125 (O_125,N_2947,N_2931);
nor UO_126 (O_126,N_2961,N_2971);
and UO_127 (O_127,N_2994,N_2979);
nor UO_128 (O_128,N_2969,N_2935);
and UO_129 (O_129,N_2961,N_2938);
or UO_130 (O_130,N_2954,N_2929);
or UO_131 (O_131,N_2937,N_2953);
nand UO_132 (O_132,N_2945,N_2964);
or UO_133 (O_133,N_2936,N_2931);
nor UO_134 (O_134,N_2988,N_2968);
nand UO_135 (O_135,N_2950,N_2972);
and UO_136 (O_136,N_2979,N_2990);
xnor UO_137 (O_137,N_2938,N_2959);
or UO_138 (O_138,N_2925,N_2946);
and UO_139 (O_139,N_2954,N_2941);
and UO_140 (O_140,N_2975,N_2934);
and UO_141 (O_141,N_2955,N_2987);
or UO_142 (O_142,N_2937,N_2995);
nor UO_143 (O_143,N_2994,N_2951);
or UO_144 (O_144,N_2989,N_2976);
nor UO_145 (O_145,N_2934,N_2947);
nand UO_146 (O_146,N_2988,N_2986);
or UO_147 (O_147,N_2978,N_2987);
or UO_148 (O_148,N_2941,N_2943);
or UO_149 (O_149,N_2989,N_2945);
or UO_150 (O_150,N_2934,N_2970);
nand UO_151 (O_151,N_2936,N_2929);
or UO_152 (O_152,N_2949,N_2947);
nand UO_153 (O_153,N_2942,N_2957);
and UO_154 (O_154,N_2951,N_2967);
or UO_155 (O_155,N_2996,N_2960);
xnor UO_156 (O_156,N_2992,N_2946);
xnor UO_157 (O_157,N_2939,N_2953);
or UO_158 (O_158,N_2984,N_2950);
or UO_159 (O_159,N_2991,N_2949);
nor UO_160 (O_160,N_2983,N_2970);
and UO_161 (O_161,N_2978,N_2928);
and UO_162 (O_162,N_2936,N_2955);
nand UO_163 (O_163,N_2955,N_2957);
or UO_164 (O_164,N_2958,N_2957);
and UO_165 (O_165,N_2996,N_2984);
and UO_166 (O_166,N_2996,N_2974);
xnor UO_167 (O_167,N_2928,N_2966);
nand UO_168 (O_168,N_2997,N_2949);
nand UO_169 (O_169,N_2988,N_2929);
nor UO_170 (O_170,N_2985,N_2967);
or UO_171 (O_171,N_2926,N_2937);
or UO_172 (O_172,N_2981,N_2973);
and UO_173 (O_173,N_2940,N_2982);
and UO_174 (O_174,N_2935,N_2960);
and UO_175 (O_175,N_2986,N_2950);
and UO_176 (O_176,N_2937,N_2956);
or UO_177 (O_177,N_2947,N_2942);
nor UO_178 (O_178,N_2942,N_2978);
nor UO_179 (O_179,N_2936,N_2945);
and UO_180 (O_180,N_2971,N_2936);
nor UO_181 (O_181,N_2946,N_2953);
xnor UO_182 (O_182,N_2931,N_2939);
nor UO_183 (O_183,N_2976,N_2956);
nand UO_184 (O_184,N_2940,N_2977);
nor UO_185 (O_185,N_2940,N_2978);
and UO_186 (O_186,N_2930,N_2972);
or UO_187 (O_187,N_2961,N_2942);
or UO_188 (O_188,N_2990,N_2974);
nor UO_189 (O_189,N_2964,N_2961);
nand UO_190 (O_190,N_2968,N_2997);
nand UO_191 (O_191,N_2940,N_2971);
or UO_192 (O_192,N_2997,N_2927);
and UO_193 (O_193,N_2933,N_2983);
and UO_194 (O_194,N_2976,N_2966);
nand UO_195 (O_195,N_2950,N_2960);
nand UO_196 (O_196,N_2990,N_2960);
and UO_197 (O_197,N_2936,N_2964);
and UO_198 (O_198,N_2929,N_2945);
nor UO_199 (O_199,N_2980,N_2998);
and UO_200 (O_200,N_2963,N_2979);
xor UO_201 (O_201,N_2969,N_2948);
and UO_202 (O_202,N_2959,N_2968);
nand UO_203 (O_203,N_2931,N_2956);
xnor UO_204 (O_204,N_2965,N_2964);
or UO_205 (O_205,N_2925,N_2989);
nor UO_206 (O_206,N_2964,N_2926);
xnor UO_207 (O_207,N_2968,N_2966);
nor UO_208 (O_208,N_2976,N_2970);
or UO_209 (O_209,N_2988,N_2957);
or UO_210 (O_210,N_2931,N_2993);
nand UO_211 (O_211,N_2946,N_2934);
nor UO_212 (O_212,N_2995,N_2961);
or UO_213 (O_213,N_2980,N_2975);
or UO_214 (O_214,N_2969,N_2942);
nor UO_215 (O_215,N_2984,N_2986);
xnor UO_216 (O_216,N_2993,N_2977);
nand UO_217 (O_217,N_2929,N_2969);
or UO_218 (O_218,N_2961,N_2927);
or UO_219 (O_219,N_2993,N_2994);
xor UO_220 (O_220,N_2987,N_2990);
nand UO_221 (O_221,N_2967,N_2968);
or UO_222 (O_222,N_2986,N_2947);
nor UO_223 (O_223,N_2958,N_2997);
and UO_224 (O_224,N_2980,N_2984);
or UO_225 (O_225,N_2961,N_2943);
or UO_226 (O_226,N_2980,N_2982);
nor UO_227 (O_227,N_2925,N_2926);
or UO_228 (O_228,N_2942,N_2964);
and UO_229 (O_229,N_2925,N_2969);
nand UO_230 (O_230,N_2995,N_2981);
nor UO_231 (O_231,N_2934,N_2944);
or UO_232 (O_232,N_2997,N_2981);
or UO_233 (O_233,N_2927,N_2968);
nand UO_234 (O_234,N_2985,N_2998);
or UO_235 (O_235,N_2956,N_2948);
xor UO_236 (O_236,N_2966,N_2985);
or UO_237 (O_237,N_2965,N_2946);
nor UO_238 (O_238,N_2949,N_2976);
and UO_239 (O_239,N_2993,N_2936);
or UO_240 (O_240,N_2955,N_2992);
xor UO_241 (O_241,N_2991,N_2995);
nand UO_242 (O_242,N_2929,N_2931);
and UO_243 (O_243,N_2941,N_2980);
nand UO_244 (O_244,N_2961,N_2997);
nand UO_245 (O_245,N_2978,N_2984);
nor UO_246 (O_246,N_2982,N_2944);
and UO_247 (O_247,N_2962,N_2988);
and UO_248 (O_248,N_2995,N_2998);
nor UO_249 (O_249,N_2926,N_2934);
and UO_250 (O_250,N_2942,N_2977);
and UO_251 (O_251,N_2978,N_2958);
and UO_252 (O_252,N_2932,N_2980);
nand UO_253 (O_253,N_2955,N_2991);
xnor UO_254 (O_254,N_2982,N_2941);
or UO_255 (O_255,N_2942,N_2979);
nor UO_256 (O_256,N_2982,N_2992);
nand UO_257 (O_257,N_2947,N_2977);
nor UO_258 (O_258,N_2958,N_2964);
nand UO_259 (O_259,N_2928,N_2987);
nand UO_260 (O_260,N_2960,N_2972);
xor UO_261 (O_261,N_2954,N_2978);
or UO_262 (O_262,N_2988,N_2964);
or UO_263 (O_263,N_2925,N_2984);
or UO_264 (O_264,N_2998,N_2967);
or UO_265 (O_265,N_2941,N_2942);
xor UO_266 (O_266,N_2994,N_2955);
xnor UO_267 (O_267,N_2936,N_2990);
nor UO_268 (O_268,N_2986,N_2942);
nand UO_269 (O_269,N_2975,N_2962);
nor UO_270 (O_270,N_2939,N_2933);
and UO_271 (O_271,N_2936,N_2952);
nand UO_272 (O_272,N_2990,N_2948);
or UO_273 (O_273,N_2997,N_2951);
and UO_274 (O_274,N_2981,N_2953);
nor UO_275 (O_275,N_2984,N_2967);
nor UO_276 (O_276,N_2998,N_2993);
or UO_277 (O_277,N_2953,N_2945);
and UO_278 (O_278,N_2933,N_2962);
nand UO_279 (O_279,N_2999,N_2990);
and UO_280 (O_280,N_2961,N_2947);
nor UO_281 (O_281,N_2956,N_2999);
xnor UO_282 (O_282,N_2982,N_2955);
nand UO_283 (O_283,N_2942,N_2940);
or UO_284 (O_284,N_2947,N_2959);
and UO_285 (O_285,N_2994,N_2940);
and UO_286 (O_286,N_2938,N_2986);
or UO_287 (O_287,N_2974,N_2985);
nand UO_288 (O_288,N_2996,N_2964);
or UO_289 (O_289,N_2950,N_2954);
or UO_290 (O_290,N_2954,N_2927);
xnor UO_291 (O_291,N_2964,N_2974);
or UO_292 (O_292,N_2954,N_2939);
and UO_293 (O_293,N_2951,N_2930);
or UO_294 (O_294,N_2976,N_2990);
or UO_295 (O_295,N_2965,N_2999);
nor UO_296 (O_296,N_2968,N_2930);
or UO_297 (O_297,N_2963,N_2993);
and UO_298 (O_298,N_2935,N_2980);
nand UO_299 (O_299,N_2958,N_2952);
and UO_300 (O_300,N_2966,N_2987);
nor UO_301 (O_301,N_2986,N_2979);
nand UO_302 (O_302,N_2990,N_2998);
and UO_303 (O_303,N_2938,N_2941);
or UO_304 (O_304,N_2988,N_2943);
or UO_305 (O_305,N_2969,N_2989);
nor UO_306 (O_306,N_2959,N_2972);
or UO_307 (O_307,N_2950,N_2955);
or UO_308 (O_308,N_2982,N_2999);
nor UO_309 (O_309,N_2996,N_2947);
nor UO_310 (O_310,N_2952,N_2966);
nor UO_311 (O_311,N_2975,N_2979);
or UO_312 (O_312,N_2991,N_2987);
or UO_313 (O_313,N_2938,N_2937);
nor UO_314 (O_314,N_2973,N_2929);
nand UO_315 (O_315,N_2979,N_2944);
nand UO_316 (O_316,N_2927,N_2970);
nand UO_317 (O_317,N_2930,N_2962);
nor UO_318 (O_318,N_2960,N_2999);
xor UO_319 (O_319,N_2999,N_2997);
or UO_320 (O_320,N_2931,N_2979);
or UO_321 (O_321,N_2963,N_2980);
and UO_322 (O_322,N_2934,N_2993);
nand UO_323 (O_323,N_2941,N_2991);
and UO_324 (O_324,N_2973,N_2972);
or UO_325 (O_325,N_2937,N_2933);
nand UO_326 (O_326,N_2998,N_2932);
and UO_327 (O_327,N_2982,N_2962);
or UO_328 (O_328,N_2966,N_2967);
nor UO_329 (O_329,N_2974,N_2960);
xnor UO_330 (O_330,N_2986,N_2940);
or UO_331 (O_331,N_2975,N_2994);
nor UO_332 (O_332,N_2978,N_2985);
nor UO_333 (O_333,N_2925,N_2941);
or UO_334 (O_334,N_2953,N_2985);
xnor UO_335 (O_335,N_2973,N_2990);
xor UO_336 (O_336,N_2961,N_2987);
nor UO_337 (O_337,N_2981,N_2965);
or UO_338 (O_338,N_2980,N_2927);
or UO_339 (O_339,N_2983,N_2990);
nor UO_340 (O_340,N_2993,N_2989);
and UO_341 (O_341,N_2968,N_2962);
and UO_342 (O_342,N_2961,N_2940);
nand UO_343 (O_343,N_2926,N_2986);
or UO_344 (O_344,N_2990,N_2961);
or UO_345 (O_345,N_2987,N_2948);
or UO_346 (O_346,N_2952,N_2935);
and UO_347 (O_347,N_2980,N_2991);
and UO_348 (O_348,N_2928,N_2980);
nand UO_349 (O_349,N_2948,N_2955);
or UO_350 (O_350,N_2957,N_2950);
or UO_351 (O_351,N_2976,N_2999);
nand UO_352 (O_352,N_2930,N_2955);
and UO_353 (O_353,N_2962,N_2983);
or UO_354 (O_354,N_2978,N_2983);
nor UO_355 (O_355,N_2996,N_2998);
or UO_356 (O_356,N_2930,N_2958);
nor UO_357 (O_357,N_2978,N_2970);
nand UO_358 (O_358,N_2999,N_2929);
and UO_359 (O_359,N_2930,N_2987);
or UO_360 (O_360,N_2956,N_2955);
nand UO_361 (O_361,N_2970,N_2942);
nand UO_362 (O_362,N_2992,N_2980);
nor UO_363 (O_363,N_2971,N_2985);
and UO_364 (O_364,N_2968,N_2949);
nand UO_365 (O_365,N_2987,N_2965);
xor UO_366 (O_366,N_2971,N_2954);
nand UO_367 (O_367,N_2939,N_2999);
and UO_368 (O_368,N_2975,N_2977);
and UO_369 (O_369,N_2935,N_2988);
nor UO_370 (O_370,N_2950,N_2925);
and UO_371 (O_371,N_2925,N_2980);
and UO_372 (O_372,N_2926,N_2941);
and UO_373 (O_373,N_2927,N_2935);
nor UO_374 (O_374,N_2998,N_2937);
xnor UO_375 (O_375,N_2926,N_2961);
or UO_376 (O_376,N_2977,N_2925);
or UO_377 (O_377,N_2930,N_2933);
or UO_378 (O_378,N_2946,N_2943);
or UO_379 (O_379,N_2996,N_2995);
xnor UO_380 (O_380,N_2957,N_2926);
or UO_381 (O_381,N_2928,N_2945);
or UO_382 (O_382,N_2945,N_2973);
and UO_383 (O_383,N_2958,N_2939);
and UO_384 (O_384,N_2969,N_2933);
nand UO_385 (O_385,N_2950,N_2976);
xnor UO_386 (O_386,N_2972,N_2944);
and UO_387 (O_387,N_2930,N_2990);
nand UO_388 (O_388,N_2969,N_2995);
or UO_389 (O_389,N_2985,N_2925);
xnor UO_390 (O_390,N_2956,N_2927);
and UO_391 (O_391,N_2955,N_2976);
nor UO_392 (O_392,N_2952,N_2951);
nor UO_393 (O_393,N_2956,N_2971);
xor UO_394 (O_394,N_2973,N_2947);
and UO_395 (O_395,N_2965,N_2985);
and UO_396 (O_396,N_2956,N_2969);
and UO_397 (O_397,N_2991,N_2942);
or UO_398 (O_398,N_2982,N_2984);
nand UO_399 (O_399,N_2971,N_2965);
or UO_400 (O_400,N_2927,N_2940);
or UO_401 (O_401,N_2949,N_2946);
xnor UO_402 (O_402,N_2971,N_2946);
nor UO_403 (O_403,N_2970,N_2967);
nand UO_404 (O_404,N_2974,N_2992);
or UO_405 (O_405,N_2936,N_2958);
or UO_406 (O_406,N_2954,N_2977);
or UO_407 (O_407,N_2991,N_2959);
nor UO_408 (O_408,N_2945,N_2933);
and UO_409 (O_409,N_2931,N_2990);
nor UO_410 (O_410,N_2946,N_2962);
and UO_411 (O_411,N_2944,N_2998);
nor UO_412 (O_412,N_2979,N_2962);
nor UO_413 (O_413,N_2950,N_2992);
nand UO_414 (O_414,N_2966,N_2991);
nand UO_415 (O_415,N_2961,N_2958);
xor UO_416 (O_416,N_2951,N_2948);
nand UO_417 (O_417,N_2952,N_2949);
or UO_418 (O_418,N_2938,N_2985);
or UO_419 (O_419,N_2936,N_2986);
and UO_420 (O_420,N_2936,N_2934);
nor UO_421 (O_421,N_2977,N_2983);
nor UO_422 (O_422,N_2986,N_2983);
nor UO_423 (O_423,N_2933,N_2963);
nor UO_424 (O_424,N_2958,N_2927);
and UO_425 (O_425,N_2941,N_2936);
and UO_426 (O_426,N_2971,N_2957);
and UO_427 (O_427,N_2971,N_2962);
nor UO_428 (O_428,N_2936,N_2988);
and UO_429 (O_429,N_2953,N_2933);
and UO_430 (O_430,N_2990,N_2966);
or UO_431 (O_431,N_2960,N_2951);
and UO_432 (O_432,N_2933,N_2942);
nand UO_433 (O_433,N_2950,N_2964);
or UO_434 (O_434,N_2992,N_2953);
nand UO_435 (O_435,N_2942,N_2980);
xor UO_436 (O_436,N_2992,N_2966);
or UO_437 (O_437,N_2931,N_2930);
nand UO_438 (O_438,N_2979,N_2925);
or UO_439 (O_439,N_2985,N_2932);
nor UO_440 (O_440,N_2954,N_2959);
xor UO_441 (O_441,N_2972,N_2947);
nand UO_442 (O_442,N_2951,N_2976);
nor UO_443 (O_443,N_2963,N_2941);
nand UO_444 (O_444,N_2939,N_2962);
and UO_445 (O_445,N_2930,N_2952);
nor UO_446 (O_446,N_2931,N_2961);
nor UO_447 (O_447,N_2981,N_2925);
xor UO_448 (O_448,N_2998,N_2952);
and UO_449 (O_449,N_2948,N_2964);
or UO_450 (O_450,N_2963,N_2952);
or UO_451 (O_451,N_2936,N_2946);
nand UO_452 (O_452,N_2937,N_2967);
or UO_453 (O_453,N_2981,N_2970);
and UO_454 (O_454,N_2974,N_2948);
or UO_455 (O_455,N_2976,N_2943);
nor UO_456 (O_456,N_2932,N_2947);
nor UO_457 (O_457,N_2947,N_2955);
nor UO_458 (O_458,N_2990,N_2958);
or UO_459 (O_459,N_2932,N_2952);
xor UO_460 (O_460,N_2971,N_2968);
or UO_461 (O_461,N_2991,N_2954);
nor UO_462 (O_462,N_2990,N_2981);
xor UO_463 (O_463,N_2932,N_2953);
and UO_464 (O_464,N_2987,N_2927);
nand UO_465 (O_465,N_2950,N_2930);
and UO_466 (O_466,N_2973,N_2940);
xnor UO_467 (O_467,N_2999,N_2944);
nand UO_468 (O_468,N_2998,N_2988);
nor UO_469 (O_469,N_2991,N_2931);
and UO_470 (O_470,N_2965,N_2930);
or UO_471 (O_471,N_2998,N_2936);
nor UO_472 (O_472,N_2957,N_2977);
nor UO_473 (O_473,N_2981,N_2980);
nor UO_474 (O_474,N_2972,N_2976);
nor UO_475 (O_475,N_2993,N_2991);
or UO_476 (O_476,N_2977,N_2962);
nor UO_477 (O_477,N_2966,N_2950);
or UO_478 (O_478,N_2938,N_2956);
xnor UO_479 (O_479,N_2930,N_2943);
or UO_480 (O_480,N_2954,N_2993);
nor UO_481 (O_481,N_2995,N_2955);
nand UO_482 (O_482,N_2948,N_2929);
or UO_483 (O_483,N_2931,N_2953);
nand UO_484 (O_484,N_2995,N_2958);
or UO_485 (O_485,N_2933,N_2944);
and UO_486 (O_486,N_2990,N_2991);
and UO_487 (O_487,N_2984,N_2926);
and UO_488 (O_488,N_2971,N_2963);
nand UO_489 (O_489,N_2980,N_2939);
and UO_490 (O_490,N_2930,N_2926);
xor UO_491 (O_491,N_2940,N_2946);
and UO_492 (O_492,N_2957,N_2997);
or UO_493 (O_493,N_2950,N_2962);
nor UO_494 (O_494,N_2966,N_2941);
xor UO_495 (O_495,N_2980,N_2986);
nand UO_496 (O_496,N_2926,N_2983);
or UO_497 (O_497,N_2977,N_2994);
nand UO_498 (O_498,N_2982,N_2957);
and UO_499 (O_499,N_2975,N_2973);
endmodule