module basic_1000_10000_1500_20_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_429,In_244);
nand U1 (N_1,In_87,In_631);
nor U2 (N_2,In_746,In_906);
xor U3 (N_3,In_627,In_662);
and U4 (N_4,In_107,In_865);
nand U5 (N_5,In_79,In_361);
or U6 (N_6,In_22,In_702);
nor U7 (N_7,In_4,In_656);
xnor U8 (N_8,In_329,In_929);
nand U9 (N_9,In_667,In_949);
and U10 (N_10,In_821,In_710);
nand U11 (N_11,In_278,In_80);
or U12 (N_12,In_208,In_103);
and U13 (N_13,In_486,In_445);
nor U14 (N_14,In_143,In_831);
nor U15 (N_15,In_636,In_468);
nor U16 (N_16,In_839,In_705);
nor U17 (N_17,In_150,In_653);
nand U18 (N_18,In_98,In_297);
nand U19 (N_19,In_158,In_372);
nor U20 (N_20,In_265,In_47);
and U21 (N_21,In_401,In_536);
nand U22 (N_22,In_780,In_398);
or U23 (N_23,In_460,In_211);
and U24 (N_24,In_266,In_320);
nor U25 (N_25,In_779,In_454);
nand U26 (N_26,In_415,In_974);
nor U27 (N_27,In_583,In_584);
nand U28 (N_28,In_254,In_609);
and U29 (N_29,In_983,In_168);
and U30 (N_30,In_255,In_473);
nand U31 (N_31,In_748,In_531);
or U32 (N_32,In_26,In_959);
nor U33 (N_33,In_623,In_451);
or U34 (N_34,In_840,In_160);
and U35 (N_35,In_901,In_695);
nor U36 (N_36,In_835,In_61);
nand U37 (N_37,In_194,In_503);
or U38 (N_38,In_802,In_992);
or U39 (N_39,In_533,In_170);
and U40 (N_40,In_961,In_355);
nand U41 (N_41,In_784,In_389);
or U42 (N_42,In_875,In_55);
and U43 (N_43,In_792,In_326);
or U44 (N_44,In_562,In_616);
and U45 (N_45,In_210,In_152);
and U46 (N_46,In_50,In_76);
nand U47 (N_47,In_713,In_427);
nor U48 (N_48,In_387,In_546);
and U49 (N_49,In_809,In_847);
xnor U50 (N_50,In_359,In_89);
xnor U51 (N_51,In_595,In_6);
or U52 (N_52,In_153,In_880);
or U53 (N_53,In_733,In_947);
and U54 (N_54,In_505,In_5);
or U55 (N_55,In_925,In_741);
nand U56 (N_56,In_159,In_393);
and U57 (N_57,In_338,In_491);
and U58 (N_58,In_969,In_514);
xnor U59 (N_59,In_485,In_140);
and U60 (N_60,In_30,In_314);
nand U61 (N_61,In_467,In_489);
nand U62 (N_62,In_722,In_442);
xnor U63 (N_63,In_275,In_568);
and U64 (N_64,In_664,In_180);
nor U65 (N_65,In_206,In_414);
and U66 (N_66,In_866,In_330);
nand U67 (N_67,In_367,In_758);
nor U68 (N_68,In_498,In_948);
xor U69 (N_69,In_85,In_776);
or U70 (N_70,In_321,In_986);
or U71 (N_71,In_692,In_886);
nand U72 (N_72,In_296,In_812);
xnor U73 (N_73,In_714,In_214);
and U74 (N_74,In_997,In_663);
and U75 (N_75,In_262,In_870);
nand U76 (N_76,In_859,In_786);
nor U77 (N_77,In_551,In_785);
and U78 (N_78,In_704,In_224);
nand U79 (N_79,In_896,In_370);
and U80 (N_80,In_680,In_417);
nor U81 (N_81,In_69,In_665);
and U82 (N_82,In_548,In_298);
nand U83 (N_83,In_299,In_543);
nand U84 (N_84,In_365,In_773);
or U85 (N_85,In_540,In_783);
xor U86 (N_86,In_340,In_71);
or U87 (N_87,In_617,In_962);
nor U88 (N_88,In_286,In_926);
or U89 (N_89,In_226,In_407);
xor U90 (N_90,In_237,In_698);
xnor U91 (N_91,In_577,In_761);
nand U92 (N_92,In_283,In_918);
and U93 (N_93,In_893,In_753);
nand U94 (N_94,In_911,In_432);
or U95 (N_95,In_131,In_256);
and U96 (N_96,In_740,In_440);
nand U97 (N_97,In_317,In_234);
or U98 (N_98,In_894,In_149);
nor U99 (N_99,In_720,In_198);
and U100 (N_100,In_905,In_300);
and U101 (N_101,In_322,In_112);
nand U102 (N_102,In_466,In_731);
and U103 (N_103,In_556,In_304);
and U104 (N_104,In_481,In_878);
or U105 (N_105,In_825,In_479);
and U106 (N_106,In_204,In_520);
or U107 (N_107,In_411,In_738);
and U108 (N_108,In_476,In_483);
xnor U109 (N_109,In_110,In_899);
nand U110 (N_110,In_789,In_348);
or U111 (N_111,In_449,In_328);
xor U112 (N_112,In_100,In_666);
or U113 (N_113,In_176,In_890);
or U114 (N_114,In_989,In_693);
and U115 (N_115,In_601,In_646);
nor U116 (N_116,In_537,In_426);
and U117 (N_117,In_225,In_209);
and U118 (N_118,In_579,In_67);
and U119 (N_119,In_567,In_863);
or U120 (N_120,In_308,In_86);
nor U121 (N_121,In_566,In_178);
xnor U122 (N_122,In_757,In_815);
nand U123 (N_123,In_988,In_645);
xnor U124 (N_124,In_124,In_516);
nor U125 (N_125,In_220,In_174);
nor U126 (N_126,In_72,In_655);
nor U127 (N_127,In_288,In_972);
and U128 (N_128,In_597,In_238);
or U129 (N_129,In_324,In_826);
nand U130 (N_130,In_38,In_25);
or U131 (N_131,In_724,In_276);
nor U132 (N_132,In_74,In_223);
nor U133 (N_133,In_699,In_844);
xor U134 (N_134,In_712,In_356);
nor U135 (N_135,In_795,In_763);
nand U136 (N_136,In_381,In_767);
xor U137 (N_137,In_438,In_343);
xnor U138 (N_138,In_626,In_569);
and U139 (N_139,In_777,In_943);
nand U140 (N_140,In_728,In_790);
or U141 (N_141,In_129,In_325);
xnor U142 (N_142,In_0,In_212);
nor U143 (N_143,In_694,In_11);
nand U144 (N_144,In_251,In_990);
or U145 (N_145,In_994,In_402);
and U146 (N_146,In_654,In_121);
xnor U147 (N_147,In_690,In_35);
nand U148 (N_148,In_871,In_574);
nand U149 (N_149,In_145,In_135);
or U150 (N_150,In_669,In_412);
nor U151 (N_151,In_49,In_205);
or U152 (N_152,In_778,In_227);
xnor U153 (N_153,In_147,In_599);
nor U154 (N_154,In_33,In_719);
nor U155 (N_155,In_727,In_456);
and U156 (N_156,In_165,In_846);
xnor U157 (N_157,In_382,In_788);
and U158 (N_158,In_101,In_104);
nand U159 (N_159,In_782,In_682);
nor U160 (N_160,In_315,In_855);
nand U161 (N_161,In_162,In_993);
or U162 (N_162,In_106,In_29);
nor U163 (N_163,In_512,In_109);
nand U164 (N_164,In_43,In_7);
or U165 (N_165,In_68,In_120);
xnor U166 (N_166,In_229,In_130);
or U167 (N_167,In_923,In_84);
nor U168 (N_168,In_903,In_399);
and U169 (N_169,In_292,In_658);
and U170 (N_170,In_751,In_183);
or U171 (N_171,In_290,In_632);
and U172 (N_172,In_916,In_824);
xnor U173 (N_173,In_629,In_587);
and U174 (N_174,In_277,In_798);
or U175 (N_175,In_388,In_671);
nor U176 (N_176,In_478,In_346);
xor U177 (N_177,In_799,In_917);
or U178 (N_178,In_607,In_138);
or U179 (N_179,In_810,In_676);
and U180 (N_180,In_827,In_832);
and U181 (N_181,In_708,In_358);
nor U182 (N_182,In_873,In_884);
nand U183 (N_183,In_703,In_122);
nand U184 (N_184,In_634,In_900);
nor U185 (N_185,In_697,In_557);
xnor U186 (N_186,In_439,In_58);
and U187 (N_187,In_615,In_218);
nand U188 (N_188,In_726,In_681);
xor U189 (N_189,In_527,In_549);
and U190 (N_190,In_700,In_369);
and U191 (N_191,In_435,In_497);
and U192 (N_192,In_858,In_806);
and U193 (N_193,In_443,In_270);
and U194 (N_194,In_199,In_133);
or U195 (N_195,In_685,In_553);
nand U196 (N_196,In_572,In_334);
nand U197 (N_197,In_307,In_24);
xor U198 (N_198,In_633,In_219);
and U199 (N_199,In_570,In_97);
xor U200 (N_200,In_960,In_602);
and U201 (N_201,In_725,In_189);
and U202 (N_202,In_215,In_472);
xor U203 (N_203,In_613,In_269);
and U204 (N_204,In_446,In_172);
and U205 (N_205,In_544,In_987);
nand U206 (N_206,In_425,In_213);
or U207 (N_207,In_507,In_196);
and U208 (N_208,In_457,In_157);
nand U209 (N_209,In_876,In_813);
nand U210 (N_210,In_93,In_768);
nor U211 (N_211,In_822,In_181);
and U212 (N_212,In_828,In_965);
nand U213 (N_213,In_953,In_892);
and U214 (N_214,In_921,In_21);
nand U215 (N_215,In_829,In_762);
and U216 (N_216,In_709,In_848);
and U217 (N_217,In_316,In_715);
and U218 (N_218,In_409,In_56);
or U219 (N_219,In_868,In_596);
or U220 (N_220,In_590,In_464);
or U221 (N_221,In_838,In_955);
or U222 (N_222,In_281,In_999);
xor U223 (N_223,In_766,In_267);
nor U224 (N_224,In_547,In_462);
and U225 (N_225,In_380,In_524);
xnor U226 (N_226,In_877,In_723);
nand U227 (N_227,In_854,In_470);
nand U228 (N_228,In_554,In_287);
nor U229 (N_229,In_657,In_18);
nor U230 (N_230,In_650,In_15);
nor U231 (N_231,In_60,In_352);
nor U232 (N_232,In_578,In_236);
nand U233 (N_233,In_985,In_23);
or U234 (N_234,In_430,In_593);
and U235 (N_235,In_530,In_418);
nor U236 (N_236,In_408,In_672);
nand U237 (N_237,In_353,In_744);
nor U238 (N_238,In_115,In_771);
nor U239 (N_239,In_250,In_175);
and U240 (N_240,In_336,In_461);
and U241 (N_241,In_83,In_207);
and U242 (N_242,In_291,In_200);
and U243 (N_243,In_689,In_621);
nand U244 (N_244,In_141,In_874);
and U245 (N_245,In_19,In_711);
and U246 (N_246,In_273,In_630);
and U247 (N_247,In_63,In_431);
nor U248 (N_248,In_13,In_339);
nand U249 (N_249,In_573,In_332);
and U250 (N_250,In_309,In_444);
nor U251 (N_251,In_306,In_560);
nor U252 (N_252,In_357,In_8);
nor U253 (N_253,In_919,In_44);
nand U254 (N_254,In_635,In_319);
and U255 (N_255,In_259,In_469);
nor U256 (N_256,In_834,In_898);
nand U257 (N_257,In_729,In_217);
nor U258 (N_258,In_484,In_743);
nor U259 (N_259,In_752,In_395);
nand U260 (N_260,In_707,In_248);
nand U261 (N_261,In_622,In_78);
xor U262 (N_262,In_849,In_881);
nand U263 (N_263,In_842,In_862);
nor U264 (N_264,In_661,In_542);
nor U265 (N_265,In_113,In_750);
and U266 (N_266,In_730,In_561);
nor U267 (N_267,In_364,In_995);
nand U268 (N_268,In_749,In_920);
nor U269 (N_269,In_240,In_294);
and U270 (N_270,In_614,In_608);
and U271 (N_271,In_808,In_800);
xnor U272 (N_272,In_241,In_957);
xor U273 (N_273,In_742,In_591);
nor U274 (N_274,In_327,In_111);
nand U275 (N_275,In_935,In_677);
nor U276 (N_276,In_302,In_539);
nor U277 (N_277,In_57,In_747);
nor U278 (N_278,In_774,In_144);
and U279 (N_279,In_450,In_154);
and U280 (N_280,In_490,In_745);
and U281 (N_281,In_619,In_390);
and U282 (N_282,In_437,In_134);
and U283 (N_283,In_769,In_592);
nand U284 (N_284,In_126,In_375);
or U285 (N_285,In_869,In_642);
or U286 (N_286,In_518,In_192);
nor U287 (N_287,In_252,In_679);
and U288 (N_288,In_264,In_879);
nand U289 (N_289,In_979,In_167);
xnor U290 (N_290,In_797,In_860);
nand U291 (N_291,In_804,In_305);
or U292 (N_292,In_41,In_717);
nand U293 (N_293,In_515,In_413);
or U294 (N_294,In_421,In_754);
nor U295 (N_295,In_787,In_504);
xnor U296 (N_296,In_648,In_934);
or U297 (N_297,In_216,In_366);
or U298 (N_298,In_851,In_155);
or U299 (N_299,In_966,In_163);
nand U300 (N_300,In_423,In_529);
xor U301 (N_301,In_34,In_924);
nand U302 (N_302,In_90,In_760);
nor U303 (N_303,In_465,In_51);
or U304 (N_304,In_830,In_998);
nand U305 (N_305,In_54,In_952);
nand U306 (N_306,In_173,In_70);
nor U307 (N_307,In_558,In_996);
or U308 (N_308,In_624,In_818);
and U309 (N_309,In_96,In_659);
or U310 (N_310,In_436,In_239);
or U311 (N_311,In_66,In_600);
xor U312 (N_312,In_973,In_541);
or U313 (N_313,In_867,In_179);
xor U314 (N_314,In_885,In_45);
and U315 (N_315,In_493,In_670);
or U316 (N_316,In_123,In_374);
nor U317 (N_317,In_891,In_403);
and U318 (N_318,In_494,In_936);
and U319 (N_319,In_499,In_563);
or U320 (N_320,In_17,In_397);
and U321 (N_321,In_202,In_837);
nand U322 (N_322,In_908,In_161);
or U323 (N_323,In_243,In_52);
or U324 (N_324,In_950,In_734);
nor U325 (N_325,In_736,In_564);
or U326 (N_326,In_349,In_687);
nor U327 (N_327,In_416,In_521);
xor U328 (N_328,In_95,In_801);
nand U329 (N_329,In_221,In_233);
and U330 (N_330,In_803,In_586);
or U331 (N_331,In_193,In_384);
nand U332 (N_332,In_625,In_53);
nor U333 (N_333,In_222,In_448);
nand U334 (N_334,In_280,In_9);
xor U335 (N_335,In_639,In_303);
nor U336 (N_336,In_362,In_649);
and U337 (N_337,In_2,In_605);
xnor U338 (N_338,In_301,In_718);
nor U339 (N_339,In_39,In_668);
and U340 (N_340,In_678,In_756);
xnor U341 (N_341,In_883,In_142);
nand U342 (N_342,In_404,In_257);
or U343 (N_343,In_978,In_42);
xnor U344 (N_344,In_184,In_637);
or U345 (N_345,In_139,In_360);
and U346 (N_346,In_495,In_247);
and U347 (N_347,In_555,In_984);
and U348 (N_348,In_807,In_428);
nand U349 (N_349,In_48,In_171);
or U350 (N_350,In_116,In_246);
xor U351 (N_351,In_253,In_598);
xor U352 (N_352,In_311,In_968);
xor U353 (N_353,In_31,In_930);
or U354 (N_354,In_611,In_156);
or U355 (N_355,In_958,In_843);
nand U356 (N_356,In_410,In_10);
and U357 (N_357,In_125,In_647);
and U358 (N_358,In_32,In_105);
nor U359 (N_359,In_82,In_166);
nand U360 (N_360,In_823,In_487);
xnor U361 (N_361,In_376,In_535);
and U362 (N_362,In_833,In_982);
xnor U363 (N_363,In_660,In_27);
and U364 (N_364,In_971,In_201);
or U365 (N_365,In_271,In_791);
nor U366 (N_366,In_459,In_433);
nand U367 (N_367,In_852,In_907);
nand U368 (N_368,In_706,In_312);
or U369 (N_369,In_981,In_261);
xor U370 (N_370,In_391,In_857);
xnor U371 (N_371,In_177,In_914);
nor U372 (N_372,In_528,In_517);
nor U373 (N_373,In_508,In_386);
nand U374 (N_374,In_345,In_463);
or U375 (N_375,In_419,In_268);
nand U376 (N_376,In_151,In_581);
nand U377 (N_377,In_571,In_14);
xor U378 (N_378,In_148,In_559);
nor U379 (N_379,In_604,In_913);
or U380 (N_380,In_552,In_46);
nand U381 (N_381,In_351,In_509);
nor U382 (N_382,In_137,In_912);
xor U383 (N_383,In_169,In_64);
or U384 (N_384,In_347,In_940);
and U385 (N_385,In_931,In_675);
and U386 (N_386,In_861,In_190);
nor U387 (N_387,In_612,In_550);
or U388 (N_388,In_263,In_127);
nand U389 (N_389,In_182,In_575);
and U390 (N_390,In_895,In_405);
nand U391 (N_391,In_455,In_618);
nand U392 (N_392,In_164,In_887);
and U393 (N_393,In_128,In_453);
xnor U394 (N_394,In_40,In_526);
and U395 (N_395,In_770,In_970);
or U396 (N_396,In_458,In_81);
nor U397 (N_397,In_684,In_434);
or U398 (N_398,In_939,In_938);
or U399 (N_399,In_249,In_816);
xor U400 (N_400,In_820,In_963);
nand U401 (N_401,In_941,In_942);
or U402 (N_402,In_817,In_260);
nor U403 (N_403,In_696,In_764);
nor U404 (N_404,In_576,In_651);
or U405 (N_405,In_378,In_580);
xor U406 (N_406,In_132,In_337);
nand U407 (N_407,In_500,In_836);
and U408 (N_408,In_295,In_373);
or U409 (N_409,In_394,In_641);
xnor U410 (N_410,In_927,In_235);
xor U411 (N_411,In_77,In_951);
and U412 (N_412,In_335,In_932);
xor U413 (N_413,In_980,In_937);
and U414 (N_414,In_114,In_354);
and U415 (N_415,In_310,In_475);
and U416 (N_416,In_331,In_610);
xor U417 (N_417,In_796,In_102);
or U418 (N_418,In_377,In_62);
xor U419 (N_419,In_282,In_272);
nand U420 (N_420,In_850,In_793);
nor U421 (N_421,In_37,In_99);
and U422 (N_422,In_91,In_565);
and U423 (N_423,In_673,In_28);
and U424 (N_424,In_88,In_197);
nand U425 (N_425,In_65,In_371);
or U426 (N_426,In_882,In_522);
or U427 (N_427,In_819,In_721);
and U428 (N_428,In_20,In_954);
xnor U429 (N_429,In_258,In_400);
nor U430 (N_430,In_36,In_289);
nand U431 (N_431,In_643,In_805);
or U432 (N_432,In_652,In_392);
or U433 (N_433,In_732,In_946);
and U434 (N_434,In_187,In_933);
xnor U435 (N_435,In_480,In_333);
or U436 (N_436,In_279,In_686);
and U437 (N_437,In_638,In_606);
and U438 (N_438,In_342,In_928);
nor U439 (N_439,In_735,In_452);
and U440 (N_440,In_588,In_496);
or U441 (N_441,In_274,In_92);
nor U442 (N_442,In_691,In_739);
or U443 (N_443,In_119,In_406);
xor U444 (N_444,In_910,In_231);
or U445 (N_445,In_363,In_977);
nor U446 (N_446,In_12,In_775);
nor U447 (N_447,In_368,In_422);
or U448 (N_448,In_944,In_242);
nor U449 (N_449,In_1,In_73);
nand U450 (N_450,In_501,In_188);
nand U451 (N_451,In_471,In_341);
nor U452 (N_452,In_701,In_506);
nand U453 (N_453,In_477,In_853);
or U454 (N_454,In_964,In_975);
and U455 (N_455,In_186,In_245);
and U456 (N_456,In_441,In_523);
or U457 (N_457,In_582,In_915);
and U458 (N_458,In_488,In_856);
xor U459 (N_459,In_589,In_814);
nor U460 (N_460,In_688,In_318);
or U461 (N_461,In_755,In_117);
or U462 (N_462,In_293,In_781);
nand U463 (N_463,In_118,In_888);
xnor U464 (N_464,In_519,In_474);
xnor U465 (N_465,In_845,In_511);
nor U466 (N_466,In_909,In_59);
and U467 (N_467,In_3,In_228);
xor U468 (N_468,In_420,In_146);
nand U469 (N_469,In_737,In_230);
nand U470 (N_470,In_492,In_75);
and U471 (N_471,In_344,In_716);
xnor U472 (N_472,In_313,In_396);
nand U473 (N_473,In_284,In_640);
nand U474 (N_474,In_16,In_864);
and U475 (N_475,In_136,In_872);
nand U476 (N_476,In_603,In_379);
nor U477 (N_477,In_424,In_956);
or U478 (N_478,In_185,In_594);
xnor U479 (N_479,In_94,In_765);
nor U480 (N_480,In_794,In_385);
or U481 (N_481,In_967,In_350);
or U482 (N_482,In_945,In_922);
or U483 (N_483,In_628,In_545);
and U484 (N_484,In_683,In_323);
xnor U485 (N_485,In_538,In_976);
or U486 (N_486,In_534,In_585);
nor U487 (N_487,In_285,In_811);
or U488 (N_488,In_203,In_502);
and U489 (N_489,In_759,In_897);
nor U490 (N_490,In_447,In_195);
nand U491 (N_491,In_513,In_383);
nor U492 (N_492,In_191,In_674);
xor U493 (N_493,In_232,In_902);
and U494 (N_494,In_482,In_644);
or U495 (N_495,In_904,In_841);
and U496 (N_496,In_108,In_620);
nor U497 (N_497,In_889,In_991);
or U498 (N_498,In_772,In_532);
or U499 (N_499,In_510,In_525);
nor U500 (N_500,N_75,N_62);
nand U501 (N_501,N_83,N_482);
xnor U502 (N_502,N_76,N_361);
and U503 (N_503,N_46,N_403);
nor U504 (N_504,N_344,N_201);
xnor U505 (N_505,N_276,N_26);
nand U506 (N_506,N_396,N_398);
and U507 (N_507,N_366,N_326);
and U508 (N_508,N_7,N_16);
xnor U509 (N_509,N_102,N_212);
nor U510 (N_510,N_321,N_112);
nand U511 (N_511,N_110,N_134);
nor U512 (N_512,N_91,N_342);
xor U513 (N_513,N_185,N_178);
nand U514 (N_514,N_260,N_8);
xor U515 (N_515,N_303,N_343);
nand U516 (N_516,N_136,N_52);
or U517 (N_517,N_429,N_411);
xor U518 (N_518,N_200,N_419);
nor U519 (N_519,N_440,N_17);
and U520 (N_520,N_473,N_117);
xor U521 (N_521,N_494,N_157);
nor U522 (N_522,N_160,N_35);
nand U523 (N_523,N_446,N_277);
xnor U524 (N_524,N_124,N_44);
or U525 (N_525,N_232,N_427);
xor U526 (N_526,N_229,N_324);
xor U527 (N_527,N_376,N_196);
or U528 (N_528,N_262,N_491);
and U529 (N_529,N_240,N_489);
and U530 (N_530,N_441,N_413);
xnor U531 (N_531,N_54,N_351);
and U532 (N_532,N_292,N_369);
and U533 (N_533,N_152,N_51);
and U534 (N_534,N_367,N_392);
nand U535 (N_535,N_358,N_363);
and U536 (N_536,N_356,N_364);
nand U537 (N_537,N_123,N_250);
nor U538 (N_538,N_132,N_495);
xnor U539 (N_539,N_158,N_450);
nand U540 (N_540,N_488,N_273);
nor U541 (N_541,N_225,N_312);
xnor U542 (N_542,N_439,N_288);
and U543 (N_543,N_255,N_470);
or U544 (N_544,N_352,N_395);
nand U545 (N_545,N_252,N_498);
nand U546 (N_546,N_202,N_329);
nand U547 (N_547,N_426,N_345);
nor U548 (N_548,N_462,N_453);
and U549 (N_549,N_221,N_448);
nor U550 (N_550,N_80,N_12);
or U551 (N_551,N_25,N_92);
xor U552 (N_552,N_301,N_454);
or U553 (N_553,N_140,N_139);
xor U554 (N_554,N_320,N_207);
and U555 (N_555,N_438,N_71);
nor U556 (N_556,N_49,N_173);
and U557 (N_557,N_332,N_341);
nand U558 (N_558,N_282,N_267);
and U559 (N_559,N_218,N_258);
xnor U560 (N_560,N_99,N_302);
or U561 (N_561,N_349,N_228);
and U562 (N_562,N_456,N_327);
nand U563 (N_563,N_129,N_161);
xor U564 (N_564,N_304,N_457);
or U565 (N_565,N_235,N_325);
nand U566 (N_566,N_348,N_154);
nor U567 (N_567,N_298,N_314);
nor U568 (N_568,N_111,N_472);
xor U569 (N_569,N_407,N_29);
and U570 (N_570,N_399,N_391);
or U571 (N_571,N_30,N_318);
xor U572 (N_572,N_50,N_170);
xnor U573 (N_573,N_108,N_121);
nand U574 (N_574,N_171,N_245);
and U575 (N_575,N_452,N_257);
and U576 (N_576,N_346,N_45);
and U577 (N_577,N_82,N_233);
nand U578 (N_578,N_469,N_291);
xor U579 (N_579,N_217,N_485);
or U580 (N_580,N_434,N_353);
nand U581 (N_581,N_184,N_3);
and U582 (N_582,N_143,N_425);
nand U583 (N_583,N_116,N_179);
nand U584 (N_584,N_477,N_105);
or U585 (N_585,N_307,N_204);
xnor U586 (N_586,N_4,N_360);
or U587 (N_587,N_219,N_23);
nor U588 (N_588,N_86,N_85);
nor U589 (N_589,N_265,N_382);
and U590 (N_590,N_97,N_374);
nor U591 (N_591,N_96,N_115);
and U592 (N_592,N_34,N_205);
xor U593 (N_593,N_404,N_194);
and U594 (N_594,N_445,N_471);
nand U595 (N_595,N_107,N_84);
and U596 (N_596,N_79,N_417);
nand U597 (N_597,N_406,N_131);
xor U598 (N_598,N_174,N_64);
and U599 (N_599,N_15,N_19);
and U600 (N_600,N_493,N_21);
or U601 (N_601,N_141,N_101);
and U602 (N_602,N_78,N_31);
and U603 (N_603,N_58,N_316);
and U604 (N_604,N_447,N_295);
and U605 (N_605,N_283,N_135);
nand U606 (N_606,N_106,N_323);
and U607 (N_607,N_336,N_10);
xor U608 (N_608,N_371,N_313);
xor U609 (N_609,N_133,N_216);
and U610 (N_610,N_32,N_284);
and U611 (N_611,N_241,N_74);
xnor U612 (N_612,N_213,N_168);
and U613 (N_613,N_0,N_455);
xnor U614 (N_614,N_43,N_490);
and U615 (N_615,N_113,N_39);
or U616 (N_616,N_224,N_146);
or U617 (N_617,N_210,N_308);
and U618 (N_618,N_259,N_22);
nand U619 (N_619,N_460,N_188);
xor U620 (N_620,N_333,N_211);
or U621 (N_621,N_95,N_209);
nor U622 (N_622,N_195,N_484);
nor U623 (N_623,N_414,N_145);
and U624 (N_624,N_128,N_300);
nor U625 (N_625,N_169,N_381);
nor U626 (N_626,N_67,N_483);
or U627 (N_627,N_256,N_408);
xor U628 (N_628,N_56,N_165);
nor U629 (N_629,N_226,N_465);
nand U630 (N_630,N_389,N_442);
xor U631 (N_631,N_127,N_377);
xor U632 (N_632,N_66,N_68);
nor U633 (N_633,N_286,N_280);
nor U634 (N_634,N_443,N_192);
or U635 (N_635,N_272,N_42);
nand U636 (N_636,N_478,N_476);
nor U637 (N_637,N_474,N_148);
and U638 (N_638,N_335,N_1);
nor U639 (N_639,N_6,N_458);
and U640 (N_640,N_230,N_350);
or U641 (N_641,N_285,N_379);
or U642 (N_642,N_13,N_357);
or U643 (N_643,N_278,N_93);
nor U644 (N_644,N_370,N_311);
nand U645 (N_645,N_5,N_290);
nand U646 (N_646,N_130,N_415);
nor U647 (N_647,N_365,N_150);
xor U648 (N_648,N_299,N_138);
nor U649 (N_649,N_479,N_215);
and U650 (N_650,N_263,N_334);
nand U651 (N_651,N_53,N_94);
or U652 (N_652,N_191,N_14);
or U653 (N_653,N_147,N_492);
and U654 (N_654,N_317,N_40);
or U655 (N_655,N_499,N_422);
nor U656 (N_656,N_187,N_223);
xnor U657 (N_657,N_144,N_340);
xnor U658 (N_658,N_387,N_36);
and U659 (N_659,N_467,N_88);
nand U660 (N_660,N_430,N_373);
nand U661 (N_661,N_47,N_338);
or U662 (N_662,N_297,N_281);
or U663 (N_663,N_261,N_61);
nor U664 (N_664,N_459,N_461);
or U665 (N_665,N_444,N_163);
xnor U666 (N_666,N_378,N_397);
xor U667 (N_667,N_423,N_151);
xor U668 (N_668,N_322,N_436);
nor U669 (N_669,N_72,N_176);
nand U670 (N_670,N_264,N_103);
xnor U671 (N_671,N_162,N_149);
nor U672 (N_672,N_98,N_435);
nor U673 (N_673,N_354,N_331);
nand U674 (N_674,N_339,N_186);
nor U675 (N_675,N_475,N_247);
nor U676 (N_676,N_28,N_11);
nor U677 (N_677,N_87,N_294);
xnor U678 (N_678,N_287,N_388);
and U679 (N_679,N_220,N_412);
and U680 (N_680,N_198,N_77);
and U681 (N_681,N_305,N_362);
nor U682 (N_682,N_208,N_27);
xnor U683 (N_683,N_109,N_69);
xnor U684 (N_684,N_401,N_203);
and U685 (N_685,N_310,N_497);
or U686 (N_686,N_20,N_296);
and U687 (N_687,N_222,N_463);
xnor U688 (N_688,N_437,N_409);
or U689 (N_689,N_167,N_432);
nor U690 (N_690,N_253,N_380);
nand U691 (N_691,N_183,N_268);
or U692 (N_692,N_120,N_393);
nor U693 (N_693,N_182,N_237);
nand U694 (N_694,N_418,N_315);
xnor U695 (N_695,N_114,N_60);
nand U696 (N_696,N_486,N_306);
xnor U697 (N_697,N_100,N_416);
or U698 (N_698,N_122,N_420);
xor U699 (N_699,N_246,N_33);
nor U700 (N_700,N_464,N_37);
xor U701 (N_701,N_421,N_9);
and U702 (N_702,N_231,N_275);
nand U703 (N_703,N_289,N_55);
and U704 (N_704,N_355,N_159);
and U705 (N_705,N_243,N_251);
nand U706 (N_706,N_63,N_372);
xor U707 (N_707,N_164,N_118);
and U708 (N_708,N_70,N_81);
nand U709 (N_709,N_394,N_359);
or U710 (N_710,N_496,N_90);
xnor U711 (N_711,N_309,N_206);
nor U712 (N_712,N_18,N_189);
xnor U713 (N_713,N_270,N_38);
nor U714 (N_714,N_384,N_271);
nor U715 (N_715,N_238,N_48);
or U716 (N_716,N_156,N_190);
nand U717 (N_717,N_73,N_274);
or U718 (N_718,N_125,N_244);
xor U719 (N_719,N_126,N_59);
xnor U720 (N_720,N_180,N_254);
nand U721 (N_721,N_424,N_368);
or U722 (N_722,N_172,N_428);
xor U723 (N_723,N_197,N_2);
or U724 (N_724,N_269,N_293);
nor U725 (N_725,N_375,N_175);
nand U726 (N_726,N_239,N_337);
nand U727 (N_727,N_347,N_234);
nand U728 (N_728,N_431,N_249);
nand U729 (N_729,N_89,N_400);
nor U730 (N_730,N_155,N_402);
nor U731 (N_731,N_390,N_166);
nor U732 (N_732,N_104,N_386);
xor U733 (N_733,N_433,N_279);
xnor U734 (N_734,N_248,N_481);
and U735 (N_735,N_383,N_242);
and U736 (N_736,N_65,N_24);
and U737 (N_737,N_449,N_487);
nor U738 (N_738,N_142,N_410);
and U739 (N_739,N_266,N_451);
and U740 (N_740,N_193,N_468);
or U741 (N_741,N_328,N_480);
nor U742 (N_742,N_153,N_319);
and U743 (N_743,N_137,N_405);
and U744 (N_744,N_57,N_199);
and U745 (N_745,N_177,N_119);
and U746 (N_746,N_385,N_330);
nor U747 (N_747,N_214,N_236);
nor U748 (N_748,N_181,N_466);
nand U749 (N_749,N_41,N_227);
xor U750 (N_750,N_246,N_312);
or U751 (N_751,N_235,N_266);
nand U752 (N_752,N_239,N_278);
nand U753 (N_753,N_186,N_359);
xnor U754 (N_754,N_362,N_432);
nand U755 (N_755,N_291,N_182);
xor U756 (N_756,N_486,N_11);
xor U757 (N_757,N_32,N_154);
xnor U758 (N_758,N_434,N_339);
and U759 (N_759,N_13,N_217);
nor U760 (N_760,N_352,N_148);
or U761 (N_761,N_440,N_56);
nor U762 (N_762,N_135,N_291);
nand U763 (N_763,N_435,N_453);
xor U764 (N_764,N_344,N_385);
nand U765 (N_765,N_103,N_294);
or U766 (N_766,N_21,N_309);
nand U767 (N_767,N_148,N_451);
xor U768 (N_768,N_112,N_262);
nand U769 (N_769,N_256,N_432);
and U770 (N_770,N_382,N_164);
nand U771 (N_771,N_134,N_74);
xnor U772 (N_772,N_108,N_356);
and U773 (N_773,N_54,N_425);
and U774 (N_774,N_330,N_298);
nor U775 (N_775,N_40,N_137);
nand U776 (N_776,N_96,N_389);
nor U777 (N_777,N_312,N_240);
nand U778 (N_778,N_10,N_473);
nor U779 (N_779,N_98,N_429);
or U780 (N_780,N_169,N_288);
and U781 (N_781,N_482,N_283);
nor U782 (N_782,N_122,N_380);
nand U783 (N_783,N_498,N_157);
nor U784 (N_784,N_73,N_20);
nand U785 (N_785,N_214,N_273);
nor U786 (N_786,N_258,N_92);
nor U787 (N_787,N_272,N_176);
xor U788 (N_788,N_496,N_322);
xnor U789 (N_789,N_376,N_110);
nor U790 (N_790,N_118,N_326);
xor U791 (N_791,N_416,N_191);
xor U792 (N_792,N_113,N_173);
and U793 (N_793,N_87,N_90);
nor U794 (N_794,N_492,N_432);
and U795 (N_795,N_377,N_267);
nor U796 (N_796,N_79,N_2);
or U797 (N_797,N_83,N_406);
and U798 (N_798,N_35,N_458);
or U799 (N_799,N_115,N_25);
nand U800 (N_800,N_198,N_74);
xnor U801 (N_801,N_11,N_173);
nand U802 (N_802,N_440,N_24);
and U803 (N_803,N_306,N_368);
nand U804 (N_804,N_146,N_345);
nand U805 (N_805,N_345,N_7);
or U806 (N_806,N_168,N_445);
nor U807 (N_807,N_355,N_172);
nand U808 (N_808,N_61,N_177);
xor U809 (N_809,N_134,N_104);
and U810 (N_810,N_318,N_57);
xnor U811 (N_811,N_368,N_270);
nand U812 (N_812,N_153,N_82);
xnor U813 (N_813,N_242,N_399);
and U814 (N_814,N_101,N_428);
nor U815 (N_815,N_276,N_140);
or U816 (N_816,N_186,N_234);
or U817 (N_817,N_497,N_320);
xor U818 (N_818,N_113,N_219);
xor U819 (N_819,N_352,N_24);
or U820 (N_820,N_368,N_396);
xor U821 (N_821,N_273,N_203);
nor U822 (N_822,N_76,N_478);
or U823 (N_823,N_430,N_230);
nand U824 (N_824,N_173,N_397);
xor U825 (N_825,N_329,N_159);
xnor U826 (N_826,N_195,N_421);
xor U827 (N_827,N_173,N_156);
or U828 (N_828,N_398,N_340);
xnor U829 (N_829,N_180,N_272);
nor U830 (N_830,N_197,N_163);
nor U831 (N_831,N_366,N_299);
xnor U832 (N_832,N_363,N_271);
and U833 (N_833,N_437,N_476);
nor U834 (N_834,N_480,N_25);
nor U835 (N_835,N_349,N_30);
and U836 (N_836,N_145,N_100);
xor U837 (N_837,N_226,N_71);
and U838 (N_838,N_63,N_329);
xor U839 (N_839,N_33,N_372);
xnor U840 (N_840,N_115,N_372);
nor U841 (N_841,N_210,N_1);
xor U842 (N_842,N_0,N_311);
xor U843 (N_843,N_361,N_276);
nor U844 (N_844,N_25,N_159);
xnor U845 (N_845,N_228,N_191);
nand U846 (N_846,N_388,N_125);
nor U847 (N_847,N_406,N_275);
nor U848 (N_848,N_128,N_119);
nand U849 (N_849,N_265,N_91);
xor U850 (N_850,N_134,N_337);
xnor U851 (N_851,N_207,N_211);
or U852 (N_852,N_181,N_277);
and U853 (N_853,N_234,N_380);
and U854 (N_854,N_367,N_3);
or U855 (N_855,N_249,N_330);
xnor U856 (N_856,N_21,N_244);
and U857 (N_857,N_136,N_399);
xor U858 (N_858,N_133,N_424);
nor U859 (N_859,N_365,N_202);
nor U860 (N_860,N_491,N_270);
xnor U861 (N_861,N_98,N_418);
nand U862 (N_862,N_25,N_43);
xor U863 (N_863,N_254,N_46);
and U864 (N_864,N_13,N_412);
nor U865 (N_865,N_197,N_418);
xnor U866 (N_866,N_191,N_73);
or U867 (N_867,N_244,N_97);
xnor U868 (N_868,N_271,N_401);
and U869 (N_869,N_100,N_334);
or U870 (N_870,N_353,N_455);
nand U871 (N_871,N_64,N_24);
xor U872 (N_872,N_12,N_208);
nor U873 (N_873,N_97,N_373);
or U874 (N_874,N_174,N_373);
and U875 (N_875,N_120,N_428);
nand U876 (N_876,N_428,N_308);
xor U877 (N_877,N_429,N_372);
and U878 (N_878,N_376,N_149);
nor U879 (N_879,N_113,N_79);
and U880 (N_880,N_413,N_341);
or U881 (N_881,N_448,N_167);
nand U882 (N_882,N_74,N_223);
or U883 (N_883,N_311,N_18);
and U884 (N_884,N_24,N_146);
nand U885 (N_885,N_423,N_342);
and U886 (N_886,N_107,N_218);
nand U887 (N_887,N_353,N_390);
and U888 (N_888,N_351,N_256);
xnor U889 (N_889,N_443,N_178);
xnor U890 (N_890,N_313,N_355);
xor U891 (N_891,N_393,N_360);
nand U892 (N_892,N_154,N_222);
xor U893 (N_893,N_288,N_389);
and U894 (N_894,N_153,N_353);
and U895 (N_895,N_79,N_115);
or U896 (N_896,N_345,N_92);
xor U897 (N_897,N_45,N_305);
and U898 (N_898,N_437,N_387);
xor U899 (N_899,N_343,N_128);
nand U900 (N_900,N_15,N_330);
or U901 (N_901,N_60,N_358);
or U902 (N_902,N_186,N_281);
and U903 (N_903,N_233,N_37);
or U904 (N_904,N_323,N_377);
nor U905 (N_905,N_200,N_344);
xor U906 (N_906,N_383,N_82);
nand U907 (N_907,N_297,N_29);
or U908 (N_908,N_369,N_164);
nand U909 (N_909,N_210,N_75);
and U910 (N_910,N_322,N_443);
xnor U911 (N_911,N_109,N_381);
nor U912 (N_912,N_278,N_336);
nor U913 (N_913,N_379,N_450);
xor U914 (N_914,N_343,N_404);
or U915 (N_915,N_295,N_328);
and U916 (N_916,N_90,N_81);
nand U917 (N_917,N_38,N_376);
nand U918 (N_918,N_311,N_420);
nand U919 (N_919,N_119,N_158);
and U920 (N_920,N_381,N_490);
xnor U921 (N_921,N_456,N_66);
nor U922 (N_922,N_400,N_191);
and U923 (N_923,N_429,N_53);
nand U924 (N_924,N_454,N_132);
and U925 (N_925,N_448,N_227);
or U926 (N_926,N_369,N_56);
nand U927 (N_927,N_403,N_38);
and U928 (N_928,N_31,N_440);
nor U929 (N_929,N_416,N_493);
xnor U930 (N_930,N_346,N_189);
or U931 (N_931,N_289,N_441);
and U932 (N_932,N_292,N_222);
nand U933 (N_933,N_447,N_453);
xnor U934 (N_934,N_411,N_145);
and U935 (N_935,N_329,N_354);
nand U936 (N_936,N_18,N_378);
and U937 (N_937,N_218,N_181);
nor U938 (N_938,N_236,N_279);
nor U939 (N_939,N_320,N_352);
nor U940 (N_940,N_361,N_443);
nor U941 (N_941,N_493,N_52);
and U942 (N_942,N_30,N_259);
xnor U943 (N_943,N_53,N_258);
xor U944 (N_944,N_420,N_315);
or U945 (N_945,N_220,N_7);
or U946 (N_946,N_384,N_141);
or U947 (N_947,N_109,N_181);
or U948 (N_948,N_365,N_275);
and U949 (N_949,N_461,N_369);
nand U950 (N_950,N_309,N_398);
or U951 (N_951,N_277,N_88);
nor U952 (N_952,N_418,N_118);
and U953 (N_953,N_374,N_316);
xor U954 (N_954,N_308,N_344);
nand U955 (N_955,N_461,N_427);
nor U956 (N_956,N_200,N_253);
nor U957 (N_957,N_20,N_286);
and U958 (N_958,N_221,N_449);
nor U959 (N_959,N_328,N_492);
or U960 (N_960,N_316,N_21);
nand U961 (N_961,N_76,N_264);
xnor U962 (N_962,N_361,N_191);
nand U963 (N_963,N_425,N_103);
nor U964 (N_964,N_207,N_265);
nand U965 (N_965,N_344,N_212);
nor U966 (N_966,N_188,N_189);
nor U967 (N_967,N_290,N_220);
and U968 (N_968,N_331,N_426);
nor U969 (N_969,N_295,N_321);
nand U970 (N_970,N_442,N_422);
and U971 (N_971,N_41,N_370);
xor U972 (N_972,N_139,N_406);
and U973 (N_973,N_81,N_379);
or U974 (N_974,N_384,N_359);
xnor U975 (N_975,N_341,N_462);
nor U976 (N_976,N_133,N_335);
nor U977 (N_977,N_320,N_461);
nor U978 (N_978,N_140,N_300);
nand U979 (N_979,N_130,N_47);
and U980 (N_980,N_92,N_418);
and U981 (N_981,N_265,N_485);
nand U982 (N_982,N_336,N_442);
nor U983 (N_983,N_496,N_143);
or U984 (N_984,N_249,N_361);
nand U985 (N_985,N_490,N_1);
nand U986 (N_986,N_189,N_369);
and U987 (N_987,N_449,N_361);
xnor U988 (N_988,N_269,N_255);
nand U989 (N_989,N_73,N_376);
nand U990 (N_990,N_377,N_131);
xor U991 (N_991,N_322,N_31);
or U992 (N_992,N_105,N_75);
and U993 (N_993,N_134,N_76);
and U994 (N_994,N_419,N_441);
or U995 (N_995,N_278,N_185);
nand U996 (N_996,N_470,N_252);
xor U997 (N_997,N_44,N_412);
and U998 (N_998,N_163,N_83);
xor U999 (N_999,N_465,N_86);
or U1000 (N_1000,N_516,N_597);
nand U1001 (N_1001,N_654,N_792);
and U1002 (N_1002,N_935,N_598);
and U1003 (N_1003,N_615,N_876);
xor U1004 (N_1004,N_774,N_582);
xor U1005 (N_1005,N_624,N_603);
or U1006 (N_1006,N_874,N_656);
or U1007 (N_1007,N_943,N_873);
xor U1008 (N_1008,N_541,N_613);
xnor U1009 (N_1009,N_545,N_894);
or U1010 (N_1010,N_675,N_709);
or U1011 (N_1011,N_665,N_992);
or U1012 (N_1012,N_523,N_795);
nor U1013 (N_1013,N_849,N_946);
nand U1014 (N_1014,N_825,N_672);
nand U1015 (N_1015,N_855,N_738);
or U1016 (N_1016,N_852,N_560);
xnor U1017 (N_1017,N_923,N_682);
nor U1018 (N_1018,N_879,N_844);
nand U1019 (N_1019,N_890,N_776);
nor U1020 (N_1020,N_594,N_911);
nand U1021 (N_1021,N_987,N_956);
nor U1022 (N_1022,N_532,N_700);
xor U1023 (N_1023,N_962,N_881);
or U1024 (N_1024,N_534,N_864);
or U1025 (N_1025,N_637,N_659);
nor U1026 (N_1026,N_801,N_674);
nand U1027 (N_1027,N_889,N_780);
and U1028 (N_1028,N_908,N_918);
nand U1029 (N_1029,N_737,N_689);
xnor U1030 (N_1030,N_998,N_677);
nor U1031 (N_1031,N_954,N_952);
nand U1032 (N_1032,N_745,N_566);
nor U1033 (N_1033,N_818,N_501);
nand U1034 (N_1034,N_502,N_642);
and U1035 (N_1035,N_891,N_932);
nor U1036 (N_1036,N_939,N_683);
xor U1037 (N_1037,N_673,N_607);
xor U1038 (N_1038,N_666,N_871);
and U1039 (N_1039,N_937,N_590);
nor U1040 (N_1040,N_551,N_726);
xor U1041 (N_1041,N_870,N_629);
and U1042 (N_1042,N_805,N_733);
or U1043 (N_1043,N_605,N_741);
or U1044 (N_1044,N_627,N_841);
or U1045 (N_1045,N_503,N_595);
nor U1046 (N_1046,N_620,N_657);
nor U1047 (N_1047,N_899,N_611);
or U1048 (N_1048,N_513,N_730);
xnor U1049 (N_1049,N_508,N_797);
nand U1050 (N_1050,N_925,N_647);
and U1051 (N_1051,N_972,N_616);
and U1052 (N_1052,N_802,N_658);
xor U1053 (N_1053,N_989,N_552);
and U1054 (N_1054,N_866,N_628);
nor U1055 (N_1055,N_951,N_934);
and U1056 (N_1056,N_589,N_839);
nand U1057 (N_1057,N_751,N_717);
and U1058 (N_1058,N_572,N_617);
nand U1059 (N_1059,N_840,N_707);
and U1060 (N_1060,N_978,N_878);
nor U1061 (N_1061,N_696,N_555);
xnor U1062 (N_1062,N_847,N_524);
nand U1063 (N_1063,N_980,N_526);
xnor U1064 (N_1064,N_529,N_718);
nand U1065 (N_1065,N_569,N_655);
or U1066 (N_1066,N_591,N_814);
or U1067 (N_1067,N_957,N_808);
xor U1068 (N_1068,N_568,N_875);
nor U1069 (N_1069,N_900,N_710);
or U1070 (N_1070,N_688,N_521);
xor U1071 (N_1071,N_893,N_650);
or U1072 (N_1072,N_888,N_817);
nand U1073 (N_1073,N_877,N_820);
nor U1074 (N_1074,N_942,N_967);
nor U1075 (N_1075,N_563,N_606);
nor U1076 (N_1076,N_662,N_760);
xor U1077 (N_1077,N_693,N_621);
nor U1078 (N_1078,N_511,N_567);
and U1079 (N_1079,N_869,N_544);
nand U1080 (N_1080,N_610,N_515);
nand U1081 (N_1081,N_525,N_858);
nor U1082 (N_1082,N_921,N_885);
xor U1083 (N_1083,N_507,N_807);
nor U1084 (N_1084,N_638,N_625);
and U1085 (N_1085,N_732,N_540);
nand U1086 (N_1086,N_531,N_542);
nand U1087 (N_1087,N_680,N_549);
nor U1088 (N_1088,N_764,N_559);
nor U1089 (N_1089,N_846,N_781);
and U1090 (N_1090,N_955,N_931);
or U1091 (N_1091,N_828,N_916);
nor U1092 (N_1092,N_699,N_974);
and U1093 (N_1093,N_768,N_588);
or U1094 (N_1094,N_853,N_915);
nand U1095 (N_1095,N_695,N_671);
or U1096 (N_1096,N_772,N_535);
or U1097 (N_1097,N_720,N_822);
and U1098 (N_1098,N_810,N_635);
nor U1099 (N_1099,N_639,N_510);
nor U1100 (N_1100,N_993,N_714);
or U1101 (N_1101,N_796,N_653);
xnor U1102 (N_1102,N_632,N_593);
xor U1103 (N_1103,N_547,N_984);
nor U1104 (N_1104,N_819,N_773);
xnor U1105 (N_1105,N_652,N_729);
nand U1106 (N_1106,N_880,N_767);
nand U1107 (N_1107,N_948,N_766);
and U1108 (N_1108,N_743,N_790);
nand U1109 (N_1109,N_602,N_527);
xnor U1110 (N_1110,N_645,N_669);
and U1111 (N_1111,N_500,N_701);
nor U1112 (N_1112,N_811,N_933);
or U1113 (N_1113,N_756,N_755);
nor U1114 (N_1114,N_960,N_578);
and U1115 (N_1115,N_836,N_920);
nand U1116 (N_1116,N_571,N_986);
or U1117 (N_1117,N_583,N_731);
or U1118 (N_1118,N_977,N_860);
nor U1119 (N_1119,N_982,N_608);
and U1120 (N_1120,N_641,N_827);
nor U1121 (N_1121,N_570,N_973);
nor U1122 (N_1122,N_600,N_787);
nand U1123 (N_1123,N_599,N_765);
and U1124 (N_1124,N_834,N_636);
nor U1125 (N_1125,N_519,N_504);
xnor U1126 (N_1126,N_830,N_754);
xnor U1127 (N_1127,N_944,N_612);
and U1128 (N_1128,N_661,N_678);
xnor U1129 (N_1129,N_660,N_927);
or U1130 (N_1130,N_848,N_835);
xor U1131 (N_1131,N_929,N_771);
nand U1132 (N_1132,N_850,N_961);
nand U1133 (N_1133,N_812,N_904);
xor U1134 (N_1134,N_882,N_966);
xor U1135 (N_1135,N_821,N_575);
and U1136 (N_1136,N_919,N_905);
and U1137 (N_1137,N_579,N_685);
and U1138 (N_1138,N_994,N_528);
nand U1139 (N_1139,N_775,N_783);
xor U1140 (N_1140,N_705,N_975);
nand U1141 (N_1141,N_988,N_564);
and U1142 (N_1142,N_522,N_788);
and U1143 (N_1143,N_649,N_803);
and U1144 (N_1144,N_862,N_845);
xor U1145 (N_1145,N_520,N_763);
or U1146 (N_1146,N_562,N_884);
xor U1147 (N_1147,N_762,N_712);
or U1148 (N_1148,N_981,N_727);
and U1149 (N_1149,N_902,N_861);
nor U1150 (N_1150,N_995,N_901);
xor U1151 (N_1151,N_722,N_630);
and U1152 (N_1152,N_663,N_643);
or U1153 (N_1153,N_719,N_711);
or U1154 (N_1154,N_785,N_909);
nor U1155 (N_1155,N_843,N_736);
nor U1156 (N_1156,N_794,N_757);
xnor U1157 (N_1157,N_786,N_681);
or U1158 (N_1158,N_958,N_910);
nor U1159 (N_1159,N_815,N_859);
xor U1160 (N_1160,N_748,N_561);
xor U1161 (N_1161,N_609,N_577);
nand U1162 (N_1162,N_576,N_930);
or U1163 (N_1163,N_753,N_644);
or U1164 (N_1164,N_959,N_536);
or U1165 (N_1165,N_907,N_668);
xnor U1166 (N_1166,N_883,N_799);
nor U1167 (N_1167,N_704,N_618);
nor U1168 (N_1168,N_979,N_823);
nand U1169 (N_1169,N_505,N_546);
nor U1170 (N_1170,N_758,N_777);
and U1171 (N_1171,N_514,N_554);
xor U1172 (N_1172,N_747,N_865);
nand U1173 (N_1173,N_537,N_557);
xnor U1174 (N_1174,N_964,N_917);
xnor U1175 (N_1175,N_596,N_976);
xnor U1176 (N_1176,N_770,N_945);
nand U1177 (N_1177,N_970,N_581);
nand U1178 (N_1178,N_914,N_530);
or U1179 (N_1179,N_903,N_724);
nand U1180 (N_1180,N_990,N_713);
nor U1181 (N_1181,N_728,N_640);
xor U1182 (N_1182,N_744,N_831);
or U1183 (N_1183,N_580,N_906);
nand U1184 (N_1184,N_543,N_867);
nor U1185 (N_1185,N_587,N_623);
nand U1186 (N_1186,N_968,N_721);
xnor U1187 (N_1187,N_698,N_604);
xor U1188 (N_1188,N_833,N_912);
and U1189 (N_1189,N_851,N_838);
xor U1190 (N_1190,N_651,N_558);
or U1191 (N_1191,N_953,N_703);
xor U1192 (N_1192,N_574,N_971);
or U1193 (N_1193,N_897,N_533);
or U1194 (N_1194,N_592,N_619);
and U1195 (N_1195,N_793,N_631);
or U1196 (N_1196,N_518,N_538);
nor U1197 (N_1197,N_739,N_667);
or U1198 (N_1198,N_676,N_742);
nor U1199 (N_1199,N_517,N_702);
nor U1200 (N_1200,N_708,N_556);
nand U1201 (N_1201,N_697,N_997);
or U1202 (N_1202,N_715,N_806);
nor U1203 (N_1203,N_832,N_684);
and U1204 (N_1204,N_872,N_778);
or U1205 (N_1205,N_922,N_829);
xor U1206 (N_1206,N_863,N_940);
and U1207 (N_1207,N_800,N_664);
nor U1208 (N_1208,N_735,N_553);
nand U1209 (N_1209,N_694,N_679);
xnor U1210 (N_1210,N_692,N_750);
xor U1211 (N_1211,N_936,N_924);
nor U1212 (N_1212,N_868,N_854);
and U1213 (N_1213,N_813,N_913);
xor U1214 (N_1214,N_969,N_512);
nand U1215 (N_1215,N_734,N_723);
xnor U1216 (N_1216,N_565,N_965);
or U1217 (N_1217,N_686,N_752);
and U1218 (N_1218,N_782,N_824);
nor U1219 (N_1219,N_746,N_809);
xnor U1220 (N_1220,N_856,N_816);
or U1221 (N_1221,N_926,N_999);
or U1222 (N_1222,N_548,N_622);
xor U1223 (N_1223,N_928,N_725);
or U1224 (N_1224,N_648,N_716);
nand U1225 (N_1225,N_633,N_963);
nand U1226 (N_1226,N_784,N_898);
nor U1227 (N_1227,N_991,N_769);
xnor U1228 (N_1228,N_892,N_740);
nor U1229 (N_1229,N_601,N_626);
or U1230 (N_1230,N_506,N_983);
xor U1231 (N_1231,N_779,N_941);
and U1232 (N_1232,N_798,N_614);
xnor U1233 (N_1233,N_938,N_950);
xnor U1234 (N_1234,N_895,N_837);
or U1235 (N_1235,N_573,N_584);
xor U1236 (N_1236,N_887,N_791);
xnor U1237 (N_1237,N_749,N_761);
nor U1238 (N_1238,N_759,N_949);
and U1239 (N_1239,N_789,N_706);
nor U1240 (N_1240,N_985,N_857);
nand U1241 (N_1241,N_996,N_886);
nand U1242 (N_1242,N_634,N_842);
or U1243 (N_1243,N_687,N_690);
nor U1244 (N_1244,N_646,N_550);
and U1245 (N_1245,N_896,N_670);
or U1246 (N_1246,N_691,N_947);
or U1247 (N_1247,N_804,N_539);
xor U1248 (N_1248,N_509,N_826);
nor U1249 (N_1249,N_585,N_586);
xnor U1250 (N_1250,N_998,N_891);
and U1251 (N_1251,N_629,N_696);
nand U1252 (N_1252,N_507,N_970);
or U1253 (N_1253,N_799,N_551);
nand U1254 (N_1254,N_856,N_997);
xnor U1255 (N_1255,N_982,N_960);
or U1256 (N_1256,N_791,N_906);
xor U1257 (N_1257,N_756,N_667);
nor U1258 (N_1258,N_853,N_970);
or U1259 (N_1259,N_633,N_993);
xor U1260 (N_1260,N_645,N_884);
and U1261 (N_1261,N_586,N_707);
and U1262 (N_1262,N_526,N_544);
nand U1263 (N_1263,N_933,N_683);
and U1264 (N_1264,N_705,N_533);
and U1265 (N_1265,N_877,N_838);
xor U1266 (N_1266,N_925,N_649);
nand U1267 (N_1267,N_869,N_778);
xnor U1268 (N_1268,N_751,N_853);
nor U1269 (N_1269,N_946,N_810);
xor U1270 (N_1270,N_517,N_856);
or U1271 (N_1271,N_933,N_731);
and U1272 (N_1272,N_979,N_518);
nor U1273 (N_1273,N_564,N_740);
and U1274 (N_1274,N_744,N_922);
or U1275 (N_1275,N_656,N_657);
and U1276 (N_1276,N_922,N_679);
xor U1277 (N_1277,N_627,N_806);
and U1278 (N_1278,N_987,N_943);
nor U1279 (N_1279,N_588,N_673);
and U1280 (N_1280,N_637,N_525);
xor U1281 (N_1281,N_613,N_711);
and U1282 (N_1282,N_919,N_509);
nor U1283 (N_1283,N_820,N_823);
or U1284 (N_1284,N_704,N_696);
and U1285 (N_1285,N_843,N_931);
nor U1286 (N_1286,N_666,N_789);
nand U1287 (N_1287,N_501,N_557);
or U1288 (N_1288,N_893,N_536);
nand U1289 (N_1289,N_910,N_951);
and U1290 (N_1290,N_881,N_733);
or U1291 (N_1291,N_942,N_975);
nand U1292 (N_1292,N_878,N_926);
and U1293 (N_1293,N_653,N_768);
xnor U1294 (N_1294,N_656,N_700);
xnor U1295 (N_1295,N_774,N_583);
nand U1296 (N_1296,N_984,N_930);
nor U1297 (N_1297,N_567,N_618);
nor U1298 (N_1298,N_821,N_601);
xnor U1299 (N_1299,N_535,N_724);
xor U1300 (N_1300,N_663,N_631);
nand U1301 (N_1301,N_817,N_860);
nand U1302 (N_1302,N_823,N_540);
and U1303 (N_1303,N_820,N_765);
and U1304 (N_1304,N_971,N_578);
nor U1305 (N_1305,N_961,N_614);
and U1306 (N_1306,N_986,N_782);
nand U1307 (N_1307,N_716,N_686);
or U1308 (N_1308,N_604,N_530);
nand U1309 (N_1309,N_830,N_842);
or U1310 (N_1310,N_794,N_937);
and U1311 (N_1311,N_629,N_822);
or U1312 (N_1312,N_843,N_911);
or U1313 (N_1313,N_796,N_710);
or U1314 (N_1314,N_733,N_761);
or U1315 (N_1315,N_920,N_504);
nor U1316 (N_1316,N_674,N_666);
nand U1317 (N_1317,N_552,N_545);
nor U1318 (N_1318,N_836,N_774);
or U1319 (N_1319,N_805,N_546);
xnor U1320 (N_1320,N_854,N_719);
and U1321 (N_1321,N_803,N_695);
nor U1322 (N_1322,N_653,N_720);
xnor U1323 (N_1323,N_550,N_845);
xnor U1324 (N_1324,N_797,N_820);
or U1325 (N_1325,N_729,N_899);
nor U1326 (N_1326,N_988,N_961);
and U1327 (N_1327,N_972,N_629);
nor U1328 (N_1328,N_983,N_921);
or U1329 (N_1329,N_557,N_712);
or U1330 (N_1330,N_799,N_550);
or U1331 (N_1331,N_519,N_838);
or U1332 (N_1332,N_608,N_854);
nand U1333 (N_1333,N_765,N_978);
and U1334 (N_1334,N_708,N_501);
xnor U1335 (N_1335,N_906,N_585);
nand U1336 (N_1336,N_705,N_677);
nand U1337 (N_1337,N_780,N_895);
nand U1338 (N_1338,N_961,N_875);
and U1339 (N_1339,N_644,N_741);
xor U1340 (N_1340,N_560,N_680);
nand U1341 (N_1341,N_568,N_774);
and U1342 (N_1342,N_593,N_908);
or U1343 (N_1343,N_906,N_899);
nand U1344 (N_1344,N_835,N_992);
nor U1345 (N_1345,N_876,N_740);
nand U1346 (N_1346,N_755,N_802);
xor U1347 (N_1347,N_505,N_858);
or U1348 (N_1348,N_897,N_851);
nand U1349 (N_1349,N_615,N_962);
nor U1350 (N_1350,N_899,N_767);
xor U1351 (N_1351,N_511,N_843);
nand U1352 (N_1352,N_547,N_772);
or U1353 (N_1353,N_569,N_572);
nor U1354 (N_1354,N_936,N_544);
and U1355 (N_1355,N_754,N_698);
or U1356 (N_1356,N_862,N_786);
nor U1357 (N_1357,N_701,N_730);
or U1358 (N_1358,N_827,N_875);
and U1359 (N_1359,N_836,N_763);
or U1360 (N_1360,N_669,N_779);
and U1361 (N_1361,N_665,N_501);
xnor U1362 (N_1362,N_633,N_893);
or U1363 (N_1363,N_784,N_607);
xor U1364 (N_1364,N_801,N_601);
xor U1365 (N_1365,N_829,N_747);
and U1366 (N_1366,N_996,N_988);
and U1367 (N_1367,N_800,N_791);
nand U1368 (N_1368,N_798,N_902);
nor U1369 (N_1369,N_531,N_944);
nand U1370 (N_1370,N_955,N_567);
xnor U1371 (N_1371,N_504,N_960);
nor U1372 (N_1372,N_647,N_740);
or U1373 (N_1373,N_554,N_848);
nor U1374 (N_1374,N_977,N_738);
and U1375 (N_1375,N_799,N_848);
xor U1376 (N_1376,N_630,N_726);
nor U1377 (N_1377,N_632,N_823);
or U1378 (N_1378,N_646,N_733);
nand U1379 (N_1379,N_525,N_802);
and U1380 (N_1380,N_675,N_889);
xnor U1381 (N_1381,N_848,N_927);
xor U1382 (N_1382,N_772,N_965);
nor U1383 (N_1383,N_944,N_895);
nor U1384 (N_1384,N_836,N_938);
xor U1385 (N_1385,N_719,N_784);
or U1386 (N_1386,N_726,N_612);
nor U1387 (N_1387,N_573,N_525);
or U1388 (N_1388,N_568,N_636);
nand U1389 (N_1389,N_740,N_838);
nand U1390 (N_1390,N_788,N_524);
nor U1391 (N_1391,N_846,N_738);
xnor U1392 (N_1392,N_958,N_742);
or U1393 (N_1393,N_523,N_611);
xor U1394 (N_1394,N_639,N_751);
nor U1395 (N_1395,N_583,N_640);
or U1396 (N_1396,N_756,N_625);
xor U1397 (N_1397,N_692,N_501);
nor U1398 (N_1398,N_601,N_569);
and U1399 (N_1399,N_760,N_704);
nor U1400 (N_1400,N_653,N_602);
and U1401 (N_1401,N_857,N_640);
and U1402 (N_1402,N_619,N_561);
xnor U1403 (N_1403,N_849,N_505);
and U1404 (N_1404,N_562,N_535);
and U1405 (N_1405,N_545,N_546);
xnor U1406 (N_1406,N_667,N_703);
xor U1407 (N_1407,N_888,N_561);
nand U1408 (N_1408,N_985,N_503);
and U1409 (N_1409,N_988,N_703);
nor U1410 (N_1410,N_749,N_680);
xnor U1411 (N_1411,N_912,N_594);
and U1412 (N_1412,N_982,N_777);
nand U1413 (N_1413,N_791,N_830);
or U1414 (N_1414,N_831,N_668);
and U1415 (N_1415,N_538,N_719);
and U1416 (N_1416,N_969,N_505);
xnor U1417 (N_1417,N_538,N_744);
and U1418 (N_1418,N_520,N_741);
or U1419 (N_1419,N_885,N_552);
nand U1420 (N_1420,N_756,N_983);
xor U1421 (N_1421,N_931,N_861);
nor U1422 (N_1422,N_835,N_906);
nor U1423 (N_1423,N_750,N_726);
nor U1424 (N_1424,N_801,N_821);
and U1425 (N_1425,N_926,N_953);
nand U1426 (N_1426,N_804,N_847);
xnor U1427 (N_1427,N_753,N_625);
or U1428 (N_1428,N_675,N_777);
xor U1429 (N_1429,N_924,N_810);
nor U1430 (N_1430,N_591,N_583);
and U1431 (N_1431,N_865,N_643);
xor U1432 (N_1432,N_777,N_970);
nor U1433 (N_1433,N_762,N_536);
xor U1434 (N_1434,N_939,N_900);
xor U1435 (N_1435,N_782,N_928);
and U1436 (N_1436,N_539,N_805);
nand U1437 (N_1437,N_644,N_849);
or U1438 (N_1438,N_613,N_944);
nand U1439 (N_1439,N_533,N_636);
xnor U1440 (N_1440,N_580,N_943);
nor U1441 (N_1441,N_604,N_927);
xnor U1442 (N_1442,N_648,N_524);
or U1443 (N_1443,N_509,N_548);
nand U1444 (N_1444,N_783,N_500);
nand U1445 (N_1445,N_749,N_937);
nand U1446 (N_1446,N_912,N_760);
nand U1447 (N_1447,N_554,N_929);
nand U1448 (N_1448,N_936,N_612);
nor U1449 (N_1449,N_552,N_770);
or U1450 (N_1450,N_508,N_550);
nand U1451 (N_1451,N_717,N_617);
and U1452 (N_1452,N_623,N_919);
xnor U1453 (N_1453,N_709,N_824);
nand U1454 (N_1454,N_525,N_959);
nor U1455 (N_1455,N_959,N_705);
xor U1456 (N_1456,N_701,N_769);
nand U1457 (N_1457,N_630,N_959);
or U1458 (N_1458,N_908,N_927);
xor U1459 (N_1459,N_924,N_802);
or U1460 (N_1460,N_885,N_560);
nand U1461 (N_1461,N_503,N_619);
xnor U1462 (N_1462,N_946,N_913);
nand U1463 (N_1463,N_985,N_973);
xnor U1464 (N_1464,N_690,N_583);
xor U1465 (N_1465,N_756,N_518);
or U1466 (N_1466,N_655,N_742);
nor U1467 (N_1467,N_722,N_713);
nor U1468 (N_1468,N_602,N_918);
or U1469 (N_1469,N_651,N_602);
and U1470 (N_1470,N_769,N_961);
nor U1471 (N_1471,N_510,N_994);
xor U1472 (N_1472,N_520,N_863);
nand U1473 (N_1473,N_890,N_922);
nand U1474 (N_1474,N_954,N_658);
and U1475 (N_1475,N_631,N_685);
nand U1476 (N_1476,N_861,N_534);
nand U1477 (N_1477,N_534,N_868);
nand U1478 (N_1478,N_953,N_544);
nand U1479 (N_1479,N_526,N_728);
and U1480 (N_1480,N_678,N_641);
xor U1481 (N_1481,N_975,N_674);
nor U1482 (N_1482,N_947,N_702);
nor U1483 (N_1483,N_776,N_883);
or U1484 (N_1484,N_815,N_862);
nor U1485 (N_1485,N_681,N_600);
xor U1486 (N_1486,N_557,N_538);
nand U1487 (N_1487,N_661,N_615);
and U1488 (N_1488,N_819,N_741);
and U1489 (N_1489,N_628,N_609);
xor U1490 (N_1490,N_851,N_834);
xnor U1491 (N_1491,N_735,N_830);
xor U1492 (N_1492,N_856,N_609);
nor U1493 (N_1493,N_889,N_778);
xor U1494 (N_1494,N_744,N_535);
xnor U1495 (N_1495,N_780,N_934);
and U1496 (N_1496,N_931,N_560);
xor U1497 (N_1497,N_865,N_765);
or U1498 (N_1498,N_932,N_815);
nand U1499 (N_1499,N_538,N_983);
or U1500 (N_1500,N_1212,N_1474);
and U1501 (N_1501,N_1023,N_1391);
and U1502 (N_1502,N_1339,N_1043);
xor U1503 (N_1503,N_1269,N_1187);
nor U1504 (N_1504,N_1238,N_1007);
and U1505 (N_1505,N_1283,N_1094);
nor U1506 (N_1506,N_1164,N_1211);
nand U1507 (N_1507,N_1114,N_1080);
and U1508 (N_1508,N_1086,N_1268);
xor U1509 (N_1509,N_1064,N_1001);
and U1510 (N_1510,N_1360,N_1173);
or U1511 (N_1511,N_1150,N_1319);
or U1512 (N_1512,N_1108,N_1146);
or U1513 (N_1513,N_1099,N_1200);
nand U1514 (N_1514,N_1247,N_1366);
nand U1515 (N_1515,N_1470,N_1324);
or U1516 (N_1516,N_1098,N_1165);
nor U1517 (N_1517,N_1465,N_1447);
nor U1518 (N_1518,N_1184,N_1107);
nor U1519 (N_1519,N_1275,N_1198);
or U1520 (N_1520,N_1091,N_1393);
and U1521 (N_1521,N_1049,N_1430);
and U1522 (N_1522,N_1399,N_1125);
or U1523 (N_1523,N_1045,N_1398);
or U1524 (N_1524,N_1051,N_1496);
nand U1525 (N_1525,N_1300,N_1264);
and U1526 (N_1526,N_1342,N_1403);
nand U1527 (N_1527,N_1185,N_1016);
or U1528 (N_1528,N_1374,N_1149);
and U1529 (N_1529,N_1229,N_1303);
xor U1530 (N_1530,N_1156,N_1097);
and U1531 (N_1531,N_1239,N_1122);
xor U1532 (N_1532,N_1132,N_1490);
xor U1533 (N_1533,N_1231,N_1009);
and U1534 (N_1534,N_1261,N_1371);
xor U1535 (N_1535,N_1406,N_1158);
nor U1536 (N_1536,N_1116,N_1127);
xor U1537 (N_1537,N_1473,N_1380);
nor U1538 (N_1538,N_1110,N_1040);
nor U1539 (N_1539,N_1224,N_1359);
nand U1540 (N_1540,N_1218,N_1081);
xor U1541 (N_1541,N_1017,N_1196);
or U1542 (N_1542,N_1178,N_1208);
nor U1543 (N_1543,N_1452,N_1401);
nand U1544 (N_1544,N_1139,N_1028);
and U1545 (N_1545,N_1278,N_1032);
nor U1546 (N_1546,N_1070,N_1498);
nand U1547 (N_1547,N_1281,N_1256);
nor U1548 (N_1548,N_1321,N_1460);
nor U1549 (N_1549,N_1076,N_1355);
xnor U1550 (N_1550,N_1249,N_1482);
or U1551 (N_1551,N_1134,N_1159);
nand U1552 (N_1552,N_1414,N_1033);
nor U1553 (N_1553,N_1083,N_1135);
nor U1554 (N_1554,N_1320,N_1318);
nor U1555 (N_1555,N_1075,N_1004);
nor U1556 (N_1556,N_1106,N_1494);
xor U1557 (N_1557,N_1217,N_1453);
nand U1558 (N_1558,N_1464,N_1332);
xor U1559 (N_1559,N_1069,N_1000);
nor U1560 (N_1560,N_1243,N_1432);
xnor U1561 (N_1561,N_1216,N_1109);
or U1562 (N_1562,N_1499,N_1410);
nand U1563 (N_1563,N_1316,N_1126);
or U1564 (N_1564,N_1131,N_1307);
nor U1565 (N_1565,N_1455,N_1423);
xnor U1566 (N_1566,N_1317,N_1351);
or U1567 (N_1567,N_1129,N_1044);
xnor U1568 (N_1568,N_1330,N_1199);
xor U1569 (N_1569,N_1133,N_1101);
and U1570 (N_1570,N_1357,N_1444);
nand U1571 (N_1571,N_1246,N_1367);
nor U1572 (N_1572,N_1345,N_1331);
xnor U1573 (N_1573,N_1215,N_1418);
or U1574 (N_1574,N_1475,N_1119);
or U1575 (N_1575,N_1191,N_1334);
and U1576 (N_1576,N_1308,N_1435);
and U1577 (N_1577,N_1036,N_1120);
and U1578 (N_1578,N_1412,N_1177);
xor U1579 (N_1579,N_1195,N_1483);
and U1580 (N_1580,N_1188,N_1254);
or U1581 (N_1581,N_1221,N_1061);
xnor U1582 (N_1582,N_1244,N_1388);
nor U1583 (N_1583,N_1370,N_1118);
and U1584 (N_1584,N_1287,N_1011);
nor U1585 (N_1585,N_1271,N_1006);
xnor U1586 (N_1586,N_1207,N_1486);
and U1587 (N_1587,N_1192,N_1458);
or U1588 (N_1588,N_1340,N_1030);
or U1589 (N_1589,N_1258,N_1492);
xor U1590 (N_1590,N_1471,N_1230);
nor U1591 (N_1591,N_1142,N_1143);
and U1592 (N_1592,N_1089,N_1273);
nor U1593 (N_1593,N_1111,N_1136);
nor U1594 (N_1594,N_1093,N_1379);
nor U1595 (N_1595,N_1445,N_1270);
or U1596 (N_1596,N_1301,N_1228);
nand U1597 (N_1597,N_1404,N_1209);
nor U1598 (N_1598,N_1052,N_1341);
nor U1599 (N_1599,N_1441,N_1042);
nor U1600 (N_1600,N_1087,N_1297);
and U1601 (N_1601,N_1197,N_1488);
xor U1602 (N_1602,N_1237,N_1123);
nand U1603 (N_1603,N_1480,N_1153);
and U1604 (N_1604,N_1227,N_1276);
and U1605 (N_1605,N_1395,N_1233);
and U1606 (N_1606,N_1425,N_1053);
nand U1607 (N_1607,N_1020,N_1364);
xor U1608 (N_1608,N_1299,N_1124);
nand U1609 (N_1609,N_1417,N_1386);
or U1610 (N_1610,N_1206,N_1013);
nand U1611 (N_1611,N_1409,N_1223);
xnor U1612 (N_1612,N_1434,N_1257);
or U1613 (N_1613,N_1008,N_1151);
nor U1614 (N_1614,N_1189,N_1012);
and U1615 (N_1615,N_1282,N_1429);
xnor U1616 (N_1616,N_1352,N_1362);
nand U1617 (N_1617,N_1039,N_1161);
nor U1618 (N_1618,N_1067,N_1346);
nor U1619 (N_1619,N_1183,N_1497);
and U1620 (N_1620,N_1438,N_1493);
nand U1621 (N_1621,N_1066,N_1427);
or U1622 (N_1622,N_1433,N_1495);
and U1623 (N_1623,N_1236,N_1251);
nor U1624 (N_1624,N_1400,N_1485);
nand U1625 (N_1625,N_1377,N_1446);
nand U1626 (N_1626,N_1029,N_1112);
and U1627 (N_1627,N_1113,N_1288);
and U1628 (N_1628,N_1085,N_1137);
nand U1629 (N_1629,N_1226,N_1448);
nand U1630 (N_1630,N_1130,N_1372);
nand U1631 (N_1631,N_1103,N_1296);
nor U1632 (N_1632,N_1079,N_1078);
xor U1633 (N_1633,N_1356,N_1484);
xnor U1634 (N_1634,N_1267,N_1387);
or U1635 (N_1635,N_1326,N_1385);
xnor U1636 (N_1636,N_1344,N_1263);
nor U1637 (N_1637,N_1163,N_1337);
xor U1638 (N_1638,N_1477,N_1375);
xnor U1639 (N_1639,N_1424,N_1059);
xnor U1640 (N_1640,N_1478,N_1312);
nor U1641 (N_1641,N_1408,N_1095);
and U1642 (N_1642,N_1309,N_1396);
or U1643 (N_1643,N_1071,N_1462);
xnor U1644 (N_1644,N_1201,N_1411);
or U1645 (N_1645,N_1304,N_1284);
nor U1646 (N_1646,N_1280,N_1181);
nand U1647 (N_1647,N_1214,N_1128);
or U1648 (N_1648,N_1358,N_1294);
xor U1649 (N_1649,N_1290,N_1219);
nand U1650 (N_1650,N_1415,N_1186);
and U1651 (N_1651,N_1378,N_1323);
or U1652 (N_1652,N_1003,N_1402);
nand U1653 (N_1653,N_1073,N_1147);
xor U1654 (N_1654,N_1274,N_1353);
nor U1655 (N_1655,N_1234,N_1428);
and U1656 (N_1656,N_1056,N_1327);
and U1657 (N_1657,N_1397,N_1157);
and U1658 (N_1658,N_1363,N_1205);
and U1659 (N_1659,N_1407,N_1361);
nor U1660 (N_1660,N_1382,N_1384);
or U1661 (N_1661,N_1333,N_1048);
or U1662 (N_1662,N_1405,N_1311);
nand U1663 (N_1663,N_1390,N_1381);
and U1664 (N_1664,N_1060,N_1027);
xor U1665 (N_1665,N_1015,N_1115);
and U1666 (N_1666,N_1065,N_1176);
xor U1667 (N_1667,N_1014,N_1459);
and U1668 (N_1668,N_1072,N_1285);
and U1669 (N_1669,N_1062,N_1487);
xnor U1670 (N_1670,N_1148,N_1437);
xnor U1671 (N_1671,N_1350,N_1225);
xnor U1672 (N_1672,N_1169,N_1456);
or U1673 (N_1673,N_1038,N_1373);
xor U1674 (N_1674,N_1266,N_1063);
nor U1675 (N_1675,N_1343,N_1250);
nand U1676 (N_1676,N_1240,N_1140);
xnor U1677 (N_1677,N_1325,N_1025);
or U1678 (N_1678,N_1489,N_1092);
or U1679 (N_1679,N_1175,N_1138);
nand U1680 (N_1680,N_1431,N_1041);
nor U1681 (N_1681,N_1252,N_1024);
xor U1682 (N_1682,N_1248,N_1315);
nor U1683 (N_1683,N_1210,N_1174);
or U1684 (N_1684,N_1467,N_1034);
and U1685 (N_1685,N_1102,N_1213);
nor U1686 (N_1686,N_1348,N_1117);
nand U1687 (N_1687,N_1232,N_1292);
or U1688 (N_1688,N_1472,N_1259);
nor U1689 (N_1689,N_1277,N_1298);
nor U1690 (N_1690,N_1194,N_1204);
xnor U1691 (N_1691,N_1104,N_1160);
and U1692 (N_1692,N_1466,N_1416);
or U1693 (N_1693,N_1295,N_1255);
xor U1694 (N_1694,N_1121,N_1260);
and U1695 (N_1695,N_1152,N_1105);
nand U1696 (N_1696,N_1306,N_1293);
and U1697 (N_1697,N_1057,N_1026);
or U1698 (N_1698,N_1481,N_1180);
nor U1699 (N_1699,N_1328,N_1368);
nand U1700 (N_1700,N_1154,N_1421);
nor U1701 (N_1701,N_1253,N_1338);
nand U1702 (N_1702,N_1235,N_1439);
and U1703 (N_1703,N_1171,N_1347);
and U1704 (N_1704,N_1422,N_1469);
nor U1705 (N_1705,N_1090,N_1047);
nand U1706 (N_1706,N_1286,N_1389);
xnor U1707 (N_1707,N_1335,N_1037);
and U1708 (N_1708,N_1005,N_1426);
xor U1709 (N_1709,N_1021,N_1443);
nor U1710 (N_1710,N_1454,N_1450);
or U1711 (N_1711,N_1245,N_1449);
xnor U1712 (N_1712,N_1322,N_1084);
nand U1713 (N_1713,N_1461,N_1050);
or U1714 (N_1714,N_1310,N_1167);
or U1715 (N_1715,N_1046,N_1314);
xnor U1716 (N_1716,N_1182,N_1336);
nand U1717 (N_1717,N_1010,N_1365);
xor U1718 (N_1718,N_1100,N_1088);
or U1719 (N_1719,N_1272,N_1468);
xnor U1720 (N_1720,N_1442,N_1162);
nor U1721 (N_1721,N_1383,N_1222);
and U1722 (N_1722,N_1436,N_1220);
nor U1723 (N_1723,N_1068,N_1190);
or U1724 (N_1724,N_1392,N_1313);
nand U1725 (N_1725,N_1203,N_1262);
nand U1726 (N_1726,N_1420,N_1058);
nor U1727 (N_1727,N_1394,N_1242);
or U1728 (N_1728,N_1413,N_1265);
or U1729 (N_1729,N_1369,N_1141);
nor U1730 (N_1730,N_1166,N_1022);
nand U1731 (N_1731,N_1054,N_1031);
nor U1732 (N_1732,N_1074,N_1055);
nor U1733 (N_1733,N_1241,N_1155);
or U1734 (N_1734,N_1279,N_1305);
nor U1735 (N_1735,N_1144,N_1376);
or U1736 (N_1736,N_1302,N_1035);
nand U1737 (N_1737,N_1289,N_1179);
xnor U1738 (N_1738,N_1329,N_1202);
xor U1739 (N_1739,N_1354,N_1018);
nor U1740 (N_1740,N_1170,N_1019);
xor U1741 (N_1741,N_1291,N_1168);
nand U1742 (N_1742,N_1457,N_1077);
and U1743 (N_1743,N_1082,N_1002);
nand U1744 (N_1744,N_1193,N_1476);
or U1745 (N_1745,N_1349,N_1479);
and U1746 (N_1746,N_1451,N_1440);
or U1747 (N_1747,N_1145,N_1419);
or U1748 (N_1748,N_1172,N_1096);
and U1749 (N_1749,N_1463,N_1491);
xnor U1750 (N_1750,N_1049,N_1102);
or U1751 (N_1751,N_1055,N_1275);
or U1752 (N_1752,N_1397,N_1058);
nor U1753 (N_1753,N_1056,N_1039);
and U1754 (N_1754,N_1282,N_1165);
xnor U1755 (N_1755,N_1266,N_1322);
nand U1756 (N_1756,N_1397,N_1428);
and U1757 (N_1757,N_1089,N_1246);
xor U1758 (N_1758,N_1107,N_1208);
nand U1759 (N_1759,N_1357,N_1487);
or U1760 (N_1760,N_1131,N_1175);
or U1761 (N_1761,N_1484,N_1144);
and U1762 (N_1762,N_1376,N_1212);
nand U1763 (N_1763,N_1123,N_1161);
or U1764 (N_1764,N_1187,N_1439);
nor U1765 (N_1765,N_1277,N_1043);
nand U1766 (N_1766,N_1297,N_1222);
nand U1767 (N_1767,N_1298,N_1386);
nor U1768 (N_1768,N_1291,N_1127);
xnor U1769 (N_1769,N_1309,N_1220);
xnor U1770 (N_1770,N_1383,N_1240);
nor U1771 (N_1771,N_1394,N_1386);
xnor U1772 (N_1772,N_1433,N_1165);
xnor U1773 (N_1773,N_1299,N_1414);
or U1774 (N_1774,N_1291,N_1220);
xnor U1775 (N_1775,N_1137,N_1171);
or U1776 (N_1776,N_1358,N_1181);
nand U1777 (N_1777,N_1235,N_1031);
and U1778 (N_1778,N_1038,N_1012);
or U1779 (N_1779,N_1236,N_1011);
and U1780 (N_1780,N_1065,N_1044);
nand U1781 (N_1781,N_1209,N_1393);
or U1782 (N_1782,N_1436,N_1036);
and U1783 (N_1783,N_1169,N_1093);
nor U1784 (N_1784,N_1300,N_1031);
and U1785 (N_1785,N_1197,N_1181);
and U1786 (N_1786,N_1046,N_1254);
xnor U1787 (N_1787,N_1467,N_1322);
nor U1788 (N_1788,N_1384,N_1005);
or U1789 (N_1789,N_1185,N_1398);
and U1790 (N_1790,N_1000,N_1083);
or U1791 (N_1791,N_1006,N_1160);
or U1792 (N_1792,N_1331,N_1400);
and U1793 (N_1793,N_1317,N_1322);
nand U1794 (N_1794,N_1166,N_1155);
or U1795 (N_1795,N_1114,N_1295);
nor U1796 (N_1796,N_1330,N_1452);
nor U1797 (N_1797,N_1082,N_1125);
nand U1798 (N_1798,N_1230,N_1413);
xnor U1799 (N_1799,N_1317,N_1175);
and U1800 (N_1800,N_1166,N_1045);
xor U1801 (N_1801,N_1330,N_1329);
nand U1802 (N_1802,N_1474,N_1332);
or U1803 (N_1803,N_1233,N_1154);
nand U1804 (N_1804,N_1116,N_1146);
nor U1805 (N_1805,N_1259,N_1019);
xor U1806 (N_1806,N_1160,N_1251);
nor U1807 (N_1807,N_1430,N_1213);
xor U1808 (N_1808,N_1070,N_1270);
or U1809 (N_1809,N_1471,N_1048);
and U1810 (N_1810,N_1321,N_1436);
nor U1811 (N_1811,N_1416,N_1321);
nor U1812 (N_1812,N_1405,N_1186);
or U1813 (N_1813,N_1072,N_1379);
and U1814 (N_1814,N_1361,N_1302);
nor U1815 (N_1815,N_1144,N_1277);
nor U1816 (N_1816,N_1275,N_1123);
nor U1817 (N_1817,N_1067,N_1297);
nor U1818 (N_1818,N_1138,N_1497);
nand U1819 (N_1819,N_1075,N_1165);
nor U1820 (N_1820,N_1360,N_1330);
nand U1821 (N_1821,N_1421,N_1220);
nand U1822 (N_1822,N_1393,N_1017);
or U1823 (N_1823,N_1423,N_1258);
xor U1824 (N_1824,N_1011,N_1451);
and U1825 (N_1825,N_1348,N_1122);
nor U1826 (N_1826,N_1245,N_1020);
and U1827 (N_1827,N_1237,N_1179);
or U1828 (N_1828,N_1247,N_1022);
xor U1829 (N_1829,N_1325,N_1010);
nor U1830 (N_1830,N_1413,N_1267);
nor U1831 (N_1831,N_1292,N_1007);
and U1832 (N_1832,N_1388,N_1039);
xnor U1833 (N_1833,N_1411,N_1195);
nor U1834 (N_1834,N_1165,N_1474);
nand U1835 (N_1835,N_1261,N_1287);
and U1836 (N_1836,N_1413,N_1185);
nor U1837 (N_1837,N_1292,N_1008);
xor U1838 (N_1838,N_1056,N_1014);
xor U1839 (N_1839,N_1175,N_1413);
xnor U1840 (N_1840,N_1085,N_1284);
nor U1841 (N_1841,N_1202,N_1021);
nand U1842 (N_1842,N_1124,N_1230);
and U1843 (N_1843,N_1174,N_1242);
and U1844 (N_1844,N_1384,N_1453);
nor U1845 (N_1845,N_1051,N_1184);
and U1846 (N_1846,N_1360,N_1497);
nor U1847 (N_1847,N_1380,N_1079);
and U1848 (N_1848,N_1109,N_1425);
and U1849 (N_1849,N_1281,N_1199);
nand U1850 (N_1850,N_1189,N_1382);
nand U1851 (N_1851,N_1110,N_1268);
and U1852 (N_1852,N_1063,N_1012);
xnor U1853 (N_1853,N_1366,N_1365);
and U1854 (N_1854,N_1310,N_1240);
xnor U1855 (N_1855,N_1080,N_1021);
and U1856 (N_1856,N_1107,N_1158);
or U1857 (N_1857,N_1414,N_1352);
nor U1858 (N_1858,N_1316,N_1142);
xor U1859 (N_1859,N_1127,N_1040);
nor U1860 (N_1860,N_1151,N_1075);
xnor U1861 (N_1861,N_1234,N_1171);
nand U1862 (N_1862,N_1425,N_1066);
or U1863 (N_1863,N_1225,N_1338);
xor U1864 (N_1864,N_1189,N_1237);
nor U1865 (N_1865,N_1320,N_1490);
or U1866 (N_1866,N_1156,N_1121);
xor U1867 (N_1867,N_1263,N_1005);
xor U1868 (N_1868,N_1403,N_1490);
nand U1869 (N_1869,N_1045,N_1338);
xor U1870 (N_1870,N_1298,N_1306);
xor U1871 (N_1871,N_1023,N_1220);
xnor U1872 (N_1872,N_1490,N_1478);
and U1873 (N_1873,N_1130,N_1406);
or U1874 (N_1874,N_1190,N_1114);
nand U1875 (N_1875,N_1234,N_1161);
xnor U1876 (N_1876,N_1030,N_1058);
nand U1877 (N_1877,N_1478,N_1462);
xnor U1878 (N_1878,N_1151,N_1095);
nand U1879 (N_1879,N_1374,N_1369);
and U1880 (N_1880,N_1140,N_1368);
xor U1881 (N_1881,N_1108,N_1372);
nor U1882 (N_1882,N_1178,N_1456);
nor U1883 (N_1883,N_1436,N_1397);
or U1884 (N_1884,N_1154,N_1035);
and U1885 (N_1885,N_1133,N_1155);
or U1886 (N_1886,N_1203,N_1416);
and U1887 (N_1887,N_1072,N_1433);
nand U1888 (N_1888,N_1329,N_1222);
or U1889 (N_1889,N_1146,N_1485);
and U1890 (N_1890,N_1017,N_1179);
and U1891 (N_1891,N_1053,N_1198);
and U1892 (N_1892,N_1102,N_1300);
nor U1893 (N_1893,N_1215,N_1317);
nand U1894 (N_1894,N_1497,N_1399);
or U1895 (N_1895,N_1378,N_1107);
nand U1896 (N_1896,N_1377,N_1480);
xor U1897 (N_1897,N_1213,N_1258);
nor U1898 (N_1898,N_1045,N_1288);
xnor U1899 (N_1899,N_1257,N_1243);
nor U1900 (N_1900,N_1452,N_1472);
xnor U1901 (N_1901,N_1315,N_1478);
and U1902 (N_1902,N_1433,N_1304);
and U1903 (N_1903,N_1079,N_1421);
nand U1904 (N_1904,N_1280,N_1145);
and U1905 (N_1905,N_1384,N_1006);
or U1906 (N_1906,N_1413,N_1025);
nand U1907 (N_1907,N_1284,N_1486);
xor U1908 (N_1908,N_1315,N_1310);
and U1909 (N_1909,N_1094,N_1251);
and U1910 (N_1910,N_1166,N_1364);
or U1911 (N_1911,N_1435,N_1260);
xor U1912 (N_1912,N_1494,N_1229);
xor U1913 (N_1913,N_1139,N_1374);
nand U1914 (N_1914,N_1385,N_1254);
xor U1915 (N_1915,N_1032,N_1334);
and U1916 (N_1916,N_1320,N_1200);
or U1917 (N_1917,N_1049,N_1048);
nand U1918 (N_1918,N_1168,N_1126);
nor U1919 (N_1919,N_1423,N_1259);
or U1920 (N_1920,N_1223,N_1424);
nor U1921 (N_1921,N_1104,N_1496);
and U1922 (N_1922,N_1219,N_1472);
and U1923 (N_1923,N_1203,N_1283);
nand U1924 (N_1924,N_1189,N_1066);
nor U1925 (N_1925,N_1441,N_1296);
nor U1926 (N_1926,N_1051,N_1000);
and U1927 (N_1927,N_1073,N_1403);
or U1928 (N_1928,N_1254,N_1073);
nand U1929 (N_1929,N_1353,N_1322);
or U1930 (N_1930,N_1136,N_1330);
xnor U1931 (N_1931,N_1288,N_1056);
xor U1932 (N_1932,N_1240,N_1264);
xor U1933 (N_1933,N_1452,N_1005);
xor U1934 (N_1934,N_1208,N_1130);
nor U1935 (N_1935,N_1322,N_1487);
and U1936 (N_1936,N_1443,N_1483);
and U1937 (N_1937,N_1442,N_1409);
nand U1938 (N_1938,N_1081,N_1315);
nor U1939 (N_1939,N_1100,N_1340);
and U1940 (N_1940,N_1349,N_1137);
nand U1941 (N_1941,N_1389,N_1014);
nand U1942 (N_1942,N_1134,N_1408);
or U1943 (N_1943,N_1146,N_1328);
xor U1944 (N_1944,N_1019,N_1348);
nand U1945 (N_1945,N_1236,N_1197);
nand U1946 (N_1946,N_1193,N_1479);
nor U1947 (N_1947,N_1146,N_1185);
and U1948 (N_1948,N_1275,N_1359);
nand U1949 (N_1949,N_1283,N_1366);
nand U1950 (N_1950,N_1186,N_1235);
nor U1951 (N_1951,N_1222,N_1133);
nand U1952 (N_1952,N_1020,N_1163);
xor U1953 (N_1953,N_1023,N_1124);
or U1954 (N_1954,N_1011,N_1395);
nand U1955 (N_1955,N_1096,N_1372);
nand U1956 (N_1956,N_1388,N_1442);
nor U1957 (N_1957,N_1038,N_1382);
nand U1958 (N_1958,N_1103,N_1281);
and U1959 (N_1959,N_1292,N_1088);
nor U1960 (N_1960,N_1334,N_1212);
nor U1961 (N_1961,N_1037,N_1426);
nand U1962 (N_1962,N_1143,N_1279);
or U1963 (N_1963,N_1148,N_1052);
nand U1964 (N_1964,N_1452,N_1419);
xnor U1965 (N_1965,N_1090,N_1276);
nand U1966 (N_1966,N_1195,N_1156);
or U1967 (N_1967,N_1437,N_1176);
nand U1968 (N_1968,N_1421,N_1218);
and U1969 (N_1969,N_1135,N_1438);
nand U1970 (N_1970,N_1032,N_1399);
nor U1971 (N_1971,N_1000,N_1275);
nand U1972 (N_1972,N_1402,N_1004);
nand U1973 (N_1973,N_1483,N_1065);
nand U1974 (N_1974,N_1255,N_1279);
nand U1975 (N_1975,N_1423,N_1158);
xor U1976 (N_1976,N_1248,N_1053);
nand U1977 (N_1977,N_1306,N_1375);
and U1978 (N_1978,N_1416,N_1317);
nand U1979 (N_1979,N_1227,N_1321);
nor U1980 (N_1980,N_1164,N_1204);
or U1981 (N_1981,N_1430,N_1078);
and U1982 (N_1982,N_1438,N_1398);
or U1983 (N_1983,N_1292,N_1072);
nand U1984 (N_1984,N_1279,N_1308);
or U1985 (N_1985,N_1220,N_1324);
xor U1986 (N_1986,N_1415,N_1069);
nor U1987 (N_1987,N_1209,N_1172);
nor U1988 (N_1988,N_1461,N_1078);
nand U1989 (N_1989,N_1361,N_1386);
or U1990 (N_1990,N_1085,N_1377);
xor U1991 (N_1991,N_1388,N_1365);
nand U1992 (N_1992,N_1324,N_1465);
xor U1993 (N_1993,N_1280,N_1315);
or U1994 (N_1994,N_1320,N_1278);
nor U1995 (N_1995,N_1448,N_1440);
nor U1996 (N_1996,N_1065,N_1073);
xnor U1997 (N_1997,N_1190,N_1253);
xor U1998 (N_1998,N_1412,N_1362);
or U1999 (N_1999,N_1324,N_1081);
and U2000 (N_2000,N_1629,N_1807);
or U2001 (N_2001,N_1533,N_1923);
xor U2002 (N_2002,N_1635,N_1858);
or U2003 (N_2003,N_1738,N_1996);
nor U2004 (N_2004,N_1985,N_1731);
nand U2005 (N_2005,N_1880,N_1943);
or U2006 (N_2006,N_1556,N_1568);
nor U2007 (N_2007,N_1976,N_1619);
and U2008 (N_2008,N_1925,N_1734);
nand U2009 (N_2009,N_1674,N_1566);
nand U2010 (N_2010,N_1979,N_1969);
or U2011 (N_2011,N_1602,N_1643);
xnor U2012 (N_2012,N_1912,N_1722);
nand U2013 (N_2013,N_1820,N_1961);
nor U2014 (N_2014,N_1816,N_1636);
xor U2015 (N_2015,N_1641,N_1878);
nor U2016 (N_2016,N_1642,N_1649);
xnor U2017 (N_2017,N_1669,N_1841);
nor U2018 (N_2018,N_1606,N_1758);
nor U2019 (N_2019,N_1813,N_1711);
nand U2020 (N_2020,N_1767,N_1599);
nand U2021 (N_2021,N_1988,N_1920);
or U2022 (N_2022,N_1671,N_1709);
nand U2023 (N_2023,N_1875,N_1561);
nand U2024 (N_2024,N_1865,N_1862);
xnor U2025 (N_2025,N_1890,N_1924);
or U2026 (N_2026,N_1622,N_1938);
xnor U2027 (N_2027,N_1684,N_1777);
and U2028 (N_2028,N_1967,N_1661);
xor U2029 (N_2029,N_1978,N_1888);
nand U2030 (N_2030,N_1630,N_1830);
xnor U2031 (N_2031,N_1743,N_1680);
nor U2032 (N_2032,N_1632,N_1797);
xnor U2033 (N_2033,N_1785,N_1626);
nand U2034 (N_2034,N_1523,N_1932);
nand U2035 (N_2035,N_1745,N_1952);
or U2036 (N_2036,N_1717,N_1853);
or U2037 (N_2037,N_1735,N_1819);
nor U2038 (N_2038,N_1686,N_1627);
nor U2039 (N_2039,N_1915,N_1935);
or U2040 (N_2040,N_1927,N_1727);
and U2041 (N_2041,N_1585,N_1665);
or U2042 (N_2042,N_1538,N_1838);
and U2043 (N_2043,N_1729,N_1775);
or U2044 (N_2044,N_1748,N_1590);
nand U2045 (N_2045,N_1675,N_1774);
nand U2046 (N_2046,N_1866,N_1605);
nor U2047 (N_2047,N_1965,N_1895);
xnor U2048 (N_2048,N_1571,N_1576);
nand U2049 (N_2049,N_1874,N_1608);
nor U2050 (N_2050,N_1582,N_1908);
nand U2051 (N_2051,N_1826,N_1871);
xor U2052 (N_2052,N_1714,N_1963);
nor U2053 (N_2053,N_1739,N_1614);
xor U2054 (N_2054,N_1740,N_1609);
or U2055 (N_2055,N_1956,N_1589);
nand U2056 (N_2056,N_1601,N_1995);
and U2057 (N_2057,N_1966,N_1870);
nand U2058 (N_2058,N_1771,N_1668);
nor U2059 (N_2059,N_1986,N_1696);
and U2060 (N_2060,N_1733,N_1793);
xor U2061 (N_2061,N_1896,N_1531);
or U2062 (N_2062,N_1579,N_1863);
xnor U2063 (N_2063,N_1512,N_1984);
nor U2064 (N_2064,N_1980,N_1509);
or U2065 (N_2065,N_1683,N_1603);
nand U2066 (N_2066,N_1719,N_1891);
xnor U2067 (N_2067,N_1919,N_1573);
nand U2068 (N_2068,N_1581,N_1882);
or U2069 (N_2069,N_1744,N_1558);
or U2070 (N_2070,N_1840,N_1913);
or U2071 (N_2071,N_1993,N_1712);
xor U2072 (N_2072,N_1543,N_1886);
nand U2073 (N_2073,N_1689,N_1849);
nand U2074 (N_2074,N_1836,N_1947);
or U2075 (N_2075,N_1945,N_1657);
xor U2076 (N_2076,N_1968,N_1726);
or U2077 (N_2077,N_1818,N_1842);
or U2078 (N_2078,N_1699,N_1832);
nor U2079 (N_2079,N_1939,N_1801);
and U2080 (N_2080,N_1950,N_1916);
or U2081 (N_2081,N_1904,N_1898);
nand U2082 (N_2082,N_1667,N_1994);
or U2083 (N_2083,N_1613,N_1944);
or U2084 (N_2084,N_1911,N_1542);
xor U2085 (N_2085,N_1855,N_1765);
or U2086 (N_2086,N_1781,N_1833);
nand U2087 (N_2087,N_1828,N_1577);
nor U2088 (N_2088,N_1565,N_1746);
and U2089 (N_2089,N_1715,N_1788);
or U2090 (N_2090,N_1867,N_1502);
xnor U2091 (N_2091,N_1852,N_1780);
nand U2092 (N_2092,N_1604,N_1631);
nand U2093 (N_2093,N_1755,N_1646);
and U2094 (N_2094,N_1902,N_1670);
xnor U2095 (N_2095,N_1551,N_1698);
nand U2096 (N_2096,N_1940,N_1564);
and U2097 (N_2097,N_1821,N_1666);
nand U2098 (N_2098,N_1989,N_1539);
xnor U2099 (N_2099,N_1883,N_1650);
nand U2100 (N_2100,N_1625,N_1555);
and U2101 (N_2101,N_1600,N_1757);
nand U2102 (N_2102,N_1998,N_1843);
nor U2103 (N_2103,N_1591,N_1559);
and U2104 (N_2104,N_1854,N_1706);
xnor U2105 (N_2105,N_1762,N_1595);
and U2106 (N_2106,N_1638,N_1876);
nand U2107 (N_2107,N_1955,N_1960);
or U2108 (N_2108,N_1972,N_1766);
nand U2109 (N_2109,N_1540,N_1805);
nor U2110 (N_2110,N_1574,N_1628);
nor U2111 (N_2111,N_1977,N_1872);
and U2112 (N_2112,N_1682,N_1934);
xnor U2113 (N_2113,N_1672,N_1501);
nor U2114 (N_2114,N_1537,N_1701);
and U2115 (N_2115,N_1697,N_1545);
and U2116 (N_2116,N_1514,N_1957);
and U2117 (N_2117,N_1524,N_1592);
or U2118 (N_2118,N_1897,N_1931);
or U2119 (N_2119,N_1648,N_1894);
and U2120 (N_2120,N_1983,N_1962);
nor U2121 (N_2121,N_1930,N_1784);
xor U2122 (N_2122,N_1522,N_1885);
and U2123 (N_2123,N_1829,N_1789);
nand U2124 (N_2124,N_1593,N_1663);
nor U2125 (N_2125,N_1844,N_1827);
or U2126 (N_2126,N_1804,N_1644);
and U2127 (N_2127,N_1570,N_1519);
nand U2128 (N_2128,N_1583,N_1760);
or U2129 (N_2129,N_1679,N_1685);
xor U2130 (N_2130,N_1823,N_1742);
nand U2131 (N_2131,N_1710,N_1937);
or U2132 (N_2132,N_1792,N_1612);
and U2133 (N_2133,N_1508,N_1580);
and U2134 (N_2134,N_1552,N_1700);
xor U2135 (N_2135,N_1856,N_1861);
or U2136 (N_2136,N_1521,N_1562);
or U2137 (N_2137,N_1594,N_1702);
nand U2138 (N_2138,N_1791,N_1639);
nor U2139 (N_2139,N_1811,N_1835);
nand U2140 (N_2140,N_1751,N_1812);
or U2141 (N_2141,N_1921,N_1503);
xor U2142 (N_2142,N_1554,N_1624);
nand U2143 (N_2143,N_1694,N_1730);
nor U2144 (N_2144,N_1598,N_1929);
xnor U2145 (N_2145,N_1526,N_1553);
nand U2146 (N_2146,N_1620,N_1951);
nor U2147 (N_2147,N_1759,N_1810);
and U2148 (N_2148,N_1587,N_1942);
or U2149 (N_2149,N_1954,N_1949);
nand U2150 (N_2150,N_1786,N_1907);
and U2151 (N_2151,N_1659,N_1511);
and U2152 (N_2152,N_1518,N_1504);
nor U2153 (N_2153,N_1825,N_1795);
nor U2154 (N_2154,N_1505,N_1990);
and U2155 (N_2155,N_1873,N_1536);
nand U2156 (N_2156,N_1909,N_1618);
or U2157 (N_2157,N_1704,N_1506);
or U2158 (N_2158,N_1941,N_1928);
nand U2159 (N_2159,N_1681,N_1851);
nor U2160 (N_2160,N_1658,N_1900);
nand U2161 (N_2161,N_1633,N_1987);
and U2162 (N_2162,N_1999,N_1567);
and U2163 (N_2163,N_1691,N_1814);
nor U2164 (N_2164,N_1747,N_1640);
and U2165 (N_2165,N_1837,N_1721);
and U2166 (N_2166,N_1899,N_1728);
or U2167 (N_2167,N_1926,N_1936);
nand U2168 (N_2168,N_1959,N_1857);
nor U2169 (N_2169,N_1834,N_1779);
nand U2170 (N_2170,N_1586,N_1991);
and U2171 (N_2171,N_1724,N_1877);
xor U2172 (N_2172,N_1806,N_1718);
and U2173 (N_2173,N_1656,N_1845);
and U2174 (N_2174,N_1848,N_1754);
and U2175 (N_2175,N_1892,N_1881);
nand U2176 (N_2176,N_1527,N_1973);
xor U2177 (N_2177,N_1693,N_1850);
nand U2178 (N_2178,N_1803,N_1645);
or U2179 (N_2179,N_1776,N_1708);
nand U2180 (N_2180,N_1615,N_1783);
nor U2181 (N_2181,N_1953,N_1922);
and U2182 (N_2182,N_1981,N_1546);
and U2183 (N_2183,N_1749,N_1790);
nand U2184 (N_2184,N_1510,N_1532);
and U2185 (N_2185,N_1914,N_1859);
xor U2186 (N_2186,N_1596,N_1884);
or U2187 (N_2187,N_1687,N_1549);
or U2188 (N_2188,N_1794,N_1500);
or U2189 (N_2189,N_1879,N_1808);
xnor U2190 (N_2190,N_1597,N_1720);
nand U2191 (N_2191,N_1906,N_1617);
or U2192 (N_2192,N_1846,N_1800);
nor U2193 (N_2193,N_1655,N_1918);
xnor U2194 (N_2194,N_1887,N_1541);
nand U2195 (N_2195,N_1917,N_1548);
nand U2196 (N_2196,N_1705,N_1572);
and U2197 (N_2197,N_1753,N_1773);
xnor U2198 (N_2198,N_1544,N_1889);
and U2199 (N_2199,N_1737,N_1992);
or U2200 (N_2200,N_1933,N_1893);
nor U2201 (N_2201,N_1578,N_1847);
nor U2202 (N_2202,N_1860,N_1725);
nand U2203 (N_2203,N_1634,N_1815);
nor U2204 (N_2204,N_1910,N_1677);
xnor U2205 (N_2205,N_1764,N_1695);
and U2206 (N_2206,N_1864,N_1652);
or U2207 (N_2207,N_1588,N_1778);
nand U2208 (N_2208,N_1741,N_1557);
and U2209 (N_2209,N_1654,N_1903);
nor U2210 (N_2210,N_1770,N_1964);
nor U2211 (N_2211,N_1678,N_1550);
nor U2212 (N_2212,N_1707,N_1517);
nand U2213 (N_2213,N_1817,N_1607);
nor U2214 (N_2214,N_1868,N_1621);
nand U2215 (N_2215,N_1690,N_1584);
and U2216 (N_2216,N_1736,N_1525);
nand U2217 (N_2217,N_1796,N_1782);
nor U2218 (N_2218,N_1529,N_1653);
or U2219 (N_2219,N_1647,N_1905);
nor U2220 (N_2220,N_1809,N_1869);
nand U2221 (N_2221,N_1662,N_1901);
and U2222 (N_2222,N_1970,N_1768);
xor U2223 (N_2223,N_1560,N_1769);
nor U2224 (N_2224,N_1831,N_1530);
and U2225 (N_2225,N_1660,N_1822);
and U2226 (N_2226,N_1772,N_1975);
or U2227 (N_2227,N_1982,N_1799);
nand U2228 (N_2228,N_1507,N_1958);
xor U2229 (N_2229,N_1732,N_1563);
or U2230 (N_2230,N_1703,N_1713);
nand U2231 (N_2231,N_1569,N_1716);
nand U2232 (N_2232,N_1997,N_1839);
or U2233 (N_2233,N_1547,N_1946);
nor U2234 (N_2234,N_1761,N_1763);
or U2235 (N_2235,N_1798,N_1623);
or U2236 (N_2236,N_1651,N_1756);
xor U2237 (N_2237,N_1673,N_1750);
nor U2238 (N_2238,N_1610,N_1616);
nor U2239 (N_2239,N_1534,N_1611);
and U2240 (N_2240,N_1974,N_1688);
xnor U2241 (N_2241,N_1676,N_1528);
nor U2242 (N_2242,N_1515,N_1513);
xnor U2243 (N_2243,N_1516,N_1787);
nand U2244 (N_2244,N_1948,N_1752);
or U2245 (N_2245,N_1575,N_1723);
xnor U2246 (N_2246,N_1637,N_1692);
and U2247 (N_2247,N_1802,N_1664);
and U2248 (N_2248,N_1824,N_1520);
nor U2249 (N_2249,N_1971,N_1535);
or U2250 (N_2250,N_1611,N_1549);
nor U2251 (N_2251,N_1784,N_1941);
and U2252 (N_2252,N_1754,N_1565);
nand U2253 (N_2253,N_1928,N_1997);
nor U2254 (N_2254,N_1563,N_1741);
and U2255 (N_2255,N_1924,N_1867);
nand U2256 (N_2256,N_1924,N_1970);
nor U2257 (N_2257,N_1636,N_1691);
nand U2258 (N_2258,N_1839,N_1771);
nand U2259 (N_2259,N_1857,N_1659);
nor U2260 (N_2260,N_1554,N_1724);
or U2261 (N_2261,N_1604,N_1960);
and U2262 (N_2262,N_1957,N_1976);
or U2263 (N_2263,N_1683,N_1977);
nor U2264 (N_2264,N_1714,N_1892);
xnor U2265 (N_2265,N_1525,N_1622);
or U2266 (N_2266,N_1682,N_1727);
xnor U2267 (N_2267,N_1947,N_1626);
nand U2268 (N_2268,N_1980,N_1944);
nor U2269 (N_2269,N_1647,N_1540);
nand U2270 (N_2270,N_1827,N_1574);
nand U2271 (N_2271,N_1577,N_1992);
xor U2272 (N_2272,N_1579,N_1866);
and U2273 (N_2273,N_1505,N_1604);
xor U2274 (N_2274,N_1585,N_1971);
and U2275 (N_2275,N_1902,N_1762);
or U2276 (N_2276,N_1582,N_1764);
or U2277 (N_2277,N_1676,N_1774);
xnor U2278 (N_2278,N_1902,N_1823);
nand U2279 (N_2279,N_1688,N_1882);
and U2280 (N_2280,N_1787,N_1581);
nor U2281 (N_2281,N_1512,N_1908);
or U2282 (N_2282,N_1775,N_1650);
nor U2283 (N_2283,N_1731,N_1925);
or U2284 (N_2284,N_1717,N_1799);
or U2285 (N_2285,N_1741,N_1801);
or U2286 (N_2286,N_1834,N_1652);
or U2287 (N_2287,N_1719,N_1661);
nand U2288 (N_2288,N_1849,N_1857);
and U2289 (N_2289,N_1579,N_1609);
or U2290 (N_2290,N_1711,N_1644);
nor U2291 (N_2291,N_1776,N_1972);
xor U2292 (N_2292,N_1856,N_1806);
nor U2293 (N_2293,N_1738,N_1871);
or U2294 (N_2294,N_1877,N_1770);
xnor U2295 (N_2295,N_1646,N_1979);
nand U2296 (N_2296,N_1890,N_1556);
nand U2297 (N_2297,N_1914,N_1955);
or U2298 (N_2298,N_1838,N_1772);
xnor U2299 (N_2299,N_1677,N_1662);
or U2300 (N_2300,N_1548,N_1568);
xnor U2301 (N_2301,N_1626,N_1759);
or U2302 (N_2302,N_1931,N_1856);
nor U2303 (N_2303,N_1633,N_1858);
and U2304 (N_2304,N_1801,N_1643);
nor U2305 (N_2305,N_1881,N_1724);
nor U2306 (N_2306,N_1770,N_1940);
nand U2307 (N_2307,N_1749,N_1568);
nor U2308 (N_2308,N_1674,N_1871);
nand U2309 (N_2309,N_1726,N_1624);
or U2310 (N_2310,N_1674,N_1767);
nor U2311 (N_2311,N_1510,N_1781);
and U2312 (N_2312,N_1758,N_1594);
or U2313 (N_2313,N_1687,N_1603);
nand U2314 (N_2314,N_1598,N_1607);
and U2315 (N_2315,N_1791,N_1680);
nand U2316 (N_2316,N_1677,N_1853);
nand U2317 (N_2317,N_1983,N_1550);
nand U2318 (N_2318,N_1623,N_1524);
xnor U2319 (N_2319,N_1962,N_1616);
and U2320 (N_2320,N_1711,N_1568);
nor U2321 (N_2321,N_1683,N_1886);
xnor U2322 (N_2322,N_1835,N_1648);
nand U2323 (N_2323,N_1625,N_1937);
nor U2324 (N_2324,N_1703,N_1867);
nor U2325 (N_2325,N_1543,N_1583);
or U2326 (N_2326,N_1752,N_1518);
xor U2327 (N_2327,N_1626,N_1819);
and U2328 (N_2328,N_1673,N_1744);
nand U2329 (N_2329,N_1956,N_1812);
and U2330 (N_2330,N_1782,N_1557);
nor U2331 (N_2331,N_1778,N_1839);
nor U2332 (N_2332,N_1788,N_1997);
nor U2333 (N_2333,N_1604,N_1514);
or U2334 (N_2334,N_1829,N_1880);
or U2335 (N_2335,N_1530,N_1568);
and U2336 (N_2336,N_1705,N_1818);
and U2337 (N_2337,N_1643,N_1795);
or U2338 (N_2338,N_1917,N_1936);
or U2339 (N_2339,N_1629,N_1541);
nand U2340 (N_2340,N_1833,N_1568);
or U2341 (N_2341,N_1535,N_1833);
xnor U2342 (N_2342,N_1559,N_1865);
nor U2343 (N_2343,N_1836,N_1901);
nand U2344 (N_2344,N_1648,N_1603);
nand U2345 (N_2345,N_1727,N_1582);
xor U2346 (N_2346,N_1808,N_1644);
nor U2347 (N_2347,N_1576,N_1510);
xnor U2348 (N_2348,N_1875,N_1546);
or U2349 (N_2349,N_1610,N_1963);
and U2350 (N_2350,N_1827,N_1580);
and U2351 (N_2351,N_1570,N_1930);
nand U2352 (N_2352,N_1610,N_1692);
and U2353 (N_2353,N_1611,N_1941);
nor U2354 (N_2354,N_1864,N_1935);
xnor U2355 (N_2355,N_1827,N_1882);
or U2356 (N_2356,N_1856,N_1686);
and U2357 (N_2357,N_1825,N_1794);
or U2358 (N_2358,N_1828,N_1982);
nor U2359 (N_2359,N_1713,N_1505);
and U2360 (N_2360,N_1767,N_1996);
or U2361 (N_2361,N_1755,N_1601);
or U2362 (N_2362,N_1932,N_1835);
nor U2363 (N_2363,N_1694,N_1932);
and U2364 (N_2364,N_1971,N_1566);
and U2365 (N_2365,N_1507,N_1594);
nor U2366 (N_2366,N_1805,N_1818);
nand U2367 (N_2367,N_1870,N_1936);
or U2368 (N_2368,N_1612,N_1589);
and U2369 (N_2369,N_1973,N_1532);
nand U2370 (N_2370,N_1862,N_1815);
and U2371 (N_2371,N_1941,N_1700);
xor U2372 (N_2372,N_1947,N_1537);
xor U2373 (N_2373,N_1897,N_1663);
xnor U2374 (N_2374,N_1746,N_1795);
or U2375 (N_2375,N_1766,N_1929);
nand U2376 (N_2376,N_1615,N_1510);
or U2377 (N_2377,N_1642,N_1677);
nand U2378 (N_2378,N_1532,N_1660);
nor U2379 (N_2379,N_1950,N_1765);
and U2380 (N_2380,N_1685,N_1584);
xnor U2381 (N_2381,N_1633,N_1639);
nand U2382 (N_2382,N_1520,N_1914);
xnor U2383 (N_2383,N_1542,N_1599);
xor U2384 (N_2384,N_1637,N_1845);
nor U2385 (N_2385,N_1706,N_1908);
and U2386 (N_2386,N_1502,N_1823);
xor U2387 (N_2387,N_1867,N_1591);
nor U2388 (N_2388,N_1782,N_1719);
nand U2389 (N_2389,N_1533,N_1788);
xor U2390 (N_2390,N_1838,N_1804);
xor U2391 (N_2391,N_1614,N_1645);
and U2392 (N_2392,N_1682,N_1515);
or U2393 (N_2393,N_1522,N_1627);
and U2394 (N_2394,N_1744,N_1840);
nor U2395 (N_2395,N_1661,N_1588);
and U2396 (N_2396,N_1815,N_1838);
or U2397 (N_2397,N_1591,N_1640);
nor U2398 (N_2398,N_1519,N_1535);
and U2399 (N_2399,N_1897,N_1657);
or U2400 (N_2400,N_1744,N_1735);
nand U2401 (N_2401,N_1643,N_1784);
nand U2402 (N_2402,N_1984,N_1985);
or U2403 (N_2403,N_1759,N_1693);
nor U2404 (N_2404,N_1631,N_1663);
or U2405 (N_2405,N_1996,N_1822);
or U2406 (N_2406,N_1946,N_1864);
xnor U2407 (N_2407,N_1962,N_1719);
and U2408 (N_2408,N_1943,N_1984);
or U2409 (N_2409,N_1769,N_1826);
nor U2410 (N_2410,N_1640,N_1913);
xor U2411 (N_2411,N_1831,N_1579);
nor U2412 (N_2412,N_1618,N_1961);
and U2413 (N_2413,N_1604,N_1519);
and U2414 (N_2414,N_1701,N_1589);
and U2415 (N_2415,N_1918,N_1575);
or U2416 (N_2416,N_1630,N_1853);
or U2417 (N_2417,N_1973,N_1639);
xnor U2418 (N_2418,N_1516,N_1894);
nor U2419 (N_2419,N_1584,N_1877);
nor U2420 (N_2420,N_1604,N_1577);
xor U2421 (N_2421,N_1802,N_1591);
and U2422 (N_2422,N_1757,N_1561);
nand U2423 (N_2423,N_1637,N_1996);
and U2424 (N_2424,N_1929,N_1949);
nor U2425 (N_2425,N_1515,N_1582);
and U2426 (N_2426,N_1657,N_1723);
nand U2427 (N_2427,N_1934,N_1507);
xnor U2428 (N_2428,N_1681,N_1863);
or U2429 (N_2429,N_1948,N_1514);
xor U2430 (N_2430,N_1891,N_1713);
or U2431 (N_2431,N_1539,N_1701);
nor U2432 (N_2432,N_1745,N_1924);
nand U2433 (N_2433,N_1517,N_1532);
nor U2434 (N_2434,N_1989,N_1927);
and U2435 (N_2435,N_1824,N_1517);
or U2436 (N_2436,N_1957,N_1962);
and U2437 (N_2437,N_1529,N_1701);
xor U2438 (N_2438,N_1776,N_1865);
or U2439 (N_2439,N_1899,N_1898);
xnor U2440 (N_2440,N_1726,N_1978);
xor U2441 (N_2441,N_1711,N_1680);
nor U2442 (N_2442,N_1562,N_1700);
nor U2443 (N_2443,N_1661,N_1855);
or U2444 (N_2444,N_1891,N_1992);
nor U2445 (N_2445,N_1589,N_1703);
nand U2446 (N_2446,N_1894,N_1971);
nor U2447 (N_2447,N_1972,N_1911);
nor U2448 (N_2448,N_1528,N_1877);
nand U2449 (N_2449,N_1847,N_1909);
or U2450 (N_2450,N_1956,N_1651);
and U2451 (N_2451,N_1887,N_1695);
or U2452 (N_2452,N_1524,N_1573);
nand U2453 (N_2453,N_1585,N_1560);
or U2454 (N_2454,N_1556,N_1662);
nand U2455 (N_2455,N_1637,N_1932);
and U2456 (N_2456,N_1991,N_1579);
and U2457 (N_2457,N_1991,N_1821);
and U2458 (N_2458,N_1881,N_1968);
or U2459 (N_2459,N_1718,N_1725);
nand U2460 (N_2460,N_1952,N_1789);
nand U2461 (N_2461,N_1523,N_1521);
or U2462 (N_2462,N_1590,N_1998);
and U2463 (N_2463,N_1857,N_1575);
xnor U2464 (N_2464,N_1682,N_1648);
xor U2465 (N_2465,N_1706,N_1949);
and U2466 (N_2466,N_1897,N_1915);
xnor U2467 (N_2467,N_1905,N_1951);
or U2468 (N_2468,N_1664,N_1954);
xnor U2469 (N_2469,N_1996,N_1970);
or U2470 (N_2470,N_1981,N_1755);
nand U2471 (N_2471,N_1768,N_1875);
and U2472 (N_2472,N_1648,N_1944);
and U2473 (N_2473,N_1544,N_1934);
nand U2474 (N_2474,N_1983,N_1865);
and U2475 (N_2475,N_1572,N_1511);
and U2476 (N_2476,N_1579,N_1671);
nand U2477 (N_2477,N_1746,N_1991);
nor U2478 (N_2478,N_1805,N_1629);
and U2479 (N_2479,N_1597,N_1944);
nand U2480 (N_2480,N_1819,N_1505);
xor U2481 (N_2481,N_1821,N_1866);
and U2482 (N_2482,N_1799,N_1644);
nor U2483 (N_2483,N_1868,N_1926);
nand U2484 (N_2484,N_1505,N_1878);
nor U2485 (N_2485,N_1591,N_1682);
nor U2486 (N_2486,N_1523,N_1771);
and U2487 (N_2487,N_1819,N_1899);
nand U2488 (N_2488,N_1616,N_1919);
nand U2489 (N_2489,N_1545,N_1999);
nand U2490 (N_2490,N_1753,N_1675);
and U2491 (N_2491,N_1947,N_1900);
or U2492 (N_2492,N_1716,N_1626);
or U2493 (N_2493,N_1710,N_1805);
nor U2494 (N_2494,N_1775,N_1537);
nor U2495 (N_2495,N_1762,N_1525);
xnor U2496 (N_2496,N_1910,N_1500);
or U2497 (N_2497,N_1845,N_1915);
or U2498 (N_2498,N_1839,N_1563);
or U2499 (N_2499,N_1655,N_1797);
or U2500 (N_2500,N_2492,N_2058);
nand U2501 (N_2501,N_2246,N_2237);
xor U2502 (N_2502,N_2038,N_2366);
nor U2503 (N_2503,N_2461,N_2108);
or U2504 (N_2504,N_2229,N_2358);
and U2505 (N_2505,N_2422,N_2399);
or U2506 (N_2506,N_2306,N_2021);
and U2507 (N_2507,N_2334,N_2064);
nand U2508 (N_2508,N_2078,N_2485);
nor U2509 (N_2509,N_2091,N_2333);
and U2510 (N_2510,N_2070,N_2139);
xnor U2511 (N_2511,N_2228,N_2127);
and U2512 (N_2512,N_2392,N_2030);
nand U2513 (N_2513,N_2075,N_2217);
nand U2514 (N_2514,N_2491,N_2288);
nor U2515 (N_2515,N_2293,N_2397);
xor U2516 (N_2516,N_2478,N_2322);
and U2517 (N_2517,N_2088,N_2136);
nor U2518 (N_2518,N_2182,N_2481);
and U2519 (N_2519,N_2126,N_2351);
nor U2520 (N_2520,N_2313,N_2028);
nor U2521 (N_2521,N_2036,N_2227);
nand U2522 (N_2522,N_2270,N_2157);
xor U2523 (N_2523,N_2235,N_2455);
or U2524 (N_2524,N_2381,N_2471);
xor U2525 (N_2525,N_2209,N_2301);
and U2526 (N_2526,N_2375,N_2224);
nand U2527 (N_2527,N_2155,N_2460);
xor U2528 (N_2528,N_2051,N_2158);
nand U2529 (N_2529,N_2274,N_2403);
nor U2530 (N_2530,N_2465,N_2437);
xnor U2531 (N_2531,N_2286,N_2277);
or U2532 (N_2532,N_2247,N_2014);
xor U2533 (N_2533,N_2476,N_2410);
xor U2534 (N_2534,N_2242,N_2419);
or U2535 (N_2535,N_2303,N_2206);
xnor U2536 (N_2536,N_2102,N_2362);
nor U2537 (N_2537,N_2211,N_2387);
or U2538 (N_2538,N_2119,N_2386);
nor U2539 (N_2539,N_2141,N_2407);
xor U2540 (N_2540,N_2121,N_2384);
or U2541 (N_2541,N_2018,N_2068);
nand U2542 (N_2542,N_2061,N_2077);
nor U2543 (N_2543,N_2219,N_2218);
xnor U2544 (N_2544,N_2198,N_2369);
nor U2545 (N_2545,N_2200,N_2100);
nand U2546 (N_2546,N_2111,N_2166);
nor U2547 (N_2547,N_2454,N_2340);
or U2548 (N_2548,N_2378,N_2368);
xor U2549 (N_2549,N_2412,N_2231);
nand U2550 (N_2550,N_2284,N_2307);
nand U2551 (N_2551,N_2025,N_2353);
or U2552 (N_2552,N_2262,N_2453);
nor U2553 (N_2553,N_2201,N_2110);
nor U2554 (N_2554,N_2269,N_2092);
and U2555 (N_2555,N_2005,N_2096);
or U2556 (N_2556,N_2440,N_2469);
or U2557 (N_2557,N_2052,N_2470);
and U2558 (N_2558,N_2196,N_2221);
nand U2559 (N_2559,N_2299,N_2199);
nor U2560 (N_2560,N_2330,N_2389);
nor U2561 (N_2561,N_2382,N_2148);
nor U2562 (N_2562,N_2281,N_2029);
nor U2563 (N_2563,N_2167,N_2041);
and U2564 (N_2564,N_2006,N_2483);
xor U2565 (N_2565,N_2304,N_2479);
and U2566 (N_2566,N_2486,N_2011);
xnor U2567 (N_2567,N_2035,N_2054);
nor U2568 (N_2568,N_2271,N_2405);
nor U2569 (N_2569,N_2464,N_2423);
nor U2570 (N_2570,N_2050,N_2380);
nand U2571 (N_2571,N_2310,N_2365);
or U2572 (N_2572,N_2335,N_2193);
or U2573 (N_2573,N_2426,N_2215);
and U2574 (N_2574,N_2431,N_2189);
nor U2575 (N_2575,N_2266,N_2142);
and U2576 (N_2576,N_2482,N_2402);
or U2577 (N_2577,N_2245,N_2095);
nand U2578 (N_2578,N_2164,N_2255);
xor U2579 (N_2579,N_2261,N_2116);
nand U2580 (N_2580,N_2249,N_2377);
nor U2581 (N_2581,N_2001,N_2241);
nand U2582 (N_2582,N_2212,N_2390);
nor U2583 (N_2583,N_2393,N_2012);
or U2584 (N_2584,N_2066,N_2207);
nor U2585 (N_2585,N_2019,N_2364);
nand U2586 (N_2586,N_2298,N_2106);
nand U2587 (N_2587,N_2093,N_2244);
or U2588 (N_2588,N_2177,N_2394);
or U2589 (N_2589,N_2406,N_2002);
xor U2590 (N_2590,N_2357,N_2162);
and U2591 (N_2591,N_2067,N_2183);
xnor U2592 (N_2592,N_2133,N_2250);
or U2593 (N_2593,N_2264,N_2265);
nand U2594 (N_2594,N_2278,N_2473);
or U2595 (N_2595,N_2466,N_2356);
nor U2596 (N_2596,N_2230,N_2020);
or U2597 (N_2597,N_2395,N_2131);
xnor U2598 (N_2598,N_2056,N_2226);
and U2599 (N_2599,N_2272,N_2371);
xor U2600 (N_2600,N_2031,N_2022);
or U2601 (N_2601,N_2101,N_2490);
nor U2602 (N_2602,N_2083,N_2442);
nor U2603 (N_2603,N_2147,N_2034);
nand U2604 (N_2604,N_2263,N_2416);
or U2605 (N_2605,N_2370,N_2169);
and U2606 (N_2606,N_2007,N_2421);
xnor U2607 (N_2607,N_2239,N_2458);
xnor U2608 (N_2608,N_2346,N_2477);
xnor U2609 (N_2609,N_2452,N_2178);
nor U2610 (N_2610,N_2137,N_2396);
nand U2611 (N_2611,N_2062,N_2444);
nand U2612 (N_2612,N_2191,N_2023);
or U2613 (N_2613,N_2385,N_2287);
nand U2614 (N_2614,N_2117,N_2197);
nor U2615 (N_2615,N_2360,N_2383);
nor U2616 (N_2616,N_2309,N_2190);
nand U2617 (N_2617,N_2374,N_2071);
and U2618 (N_2618,N_2185,N_2257);
or U2619 (N_2619,N_2123,N_2339);
nand U2620 (N_2620,N_2295,N_2084);
or U2621 (N_2621,N_2016,N_2172);
xor U2622 (N_2622,N_2240,N_2079);
xnor U2623 (N_2623,N_2149,N_2194);
nor U2624 (N_2624,N_2338,N_2128);
nand U2625 (N_2625,N_2325,N_2176);
and U2626 (N_2626,N_2138,N_2109);
nor U2627 (N_2627,N_2499,N_2343);
or U2628 (N_2628,N_2152,N_2163);
xor U2629 (N_2629,N_2049,N_2180);
xor U2630 (N_2630,N_2174,N_2297);
and U2631 (N_2631,N_2498,N_2008);
or U2632 (N_2632,N_2175,N_2063);
nor U2633 (N_2633,N_2415,N_2398);
nor U2634 (N_2634,N_2216,N_2044);
and U2635 (N_2635,N_2355,N_2475);
nor U2636 (N_2636,N_2292,N_2424);
nand U2637 (N_2637,N_2009,N_2451);
and U2638 (N_2638,N_2140,N_2420);
xnor U2639 (N_2639,N_2143,N_2457);
xor U2640 (N_2640,N_2214,N_2130);
and U2641 (N_2641,N_2291,N_2081);
or U2642 (N_2642,N_2345,N_2436);
and U2643 (N_2643,N_2379,N_2236);
nor U2644 (N_2644,N_2113,N_2296);
nand U2645 (N_2645,N_2072,N_2042);
nor U2646 (N_2646,N_2497,N_2459);
and U2647 (N_2647,N_2429,N_2467);
or U2648 (N_2648,N_2258,N_2047);
nand U2649 (N_2649,N_2487,N_2474);
and U2650 (N_2650,N_2275,N_2048);
nand U2651 (N_2651,N_2060,N_2074);
nor U2652 (N_2652,N_2408,N_2238);
and U2653 (N_2653,N_2332,N_2268);
nand U2654 (N_2654,N_2188,N_2192);
or U2655 (N_2655,N_2220,N_2326);
xnor U2656 (N_2656,N_2181,N_2449);
xnor U2657 (N_2657,N_2210,N_2195);
nand U2658 (N_2658,N_2114,N_2129);
or U2659 (N_2659,N_2087,N_2225);
and U2660 (N_2660,N_2057,N_2443);
nor U2661 (N_2661,N_2279,N_2352);
or U2662 (N_2662,N_2373,N_2363);
and U2663 (N_2663,N_2124,N_2232);
or U2664 (N_2664,N_2289,N_2341);
nand U2665 (N_2665,N_2187,N_2348);
and U2666 (N_2666,N_2097,N_2003);
nand U2667 (N_2667,N_2076,N_2305);
or U2668 (N_2668,N_2488,N_2361);
nand U2669 (N_2669,N_2099,N_2103);
and U2670 (N_2670,N_2290,N_2118);
nor U2671 (N_2671,N_2145,N_2135);
nor U2672 (N_2672,N_2480,N_2089);
xor U2673 (N_2673,N_2132,N_2337);
xnor U2674 (N_2674,N_2010,N_2046);
nand U2675 (N_2675,N_2125,N_2350);
xnor U2676 (N_2676,N_2349,N_2248);
or U2677 (N_2677,N_2401,N_2446);
nand U2678 (N_2678,N_2256,N_2045);
xnor U2679 (N_2679,N_2017,N_2086);
or U2680 (N_2680,N_2202,N_2328);
nand U2681 (N_2681,N_2445,N_2065);
nand U2682 (N_2682,N_2462,N_2425);
or U2683 (N_2683,N_2324,N_2153);
nand U2684 (N_2684,N_2347,N_2427);
and U2685 (N_2685,N_2186,N_2450);
nand U2686 (N_2686,N_2094,N_2300);
nand U2687 (N_2687,N_2260,N_2205);
xor U2688 (N_2688,N_2073,N_2168);
xnor U2689 (N_2689,N_2434,N_2098);
and U2690 (N_2690,N_2160,N_2043);
or U2691 (N_2691,N_2439,N_2463);
and U2692 (N_2692,N_2024,N_2000);
xor U2693 (N_2693,N_2321,N_2122);
xnor U2694 (N_2694,N_2468,N_2282);
or U2695 (N_2695,N_2418,N_2204);
nand U2696 (N_2696,N_2253,N_2302);
nor U2697 (N_2697,N_2312,N_2400);
nor U2698 (N_2698,N_2090,N_2448);
nand U2699 (N_2699,N_2134,N_2311);
xnor U2700 (N_2700,N_2319,N_2161);
nand U2701 (N_2701,N_2376,N_2150);
xor U2702 (N_2702,N_2359,N_2069);
and U2703 (N_2703,N_2285,N_2409);
or U2704 (N_2704,N_2489,N_2223);
and U2705 (N_2705,N_2280,N_2179);
or U2706 (N_2706,N_2495,N_2233);
xor U2707 (N_2707,N_2115,N_2435);
nor U2708 (N_2708,N_2170,N_2027);
and U2709 (N_2709,N_2494,N_2354);
xor U2710 (N_2710,N_2203,N_2208);
or U2711 (N_2711,N_2107,N_2294);
or U2712 (N_2712,N_2154,N_2267);
or U2713 (N_2713,N_2404,N_2336);
xor U2714 (N_2714,N_2493,N_2308);
nand U2715 (N_2715,N_2417,N_2414);
nor U2716 (N_2716,N_2173,N_2254);
or U2717 (N_2717,N_2252,N_2441);
and U2718 (N_2718,N_2472,N_2105);
or U2719 (N_2719,N_2430,N_2273);
and U2720 (N_2720,N_2055,N_2320);
xor U2721 (N_2721,N_2428,N_2171);
nor U2722 (N_2722,N_2156,N_2447);
nor U2723 (N_2723,N_2413,N_2411);
nand U2724 (N_2724,N_2331,N_2032);
xor U2725 (N_2725,N_2004,N_2314);
nor U2726 (N_2726,N_2327,N_2080);
or U2727 (N_2727,N_2146,N_2438);
or U2728 (N_2728,N_2317,N_2323);
nor U2729 (N_2729,N_2315,N_2104);
nand U2730 (N_2730,N_2276,N_2165);
or U2731 (N_2731,N_2318,N_2112);
nor U2732 (N_2732,N_2329,N_2433);
nor U2733 (N_2733,N_2151,N_2159);
nor U2734 (N_2734,N_2391,N_2037);
xnor U2735 (N_2735,N_2026,N_2456);
and U2736 (N_2736,N_2484,N_2283);
nor U2737 (N_2737,N_2033,N_2082);
nor U2738 (N_2738,N_2388,N_2496);
and U2739 (N_2739,N_2432,N_2120);
nor U2740 (N_2740,N_2015,N_2013);
xor U2741 (N_2741,N_2059,N_2243);
and U2742 (N_2742,N_2372,N_2342);
nor U2743 (N_2743,N_2039,N_2053);
and U2744 (N_2744,N_2367,N_2222);
nor U2745 (N_2745,N_2184,N_2251);
xor U2746 (N_2746,N_2344,N_2040);
and U2747 (N_2747,N_2213,N_2085);
nand U2748 (N_2748,N_2144,N_2316);
nand U2749 (N_2749,N_2259,N_2234);
xnor U2750 (N_2750,N_2416,N_2034);
nor U2751 (N_2751,N_2040,N_2280);
xor U2752 (N_2752,N_2324,N_2360);
nand U2753 (N_2753,N_2037,N_2249);
xnor U2754 (N_2754,N_2290,N_2033);
nor U2755 (N_2755,N_2140,N_2399);
xor U2756 (N_2756,N_2163,N_2009);
xor U2757 (N_2757,N_2341,N_2104);
or U2758 (N_2758,N_2288,N_2342);
nor U2759 (N_2759,N_2073,N_2493);
and U2760 (N_2760,N_2240,N_2218);
nand U2761 (N_2761,N_2346,N_2445);
and U2762 (N_2762,N_2167,N_2277);
or U2763 (N_2763,N_2258,N_2290);
or U2764 (N_2764,N_2186,N_2180);
and U2765 (N_2765,N_2081,N_2006);
nor U2766 (N_2766,N_2325,N_2358);
nand U2767 (N_2767,N_2084,N_2257);
and U2768 (N_2768,N_2370,N_2251);
and U2769 (N_2769,N_2294,N_2399);
nand U2770 (N_2770,N_2267,N_2025);
and U2771 (N_2771,N_2360,N_2196);
or U2772 (N_2772,N_2292,N_2165);
and U2773 (N_2773,N_2271,N_2412);
or U2774 (N_2774,N_2328,N_2337);
nor U2775 (N_2775,N_2111,N_2092);
xnor U2776 (N_2776,N_2264,N_2448);
or U2777 (N_2777,N_2351,N_2214);
xor U2778 (N_2778,N_2397,N_2146);
nand U2779 (N_2779,N_2064,N_2315);
or U2780 (N_2780,N_2432,N_2260);
nand U2781 (N_2781,N_2126,N_2174);
nand U2782 (N_2782,N_2291,N_2042);
nor U2783 (N_2783,N_2043,N_2145);
xnor U2784 (N_2784,N_2183,N_2487);
nand U2785 (N_2785,N_2093,N_2256);
or U2786 (N_2786,N_2433,N_2089);
nand U2787 (N_2787,N_2126,N_2141);
or U2788 (N_2788,N_2012,N_2277);
xnor U2789 (N_2789,N_2392,N_2295);
nor U2790 (N_2790,N_2262,N_2266);
or U2791 (N_2791,N_2080,N_2002);
nor U2792 (N_2792,N_2142,N_2344);
xor U2793 (N_2793,N_2053,N_2334);
or U2794 (N_2794,N_2090,N_2493);
nor U2795 (N_2795,N_2286,N_2232);
nand U2796 (N_2796,N_2056,N_2292);
nand U2797 (N_2797,N_2185,N_2068);
or U2798 (N_2798,N_2422,N_2017);
xor U2799 (N_2799,N_2190,N_2179);
nand U2800 (N_2800,N_2319,N_2429);
nor U2801 (N_2801,N_2148,N_2268);
xnor U2802 (N_2802,N_2480,N_2250);
or U2803 (N_2803,N_2427,N_2251);
or U2804 (N_2804,N_2184,N_2093);
nand U2805 (N_2805,N_2103,N_2021);
and U2806 (N_2806,N_2155,N_2087);
nor U2807 (N_2807,N_2002,N_2499);
xnor U2808 (N_2808,N_2365,N_2410);
nand U2809 (N_2809,N_2024,N_2243);
or U2810 (N_2810,N_2306,N_2005);
or U2811 (N_2811,N_2307,N_2491);
nand U2812 (N_2812,N_2369,N_2375);
and U2813 (N_2813,N_2449,N_2401);
nand U2814 (N_2814,N_2429,N_2161);
or U2815 (N_2815,N_2142,N_2220);
nor U2816 (N_2816,N_2299,N_2377);
and U2817 (N_2817,N_2297,N_2387);
nand U2818 (N_2818,N_2300,N_2491);
and U2819 (N_2819,N_2474,N_2298);
nand U2820 (N_2820,N_2040,N_2430);
xor U2821 (N_2821,N_2254,N_2031);
nor U2822 (N_2822,N_2259,N_2441);
nand U2823 (N_2823,N_2102,N_2331);
nor U2824 (N_2824,N_2208,N_2188);
or U2825 (N_2825,N_2132,N_2023);
nand U2826 (N_2826,N_2106,N_2343);
nand U2827 (N_2827,N_2448,N_2435);
or U2828 (N_2828,N_2486,N_2196);
or U2829 (N_2829,N_2439,N_2177);
or U2830 (N_2830,N_2042,N_2019);
xor U2831 (N_2831,N_2439,N_2230);
or U2832 (N_2832,N_2445,N_2389);
and U2833 (N_2833,N_2467,N_2477);
nand U2834 (N_2834,N_2357,N_2156);
xor U2835 (N_2835,N_2300,N_2061);
nor U2836 (N_2836,N_2035,N_2008);
and U2837 (N_2837,N_2373,N_2396);
nor U2838 (N_2838,N_2434,N_2114);
nand U2839 (N_2839,N_2032,N_2386);
xnor U2840 (N_2840,N_2114,N_2248);
and U2841 (N_2841,N_2152,N_2373);
xor U2842 (N_2842,N_2475,N_2209);
xnor U2843 (N_2843,N_2328,N_2167);
and U2844 (N_2844,N_2213,N_2455);
nor U2845 (N_2845,N_2468,N_2460);
nor U2846 (N_2846,N_2308,N_2423);
and U2847 (N_2847,N_2234,N_2213);
xor U2848 (N_2848,N_2460,N_2323);
nor U2849 (N_2849,N_2418,N_2353);
and U2850 (N_2850,N_2287,N_2011);
nor U2851 (N_2851,N_2010,N_2433);
and U2852 (N_2852,N_2285,N_2350);
nor U2853 (N_2853,N_2092,N_2139);
xnor U2854 (N_2854,N_2135,N_2078);
and U2855 (N_2855,N_2456,N_2393);
nand U2856 (N_2856,N_2334,N_2263);
nand U2857 (N_2857,N_2052,N_2151);
nand U2858 (N_2858,N_2091,N_2031);
and U2859 (N_2859,N_2102,N_2486);
xnor U2860 (N_2860,N_2024,N_2152);
or U2861 (N_2861,N_2056,N_2123);
nor U2862 (N_2862,N_2052,N_2323);
nand U2863 (N_2863,N_2061,N_2156);
nor U2864 (N_2864,N_2254,N_2399);
xor U2865 (N_2865,N_2374,N_2419);
xnor U2866 (N_2866,N_2412,N_2432);
and U2867 (N_2867,N_2153,N_2218);
nand U2868 (N_2868,N_2316,N_2453);
xor U2869 (N_2869,N_2466,N_2091);
and U2870 (N_2870,N_2009,N_2139);
xnor U2871 (N_2871,N_2077,N_2053);
and U2872 (N_2872,N_2215,N_2339);
and U2873 (N_2873,N_2112,N_2423);
xnor U2874 (N_2874,N_2101,N_2044);
or U2875 (N_2875,N_2054,N_2376);
and U2876 (N_2876,N_2439,N_2285);
nor U2877 (N_2877,N_2050,N_2483);
and U2878 (N_2878,N_2193,N_2445);
or U2879 (N_2879,N_2466,N_2112);
or U2880 (N_2880,N_2251,N_2193);
nor U2881 (N_2881,N_2180,N_2258);
nor U2882 (N_2882,N_2309,N_2413);
nand U2883 (N_2883,N_2407,N_2312);
and U2884 (N_2884,N_2297,N_2130);
and U2885 (N_2885,N_2228,N_2129);
or U2886 (N_2886,N_2044,N_2432);
or U2887 (N_2887,N_2442,N_2432);
nand U2888 (N_2888,N_2224,N_2437);
nor U2889 (N_2889,N_2137,N_2447);
nand U2890 (N_2890,N_2314,N_2406);
and U2891 (N_2891,N_2494,N_2499);
xor U2892 (N_2892,N_2211,N_2474);
and U2893 (N_2893,N_2065,N_2151);
and U2894 (N_2894,N_2490,N_2394);
nand U2895 (N_2895,N_2310,N_2123);
and U2896 (N_2896,N_2388,N_2143);
nor U2897 (N_2897,N_2069,N_2021);
nor U2898 (N_2898,N_2313,N_2370);
xnor U2899 (N_2899,N_2196,N_2381);
or U2900 (N_2900,N_2301,N_2249);
and U2901 (N_2901,N_2372,N_2181);
xnor U2902 (N_2902,N_2402,N_2337);
nand U2903 (N_2903,N_2203,N_2256);
nor U2904 (N_2904,N_2299,N_2491);
xnor U2905 (N_2905,N_2103,N_2306);
nand U2906 (N_2906,N_2367,N_2382);
xor U2907 (N_2907,N_2187,N_2313);
xor U2908 (N_2908,N_2074,N_2231);
nand U2909 (N_2909,N_2317,N_2255);
or U2910 (N_2910,N_2195,N_2372);
and U2911 (N_2911,N_2294,N_2401);
nand U2912 (N_2912,N_2005,N_2434);
and U2913 (N_2913,N_2299,N_2463);
nor U2914 (N_2914,N_2022,N_2299);
or U2915 (N_2915,N_2397,N_2263);
or U2916 (N_2916,N_2492,N_2119);
xnor U2917 (N_2917,N_2372,N_2421);
xnor U2918 (N_2918,N_2255,N_2208);
and U2919 (N_2919,N_2064,N_2451);
nor U2920 (N_2920,N_2232,N_2477);
or U2921 (N_2921,N_2113,N_2356);
and U2922 (N_2922,N_2141,N_2208);
xnor U2923 (N_2923,N_2105,N_2365);
and U2924 (N_2924,N_2137,N_2145);
xnor U2925 (N_2925,N_2230,N_2334);
and U2926 (N_2926,N_2238,N_2233);
nand U2927 (N_2927,N_2276,N_2189);
nand U2928 (N_2928,N_2433,N_2375);
nand U2929 (N_2929,N_2307,N_2173);
nand U2930 (N_2930,N_2176,N_2317);
nor U2931 (N_2931,N_2462,N_2221);
nor U2932 (N_2932,N_2461,N_2380);
xor U2933 (N_2933,N_2389,N_2191);
and U2934 (N_2934,N_2283,N_2325);
xnor U2935 (N_2935,N_2140,N_2078);
and U2936 (N_2936,N_2081,N_2017);
nand U2937 (N_2937,N_2256,N_2375);
or U2938 (N_2938,N_2110,N_2397);
nand U2939 (N_2939,N_2466,N_2280);
nand U2940 (N_2940,N_2264,N_2178);
nor U2941 (N_2941,N_2073,N_2155);
nor U2942 (N_2942,N_2357,N_2247);
xnor U2943 (N_2943,N_2259,N_2201);
and U2944 (N_2944,N_2153,N_2264);
nor U2945 (N_2945,N_2459,N_2010);
xor U2946 (N_2946,N_2261,N_2264);
or U2947 (N_2947,N_2276,N_2324);
nor U2948 (N_2948,N_2409,N_2364);
nand U2949 (N_2949,N_2138,N_2443);
xor U2950 (N_2950,N_2052,N_2358);
or U2951 (N_2951,N_2101,N_2442);
nor U2952 (N_2952,N_2338,N_2180);
xor U2953 (N_2953,N_2099,N_2462);
or U2954 (N_2954,N_2485,N_2298);
xnor U2955 (N_2955,N_2490,N_2264);
nand U2956 (N_2956,N_2203,N_2141);
nand U2957 (N_2957,N_2024,N_2195);
and U2958 (N_2958,N_2496,N_2442);
xor U2959 (N_2959,N_2332,N_2059);
and U2960 (N_2960,N_2021,N_2110);
nor U2961 (N_2961,N_2206,N_2435);
nor U2962 (N_2962,N_2036,N_2400);
nand U2963 (N_2963,N_2022,N_2467);
nor U2964 (N_2964,N_2457,N_2270);
xor U2965 (N_2965,N_2348,N_2131);
or U2966 (N_2966,N_2075,N_2178);
nor U2967 (N_2967,N_2113,N_2368);
xor U2968 (N_2968,N_2048,N_2157);
nand U2969 (N_2969,N_2004,N_2393);
and U2970 (N_2970,N_2452,N_2374);
nand U2971 (N_2971,N_2109,N_2436);
or U2972 (N_2972,N_2097,N_2060);
xnor U2973 (N_2973,N_2363,N_2487);
or U2974 (N_2974,N_2443,N_2258);
nor U2975 (N_2975,N_2421,N_2091);
nand U2976 (N_2976,N_2316,N_2055);
nor U2977 (N_2977,N_2001,N_2253);
nor U2978 (N_2978,N_2397,N_2211);
xor U2979 (N_2979,N_2434,N_2429);
and U2980 (N_2980,N_2176,N_2306);
nor U2981 (N_2981,N_2301,N_2148);
or U2982 (N_2982,N_2262,N_2293);
or U2983 (N_2983,N_2023,N_2216);
or U2984 (N_2984,N_2182,N_2293);
and U2985 (N_2985,N_2410,N_2051);
xor U2986 (N_2986,N_2216,N_2318);
nor U2987 (N_2987,N_2076,N_2475);
xor U2988 (N_2988,N_2364,N_2340);
xnor U2989 (N_2989,N_2246,N_2266);
nand U2990 (N_2990,N_2308,N_2341);
and U2991 (N_2991,N_2212,N_2198);
xor U2992 (N_2992,N_2354,N_2380);
and U2993 (N_2993,N_2429,N_2385);
xor U2994 (N_2994,N_2413,N_2062);
xnor U2995 (N_2995,N_2317,N_2064);
and U2996 (N_2996,N_2175,N_2290);
and U2997 (N_2997,N_2379,N_2391);
nor U2998 (N_2998,N_2451,N_2299);
or U2999 (N_2999,N_2296,N_2071);
nor U3000 (N_3000,N_2723,N_2551);
and U3001 (N_3001,N_2704,N_2757);
xor U3002 (N_3002,N_2534,N_2839);
and U3003 (N_3003,N_2556,N_2832);
nand U3004 (N_3004,N_2781,N_2697);
nor U3005 (N_3005,N_2884,N_2696);
nand U3006 (N_3006,N_2703,N_2528);
nor U3007 (N_3007,N_2974,N_2867);
nand U3008 (N_3008,N_2898,N_2956);
and U3009 (N_3009,N_2519,N_2661);
and U3010 (N_3010,N_2613,N_2773);
nor U3011 (N_3011,N_2564,N_2973);
xor U3012 (N_3012,N_2560,N_2550);
nand U3013 (N_3013,N_2817,N_2855);
or U3014 (N_3014,N_2951,N_2758);
nor U3015 (N_3015,N_2657,N_2744);
or U3016 (N_3016,N_2761,N_2920);
or U3017 (N_3017,N_2529,N_2507);
or U3018 (N_3018,N_2796,N_2578);
nor U3019 (N_3019,N_2607,N_2577);
or U3020 (N_3020,N_2522,N_2909);
nor U3021 (N_3021,N_2666,N_2615);
xnor U3022 (N_3022,N_2640,N_2732);
or U3023 (N_3023,N_2769,N_2838);
and U3024 (N_3024,N_2901,N_2617);
nand U3025 (N_3025,N_2902,N_2997);
xnor U3026 (N_3026,N_2962,N_2824);
or U3027 (N_3027,N_2558,N_2970);
nor U3028 (N_3028,N_2503,N_2934);
xor U3029 (N_3029,N_2881,N_2953);
nor U3030 (N_3030,N_2853,N_2561);
nor U3031 (N_3031,N_2795,N_2592);
nor U3032 (N_3032,N_2699,N_2762);
or U3033 (N_3033,N_2848,N_2642);
nand U3034 (N_3034,N_2656,N_2980);
or U3035 (N_3035,N_2771,N_2683);
xor U3036 (N_3036,N_2739,N_2584);
nand U3037 (N_3037,N_2768,N_2552);
nor U3038 (N_3038,N_2882,N_2897);
and U3039 (N_3039,N_2525,N_2767);
nand U3040 (N_3040,N_2601,N_2943);
or U3041 (N_3041,N_2931,N_2567);
or U3042 (N_3042,N_2537,N_2936);
and U3043 (N_3043,N_2527,N_2856);
or U3044 (N_3044,N_2994,N_2983);
or U3045 (N_3045,N_2581,N_2937);
xnor U3046 (N_3046,N_2738,N_2665);
and U3047 (N_3047,N_2565,N_2634);
and U3048 (N_3048,N_2646,N_2643);
nand U3049 (N_3049,N_2857,N_2804);
or U3050 (N_3050,N_2500,N_2921);
xor U3051 (N_3051,N_2737,N_2830);
nor U3052 (N_3052,N_2576,N_2506);
nor U3053 (N_3053,N_2833,N_2981);
and U3054 (N_3054,N_2978,N_2850);
nor U3055 (N_3055,N_2915,N_2653);
and U3056 (N_3056,N_2835,N_2521);
and U3057 (N_3057,N_2972,N_2539);
and U3058 (N_3058,N_2698,N_2549);
and U3059 (N_3059,N_2952,N_2783);
nor U3060 (N_3060,N_2545,N_2533);
xnor U3061 (N_3061,N_2518,N_2892);
or U3062 (N_3062,N_2711,N_2676);
and U3063 (N_3063,N_2818,N_2582);
or U3064 (N_3064,N_2861,N_2509);
nand U3065 (N_3065,N_2919,N_2886);
nand U3066 (N_3066,N_2928,N_2787);
xnor U3067 (N_3067,N_2664,N_2627);
nand U3068 (N_3068,N_2825,N_2917);
and U3069 (N_3069,N_2680,N_2786);
and U3070 (N_3070,N_2714,N_2930);
nand U3071 (N_3071,N_2932,N_2942);
or U3072 (N_3072,N_2712,N_2692);
nand U3073 (N_3073,N_2702,N_2979);
nand U3074 (N_3074,N_2910,N_2988);
nand U3075 (N_3075,N_2846,N_2587);
nand U3076 (N_3076,N_2730,N_2555);
and U3077 (N_3077,N_2645,N_2879);
nor U3078 (N_3078,N_2746,N_2517);
or U3079 (N_3079,N_2831,N_2700);
and U3080 (N_3080,N_2829,N_2905);
or U3081 (N_3081,N_2961,N_2514);
and U3082 (N_3082,N_2733,N_2624);
nor U3083 (N_3083,N_2605,N_2793);
nor U3084 (N_3084,N_2826,N_2914);
nor U3085 (N_3085,N_2508,N_2754);
and U3086 (N_3086,N_2990,N_2992);
xor U3087 (N_3087,N_2625,N_2669);
or U3088 (N_3088,N_2513,N_2718);
xnor U3089 (N_3089,N_2899,N_2784);
nand U3090 (N_3090,N_2925,N_2659);
xor U3091 (N_3091,N_2976,N_2885);
and U3092 (N_3092,N_2893,N_2713);
nand U3093 (N_3093,N_2594,N_2929);
and U3094 (N_3094,N_2690,N_2864);
nor U3095 (N_3095,N_2707,N_2996);
nand U3096 (N_3096,N_2782,N_2819);
nand U3097 (N_3097,N_2862,N_2858);
nand U3098 (N_3098,N_2541,N_2721);
nor U3099 (N_3099,N_2619,N_2540);
and U3100 (N_3100,N_2751,N_2610);
nand U3101 (N_3101,N_2759,N_2868);
nand U3102 (N_3102,N_2637,N_2750);
xnor U3103 (N_3103,N_2741,N_2623);
xor U3104 (N_3104,N_2671,N_2851);
xor U3105 (N_3105,N_2877,N_2570);
xnor U3106 (N_3106,N_2844,N_2821);
and U3107 (N_3107,N_2789,N_2938);
nand U3108 (N_3108,N_2719,N_2860);
nand U3109 (N_3109,N_2810,N_2559);
or U3110 (N_3110,N_2813,N_2675);
and U3111 (N_3111,N_2922,N_2583);
nor U3112 (N_3112,N_2725,N_2621);
or U3113 (N_3113,N_2799,N_2672);
nor U3114 (N_3114,N_2775,N_2971);
and U3115 (N_3115,N_2889,N_2542);
and U3116 (N_3116,N_2984,N_2691);
nand U3117 (N_3117,N_2964,N_2635);
and U3118 (N_3118,N_2599,N_2535);
nor U3119 (N_3119,N_2797,N_2989);
or U3120 (N_3120,N_2727,N_2842);
or U3121 (N_3121,N_2650,N_2536);
or U3122 (N_3122,N_2674,N_2742);
xnor U3123 (N_3123,N_2710,N_2649);
and U3124 (N_3124,N_2986,N_2816);
and U3125 (N_3125,N_2532,N_2798);
or U3126 (N_3126,N_2945,N_2572);
and U3127 (N_3127,N_2566,N_2652);
xor U3128 (N_3128,N_2631,N_2597);
and U3129 (N_3129,N_2553,N_2622);
and U3130 (N_3130,N_2809,N_2734);
xnor U3131 (N_3131,N_2852,N_2726);
nor U3132 (N_3132,N_2579,N_2959);
nor U3133 (N_3133,N_2903,N_2632);
or U3134 (N_3134,N_2965,N_2554);
nand U3135 (N_3135,N_2593,N_2891);
and U3136 (N_3136,N_2684,N_2590);
or U3137 (N_3137,N_2695,N_2763);
nor U3138 (N_3138,N_2926,N_2620);
xor U3139 (N_3139,N_2717,N_2505);
and U3140 (N_3140,N_2548,N_2849);
or U3141 (N_3141,N_2686,N_2639);
and U3142 (N_3142,N_2985,N_2569);
or U3143 (N_3143,N_2894,N_2526);
and U3144 (N_3144,N_2870,N_2629);
nand U3145 (N_3145,N_2792,N_2504);
xor U3146 (N_3146,N_2820,N_2907);
nor U3147 (N_3147,N_2764,N_2944);
nand U3148 (N_3148,N_2600,N_2557);
nor U3149 (N_3149,N_2801,N_2573);
or U3150 (N_3150,N_2955,N_2766);
nand U3151 (N_3151,N_2606,N_2644);
nand U3152 (N_3152,N_2512,N_2747);
nor U3153 (N_3153,N_2777,N_2854);
and U3154 (N_3154,N_2982,N_2918);
nor U3155 (N_3155,N_2511,N_2654);
nor U3156 (N_3156,N_2682,N_2840);
xor U3157 (N_3157,N_2681,N_2660);
and U3158 (N_3158,N_2641,N_2628);
or U3159 (N_3159,N_2941,N_2589);
or U3160 (N_3160,N_2515,N_2823);
and U3161 (N_3161,N_2706,N_2872);
and U3162 (N_3162,N_2688,N_2720);
and U3163 (N_3163,N_2633,N_2626);
xor U3164 (N_3164,N_2999,N_2608);
and U3165 (N_3165,N_2603,N_2794);
nor U3166 (N_3166,N_2591,N_2586);
or U3167 (N_3167,N_2708,N_2845);
nand U3168 (N_3168,N_2687,N_2602);
nor U3169 (N_3169,N_2729,N_2563);
nor U3170 (N_3170,N_2568,N_2803);
nor U3171 (N_3171,N_2724,N_2800);
or U3172 (N_3172,N_2812,N_2530);
and U3173 (N_3173,N_2960,N_2774);
or U3174 (N_3174,N_2736,N_2531);
and U3175 (N_3175,N_2836,N_2655);
xor U3176 (N_3176,N_2705,N_2651);
nand U3177 (N_3177,N_2940,N_2895);
xnor U3178 (N_3178,N_2807,N_2874);
nor U3179 (N_3179,N_2806,N_2957);
nand U3180 (N_3180,N_2662,N_2866);
or U3181 (N_3181,N_2544,N_2574);
xor U3182 (N_3182,N_2906,N_2614);
nor U3183 (N_3183,N_2948,N_2547);
or U3184 (N_3184,N_2752,N_2811);
nand U3185 (N_3185,N_2648,N_2735);
or U3186 (N_3186,N_2760,N_2876);
xor U3187 (N_3187,N_2828,N_2896);
xnor U3188 (N_3188,N_2880,N_2949);
or U3189 (N_3189,N_2638,N_2658);
or U3190 (N_3190,N_2679,N_2841);
nand U3191 (N_3191,N_2731,N_2967);
or U3192 (N_3192,N_2950,N_2670);
and U3193 (N_3193,N_2749,N_2709);
or U3194 (N_3194,N_2755,N_2791);
xor U3195 (N_3195,N_2743,N_2993);
nand U3196 (N_3196,N_2543,N_2701);
and U3197 (N_3197,N_2822,N_2745);
nand U3198 (N_3198,N_2588,N_2609);
and U3199 (N_3199,N_2693,N_2788);
nand U3200 (N_3200,N_2770,N_2916);
nor U3201 (N_3201,N_2923,N_2611);
or U3202 (N_3202,N_2875,N_2524);
and U3203 (N_3203,N_2668,N_2685);
nor U3204 (N_3204,N_2636,N_2785);
and U3205 (N_3205,N_2677,N_2694);
or U3206 (N_3206,N_2562,N_2673);
xor U3207 (N_3207,N_2888,N_2900);
and U3208 (N_3208,N_2630,N_2502);
nand U3209 (N_3209,N_2616,N_2538);
and U3210 (N_3210,N_2596,N_2969);
and U3211 (N_3211,N_2748,N_2779);
xor U3212 (N_3212,N_2546,N_2924);
nand U3213 (N_3213,N_2865,N_2501);
and U3214 (N_3214,N_2520,N_2756);
nor U3215 (N_3215,N_2523,N_2808);
or U3216 (N_3216,N_2998,N_2753);
and U3217 (N_3217,N_2991,N_2716);
and U3218 (N_3218,N_2618,N_2933);
nor U3219 (N_3219,N_2966,N_2667);
nor U3220 (N_3220,N_2663,N_2689);
or U3221 (N_3221,N_2847,N_2935);
or U3222 (N_3222,N_2968,N_2975);
xnor U3223 (N_3223,N_2987,N_2927);
and U3224 (N_3224,N_2604,N_2887);
xor U3225 (N_3225,N_2871,N_2571);
or U3226 (N_3226,N_2805,N_2575);
xnor U3227 (N_3227,N_2834,N_2977);
and U3228 (N_3228,N_2647,N_2814);
and U3229 (N_3229,N_2815,N_2963);
or U3230 (N_3230,N_2912,N_2790);
xnor U3231 (N_3231,N_2802,N_2780);
and U3232 (N_3232,N_2772,N_2612);
xnor U3233 (N_3233,N_2837,N_2740);
nand U3234 (N_3234,N_2765,N_2904);
nor U3235 (N_3235,N_2776,N_2946);
nand U3236 (N_3236,N_2843,N_2715);
nor U3237 (N_3237,N_2585,N_2995);
xor U3238 (N_3238,N_2869,N_2516);
xnor U3239 (N_3239,N_2580,N_2722);
nand U3240 (N_3240,N_2908,N_2859);
nor U3241 (N_3241,N_2778,N_2873);
or U3242 (N_3242,N_2883,N_2595);
xnor U3243 (N_3243,N_2678,N_2827);
or U3244 (N_3244,N_2878,N_2954);
or U3245 (N_3245,N_2913,N_2947);
xnor U3246 (N_3246,N_2911,N_2510);
xnor U3247 (N_3247,N_2728,N_2958);
xor U3248 (N_3248,N_2939,N_2890);
nor U3249 (N_3249,N_2863,N_2598);
xor U3250 (N_3250,N_2706,N_2895);
nand U3251 (N_3251,N_2634,N_2754);
nand U3252 (N_3252,N_2966,N_2761);
nand U3253 (N_3253,N_2723,N_2912);
nand U3254 (N_3254,N_2520,N_2805);
nor U3255 (N_3255,N_2642,N_2665);
nand U3256 (N_3256,N_2840,N_2645);
and U3257 (N_3257,N_2874,N_2765);
nor U3258 (N_3258,N_2934,N_2615);
nand U3259 (N_3259,N_2977,N_2979);
xor U3260 (N_3260,N_2924,N_2550);
xor U3261 (N_3261,N_2657,N_2538);
or U3262 (N_3262,N_2914,N_2700);
nand U3263 (N_3263,N_2633,N_2817);
xnor U3264 (N_3264,N_2618,N_2776);
nand U3265 (N_3265,N_2716,N_2592);
and U3266 (N_3266,N_2924,N_2772);
or U3267 (N_3267,N_2821,N_2985);
and U3268 (N_3268,N_2518,N_2820);
or U3269 (N_3269,N_2550,N_2723);
or U3270 (N_3270,N_2667,N_2688);
and U3271 (N_3271,N_2826,N_2908);
nand U3272 (N_3272,N_2661,N_2507);
or U3273 (N_3273,N_2964,N_2757);
and U3274 (N_3274,N_2777,N_2832);
xor U3275 (N_3275,N_2610,N_2872);
xor U3276 (N_3276,N_2627,N_2899);
or U3277 (N_3277,N_2682,N_2593);
nor U3278 (N_3278,N_2686,N_2673);
nor U3279 (N_3279,N_2539,N_2585);
nor U3280 (N_3280,N_2845,N_2762);
or U3281 (N_3281,N_2967,N_2595);
nor U3282 (N_3282,N_2966,N_2794);
and U3283 (N_3283,N_2900,N_2992);
xor U3284 (N_3284,N_2861,N_2645);
xnor U3285 (N_3285,N_2962,N_2590);
nand U3286 (N_3286,N_2847,N_2998);
nand U3287 (N_3287,N_2755,N_2938);
or U3288 (N_3288,N_2722,N_2649);
nor U3289 (N_3289,N_2962,N_2949);
nor U3290 (N_3290,N_2827,N_2956);
xor U3291 (N_3291,N_2672,N_2563);
and U3292 (N_3292,N_2760,N_2735);
or U3293 (N_3293,N_2965,N_2808);
nand U3294 (N_3294,N_2638,N_2896);
nand U3295 (N_3295,N_2828,N_2668);
or U3296 (N_3296,N_2840,N_2671);
and U3297 (N_3297,N_2993,N_2880);
and U3298 (N_3298,N_2973,N_2763);
and U3299 (N_3299,N_2840,N_2750);
xor U3300 (N_3300,N_2817,N_2742);
or U3301 (N_3301,N_2819,N_2663);
or U3302 (N_3302,N_2948,N_2856);
or U3303 (N_3303,N_2532,N_2801);
or U3304 (N_3304,N_2572,N_2990);
xor U3305 (N_3305,N_2761,N_2982);
and U3306 (N_3306,N_2876,N_2657);
nand U3307 (N_3307,N_2838,N_2730);
xor U3308 (N_3308,N_2825,N_2850);
nand U3309 (N_3309,N_2652,N_2663);
nand U3310 (N_3310,N_2746,N_2587);
nand U3311 (N_3311,N_2528,N_2717);
nor U3312 (N_3312,N_2944,N_2607);
and U3313 (N_3313,N_2586,N_2995);
nor U3314 (N_3314,N_2800,N_2656);
or U3315 (N_3315,N_2775,N_2772);
nand U3316 (N_3316,N_2596,N_2920);
nand U3317 (N_3317,N_2882,N_2516);
or U3318 (N_3318,N_2656,N_2974);
xor U3319 (N_3319,N_2976,N_2894);
nor U3320 (N_3320,N_2916,N_2640);
xor U3321 (N_3321,N_2722,N_2600);
nor U3322 (N_3322,N_2689,N_2528);
nand U3323 (N_3323,N_2730,N_2729);
nor U3324 (N_3324,N_2782,N_2783);
xnor U3325 (N_3325,N_2584,N_2773);
nor U3326 (N_3326,N_2878,N_2578);
nand U3327 (N_3327,N_2567,N_2543);
xnor U3328 (N_3328,N_2755,N_2902);
nand U3329 (N_3329,N_2639,N_2895);
nand U3330 (N_3330,N_2573,N_2994);
or U3331 (N_3331,N_2569,N_2766);
xor U3332 (N_3332,N_2591,N_2746);
xor U3333 (N_3333,N_2803,N_2559);
or U3334 (N_3334,N_2742,N_2765);
or U3335 (N_3335,N_2962,N_2928);
xnor U3336 (N_3336,N_2821,N_2834);
nand U3337 (N_3337,N_2776,N_2633);
or U3338 (N_3338,N_2644,N_2871);
nand U3339 (N_3339,N_2569,N_2773);
and U3340 (N_3340,N_2707,N_2580);
nand U3341 (N_3341,N_2688,N_2969);
or U3342 (N_3342,N_2902,N_2912);
and U3343 (N_3343,N_2539,N_2657);
and U3344 (N_3344,N_2556,N_2647);
nor U3345 (N_3345,N_2988,N_2659);
nor U3346 (N_3346,N_2599,N_2744);
nor U3347 (N_3347,N_2587,N_2555);
or U3348 (N_3348,N_2772,N_2586);
and U3349 (N_3349,N_2504,N_2999);
nand U3350 (N_3350,N_2622,N_2884);
xor U3351 (N_3351,N_2893,N_2578);
nand U3352 (N_3352,N_2688,N_2531);
nor U3353 (N_3353,N_2727,N_2725);
nor U3354 (N_3354,N_2989,N_2899);
nor U3355 (N_3355,N_2640,N_2668);
xnor U3356 (N_3356,N_2821,N_2796);
xnor U3357 (N_3357,N_2991,N_2597);
and U3358 (N_3358,N_2940,N_2816);
nand U3359 (N_3359,N_2925,N_2877);
or U3360 (N_3360,N_2878,N_2619);
or U3361 (N_3361,N_2596,N_2981);
xnor U3362 (N_3362,N_2799,N_2900);
or U3363 (N_3363,N_2822,N_2960);
nor U3364 (N_3364,N_2980,N_2855);
xor U3365 (N_3365,N_2778,N_2618);
xnor U3366 (N_3366,N_2913,N_2827);
xnor U3367 (N_3367,N_2626,N_2517);
or U3368 (N_3368,N_2711,N_2990);
nor U3369 (N_3369,N_2982,N_2666);
and U3370 (N_3370,N_2769,N_2682);
xor U3371 (N_3371,N_2686,N_2608);
nor U3372 (N_3372,N_2769,N_2766);
and U3373 (N_3373,N_2840,N_2991);
nor U3374 (N_3374,N_2517,N_2624);
nand U3375 (N_3375,N_2590,N_2571);
and U3376 (N_3376,N_2915,N_2998);
or U3377 (N_3377,N_2803,N_2887);
xor U3378 (N_3378,N_2773,N_2868);
xor U3379 (N_3379,N_2634,N_2840);
nand U3380 (N_3380,N_2972,N_2562);
and U3381 (N_3381,N_2629,N_2929);
or U3382 (N_3382,N_2752,N_2545);
xor U3383 (N_3383,N_2874,N_2841);
nand U3384 (N_3384,N_2554,N_2611);
and U3385 (N_3385,N_2860,N_2811);
or U3386 (N_3386,N_2912,N_2956);
nor U3387 (N_3387,N_2867,N_2727);
xnor U3388 (N_3388,N_2970,N_2667);
nand U3389 (N_3389,N_2766,N_2847);
nor U3390 (N_3390,N_2597,N_2959);
or U3391 (N_3391,N_2729,N_2503);
or U3392 (N_3392,N_2977,N_2535);
nand U3393 (N_3393,N_2570,N_2913);
or U3394 (N_3394,N_2924,N_2654);
and U3395 (N_3395,N_2827,N_2914);
and U3396 (N_3396,N_2859,N_2833);
xor U3397 (N_3397,N_2834,N_2940);
xor U3398 (N_3398,N_2756,N_2933);
and U3399 (N_3399,N_2623,N_2996);
and U3400 (N_3400,N_2668,N_2991);
and U3401 (N_3401,N_2510,N_2881);
nand U3402 (N_3402,N_2779,N_2688);
or U3403 (N_3403,N_2535,N_2678);
and U3404 (N_3404,N_2830,N_2996);
nor U3405 (N_3405,N_2503,N_2703);
xnor U3406 (N_3406,N_2868,N_2782);
nand U3407 (N_3407,N_2741,N_2571);
and U3408 (N_3408,N_2811,N_2639);
nand U3409 (N_3409,N_2670,N_2925);
or U3410 (N_3410,N_2830,N_2901);
and U3411 (N_3411,N_2768,N_2585);
nand U3412 (N_3412,N_2705,N_2795);
xor U3413 (N_3413,N_2679,N_2635);
and U3414 (N_3414,N_2944,N_2538);
nor U3415 (N_3415,N_2980,N_2580);
xor U3416 (N_3416,N_2776,N_2690);
xnor U3417 (N_3417,N_2950,N_2875);
xor U3418 (N_3418,N_2969,N_2754);
or U3419 (N_3419,N_2660,N_2795);
or U3420 (N_3420,N_2795,N_2632);
and U3421 (N_3421,N_2934,N_2576);
nand U3422 (N_3422,N_2508,N_2538);
or U3423 (N_3423,N_2665,N_2744);
nor U3424 (N_3424,N_2831,N_2838);
and U3425 (N_3425,N_2806,N_2903);
and U3426 (N_3426,N_2756,N_2757);
xor U3427 (N_3427,N_2830,N_2878);
and U3428 (N_3428,N_2811,N_2588);
or U3429 (N_3429,N_2936,N_2686);
nand U3430 (N_3430,N_2516,N_2583);
and U3431 (N_3431,N_2759,N_2912);
xnor U3432 (N_3432,N_2910,N_2664);
xor U3433 (N_3433,N_2885,N_2861);
xnor U3434 (N_3434,N_2816,N_2616);
xor U3435 (N_3435,N_2843,N_2674);
and U3436 (N_3436,N_2641,N_2759);
xnor U3437 (N_3437,N_2741,N_2539);
xnor U3438 (N_3438,N_2569,N_2977);
xor U3439 (N_3439,N_2620,N_2792);
or U3440 (N_3440,N_2735,N_2738);
xnor U3441 (N_3441,N_2529,N_2617);
xor U3442 (N_3442,N_2862,N_2504);
nor U3443 (N_3443,N_2818,N_2561);
or U3444 (N_3444,N_2764,N_2644);
nand U3445 (N_3445,N_2553,N_2818);
or U3446 (N_3446,N_2863,N_2647);
and U3447 (N_3447,N_2919,N_2699);
or U3448 (N_3448,N_2633,N_2923);
nand U3449 (N_3449,N_2527,N_2682);
xor U3450 (N_3450,N_2573,N_2625);
nand U3451 (N_3451,N_2975,N_2587);
xnor U3452 (N_3452,N_2578,N_2937);
and U3453 (N_3453,N_2527,N_2992);
nor U3454 (N_3454,N_2602,N_2638);
xor U3455 (N_3455,N_2962,N_2520);
or U3456 (N_3456,N_2513,N_2979);
or U3457 (N_3457,N_2692,N_2640);
xnor U3458 (N_3458,N_2965,N_2916);
and U3459 (N_3459,N_2698,N_2516);
or U3460 (N_3460,N_2869,N_2703);
nand U3461 (N_3461,N_2503,N_2635);
and U3462 (N_3462,N_2887,N_2569);
xor U3463 (N_3463,N_2708,N_2846);
or U3464 (N_3464,N_2661,N_2775);
xor U3465 (N_3465,N_2833,N_2806);
or U3466 (N_3466,N_2866,N_2896);
nor U3467 (N_3467,N_2987,N_2843);
nor U3468 (N_3468,N_2829,N_2933);
nand U3469 (N_3469,N_2739,N_2769);
nand U3470 (N_3470,N_2747,N_2503);
and U3471 (N_3471,N_2875,N_2901);
xnor U3472 (N_3472,N_2756,N_2892);
nand U3473 (N_3473,N_2533,N_2568);
and U3474 (N_3474,N_2699,N_2796);
xor U3475 (N_3475,N_2870,N_2552);
and U3476 (N_3476,N_2546,N_2739);
nand U3477 (N_3477,N_2702,N_2690);
or U3478 (N_3478,N_2818,N_2573);
nand U3479 (N_3479,N_2989,N_2831);
nand U3480 (N_3480,N_2618,N_2703);
nand U3481 (N_3481,N_2684,N_2969);
nor U3482 (N_3482,N_2705,N_2803);
or U3483 (N_3483,N_2681,N_2688);
or U3484 (N_3484,N_2589,N_2658);
xnor U3485 (N_3485,N_2909,N_2980);
nor U3486 (N_3486,N_2552,N_2756);
nand U3487 (N_3487,N_2687,N_2917);
nand U3488 (N_3488,N_2618,N_2870);
nor U3489 (N_3489,N_2786,N_2673);
xor U3490 (N_3490,N_2922,N_2699);
and U3491 (N_3491,N_2587,N_2682);
and U3492 (N_3492,N_2800,N_2695);
xnor U3493 (N_3493,N_2561,N_2944);
and U3494 (N_3494,N_2877,N_2707);
nor U3495 (N_3495,N_2620,N_2671);
nor U3496 (N_3496,N_2531,N_2775);
or U3497 (N_3497,N_2808,N_2810);
nor U3498 (N_3498,N_2614,N_2815);
nor U3499 (N_3499,N_2589,N_2695);
nand U3500 (N_3500,N_3223,N_3110);
nor U3501 (N_3501,N_3403,N_3211);
or U3502 (N_3502,N_3380,N_3362);
nand U3503 (N_3503,N_3332,N_3202);
and U3504 (N_3504,N_3348,N_3026);
nor U3505 (N_3505,N_3129,N_3323);
xor U3506 (N_3506,N_3014,N_3391);
nor U3507 (N_3507,N_3250,N_3133);
or U3508 (N_3508,N_3056,N_3327);
nand U3509 (N_3509,N_3141,N_3020);
xnor U3510 (N_3510,N_3143,N_3363);
nor U3511 (N_3511,N_3285,N_3090);
nor U3512 (N_3512,N_3075,N_3262);
or U3513 (N_3513,N_3464,N_3140);
or U3514 (N_3514,N_3063,N_3466);
nor U3515 (N_3515,N_3207,N_3259);
or U3516 (N_3516,N_3209,N_3032);
and U3517 (N_3517,N_3389,N_3443);
nor U3518 (N_3518,N_3196,N_3089);
and U3519 (N_3519,N_3491,N_3031);
nand U3520 (N_3520,N_3379,N_3038);
xor U3521 (N_3521,N_3481,N_3122);
and U3522 (N_3522,N_3385,N_3359);
xor U3523 (N_3523,N_3153,N_3247);
or U3524 (N_3524,N_3213,N_3434);
xor U3525 (N_3525,N_3203,N_3084);
or U3526 (N_3526,N_3286,N_3409);
nor U3527 (N_3527,N_3103,N_3139);
or U3528 (N_3528,N_3127,N_3119);
and U3529 (N_3529,N_3179,N_3463);
nor U3530 (N_3530,N_3057,N_3473);
or U3531 (N_3531,N_3137,N_3155);
or U3532 (N_3532,N_3373,N_3046);
nor U3533 (N_3533,N_3219,N_3293);
xnor U3534 (N_3534,N_3030,N_3036);
and U3535 (N_3535,N_3436,N_3192);
nand U3536 (N_3536,N_3483,N_3218);
and U3537 (N_3537,N_3324,N_3414);
and U3538 (N_3538,N_3017,N_3073);
or U3539 (N_3539,N_3095,N_3190);
or U3540 (N_3540,N_3315,N_3292);
and U3541 (N_3541,N_3330,N_3043);
or U3542 (N_3542,N_3333,N_3069);
nor U3543 (N_3543,N_3494,N_3042);
xnor U3544 (N_3544,N_3281,N_3401);
nor U3545 (N_3545,N_3307,N_3412);
nor U3546 (N_3546,N_3449,N_3168);
or U3547 (N_3547,N_3024,N_3260);
nand U3548 (N_3548,N_3461,N_3265);
xnor U3549 (N_3549,N_3462,N_3297);
and U3550 (N_3550,N_3430,N_3130);
or U3551 (N_3551,N_3460,N_3270);
nand U3552 (N_3552,N_3425,N_3134);
nand U3553 (N_3553,N_3033,N_3397);
and U3554 (N_3554,N_3342,N_3275);
or U3555 (N_3555,N_3079,N_3239);
nor U3556 (N_3556,N_3006,N_3337);
nor U3557 (N_3557,N_3244,N_3195);
and U3558 (N_3558,N_3357,N_3156);
and U3559 (N_3559,N_3199,N_3317);
nor U3560 (N_3560,N_3086,N_3162);
nor U3561 (N_3561,N_3366,N_3147);
nand U3562 (N_3562,N_3041,N_3471);
nand U3563 (N_3563,N_3167,N_3375);
xor U3564 (N_3564,N_3496,N_3051);
or U3565 (N_3565,N_3170,N_3116);
nand U3566 (N_3566,N_3040,N_3085);
nor U3567 (N_3567,N_3083,N_3109);
or U3568 (N_3568,N_3393,N_3263);
or U3569 (N_3569,N_3191,N_3115);
or U3570 (N_3570,N_3186,N_3325);
xnor U3571 (N_3571,N_3480,N_3048);
or U3572 (N_3572,N_3182,N_3187);
and U3573 (N_3573,N_3248,N_3231);
or U3574 (N_3574,N_3125,N_3001);
xnor U3575 (N_3575,N_3427,N_3246);
nor U3576 (N_3576,N_3088,N_3451);
or U3577 (N_3577,N_3268,N_3445);
and U3578 (N_3578,N_3124,N_3349);
or U3579 (N_3579,N_3055,N_3234);
xor U3580 (N_3580,N_3012,N_3309);
and U3581 (N_3581,N_3453,N_3291);
and U3582 (N_3582,N_3264,N_3082);
and U3583 (N_3583,N_3267,N_3052);
nand U3584 (N_3584,N_3230,N_3321);
and U3585 (N_3585,N_3238,N_3037);
or U3586 (N_3586,N_3489,N_3128);
xnor U3587 (N_3587,N_3080,N_3365);
and U3588 (N_3588,N_3099,N_3402);
xor U3589 (N_3589,N_3126,N_3013);
and U3590 (N_3590,N_3256,N_3101);
and U3591 (N_3591,N_3484,N_3336);
nand U3592 (N_3592,N_3433,N_3008);
or U3593 (N_3593,N_3132,N_3205);
nor U3594 (N_3594,N_3004,N_3372);
nand U3595 (N_3595,N_3479,N_3396);
or U3596 (N_3596,N_3346,N_3157);
or U3597 (N_3597,N_3197,N_3428);
xnor U3598 (N_3598,N_3354,N_3470);
nor U3599 (N_3599,N_3440,N_3242);
nor U3600 (N_3600,N_3023,N_3229);
nor U3601 (N_3601,N_3065,N_3228);
and U3602 (N_3602,N_3296,N_3169);
and U3603 (N_3603,N_3455,N_3314);
nor U3604 (N_3604,N_3148,N_3039);
xnor U3605 (N_3605,N_3497,N_3111);
xnor U3606 (N_3606,N_3355,N_3255);
xor U3607 (N_3607,N_3283,N_3395);
nor U3608 (N_3608,N_3097,N_3025);
or U3609 (N_3609,N_3261,N_3413);
and U3610 (N_3610,N_3236,N_3439);
nor U3611 (N_3611,N_3353,N_3294);
nand U3612 (N_3612,N_3108,N_3174);
nand U3613 (N_3613,N_3245,N_3383);
or U3614 (N_3614,N_3009,N_3171);
xor U3615 (N_3615,N_3347,N_3107);
nor U3616 (N_3616,N_3341,N_3163);
nor U3617 (N_3617,N_3426,N_3416);
or U3618 (N_3618,N_3210,N_3368);
xnor U3619 (N_3619,N_3176,N_3388);
and U3620 (N_3620,N_3432,N_3422);
xnor U3621 (N_3621,N_3217,N_3257);
or U3622 (N_3622,N_3194,N_3007);
xnor U3623 (N_3623,N_3300,N_3420);
nand U3624 (N_3624,N_3326,N_3472);
xnor U3625 (N_3625,N_3118,N_3058);
xor U3626 (N_3626,N_3266,N_3322);
nor U3627 (N_3627,N_3310,N_3121);
xnor U3628 (N_3628,N_3417,N_3456);
nand U3629 (N_3629,N_3382,N_3328);
xnor U3630 (N_3630,N_3145,N_3295);
or U3631 (N_3631,N_3222,N_3361);
and U3632 (N_3632,N_3374,N_3100);
xnor U3633 (N_3633,N_3165,N_3044);
nor U3634 (N_3634,N_3467,N_3214);
nor U3635 (N_3635,N_3181,N_3068);
and U3636 (N_3636,N_3301,N_3423);
nand U3637 (N_3637,N_3406,N_3486);
and U3638 (N_3638,N_3215,N_3492);
xnor U3639 (N_3639,N_3334,N_3356);
xnor U3640 (N_3640,N_3476,N_3411);
xnor U3641 (N_3641,N_3078,N_3482);
and U3642 (N_3642,N_3367,N_3410);
nor U3643 (N_3643,N_3352,N_3166);
nand U3644 (N_3644,N_3477,N_3272);
nand U3645 (N_3645,N_3340,N_3490);
nor U3646 (N_3646,N_3384,N_3343);
nand U3647 (N_3647,N_3290,N_3399);
or U3648 (N_3648,N_3198,N_3235);
or U3649 (N_3649,N_3249,N_3319);
nand U3650 (N_3650,N_3378,N_3287);
or U3651 (N_3651,N_3370,N_3308);
nand U3652 (N_3652,N_3271,N_3320);
nor U3653 (N_3653,N_3339,N_3240);
and U3654 (N_3654,N_3011,N_3232);
and U3655 (N_3655,N_3488,N_3298);
nand U3656 (N_3656,N_3104,N_3233);
and U3657 (N_3657,N_3050,N_3159);
nor U3658 (N_3658,N_3364,N_3446);
or U3659 (N_3659,N_3421,N_3193);
xor U3660 (N_3660,N_3474,N_3302);
and U3661 (N_3661,N_3431,N_3350);
and U3662 (N_3662,N_3183,N_3276);
xnor U3663 (N_3663,N_3499,N_3028);
nand U3664 (N_3664,N_3498,N_3206);
and U3665 (N_3665,N_3201,N_3180);
nor U3666 (N_3666,N_3220,N_3208);
nand U3667 (N_3667,N_3062,N_3468);
nand U3668 (N_3668,N_3335,N_3096);
nand U3669 (N_3669,N_3120,N_3419);
or U3670 (N_3670,N_3072,N_3151);
nand U3671 (N_3671,N_3149,N_3237);
or U3672 (N_3672,N_3029,N_3304);
nand U3673 (N_3673,N_3243,N_3172);
and U3674 (N_3674,N_3067,N_3369);
or U3675 (N_3675,N_3173,N_3034);
xor U3676 (N_3676,N_3273,N_3282);
and U3677 (N_3677,N_3142,N_3113);
xnor U3678 (N_3678,N_3386,N_3066);
or U3679 (N_3679,N_3061,N_3278);
nand U3680 (N_3680,N_3253,N_3081);
and U3681 (N_3681,N_3241,N_3442);
and U3682 (N_3682,N_3465,N_3459);
nor U3683 (N_3683,N_3478,N_3138);
or U3684 (N_3684,N_3093,N_3010);
or U3685 (N_3685,N_3212,N_3064);
or U3686 (N_3686,N_3105,N_3164);
nand U3687 (N_3687,N_3131,N_3224);
nor U3688 (N_3688,N_3189,N_3071);
xnor U3689 (N_3689,N_3457,N_3152);
xor U3690 (N_3690,N_3398,N_3289);
xnor U3691 (N_3691,N_3252,N_3448);
nor U3692 (N_3692,N_3303,N_3495);
and U3693 (N_3693,N_3318,N_3200);
and U3694 (N_3694,N_3188,N_3150);
or U3695 (N_3695,N_3022,N_3312);
nor U3696 (N_3696,N_3178,N_3184);
nor U3697 (N_3697,N_3076,N_3000);
and U3698 (N_3698,N_3279,N_3280);
nor U3699 (N_3699,N_3005,N_3429);
xor U3700 (N_3700,N_3204,N_3377);
xnor U3701 (N_3701,N_3437,N_3060);
xnor U3702 (N_3702,N_3329,N_3405);
nor U3703 (N_3703,N_3400,N_3035);
nor U3704 (N_3704,N_3216,N_3112);
and U3705 (N_3705,N_3015,N_3049);
or U3706 (N_3706,N_3175,N_3098);
and U3707 (N_3707,N_3311,N_3021);
xor U3708 (N_3708,N_3424,N_3258);
or U3709 (N_3709,N_3381,N_3185);
nand U3710 (N_3710,N_3227,N_3441);
or U3711 (N_3711,N_3158,N_3226);
xnor U3712 (N_3712,N_3387,N_3114);
nor U3713 (N_3713,N_3135,N_3077);
xor U3714 (N_3714,N_3418,N_3092);
or U3715 (N_3715,N_3160,N_3102);
nor U3716 (N_3716,N_3123,N_3117);
xnor U3717 (N_3717,N_3177,N_3018);
nor U3718 (N_3718,N_3094,N_3254);
or U3719 (N_3719,N_3438,N_3392);
nand U3720 (N_3720,N_3091,N_3371);
nor U3721 (N_3721,N_3045,N_3106);
nor U3722 (N_3722,N_3444,N_3306);
nand U3723 (N_3723,N_3344,N_3475);
and U3724 (N_3724,N_3493,N_3313);
nand U3725 (N_3725,N_3435,N_3274);
xnor U3726 (N_3726,N_3415,N_3450);
xnor U3727 (N_3727,N_3408,N_3154);
xnor U3728 (N_3728,N_3338,N_3027);
nor U3729 (N_3729,N_3316,N_3345);
xor U3730 (N_3730,N_3331,N_3146);
and U3731 (N_3731,N_3144,N_3070);
nand U3732 (N_3732,N_3221,N_3269);
and U3733 (N_3733,N_3452,N_3019);
and U3734 (N_3734,N_3251,N_3161);
xnor U3735 (N_3735,N_3284,N_3469);
nor U3736 (N_3736,N_3407,N_3059);
or U3737 (N_3737,N_3458,N_3376);
xor U3738 (N_3738,N_3351,N_3136);
or U3739 (N_3739,N_3074,N_3054);
xnor U3740 (N_3740,N_3277,N_3390);
xor U3741 (N_3741,N_3447,N_3087);
nor U3742 (N_3742,N_3358,N_3404);
nand U3743 (N_3743,N_3002,N_3299);
xor U3744 (N_3744,N_3305,N_3487);
and U3745 (N_3745,N_3003,N_3288);
or U3746 (N_3746,N_3016,N_3394);
xnor U3747 (N_3747,N_3454,N_3053);
nand U3748 (N_3748,N_3225,N_3360);
or U3749 (N_3749,N_3485,N_3047);
nand U3750 (N_3750,N_3149,N_3360);
or U3751 (N_3751,N_3271,N_3340);
xnor U3752 (N_3752,N_3130,N_3056);
nand U3753 (N_3753,N_3077,N_3219);
nor U3754 (N_3754,N_3480,N_3412);
or U3755 (N_3755,N_3082,N_3086);
or U3756 (N_3756,N_3420,N_3044);
xnor U3757 (N_3757,N_3129,N_3211);
and U3758 (N_3758,N_3338,N_3070);
nor U3759 (N_3759,N_3387,N_3218);
nor U3760 (N_3760,N_3349,N_3188);
nand U3761 (N_3761,N_3494,N_3116);
nor U3762 (N_3762,N_3292,N_3009);
nand U3763 (N_3763,N_3471,N_3466);
xnor U3764 (N_3764,N_3423,N_3420);
xor U3765 (N_3765,N_3203,N_3298);
nand U3766 (N_3766,N_3308,N_3040);
or U3767 (N_3767,N_3369,N_3263);
xnor U3768 (N_3768,N_3214,N_3279);
nor U3769 (N_3769,N_3290,N_3163);
or U3770 (N_3770,N_3150,N_3233);
or U3771 (N_3771,N_3373,N_3268);
and U3772 (N_3772,N_3100,N_3431);
or U3773 (N_3773,N_3408,N_3265);
and U3774 (N_3774,N_3324,N_3341);
and U3775 (N_3775,N_3260,N_3317);
nand U3776 (N_3776,N_3475,N_3261);
nand U3777 (N_3777,N_3370,N_3477);
or U3778 (N_3778,N_3433,N_3080);
nor U3779 (N_3779,N_3309,N_3341);
or U3780 (N_3780,N_3219,N_3012);
nor U3781 (N_3781,N_3377,N_3347);
and U3782 (N_3782,N_3376,N_3021);
and U3783 (N_3783,N_3001,N_3430);
xor U3784 (N_3784,N_3225,N_3371);
and U3785 (N_3785,N_3069,N_3302);
and U3786 (N_3786,N_3209,N_3291);
or U3787 (N_3787,N_3288,N_3070);
and U3788 (N_3788,N_3026,N_3174);
and U3789 (N_3789,N_3314,N_3296);
xnor U3790 (N_3790,N_3407,N_3377);
nor U3791 (N_3791,N_3053,N_3254);
xor U3792 (N_3792,N_3186,N_3212);
nor U3793 (N_3793,N_3124,N_3239);
nor U3794 (N_3794,N_3421,N_3004);
nor U3795 (N_3795,N_3021,N_3477);
and U3796 (N_3796,N_3023,N_3458);
nand U3797 (N_3797,N_3098,N_3328);
or U3798 (N_3798,N_3371,N_3323);
and U3799 (N_3799,N_3012,N_3083);
and U3800 (N_3800,N_3483,N_3374);
or U3801 (N_3801,N_3458,N_3208);
nand U3802 (N_3802,N_3338,N_3186);
or U3803 (N_3803,N_3198,N_3096);
xnor U3804 (N_3804,N_3254,N_3179);
nor U3805 (N_3805,N_3098,N_3289);
or U3806 (N_3806,N_3414,N_3294);
xnor U3807 (N_3807,N_3205,N_3101);
nor U3808 (N_3808,N_3468,N_3311);
and U3809 (N_3809,N_3415,N_3042);
xnor U3810 (N_3810,N_3127,N_3095);
or U3811 (N_3811,N_3480,N_3124);
nor U3812 (N_3812,N_3307,N_3322);
or U3813 (N_3813,N_3331,N_3190);
nand U3814 (N_3814,N_3133,N_3375);
and U3815 (N_3815,N_3266,N_3260);
and U3816 (N_3816,N_3439,N_3469);
and U3817 (N_3817,N_3247,N_3180);
or U3818 (N_3818,N_3225,N_3108);
nor U3819 (N_3819,N_3297,N_3185);
and U3820 (N_3820,N_3205,N_3366);
xnor U3821 (N_3821,N_3392,N_3354);
xnor U3822 (N_3822,N_3041,N_3375);
nand U3823 (N_3823,N_3191,N_3425);
or U3824 (N_3824,N_3111,N_3179);
or U3825 (N_3825,N_3106,N_3089);
xor U3826 (N_3826,N_3312,N_3105);
xor U3827 (N_3827,N_3135,N_3382);
nor U3828 (N_3828,N_3415,N_3156);
nor U3829 (N_3829,N_3069,N_3349);
xor U3830 (N_3830,N_3220,N_3326);
xnor U3831 (N_3831,N_3460,N_3394);
nand U3832 (N_3832,N_3413,N_3410);
and U3833 (N_3833,N_3427,N_3251);
and U3834 (N_3834,N_3399,N_3023);
nor U3835 (N_3835,N_3194,N_3256);
nor U3836 (N_3836,N_3198,N_3119);
or U3837 (N_3837,N_3092,N_3001);
or U3838 (N_3838,N_3056,N_3486);
or U3839 (N_3839,N_3156,N_3378);
or U3840 (N_3840,N_3389,N_3069);
nor U3841 (N_3841,N_3253,N_3298);
and U3842 (N_3842,N_3134,N_3329);
nor U3843 (N_3843,N_3480,N_3204);
xnor U3844 (N_3844,N_3306,N_3063);
xor U3845 (N_3845,N_3395,N_3080);
xor U3846 (N_3846,N_3330,N_3211);
nor U3847 (N_3847,N_3231,N_3052);
or U3848 (N_3848,N_3223,N_3038);
or U3849 (N_3849,N_3000,N_3399);
and U3850 (N_3850,N_3078,N_3040);
nand U3851 (N_3851,N_3331,N_3127);
nor U3852 (N_3852,N_3295,N_3174);
or U3853 (N_3853,N_3402,N_3138);
nor U3854 (N_3854,N_3172,N_3038);
nor U3855 (N_3855,N_3009,N_3236);
nand U3856 (N_3856,N_3049,N_3254);
nor U3857 (N_3857,N_3146,N_3317);
and U3858 (N_3858,N_3179,N_3326);
nand U3859 (N_3859,N_3184,N_3248);
or U3860 (N_3860,N_3368,N_3367);
nor U3861 (N_3861,N_3276,N_3262);
nor U3862 (N_3862,N_3471,N_3207);
and U3863 (N_3863,N_3491,N_3403);
xor U3864 (N_3864,N_3276,N_3255);
or U3865 (N_3865,N_3156,N_3435);
nor U3866 (N_3866,N_3327,N_3291);
nor U3867 (N_3867,N_3146,N_3203);
nor U3868 (N_3868,N_3476,N_3444);
nand U3869 (N_3869,N_3020,N_3362);
and U3870 (N_3870,N_3273,N_3428);
xnor U3871 (N_3871,N_3293,N_3350);
or U3872 (N_3872,N_3046,N_3008);
nor U3873 (N_3873,N_3420,N_3437);
or U3874 (N_3874,N_3205,N_3480);
and U3875 (N_3875,N_3232,N_3472);
or U3876 (N_3876,N_3462,N_3361);
or U3877 (N_3877,N_3484,N_3122);
xnor U3878 (N_3878,N_3276,N_3179);
or U3879 (N_3879,N_3421,N_3207);
xor U3880 (N_3880,N_3412,N_3163);
xor U3881 (N_3881,N_3092,N_3450);
nor U3882 (N_3882,N_3396,N_3433);
xor U3883 (N_3883,N_3220,N_3144);
nor U3884 (N_3884,N_3364,N_3013);
nor U3885 (N_3885,N_3077,N_3067);
and U3886 (N_3886,N_3029,N_3161);
nand U3887 (N_3887,N_3026,N_3415);
nor U3888 (N_3888,N_3494,N_3072);
or U3889 (N_3889,N_3003,N_3100);
or U3890 (N_3890,N_3025,N_3360);
nand U3891 (N_3891,N_3353,N_3330);
nor U3892 (N_3892,N_3358,N_3060);
nand U3893 (N_3893,N_3151,N_3424);
and U3894 (N_3894,N_3411,N_3048);
nor U3895 (N_3895,N_3423,N_3286);
nand U3896 (N_3896,N_3334,N_3142);
xor U3897 (N_3897,N_3225,N_3207);
xor U3898 (N_3898,N_3239,N_3378);
or U3899 (N_3899,N_3442,N_3087);
and U3900 (N_3900,N_3388,N_3480);
nand U3901 (N_3901,N_3443,N_3396);
and U3902 (N_3902,N_3191,N_3335);
nor U3903 (N_3903,N_3293,N_3168);
xor U3904 (N_3904,N_3097,N_3046);
nor U3905 (N_3905,N_3397,N_3011);
and U3906 (N_3906,N_3275,N_3401);
or U3907 (N_3907,N_3226,N_3377);
or U3908 (N_3908,N_3368,N_3204);
nor U3909 (N_3909,N_3290,N_3058);
and U3910 (N_3910,N_3146,N_3496);
xor U3911 (N_3911,N_3263,N_3380);
or U3912 (N_3912,N_3000,N_3281);
nand U3913 (N_3913,N_3310,N_3466);
and U3914 (N_3914,N_3206,N_3395);
nor U3915 (N_3915,N_3159,N_3446);
or U3916 (N_3916,N_3265,N_3455);
xor U3917 (N_3917,N_3332,N_3134);
nor U3918 (N_3918,N_3436,N_3307);
nand U3919 (N_3919,N_3188,N_3412);
and U3920 (N_3920,N_3052,N_3172);
xor U3921 (N_3921,N_3406,N_3169);
nand U3922 (N_3922,N_3062,N_3035);
nor U3923 (N_3923,N_3363,N_3379);
nor U3924 (N_3924,N_3149,N_3476);
nor U3925 (N_3925,N_3155,N_3346);
nor U3926 (N_3926,N_3116,N_3277);
or U3927 (N_3927,N_3448,N_3136);
xnor U3928 (N_3928,N_3456,N_3074);
nand U3929 (N_3929,N_3177,N_3351);
nor U3930 (N_3930,N_3066,N_3188);
or U3931 (N_3931,N_3205,N_3214);
nand U3932 (N_3932,N_3034,N_3386);
or U3933 (N_3933,N_3117,N_3208);
and U3934 (N_3934,N_3047,N_3386);
nor U3935 (N_3935,N_3352,N_3243);
and U3936 (N_3936,N_3081,N_3463);
xor U3937 (N_3937,N_3214,N_3272);
or U3938 (N_3938,N_3420,N_3485);
nor U3939 (N_3939,N_3359,N_3025);
xnor U3940 (N_3940,N_3279,N_3067);
and U3941 (N_3941,N_3382,N_3039);
xor U3942 (N_3942,N_3114,N_3046);
or U3943 (N_3943,N_3463,N_3056);
and U3944 (N_3944,N_3367,N_3454);
and U3945 (N_3945,N_3222,N_3429);
nand U3946 (N_3946,N_3469,N_3093);
nor U3947 (N_3947,N_3226,N_3095);
and U3948 (N_3948,N_3220,N_3327);
nor U3949 (N_3949,N_3015,N_3444);
or U3950 (N_3950,N_3300,N_3495);
xor U3951 (N_3951,N_3045,N_3120);
or U3952 (N_3952,N_3268,N_3086);
nor U3953 (N_3953,N_3162,N_3289);
nand U3954 (N_3954,N_3498,N_3406);
nor U3955 (N_3955,N_3209,N_3415);
or U3956 (N_3956,N_3238,N_3464);
and U3957 (N_3957,N_3334,N_3352);
and U3958 (N_3958,N_3325,N_3141);
or U3959 (N_3959,N_3306,N_3115);
xor U3960 (N_3960,N_3136,N_3271);
nand U3961 (N_3961,N_3237,N_3075);
nand U3962 (N_3962,N_3035,N_3299);
nor U3963 (N_3963,N_3256,N_3403);
nor U3964 (N_3964,N_3378,N_3003);
or U3965 (N_3965,N_3005,N_3249);
or U3966 (N_3966,N_3142,N_3357);
nor U3967 (N_3967,N_3469,N_3379);
nor U3968 (N_3968,N_3258,N_3010);
or U3969 (N_3969,N_3134,N_3178);
nand U3970 (N_3970,N_3451,N_3236);
and U3971 (N_3971,N_3287,N_3208);
nor U3972 (N_3972,N_3487,N_3457);
nand U3973 (N_3973,N_3216,N_3102);
xnor U3974 (N_3974,N_3273,N_3043);
and U3975 (N_3975,N_3490,N_3262);
and U3976 (N_3976,N_3431,N_3189);
xnor U3977 (N_3977,N_3172,N_3005);
xnor U3978 (N_3978,N_3356,N_3243);
and U3979 (N_3979,N_3305,N_3286);
and U3980 (N_3980,N_3274,N_3163);
and U3981 (N_3981,N_3232,N_3411);
and U3982 (N_3982,N_3089,N_3117);
and U3983 (N_3983,N_3057,N_3242);
nand U3984 (N_3984,N_3077,N_3447);
nor U3985 (N_3985,N_3139,N_3288);
xor U3986 (N_3986,N_3353,N_3150);
nand U3987 (N_3987,N_3063,N_3061);
or U3988 (N_3988,N_3209,N_3223);
and U3989 (N_3989,N_3423,N_3022);
nor U3990 (N_3990,N_3460,N_3483);
or U3991 (N_3991,N_3402,N_3280);
or U3992 (N_3992,N_3406,N_3467);
and U3993 (N_3993,N_3174,N_3366);
or U3994 (N_3994,N_3363,N_3055);
and U3995 (N_3995,N_3120,N_3124);
and U3996 (N_3996,N_3388,N_3103);
or U3997 (N_3997,N_3185,N_3452);
or U3998 (N_3998,N_3232,N_3488);
and U3999 (N_3999,N_3269,N_3188);
nand U4000 (N_4000,N_3776,N_3886);
nand U4001 (N_4001,N_3676,N_3868);
nor U4002 (N_4002,N_3936,N_3576);
nand U4003 (N_4003,N_3779,N_3536);
nand U4004 (N_4004,N_3512,N_3574);
xnor U4005 (N_4005,N_3685,N_3882);
and U4006 (N_4006,N_3708,N_3567);
or U4007 (N_4007,N_3553,N_3570);
nand U4008 (N_4008,N_3797,N_3781);
or U4009 (N_4009,N_3627,N_3907);
nor U4010 (N_4010,N_3753,N_3757);
nand U4011 (N_4011,N_3758,N_3878);
and U4012 (N_4012,N_3656,N_3552);
nor U4013 (N_4013,N_3864,N_3510);
or U4014 (N_4014,N_3824,N_3823);
xnor U4015 (N_4015,N_3979,N_3584);
nand U4016 (N_4016,N_3546,N_3730);
or U4017 (N_4017,N_3673,N_3923);
nand U4018 (N_4018,N_3622,N_3952);
and U4019 (N_4019,N_3983,N_3514);
or U4020 (N_4020,N_3648,N_3654);
and U4021 (N_4021,N_3680,N_3598);
xor U4022 (N_4022,N_3586,N_3606);
nor U4023 (N_4023,N_3630,N_3812);
or U4024 (N_4024,N_3847,N_3624);
and U4025 (N_4025,N_3919,N_3926);
nand U4026 (N_4026,N_3711,N_3960);
xor U4027 (N_4027,N_3772,N_3808);
xnor U4028 (N_4028,N_3600,N_3653);
and U4029 (N_4029,N_3703,N_3597);
or U4030 (N_4030,N_3783,N_3671);
or U4031 (N_4031,N_3532,N_3924);
nand U4032 (N_4032,N_3935,N_3846);
nand U4033 (N_4033,N_3592,N_3658);
or U4034 (N_4034,N_3811,N_3617);
or U4035 (N_4035,N_3702,N_3799);
nor U4036 (N_4036,N_3647,N_3707);
and U4037 (N_4037,N_3740,N_3918);
xor U4038 (N_4038,N_3761,N_3986);
or U4039 (N_4039,N_3726,N_3844);
nor U4040 (N_4040,N_3564,N_3714);
or U4041 (N_4041,N_3791,N_3858);
and U4042 (N_4042,N_3501,N_3667);
and U4043 (N_4043,N_3975,N_3665);
and U4044 (N_4044,N_3523,N_3749);
or U4045 (N_4045,N_3742,N_3655);
nor U4046 (N_4046,N_3769,N_3838);
or U4047 (N_4047,N_3717,N_3992);
and U4048 (N_4048,N_3644,N_3976);
and U4049 (N_4049,N_3883,N_3745);
nor U4050 (N_4050,N_3694,N_3977);
nand U4051 (N_4051,N_3659,N_3775);
nor U4052 (N_4052,N_3618,N_3712);
or U4053 (N_4053,N_3569,N_3911);
nand U4054 (N_4054,N_3966,N_3943);
nand U4055 (N_4055,N_3932,N_3848);
and U4056 (N_4056,N_3785,N_3639);
or U4057 (N_4057,N_3596,N_3601);
nand U4058 (N_4058,N_3610,N_3965);
xnor U4059 (N_4059,N_3526,N_3857);
and U4060 (N_4060,N_3841,N_3732);
nor U4061 (N_4061,N_3879,N_3652);
xor U4062 (N_4062,N_3669,N_3743);
xor U4063 (N_4063,N_3651,N_3921);
nor U4064 (N_4064,N_3603,N_3562);
and U4065 (N_4065,N_3831,N_3663);
and U4066 (N_4066,N_3575,N_3794);
xor U4067 (N_4067,N_3987,N_3689);
xnor U4068 (N_4068,N_3942,N_3503);
nor U4069 (N_4069,N_3660,N_3643);
nor U4070 (N_4070,N_3578,N_3525);
nor U4071 (N_4071,N_3710,N_3507);
or U4072 (N_4072,N_3609,N_3733);
and U4073 (N_4073,N_3833,N_3922);
nor U4074 (N_4074,N_3716,N_3690);
nand U4075 (N_4075,N_3937,N_3566);
xnor U4076 (N_4076,N_3941,N_3642);
nand U4077 (N_4077,N_3884,N_3997);
or U4078 (N_4078,N_3538,N_3701);
nand U4079 (N_4079,N_3559,N_3688);
nor U4080 (N_4080,N_3885,N_3947);
xor U4081 (N_4081,N_3820,N_3551);
nor U4082 (N_4082,N_3756,N_3585);
nor U4083 (N_4083,N_3920,N_3563);
and U4084 (N_4084,N_3961,N_3777);
or U4085 (N_4085,N_3682,N_3678);
or U4086 (N_4086,N_3829,N_3948);
or U4087 (N_4087,N_3876,N_3872);
and U4088 (N_4088,N_3637,N_3500);
nand U4089 (N_4089,N_3780,N_3696);
or U4090 (N_4090,N_3999,N_3674);
and U4091 (N_4091,N_3891,N_3657);
nand U4092 (N_4092,N_3807,N_3955);
or U4093 (N_4093,N_3865,N_3721);
nand U4094 (N_4094,N_3629,N_3851);
or U4095 (N_4095,N_3543,N_3871);
nand U4096 (N_4096,N_3747,N_3760);
xnor U4097 (N_4097,N_3534,N_3905);
nand U4098 (N_4098,N_3778,N_3612);
or U4099 (N_4099,N_3593,N_3852);
and U4100 (N_4100,N_3684,N_3895);
nand U4101 (N_4101,N_3875,N_3813);
xor U4102 (N_4102,N_3902,N_3819);
nand U4103 (N_4103,N_3989,N_3542);
or U4104 (N_4104,N_3621,N_3560);
and U4105 (N_4105,N_3614,N_3509);
xor U4106 (N_4106,N_3513,N_3774);
nor U4107 (N_4107,N_3594,N_3540);
or U4108 (N_4108,N_3801,N_3832);
and U4109 (N_4109,N_3839,N_3927);
nor U4110 (N_4110,N_3615,N_3723);
and U4111 (N_4111,N_3754,N_3970);
nand U4112 (N_4112,N_3899,N_3972);
xnor U4113 (N_4113,N_3699,N_3840);
nor U4114 (N_4114,N_3530,N_3686);
xor U4115 (N_4115,N_3763,N_3539);
or U4116 (N_4116,N_3764,N_3816);
and U4117 (N_4117,N_3788,N_3632);
or U4118 (N_4118,N_3544,N_3913);
nand U4119 (N_4119,N_3928,N_3697);
xor U4120 (N_4120,N_3954,N_3693);
or U4121 (N_4121,N_3565,N_3555);
or U4122 (N_4122,N_3640,N_3504);
nand U4123 (N_4123,N_3963,N_3964);
nand U4124 (N_4124,N_3800,N_3611);
xor U4125 (N_4125,N_3568,N_3650);
or U4126 (N_4126,N_3589,N_3626);
nor U4127 (N_4127,N_3722,N_3587);
nor U4128 (N_4128,N_3623,N_3985);
or U4129 (N_4129,N_3825,N_3580);
xnor U4130 (N_4130,N_3641,N_3581);
nand U4131 (N_4131,N_3842,N_3925);
or U4132 (N_4132,N_3515,N_3725);
or U4133 (N_4133,N_3861,N_3616);
xor U4134 (N_4134,N_3815,N_3853);
nand U4135 (N_4135,N_3731,N_3765);
and U4136 (N_4136,N_3880,N_3636);
xnor U4137 (N_4137,N_3901,N_3933);
and U4138 (N_4138,N_3877,N_3506);
and U4139 (N_4139,N_3856,N_3792);
xnor U4140 (N_4140,N_3604,N_3508);
and U4141 (N_4141,N_3528,N_3670);
and U4142 (N_4142,N_3548,N_3784);
or U4143 (N_4143,N_3789,N_3962);
and U4144 (N_4144,N_3751,N_3531);
or U4145 (N_4145,N_3810,N_3557);
nand U4146 (N_4146,N_3634,N_3843);
xor U4147 (N_4147,N_3796,N_3571);
and U4148 (N_4148,N_3628,N_3599);
xnor U4149 (N_4149,N_3527,N_3958);
xnor U4150 (N_4150,N_3859,N_3991);
and U4151 (N_4151,N_3957,N_3638);
or U4152 (N_4152,N_3645,N_3524);
or U4153 (N_4153,N_3705,N_3582);
and U4154 (N_4154,N_3649,N_3625);
or U4155 (N_4155,N_3537,N_3814);
nand U4156 (N_4156,N_3519,N_3768);
or U4157 (N_4157,N_3967,N_3854);
or U4158 (N_4158,N_3945,N_3826);
or U4159 (N_4159,N_3698,N_3956);
nand U4160 (N_4160,N_3912,N_3520);
and U4161 (N_4161,N_3521,N_3862);
xnor U4162 (N_4162,N_3605,N_3929);
nand U4163 (N_4163,N_3867,N_3821);
nand U4164 (N_4164,N_3830,N_3556);
nand U4165 (N_4165,N_3770,N_3728);
xor U4166 (N_4166,N_3887,N_3809);
or U4167 (N_4167,N_3607,N_3909);
or U4168 (N_4168,N_3541,N_3619);
and U4169 (N_4169,N_3683,N_3974);
nand U4170 (N_4170,N_3720,N_3771);
nand U4171 (N_4171,N_3870,N_3904);
nand U4172 (N_4172,N_3767,N_3995);
and U4173 (N_4173,N_3662,N_3805);
nor U4174 (N_4174,N_3573,N_3668);
nor U4175 (N_4175,N_3817,N_3734);
xnor U4176 (N_4176,N_3691,N_3903);
nand U4177 (N_4177,N_3675,N_3822);
nand U4178 (N_4178,N_3836,N_3577);
nor U4179 (N_4179,N_3518,N_3969);
and U4180 (N_4180,N_3900,N_3971);
nor U4181 (N_4181,N_3939,N_3561);
and U4182 (N_4182,N_3766,N_3620);
nand U4183 (N_4183,N_3881,N_3549);
xnor U4184 (N_4184,N_3953,N_3572);
or U4185 (N_4185,N_3715,N_3511);
xnor U4186 (N_4186,N_3631,N_3738);
xor U4187 (N_4187,N_3994,N_3545);
nand U4188 (N_4188,N_3938,N_3874);
nor U4189 (N_4189,N_3984,N_3535);
and U4190 (N_4190,N_3746,N_3908);
nor U4191 (N_4191,N_3998,N_3661);
or U4192 (N_4192,N_3748,N_3798);
or U4193 (N_4193,N_3739,N_3752);
or U4194 (N_4194,N_3679,N_3906);
and U4195 (N_4195,N_3595,N_3827);
nor U4196 (N_4196,N_3635,N_3973);
and U4197 (N_4197,N_3773,N_3897);
and U4198 (N_4198,N_3550,N_3713);
xnor U4199 (N_4199,N_3672,N_3505);
xor U4200 (N_4200,N_3980,N_3898);
or U4201 (N_4201,N_3866,N_3759);
nand U4202 (N_4202,N_3978,N_3950);
or U4203 (N_4203,N_3529,N_3795);
xor U4204 (N_4204,N_3704,N_3804);
xnor U4205 (N_4205,N_3695,N_3949);
and U4206 (N_4206,N_3706,N_3516);
or U4207 (N_4207,N_3890,N_3588);
or U4208 (N_4208,N_3793,N_3522);
nor U4209 (N_4209,N_3646,N_3692);
and U4210 (N_4210,N_3786,N_3755);
nor U4211 (N_4211,N_3583,N_3931);
and U4212 (N_4212,N_3869,N_3737);
nand U4213 (N_4213,N_3934,N_3666);
nor U4214 (N_4214,N_3828,N_3762);
and U4215 (N_4215,N_3845,N_3888);
or U4216 (N_4216,N_3896,N_3996);
and U4217 (N_4217,N_3750,N_3835);
xnor U4218 (N_4218,N_3837,N_3802);
nand U4219 (N_4219,N_3893,N_3892);
nand U4220 (N_4220,N_3894,N_3917);
nor U4221 (N_4221,N_3944,N_3700);
and U4222 (N_4222,N_3787,N_3517);
or U4223 (N_4223,N_3993,N_3959);
xnor U4224 (N_4224,N_3803,N_3608);
xor U4225 (N_4225,N_3664,N_3554);
and U4226 (N_4226,N_3863,N_3834);
and U4227 (N_4227,N_3930,N_3736);
nor U4228 (N_4228,N_3790,N_3724);
and U4229 (N_4229,N_3744,N_3946);
or U4230 (N_4230,N_3613,N_3981);
nand U4231 (N_4231,N_3914,N_3602);
nand U4232 (N_4232,N_3849,N_3687);
or U4233 (N_4233,N_3855,N_3719);
and U4234 (N_4234,N_3533,N_3727);
xnor U4235 (N_4235,N_3677,N_3735);
nand U4236 (N_4236,N_3889,N_3579);
nand U4237 (N_4237,N_3633,N_3910);
nand U4238 (N_4238,N_3591,N_3502);
and U4239 (N_4239,N_3850,N_3915);
nor U4240 (N_4240,N_3982,N_3968);
and U4241 (N_4241,N_3709,N_3818);
xor U4242 (N_4242,N_3940,N_3718);
and U4243 (N_4243,N_3741,N_3729);
xor U4244 (N_4244,N_3681,N_3806);
nor U4245 (N_4245,N_3988,N_3873);
and U4246 (N_4246,N_3951,N_3547);
nand U4247 (N_4247,N_3990,N_3590);
xor U4248 (N_4248,N_3916,N_3860);
nand U4249 (N_4249,N_3558,N_3782);
xnor U4250 (N_4250,N_3922,N_3594);
nand U4251 (N_4251,N_3770,N_3734);
nand U4252 (N_4252,N_3769,N_3846);
xor U4253 (N_4253,N_3823,N_3936);
and U4254 (N_4254,N_3932,N_3761);
nor U4255 (N_4255,N_3705,N_3731);
and U4256 (N_4256,N_3839,N_3909);
and U4257 (N_4257,N_3711,N_3970);
nand U4258 (N_4258,N_3781,N_3922);
and U4259 (N_4259,N_3626,N_3635);
and U4260 (N_4260,N_3526,N_3675);
or U4261 (N_4261,N_3655,N_3769);
and U4262 (N_4262,N_3685,N_3503);
nand U4263 (N_4263,N_3952,N_3916);
xor U4264 (N_4264,N_3658,N_3551);
and U4265 (N_4265,N_3833,N_3865);
and U4266 (N_4266,N_3678,N_3616);
nor U4267 (N_4267,N_3759,N_3586);
xnor U4268 (N_4268,N_3925,N_3966);
xor U4269 (N_4269,N_3680,N_3685);
nand U4270 (N_4270,N_3699,N_3827);
nor U4271 (N_4271,N_3778,N_3905);
xnor U4272 (N_4272,N_3679,N_3977);
nand U4273 (N_4273,N_3721,N_3658);
nand U4274 (N_4274,N_3613,N_3859);
or U4275 (N_4275,N_3712,N_3884);
nor U4276 (N_4276,N_3536,N_3658);
xnor U4277 (N_4277,N_3571,N_3529);
xnor U4278 (N_4278,N_3509,N_3741);
nor U4279 (N_4279,N_3928,N_3631);
nand U4280 (N_4280,N_3786,N_3505);
nor U4281 (N_4281,N_3842,N_3593);
nor U4282 (N_4282,N_3630,N_3613);
nand U4283 (N_4283,N_3576,N_3540);
nor U4284 (N_4284,N_3620,N_3782);
xor U4285 (N_4285,N_3573,N_3809);
nor U4286 (N_4286,N_3677,N_3549);
nand U4287 (N_4287,N_3779,N_3781);
or U4288 (N_4288,N_3504,N_3935);
xor U4289 (N_4289,N_3879,N_3553);
nor U4290 (N_4290,N_3562,N_3757);
nand U4291 (N_4291,N_3899,N_3928);
nand U4292 (N_4292,N_3828,N_3900);
nand U4293 (N_4293,N_3930,N_3941);
nor U4294 (N_4294,N_3899,N_3525);
xnor U4295 (N_4295,N_3925,N_3623);
or U4296 (N_4296,N_3584,N_3524);
nor U4297 (N_4297,N_3675,N_3586);
or U4298 (N_4298,N_3504,N_3982);
xnor U4299 (N_4299,N_3577,N_3889);
nor U4300 (N_4300,N_3569,N_3913);
nor U4301 (N_4301,N_3662,N_3726);
or U4302 (N_4302,N_3578,N_3897);
and U4303 (N_4303,N_3927,N_3651);
or U4304 (N_4304,N_3936,N_3826);
nor U4305 (N_4305,N_3591,N_3853);
nor U4306 (N_4306,N_3682,N_3597);
xnor U4307 (N_4307,N_3805,N_3635);
or U4308 (N_4308,N_3794,N_3534);
or U4309 (N_4309,N_3892,N_3505);
or U4310 (N_4310,N_3955,N_3882);
nor U4311 (N_4311,N_3590,N_3910);
nand U4312 (N_4312,N_3882,N_3562);
nor U4313 (N_4313,N_3548,N_3968);
and U4314 (N_4314,N_3828,N_3731);
or U4315 (N_4315,N_3833,N_3885);
nor U4316 (N_4316,N_3664,N_3869);
or U4317 (N_4317,N_3561,N_3679);
nor U4318 (N_4318,N_3517,N_3506);
and U4319 (N_4319,N_3620,N_3745);
nor U4320 (N_4320,N_3514,N_3565);
or U4321 (N_4321,N_3709,N_3908);
or U4322 (N_4322,N_3697,N_3598);
nand U4323 (N_4323,N_3830,N_3581);
nand U4324 (N_4324,N_3809,N_3668);
xor U4325 (N_4325,N_3914,N_3833);
nor U4326 (N_4326,N_3993,N_3587);
or U4327 (N_4327,N_3717,N_3660);
nor U4328 (N_4328,N_3566,N_3876);
xor U4329 (N_4329,N_3901,N_3950);
nor U4330 (N_4330,N_3864,N_3807);
or U4331 (N_4331,N_3826,N_3873);
xnor U4332 (N_4332,N_3864,N_3550);
and U4333 (N_4333,N_3731,N_3853);
and U4334 (N_4334,N_3945,N_3916);
or U4335 (N_4335,N_3654,N_3792);
nor U4336 (N_4336,N_3643,N_3964);
nand U4337 (N_4337,N_3990,N_3748);
or U4338 (N_4338,N_3802,N_3944);
nand U4339 (N_4339,N_3850,N_3745);
nor U4340 (N_4340,N_3690,N_3659);
xor U4341 (N_4341,N_3894,N_3612);
xnor U4342 (N_4342,N_3980,N_3803);
nor U4343 (N_4343,N_3621,N_3968);
xnor U4344 (N_4344,N_3839,N_3798);
and U4345 (N_4345,N_3595,N_3677);
or U4346 (N_4346,N_3963,N_3992);
xor U4347 (N_4347,N_3805,N_3855);
and U4348 (N_4348,N_3815,N_3870);
nor U4349 (N_4349,N_3645,N_3985);
or U4350 (N_4350,N_3742,N_3582);
nand U4351 (N_4351,N_3581,N_3892);
nor U4352 (N_4352,N_3661,N_3773);
xor U4353 (N_4353,N_3618,N_3981);
and U4354 (N_4354,N_3688,N_3779);
nor U4355 (N_4355,N_3942,N_3665);
and U4356 (N_4356,N_3546,N_3758);
xor U4357 (N_4357,N_3999,N_3847);
nor U4358 (N_4358,N_3835,N_3738);
and U4359 (N_4359,N_3531,N_3905);
nand U4360 (N_4360,N_3540,N_3546);
nor U4361 (N_4361,N_3603,N_3647);
nand U4362 (N_4362,N_3700,N_3891);
nand U4363 (N_4363,N_3559,N_3584);
and U4364 (N_4364,N_3687,N_3789);
and U4365 (N_4365,N_3904,N_3766);
nor U4366 (N_4366,N_3753,N_3885);
or U4367 (N_4367,N_3634,N_3616);
or U4368 (N_4368,N_3631,N_3624);
xor U4369 (N_4369,N_3784,N_3852);
nor U4370 (N_4370,N_3502,N_3598);
or U4371 (N_4371,N_3542,N_3614);
xnor U4372 (N_4372,N_3586,N_3884);
nand U4373 (N_4373,N_3842,N_3733);
or U4374 (N_4374,N_3567,N_3533);
or U4375 (N_4375,N_3814,N_3918);
xor U4376 (N_4376,N_3611,N_3523);
xnor U4377 (N_4377,N_3824,N_3838);
or U4378 (N_4378,N_3874,N_3527);
nand U4379 (N_4379,N_3533,N_3873);
xnor U4380 (N_4380,N_3508,N_3531);
xor U4381 (N_4381,N_3926,N_3673);
and U4382 (N_4382,N_3750,N_3849);
xor U4383 (N_4383,N_3980,N_3845);
and U4384 (N_4384,N_3742,N_3626);
or U4385 (N_4385,N_3532,N_3553);
or U4386 (N_4386,N_3828,N_3775);
nand U4387 (N_4387,N_3694,N_3701);
nand U4388 (N_4388,N_3820,N_3713);
xor U4389 (N_4389,N_3585,N_3613);
and U4390 (N_4390,N_3786,N_3959);
or U4391 (N_4391,N_3946,N_3716);
and U4392 (N_4392,N_3562,N_3650);
nor U4393 (N_4393,N_3516,N_3736);
and U4394 (N_4394,N_3606,N_3667);
xor U4395 (N_4395,N_3687,N_3728);
and U4396 (N_4396,N_3607,N_3945);
nand U4397 (N_4397,N_3709,N_3937);
or U4398 (N_4398,N_3558,N_3905);
xnor U4399 (N_4399,N_3525,N_3685);
xor U4400 (N_4400,N_3844,N_3918);
xnor U4401 (N_4401,N_3609,N_3787);
nor U4402 (N_4402,N_3800,N_3725);
nor U4403 (N_4403,N_3648,N_3686);
nor U4404 (N_4404,N_3691,N_3538);
nand U4405 (N_4405,N_3550,N_3704);
nand U4406 (N_4406,N_3805,N_3786);
and U4407 (N_4407,N_3552,N_3678);
and U4408 (N_4408,N_3971,N_3567);
and U4409 (N_4409,N_3613,N_3958);
nor U4410 (N_4410,N_3999,N_3844);
or U4411 (N_4411,N_3863,N_3680);
nor U4412 (N_4412,N_3957,N_3892);
or U4413 (N_4413,N_3967,N_3549);
and U4414 (N_4414,N_3741,N_3604);
and U4415 (N_4415,N_3965,N_3982);
and U4416 (N_4416,N_3700,N_3536);
and U4417 (N_4417,N_3828,N_3623);
nand U4418 (N_4418,N_3609,N_3867);
or U4419 (N_4419,N_3796,N_3582);
or U4420 (N_4420,N_3816,N_3681);
and U4421 (N_4421,N_3504,N_3683);
xor U4422 (N_4422,N_3761,N_3701);
and U4423 (N_4423,N_3674,N_3776);
nor U4424 (N_4424,N_3565,N_3897);
or U4425 (N_4425,N_3945,N_3619);
xnor U4426 (N_4426,N_3902,N_3594);
nand U4427 (N_4427,N_3510,N_3937);
nand U4428 (N_4428,N_3637,N_3549);
nor U4429 (N_4429,N_3888,N_3954);
and U4430 (N_4430,N_3902,N_3658);
nand U4431 (N_4431,N_3976,N_3761);
and U4432 (N_4432,N_3714,N_3529);
xor U4433 (N_4433,N_3790,N_3661);
nand U4434 (N_4434,N_3724,N_3965);
or U4435 (N_4435,N_3506,N_3727);
nand U4436 (N_4436,N_3593,N_3723);
nor U4437 (N_4437,N_3989,N_3852);
or U4438 (N_4438,N_3717,N_3513);
and U4439 (N_4439,N_3524,N_3651);
xnor U4440 (N_4440,N_3518,N_3763);
nor U4441 (N_4441,N_3898,N_3873);
nor U4442 (N_4442,N_3765,N_3789);
nand U4443 (N_4443,N_3604,N_3693);
nand U4444 (N_4444,N_3880,N_3833);
nand U4445 (N_4445,N_3847,N_3833);
xnor U4446 (N_4446,N_3605,N_3871);
xnor U4447 (N_4447,N_3874,N_3606);
nand U4448 (N_4448,N_3833,N_3784);
nor U4449 (N_4449,N_3805,N_3529);
nand U4450 (N_4450,N_3704,N_3730);
xor U4451 (N_4451,N_3639,N_3931);
xor U4452 (N_4452,N_3685,N_3930);
nand U4453 (N_4453,N_3736,N_3982);
nand U4454 (N_4454,N_3572,N_3567);
or U4455 (N_4455,N_3732,N_3650);
nand U4456 (N_4456,N_3951,N_3716);
nor U4457 (N_4457,N_3726,N_3978);
nor U4458 (N_4458,N_3919,N_3523);
and U4459 (N_4459,N_3794,N_3868);
or U4460 (N_4460,N_3577,N_3533);
nand U4461 (N_4461,N_3779,N_3806);
xor U4462 (N_4462,N_3897,N_3651);
nand U4463 (N_4463,N_3839,N_3836);
or U4464 (N_4464,N_3989,N_3571);
xor U4465 (N_4465,N_3849,N_3774);
and U4466 (N_4466,N_3740,N_3980);
nor U4467 (N_4467,N_3615,N_3605);
xor U4468 (N_4468,N_3866,N_3854);
nor U4469 (N_4469,N_3501,N_3932);
nand U4470 (N_4470,N_3852,N_3954);
and U4471 (N_4471,N_3596,N_3801);
or U4472 (N_4472,N_3834,N_3724);
and U4473 (N_4473,N_3752,N_3742);
and U4474 (N_4474,N_3746,N_3564);
or U4475 (N_4475,N_3824,N_3548);
nor U4476 (N_4476,N_3829,N_3745);
and U4477 (N_4477,N_3640,N_3701);
and U4478 (N_4478,N_3834,N_3707);
xor U4479 (N_4479,N_3980,N_3934);
or U4480 (N_4480,N_3966,N_3844);
and U4481 (N_4481,N_3783,N_3851);
xor U4482 (N_4482,N_3538,N_3850);
nor U4483 (N_4483,N_3550,N_3722);
nor U4484 (N_4484,N_3533,N_3913);
and U4485 (N_4485,N_3699,N_3647);
xnor U4486 (N_4486,N_3595,N_3729);
nor U4487 (N_4487,N_3901,N_3982);
nor U4488 (N_4488,N_3849,N_3685);
nor U4489 (N_4489,N_3678,N_3593);
nand U4490 (N_4490,N_3644,N_3752);
or U4491 (N_4491,N_3545,N_3561);
nand U4492 (N_4492,N_3978,N_3793);
nor U4493 (N_4493,N_3666,N_3858);
xor U4494 (N_4494,N_3536,N_3528);
nand U4495 (N_4495,N_3507,N_3748);
nor U4496 (N_4496,N_3811,N_3910);
nand U4497 (N_4497,N_3735,N_3803);
nand U4498 (N_4498,N_3572,N_3800);
or U4499 (N_4499,N_3974,N_3680);
and U4500 (N_4500,N_4271,N_4483);
nand U4501 (N_4501,N_4036,N_4015);
or U4502 (N_4502,N_4112,N_4218);
nor U4503 (N_4503,N_4441,N_4259);
nor U4504 (N_4504,N_4233,N_4337);
nor U4505 (N_4505,N_4089,N_4330);
nand U4506 (N_4506,N_4003,N_4030);
and U4507 (N_4507,N_4047,N_4090);
xnor U4508 (N_4508,N_4215,N_4053);
nor U4509 (N_4509,N_4351,N_4202);
and U4510 (N_4510,N_4173,N_4125);
nor U4511 (N_4511,N_4139,N_4447);
and U4512 (N_4512,N_4050,N_4136);
or U4513 (N_4513,N_4087,N_4035);
nand U4514 (N_4514,N_4397,N_4041);
nand U4515 (N_4515,N_4379,N_4460);
and U4516 (N_4516,N_4414,N_4205);
or U4517 (N_4517,N_4170,N_4316);
or U4518 (N_4518,N_4282,N_4428);
or U4519 (N_4519,N_4383,N_4124);
xnor U4520 (N_4520,N_4308,N_4022);
xor U4521 (N_4521,N_4107,N_4189);
nor U4522 (N_4522,N_4426,N_4450);
and U4523 (N_4523,N_4115,N_4405);
and U4524 (N_4524,N_4315,N_4327);
and U4525 (N_4525,N_4048,N_4007);
xnor U4526 (N_4526,N_4395,N_4220);
or U4527 (N_4527,N_4241,N_4467);
xnor U4528 (N_4528,N_4250,N_4137);
or U4529 (N_4529,N_4438,N_4223);
and U4530 (N_4530,N_4019,N_4005);
nand U4531 (N_4531,N_4274,N_4355);
or U4532 (N_4532,N_4260,N_4341);
xnor U4533 (N_4533,N_4464,N_4208);
or U4534 (N_4534,N_4336,N_4407);
or U4535 (N_4535,N_4077,N_4066);
and U4536 (N_4536,N_4060,N_4265);
or U4537 (N_4537,N_4199,N_4443);
or U4538 (N_4538,N_4437,N_4054);
nand U4539 (N_4539,N_4143,N_4335);
nand U4540 (N_4540,N_4130,N_4479);
nand U4541 (N_4541,N_4458,N_4111);
xnor U4542 (N_4542,N_4180,N_4219);
nor U4543 (N_4543,N_4348,N_4404);
and U4544 (N_4544,N_4451,N_4142);
nor U4545 (N_4545,N_4377,N_4209);
nor U4546 (N_4546,N_4453,N_4364);
and U4547 (N_4547,N_4424,N_4197);
xnor U4548 (N_4548,N_4380,N_4301);
or U4549 (N_4549,N_4435,N_4062);
and U4550 (N_4550,N_4468,N_4042);
nor U4551 (N_4551,N_4221,N_4459);
xor U4552 (N_4552,N_4409,N_4293);
and U4553 (N_4553,N_4236,N_4242);
and U4554 (N_4554,N_4068,N_4349);
xor U4555 (N_4555,N_4346,N_4210);
or U4556 (N_4556,N_4084,N_4161);
and U4557 (N_4557,N_4224,N_4285);
nand U4558 (N_4558,N_4117,N_4491);
or U4559 (N_4559,N_4227,N_4363);
xor U4560 (N_4560,N_4328,N_4126);
or U4561 (N_4561,N_4080,N_4201);
and U4562 (N_4562,N_4389,N_4001);
and U4563 (N_4563,N_4385,N_4017);
nand U4564 (N_4564,N_4446,N_4040);
nand U4565 (N_4565,N_4332,N_4345);
xor U4566 (N_4566,N_4488,N_4278);
nor U4567 (N_4567,N_4486,N_4217);
xnor U4568 (N_4568,N_4171,N_4326);
nor U4569 (N_4569,N_4299,N_4454);
xor U4570 (N_4570,N_4413,N_4166);
nand U4571 (N_4571,N_4290,N_4081);
and U4572 (N_4572,N_4411,N_4403);
xor U4573 (N_4573,N_4246,N_4333);
nor U4574 (N_4574,N_4097,N_4418);
and U4575 (N_4575,N_4248,N_4088);
nand U4576 (N_4576,N_4267,N_4325);
and U4577 (N_4577,N_4181,N_4484);
or U4578 (N_4578,N_4469,N_4184);
nor U4579 (N_4579,N_4489,N_4046);
or U4580 (N_4580,N_4400,N_4334);
xor U4581 (N_4581,N_4319,N_4318);
nand U4582 (N_4582,N_4140,N_4465);
xnor U4583 (N_4583,N_4287,N_4113);
and U4584 (N_4584,N_4471,N_4212);
and U4585 (N_4585,N_4183,N_4381);
or U4586 (N_4586,N_4421,N_4422);
and U4587 (N_4587,N_4496,N_4127);
xor U4588 (N_4588,N_4045,N_4401);
nor U4589 (N_4589,N_4141,N_4416);
and U4590 (N_4590,N_4052,N_4474);
xnor U4591 (N_4591,N_4191,N_4207);
or U4592 (N_4592,N_4275,N_4195);
and U4593 (N_4593,N_4037,N_4268);
and U4594 (N_4594,N_4311,N_4371);
nand U4595 (N_4595,N_4376,N_4008);
or U4596 (N_4596,N_4024,N_4114);
and U4597 (N_4597,N_4059,N_4128);
or U4598 (N_4598,N_4091,N_4277);
and U4599 (N_4599,N_4366,N_4206);
or U4600 (N_4600,N_4235,N_4163);
or U4601 (N_4601,N_4322,N_4072);
xor U4602 (N_4602,N_4304,N_4386);
or U4603 (N_4603,N_4433,N_4432);
nand U4604 (N_4604,N_4306,N_4063);
nor U4605 (N_4605,N_4165,N_4034);
and U4606 (N_4606,N_4044,N_4070);
and U4607 (N_4607,N_4020,N_4425);
and U4608 (N_4608,N_4357,N_4211);
nand U4609 (N_4609,N_4410,N_4281);
or U4610 (N_4610,N_4300,N_4175);
xnor U4611 (N_4611,N_4495,N_4051);
nor U4612 (N_4612,N_4370,N_4138);
and U4613 (N_4613,N_4176,N_4204);
nand U4614 (N_4614,N_4382,N_4493);
nor U4615 (N_4615,N_4258,N_4134);
or U4616 (N_4616,N_4320,N_4083);
xor U4617 (N_4617,N_4058,N_4392);
and U4618 (N_4618,N_4384,N_4239);
xor U4619 (N_4619,N_4200,N_4093);
xor U4620 (N_4620,N_4490,N_4412);
or U4621 (N_4621,N_4192,N_4095);
nand U4622 (N_4622,N_4402,N_4108);
nand U4623 (N_4623,N_4198,N_4477);
xnor U4624 (N_4624,N_4359,N_4014);
and U4625 (N_4625,N_4261,N_4276);
nand U4626 (N_4626,N_4237,N_4043);
xnor U4627 (N_4627,N_4247,N_4478);
or U4628 (N_4628,N_4031,N_4156);
or U4629 (N_4629,N_4396,N_4362);
and U4630 (N_4630,N_4251,N_4073);
and U4631 (N_4631,N_4406,N_4029);
nor U4632 (N_4632,N_4178,N_4010);
xor U4633 (N_4633,N_4273,N_4360);
xnor U4634 (N_4634,N_4011,N_4297);
nor U4635 (N_4635,N_4427,N_4347);
nor U4636 (N_4636,N_4185,N_4481);
nor U4637 (N_4637,N_4436,N_4434);
xnor U4638 (N_4638,N_4033,N_4025);
nor U4639 (N_4639,N_4372,N_4118);
and U4640 (N_4640,N_4388,N_4155);
and U4641 (N_4641,N_4494,N_4294);
xnor U4642 (N_4642,N_4240,N_4172);
and U4643 (N_4643,N_4466,N_4309);
nand U4644 (N_4644,N_4295,N_4131);
nor U4645 (N_4645,N_4075,N_4462);
nand U4646 (N_4646,N_4016,N_4105);
xor U4647 (N_4647,N_4292,N_4196);
nand U4648 (N_4648,N_4028,N_4187);
nor U4649 (N_4649,N_4356,N_4009);
nand U4650 (N_4650,N_4120,N_4076);
or U4651 (N_4651,N_4103,N_4289);
xor U4652 (N_4652,N_4188,N_4487);
and U4653 (N_4653,N_4110,N_4182);
xnor U4654 (N_4654,N_4055,N_4094);
and U4655 (N_4655,N_4245,N_4461);
and U4656 (N_4656,N_4116,N_4321);
nand U4657 (N_4657,N_4123,N_4279);
nor U4658 (N_4658,N_4057,N_4352);
xor U4659 (N_4659,N_4027,N_4476);
or U4660 (N_4660,N_4312,N_4092);
xnor U4661 (N_4661,N_4012,N_4038);
xor U4662 (N_4662,N_4368,N_4317);
and U4663 (N_4663,N_4456,N_4144);
xnor U4664 (N_4664,N_4065,N_4106);
xor U4665 (N_4665,N_4148,N_4393);
and U4666 (N_4666,N_4339,N_4064);
nand U4667 (N_4667,N_4049,N_4067);
or U4668 (N_4668,N_4129,N_4152);
or U4669 (N_4669,N_4203,N_4169);
nand U4670 (N_4670,N_4498,N_4228);
nor U4671 (N_4671,N_4313,N_4154);
xor U4672 (N_4672,N_4291,N_4056);
xnor U4673 (N_4673,N_4442,N_4153);
or U4674 (N_4674,N_4002,N_4069);
or U4675 (N_4675,N_4249,N_4135);
or U4676 (N_4676,N_4305,N_4102);
or U4677 (N_4677,N_4263,N_4174);
nor U4678 (N_4678,N_4280,N_4485);
nor U4679 (N_4679,N_4415,N_4229);
nor U4680 (N_4680,N_4032,N_4082);
or U4681 (N_4681,N_4119,N_4147);
nor U4682 (N_4682,N_4146,N_4497);
xnor U4683 (N_4683,N_4096,N_4298);
and U4684 (N_4684,N_4310,N_4222);
nor U4685 (N_4685,N_4004,N_4071);
xnor U4686 (N_4686,N_4445,N_4286);
xnor U4687 (N_4687,N_4475,N_4365);
nor U4688 (N_4688,N_4499,N_4369);
or U4689 (N_4689,N_4225,N_4252);
xor U4690 (N_4690,N_4213,N_4344);
xor U4691 (N_4691,N_4266,N_4121);
or U4692 (N_4692,N_4230,N_4216);
and U4693 (N_4693,N_4018,N_4133);
nand U4694 (N_4694,N_4086,N_4100);
nor U4695 (N_4695,N_4079,N_4343);
xor U4696 (N_4696,N_4457,N_4423);
xor U4697 (N_4697,N_4440,N_4149);
xnor U4698 (N_4698,N_4253,N_4023);
and U4699 (N_4699,N_4179,N_4387);
xnor U4700 (N_4700,N_4394,N_4160);
xnor U4701 (N_4701,N_4162,N_4419);
xor U4702 (N_4702,N_4367,N_4270);
and U4703 (N_4703,N_4284,N_4302);
xor U4704 (N_4704,N_4000,N_4269);
nand U4705 (N_4705,N_4262,N_4323);
or U4706 (N_4706,N_4244,N_4391);
and U4707 (N_4707,N_4472,N_4439);
or U4708 (N_4708,N_4085,N_4420);
nor U4709 (N_4709,N_4303,N_4256);
or U4710 (N_4710,N_4482,N_4449);
nand U4711 (N_4711,N_4061,N_4272);
nor U4712 (N_4712,N_4296,N_4021);
or U4713 (N_4713,N_4340,N_4190);
and U4714 (N_4714,N_4226,N_4104);
or U4715 (N_4715,N_4350,N_4480);
xnor U4716 (N_4716,N_4399,N_4429);
or U4717 (N_4717,N_4232,N_4013);
and U4718 (N_4718,N_4492,N_4168);
nand U4719 (N_4719,N_4231,N_4452);
xnor U4720 (N_4720,N_4314,N_4238);
nor U4721 (N_4721,N_4358,N_4417);
or U4722 (N_4722,N_4448,N_4431);
nand U4723 (N_4723,N_4378,N_4444);
nand U4724 (N_4724,N_4074,N_4374);
nand U4725 (N_4725,N_4473,N_4283);
nand U4726 (N_4726,N_4157,N_4324);
nor U4727 (N_4727,N_4132,N_4194);
xnor U4728 (N_4728,N_4331,N_4122);
or U4729 (N_4729,N_4329,N_4430);
nand U4730 (N_4730,N_4307,N_4255);
or U4731 (N_4731,N_4158,N_4145);
nor U4732 (N_4732,N_4026,N_4234);
and U4733 (N_4733,N_4463,N_4455);
or U4734 (N_4734,N_4098,N_4159);
or U4735 (N_4735,N_4257,N_4109);
xnor U4736 (N_4736,N_4470,N_4186);
nand U4737 (N_4737,N_4078,N_4164);
nand U4738 (N_4738,N_4398,N_4193);
and U4739 (N_4739,N_4151,N_4264);
and U4740 (N_4740,N_4375,N_4243);
nand U4741 (N_4741,N_4150,N_4214);
or U4742 (N_4742,N_4361,N_4099);
nor U4743 (N_4743,N_4101,N_4254);
and U4744 (N_4744,N_4373,N_4342);
and U4745 (N_4745,N_4408,N_4006);
or U4746 (N_4746,N_4167,N_4338);
nand U4747 (N_4747,N_4390,N_4353);
xor U4748 (N_4748,N_4288,N_4354);
nand U4749 (N_4749,N_4177,N_4039);
or U4750 (N_4750,N_4366,N_4155);
nand U4751 (N_4751,N_4144,N_4196);
nor U4752 (N_4752,N_4000,N_4338);
or U4753 (N_4753,N_4381,N_4186);
or U4754 (N_4754,N_4082,N_4415);
nor U4755 (N_4755,N_4214,N_4266);
nand U4756 (N_4756,N_4471,N_4063);
nand U4757 (N_4757,N_4021,N_4346);
nand U4758 (N_4758,N_4049,N_4327);
nand U4759 (N_4759,N_4367,N_4491);
xor U4760 (N_4760,N_4193,N_4373);
xor U4761 (N_4761,N_4327,N_4121);
xor U4762 (N_4762,N_4326,N_4057);
xor U4763 (N_4763,N_4002,N_4429);
nand U4764 (N_4764,N_4320,N_4042);
nand U4765 (N_4765,N_4051,N_4228);
xor U4766 (N_4766,N_4347,N_4352);
nor U4767 (N_4767,N_4171,N_4460);
or U4768 (N_4768,N_4405,N_4439);
and U4769 (N_4769,N_4019,N_4412);
nand U4770 (N_4770,N_4080,N_4215);
xnor U4771 (N_4771,N_4094,N_4266);
nand U4772 (N_4772,N_4000,N_4212);
xor U4773 (N_4773,N_4474,N_4082);
nand U4774 (N_4774,N_4482,N_4293);
nor U4775 (N_4775,N_4040,N_4051);
xnor U4776 (N_4776,N_4331,N_4378);
xor U4777 (N_4777,N_4124,N_4259);
and U4778 (N_4778,N_4002,N_4062);
xnor U4779 (N_4779,N_4005,N_4122);
or U4780 (N_4780,N_4436,N_4002);
and U4781 (N_4781,N_4331,N_4189);
and U4782 (N_4782,N_4266,N_4287);
xnor U4783 (N_4783,N_4442,N_4018);
nand U4784 (N_4784,N_4145,N_4142);
nor U4785 (N_4785,N_4468,N_4203);
and U4786 (N_4786,N_4328,N_4285);
nand U4787 (N_4787,N_4194,N_4482);
or U4788 (N_4788,N_4495,N_4163);
or U4789 (N_4789,N_4439,N_4373);
or U4790 (N_4790,N_4295,N_4406);
nor U4791 (N_4791,N_4088,N_4145);
nor U4792 (N_4792,N_4060,N_4020);
or U4793 (N_4793,N_4401,N_4119);
nor U4794 (N_4794,N_4124,N_4353);
nor U4795 (N_4795,N_4362,N_4322);
nor U4796 (N_4796,N_4302,N_4211);
nor U4797 (N_4797,N_4138,N_4342);
nor U4798 (N_4798,N_4184,N_4444);
and U4799 (N_4799,N_4122,N_4475);
nor U4800 (N_4800,N_4183,N_4125);
nand U4801 (N_4801,N_4320,N_4466);
or U4802 (N_4802,N_4328,N_4037);
nand U4803 (N_4803,N_4331,N_4016);
or U4804 (N_4804,N_4242,N_4363);
or U4805 (N_4805,N_4478,N_4466);
nand U4806 (N_4806,N_4270,N_4146);
nand U4807 (N_4807,N_4246,N_4496);
xor U4808 (N_4808,N_4085,N_4320);
or U4809 (N_4809,N_4181,N_4492);
xnor U4810 (N_4810,N_4499,N_4341);
or U4811 (N_4811,N_4170,N_4078);
xnor U4812 (N_4812,N_4007,N_4292);
nor U4813 (N_4813,N_4287,N_4227);
and U4814 (N_4814,N_4229,N_4395);
nand U4815 (N_4815,N_4390,N_4239);
xnor U4816 (N_4816,N_4280,N_4168);
nand U4817 (N_4817,N_4196,N_4299);
nor U4818 (N_4818,N_4035,N_4386);
and U4819 (N_4819,N_4262,N_4472);
and U4820 (N_4820,N_4076,N_4073);
xnor U4821 (N_4821,N_4132,N_4471);
and U4822 (N_4822,N_4084,N_4284);
or U4823 (N_4823,N_4182,N_4119);
or U4824 (N_4824,N_4288,N_4215);
nor U4825 (N_4825,N_4426,N_4274);
and U4826 (N_4826,N_4253,N_4347);
or U4827 (N_4827,N_4211,N_4231);
and U4828 (N_4828,N_4354,N_4048);
or U4829 (N_4829,N_4002,N_4294);
or U4830 (N_4830,N_4467,N_4239);
nand U4831 (N_4831,N_4084,N_4268);
nand U4832 (N_4832,N_4215,N_4164);
or U4833 (N_4833,N_4099,N_4089);
xnor U4834 (N_4834,N_4169,N_4477);
or U4835 (N_4835,N_4359,N_4008);
nor U4836 (N_4836,N_4147,N_4380);
nor U4837 (N_4837,N_4027,N_4370);
nand U4838 (N_4838,N_4015,N_4441);
nand U4839 (N_4839,N_4204,N_4215);
nand U4840 (N_4840,N_4300,N_4162);
and U4841 (N_4841,N_4209,N_4397);
xor U4842 (N_4842,N_4019,N_4227);
and U4843 (N_4843,N_4317,N_4486);
or U4844 (N_4844,N_4189,N_4208);
nor U4845 (N_4845,N_4314,N_4215);
nor U4846 (N_4846,N_4071,N_4272);
nand U4847 (N_4847,N_4141,N_4160);
or U4848 (N_4848,N_4100,N_4418);
nor U4849 (N_4849,N_4066,N_4091);
or U4850 (N_4850,N_4354,N_4200);
xor U4851 (N_4851,N_4404,N_4468);
xor U4852 (N_4852,N_4053,N_4018);
nand U4853 (N_4853,N_4128,N_4380);
and U4854 (N_4854,N_4076,N_4272);
nor U4855 (N_4855,N_4299,N_4338);
nand U4856 (N_4856,N_4392,N_4247);
nand U4857 (N_4857,N_4447,N_4019);
xor U4858 (N_4858,N_4155,N_4295);
and U4859 (N_4859,N_4491,N_4334);
nand U4860 (N_4860,N_4192,N_4273);
xnor U4861 (N_4861,N_4167,N_4381);
xor U4862 (N_4862,N_4133,N_4303);
nand U4863 (N_4863,N_4433,N_4097);
xor U4864 (N_4864,N_4054,N_4112);
xor U4865 (N_4865,N_4218,N_4290);
nor U4866 (N_4866,N_4288,N_4253);
and U4867 (N_4867,N_4144,N_4411);
nor U4868 (N_4868,N_4269,N_4346);
nor U4869 (N_4869,N_4042,N_4325);
and U4870 (N_4870,N_4201,N_4271);
xor U4871 (N_4871,N_4167,N_4173);
and U4872 (N_4872,N_4385,N_4214);
xor U4873 (N_4873,N_4207,N_4441);
nand U4874 (N_4874,N_4009,N_4446);
nor U4875 (N_4875,N_4008,N_4444);
and U4876 (N_4876,N_4051,N_4431);
and U4877 (N_4877,N_4103,N_4431);
nand U4878 (N_4878,N_4203,N_4478);
and U4879 (N_4879,N_4066,N_4035);
nor U4880 (N_4880,N_4095,N_4234);
or U4881 (N_4881,N_4467,N_4381);
nand U4882 (N_4882,N_4217,N_4352);
or U4883 (N_4883,N_4273,N_4260);
or U4884 (N_4884,N_4334,N_4398);
nor U4885 (N_4885,N_4264,N_4043);
or U4886 (N_4886,N_4306,N_4266);
xnor U4887 (N_4887,N_4308,N_4366);
nor U4888 (N_4888,N_4008,N_4193);
nand U4889 (N_4889,N_4377,N_4314);
nand U4890 (N_4890,N_4414,N_4166);
nand U4891 (N_4891,N_4210,N_4156);
nor U4892 (N_4892,N_4156,N_4074);
nor U4893 (N_4893,N_4175,N_4059);
and U4894 (N_4894,N_4137,N_4315);
and U4895 (N_4895,N_4262,N_4008);
nand U4896 (N_4896,N_4436,N_4199);
nand U4897 (N_4897,N_4244,N_4394);
or U4898 (N_4898,N_4062,N_4175);
nor U4899 (N_4899,N_4230,N_4187);
xor U4900 (N_4900,N_4221,N_4097);
nor U4901 (N_4901,N_4389,N_4032);
nor U4902 (N_4902,N_4235,N_4275);
or U4903 (N_4903,N_4167,N_4388);
xnor U4904 (N_4904,N_4010,N_4482);
nand U4905 (N_4905,N_4089,N_4148);
or U4906 (N_4906,N_4170,N_4167);
or U4907 (N_4907,N_4067,N_4043);
and U4908 (N_4908,N_4433,N_4166);
and U4909 (N_4909,N_4346,N_4133);
nand U4910 (N_4910,N_4114,N_4067);
nand U4911 (N_4911,N_4336,N_4428);
xnor U4912 (N_4912,N_4190,N_4325);
nand U4913 (N_4913,N_4391,N_4073);
nand U4914 (N_4914,N_4098,N_4490);
and U4915 (N_4915,N_4373,N_4323);
nor U4916 (N_4916,N_4293,N_4233);
xor U4917 (N_4917,N_4374,N_4045);
or U4918 (N_4918,N_4373,N_4028);
and U4919 (N_4919,N_4118,N_4367);
and U4920 (N_4920,N_4200,N_4276);
and U4921 (N_4921,N_4435,N_4042);
nand U4922 (N_4922,N_4044,N_4065);
and U4923 (N_4923,N_4447,N_4131);
nor U4924 (N_4924,N_4250,N_4309);
xor U4925 (N_4925,N_4225,N_4103);
xnor U4926 (N_4926,N_4043,N_4330);
nand U4927 (N_4927,N_4088,N_4487);
and U4928 (N_4928,N_4282,N_4165);
nor U4929 (N_4929,N_4184,N_4426);
nand U4930 (N_4930,N_4044,N_4407);
xor U4931 (N_4931,N_4247,N_4464);
or U4932 (N_4932,N_4219,N_4431);
and U4933 (N_4933,N_4121,N_4412);
xnor U4934 (N_4934,N_4409,N_4392);
or U4935 (N_4935,N_4127,N_4409);
xnor U4936 (N_4936,N_4136,N_4478);
nor U4937 (N_4937,N_4347,N_4368);
xor U4938 (N_4938,N_4259,N_4063);
or U4939 (N_4939,N_4267,N_4329);
xor U4940 (N_4940,N_4308,N_4293);
and U4941 (N_4941,N_4093,N_4283);
xnor U4942 (N_4942,N_4105,N_4109);
or U4943 (N_4943,N_4303,N_4062);
xnor U4944 (N_4944,N_4308,N_4075);
xnor U4945 (N_4945,N_4168,N_4230);
xnor U4946 (N_4946,N_4009,N_4132);
and U4947 (N_4947,N_4315,N_4130);
and U4948 (N_4948,N_4436,N_4112);
or U4949 (N_4949,N_4375,N_4073);
nand U4950 (N_4950,N_4287,N_4148);
xnor U4951 (N_4951,N_4136,N_4185);
xnor U4952 (N_4952,N_4283,N_4155);
nand U4953 (N_4953,N_4348,N_4442);
nand U4954 (N_4954,N_4463,N_4307);
or U4955 (N_4955,N_4473,N_4135);
nand U4956 (N_4956,N_4057,N_4257);
xnor U4957 (N_4957,N_4405,N_4381);
or U4958 (N_4958,N_4153,N_4411);
and U4959 (N_4959,N_4277,N_4027);
or U4960 (N_4960,N_4126,N_4425);
or U4961 (N_4961,N_4091,N_4144);
nand U4962 (N_4962,N_4306,N_4369);
nor U4963 (N_4963,N_4433,N_4389);
and U4964 (N_4964,N_4244,N_4468);
nor U4965 (N_4965,N_4071,N_4396);
xor U4966 (N_4966,N_4061,N_4337);
and U4967 (N_4967,N_4252,N_4033);
nor U4968 (N_4968,N_4031,N_4003);
and U4969 (N_4969,N_4105,N_4432);
xor U4970 (N_4970,N_4280,N_4161);
nand U4971 (N_4971,N_4312,N_4216);
and U4972 (N_4972,N_4194,N_4315);
nand U4973 (N_4973,N_4305,N_4071);
nor U4974 (N_4974,N_4258,N_4066);
nor U4975 (N_4975,N_4128,N_4034);
and U4976 (N_4976,N_4348,N_4131);
and U4977 (N_4977,N_4442,N_4036);
nand U4978 (N_4978,N_4043,N_4462);
or U4979 (N_4979,N_4109,N_4172);
nand U4980 (N_4980,N_4429,N_4080);
nor U4981 (N_4981,N_4287,N_4338);
or U4982 (N_4982,N_4164,N_4200);
nor U4983 (N_4983,N_4335,N_4258);
nand U4984 (N_4984,N_4170,N_4123);
nand U4985 (N_4985,N_4368,N_4190);
or U4986 (N_4986,N_4331,N_4134);
xnor U4987 (N_4987,N_4368,N_4137);
and U4988 (N_4988,N_4226,N_4148);
and U4989 (N_4989,N_4128,N_4422);
nand U4990 (N_4990,N_4345,N_4160);
xnor U4991 (N_4991,N_4274,N_4074);
nor U4992 (N_4992,N_4102,N_4093);
or U4993 (N_4993,N_4218,N_4375);
and U4994 (N_4994,N_4014,N_4367);
xnor U4995 (N_4995,N_4387,N_4039);
or U4996 (N_4996,N_4318,N_4383);
and U4997 (N_4997,N_4345,N_4479);
xor U4998 (N_4998,N_4013,N_4149);
or U4999 (N_4999,N_4110,N_4444);
and U5000 (N_5000,N_4655,N_4812);
and U5001 (N_5001,N_4551,N_4708);
nor U5002 (N_5002,N_4790,N_4933);
and U5003 (N_5003,N_4903,N_4908);
and U5004 (N_5004,N_4777,N_4578);
nor U5005 (N_5005,N_4746,N_4773);
and U5006 (N_5006,N_4756,N_4536);
or U5007 (N_5007,N_4652,N_4709);
or U5008 (N_5008,N_4909,N_4654);
nand U5009 (N_5009,N_4723,N_4891);
nor U5010 (N_5010,N_4555,N_4695);
or U5011 (N_5011,N_4941,N_4711);
nor U5012 (N_5012,N_4693,N_4775);
xor U5013 (N_5013,N_4576,N_4607);
xor U5014 (N_5014,N_4680,N_4798);
and U5015 (N_5015,N_4806,N_4947);
nor U5016 (N_5016,N_4960,N_4689);
and U5017 (N_5017,N_4519,N_4651);
nor U5018 (N_5018,N_4615,N_4575);
xor U5019 (N_5019,N_4939,N_4946);
nor U5020 (N_5020,N_4740,N_4841);
and U5021 (N_5021,N_4938,N_4915);
nor U5022 (N_5022,N_4787,N_4727);
nor U5023 (N_5023,N_4610,N_4818);
xnor U5024 (N_5024,N_4816,N_4644);
and U5025 (N_5025,N_4601,N_4596);
nor U5026 (N_5026,N_4882,N_4999);
xor U5027 (N_5027,N_4843,N_4801);
nand U5028 (N_5028,N_4972,N_4686);
or U5029 (N_5029,N_4511,N_4623);
xnor U5030 (N_5030,N_4550,N_4949);
and U5031 (N_5031,N_4640,N_4966);
and U5032 (N_5032,N_4823,N_4774);
and U5033 (N_5033,N_4910,N_4572);
and U5034 (N_5034,N_4687,N_4547);
and U5035 (N_5035,N_4884,N_4921);
nor U5036 (N_5036,N_4898,N_4600);
nor U5037 (N_5037,N_4760,N_4870);
xnor U5038 (N_5038,N_4864,N_4824);
nor U5039 (N_5039,N_4763,N_4583);
nand U5040 (N_5040,N_4735,N_4957);
nor U5041 (N_5041,N_4567,N_4769);
nand U5042 (N_5042,N_4524,N_4937);
and U5043 (N_5043,N_4795,N_4671);
and U5044 (N_5044,N_4805,N_4876);
or U5045 (N_5045,N_4704,N_4764);
and U5046 (N_5046,N_4803,N_4815);
nor U5047 (N_5047,N_4720,N_4762);
and U5048 (N_5048,N_4565,N_4658);
xnor U5049 (N_5049,N_4842,N_4588);
xnor U5050 (N_5050,N_4845,N_4566);
and U5051 (N_5051,N_4526,N_4712);
and U5052 (N_5052,N_4970,N_4594);
nand U5053 (N_5053,N_4512,N_4827);
nand U5054 (N_5054,N_4800,N_4617);
xor U5055 (N_5055,N_4584,N_4962);
nor U5056 (N_5056,N_4643,N_4673);
nand U5057 (N_5057,N_4901,N_4974);
nor U5058 (N_5058,N_4515,N_4809);
xnor U5059 (N_5059,N_4782,N_4753);
xor U5060 (N_5060,N_4859,N_4563);
or U5061 (N_5061,N_4589,N_4844);
and U5062 (N_5062,N_4622,N_4544);
and U5063 (N_5063,N_4558,N_4825);
nand U5064 (N_5064,N_4591,N_4685);
nor U5065 (N_5065,N_4675,N_4948);
nand U5066 (N_5066,N_4540,N_4732);
and U5067 (N_5067,N_4579,N_4721);
nand U5068 (N_5068,N_4635,N_4819);
xnor U5069 (N_5069,N_4885,N_4913);
or U5070 (N_5070,N_4780,N_4666);
nor U5071 (N_5071,N_4715,N_4742);
or U5072 (N_5072,N_4877,N_4771);
nor U5073 (N_5073,N_4923,N_4628);
xor U5074 (N_5074,N_4724,N_4697);
xnor U5075 (N_5075,N_4706,N_4902);
nor U5076 (N_5076,N_4860,N_4595);
nand U5077 (N_5077,N_4924,N_4976);
nand U5078 (N_5078,N_4945,N_4529);
nor U5079 (N_5079,N_4552,N_4707);
nand U5080 (N_5080,N_4837,N_4872);
nor U5081 (N_5081,N_4821,N_4955);
nor U5082 (N_5082,N_4922,N_4883);
or U5083 (N_5083,N_4672,N_4678);
and U5084 (N_5084,N_4919,N_4554);
and U5085 (N_5085,N_4832,N_4730);
nor U5086 (N_5086,N_4533,N_4621);
nor U5087 (N_5087,N_4772,N_4839);
and U5088 (N_5088,N_4814,N_4692);
nor U5089 (N_5089,N_4542,N_4779);
nand U5090 (N_5090,N_4630,N_4609);
and U5091 (N_5091,N_4887,N_4703);
and U5092 (N_5092,N_4810,N_4507);
and U5093 (N_5093,N_4574,N_4875);
xnor U5094 (N_5094,N_4789,N_4766);
and U5095 (N_5095,N_4690,N_4797);
or U5096 (N_5096,N_4539,N_4549);
xnor U5097 (N_5097,N_4684,N_4513);
or U5098 (N_5098,N_4835,N_4577);
or U5099 (N_5099,N_4783,N_4784);
or U5100 (N_5100,N_4562,N_4770);
nand U5101 (N_5101,N_4995,N_4627);
nor U5102 (N_5102,N_4696,N_4954);
and U5103 (N_5103,N_4855,N_4847);
nand U5104 (N_5104,N_4699,N_4604);
or U5105 (N_5105,N_4813,N_4722);
or U5106 (N_5106,N_4889,N_4647);
and U5107 (N_5107,N_4807,N_4664);
or U5108 (N_5108,N_4639,N_4556);
or U5109 (N_5109,N_4571,N_4603);
xnor U5110 (N_5110,N_4765,N_4940);
xor U5111 (N_5111,N_4900,N_4679);
nand U5112 (N_5112,N_4963,N_4811);
nor U5113 (N_5113,N_4713,N_4971);
nand U5114 (N_5114,N_4525,N_4527);
or U5115 (N_5115,N_4590,N_4659);
and U5116 (N_5116,N_4920,N_4633);
nand U5117 (N_5117,N_4848,N_4657);
nand U5118 (N_5118,N_4983,N_4642);
nand U5119 (N_5119,N_4904,N_4559);
or U5120 (N_5120,N_4869,N_4934);
nor U5121 (N_5121,N_4616,N_4613);
nand U5122 (N_5122,N_4698,N_4858);
and U5123 (N_5123,N_4660,N_4996);
xnor U5124 (N_5124,N_4873,N_4820);
nor U5125 (N_5125,N_4614,N_4984);
nand U5126 (N_5126,N_4865,N_4881);
nor U5127 (N_5127,N_4737,N_4880);
or U5128 (N_5128,N_4896,N_4978);
nand U5129 (N_5129,N_4537,N_4929);
nand U5130 (N_5130,N_4928,N_4927);
or U5131 (N_5131,N_4592,N_4907);
nand U5132 (N_5132,N_4930,N_4850);
or U5133 (N_5133,N_4674,N_4528);
or U5134 (N_5134,N_4761,N_4667);
nand U5135 (N_5135,N_4645,N_4629);
nor U5136 (N_5136,N_4638,N_4759);
or U5137 (N_5137,N_4582,N_4767);
or U5138 (N_5138,N_4943,N_4854);
or U5139 (N_5139,N_4662,N_4979);
and U5140 (N_5140,N_4743,N_4866);
or U5141 (N_5141,N_4799,N_4792);
or U5142 (N_5142,N_4535,N_4980);
nand U5143 (N_5143,N_4653,N_4997);
or U5144 (N_5144,N_4606,N_4951);
nand U5145 (N_5145,N_4977,N_4959);
or U5146 (N_5146,N_4874,N_4998);
xor U5147 (N_5147,N_4969,N_4587);
or U5148 (N_5148,N_4681,N_4822);
nor U5149 (N_5149,N_4916,N_4586);
nand U5150 (N_5150,N_4833,N_4725);
nand U5151 (N_5151,N_4729,N_4502);
or U5152 (N_5152,N_4936,N_4501);
xor U5153 (N_5153,N_4736,N_4534);
nand U5154 (N_5154,N_4700,N_4856);
or U5155 (N_5155,N_4750,N_4619);
and U5156 (N_5156,N_4669,N_4993);
xor U5157 (N_5157,N_4776,N_4986);
nor U5158 (N_5158,N_4985,N_4961);
or U5159 (N_5159,N_4744,N_4503);
and U5160 (N_5160,N_4702,N_4905);
and U5161 (N_5161,N_4925,N_4718);
xor U5162 (N_5162,N_4886,N_4989);
and U5163 (N_5163,N_4830,N_4620);
nor U5164 (N_5164,N_4516,N_4717);
nor U5165 (N_5165,N_4863,N_4661);
xor U5166 (N_5166,N_4768,N_4817);
and U5167 (N_5167,N_4836,N_4500);
nor U5168 (N_5168,N_4530,N_4808);
xor U5169 (N_5169,N_4625,N_4935);
nand U5170 (N_5170,N_4705,N_4506);
nor U5171 (N_5171,N_4982,N_4593);
or U5172 (N_5172,N_4992,N_4981);
nor U5173 (N_5173,N_4612,N_4701);
or U5174 (N_5174,N_4747,N_4597);
nor U5175 (N_5175,N_4553,N_4714);
nand U5176 (N_5176,N_4758,N_4520);
and U5177 (N_5177,N_4911,N_4650);
and U5178 (N_5178,N_4956,N_4605);
nor U5179 (N_5179,N_4531,N_4670);
or U5180 (N_5180,N_4560,N_4570);
xnor U5181 (N_5181,N_4975,N_4888);
nor U5182 (N_5182,N_4508,N_4834);
nor U5183 (N_5183,N_4726,N_4788);
or U5184 (N_5184,N_4716,N_4546);
nand U5185 (N_5185,N_4942,N_4548);
xnor U5186 (N_5186,N_4990,N_4618);
or U5187 (N_5187,N_4853,N_4755);
nand U5188 (N_5188,N_4794,N_4532);
and U5189 (N_5189,N_4682,N_4781);
nor U5190 (N_5190,N_4741,N_4793);
nand U5191 (N_5191,N_4646,N_4879);
xnor U5192 (N_5192,N_4912,N_4523);
or U5193 (N_5193,N_4757,N_4624);
nor U5194 (N_5194,N_4867,N_4778);
or U5195 (N_5195,N_4952,N_4611);
or U5196 (N_5196,N_4663,N_4829);
nor U5197 (N_5197,N_4892,N_4688);
or U5198 (N_5198,N_4656,N_4754);
nor U5199 (N_5199,N_4958,N_4917);
nand U5200 (N_5200,N_4973,N_4895);
nand U5201 (N_5201,N_4918,N_4564);
and U5202 (N_5202,N_4668,N_4541);
nand U5203 (N_5203,N_4505,N_4846);
nor U5204 (N_5204,N_4509,N_4849);
nand U5205 (N_5205,N_4994,N_4878);
nand U5206 (N_5206,N_4785,N_4950);
nor U5207 (N_5207,N_4944,N_4521);
nor U5208 (N_5208,N_4557,N_4738);
xor U5209 (N_5209,N_4862,N_4665);
xor U5210 (N_5210,N_4648,N_4828);
and U5211 (N_5211,N_4719,N_4899);
xor U5212 (N_5212,N_4522,N_4691);
or U5213 (N_5213,N_4634,N_4510);
or U5214 (N_5214,N_4641,N_4987);
xnor U5215 (N_5215,N_4517,N_4840);
and U5216 (N_5216,N_4677,N_4543);
or U5217 (N_5217,N_4804,N_4857);
xnor U5218 (N_5218,N_4599,N_4893);
nor U5219 (N_5219,N_4626,N_4752);
and U5220 (N_5220,N_4731,N_4632);
xor U5221 (N_5221,N_4964,N_4580);
xnor U5222 (N_5222,N_4561,N_4897);
nor U5223 (N_5223,N_4676,N_4786);
nor U5224 (N_5224,N_4637,N_4868);
nand U5225 (N_5225,N_4796,N_4991);
nor U5226 (N_5226,N_4728,N_4545);
xor U5227 (N_5227,N_4852,N_4931);
and U5228 (N_5228,N_4926,N_4733);
or U5229 (N_5229,N_4710,N_4518);
nor U5230 (N_5230,N_4802,N_4636);
xnor U5231 (N_5231,N_4683,N_4861);
and U5232 (N_5232,N_4838,N_4932);
and U5233 (N_5233,N_4953,N_4608);
and U5234 (N_5234,N_4631,N_4649);
and U5235 (N_5235,N_4573,N_4514);
and U5236 (N_5236,N_4748,N_4890);
nand U5237 (N_5237,N_4826,N_4967);
nor U5238 (N_5238,N_4569,N_4585);
nand U5239 (N_5239,N_4851,N_4504);
nor U5240 (N_5240,N_4751,N_4739);
nor U5241 (N_5241,N_4749,N_4538);
or U5242 (N_5242,N_4602,N_4871);
and U5243 (N_5243,N_4894,N_4968);
and U5244 (N_5244,N_4598,N_4694);
xnor U5245 (N_5245,N_4988,N_4914);
and U5246 (N_5246,N_4791,N_4568);
or U5247 (N_5247,N_4965,N_4745);
and U5248 (N_5248,N_4581,N_4831);
and U5249 (N_5249,N_4906,N_4734);
nand U5250 (N_5250,N_4901,N_4804);
and U5251 (N_5251,N_4587,N_4875);
nor U5252 (N_5252,N_4976,N_4831);
and U5253 (N_5253,N_4697,N_4763);
xnor U5254 (N_5254,N_4806,N_4812);
nand U5255 (N_5255,N_4536,N_4939);
nand U5256 (N_5256,N_4597,N_4907);
nand U5257 (N_5257,N_4851,N_4828);
xnor U5258 (N_5258,N_4843,N_4900);
nand U5259 (N_5259,N_4574,N_4605);
xnor U5260 (N_5260,N_4660,N_4569);
nand U5261 (N_5261,N_4657,N_4591);
and U5262 (N_5262,N_4936,N_4945);
and U5263 (N_5263,N_4839,N_4757);
and U5264 (N_5264,N_4922,N_4758);
nor U5265 (N_5265,N_4765,N_4950);
xor U5266 (N_5266,N_4942,N_4975);
and U5267 (N_5267,N_4827,N_4899);
xnor U5268 (N_5268,N_4799,N_4806);
xnor U5269 (N_5269,N_4571,N_4977);
and U5270 (N_5270,N_4668,N_4589);
xnor U5271 (N_5271,N_4844,N_4559);
nand U5272 (N_5272,N_4724,N_4548);
and U5273 (N_5273,N_4730,N_4662);
or U5274 (N_5274,N_4602,N_4874);
xnor U5275 (N_5275,N_4961,N_4595);
nor U5276 (N_5276,N_4772,N_4656);
or U5277 (N_5277,N_4801,N_4946);
and U5278 (N_5278,N_4888,N_4704);
xor U5279 (N_5279,N_4603,N_4709);
xnor U5280 (N_5280,N_4527,N_4669);
and U5281 (N_5281,N_4868,N_4556);
nand U5282 (N_5282,N_4767,N_4540);
or U5283 (N_5283,N_4582,N_4835);
and U5284 (N_5284,N_4793,N_4592);
or U5285 (N_5285,N_4748,N_4625);
nor U5286 (N_5286,N_4663,N_4560);
or U5287 (N_5287,N_4500,N_4684);
xor U5288 (N_5288,N_4788,N_4786);
nor U5289 (N_5289,N_4558,N_4845);
and U5290 (N_5290,N_4830,N_4713);
and U5291 (N_5291,N_4901,N_4559);
or U5292 (N_5292,N_4657,N_4514);
or U5293 (N_5293,N_4661,N_4681);
nand U5294 (N_5294,N_4652,N_4571);
nor U5295 (N_5295,N_4661,N_4608);
nor U5296 (N_5296,N_4836,N_4922);
and U5297 (N_5297,N_4921,N_4585);
xor U5298 (N_5298,N_4919,N_4905);
and U5299 (N_5299,N_4978,N_4680);
nand U5300 (N_5300,N_4814,N_4773);
nor U5301 (N_5301,N_4760,N_4753);
and U5302 (N_5302,N_4994,N_4762);
nor U5303 (N_5303,N_4904,N_4917);
nor U5304 (N_5304,N_4797,N_4761);
nand U5305 (N_5305,N_4702,N_4647);
xnor U5306 (N_5306,N_4973,N_4787);
and U5307 (N_5307,N_4728,N_4702);
nor U5308 (N_5308,N_4789,N_4811);
xnor U5309 (N_5309,N_4850,N_4546);
xor U5310 (N_5310,N_4856,N_4847);
and U5311 (N_5311,N_4990,N_4665);
nand U5312 (N_5312,N_4871,N_4804);
and U5313 (N_5313,N_4654,N_4921);
xor U5314 (N_5314,N_4503,N_4754);
or U5315 (N_5315,N_4551,N_4980);
nand U5316 (N_5316,N_4845,N_4736);
or U5317 (N_5317,N_4781,N_4958);
and U5318 (N_5318,N_4658,N_4970);
nor U5319 (N_5319,N_4841,N_4902);
nor U5320 (N_5320,N_4892,N_4998);
xor U5321 (N_5321,N_4893,N_4885);
nand U5322 (N_5322,N_4797,N_4560);
nor U5323 (N_5323,N_4689,N_4707);
and U5324 (N_5324,N_4636,N_4979);
or U5325 (N_5325,N_4902,N_4548);
nand U5326 (N_5326,N_4720,N_4969);
and U5327 (N_5327,N_4536,N_4914);
and U5328 (N_5328,N_4802,N_4911);
nor U5329 (N_5329,N_4876,N_4954);
or U5330 (N_5330,N_4928,N_4931);
or U5331 (N_5331,N_4519,N_4828);
nor U5332 (N_5332,N_4943,N_4675);
xor U5333 (N_5333,N_4697,N_4576);
xor U5334 (N_5334,N_4605,N_4878);
xor U5335 (N_5335,N_4508,N_4908);
xnor U5336 (N_5336,N_4586,N_4530);
or U5337 (N_5337,N_4605,N_4704);
xnor U5338 (N_5338,N_4946,N_4927);
or U5339 (N_5339,N_4757,N_4592);
nor U5340 (N_5340,N_4544,N_4745);
xnor U5341 (N_5341,N_4934,N_4898);
xnor U5342 (N_5342,N_4541,N_4885);
or U5343 (N_5343,N_4683,N_4782);
or U5344 (N_5344,N_4644,N_4578);
nor U5345 (N_5345,N_4993,N_4989);
xor U5346 (N_5346,N_4768,N_4941);
or U5347 (N_5347,N_4611,N_4713);
and U5348 (N_5348,N_4908,N_4562);
and U5349 (N_5349,N_4596,N_4944);
nor U5350 (N_5350,N_4692,N_4800);
nor U5351 (N_5351,N_4931,N_4881);
nor U5352 (N_5352,N_4966,N_4814);
nand U5353 (N_5353,N_4956,N_4940);
nand U5354 (N_5354,N_4709,N_4606);
xnor U5355 (N_5355,N_4870,N_4976);
nor U5356 (N_5356,N_4537,N_4782);
nor U5357 (N_5357,N_4617,N_4860);
xor U5358 (N_5358,N_4580,N_4671);
and U5359 (N_5359,N_4678,N_4865);
xor U5360 (N_5360,N_4546,N_4889);
nand U5361 (N_5361,N_4648,N_4940);
xnor U5362 (N_5362,N_4672,N_4515);
nor U5363 (N_5363,N_4682,N_4848);
or U5364 (N_5364,N_4772,N_4986);
nand U5365 (N_5365,N_4718,N_4997);
nor U5366 (N_5366,N_4889,N_4855);
xor U5367 (N_5367,N_4544,N_4829);
or U5368 (N_5368,N_4727,N_4792);
or U5369 (N_5369,N_4870,N_4659);
nand U5370 (N_5370,N_4620,N_4534);
or U5371 (N_5371,N_4861,N_4520);
xnor U5372 (N_5372,N_4733,N_4564);
or U5373 (N_5373,N_4767,N_4528);
nor U5374 (N_5374,N_4646,N_4514);
xor U5375 (N_5375,N_4883,N_4869);
xnor U5376 (N_5376,N_4973,N_4910);
xor U5377 (N_5377,N_4551,N_4804);
xor U5378 (N_5378,N_4735,N_4949);
and U5379 (N_5379,N_4931,N_4544);
xnor U5380 (N_5380,N_4893,N_4695);
or U5381 (N_5381,N_4575,N_4604);
and U5382 (N_5382,N_4999,N_4610);
nand U5383 (N_5383,N_4801,N_4738);
and U5384 (N_5384,N_4574,N_4900);
nor U5385 (N_5385,N_4608,N_4676);
or U5386 (N_5386,N_4809,N_4697);
or U5387 (N_5387,N_4810,N_4777);
nor U5388 (N_5388,N_4710,N_4924);
nor U5389 (N_5389,N_4738,N_4701);
and U5390 (N_5390,N_4939,N_4728);
xnor U5391 (N_5391,N_4531,N_4612);
nand U5392 (N_5392,N_4886,N_4960);
and U5393 (N_5393,N_4885,N_4725);
nor U5394 (N_5394,N_4898,N_4649);
nor U5395 (N_5395,N_4851,N_4804);
or U5396 (N_5396,N_4888,N_4781);
nor U5397 (N_5397,N_4729,N_4985);
and U5398 (N_5398,N_4667,N_4549);
nand U5399 (N_5399,N_4959,N_4818);
nand U5400 (N_5400,N_4776,N_4992);
and U5401 (N_5401,N_4902,N_4850);
and U5402 (N_5402,N_4665,N_4864);
or U5403 (N_5403,N_4700,N_4966);
nor U5404 (N_5404,N_4843,N_4677);
or U5405 (N_5405,N_4726,N_4817);
and U5406 (N_5406,N_4982,N_4633);
and U5407 (N_5407,N_4831,N_4991);
nor U5408 (N_5408,N_4559,N_4856);
nand U5409 (N_5409,N_4968,N_4595);
xor U5410 (N_5410,N_4979,N_4771);
nand U5411 (N_5411,N_4653,N_4717);
nand U5412 (N_5412,N_4652,N_4925);
nor U5413 (N_5413,N_4669,N_4999);
or U5414 (N_5414,N_4525,N_4696);
nand U5415 (N_5415,N_4980,N_4708);
xnor U5416 (N_5416,N_4893,N_4716);
nor U5417 (N_5417,N_4719,N_4723);
xnor U5418 (N_5418,N_4754,N_4788);
nand U5419 (N_5419,N_4952,N_4500);
nand U5420 (N_5420,N_4738,N_4759);
and U5421 (N_5421,N_4650,N_4974);
and U5422 (N_5422,N_4795,N_4528);
and U5423 (N_5423,N_4928,N_4997);
and U5424 (N_5424,N_4631,N_4787);
nand U5425 (N_5425,N_4671,N_4817);
or U5426 (N_5426,N_4707,N_4714);
xnor U5427 (N_5427,N_4827,N_4624);
and U5428 (N_5428,N_4630,N_4571);
nand U5429 (N_5429,N_4961,N_4694);
or U5430 (N_5430,N_4591,N_4942);
or U5431 (N_5431,N_4946,N_4979);
or U5432 (N_5432,N_4654,N_4742);
xnor U5433 (N_5433,N_4873,N_4807);
and U5434 (N_5434,N_4512,N_4831);
or U5435 (N_5435,N_4646,N_4869);
xnor U5436 (N_5436,N_4504,N_4674);
and U5437 (N_5437,N_4522,N_4753);
and U5438 (N_5438,N_4505,N_4926);
and U5439 (N_5439,N_4956,N_4925);
and U5440 (N_5440,N_4947,N_4652);
nor U5441 (N_5441,N_4507,N_4943);
xor U5442 (N_5442,N_4961,N_4518);
nor U5443 (N_5443,N_4543,N_4894);
xor U5444 (N_5444,N_4601,N_4856);
nand U5445 (N_5445,N_4905,N_4520);
xnor U5446 (N_5446,N_4994,N_4739);
or U5447 (N_5447,N_4721,N_4543);
nand U5448 (N_5448,N_4607,N_4546);
xnor U5449 (N_5449,N_4672,N_4530);
or U5450 (N_5450,N_4766,N_4910);
or U5451 (N_5451,N_4762,N_4814);
xor U5452 (N_5452,N_4685,N_4937);
and U5453 (N_5453,N_4523,N_4939);
nor U5454 (N_5454,N_4973,N_4775);
or U5455 (N_5455,N_4869,N_4912);
nand U5456 (N_5456,N_4981,N_4945);
or U5457 (N_5457,N_4953,N_4651);
xnor U5458 (N_5458,N_4743,N_4557);
xnor U5459 (N_5459,N_4971,N_4785);
nand U5460 (N_5460,N_4585,N_4711);
nand U5461 (N_5461,N_4819,N_4606);
nand U5462 (N_5462,N_4990,N_4929);
nand U5463 (N_5463,N_4777,N_4511);
or U5464 (N_5464,N_4585,N_4835);
or U5465 (N_5465,N_4504,N_4511);
xnor U5466 (N_5466,N_4679,N_4717);
or U5467 (N_5467,N_4789,N_4747);
nor U5468 (N_5468,N_4738,N_4910);
nor U5469 (N_5469,N_4756,N_4835);
or U5470 (N_5470,N_4898,N_4967);
or U5471 (N_5471,N_4733,N_4825);
or U5472 (N_5472,N_4949,N_4620);
nand U5473 (N_5473,N_4715,N_4600);
nor U5474 (N_5474,N_4572,N_4940);
xnor U5475 (N_5475,N_4773,N_4977);
nand U5476 (N_5476,N_4670,N_4574);
xnor U5477 (N_5477,N_4688,N_4746);
and U5478 (N_5478,N_4935,N_4833);
xnor U5479 (N_5479,N_4646,N_4904);
nand U5480 (N_5480,N_4687,N_4669);
nor U5481 (N_5481,N_4721,N_4539);
nor U5482 (N_5482,N_4959,N_4621);
nor U5483 (N_5483,N_4820,N_4846);
and U5484 (N_5484,N_4785,N_4746);
xnor U5485 (N_5485,N_4559,N_4688);
or U5486 (N_5486,N_4697,N_4543);
xnor U5487 (N_5487,N_4580,N_4935);
nand U5488 (N_5488,N_4816,N_4945);
or U5489 (N_5489,N_4524,N_4656);
or U5490 (N_5490,N_4933,N_4764);
xor U5491 (N_5491,N_4952,N_4928);
nand U5492 (N_5492,N_4581,N_4621);
xnor U5493 (N_5493,N_4662,N_4782);
nor U5494 (N_5494,N_4949,N_4788);
and U5495 (N_5495,N_4746,N_4630);
nor U5496 (N_5496,N_4776,N_4973);
nand U5497 (N_5497,N_4852,N_4611);
nand U5498 (N_5498,N_4985,N_4845);
xor U5499 (N_5499,N_4550,N_4925);
nand U5500 (N_5500,N_5491,N_5332);
or U5501 (N_5501,N_5150,N_5251);
nor U5502 (N_5502,N_5164,N_5076);
xnor U5503 (N_5503,N_5234,N_5147);
or U5504 (N_5504,N_5123,N_5338);
nor U5505 (N_5505,N_5402,N_5373);
and U5506 (N_5506,N_5378,N_5364);
and U5507 (N_5507,N_5356,N_5268);
and U5508 (N_5508,N_5056,N_5448);
nand U5509 (N_5509,N_5270,N_5028);
or U5510 (N_5510,N_5274,N_5452);
or U5511 (N_5511,N_5118,N_5249);
nand U5512 (N_5512,N_5021,N_5325);
nand U5513 (N_5513,N_5361,N_5167);
xor U5514 (N_5514,N_5066,N_5026);
and U5515 (N_5515,N_5273,N_5357);
or U5516 (N_5516,N_5137,N_5453);
and U5517 (N_5517,N_5319,N_5433);
and U5518 (N_5518,N_5467,N_5132);
xnor U5519 (N_5519,N_5005,N_5475);
xor U5520 (N_5520,N_5352,N_5027);
or U5521 (N_5521,N_5488,N_5033);
and U5522 (N_5522,N_5174,N_5183);
xor U5523 (N_5523,N_5444,N_5406);
xor U5524 (N_5524,N_5483,N_5176);
nand U5525 (N_5525,N_5387,N_5204);
nand U5526 (N_5526,N_5261,N_5257);
or U5527 (N_5527,N_5271,N_5469);
xor U5528 (N_5528,N_5052,N_5473);
and U5529 (N_5529,N_5342,N_5278);
xnor U5530 (N_5530,N_5457,N_5219);
nor U5531 (N_5531,N_5163,N_5161);
xor U5532 (N_5532,N_5039,N_5388);
and U5533 (N_5533,N_5366,N_5272);
and U5534 (N_5534,N_5263,N_5086);
nand U5535 (N_5535,N_5288,N_5030);
or U5536 (N_5536,N_5193,N_5220);
nor U5537 (N_5537,N_5133,N_5470);
nor U5538 (N_5538,N_5210,N_5187);
or U5539 (N_5539,N_5228,N_5354);
and U5540 (N_5540,N_5074,N_5472);
and U5541 (N_5541,N_5148,N_5016);
nand U5542 (N_5542,N_5159,N_5317);
xnor U5543 (N_5543,N_5367,N_5432);
xor U5544 (N_5544,N_5061,N_5313);
nand U5545 (N_5545,N_5018,N_5348);
or U5546 (N_5546,N_5060,N_5478);
nor U5547 (N_5547,N_5434,N_5405);
nor U5548 (N_5548,N_5360,N_5409);
or U5549 (N_5549,N_5421,N_5276);
nand U5550 (N_5550,N_5185,N_5068);
or U5551 (N_5551,N_5291,N_5498);
or U5552 (N_5552,N_5394,N_5374);
xnor U5553 (N_5553,N_5485,N_5145);
xor U5554 (N_5554,N_5011,N_5128);
nand U5555 (N_5555,N_5430,N_5031);
and U5556 (N_5556,N_5098,N_5264);
nand U5557 (N_5557,N_5215,N_5486);
nand U5558 (N_5558,N_5427,N_5200);
xnor U5559 (N_5559,N_5397,N_5194);
and U5560 (N_5560,N_5492,N_5113);
or U5561 (N_5561,N_5152,N_5064);
nand U5562 (N_5562,N_5019,N_5480);
and U5563 (N_5563,N_5139,N_5192);
and U5564 (N_5564,N_5017,N_5496);
xor U5565 (N_5565,N_5410,N_5114);
or U5566 (N_5566,N_5445,N_5247);
nand U5567 (N_5567,N_5260,N_5230);
and U5568 (N_5568,N_5236,N_5283);
nand U5569 (N_5569,N_5300,N_5450);
or U5570 (N_5570,N_5043,N_5059);
nand U5571 (N_5571,N_5262,N_5310);
xor U5572 (N_5572,N_5135,N_5350);
or U5573 (N_5573,N_5381,N_5281);
xnor U5574 (N_5574,N_5315,N_5329);
and U5575 (N_5575,N_5437,N_5004);
nand U5576 (N_5576,N_5438,N_5321);
xnor U5577 (N_5577,N_5070,N_5013);
and U5578 (N_5578,N_5136,N_5180);
xor U5579 (N_5579,N_5385,N_5181);
nor U5580 (N_5580,N_5002,N_5463);
xor U5581 (N_5581,N_5051,N_5223);
nor U5582 (N_5582,N_5391,N_5464);
nand U5583 (N_5583,N_5454,N_5049);
xor U5584 (N_5584,N_5142,N_5412);
and U5585 (N_5585,N_5442,N_5138);
and U5586 (N_5586,N_5490,N_5117);
nor U5587 (N_5587,N_5435,N_5429);
nor U5588 (N_5588,N_5337,N_5462);
and U5589 (N_5589,N_5156,N_5116);
or U5590 (N_5590,N_5399,N_5447);
or U5591 (N_5591,N_5349,N_5363);
nand U5592 (N_5592,N_5379,N_5170);
or U5593 (N_5593,N_5158,N_5034);
and U5594 (N_5594,N_5376,N_5330);
and U5595 (N_5595,N_5422,N_5111);
nor U5596 (N_5596,N_5252,N_5112);
nor U5597 (N_5597,N_5071,N_5221);
or U5598 (N_5598,N_5022,N_5245);
and U5599 (N_5599,N_5400,N_5110);
nor U5600 (N_5600,N_5050,N_5203);
nand U5601 (N_5601,N_5045,N_5372);
xor U5602 (N_5602,N_5331,N_5216);
nor U5603 (N_5603,N_5006,N_5370);
and U5604 (N_5604,N_5202,N_5208);
or U5605 (N_5605,N_5108,N_5091);
nor U5606 (N_5606,N_5308,N_5171);
nand U5607 (N_5607,N_5062,N_5044);
and U5608 (N_5608,N_5380,N_5250);
nand U5609 (N_5609,N_5449,N_5189);
nand U5610 (N_5610,N_5286,N_5067);
nand U5611 (N_5611,N_5355,N_5100);
xor U5612 (N_5612,N_5065,N_5392);
xor U5613 (N_5613,N_5127,N_5382);
nand U5614 (N_5614,N_5347,N_5015);
nor U5615 (N_5615,N_5201,N_5466);
or U5616 (N_5616,N_5009,N_5107);
nand U5617 (N_5617,N_5431,N_5130);
nand U5618 (N_5618,N_5377,N_5369);
xor U5619 (N_5619,N_5484,N_5443);
nor U5620 (N_5620,N_5259,N_5149);
nor U5621 (N_5621,N_5010,N_5477);
xor U5622 (N_5622,N_5063,N_5190);
or U5623 (N_5623,N_5253,N_5175);
and U5624 (N_5624,N_5316,N_5334);
nand U5625 (N_5625,N_5182,N_5154);
nand U5626 (N_5626,N_5155,N_5122);
and U5627 (N_5627,N_5404,N_5080);
nor U5628 (N_5628,N_5087,N_5384);
and U5629 (N_5629,N_5493,N_5375);
nand U5630 (N_5630,N_5206,N_5209);
nand U5631 (N_5631,N_5314,N_5290);
or U5632 (N_5632,N_5456,N_5126);
nor U5633 (N_5633,N_5001,N_5089);
nand U5634 (N_5634,N_5169,N_5481);
and U5635 (N_5635,N_5346,N_5362);
nand U5636 (N_5636,N_5479,N_5295);
and U5637 (N_5637,N_5151,N_5324);
nand U5638 (N_5638,N_5197,N_5320);
nor U5639 (N_5639,N_5237,N_5040);
nor U5640 (N_5640,N_5055,N_5103);
nand U5641 (N_5641,N_5396,N_5307);
nor U5642 (N_5642,N_5416,N_5419);
xor U5643 (N_5643,N_5459,N_5353);
xnor U5644 (N_5644,N_5407,N_5340);
and U5645 (N_5645,N_5032,N_5494);
nand U5646 (N_5646,N_5143,N_5012);
xor U5647 (N_5647,N_5168,N_5077);
nor U5648 (N_5648,N_5205,N_5345);
and U5649 (N_5649,N_5225,N_5440);
nor U5650 (N_5650,N_5301,N_5101);
and U5651 (N_5651,N_5037,N_5081);
and U5652 (N_5652,N_5053,N_5303);
xor U5653 (N_5653,N_5258,N_5153);
nand U5654 (N_5654,N_5038,N_5255);
xor U5655 (N_5655,N_5425,N_5172);
and U5656 (N_5656,N_5157,N_5256);
xnor U5657 (N_5657,N_5458,N_5082);
nor U5658 (N_5658,N_5306,N_5487);
or U5659 (N_5659,N_5390,N_5497);
nor U5660 (N_5660,N_5326,N_5365);
xnor U5661 (N_5661,N_5285,N_5395);
xnor U5662 (N_5662,N_5121,N_5476);
xnor U5663 (N_5663,N_5327,N_5196);
and U5664 (N_5664,N_5025,N_5146);
xor U5665 (N_5665,N_5105,N_5069);
nand U5666 (N_5666,N_5240,N_5224);
and U5667 (N_5667,N_5213,N_5333);
nor U5668 (N_5668,N_5322,N_5265);
xor U5669 (N_5669,N_5489,N_5441);
or U5670 (N_5670,N_5214,N_5403);
or U5671 (N_5671,N_5106,N_5460);
nor U5672 (N_5672,N_5289,N_5041);
nand U5673 (N_5673,N_5227,N_5162);
nor U5674 (N_5674,N_5408,N_5297);
or U5675 (N_5675,N_5014,N_5088);
nor U5676 (N_5676,N_5093,N_5401);
xor U5677 (N_5677,N_5140,N_5424);
or U5678 (N_5678,N_5244,N_5036);
xor U5679 (N_5679,N_5280,N_5092);
nor U5680 (N_5680,N_5057,N_5266);
nor U5681 (N_5681,N_5254,N_5046);
nor U5682 (N_5682,N_5131,N_5226);
nor U5683 (N_5683,N_5109,N_5436);
or U5684 (N_5684,N_5035,N_5495);
and U5685 (N_5685,N_5411,N_5420);
and U5686 (N_5686,N_5465,N_5178);
nor U5687 (N_5687,N_5212,N_5024);
xor U5688 (N_5688,N_5267,N_5241);
nor U5689 (N_5689,N_5296,N_5097);
or U5690 (N_5690,N_5343,N_5023);
xor U5691 (N_5691,N_5000,N_5104);
and U5692 (N_5692,N_5305,N_5231);
xor U5693 (N_5693,N_5222,N_5312);
and U5694 (N_5694,N_5029,N_5358);
and U5695 (N_5695,N_5042,N_5166);
nor U5696 (N_5696,N_5294,N_5047);
and U5697 (N_5697,N_5235,N_5141);
nand U5698 (N_5698,N_5302,N_5423);
or U5699 (N_5699,N_5284,N_5413);
xor U5700 (N_5700,N_5191,N_5482);
and U5701 (N_5701,N_5085,N_5398);
or U5702 (N_5702,N_5008,N_5446);
xor U5703 (N_5703,N_5229,N_5195);
nand U5704 (N_5704,N_5165,N_5177);
or U5705 (N_5705,N_5277,N_5359);
nand U5706 (N_5706,N_5003,N_5218);
xor U5707 (N_5707,N_5339,N_5242);
or U5708 (N_5708,N_5328,N_5248);
nor U5709 (N_5709,N_5318,N_5083);
nand U5710 (N_5710,N_5095,N_5134);
nor U5711 (N_5711,N_5096,N_5094);
xnor U5712 (N_5712,N_5090,N_5102);
or U5713 (N_5713,N_5298,N_5279);
and U5714 (N_5714,N_5471,N_5451);
nor U5715 (N_5715,N_5129,N_5371);
nor U5716 (N_5716,N_5239,N_5120);
or U5717 (N_5717,N_5341,N_5468);
nand U5718 (N_5718,N_5184,N_5426);
and U5719 (N_5719,N_5393,N_5428);
or U5720 (N_5720,N_5383,N_5474);
nand U5721 (N_5721,N_5417,N_5119);
xor U5722 (N_5722,N_5336,N_5054);
or U5723 (N_5723,N_5007,N_5186);
and U5724 (N_5724,N_5188,N_5455);
nand U5725 (N_5725,N_5115,N_5144);
nor U5726 (N_5726,N_5293,N_5073);
xnor U5727 (N_5727,N_5323,N_5269);
or U5728 (N_5728,N_5217,N_5415);
or U5729 (N_5729,N_5292,N_5075);
nand U5730 (N_5730,N_5173,N_5499);
nor U5731 (N_5731,N_5335,N_5389);
or U5732 (N_5732,N_5282,N_5233);
nor U5733 (N_5733,N_5238,N_5079);
nor U5734 (N_5734,N_5386,N_5311);
xor U5735 (N_5735,N_5125,N_5207);
nor U5736 (N_5736,N_5275,N_5304);
nand U5737 (N_5737,N_5246,N_5211);
nor U5738 (N_5738,N_5072,N_5084);
and U5739 (N_5739,N_5351,N_5439);
and U5740 (N_5740,N_5020,N_5368);
nor U5741 (N_5741,N_5299,N_5199);
and U5742 (N_5742,N_5309,N_5344);
nor U5743 (N_5743,N_5160,N_5243);
xnor U5744 (N_5744,N_5414,N_5418);
and U5745 (N_5745,N_5078,N_5179);
or U5746 (N_5746,N_5461,N_5058);
nand U5747 (N_5747,N_5048,N_5232);
xnor U5748 (N_5748,N_5099,N_5287);
nor U5749 (N_5749,N_5198,N_5124);
xor U5750 (N_5750,N_5340,N_5258);
nor U5751 (N_5751,N_5467,N_5078);
nand U5752 (N_5752,N_5233,N_5356);
xnor U5753 (N_5753,N_5359,N_5221);
or U5754 (N_5754,N_5120,N_5013);
nor U5755 (N_5755,N_5342,N_5478);
xor U5756 (N_5756,N_5019,N_5151);
xor U5757 (N_5757,N_5144,N_5378);
xnor U5758 (N_5758,N_5081,N_5248);
and U5759 (N_5759,N_5395,N_5306);
nor U5760 (N_5760,N_5203,N_5478);
or U5761 (N_5761,N_5077,N_5244);
nand U5762 (N_5762,N_5413,N_5391);
and U5763 (N_5763,N_5121,N_5046);
nand U5764 (N_5764,N_5150,N_5038);
xor U5765 (N_5765,N_5255,N_5383);
nand U5766 (N_5766,N_5061,N_5398);
nor U5767 (N_5767,N_5427,N_5381);
or U5768 (N_5768,N_5021,N_5236);
nor U5769 (N_5769,N_5076,N_5032);
xnor U5770 (N_5770,N_5123,N_5149);
and U5771 (N_5771,N_5142,N_5125);
nor U5772 (N_5772,N_5359,N_5405);
nor U5773 (N_5773,N_5042,N_5091);
nand U5774 (N_5774,N_5183,N_5120);
and U5775 (N_5775,N_5280,N_5034);
or U5776 (N_5776,N_5352,N_5183);
nand U5777 (N_5777,N_5009,N_5165);
nand U5778 (N_5778,N_5219,N_5258);
or U5779 (N_5779,N_5301,N_5039);
nand U5780 (N_5780,N_5130,N_5070);
and U5781 (N_5781,N_5075,N_5366);
nor U5782 (N_5782,N_5275,N_5229);
nand U5783 (N_5783,N_5329,N_5092);
or U5784 (N_5784,N_5243,N_5374);
xor U5785 (N_5785,N_5209,N_5475);
xnor U5786 (N_5786,N_5065,N_5368);
xnor U5787 (N_5787,N_5322,N_5394);
nand U5788 (N_5788,N_5442,N_5418);
or U5789 (N_5789,N_5469,N_5049);
and U5790 (N_5790,N_5355,N_5121);
nand U5791 (N_5791,N_5458,N_5427);
nor U5792 (N_5792,N_5035,N_5453);
nand U5793 (N_5793,N_5198,N_5318);
and U5794 (N_5794,N_5326,N_5472);
nand U5795 (N_5795,N_5026,N_5393);
and U5796 (N_5796,N_5052,N_5201);
and U5797 (N_5797,N_5221,N_5191);
xor U5798 (N_5798,N_5128,N_5130);
nor U5799 (N_5799,N_5470,N_5407);
and U5800 (N_5800,N_5448,N_5201);
nand U5801 (N_5801,N_5129,N_5402);
and U5802 (N_5802,N_5281,N_5058);
and U5803 (N_5803,N_5210,N_5469);
xor U5804 (N_5804,N_5143,N_5370);
nand U5805 (N_5805,N_5478,N_5360);
and U5806 (N_5806,N_5290,N_5255);
xor U5807 (N_5807,N_5320,N_5350);
and U5808 (N_5808,N_5063,N_5380);
xnor U5809 (N_5809,N_5436,N_5302);
or U5810 (N_5810,N_5199,N_5443);
xnor U5811 (N_5811,N_5393,N_5100);
or U5812 (N_5812,N_5225,N_5275);
and U5813 (N_5813,N_5267,N_5471);
nor U5814 (N_5814,N_5330,N_5479);
or U5815 (N_5815,N_5411,N_5133);
nor U5816 (N_5816,N_5390,N_5096);
or U5817 (N_5817,N_5068,N_5044);
nor U5818 (N_5818,N_5067,N_5287);
or U5819 (N_5819,N_5199,N_5027);
and U5820 (N_5820,N_5335,N_5381);
or U5821 (N_5821,N_5284,N_5150);
and U5822 (N_5822,N_5380,N_5116);
nand U5823 (N_5823,N_5396,N_5032);
and U5824 (N_5824,N_5099,N_5336);
and U5825 (N_5825,N_5012,N_5047);
and U5826 (N_5826,N_5240,N_5098);
and U5827 (N_5827,N_5474,N_5439);
or U5828 (N_5828,N_5041,N_5131);
nand U5829 (N_5829,N_5017,N_5346);
or U5830 (N_5830,N_5179,N_5095);
or U5831 (N_5831,N_5168,N_5130);
or U5832 (N_5832,N_5103,N_5294);
xor U5833 (N_5833,N_5115,N_5497);
nand U5834 (N_5834,N_5029,N_5166);
nand U5835 (N_5835,N_5362,N_5201);
nor U5836 (N_5836,N_5368,N_5076);
nand U5837 (N_5837,N_5221,N_5449);
or U5838 (N_5838,N_5086,N_5146);
xor U5839 (N_5839,N_5019,N_5010);
and U5840 (N_5840,N_5499,N_5314);
nand U5841 (N_5841,N_5242,N_5310);
or U5842 (N_5842,N_5319,N_5371);
nor U5843 (N_5843,N_5255,N_5206);
and U5844 (N_5844,N_5175,N_5038);
nor U5845 (N_5845,N_5020,N_5386);
xnor U5846 (N_5846,N_5334,N_5163);
nor U5847 (N_5847,N_5295,N_5281);
nand U5848 (N_5848,N_5340,N_5038);
nand U5849 (N_5849,N_5468,N_5252);
xnor U5850 (N_5850,N_5171,N_5081);
xor U5851 (N_5851,N_5272,N_5397);
nand U5852 (N_5852,N_5324,N_5299);
xor U5853 (N_5853,N_5074,N_5419);
xnor U5854 (N_5854,N_5240,N_5172);
nor U5855 (N_5855,N_5004,N_5215);
nand U5856 (N_5856,N_5057,N_5321);
nor U5857 (N_5857,N_5232,N_5289);
or U5858 (N_5858,N_5173,N_5140);
and U5859 (N_5859,N_5013,N_5289);
or U5860 (N_5860,N_5315,N_5296);
and U5861 (N_5861,N_5389,N_5467);
nand U5862 (N_5862,N_5009,N_5437);
xor U5863 (N_5863,N_5018,N_5388);
nand U5864 (N_5864,N_5453,N_5113);
xnor U5865 (N_5865,N_5429,N_5252);
or U5866 (N_5866,N_5093,N_5238);
or U5867 (N_5867,N_5070,N_5253);
nor U5868 (N_5868,N_5029,N_5490);
and U5869 (N_5869,N_5221,N_5274);
or U5870 (N_5870,N_5361,N_5283);
nor U5871 (N_5871,N_5450,N_5151);
nor U5872 (N_5872,N_5488,N_5167);
nor U5873 (N_5873,N_5082,N_5138);
nand U5874 (N_5874,N_5259,N_5355);
nor U5875 (N_5875,N_5499,N_5341);
nor U5876 (N_5876,N_5468,N_5460);
nor U5877 (N_5877,N_5488,N_5335);
xnor U5878 (N_5878,N_5474,N_5132);
xnor U5879 (N_5879,N_5077,N_5267);
and U5880 (N_5880,N_5335,N_5466);
and U5881 (N_5881,N_5074,N_5485);
or U5882 (N_5882,N_5280,N_5362);
nor U5883 (N_5883,N_5203,N_5451);
xnor U5884 (N_5884,N_5007,N_5428);
nor U5885 (N_5885,N_5458,N_5286);
nand U5886 (N_5886,N_5132,N_5113);
or U5887 (N_5887,N_5310,N_5007);
xnor U5888 (N_5888,N_5208,N_5319);
xnor U5889 (N_5889,N_5033,N_5244);
xnor U5890 (N_5890,N_5010,N_5488);
nand U5891 (N_5891,N_5084,N_5402);
or U5892 (N_5892,N_5058,N_5293);
and U5893 (N_5893,N_5426,N_5060);
xnor U5894 (N_5894,N_5247,N_5239);
or U5895 (N_5895,N_5344,N_5117);
and U5896 (N_5896,N_5463,N_5043);
and U5897 (N_5897,N_5245,N_5495);
nand U5898 (N_5898,N_5196,N_5145);
nor U5899 (N_5899,N_5311,N_5364);
nand U5900 (N_5900,N_5293,N_5418);
and U5901 (N_5901,N_5183,N_5324);
nand U5902 (N_5902,N_5404,N_5284);
xor U5903 (N_5903,N_5052,N_5262);
and U5904 (N_5904,N_5016,N_5463);
nand U5905 (N_5905,N_5305,N_5361);
xnor U5906 (N_5906,N_5192,N_5481);
nand U5907 (N_5907,N_5289,N_5012);
or U5908 (N_5908,N_5347,N_5354);
nor U5909 (N_5909,N_5368,N_5063);
and U5910 (N_5910,N_5442,N_5123);
nor U5911 (N_5911,N_5435,N_5366);
nor U5912 (N_5912,N_5222,N_5233);
or U5913 (N_5913,N_5372,N_5249);
or U5914 (N_5914,N_5055,N_5253);
xnor U5915 (N_5915,N_5382,N_5040);
and U5916 (N_5916,N_5190,N_5176);
nor U5917 (N_5917,N_5476,N_5331);
or U5918 (N_5918,N_5285,N_5425);
or U5919 (N_5919,N_5339,N_5215);
nor U5920 (N_5920,N_5492,N_5160);
or U5921 (N_5921,N_5476,N_5434);
xor U5922 (N_5922,N_5245,N_5006);
xnor U5923 (N_5923,N_5164,N_5054);
and U5924 (N_5924,N_5122,N_5294);
and U5925 (N_5925,N_5249,N_5109);
nor U5926 (N_5926,N_5365,N_5492);
nor U5927 (N_5927,N_5242,N_5185);
nor U5928 (N_5928,N_5341,N_5477);
and U5929 (N_5929,N_5010,N_5384);
xnor U5930 (N_5930,N_5224,N_5242);
and U5931 (N_5931,N_5140,N_5383);
and U5932 (N_5932,N_5298,N_5092);
and U5933 (N_5933,N_5102,N_5000);
nor U5934 (N_5934,N_5404,N_5081);
nand U5935 (N_5935,N_5296,N_5025);
xor U5936 (N_5936,N_5252,N_5075);
nand U5937 (N_5937,N_5017,N_5244);
xnor U5938 (N_5938,N_5271,N_5478);
nor U5939 (N_5939,N_5272,N_5104);
xor U5940 (N_5940,N_5317,N_5289);
or U5941 (N_5941,N_5198,N_5300);
or U5942 (N_5942,N_5307,N_5209);
nand U5943 (N_5943,N_5495,N_5322);
nor U5944 (N_5944,N_5401,N_5079);
xnor U5945 (N_5945,N_5318,N_5461);
xnor U5946 (N_5946,N_5199,N_5369);
or U5947 (N_5947,N_5270,N_5259);
or U5948 (N_5948,N_5469,N_5211);
nand U5949 (N_5949,N_5088,N_5481);
nand U5950 (N_5950,N_5124,N_5075);
and U5951 (N_5951,N_5035,N_5339);
xor U5952 (N_5952,N_5442,N_5244);
nor U5953 (N_5953,N_5012,N_5234);
nor U5954 (N_5954,N_5179,N_5279);
xnor U5955 (N_5955,N_5182,N_5214);
nand U5956 (N_5956,N_5040,N_5300);
and U5957 (N_5957,N_5332,N_5363);
nor U5958 (N_5958,N_5032,N_5486);
and U5959 (N_5959,N_5030,N_5172);
and U5960 (N_5960,N_5379,N_5064);
nor U5961 (N_5961,N_5302,N_5238);
and U5962 (N_5962,N_5236,N_5105);
nor U5963 (N_5963,N_5215,N_5181);
nand U5964 (N_5964,N_5050,N_5303);
nand U5965 (N_5965,N_5240,N_5128);
or U5966 (N_5966,N_5071,N_5357);
nor U5967 (N_5967,N_5105,N_5303);
xor U5968 (N_5968,N_5426,N_5355);
nand U5969 (N_5969,N_5218,N_5138);
nand U5970 (N_5970,N_5093,N_5241);
or U5971 (N_5971,N_5444,N_5077);
nand U5972 (N_5972,N_5462,N_5251);
xnor U5973 (N_5973,N_5278,N_5110);
nand U5974 (N_5974,N_5341,N_5157);
nor U5975 (N_5975,N_5137,N_5202);
and U5976 (N_5976,N_5220,N_5163);
or U5977 (N_5977,N_5421,N_5174);
nor U5978 (N_5978,N_5202,N_5256);
and U5979 (N_5979,N_5313,N_5222);
xor U5980 (N_5980,N_5265,N_5070);
and U5981 (N_5981,N_5379,N_5304);
nand U5982 (N_5982,N_5007,N_5437);
nor U5983 (N_5983,N_5010,N_5154);
and U5984 (N_5984,N_5060,N_5045);
or U5985 (N_5985,N_5328,N_5385);
or U5986 (N_5986,N_5275,N_5038);
nor U5987 (N_5987,N_5354,N_5017);
and U5988 (N_5988,N_5494,N_5015);
nand U5989 (N_5989,N_5381,N_5174);
nand U5990 (N_5990,N_5472,N_5005);
xor U5991 (N_5991,N_5288,N_5235);
nor U5992 (N_5992,N_5014,N_5400);
nand U5993 (N_5993,N_5486,N_5392);
or U5994 (N_5994,N_5214,N_5154);
and U5995 (N_5995,N_5052,N_5034);
xnor U5996 (N_5996,N_5343,N_5412);
and U5997 (N_5997,N_5455,N_5172);
or U5998 (N_5998,N_5362,N_5452);
nand U5999 (N_5999,N_5074,N_5160);
xnor U6000 (N_6000,N_5945,N_5565);
or U6001 (N_6001,N_5767,N_5720);
xnor U6002 (N_6002,N_5521,N_5686);
xnor U6003 (N_6003,N_5997,N_5782);
xnor U6004 (N_6004,N_5952,N_5645);
nor U6005 (N_6005,N_5975,N_5799);
and U6006 (N_6006,N_5712,N_5609);
or U6007 (N_6007,N_5885,N_5856);
or U6008 (N_6008,N_5536,N_5841);
nand U6009 (N_6009,N_5919,N_5633);
nor U6010 (N_6010,N_5995,N_5932);
xor U6011 (N_6011,N_5717,N_5817);
or U6012 (N_6012,N_5898,N_5958);
nor U6013 (N_6013,N_5666,N_5830);
nand U6014 (N_6014,N_5665,N_5967);
and U6015 (N_6015,N_5671,N_5766);
nand U6016 (N_6016,N_5639,N_5502);
nand U6017 (N_6017,N_5700,N_5794);
nor U6018 (N_6018,N_5744,N_5790);
nand U6019 (N_6019,N_5556,N_5520);
nand U6020 (N_6020,N_5572,N_5508);
nor U6021 (N_6021,N_5982,N_5742);
and U6022 (N_6022,N_5844,N_5542);
nor U6023 (N_6023,N_5874,N_5883);
xnor U6024 (N_6024,N_5594,N_5903);
nand U6025 (N_6025,N_5581,N_5654);
and U6026 (N_6026,N_5784,N_5636);
or U6027 (N_6027,N_5716,N_5861);
xnor U6028 (N_6028,N_5850,N_5961);
nand U6029 (N_6029,N_5657,N_5760);
and U6030 (N_6030,N_5713,N_5730);
nand U6031 (N_6031,N_5791,N_5714);
and U6032 (N_6032,N_5727,N_5756);
xor U6033 (N_6033,N_5708,N_5899);
nand U6034 (N_6034,N_5795,N_5854);
nand U6035 (N_6035,N_5765,N_5785);
xnor U6036 (N_6036,N_5815,N_5523);
nand U6037 (N_6037,N_5679,N_5925);
or U6038 (N_6038,N_5891,N_5751);
nor U6039 (N_6039,N_5543,N_5605);
and U6040 (N_6040,N_5871,N_5985);
xor U6041 (N_6041,N_5616,N_5801);
nor U6042 (N_6042,N_5753,N_5807);
nor U6043 (N_6043,N_5643,N_5610);
nor U6044 (N_6044,N_5516,N_5827);
and U6045 (N_6045,N_5526,N_5576);
and U6046 (N_6046,N_5804,N_5855);
nand U6047 (N_6047,N_5980,N_5504);
or U6048 (N_6048,N_5549,N_5793);
or U6049 (N_6049,N_5864,N_5906);
xor U6050 (N_6050,N_5986,N_5535);
or U6051 (N_6051,N_5843,N_5518);
or U6052 (N_6052,N_5877,N_5626);
and U6053 (N_6053,N_5950,N_5685);
nor U6054 (N_6054,N_5965,N_5957);
nand U6055 (N_6055,N_5746,N_5563);
nand U6056 (N_6056,N_5923,N_5709);
nor U6057 (N_6057,N_5962,N_5710);
nor U6058 (N_6058,N_5528,N_5603);
xnor U6059 (N_6059,N_5845,N_5599);
or U6060 (N_6060,N_5591,N_5771);
nand U6061 (N_6061,N_5836,N_5889);
xnor U6062 (N_6062,N_5687,N_5737);
nand U6063 (N_6063,N_5509,N_5748);
nor U6064 (N_6064,N_5693,N_5683);
or U6065 (N_6065,N_5822,N_5870);
xor U6066 (N_6066,N_5908,N_5600);
xnor U6067 (N_6067,N_5819,N_5573);
or U6068 (N_6068,N_5773,N_5637);
or U6069 (N_6069,N_5733,N_5918);
xor U6070 (N_6070,N_5992,N_5622);
nand U6071 (N_6071,N_5577,N_5690);
xnor U6072 (N_6072,N_5606,N_5506);
nand U6073 (N_6073,N_5954,N_5640);
nand U6074 (N_6074,N_5951,N_5634);
nand U6075 (N_6075,N_5552,N_5849);
nor U6076 (N_6076,N_5675,N_5983);
and U6077 (N_6077,N_5649,N_5651);
and U6078 (N_6078,N_5688,N_5575);
xnor U6079 (N_6079,N_5655,N_5711);
xnor U6080 (N_6080,N_5812,N_5648);
nor U6081 (N_6081,N_5953,N_5629);
nor U6082 (N_6082,N_5580,N_5989);
nand U6083 (N_6083,N_5544,N_5803);
and U6084 (N_6084,N_5724,N_5956);
xnor U6085 (N_6085,N_5917,N_5792);
or U6086 (N_6086,N_5761,N_5545);
nor U6087 (N_6087,N_5707,N_5993);
or U6088 (N_6088,N_5647,N_5949);
and U6089 (N_6089,N_5628,N_5659);
and U6090 (N_6090,N_5860,N_5635);
and U6091 (N_6091,N_5660,N_5532);
or U6092 (N_6092,N_5842,N_5978);
nor U6093 (N_6093,N_5846,N_5886);
or U6094 (N_6094,N_5814,N_5926);
or U6095 (N_6095,N_5630,N_5513);
or U6096 (N_6096,N_5974,N_5517);
or U6097 (N_6097,N_5596,N_5991);
nor U6098 (N_6098,N_5534,N_5680);
nand U6099 (N_6099,N_5798,N_5823);
xor U6100 (N_6100,N_5668,N_5676);
xnor U6101 (N_6101,N_5947,N_5988);
xor U6102 (N_6102,N_5584,N_5821);
and U6103 (N_6103,N_5538,N_5762);
xor U6104 (N_6104,N_5681,N_5620);
and U6105 (N_6105,N_5863,N_5833);
or U6106 (N_6106,N_5546,N_5718);
xor U6107 (N_6107,N_5808,N_5706);
nand U6108 (N_6108,N_5539,N_5745);
nor U6109 (N_6109,N_5562,N_5853);
and U6110 (N_6110,N_5946,N_5701);
nand U6111 (N_6111,N_5857,N_5557);
or U6112 (N_6112,N_5829,N_5677);
nand U6113 (N_6113,N_5922,N_5530);
nor U6114 (N_6114,N_5578,N_5757);
or U6115 (N_6115,N_5514,N_5615);
nand U6116 (N_6116,N_5831,N_5752);
xor U6117 (N_6117,N_5696,N_5939);
xor U6118 (N_6118,N_5840,N_5990);
and U6119 (N_6119,N_5558,N_5656);
or U6120 (N_6120,N_5501,N_5809);
and U6121 (N_6121,N_5694,N_5914);
and U6122 (N_6122,N_5892,N_5927);
and U6123 (N_6123,N_5828,N_5884);
or U6124 (N_6124,N_5780,N_5510);
xor U6125 (N_6125,N_5881,N_5595);
nand U6126 (N_6126,N_5623,N_5554);
or U6127 (N_6127,N_5979,N_5598);
or U6128 (N_6128,N_5678,N_5547);
and U6129 (N_6129,N_5879,N_5692);
xor U6130 (N_6130,N_5631,N_5862);
nand U6131 (N_6131,N_5811,N_5503);
or U6132 (N_6132,N_5943,N_5505);
nor U6133 (N_6133,N_5944,N_5875);
and U6134 (N_6134,N_5847,N_5796);
or U6135 (N_6135,N_5704,N_5587);
xnor U6136 (N_6136,N_5570,N_5825);
or U6137 (N_6137,N_5641,N_5848);
or U6138 (N_6138,N_5537,N_5936);
and U6139 (N_6139,N_5867,N_5749);
or U6140 (N_6140,N_5909,N_5592);
nand U6141 (N_6141,N_5673,N_5941);
nand U6142 (N_6142,N_5826,N_5916);
nor U6143 (N_6143,N_5601,N_5566);
nor U6144 (N_6144,N_5691,N_5619);
or U6145 (N_6145,N_5934,N_5866);
and U6146 (N_6146,N_5583,N_5878);
nor U6147 (N_6147,N_5969,N_5736);
xor U6148 (N_6148,N_5618,N_5984);
nand U6149 (N_6149,N_5973,N_5627);
nand U6150 (N_6150,N_5533,N_5873);
or U6151 (N_6151,N_5933,N_5588);
xnor U6152 (N_6152,N_5728,N_5894);
nor U6153 (N_6153,N_5662,N_5882);
or U6154 (N_6154,N_5838,N_5887);
nand U6155 (N_6155,N_5888,N_5865);
and U6156 (N_6156,N_5729,N_5590);
nand U6157 (N_6157,N_5859,N_5548);
xnor U6158 (N_6158,N_5999,N_5998);
nand U6159 (N_6159,N_5772,N_5820);
nand U6160 (N_6160,N_5515,N_5650);
nor U6161 (N_6161,N_5579,N_5977);
or U6162 (N_6162,N_5699,N_5754);
nand U6163 (N_6163,N_5652,N_5779);
or U6164 (N_6164,N_5868,N_5904);
and U6165 (N_6165,N_5813,N_5834);
and U6166 (N_6166,N_5763,N_5586);
nor U6167 (N_6167,N_5698,N_5511);
nand U6168 (N_6168,N_5930,N_5674);
or U6169 (N_6169,N_5597,N_5697);
nor U6170 (N_6170,N_5540,N_5938);
or U6171 (N_6171,N_5638,N_5802);
nand U6172 (N_6172,N_5722,N_5670);
and U6173 (N_6173,N_5604,N_5672);
nand U6174 (N_6174,N_5781,N_5667);
and U6175 (N_6175,N_5658,N_5527);
nor U6176 (N_6176,N_5937,N_5805);
and U6177 (N_6177,N_5774,N_5755);
nor U6178 (N_6178,N_5955,N_5703);
nand U6179 (N_6179,N_5776,N_5964);
or U6180 (N_6180,N_5726,N_5902);
nor U6181 (N_6181,N_5912,N_5719);
and U6182 (N_6182,N_5920,N_5858);
nor U6183 (N_6183,N_5738,N_5872);
or U6184 (N_6184,N_5607,N_5741);
xnor U6185 (N_6185,N_5996,N_5702);
nor U6186 (N_6186,N_5966,N_5602);
nand U6187 (N_6187,N_5735,N_5915);
xor U6188 (N_6188,N_5759,N_5743);
xor U6189 (N_6189,N_5960,N_5560);
nor U6190 (N_6190,N_5948,N_5806);
nor U6191 (N_6191,N_5529,N_5624);
nand U6192 (N_6192,N_5901,N_5642);
nand U6193 (N_6193,N_5531,N_5893);
nor U6194 (N_6194,N_5569,N_5739);
xnor U6195 (N_6195,N_5561,N_5775);
or U6196 (N_6196,N_5810,N_5608);
or U6197 (N_6197,N_5876,N_5769);
and U6198 (N_6198,N_5942,N_5921);
or U6199 (N_6199,N_5574,N_5896);
nor U6200 (N_6200,N_5907,N_5725);
and U6201 (N_6201,N_5895,N_5800);
xor U6202 (N_6202,N_5664,N_5585);
xor U6203 (N_6203,N_5525,N_5797);
nor U6204 (N_6204,N_5614,N_5522);
and U6205 (N_6205,N_5928,N_5768);
or U6206 (N_6206,N_5661,N_5519);
nor U6207 (N_6207,N_5935,N_5669);
xnor U6208 (N_6208,N_5963,N_5839);
xnor U6209 (N_6209,N_5787,N_5571);
nand U6210 (N_6210,N_5970,N_5541);
xnor U6211 (N_6211,N_5589,N_5621);
xor U6212 (N_6212,N_5976,N_5551);
nor U6213 (N_6213,N_5750,N_5911);
or U6214 (N_6214,N_5617,N_5732);
and U6215 (N_6215,N_5632,N_5924);
or U6216 (N_6216,N_5555,N_5852);
and U6217 (N_6217,N_5758,N_5880);
and U6218 (N_6218,N_5777,N_5715);
and U6219 (N_6219,N_5788,N_5684);
and U6220 (N_6220,N_5987,N_5613);
nor U6221 (N_6221,N_5981,N_5851);
or U6222 (N_6222,N_5900,N_5559);
and U6223 (N_6223,N_5567,N_5783);
xor U6224 (N_6224,N_5764,N_5835);
xor U6225 (N_6225,N_5971,N_5905);
nor U6226 (N_6226,N_5524,N_5500);
nand U6227 (N_6227,N_5816,N_5913);
xnor U6228 (N_6228,N_5695,N_5972);
or U6229 (N_6229,N_5689,N_5731);
and U6230 (N_6230,N_5890,N_5734);
xor U6231 (N_6231,N_5837,N_5994);
nand U6232 (N_6232,N_5705,N_5832);
nand U6233 (N_6233,N_5747,N_5740);
and U6234 (N_6234,N_5778,N_5568);
nand U6235 (N_6235,N_5507,N_5770);
or U6236 (N_6236,N_5897,N_5582);
nand U6237 (N_6237,N_5959,N_5653);
nand U6238 (N_6238,N_5786,N_5723);
nor U6239 (N_6239,N_5910,N_5931);
xnor U6240 (N_6240,N_5553,N_5663);
nor U6241 (N_6241,N_5940,N_5512);
nor U6242 (N_6242,N_5682,N_5968);
nand U6243 (N_6243,N_5564,N_5869);
or U6244 (N_6244,N_5721,N_5824);
or U6245 (N_6245,N_5818,N_5646);
nor U6246 (N_6246,N_5593,N_5625);
nor U6247 (N_6247,N_5789,N_5550);
nor U6248 (N_6248,N_5612,N_5611);
and U6249 (N_6249,N_5644,N_5929);
nand U6250 (N_6250,N_5779,N_5694);
and U6251 (N_6251,N_5869,N_5680);
or U6252 (N_6252,N_5660,N_5596);
nor U6253 (N_6253,N_5903,N_5784);
nor U6254 (N_6254,N_5733,N_5674);
or U6255 (N_6255,N_5716,N_5652);
nand U6256 (N_6256,N_5793,N_5559);
and U6257 (N_6257,N_5707,N_5756);
xnor U6258 (N_6258,N_5839,N_5968);
and U6259 (N_6259,N_5547,N_5541);
nand U6260 (N_6260,N_5711,N_5696);
and U6261 (N_6261,N_5732,N_5833);
nand U6262 (N_6262,N_5715,N_5932);
nand U6263 (N_6263,N_5638,N_5590);
nand U6264 (N_6264,N_5610,N_5714);
nand U6265 (N_6265,N_5744,N_5942);
nand U6266 (N_6266,N_5933,N_5776);
nand U6267 (N_6267,N_5959,N_5822);
and U6268 (N_6268,N_5700,N_5660);
xor U6269 (N_6269,N_5711,N_5927);
nand U6270 (N_6270,N_5772,N_5514);
and U6271 (N_6271,N_5583,N_5713);
and U6272 (N_6272,N_5973,N_5654);
xnor U6273 (N_6273,N_5825,N_5526);
and U6274 (N_6274,N_5842,N_5951);
or U6275 (N_6275,N_5856,N_5858);
nor U6276 (N_6276,N_5617,N_5733);
and U6277 (N_6277,N_5528,N_5723);
and U6278 (N_6278,N_5784,N_5941);
nor U6279 (N_6279,N_5610,N_5873);
or U6280 (N_6280,N_5627,N_5995);
xor U6281 (N_6281,N_5718,N_5781);
nor U6282 (N_6282,N_5587,N_5861);
xor U6283 (N_6283,N_5593,N_5707);
and U6284 (N_6284,N_5819,N_5995);
xor U6285 (N_6285,N_5594,N_5731);
nand U6286 (N_6286,N_5942,N_5630);
and U6287 (N_6287,N_5564,N_5539);
xor U6288 (N_6288,N_5695,N_5630);
xor U6289 (N_6289,N_5974,N_5550);
nand U6290 (N_6290,N_5629,N_5526);
nand U6291 (N_6291,N_5980,N_5683);
xor U6292 (N_6292,N_5826,N_5863);
xnor U6293 (N_6293,N_5893,N_5639);
nor U6294 (N_6294,N_5866,N_5718);
xnor U6295 (N_6295,N_5608,N_5790);
or U6296 (N_6296,N_5610,N_5552);
xor U6297 (N_6297,N_5972,N_5992);
or U6298 (N_6298,N_5620,N_5582);
xnor U6299 (N_6299,N_5528,N_5686);
and U6300 (N_6300,N_5590,N_5545);
nand U6301 (N_6301,N_5726,N_5827);
nor U6302 (N_6302,N_5929,N_5835);
xnor U6303 (N_6303,N_5785,N_5547);
or U6304 (N_6304,N_5677,N_5595);
and U6305 (N_6305,N_5762,N_5846);
and U6306 (N_6306,N_5527,N_5569);
or U6307 (N_6307,N_5563,N_5555);
or U6308 (N_6308,N_5591,N_5986);
or U6309 (N_6309,N_5856,N_5757);
nand U6310 (N_6310,N_5787,N_5990);
xnor U6311 (N_6311,N_5770,N_5906);
or U6312 (N_6312,N_5700,N_5758);
and U6313 (N_6313,N_5746,N_5548);
nand U6314 (N_6314,N_5841,N_5788);
xnor U6315 (N_6315,N_5788,N_5877);
nand U6316 (N_6316,N_5516,N_5758);
and U6317 (N_6317,N_5913,N_5610);
nand U6318 (N_6318,N_5819,N_5714);
and U6319 (N_6319,N_5929,N_5575);
nand U6320 (N_6320,N_5890,N_5717);
nor U6321 (N_6321,N_5898,N_5815);
nor U6322 (N_6322,N_5751,N_5697);
nor U6323 (N_6323,N_5998,N_5623);
nor U6324 (N_6324,N_5573,N_5914);
or U6325 (N_6325,N_5550,N_5902);
or U6326 (N_6326,N_5759,N_5958);
nand U6327 (N_6327,N_5690,N_5736);
or U6328 (N_6328,N_5696,N_5858);
or U6329 (N_6329,N_5579,N_5576);
and U6330 (N_6330,N_5736,N_5813);
nor U6331 (N_6331,N_5963,N_5696);
nor U6332 (N_6332,N_5769,N_5804);
or U6333 (N_6333,N_5751,N_5668);
xnor U6334 (N_6334,N_5798,N_5882);
nor U6335 (N_6335,N_5558,N_5853);
nand U6336 (N_6336,N_5829,N_5970);
nand U6337 (N_6337,N_5603,N_5561);
xor U6338 (N_6338,N_5928,N_5765);
or U6339 (N_6339,N_5820,N_5654);
nor U6340 (N_6340,N_5686,N_5911);
nand U6341 (N_6341,N_5902,N_5756);
xnor U6342 (N_6342,N_5670,N_5682);
nand U6343 (N_6343,N_5548,N_5519);
xnor U6344 (N_6344,N_5750,N_5940);
nor U6345 (N_6345,N_5807,N_5824);
nor U6346 (N_6346,N_5804,N_5789);
or U6347 (N_6347,N_5926,N_5623);
xor U6348 (N_6348,N_5770,N_5543);
nor U6349 (N_6349,N_5807,N_5927);
and U6350 (N_6350,N_5707,N_5831);
or U6351 (N_6351,N_5691,N_5596);
or U6352 (N_6352,N_5611,N_5617);
xor U6353 (N_6353,N_5975,N_5813);
xnor U6354 (N_6354,N_5882,N_5983);
nor U6355 (N_6355,N_5938,N_5884);
nand U6356 (N_6356,N_5566,N_5563);
xnor U6357 (N_6357,N_5901,N_5798);
nor U6358 (N_6358,N_5745,N_5597);
and U6359 (N_6359,N_5528,N_5501);
nor U6360 (N_6360,N_5582,N_5906);
and U6361 (N_6361,N_5984,N_5743);
nor U6362 (N_6362,N_5907,N_5889);
or U6363 (N_6363,N_5514,N_5905);
or U6364 (N_6364,N_5509,N_5691);
and U6365 (N_6365,N_5881,N_5593);
nand U6366 (N_6366,N_5663,N_5841);
nand U6367 (N_6367,N_5974,N_5863);
nor U6368 (N_6368,N_5601,N_5726);
xor U6369 (N_6369,N_5680,N_5808);
or U6370 (N_6370,N_5783,N_5888);
and U6371 (N_6371,N_5718,N_5966);
nor U6372 (N_6372,N_5945,N_5716);
or U6373 (N_6373,N_5524,N_5836);
xnor U6374 (N_6374,N_5882,N_5936);
nor U6375 (N_6375,N_5826,N_5688);
xnor U6376 (N_6376,N_5743,N_5993);
nand U6377 (N_6377,N_5722,N_5972);
and U6378 (N_6378,N_5974,N_5973);
xnor U6379 (N_6379,N_5902,N_5970);
nor U6380 (N_6380,N_5960,N_5781);
nor U6381 (N_6381,N_5523,N_5936);
and U6382 (N_6382,N_5721,N_5804);
nor U6383 (N_6383,N_5882,N_5667);
and U6384 (N_6384,N_5980,N_5661);
or U6385 (N_6385,N_5534,N_5923);
nand U6386 (N_6386,N_5689,N_5666);
nor U6387 (N_6387,N_5956,N_5639);
xnor U6388 (N_6388,N_5600,N_5944);
nand U6389 (N_6389,N_5542,N_5974);
and U6390 (N_6390,N_5556,N_5595);
nor U6391 (N_6391,N_5750,N_5989);
nand U6392 (N_6392,N_5970,N_5721);
nand U6393 (N_6393,N_5976,N_5913);
nor U6394 (N_6394,N_5563,N_5934);
and U6395 (N_6395,N_5657,N_5838);
nand U6396 (N_6396,N_5649,N_5851);
nor U6397 (N_6397,N_5584,N_5532);
nor U6398 (N_6398,N_5514,N_5957);
and U6399 (N_6399,N_5780,N_5666);
nand U6400 (N_6400,N_5588,N_5649);
and U6401 (N_6401,N_5606,N_5955);
nand U6402 (N_6402,N_5705,N_5923);
nor U6403 (N_6403,N_5705,N_5911);
nand U6404 (N_6404,N_5771,N_5904);
nand U6405 (N_6405,N_5564,N_5559);
nand U6406 (N_6406,N_5989,N_5861);
nand U6407 (N_6407,N_5798,N_5749);
nor U6408 (N_6408,N_5537,N_5891);
nor U6409 (N_6409,N_5810,N_5987);
nor U6410 (N_6410,N_5513,N_5720);
and U6411 (N_6411,N_5670,N_5950);
or U6412 (N_6412,N_5832,N_5548);
and U6413 (N_6413,N_5885,N_5561);
xor U6414 (N_6414,N_5575,N_5504);
nor U6415 (N_6415,N_5603,N_5719);
nand U6416 (N_6416,N_5921,N_5959);
and U6417 (N_6417,N_5789,N_5873);
nor U6418 (N_6418,N_5554,N_5889);
or U6419 (N_6419,N_5967,N_5991);
nor U6420 (N_6420,N_5803,N_5843);
xnor U6421 (N_6421,N_5594,N_5825);
nand U6422 (N_6422,N_5677,N_5603);
nand U6423 (N_6423,N_5923,N_5522);
xor U6424 (N_6424,N_5775,N_5515);
and U6425 (N_6425,N_5612,N_5729);
and U6426 (N_6426,N_5555,N_5614);
nor U6427 (N_6427,N_5542,N_5842);
xnor U6428 (N_6428,N_5745,N_5791);
nor U6429 (N_6429,N_5516,N_5544);
nand U6430 (N_6430,N_5960,N_5626);
or U6431 (N_6431,N_5783,N_5958);
nand U6432 (N_6432,N_5641,N_5885);
nor U6433 (N_6433,N_5835,N_5860);
or U6434 (N_6434,N_5532,N_5788);
and U6435 (N_6435,N_5723,N_5623);
xnor U6436 (N_6436,N_5888,N_5794);
nand U6437 (N_6437,N_5653,N_5870);
xnor U6438 (N_6438,N_5533,N_5557);
or U6439 (N_6439,N_5547,N_5602);
nor U6440 (N_6440,N_5692,N_5683);
nand U6441 (N_6441,N_5523,N_5566);
xnor U6442 (N_6442,N_5638,N_5787);
nor U6443 (N_6443,N_5611,N_5758);
and U6444 (N_6444,N_5651,N_5687);
nand U6445 (N_6445,N_5658,N_5734);
xor U6446 (N_6446,N_5932,N_5865);
and U6447 (N_6447,N_5892,N_5647);
or U6448 (N_6448,N_5992,N_5848);
nor U6449 (N_6449,N_5949,N_5627);
xnor U6450 (N_6450,N_5944,N_5951);
nand U6451 (N_6451,N_5755,N_5627);
or U6452 (N_6452,N_5890,N_5590);
and U6453 (N_6453,N_5514,N_5641);
nand U6454 (N_6454,N_5529,N_5822);
xnor U6455 (N_6455,N_5811,N_5975);
or U6456 (N_6456,N_5715,N_5595);
xor U6457 (N_6457,N_5964,N_5516);
and U6458 (N_6458,N_5970,N_5618);
xor U6459 (N_6459,N_5559,N_5872);
or U6460 (N_6460,N_5741,N_5654);
nor U6461 (N_6461,N_5822,N_5979);
xor U6462 (N_6462,N_5688,N_5613);
nor U6463 (N_6463,N_5756,N_5571);
nand U6464 (N_6464,N_5858,N_5907);
xnor U6465 (N_6465,N_5848,N_5594);
or U6466 (N_6466,N_5634,N_5899);
and U6467 (N_6467,N_5718,N_5694);
xor U6468 (N_6468,N_5655,N_5602);
nand U6469 (N_6469,N_5560,N_5794);
or U6470 (N_6470,N_5553,N_5924);
and U6471 (N_6471,N_5651,N_5520);
nor U6472 (N_6472,N_5718,N_5712);
and U6473 (N_6473,N_5994,N_5764);
and U6474 (N_6474,N_5628,N_5566);
nor U6475 (N_6475,N_5922,N_5643);
or U6476 (N_6476,N_5891,N_5767);
xnor U6477 (N_6477,N_5505,N_5610);
xor U6478 (N_6478,N_5808,N_5695);
xor U6479 (N_6479,N_5701,N_5961);
nand U6480 (N_6480,N_5646,N_5957);
and U6481 (N_6481,N_5866,N_5568);
and U6482 (N_6482,N_5976,N_5792);
or U6483 (N_6483,N_5647,N_5727);
or U6484 (N_6484,N_5699,N_5653);
or U6485 (N_6485,N_5900,N_5862);
xnor U6486 (N_6486,N_5591,N_5874);
nand U6487 (N_6487,N_5747,N_5512);
nor U6488 (N_6488,N_5722,N_5699);
and U6489 (N_6489,N_5813,N_5752);
nand U6490 (N_6490,N_5968,N_5551);
xor U6491 (N_6491,N_5937,N_5771);
xnor U6492 (N_6492,N_5602,N_5579);
xor U6493 (N_6493,N_5777,N_5861);
nand U6494 (N_6494,N_5741,N_5542);
nor U6495 (N_6495,N_5624,N_5761);
xor U6496 (N_6496,N_5996,N_5660);
xor U6497 (N_6497,N_5609,N_5658);
and U6498 (N_6498,N_5517,N_5607);
nand U6499 (N_6499,N_5521,N_5630);
xor U6500 (N_6500,N_6248,N_6074);
nor U6501 (N_6501,N_6049,N_6139);
xor U6502 (N_6502,N_6052,N_6107);
nand U6503 (N_6503,N_6276,N_6326);
nor U6504 (N_6504,N_6318,N_6163);
nand U6505 (N_6505,N_6366,N_6250);
and U6506 (N_6506,N_6388,N_6443);
or U6507 (N_6507,N_6297,N_6089);
or U6508 (N_6508,N_6496,N_6474);
nor U6509 (N_6509,N_6026,N_6394);
and U6510 (N_6510,N_6216,N_6386);
xor U6511 (N_6511,N_6482,N_6345);
xor U6512 (N_6512,N_6333,N_6375);
xnor U6513 (N_6513,N_6030,N_6174);
xor U6514 (N_6514,N_6494,N_6420);
nand U6515 (N_6515,N_6153,N_6398);
nand U6516 (N_6516,N_6266,N_6493);
and U6517 (N_6517,N_6035,N_6477);
xnor U6518 (N_6518,N_6077,N_6313);
xnor U6519 (N_6519,N_6237,N_6417);
nand U6520 (N_6520,N_6063,N_6135);
nor U6521 (N_6521,N_6230,N_6426);
nand U6522 (N_6522,N_6060,N_6304);
nand U6523 (N_6523,N_6179,N_6003);
xor U6524 (N_6524,N_6222,N_6041);
or U6525 (N_6525,N_6399,N_6019);
nor U6526 (N_6526,N_6460,N_6108);
and U6527 (N_6527,N_6207,N_6235);
xnor U6528 (N_6528,N_6117,N_6098);
and U6529 (N_6529,N_6129,N_6432);
and U6530 (N_6530,N_6181,N_6412);
nor U6531 (N_6531,N_6111,N_6009);
nand U6532 (N_6532,N_6152,N_6343);
nor U6533 (N_6533,N_6485,N_6404);
xor U6534 (N_6534,N_6469,N_6346);
nor U6535 (N_6535,N_6047,N_6127);
and U6536 (N_6536,N_6415,N_6273);
and U6537 (N_6537,N_6268,N_6224);
or U6538 (N_6538,N_6253,N_6450);
nor U6539 (N_6539,N_6194,N_6040);
nor U6540 (N_6540,N_6295,N_6467);
xor U6541 (N_6541,N_6440,N_6002);
xor U6542 (N_6542,N_6146,N_6159);
or U6543 (N_6543,N_6080,N_6396);
xnor U6544 (N_6544,N_6294,N_6160);
and U6545 (N_6545,N_6354,N_6185);
and U6546 (N_6546,N_6016,N_6322);
nand U6547 (N_6547,N_6122,N_6116);
nor U6548 (N_6548,N_6358,N_6286);
or U6549 (N_6549,N_6186,N_6355);
or U6550 (N_6550,N_6189,N_6184);
or U6551 (N_6551,N_6498,N_6314);
nor U6552 (N_6552,N_6448,N_6403);
and U6553 (N_6553,N_6282,N_6411);
nand U6554 (N_6554,N_6164,N_6406);
and U6555 (N_6555,N_6374,N_6102);
or U6556 (N_6556,N_6243,N_6246);
nand U6557 (N_6557,N_6439,N_6090);
nor U6558 (N_6558,N_6013,N_6337);
xnor U6559 (N_6559,N_6114,N_6381);
nor U6560 (N_6560,N_6023,N_6199);
xnor U6561 (N_6561,N_6180,N_6109);
nand U6562 (N_6562,N_6240,N_6259);
and U6563 (N_6563,N_6262,N_6414);
nand U6564 (N_6564,N_6293,N_6087);
and U6565 (N_6565,N_6225,N_6138);
nand U6566 (N_6566,N_6034,N_6303);
nor U6567 (N_6567,N_6195,N_6461);
or U6568 (N_6568,N_6490,N_6390);
and U6569 (N_6569,N_6154,N_6369);
nor U6570 (N_6570,N_6351,N_6055);
nand U6571 (N_6571,N_6226,N_6488);
nor U6572 (N_6572,N_6210,N_6070);
nand U6573 (N_6573,N_6072,N_6271);
nor U6574 (N_6574,N_6310,N_6064);
or U6575 (N_6575,N_6312,N_6274);
nor U6576 (N_6576,N_6134,N_6384);
nor U6577 (N_6577,N_6359,N_6280);
nand U6578 (N_6578,N_6104,N_6368);
nand U6579 (N_6579,N_6076,N_6370);
nand U6580 (N_6580,N_6133,N_6046);
and U6581 (N_6581,N_6042,N_6444);
and U6582 (N_6582,N_6340,N_6245);
nand U6583 (N_6583,N_6212,N_6086);
nand U6584 (N_6584,N_6476,N_6085);
and U6585 (N_6585,N_6486,N_6130);
nor U6586 (N_6586,N_6220,N_6344);
or U6587 (N_6587,N_6317,N_6115);
or U6588 (N_6588,N_6376,N_6125);
nand U6589 (N_6589,N_6020,N_6015);
nand U6590 (N_6590,N_6054,N_6097);
or U6591 (N_6591,N_6385,N_6056);
xnor U6592 (N_6592,N_6204,N_6321);
nand U6593 (N_6593,N_6362,N_6455);
nand U6594 (N_6594,N_6434,N_6397);
nand U6595 (N_6595,N_6140,N_6029);
nor U6596 (N_6596,N_6238,N_6454);
nor U6597 (N_6597,N_6437,N_6472);
nor U6598 (N_6598,N_6027,N_6378);
or U6599 (N_6599,N_6119,N_6158);
and U6600 (N_6600,N_6331,N_6229);
xor U6601 (N_6601,N_6353,N_6236);
nand U6602 (N_6602,N_6277,N_6335);
nor U6603 (N_6603,N_6323,N_6169);
nor U6604 (N_6604,N_6031,N_6330);
or U6605 (N_6605,N_6305,N_6005);
xor U6606 (N_6606,N_6188,N_6018);
and U6607 (N_6607,N_6038,N_6401);
and U6608 (N_6608,N_6288,N_6065);
or U6609 (N_6609,N_6463,N_6315);
xnor U6610 (N_6610,N_6424,N_6449);
xnor U6611 (N_6611,N_6413,N_6291);
xor U6612 (N_6612,N_6156,N_6043);
nand U6613 (N_6613,N_6400,N_6078);
xor U6614 (N_6614,N_6148,N_6082);
or U6615 (N_6615,N_6149,N_6252);
xor U6616 (N_6616,N_6126,N_6352);
nand U6617 (N_6617,N_6497,N_6100);
and U6618 (N_6618,N_6380,N_6083);
nand U6619 (N_6619,N_6059,N_6275);
and U6620 (N_6620,N_6242,N_6022);
nor U6621 (N_6621,N_6234,N_6492);
nor U6622 (N_6622,N_6228,N_6348);
nand U6623 (N_6623,N_6192,N_6435);
and U6624 (N_6624,N_6124,N_6197);
nor U6625 (N_6625,N_6096,N_6190);
and U6626 (N_6626,N_6187,N_6499);
nor U6627 (N_6627,N_6025,N_6350);
and U6628 (N_6628,N_6165,N_6254);
nand U6629 (N_6629,N_6155,N_6427);
nor U6630 (N_6630,N_6172,N_6360);
nand U6631 (N_6631,N_6132,N_6017);
xnor U6632 (N_6632,N_6162,N_6361);
xnor U6633 (N_6633,N_6298,N_6006);
and U6634 (N_6634,N_6357,N_6445);
nand U6635 (N_6635,N_6283,N_6302);
or U6636 (N_6636,N_6141,N_6481);
or U6637 (N_6637,N_6211,N_6033);
and U6638 (N_6638,N_6290,N_6021);
nor U6639 (N_6639,N_6084,N_6215);
xor U6640 (N_6640,N_6451,N_6379);
nor U6641 (N_6641,N_6136,N_6144);
nand U6642 (N_6642,N_6438,N_6145);
nor U6643 (N_6643,N_6247,N_6419);
nand U6644 (N_6644,N_6372,N_6051);
or U6645 (N_6645,N_6405,N_6170);
xnor U6646 (N_6646,N_6422,N_6263);
nand U6647 (N_6647,N_6442,N_6329);
or U6648 (N_6648,N_6284,N_6270);
or U6649 (N_6649,N_6347,N_6267);
nand U6650 (N_6650,N_6073,N_6382);
nor U6651 (N_6651,N_6342,N_6014);
xor U6652 (N_6652,N_6191,N_6068);
nor U6653 (N_6653,N_6383,N_6478);
nand U6654 (N_6654,N_6101,N_6465);
and U6655 (N_6655,N_6150,N_6428);
and U6656 (N_6656,N_6209,N_6311);
xnor U6657 (N_6657,N_6121,N_6168);
and U6658 (N_6658,N_6334,N_6473);
xor U6659 (N_6659,N_6110,N_6183);
xnor U6660 (N_6660,N_6300,N_6470);
nand U6661 (N_6661,N_6393,N_6495);
nor U6662 (N_6662,N_6447,N_6408);
nand U6663 (N_6663,N_6429,N_6249);
and U6664 (N_6664,N_6423,N_6410);
and U6665 (N_6665,N_6039,N_6241);
nand U6666 (N_6666,N_6371,N_6193);
nor U6667 (N_6667,N_6281,N_6251);
or U6668 (N_6668,N_6028,N_6024);
and U6669 (N_6669,N_6299,N_6256);
and U6670 (N_6670,N_6258,N_6218);
or U6671 (N_6671,N_6475,N_6196);
and U6672 (N_6672,N_6239,N_6319);
xor U6673 (N_6673,N_6128,N_6269);
nand U6674 (N_6674,N_6264,N_6279);
xor U6675 (N_6675,N_6480,N_6157);
nand U6676 (N_6676,N_6200,N_6198);
nand U6677 (N_6677,N_6123,N_6356);
or U6678 (N_6678,N_6471,N_6112);
and U6679 (N_6679,N_6221,N_6453);
nand U6680 (N_6680,N_6227,N_6095);
or U6681 (N_6681,N_6484,N_6306);
nand U6682 (N_6682,N_6285,N_6171);
or U6683 (N_6683,N_6456,N_6327);
nand U6684 (N_6684,N_6464,N_6416);
xnor U6685 (N_6685,N_6147,N_6071);
nand U6686 (N_6686,N_6349,N_6050);
nand U6687 (N_6687,N_6105,N_6272);
and U6688 (N_6688,N_6094,N_6131);
xor U6689 (N_6689,N_6446,N_6265);
nand U6690 (N_6690,N_6364,N_6309);
and U6691 (N_6691,N_6430,N_6395);
and U6692 (N_6692,N_6048,N_6244);
and U6693 (N_6693,N_6151,N_6436);
and U6694 (N_6694,N_6011,N_6057);
or U6695 (N_6695,N_6208,N_6387);
xnor U6696 (N_6696,N_6407,N_6301);
xor U6697 (N_6697,N_6231,N_6103);
nand U6698 (N_6698,N_6120,N_6214);
nor U6699 (N_6699,N_6166,N_6213);
nor U6700 (N_6700,N_6421,N_6489);
or U6701 (N_6701,N_6260,N_6433);
xor U6702 (N_6702,N_6233,N_6066);
nand U6703 (N_6703,N_6001,N_6173);
and U6704 (N_6704,N_6320,N_6287);
nand U6705 (N_6705,N_6363,N_6206);
xor U6706 (N_6706,N_6137,N_6201);
xor U6707 (N_6707,N_6142,N_6093);
xnor U6708 (N_6708,N_6177,N_6261);
nand U6709 (N_6709,N_6392,N_6202);
and U6710 (N_6710,N_6296,N_6167);
xnor U6711 (N_6711,N_6079,N_6069);
nand U6712 (N_6712,N_6459,N_6402);
xnor U6713 (N_6713,N_6161,N_6425);
nand U6714 (N_6714,N_6223,N_6203);
nor U6715 (N_6715,N_6088,N_6053);
or U6716 (N_6716,N_6010,N_6044);
nand U6717 (N_6717,N_6232,N_6328);
nor U6718 (N_6718,N_6418,N_6036);
and U6719 (N_6719,N_6176,N_6000);
nor U6720 (N_6720,N_6332,N_6341);
and U6721 (N_6721,N_6175,N_6178);
nand U6722 (N_6722,N_6324,N_6466);
and U6723 (N_6723,N_6289,N_6032);
and U6724 (N_6724,N_6004,N_6257);
nand U6725 (N_6725,N_6007,N_6441);
xor U6726 (N_6726,N_6118,N_6219);
nor U6727 (N_6727,N_6373,N_6391);
and U6728 (N_6728,N_6075,N_6338);
xnor U6729 (N_6729,N_6325,N_6292);
or U6730 (N_6730,N_6307,N_6339);
nor U6731 (N_6731,N_6061,N_6336);
nor U6732 (N_6732,N_6479,N_6143);
nand U6733 (N_6733,N_6458,N_6205);
xor U6734 (N_6734,N_6113,N_6008);
and U6735 (N_6735,N_6389,N_6316);
and U6736 (N_6736,N_6278,N_6462);
xnor U6737 (N_6737,N_6483,N_6452);
and U6738 (N_6738,N_6012,N_6062);
nor U6739 (N_6739,N_6431,N_6091);
or U6740 (N_6740,N_6367,N_6106);
or U6741 (N_6741,N_6037,N_6045);
nand U6742 (N_6742,N_6182,N_6255);
xnor U6743 (N_6743,N_6491,N_6409);
or U6744 (N_6744,N_6058,N_6081);
nor U6745 (N_6745,N_6217,N_6365);
xor U6746 (N_6746,N_6377,N_6308);
or U6747 (N_6747,N_6067,N_6487);
nand U6748 (N_6748,N_6468,N_6099);
nor U6749 (N_6749,N_6092,N_6457);
or U6750 (N_6750,N_6264,N_6183);
nor U6751 (N_6751,N_6144,N_6481);
and U6752 (N_6752,N_6038,N_6476);
nand U6753 (N_6753,N_6290,N_6421);
and U6754 (N_6754,N_6026,N_6465);
xor U6755 (N_6755,N_6225,N_6041);
nand U6756 (N_6756,N_6083,N_6471);
nand U6757 (N_6757,N_6005,N_6474);
nand U6758 (N_6758,N_6063,N_6320);
or U6759 (N_6759,N_6449,N_6075);
xor U6760 (N_6760,N_6108,N_6319);
nor U6761 (N_6761,N_6027,N_6373);
and U6762 (N_6762,N_6209,N_6304);
or U6763 (N_6763,N_6494,N_6261);
or U6764 (N_6764,N_6032,N_6391);
nand U6765 (N_6765,N_6170,N_6003);
nor U6766 (N_6766,N_6456,N_6414);
nor U6767 (N_6767,N_6204,N_6401);
or U6768 (N_6768,N_6403,N_6314);
xor U6769 (N_6769,N_6129,N_6405);
or U6770 (N_6770,N_6460,N_6006);
nand U6771 (N_6771,N_6071,N_6145);
and U6772 (N_6772,N_6404,N_6048);
nand U6773 (N_6773,N_6215,N_6236);
xnor U6774 (N_6774,N_6009,N_6056);
and U6775 (N_6775,N_6465,N_6273);
or U6776 (N_6776,N_6114,N_6375);
and U6777 (N_6777,N_6207,N_6379);
and U6778 (N_6778,N_6343,N_6390);
nand U6779 (N_6779,N_6446,N_6298);
nor U6780 (N_6780,N_6250,N_6078);
nor U6781 (N_6781,N_6457,N_6366);
or U6782 (N_6782,N_6278,N_6034);
and U6783 (N_6783,N_6294,N_6196);
nand U6784 (N_6784,N_6161,N_6411);
nor U6785 (N_6785,N_6123,N_6430);
nand U6786 (N_6786,N_6024,N_6043);
nor U6787 (N_6787,N_6400,N_6039);
xor U6788 (N_6788,N_6335,N_6085);
nor U6789 (N_6789,N_6220,N_6373);
nand U6790 (N_6790,N_6128,N_6462);
xnor U6791 (N_6791,N_6166,N_6139);
and U6792 (N_6792,N_6013,N_6408);
nor U6793 (N_6793,N_6086,N_6148);
and U6794 (N_6794,N_6084,N_6409);
xnor U6795 (N_6795,N_6440,N_6419);
xor U6796 (N_6796,N_6069,N_6277);
nor U6797 (N_6797,N_6447,N_6398);
or U6798 (N_6798,N_6391,N_6249);
xnor U6799 (N_6799,N_6234,N_6018);
and U6800 (N_6800,N_6430,N_6015);
xnor U6801 (N_6801,N_6024,N_6238);
or U6802 (N_6802,N_6161,N_6476);
nand U6803 (N_6803,N_6496,N_6347);
nand U6804 (N_6804,N_6386,N_6395);
nand U6805 (N_6805,N_6100,N_6418);
and U6806 (N_6806,N_6303,N_6218);
or U6807 (N_6807,N_6495,N_6089);
nor U6808 (N_6808,N_6383,N_6158);
nor U6809 (N_6809,N_6411,N_6470);
nor U6810 (N_6810,N_6096,N_6089);
and U6811 (N_6811,N_6044,N_6291);
and U6812 (N_6812,N_6336,N_6109);
or U6813 (N_6813,N_6262,N_6136);
and U6814 (N_6814,N_6348,N_6319);
and U6815 (N_6815,N_6376,N_6111);
xor U6816 (N_6816,N_6121,N_6297);
nor U6817 (N_6817,N_6374,N_6218);
nand U6818 (N_6818,N_6499,N_6049);
nand U6819 (N_6819,N_6046,N_6259);
nor U6820 (N_6820,N_6063,N_6230);
or U6821 (N_6821,N_6499,N_6342);
xor U6822 (N_6822,N_6032,N_6038);
or U6823 (N_6823,N_6143,N_6395);
xnor U6824 (N_6824,N_6407,N_6134);
xnor U6825 (N_6825,N_6109,N_6426);
or U6826 (N_6826,N_6304,N_6079);
nor U6827 (N_6827,N_6252,N_6095);
or U6828 (N_6828,N_6456,N_6210);
or U6829 (N_6829,N_6024,N_6487);
xnor U6830 (N_6830,N_6437,N_6209);
and U6831 (N_6831,N_6428,N_6154);
xor U6832 (N_6832,N_6043,N_6185);
and U6833 (N_6833,N_6299,N_6059);
nand U6834 (N_6834,N_6390,N_6209);
nor U6835 (N_6835,N_6360,N_6214);
nand U6836 (N_6836,N_6448,N_6453);
and U6837 (N_6837,N_6041,N_6285);
or U6838 (N_6838,N_6363,N_6178);
xor U6839 (N_6839,N_6494,N_6281);
nand U6840 (N_6840,N_6426,N_6288);
xor U6841 (N_6841,N_6089,N_6247);
xor U6842 (N_6842,N_6226,N_6326);
or U6843 (N_6843,N_6062,N_6211);
or U6844 (N_6844,N_6015,N_6174);
and U6845 (N_6845,N_6032,N_6418);
nand U6846 (N_6846,N_6477,N_6178);
and U6847 (N_6847,N_6095,N_6367);
and U6848 (N_6848,N_6174,N_6018);
and U6849 (N_6849,N_6436,N_6084);
and U6850 (N_6850,N_6115,N_6264);
and U6851 (N_6851,N_6274,N_6046);
nor U6852 (N_6852,N_6330,N_6144);
nand U6853 (N_6853,N_6077,N_6126);
nand U6854 (N_6854,N_6398,N_6059);
nor U6855 (N_6855,N_6478,N_6334);
or U6856 (N_6856,N_6295,N_6160);
nand U6857 (N_6857,N_6410,N_6050);
nor U6858 (N_6858,N_6328,N_6072);
and U6859 (N_6859,N_6202,N_6165);
and U6860 (N_6860,N_6395,N_6284);
xor U6861 (N_6861,N_6028,N_6191);
or U6862 (N_6862,N_6226,N_6284);
or U6863 (N_6863,N_6303,N_6380);
nor U6864 (N_6864,N_6486,N_6452);
and U6865 (N_6865,N_6244,N_6061);
or U6866 (N_6866,N_6188,N_6482);
and U6867 (N_6867,N_6400,N_6439);
or U6868 (N_6868,N_6123,N_6399);
nor U6869 (N_6869,N_6429,N_6353);
nand U6870 (N_6870,N_6471,N_6088);
xnor U6871 (N_6871,N_6264,N_6182);
nand U6872 (N_6872,N_6338,N_6155);
xor U6873 (N_6873,N_6401,N_6044);
nand U6874 (N_6874,N_6139,N_6439);
nor U6875 (N_6875,N_6384,N_6462);
or U6876 (N_6876,N_6089,N_6216);
nor U6877 (N_6877,N_6171,N_6041);
xnor U6878 (N_6878,N_6475,N_6473);
nand U6879 (N_6879,N_6388,N_6337);
or U6880 (N_6880,N_6270,N_6223);
nand U6881 (N_6881,N_6371,N_6432);
nand U6882 (N_6882,N_6478,N_6286);
and U6883 (N_6883,N_6373,N_6348);
nor U6884 (N_6884,N_6301,N_6365);
and U6885 (N_6885,N_6185,N_6262);
nand U6886 (N_6886,N_6142,N_6300);
or U6887 (N_6887,N_6452,N_6145);
nand U6888 (N_6888,N_6197,N_6020);
nor U6889 (N_6889,N_6273,N_6422);
nand U6890 (N_6890,N_6144,N_6132);
nand U6891 (N_6891,N_6074,N_6166);
xor U6892 (N_6892,N_6398,N_6070);
and U6893 (N_6893,N_6475,N_6010);
or U6894 (N_6894,N_6286,N_6281);
or U6895 (N_6895,N_6478,N_6322);
xnor U6896 (N_6896,N_6183,N_6360);
nor U6897 (N_6897,N_6262,N_6219);
and U6898 (N_6898,N_6055,N_6387);
xor U6899 (N_6899,N_6433,N_6156);
nor U6900 (N_6900,N_6059,N_6228);
nor U6901 (N_6901,N_6404,N_6219);
and U6902 (N_6902,N_6466,N_6089);
and U6903 (N_6903,N_6132,N_6143);
xor U6904 (N_6904,N_6029,N_6190);
or U6905 (N_6905,N_6438,N_6147);
nand U6906 (N_6906,N_6351,N_6377);
or U6907 (N_6907,N_6242,N_6417);
xnor U6908 (N_6908,N_6051,N_6291);
nand U6909 (N_6909,N_6325,N_6015);
xor U6910 (N_6910,N_6146,N_6440);
nand U6911 (N_6911,N_6267,N_6410);
nor U6912 (N_6912,N_6448,N_6027);
nor U6913 (N_6913,N_6415,N_6191);
nor U6914 (N_6914,N_6438,N_6471);
xor U6915 (N_6915,N_6359,N_6190);
and U6916 (N_6916,N_6240,N_6002);
nand U6917 (N_6917,N_6376,N_6049);
and U6918 (N_6918,N_6049,N_6295);
nand U6919 (N_6919,N_6188,N_6002);
xor U6920 (N_6920,N_6107,N_6102);
or U6921 (N_6921,N_6084,N_6206);
nand U6922 (N_6922,N_6234,N_6199);
xnor U6923 (N_6923,N_6320,N_6427);
and U6924 (N_6924,N_6266,N_6246);
nor U6925 (N_6925,N_6281,N_6274);
xor U6926 (N_6926,N_6006,N_6028);
or U6927 (N_6927,N_6477,N_6010);
nand U6928 (N_6928,N_6443,N_6344);
nand U6929 (N_6929,N_6236,N_6024);
and U6930 (N_6930,N_6084,N_6088);
nand U6931 (N_6931,N_6094,N_6463);
xor U6932 (N_6932,N_6289,N_6484);
nor U6933 (N_6933,N_6348,N_6070);
nand U6934 (N_6934,N_6457,N_6348);
nand U6935 (N_6935,N_6391,N_6206);
and U6936 (N_6936,N_6319,N_6122);
nor U6937 (N_6937,N_6476,N_6225);
or U6938 (N_6938,N_6195,N_6082);
nand U6939 (N_6939,N_6216,N_6428);
nor U6940 (N_6940,N_6290,N_6207);
nand U6941 (N_6941,N_6362,N_6203);
or U6942 (N_6942,N_6452,N_6052);
nor U6943 (N_6943,N_6425,N_6001);
or U6944 (N_6944,N_6136,N_6342);
xnor U6945 (N_6945,N_6234,N_6149);
xor U6946 (N_6946,N_6143,N_6105);
and U6947 (N_6947,N_6417,N_6002);
xnor U6948 (N_6948,N_6237,N_6031);
nand U6949 (N_6949,N_6475,N_6048);
xor U6950 (N_6950,N_6447,N_6407);
and U6951 (N_6951,N_6265,N_6494);
or U6952 (N_6952,N_6052,N_6303);
or U6953 (N_6953,N_6324,N_6301);
nand U6954 (N_6954,N_6216,N_6118);
and U6955 (N_6955,N_6029,N_6266);
and U6956 (N_6956,N_6205,N_6185);
nor U6957 (N_6957,N_6498,N_6483);
xnor U6958 (N_6958,N_6329,N_6127);
nand U6959 (N_6959,N_6353,N_6119);
xnor U6960 (N_6960,N_6004,N_6430);
nand U6961 (N_6961,N_6474,N_6122);
nor U6962 (N_6962,N_6085,N_6121);
nand U6963 (N_6963,N_6416,N_6187);
or U6964 (N_6964,N_6497,N_6308);
or U6965 (N_6965,N_6190,N_6478);
or U6966 (N_6966,N_6331,N_6189);
or U6967 (N_6967,N_6294,N_6490);
or U6968 (N_6968,N_6311,N_6104);
nor U6969 (N_6969,N_6471,N_6385);
nand U6970 (N_6970,N_6109,N_6411);
xor U6971 (N_6971,N_6323,N_6216);
or U6972 (N_6972,N_6464,N_6395);
nor U6973 (N_6973,N_6124,N_6178);
nor U6974 (N_6974,N_6497,N_6236);
nor U6975 (N_6975,N_6044,N_6057);
nor U6976 (N_6976,N_6068,N_6397);
xor U6977 (N_6977,N_6202,N_6452);
and U6978 (N_6978,N_6354,N_6338);
nor U6979 (N_6979,N_6317,N_6351);
nor U6980 (N_6980,N_6152,N_6209);
nand U6981 (N_6981,N_6376,N_6214);
nor U6982 (N_6982,N_6026,N_6227);
and U6983 (N_6983,N_6265,N_6032);
nor U6984 (N_6984,N_6081,N_6242);
xnor U6985 (N_6985,N_6240,N_6139);
nor U6986 (N_6986,N_6397,N_6423);
and U6987 (N_6987,N_6206,N_6113);
and U6988 (N_6988,N_6496,N_6393);
nor U6989 (N_6989,N_6429,N_6485);
or U6990 (N_6990,N_6237,N_6300);
and U6991 (N_6991,N_6082,N_6051);
nand U6992 (N_6992,N_6152,N_6403);
xor U6993 (N_6993,N_6162,N_6407);
nor U6994 (N_6994,N_6285,N_6091);
nor U6995 (N_6995,N_6230,N_6263);
and U6996 (N_6996,N_6330,N_6218);
nor U6997 (N_6997,N_6143,N_6423);
nand U6998 (N_6998,N_6308,N_6155);
xor U6999 (N_6999,N_6005,N_6232);
and U7000 (N_7000,N_6820,N_6798);
or U7001 (N_7001,N_6700,N_6924);
nor U7002 (N_7002,N_6861,N_6911);
or U7003 (N_7003,N_6819,N_6988);
or U7004 (N_7004,N_6559,N_6829);
or U7005 (N_7005,N_6893,N_6702);
or U7006 (N_7006,N_6895,N_6909);
nand U7007 (N_7007,N_6747,N_6965);
or U7008 (N_7008,N_6766,N_6512);
nor U7009 (N_7009,N_6603,N_6553);
nor U7010 (N_7010,N_6576,N_6549);
and U7011 (N_7011,N_6767,N_6502);
and U7012 (N_7012,N_6772,N_6945);
nor U7013 (N_7013,N_6606,N_6572);
and U7014 (N_7014,N_6503,N_6908);
nor U7015 (N_7015,N_6735,N_6785);
or U7016 (N_7016,N_6540,N_6511);
and U7017 (N_7017,N_6703,N_6646);
and U7018 (N_7018,N_6952,N_6532);
or U7019 (N_7019,N_6590,N_6625);
nand U7020 (N_7020,N_6964,N_6501);
or U7021 (N_7021,N_6922,N_6634);
or U7022 (N_7022,N_6726,N_6866);
and U7023 (N_7023,N_6818,N_6834);
and U7024 (N_7024,N_6942,N_6710);
nand U7025 (N_7025,N_6896,N_6867);
nand U7026 (N_7026,N_6848,N_6966);
nand U7027 (N_7027,N_6812,N_6684);
and U7028 (N_7028,N_6672,N_6890);
nor U7029 (N_7029,N_6627,N_6705);
nor U7030 (N_7030,N_6959,N_6816);
or U7031 (N_7031,N_6782,N_6529);
and U7032 (N_7032,N_6806,N_6935);
and U7033 (N_7033,N_6982,N_6611);
and U7034 (N_7034,N_6873,N_6668);
nor U7035 (N_7035,N_6915,N_6980);
and U7036 (N_7036,N_6881,N_6566);
nor U7037 (N_7037,N_6811,N_6976);
nand U7038 (N_7038,N_6530,N_6989);
or U7039 (N_7039,N_6994,N_6796);
or U7040 (N_7040,N_6738,N_6729);
xnor U7041 (N_7041,N_6904,N_6991);
or U7042 (N_7042,N_6651,N_6649);
and U7043 (N_7043,N_6712,N_6773);
and U7044 (N_7044,N_6975,N_6783);
xnor U7045 (N_7045,N_6676,N_6780);
nand U7046 (N_7046,N_6583,N_6774);
nor U7047 (N_7047,N_6762,N_6564);
nor U7048 (N_7048,N_6516,N_6968);
nor U7049 (N_7049,N_6618,N_6894);
or U7050 (N_7050,N_6734,N_6906);
nor U7051 (N_7051,N_6602,N_6521);
nor U7052 (N_7052,N_6971,N_6841);
nor U7053 (N_7053,N_6856,N_6548);
and U7054 (N_7054,N_6888,N_6830);
nand U7055 (N_7055,N_6718,N_6657);
and U7056 (N_7056,N_6872,N_6674);
nand U7057 (N_7057,N_6565,N_6750);
and U7058 (N_7058,N_6775,N_6597);
nand U7059 (N_7059,N_6949,N_6793);
xor U7060 (N_7060,N_6821,N_6510);
or U7061 (N_7061,N_6641,N_6573);
nand U7062 (N_7062,N_6876,N_6679);
and U7063 (N_7063,N_6912,N_6917);
nand U7064 (N_7064,N_6940,N_6778);
or U7065 (N_7065,N_6685,N_6822);
xor U7066 (N_7066,N_6831,N_6577);
or U7067 (N_7067,N_6507,N_6630);
nand U7068 (N_7068,N_6944,N_6687);
nor U7069 (N_7069,N_6779,N_6732);
xor U7070 (N_7070,N_6669,N_6858);
and U7071 (N_7071,N_6961,N_6561);
nand U7072 (N_7072,N_6955,N_6997);
nor U7073 (N_7073,N_6931,N_6790);
nor U7074 (N_7074,N_6616,N_6804);
nor U7075 (N_7075,N_6644,N_6595);
and U7076 (N_7076,N_6659,N_6619);
or U7077 (N_7077,N_6707,N_6531);
nand U7078 (N_7078,N_6857,N_6926);
nor U7079 (N_7079,N_6575,N_6562);
and U7080 (N_7080,N_6981,N_6607);
or U7081 (N_7081,N_6792,N_6905);
nand U7082 (N_7082,N_6675,N_6589);
nand U7083 (N_7083,N_6591,N_6621);
nand U7084 (N_7084,N_6697,N_6560);
nor U7085 (N_7085,N_6882,N_6992);
nor U7086 (N_7086,N_6826,N_6520);
nor U7087 (N_7087,N_6533,N_6862);
nand U7088 (N_7088,N_6608,N_6805);
and U7089 (N_7089,N_6626,N_6724);
nand U7090 (N_7090,N_6683,N_6835);
or U7091 (N_7091,N_6730,N_6875);
xor U7092 (N_7092,N_6728,N_6535);
or U7093 (N_7093,N_6950,N_6614);
nand U7094 (N_7094,N_6938,N_6752);
and U7095 (N_7095,N_6941,N_6787);
or U7096 (N_7096,N_6956,N_6715);
nor U7097 (N_7097,N_6693,N_6877);
or U7098 (N_7098,N_6680,N_6939);
nor U7099 (N_7099,N_6719,N_6682);
or U7100 (N_7100,N_6681,N_6943);
nand U7101 (N_7101,N_6996,N_6586);
xnor U7102 (N_7102,N_6839,N_6765);
xor U7103 (N_7103,N_6656,N_6967);
nand U7104 (N_7104,N_6517,N_6665);
and U7105 (N_7105,N_6574,N_6828);
and U7106 (N_7106,N_6901,N_6556);
nor U7107 (N_7107,N_6568,N_6593);
xnor U7108 (N_7108,N_6527,N_6654);
nor U7109 (N_7109,N_6789,N_6899);
xnor U7110 (N_7110,N_6868,N_6550);
xor U7111 (N_7111,N_6795,N_6714);
and U7112 (N_7112,N_6761,N_6689);
or U7113 (N_7113,N_6515,N_6743);
xor U7114 (N_7114,N_6701,N_6617);
nor U7115 (N_7115,N_6581,N_6716);
xor U7116 (N_7116,N_6541,N_6919);
nand U7117 (N_7117,N_6769,N_6846);
and U7118 (N_7118,N_6757,N_6628);
or U7119 (N_7119,N_6802,N_6612);
xnor U7120 (N_7120,N_6837,N_6652);
nor U7121 (N_7121,N_6889,N_6538);
nor U7122 (N_7122,N_6983,N_6690);
nor U7123 (N_7123,N_6671,N_6869);
nor U7124 (N_7124,N_6708,N_6579);
and U7125 (N_7125,N_6555,N_6933);
or U7126 (N_7126,N_6923,N_6544);
nand U7127 (N_7127,N_6797,N_6883);
nor U7128 (N_7128,N_6620,N_6963);
nand U7129 (N_7129,N_6633,N_6986);
nor U7130 (N_7130,N_6695,N_6755);
xor U7131 (N_7131,N_6648,N_6696);
nor U7132 (N_7132,N_6613,N_6918);
and U7133 (N_7133,N_6973,N_6885);
and U7134 (N_7134,N_6999,N_6760);
or U7135 (N_7135,N_6920,N_6984);
nor U7136 (N_7136,N_6998,N_6580);
nand U7137 (N_7137,N_6946,N_6892);
xor U7138 (N_7138,N_6914,N_6514);
xor U7139 (N_7139,N_6596,N_6709);
nor U7140 (N_7140,N_6523,N_6658);
nand U7141 (N_7141,N_6969,N_6592);
nand U7142 (N_7142,N_6850,N_6958);
nand U7143 (N_7143,N_6860,N_6810);
nand U7144 (N_7144,N_6957,N_6645);
nor U7145 (N_7145,N_6635,N_6666);
nor U7146 (N_7146,N_6637,N_6903);
xor U7147 (N_7147,N_6587,N_6929);
nand U7148 (N_7148,N_6836,N_6610);
nor U7149 (N_7149,N_6954,N_6542);
nor U7150 (N_7150,N_6640,N_6803);
nor U7151 (N_7151,N_6692,N_6800);
xnor U7152 (N_7152,N_6777,N_6629);
xor U7153 (N_7153,N_6642,N_6552);
or U7154 (N_7154,N_6519,N_6653);
xor U7155 (N_7155,N_6563,N_6985);
nor U7156 (N_7156,N_6878,N_6605);
and U7157 (N_7157,N_6539,N_6814);
xor U7158 (N_7158,N_6733,N_6827);
or U7159 (N_7159,N_6825,N_6739);
and U7160 (N_7160,N_6727,N_6815);
nand U7161 (N_7161,N_6849,N_6788);
nor U7162 (N_7162,N_6764,N_6809);
nand U7163 (N_7163,N_6722,N_6534);
nor U7164 (N_7164,N_6694,N_6751);
and U7165 (N_7165,N_6673,N_6887);
nand U7166 (N_7166,N_6910,N_6664);
nor U7167 (N_7167,N_6677,N_6513);
or U7168 (N_7168,N_6578,N_6742);
or U7169 (N_7169,N_6844,N_6756);
or U7170 (N_7170,N_6748,N_6691);
or U7171 (N_7171,N_6588,N_6706);
xor U7172 (N_7172,N_6737,N_6987);
nor U7173 (N_7173,N_6655,N_6522);
and U7174 (N_7174,N_6960,N_6636);
nand U7175 (N_7175,N_6855,N_6870);
or U7176 (N_7176,N_6504,N_6970);
xnor U7177 (N_7177,N_6509,N_6801);
and U7178 (N_7178,N_6604,N_6884);
nor U7179 (N_7179,N_6930,N_6643);
nand U7180 (N_7180,N_6546,N_6731);
nand U7181 (N_7181,N_6601,N_6832);
or U7182 (N_7182,N_6817,N_6907);
or U7183 (N_7183,N_6799,N_6500);
nor U7184 (N_7184,N_6662,N_6554);
nor U7185 (N_7185,N_6927,N_6528);
and U7186 (N_7186,N_6784,N_6661);
and U7187 (N_7187,N_6947,N_6854);
xnor U7188 (N_7188,N_6663,N_6928);
and U7189 (N_7189,N_6824,N_6688);
nand U7190 (N_7190,N_6660,N_6838);
nand U7191 (N_7191,N_6874,N_6741);
and U7192 (N_7192,N_6746,N_6758);
nor U7193 (N_7193,N_6537,N_6678);
nor U7194 (N_7194,N_6740,N_6686);
or U7195 (N_7195,N_6557,N_6951);
xnor U7196 (N_7196,N_6978,N_6995);
xor U7197 (N_7197,N_6768,N_6993);
or U7198 (N_7198,N_6624,N_6932);
or U7199 (N_7199,N_6979,N_6711);
and U7200 (N_7200,N_6585,N_6632);
nand U7201 (N_7201,N_6647,N_6851);
or U7202 (N_7202,N_6843,N_6536);
and U7203 (N_7203,N_6598,N_6852);
nor U7204 (N_7204,N_6865,N_6667);
nor U7205 (N_7205,N_6847,N_6582);
and U7206 (N_7206,N_6759,N_6807);
xor U7207 (N_7207,N_6545,N_6720);
nand U7208 (N_7208,N_6725,N_6921);
xnor U7209 (N_7209,N_6886,N_6753);
nand U7210 (N_7210,N_6525,N_6948);
xnor U7211 (N_7211,N_6505,N_6900);
nand U7212 (N_7212,N_6763,N_6990);
nor U7213 (N_7213,N_6571,N_6823);
and U7214 (N_7214,N_6754,N_6879);
and U7215 (N_7215,N_6615,N_6749);
xnor U7216 (N_7216,N_6526,N_6840);
xor U7217 (N_7217,N_6925,N_6853);
nor U7218 (N_7218,N_6977,N_6813);
xnor U7219 (N_7219,N_6781,N_6770);
nand U7220 (N_7220,N_6551,N_6786);
nand U7221 (N_7221,N_6639,N_6913);
or U7222 (N_7222,N_6745,N_6833);
nor U7223 (N_7223,N_6937,N_6699);
xnor U7224 (N_7224,N_6771,N_6974);
nor U7225 (N_7225,N_6736,N_6570);
nor U7226 (N_7226,N_6936,N_6808);
nor U7227 (N_7227,N_6547,N_6650);
xnor U7228 (N_7228,N_6791,N_6670);
or U7229 (N_7229,N_6622,N_6744);
nand U7230 (N_7230,N_6916,N_6569);
or U7231 (N_7231,N_6594,N_6508);
xnor U7232 (N_7232,N_6902,N_6859);
and U7233 (N_7233,N_6891,N_6543);
and U7234 (N_7234,N_6897,N_6864);
nand U7235 (N_7235,N_6623,N_6776);
nand U7236 (N_7236,N_6953,N_6972);
and U7237 (N_7237,N_6609,N_6898);
nor U7238 (N_7238,N_6845,N_6567);
and U7239 (N_7239,N_6600,N_6713);
nor U7240 (N_7240,N_6599,N_6704);
or U7241 (N_7241,N_6723,N_6717);
nand U7242 (N_7242,N_6880,N_6962);
nor U7243 (N_7243,N_6558,N_6524);
and U7244 (N_7244,N_6506,N_6871);
nand U7245 (N_7245,N_6842,N_6863);
nor U7246 (N_7246,N_6638,N_6721);
and U7247 (N_7247,N_6934,N_6631);
nand U7248 (N_7248,N_6518,N_6794);
or U7249 (N_7249,N_6698,N_6584);
xnor U7250 (N_7250,N_6659,N_6704);
and U7251 (N_7251,N_6608,N_6814);
nor U7252 (N_7252,N_6657,N_6741);
and U7253 (N_7253,N_6682,N_6981);
xnor U7254 (N_7254,N_6527,N_6851);
xor U7255 (N_7255,N_6645,N_6538);
and U7256 (N_7256,N_6555,N_6645);
nand U7257 (N_7257,N_6623,N_6920);
nor U7258 (N_7258,N_6582,N_6915);
and U7259 (N_7259,N_6983,N_6780);
nand U7260 (N_7260,N_6887,N_6967);
and U7261 (N_7261,N_6706,N_6907);
xor U7262 (N_7262,N_6673,N_6770);
nand U7263 (N_7263,N_6501,N_6724);
nand U7264 (N_7264,N_6930,N_6529);
nand U7265 (N_7265,N_6760,N_6785);
and U7266 (N_7266,N_6642,N_6878);
and U7267 (N_7267,N_6647,N_6761);
nand U7268 (N_7268,N_6913,N_6659);
or U7269 (N_7269,N_6634,N_6520);
nand U7270 (N_7270,N_6696,N_6686);
nor U7271 (N_7271,N_6741,N_6869);
and U7272 (N_7272,N_6733,N_6720);
or U7273 (N_7273,N_6605,N_6551);
nand U7274 (N_7274,N_6605,N_6675);
nor U7275 (N_7275,N_6532,N_6589);
and U7276 (N_7276,N_6727,N_6992);
xor U7277 (N_7277,N_6519,N_6831);
and U7278 (N_7278,N_6932,N_6725);
or U7279 (N_7279,N_6686,N_6866);
xnor U7280 (N_7280,N_6906,N_6893);
and U7281 (N_7281,N_6824,N_6986);
xnor U7282 (N_7282,N_6612,N_6564);
nor U7283 (N_7283,N_6754,N_6852);
nor U7284 (N_7284,N_6924,N_6746);
nand U7285 (N_7285,N_6611,N_6549);
and U7286 (N_7286,N_6561,N_6590);
nor U7287 (N_7287,N_6644,N_6964);
or U7288 (N_7288,N_6622,N_6505);
xor U7289 (N_7289,N_6921,N_6601);
or U7290 (N_7290,N_6853,N_6574);
nand U7291 (N_7291,N_6568,N_6953);
nor U7292 (N_7292,N_6815,N_6697);
or U7293 (N_7293,N_6842,N_6671);
xnor U7294 (N_7294,N_6632,N_6909);
nor U7295 (N_7295,N_6515,N_6838);
and U7296 (N_7296,N_6532,N_6500);
nand U7297 (N_7297,N_6937,N_6707);
xnor U7298 (N_7298,N_6685,N_6692);
xnor U7299 (N_7299,N_6626,N_6933);
nor U7300 (N_7300,N_6760,N_6719);
nor U7301 (N_7301,N_6665,N_6562);
xor U7302 (N_7302,N_6816,N_6521);
nand U7303 (N_7303,N_6961,N_6874);
nor U7304 (N_7304,N_6620,N_6708);
nor U7305 (N_7305,N_6732,N_6723);
and U7306 (N_7306,N_6829,N_6731);
xnor U7307 (N_7307,N_6703,N_6987);
and U7308 (N_7308,N_6516,N_6512);
and U7309 (N_7309,N_6872,N_6890);
nand U7310 (N_7310,N_6917,N_6882);
and U7311 (N_7311,N_6586,N_6697);
and U7312 (N_7312,N_6672,N_6973);
or U7313 (N_7313,N_6531,N_6891);
xor U7314 (N_7314,N_6528,N_6961);
nand U7315 (N_7315,N_6958,N_6820);
and U7316 (N_7316,N_6527,N_6769);
xor U7317 (N_7317,N_6628,N_6840);
and U7318 (N_7318,N_6557,N_6847);
xnor U7319 (N_7319,N_6924,N_6722);
xor U7320 (N_7320,N_6702,N_6935);
nor U7321 (N_7321,N_6913,N_6834);
nor U7322 (N_7322,N_6763,N_6867);
or U7323 (N_7323,N_6527,N_6932);
nand U7324 (N_7324,N_6762,N_6864);
and U7325 (N_7325,N_6899,N_6690);
nand U7326 (N_7326,N_6763,N_6613);
or U7327 (N_7327,N_6878,N_6804);
nand U7328 (N_7328,N_6875,N_6599);
xnor U7329 (N_7329,N_6641,N_6980);
nor U7330 (N_7330,N_6656,N_6812);
nor U7331 (N_7331,N_6838,N_6578);
nand U7332 (N_7332,N_6958,N_6965);
xor U7333 (N_7333,N_6571,N_6566);
or U7334 (N_7334,N_6534,N_6950);
or U7335 (N_7335,N_6745,N_6659);
or U7336 (N_7336,N_6877,N_6955);
nor U7337 (N_7337,N_6965,N_6670);
nor U7338 (N_7338,N_6929,N_6520);
or U7339 (N_7339,N_6781,N_6618);
xor U7340 (N_7340,N_6715,N_6686);
or U7341 (N_7341,N_6797,N_6944);
xor U7342 (N_7342,N_6990,N_6819);
nor U7343 (N_7343,N_6812,N_6694);
and U7344 (N_7344,N_6720,N_6852);
nor U7345 (N_7345,N_6621,N_6826);
nor U7346 (N_7346,N_6723,N_6888);
and U7347 (N_7347,N_6834,N_6752);
and U7348 (N_7348,N_6797,N_6931);
and U7349 (N_7349,N_6769,N_6819);
xor U7350 (N_7350,N_6530,N_6696);
or U7351 (N_7351,N_6503,N_6615);
nand U7352 (N_7352,N_6878,N_6624);
xnor U7353 (N_7353,N_6719,N_6750);
and U7354 (N_7354,N_6842,N_6593);
xnor U7355 (N_7355,N_6517,N_6939);
xor U7356 (N_7356,N_6544,N_6725);
or U7357 (N_7357,N_6646,N_6689);
and U7358 (N_7358,N_6507,N_6514);
nand U7359 (N_7359,N_6981,N_6879);
nand U7360 (N_7360,N_6638,N_6538);
or U7361 (N_7361,N_6559,N_6964);
nor U7362 (N_7362,N_6801,N_6925);
xnor U7363 (N_7363,N_6882,N_6896);
nor U7364 (N_7364,N_6766,N_6558);
nor U7365 (N_7365,N_6708,N_6851);
or U7366 (N_7366,N_6880,N_6845);
or U7367 (N_7367,N_6582,N_6905);
nor U7368 (N_7368,N_6794,N_6750);
and U7369 (N_7369,N_6621,N_6817);
nand U7370 (N_7370,N_6971,N_6730);
or U7371 (N_7371,N_6630,N_6861);
nand U7372 (N_7372,N_6591,N_6560);
and U7373 (N_7373,N_6910,N_6646);
or U7374 (N_7374,N_6779,N_6915);
nor U7375 (N_7375,N_6762,N_6956);
and U7376 (N_7376,N_6640,N_6586);
nand U7377 (N_7377,N_6991,N_6796);
nand U7378 (N_7378,N_6963,N_6608);
nor U7379 (N_7379,N_6872,N_6859);
and U7380 (N_7380,N_6899,N_6865);
xor U7381 (N_7381,N_6634,N_6681);
nor U7382 (N_7382,N_6808,N_6977);
and U7383 (N_7383,N_6790,N_6600);
xnor U7384 (N_7384,N_6538,N_6865);
nand U7385 (N_7385,N_6552,N_6863);
and U7386 (N_7386,N_6852,N_6914);
nand U7387 (N_7387,N_6977,N_6782);
nor U7388 (N_7388,N_6583,N_6903);
or U7389 (N_7389,N_6637,N_6717);
or U7390 (N_7390,N_6573,N_6894);
or U7391 (N_7391,N_6977,N_6510);
and U7392 (N_7392,N_6629,N_6584);
nand U7393 (N_7393,N_6603,N_6911);
and U7394 (N_7394,N_6751,N_6793);
and U7395 (N_7395,N_6800,N_6890);
nor U7396 (N_7396,N_6852,N_6984);
and U7397 (N_7397,N_6922,N_6917);
or U7398 (N_7398,N_6772,N_6550);
and U7399 (N_7399,N_6919,N_6935);
xor U7400 (N_7400,N_6749,N_6791);
xnor U7401 (N_7401,N_6941,N_6729);
xnor U7402 (N_7402,N_6638,N_6873);
xor U7403 (N_7403,N_6875,N_6989);
nor U7404 (N_7404,N_6763,N_6826);
or U7405 (N_7405,N_6765,N_6842);
or U7406 (N_7406,N_6620,N_6875);
or U7407 (N_7407,N_6968,N_6917);
or U7408 (N_7408,N_6851,N_6638);
nor U7409 (N_7409,N_6626,N_6957);
nand U7410 (N_7410,N_6825,N_6756);
or U7411 (N_7411,N_6948,N_6930);
or U7412 (N_7412,N_6860,N_6962);
and U7413 (N_7413,N_6580,N_6583);
or U7414 (N_7414,N_6936,N_6855);
and U7415 (N_7415,N_6951,N_6576);
or U7416 (N_7416,N_6531,N_6745);
nor U7417 (N_7417,N_6541,N_6884);
nand U7418 (N_7418,N_6703,N_6831);
xor U7419 (N_7419,N_6998,N_6771);
or U7420 (N_7420,N_6921,N_6552);
nand U7421 (N_7421,N_6787,N_6605);
or U7422 (N_7422,N_6993,N_6973);
or U7423 (N_7423,N_6623,N_6931);
and U7424 (N_7424,N_6944,N_6931);
and U7425 (N_7425,N_6967,N_6603);
nor U7426 (N_7426,N_6942,N_6688);
or U7427 (N_7427,N_6866,N_6848);
nor U7428 (N_7428,N_6611,N_6687);
nor U7429 (N_7429,N_6538,N_6510);
or U7430 (N_7430,N_6540,N_6876);
nor U7431 (N_7431,N_6690,N_6876);
nor U7432 (N_7432,N_6955,N_6801);
nor U7433 (N_7433,N_6619,N_6654);
or U7434 (N_7434,N_6554,N_6762);
nor U7435 (N_7435,N_6551,N_6907);
and U7436 (N_7436,N_6817,N_6859);
xor U7437 (N_7437,N_6525,N_6764);
or U7438 (N_7438,N_6712,N_6639);
nand U7439 (N_7439,N_6878,N_6601);
xor U7440 (N_7440,N_6659,N_6644);
nor U7441 (N_7441,N_6527,N_6703);
nand U7442 (N_7442,N_6854,N_6724);
nand U7443 (N_7443,N_6914,N_6570);
nor U7444 (N_7444,N_6907,N_6879);
or U7445 (N_7445,N_6890,N_6698);
xor U7446 (N_7446,N_6505,N_6944);
or U7447 (N_7447,N_6674,N_6837);
nor U7448 (N_7448,N_6956,N_6695);
nand U7449 (N_7449,N_6808,N_6943);
and U7450 (N_7450,N_6960,N_6669);
nor U7451 (N_7451,N_6712,N_6884);
or U7452 (N_7452,N_6624,N_6796);
nor U7453 (N_7453,N_6625,N_6609);
or U7454 (N_7454,N_6533,N_6763);
or U7455 (N_7455,N_6732,N_6650);
and U7456 (N_7456,N_6705,N_6903);
and U7457 (N_7457,N_6823,N_6764);
nor U7458 (N_7458,N_6603,N_6753);
nand U7459 (N_7459,N_6822,N_6836);
xnor U7460 (N_7460,N_6800,N_6954);
xnor U7461 (N_7461,N_6766,N_6519);
and U7462 (N_7462,N_6976,N_6676);
and U7463 (N_7463,N_6731,N_6508);
nand U7464 (N_7464,N_6975,N_6712);
and U7465 (N_7465,N_6687,N_6566);
xnor U7466 (N_7466,N_6812,N_6840);
nand U7467 (N_7467,N_6589,N_6812);
nor U7468 (N_7468,N_6607,N_6911);
xnor U7469 (N_7469,N_6860,N_6918);
nand U7470 (N_7470,N_6927,N_6573);
nand U7471 (N_7471,N_6934,N_6871);
and U7472 (N_7472,N_6728,N_6669);
xor U7473 (N_7473,N_6700,N_6618);
xnor U7474 (N_7474,N_6585,N_6566);
or U7475 (N_7475,N_6936,N_6600);
and U7476 (N_7476,N_6764,N_6635);
and U7477 (N_7477,N_6561,N_6674);
or U7478 (N_7478,N_6785,N_6630);
xnor U7479 (N_7479,N_6802,N_6776);
nand U7480 (N_7480,N_6702,N_6828);
and U7481 (N_7481,N_6998,N_6676);
nand U7482 (N_7482,N_6560,N_6810);
or U7483 (N_7483,N_6983,N_6501);
or U7484 (N_7484,N_6775,N_6675);
nand U7485 (N_7485,N_6986,N_6669);
nor U7486 (N_7486,N_6780,N_6716);
nor U7487 (N_7487,N_6632,N_6661);
xor U7488 (N_7488,N_6683,N_6590);
and U7489 (N_7489,N_6830,N_6799);
and U7490 (N_7490,N_6981,N_6807);
and U7491 (N_7491,N_6910,N_6573);
xnor U7492 (N_7492,N_6634,N_6851);
nand U7493 (N_7493,N_6914,N_6565);
and U7494 (N_7494,N_6755,N_6626);
or U7495 (N_7495,N_6964,N_6831);
nor U7496 (N_7496,N_6517,N_6511);
xor U7497 (N_7497,N_6973,N_6699);
or U7498 (N_7498,N_6878,N_6888);
and U7499 (N_7499,N_6729,N_6959);
nor U7500 (N_7500,N_7381,N_7492);
or U7501 (N_7501,N_7173,N_7226);
and U7502 (N_7502,N_7064,N_7227);
nor U7503 (N_7503,N_7051,N_7355);
xor U7504 (N_7504,N_7360,N_7282);
or U7505 (N_7505,N_7272,N_7228);
nand U7506 (N_7506,N_7241,N_7224);
nand U7507 (N_7507,N_7102,N_7384);
nor U7508 (N_7508,N_7373,N_7335);
and U7509 (N_7509,N_7075,N_7038);
or U7510 (N_7510,N_7089,N_7451);
and U7511 (N_7511,N_7474,N_7138);
or U7512 (N_7512,N_7086,N_7047);
nand U7513 (N_7513,N_7255,N_7434);
nand U7514 (N_7514,N_7347,N_7039);
or U7515 (N_7515,N_7178,N_7020);
or U7516 (N_7516,N_7273,N_7092);
or U7517 (N_7517,N_7033,N_7285);
nor U7518 (N_7518,N_7495,N_7036);
or U7519 (N_7519,N_7367,N_7481);
and U7520 (N_7520,N_7304,N_7187);
or U7521 (N_7521,N_7419,N_7112);
and U7522 (N_7522,N_7498,N_7058);
and U7523 (N_7523,N_7259,N_7488);
xnor U7524 (N_7524,N_7052,N_7371);
and U7525 (N_7525,N_7029,N_7490);
and U7526 (N_7526,N_7127,N_7081);
or U7527 (N_7527,N_7164,N_7264);
nor U7528 (N_7528,N_7185,N_7095);
or U7529 (N_7529,N_7357,N_7310);
nor U7530 (N_7530,N_7030,N_7414);
or U7531 (N_7531,N_7471,N_7311);
nor U7532 (N_7532,N_7125,N_7026);
and U7533 (N_7533,N_7364,N_7293);
nor U7534 (N_7534,N_7176,N_7453);
xor U7535 (N_7535,N_7231,N_7175);
or U7536 (N_7536,N_7210,N_7337);
and U7537 (N_7537,N_7115,N_7216);
nor U7538 (N_7538,N_7254,N_7197);
xnor U7539 (N_7539,N_7014,N_7324);
and U7540 (N_7540,N_7237,N_7244);
nor U7541 (N_7541,N_7374,N_7076);
or U7542 (N_7542,N_7363,N_7499);
nand U7543 (N_7543,N_7019,N_7157);
or U7544 (N_7544,N_7236,N_7274);
nand U7545 (N_7545,N_7423,N_7467);
nor U7546 (N_7546,N_7417,N_7351);
nor U7547 (N_7547,N_7439,N_7462);
nand U7548 (N_7548,N_7289,N_7126);
and U7549 (N_7549,N_7249,N_7349);
xnor U7550 (N_7550,N_7486,N_7412);
nand U7551 (N_7551,N_7158,N_7121);
nor U7552 (N_7552,N_7234,N_7422);
nor U7553 (N_7553,N_7393,N_7378);
nand U7554 (N_7554,N_7483,N_7375);
nor U7555 (N_7555,N_7040,N_7493);
xor U7556 (N_7556,N_7097,N_7362);
or U7557 (N_7557,N_7330,N_7252);
nand U7558 (N_7558,N_7426,N_7457);
xor U7559 (N_7559,N_7093,N_7180);
nand U7560 (N_7560,N_7004,N_7010);
nor U7561 (N_7561,N_7012,N_7314);
xnor U7562 (N_7562,N_7268,N_7156);
xnor U7563 (N_7563,N_7025,N_7261);
and U7564 (N_7564,N_7204,N_7421);
xor U7565 (N_7565,N_7298,N_7122);
nor U7566 (N_7566,N_7416,N_7336);
and U7567 (N_7567,N_7031,N_7059);
xnor U7568 (N_7568,N_7160,N_7331);
nand U7569 (N_7569,N_7312,N_7369);
or U7570 (N_7570,N_7464,N_7461);
nand U7571 (N_7571,N_7099,N_7191);
and U7572 (N_7572,N_7222,N_7144);
xor U7573 (N_7573,N_7395,N_7452);
xnor U7574 (N_7574,N_7430,N_7319);
nand U7575 (N_7575,N_7005,N_7056);
xor U7576 (N_7576,N_7205,N_7281);
xnor U7577 (N_7577,N_7437,N_7079);
or U7578 (N_7578,N_7350,N_7403);
or U7579 (N_7579,N_7153,N_7410);
nor U7580 (N_7580,N_7090,N_7313);
and U7581 (N_7581,N_7400,N_7401);
nand U7582 (N_7582,N_7447,N_7267);
nor U7583 (N_7583,N_7209,N_7100);
and U7584 (N_7584,N_7391,N_7308);
xor U7585 (N_7585,N_7402,N_7168);
xor U7586 (N_7586,N_7271,N_7405);
xnor U7587 (N_7587,N_7015,N_7315);
nor U7588 (N_7588,N_7262,N_7466);
and U7589 (N_7589,N_7139,N_7361);
or U7590 (N_7590,N_7368,N_7379);
nor U7591 (N_7591,N_7141,N_7062);
nand U7592 (N_7592,N_7199,N_7151);
xor U7593 (N_7593,N_7078,N_7433);
and U7594 (N_7594,N_7415,N_7494);
or U7595 (N_7595,N_7303,N_7096);
or U7596 (N_7596,N_7161,N_7297);
nand U7597 (N_7597,N_7435,N_7195);
nor U7598 (N_7598,N_7235,N_7166);
xor U7599 (N_7599,N_7109,N_7444);
nor U7600 (N_7600,N_7256,N_7491);
nand U7601 (N_7601,N_7077,N_7009);
or U7602 (N_7602,N_7060,N_7049);
nor U7603 (N_7603,N_7003,N_7117);
or U7604 (N_7604,N_7063,N_7130);
xor U7605 (N_7605,N_7203,N_7084);
and U7606 (N_7606,N_7327,N_7398);
xnor U7607 (N_7607,N_7370,N_7061);
nor U7608 (N_7608,N_7449,N_7468);
xnor U7609 (N_7609,N_7027,N_7170);
xnor U7610 (N_7610,N_7406,N_7358);
nand U7611 (N_7611,N_7008,N_7154);
xor U7612 (N_7612,N_7334,N_7057);
and U7613 (N_7613,N_7066,N_7045);
xor U7614 (N_7614,N_7283,N_7163);
xor U7615 (N_7615,N_7299,N_7294);
xnor U7616 (N_7616,N_7028,N_7287);
or U7617 (N_7617,N_7239,N_7316);
nand U7618 (N_7618,N_7142,N_7183);
nand U7619 (N_7619,N_7091,N_7372);
nand U7620 (N_7620,N_7087,N_7325);
nor U7621 (N_7621,N_7162,N_7278);
and U7622 (N_7622,N_7240,N_7290);
xor U7623 (N_7623,N_7107,N_7013);
and U7624 (N_7624,N_7306,N_7424);
nand U7625 (N_7625,N_7149,N_7346);
nor U7626 (N_7626,N_7229,N_7352);
and U7627 (N_7627,N_7409,N_7214);
xnor U7628 (N_7628,N_7365,N_7065);
and U7629 (N_7629,N_7342,N_7011);
or U7630 (N_7630,N_7456,N_7108);
nand U7631 (N_7631,N_7103,N_7390);
and U7632 (N_7632,N_7207,N_7193);
and U7633 (N_7633,N_7477,N_7192);
and U7634 (N_7634,N_7480,N_7110);
or U7635 (N_7635,N_7332,N_7418);
nor U7636 (N_7636,N_7257,N_7196);
xnor U7637 (N_7637,N_7463,N_7258);
or U7638 (N_7638,N_7399,N_7120);
or U7639 (N_7639,N_7440,N_7448);
or U7640 (N_7640,N_7174,N_7050);
xor U7641 (N_7641,N_7208,N_7221);
nor U7642 (N_7642,N_7182,N_7429);
nor U7643 (N_7643,N_7152,N_7053);
xor U7644 (N_7644,N_7250,N_7321);
nand U7645 (N_7645,N_7260,N_7106);
nor U7646 (N_7646,N_7128,N_7441);
nand U7647 (N_7647,N_7002,N_7016);
nor U7648 (N_7648,N_7171,N_7275);
and U7649 (N_7649,N_7085,N_7455);
and U7650 (N_7650,N_7386,N_7124);
nor U7651 (N_7651,N_7450,N_7253);
nand U7652 (N_7652,N_7454,N_7465);
nor U7653 (N_7653,N_7206,N_7094);
nor U7654 (N_7654,N_7497,N_7069);
and U7655 (N_7655,N_7201,N_7328);
nor U7656 (N_7656,N_7394,N_7427);
and U7657 (N_7657,N_7140,N_7213);
xnor U7658 (N_7658,N_7317,N_7083);
or U7659 (N_7659,N_7024,N_7307);
xnor U7660 (N_7660,N_7068,N_7007);
xor U7661 (N_7661,N_7202,N_7043);
nor U7662 (N_7662,N_7396,N_7323);
nor U7663 (N_7663,N_7288,N_7018);
and U7664 (N_7664,N_7366,N_7392);
xor U7665 (N_7665,N_7145,N_7088);
or U7666 (N_7666,N_7225,N_7035);
nand U7667 (N_7667,N_7022,N_7266);
nand U7668 (N_7668,N_7359,N_7105);
nor U7669 (N_7669,N_7322,N_7169);
xor U7670 (N_7670,N_7382,N_7428);
or U7671 (N_7671,N_7473,N_7230);
nor U7672 (N_7672,N_7220,N_7006);
nand U7673 (N_7673,N_7129,N_7305);
nor U7674 (N_7674,N_7217,N_7296);
or U7675 (N_7675,N_7295,N_7425);
nand U7676 (N_7676,N_7356,N_7037);
nand U7677 (N_7677,N_7080,N_7179);
xor U7678 (N_7678,N_7354,N_7136);
nor U7679 (N_7679,N_7340,N_7181);
and U7680 (N_7680,N_7133,N_7277);
nor U7681 (N_7681,N_7150,N_7291);
and U7682 (N_7682,N_7070,N_7223);
and U7683 (N_7683,N_7270,N_7318);
nand U7684 (N_7684,N_7211,N_7387);
nand U7685 (N_7685,N_7269,N_7411);
nor U7686 (N_7686,N_7438,N_7155);
and U7687 (N_7687,N_7460,N_7159);
or U7688 (N_7688,N_7242,N_7339);
nor U7689 (N_7689,N_7101,N_7082);
xor U7690 (N_7690,N_7376,N_7326);
or U7691 (N_7691,N_7489,N_7186);
and U7692 (N_7692,N_7200,N_7459);
nor U7693 (N_7693,N_7042,N_7132);
and U7694 (N_7694,N_7243,N_7263);
xor U7695 (N_7695,N_7458,N_7116);
xnor U7696 (N_7696,N_7246,N_7338);
nor U7697 (N_7697,N_7044,N_7344);
nand U7698 (N_7698,N_7284,N_7276);
and U7699 (N_7699,N_7300,N_7442);
and U7700 (N_7700,N_7188,N_7413);
xor U7701 (N_7701,N_7143,N_7397);
nor U7702 (N_7702,N_7032,N_7054);
nand U7703 (N_7703,N_7137,N_7248);
nand U7704 (N_7704,N_7218,N_7475);
or U7705 (N_7705,N_7000,N_7123);
xor U7706 (N_7706,N_7420,N_7167);
or U7707 (N_7707,N_7469,N_7048);
nor U7708 (N_7708,N_7114,N_7446);
nor U7709 (N_7709,N_7251,N_7482);
nand U7710 (N_7710,N_7098,N_7233);
and U7711 (N_7711,N_7353,N_7219);
nor U7712 (N_7712,N_7184,N_7113);
and U7713 (N_7713,N_7329,N_7104);
and U7714 (N_7714,N_7280,N_7485);
or U7715 (N_7715,N_7309,N_7443);
or U7716 (N_7716,N_7388,N_7432);
xnor U7717 (N_7717,N_7487,N_7245);
or U7718 (N_7718,N_7001,N_7470);
xnor U7719 (N_7719,N_7212,N_7148);
and U7720 (N_7720,N_7404,N_7146);
xor U7721 (N_7721,N_7478,N_7292);
or U7722 (N_7722,N_7067,N_7135);
and U7723 (N_7723,N_7431,N_7190);
xor U7724 (N_7724,N_7147,N_7445);
nand U7725 (N_7725,N_7389,N_7215);
nor U7726 (N_7726,N_7055,N_7279);
or U7727 (N_7727,N_7071,N_7265);
or U7728 (N_7728,N_7194,N_7407);
nor U7729 (N_7729,N_7072,N_7172);
nor U7730 (N_7730,N_7343,N_7320);
xor U7731 (N_7731,N_7131,N_7021);
xnor U7732 (N_7732,N_7301,N_7496);
nand U7733 (N_7733,N_7034,N_7383);
nor U7734 (N_7734,N_7118,N_7134);
nor U7735 (N_7735,N_7302,N_7479);
nand U7736 (N_7736,N_7041,N_7046);
and U7737 (N_7737,N_7189,N_7286);
xnor U7738 (N_7738,N_7380,N_7247);
or U7739 (N_7739,N_7341,N_7165);
and U7740 (N_7740,N_7377,N_7436);
nor U7741 (N_7741,N_7074,N_7238);
and U7742 (N_7742,N_7017,N_7476);
nor U7743 (N_7743,N_7408,N_7472);
nand U7744 (N_7744,N_7333,N_7232);
and U7745 (N_7745,N_7073,N_7348);
xnor U7746 (N_7746,N_7484,N_7119);
nand U7747 (N_7747,N_7111,N_7023);
nand U7748 (N_7748,N_7385,N_7177);
nor U7749 (N_7749,N_7198,N_7345);
nor U7750 (N_7750,N_7064,N_7160);
nand U7751 (N_7751,N_7111,N_7443);
xnor U7752 (N_7752,N_7027,N_7310);
or U7753 (N_7753,N_7045,N_7182);
nor U7754 (N_7754,N_7024,N_7233);
and U7755 (N_7755,N_7293,N_7139);
or U7756 (N_7756,N_7188,N_7258);
and U7757 (N_7757,N_7390,N_7024);
xor U7758 (N_7758,N_7047,N_7058);
nor U7759 (N_7759,N_7181,N_7227);
or U7760 (N_7760,N_7191,N_7064);
xor U7761 (N_7761,N_7376,N_7082);
and U7762 (N_7762,N_7337,N_7125);
nor U7763 (N_7763,N_7349,N_7152);
or U7764 (N_7764,N_7274,N_7107);
and U7765 (N_7765,N_7172,N_7339);
xnor U7766 (N_7766,N_7207,N_7192);
nand U7767 (N_7767,N_7426,N_7370);
xor U7768 (N_7768,N_7445,N_7211);
xnor U7769 (N_7769,N_7212,N_7256);
and U7770 (N_7770,N_7108,N_7000);
xnor U7771 (N_7771,N_7257,N_7118);
or U7772 (N_7772,N_7343,N_7234);
nor U7773 (N_7773,N_7338,N_7039);
nand U7774 (N_7774,N_7155,N_7493);
nand U7775 (N_7775,N_7026,N_7199);
nand U7776 (N_7776,N_7471,N_7485);
or U7777 (N_7777,N_7244,N_7209);
nor U7778 (N_7778,N_7323,N_7148);
or U7779 (N_7779,N_7475,N_7462);
nand U7780 (N_7780,N_7061,N_7495);
nor U7781 (N_7781,N_7448,N_7482);
xor U7782 (N_7782,N_7053,N_7242);
nor U7783 (N_7783,N_7093,N_7013);
xor U7784 (N_7784,N_7354,N_7245);
nor U7785 (N_7785,N_7039,N_7398);
or U7786 (N_7786,N_7195,N_7214);
and U7787 (N_7787,N_7153,N_7281);
and U7788 (N_7788,N_7016,N_7383);
or U7789 (N_7789,N_7084,N_7427);
nand U7790 (N_7790,N_7494,N_7381);
and U7791 (N_7791,N_7313,N_7298);
nor U7792 (N_7792,N_7393,N_7404);
and U7793 (N_7793,N_7458,N_7279);
and U7794 (N_7794,N_7374,N_7485);
xnor U7795 (N_7795,N_7336,N_7085);
xor U7796 (N_7796,N_7140,N_7357);
nand U7797 (N_7797,N_7332,N_7239);
or U7798 (N_7798,N_7306,N_7418);
nand U7799 (N_7799,N_7266,N_7463);
nand U7800 (N_7800,N_7113,N_7024);
nor U7801 (N_7801,N_7103,N_7431);
nand U7802 (N_7802,N_7365,N_7072);
or U7803 (N_7803,N_7097,N_7286);
nor U7804 (N_7804,N_7465,N_7430);
and U7805 (N_7805,N_7310,N_7409);
xnor U7806 (N_7806,N_7308,N_7387);
and U7807 (N_7807,N_7174,N_7181);
nor U7808 (N_7808,N_7493,N_7174);
nor U7809 (N_7809,N_7414,N_7218);
xnor U7810 (N_7810,N_7295,N_7102);
xor U7811 (N_7811,N_7343,N_7499);
and U7812 (N_7812,N_7062,N_7049);
and U7813 (N_7813,N_7039,N_7439);
or U7814 (N_7814,N_7151,N_7304);
and U7815 (N_7815,N_7130,N_7354);
nand U7816 (N_7816,N_7063,N_7222);
and U7817 (N_7817,N_7349,N_7121);
nor U7818 (N_7818,N_7468,N_7251);
or U7819 (N_7819,N_7499,N_7069);
nor U7820 (N_7820,N_7258,N_7424);
nand U7821 (N_7821,N_7402,N_7150);
and U7822 (N_7822,N_7083,N_7465);
nor U7823 (N_7823,N_7399,N_7172);
or U7824 (N_7824,N_7159,N_7314);
and U7825 (N_7825,N_7495,N_7167);
xnor U7826 (N_7826,N_7077,N_7449);
or U7827 (N_7827,N_7310,N_7084);
and U7828 (N_7828,N_7331,N_7079);
xnor U7829 (N_7829,N_7313,N_7282);
nand U7830 (N_7830,N_7155,N_7282);
xnor U7831 (N_7831,N_7352,N_7217);
nor U7832 (N_7832,N_7155,N_7027);
and U7833 (N_7833,N_7331,N_7392);
nor U7834 (N_7834,N_7235,N_7288);
nor U7835 (N_7835,N_7201,N_7144);
nand U7836 (N_7836,N_7201,N_7441);
xnor U7837 (N_7837,N_7058,N_7037);
nand U7838 (N_7838,N_7489,N_7416);
nand U7839 (N_7839,N_7392,N_7166);
xnor U7840 (N_7840,N_7221,N_7244);
or U7841 (N_7841,N_7206,N_7124);
and U7842 (N_7842,N_7239,N_7279);
nand U7843 (N_7843,N_7196,N_7428);
nand U7844 (N_7844,N_7497,N_7021);
and U7845 (N_7845,N_7388,N_7093);
or U7846 (N_7846,N_7196,N_7068);
and U7847 (N_7847,N_7408,N_7318);
and U7848 (N_7848,N_7321,N_7426);
nand U7849 (N_7849,N_7261,N_7061);
and U7850 (N_7850,N_7475,N_7437);
nand U7851 (N_7851,N_7215,N_7388);
nor U7852 (N_7852,N_7261,N_7478);
nand U7853 (N_7853,N_7321,N_7109);
xnor U7854 (N_7854,N_7239,N_7317);
nand U7855 (N_7855,N_7108,N_7360);
nor U7856 (N_7856,N_7099,N_7196);
and U7857 (N_7857,N_7196,N_7147);
and U7858 (N_7858,N_7337,N_7241);
or U7859 (N_7859,N_7223,N_7108);
nand U7860 (N_7860,N_7018,N_7177);
and U7861 (N_7861,N_7209,N_7204);
and U7862 (N_7862,N_7033,N_7372);
or U7863 (N_7863,N_7272,N_7072);
or U7864 (N_7864,N_7452,N_7352);
xnor U7865 (N_7865,N_7180,N_7224);
and U7866 (N_7866,N_7393,N_7407);
nor U7867 (N_7867,N_7164,N_7312);
nor U7868 (N_7868,N_7044,N_7299);
xor U7869 (N_7869,N_7469,N_7017);
and U7870 (N_7870,N_7465,N_7358);
or U7871 (N_7871,N_7384,N_7371);
xor U7872 (N_7872,N_7175,N_7320);
or U7873 (N_7873,N_7312,N_7070);
nand U7874 (N_7874,N_7487,N_7395);
nand U7875 (N_7875,N_7347,N_7378);
nand U7876 (N_7876,N_7244,N_7329);
or U7877 (N_7877,N_7210,N_7019);
nor U7878 (N_7878,N_7278,N_7262);
and U7879 (N_7879,N_7387,N_7370);
nand U7880 (N_7880,N_7276,N_7192);
and U7881 (N_7881,N_7253,N_7305);
nand U7882 (N_7882,N_7179,N_7104);
nor U7883 (N_7883,N_7437,N_7290);
or U7884 (N_7884,N_7463,N_7220);
nor U7885 (N_7885,N_7315,N_7239);
nand U7886 (N_7886,N_7409,N_7171);
and U7887 (N_7887,N_7408,N_7399);
nor U7888 (N_7888,N_7246,N_7462);
and U7889 (N_7889,N_7427,N_7224);
xor U7890 (N_7890,N_7010,N_7068);
or U7891 (N_7891,N_7446,N_7162);
nor U7892 (N_7892,N_7072,N_7097);
nor U7893 (N_7893,N_7048,N_7392);
or U7894 (N_7894,N_7097,N_7357);
xnor U7895 (N_7895,N_7394,N_7236);
nor U7896 (N_7896,N_7308,N_7301);
nor U7897 (N_7897,N_7437,N_7199);
nand U7898 (N_7898,N_7023,N_7154);
nand U7899 (N_7899,N_7139,N_7269);
xor U7900 (N_7900,N_7224,N_7378);
nand U7901 (N_7901,N_7492,N_7190);
or U7902 (N_7902,N_7354,N_7440);
or U7903 (N_7903,N_7068,N_7344);
xor U7904 (N_7904,N_7235,N_7068);
or U7905 (N_7905,N_7093,N_7254);
or U7906 (N_7906,N_7481,N_7083);
xor U7907 (N_7907,N_7054,N_7179);
nor U7908 (N_7908,N_7002,N_7018);
or U7909 (N_7909,N_7101,N_7038);
nor U7910 (N_7910,N_7478,N_7029);
or U7911 (N_7911,N_7176,N_7057);
and U7912 (N_7912,N_7139,N_7206);
xor U7913 (N_7913,N_7072,N_7445);
and U7914 (N_7914,N_7136,N_7067);
and U7915 (N_7915,N_7413,N_7165);
or U7916 (N_7916,N_7216,N_7453);
or U7917 (N_7917,N_7262,N_7454);
xnor U7918 (N_7918,N_7341,N_7145);
or U7919 (N_7919,N_7219,N_7455);
nand U7920 (N_7920,N_7273,N_7248);
nor U7921 (N_7921,N_7435,N_7125);
xnor U7922 (N_7922,N_7407,N_7316);
and U7923 (N_7923,N_7153,N_7289);
nor U7924 (N_7924,N_7098,N_7156);
and U7925 (N_7925,N_7133,N_7203);
nand U7926 (N_7926,N_7184,N_7084);
xor U7927 (N_7927,N_7003,N_7398);
nor U7928 (N_7928,N_7445,N_7313);
and U7929 (N_7929,N_7471,N_7468);
or U7930 (N_7930,N_7214,N_7359);
nand U7931 (N_7931,N_7090,N_7350);
or U7932 (N_7932,N_7498,N_7018);
xnor U7933 (N_7933,N_7195,N_7072);
or U7934 (N_7934,N_7286,N_7073);
and U7935 (N_7935,N_7237,N_7459);
or U7936 (N_7936,N_7069,N_7410);
xnor U7937 (N_7937,N_7258,N_7233);
or U7938 (N_7938,N_7124,N_7324);
or U7939 (N_7939,N_7117,N_7026);
nand U7940 (N_7940,N_7323,N_7494);
nand U7941 (N_7941,N_7406,N_7387);
xor U7942 (N_7942,N_7490,N_7447);
or U7943 (N_7943,N_7349,N_7386);
nor U7944 (N_7944,N_7149,N_7284);
and U7945 (N_7945,N_7302,N_7118);
xor U7946 (N_7946,N_7399,N_7089);
and U7947 (N_7947,N_7160,N_7425);
and U7948 (N_7948,N_7377,N_7461);
xnor U7949 (N_7949,N_7270,N_7020);
nor U7950 (N_7950,N_7023,N_7247);
nand U7951 (N_7951,N_7145,N_7289);
xnor U7952 (N_7952,N_7049,N_7104);
and U7953 (N_7953,N_7029,N_7184);
nand U7954 (N_7954,N_7393,N_7221);
and U7955 (N_7955,N_7200,N_7033);
nand U7956 (N_7956,N_7142,N_7368);
or U7957 (N_7957,N_7407,N_7327);
nor U7958 (N_7958,N_7193,N_7151);
and U7959 (N_7959,N_7111,N_7326);
xnor U7960 (N_7960,N_7128,N_7220);
nand U7961 (N_7961,N_7411,N_7299);
and U7962 (N_7962,N_7417,N_7376);
and U7963 (N_7963,N_7398,N_7411);
or U7964 (N_7964,N_7464,N_7061);
nor U7965 (N_7965,N_7285,N_7171);
nor U7966 (N_7966,N_7156,N_7028);
or U7967 (N_7967,N_7215,N_7099);
or U7968 (N_7968,N_7414,N_7407);
or U7969 (N_7969,N_7397,N_7427);
or U7970 (N_7970,N_7085,N_7273);
xor U7971 (N_7971,N_7347,N_7414);
or U7972 (N_7972,N_7326,N_7374);
nor U7973 (N_7973,N_7428,N_7236);
xnor U7974 (N_7974,N_7393,N_7347);
or U7975 (N_7975,N_7395,N_7446);
nand U7976 (N_7976,N_7402,N_7254);
or U7977 (N_7977,N_7478,N_7285);
xor U7978 (N_7978,N_7164,N_7296);
or U7979 (N_7979,N_7407,N_7217);
xor U7980 (N_7980,N_7478,N_7098);
or U7981 (N_7981,N_7164,N_7210);
nand U7982 (N_7982,N_7183,N_7189);
and U7983 (N_7983,N_7434,N_7254);
xor U7984 (N_7984,N_7105,N_7014);
and U7985 (N_7985,N_7296,N_7485);
and U7986 (N_7986,N_7095,N_7310);
nor U7987 (N_7987,N_7353,N_7252);
nor U7988 (N_7988,N_7404,N_7353);
nand U7989 (N_7989,N_7325,N_7211);
xnor U7990 (N_7990,N_7146,N_7431);
xor U7991 (N_7991,N_7288,N_7029);
and U7992 (N_7992,N_7218,N_7353);
nand U7993 (N_7993,N_7008,N_7086);
and U7994 (N_7994,N_7280,N_7359);
and U7995 (N_7995,N_7467,N_7172);
nand U7996 (N_7996,N_7368,N_7173);
nor U7997 (N_7997,N_7224,N_7164);
and U7998 (N_7998,N_7063,N_7450);
nand U7999 (N_7999,N_7004,N_7181);
or U8000 (N_8000,N_7533,N_7871);
and U8001 (N_8001,N_7641,N_7991);
and U8002 (N_8002,N_7684,N_7626);
xnor U8003 (N_8003,N_7678,N_7951);
nor U8004 (N_8004,N_7529,N_7781);
xnor U8005 (N_8005,N_7961,N_7592);
nand U8006 (N_8006,N_7547,N_7527);
and U8007 (N_8007,N_7865,N_7915);
nor U8008 (N_8008,N_7728,N_7758);
and U8009 (N_8009,N_7739,N_7817);
nor U8010 (N_8010,N_7856,N_7808);
nor U8011 (N_8011,N_7889,N_7909);
xor U8012 (N_8012,N_7891,N_7937);
or U8013 (N_8013,N_7510,N_7730);
nor U8014 (N_8014,N_7798,N_7890);
nand U8015 (N_8015,N_7610,N_7561);
nand U8016 (N_8016,N_7884,N_7872);
and U8017 (N_8017,N_7582,N_7974);
nor U8018 (N_8018,N_7503,N_7964);
and U8019 (N_8019,N_7908,N_7605);
nor U8020 (N_8020,N_7709,N_7824);
xnor U8021 (N_8021,N_7819,N_7789);
or U8022 (N_8022,N_7899,N_7942);
xnor U8023 (N_8023,N_7633,N_7785);
or U8024 (N_8024,N_7548,N_7946);
xor U8025 (N_8025,N_7864,N_7837);
and U8026 (N_8026,N_7540,N_7744);
nor U8027 (N_8027,N_7532,N_7702);
nor U8028 (N_8028,N_7528,N_7805);
nor U8029 (N_8029,N_7591,N_7848);
or U8030 (N_8030,N_7828,N_7793);
nor U8031 (N_8031,N_7830,N_7885);
nand U8032 (N_8032,N_7981,N_7893);
nor U8033 (N_8033,N_7657,N_7556);
xnor U8034 (N_8034,N_7635,N_7672);
nor U8035 (N_8035,N_7854,N_7863);
nand U8036 (N_8036,N_7840,N_7998);
xor U8037 (N_8037,N_7970,N_7571);
nor U8038 (N_8038,N_7751,N_7955);
xor U8039 (N_8039,N_7827,N_7584);
or U8040 (N_8040,N_7897,N_7983);
nand U8041 (N_8041,N_7901,N_7555);
nor U8042 (N_8042,N_7590,N_7883);
and U8043 (N_8043,N_7844,N_7554);
or U8044 (N_8044,N_7777,N_7741);
xnor U8045 (N_8045,N_7644,N_7782);
xor U8046 (N_8046,N_7965,N_7846);
nand U8047 (N_8047,N_7809,N_7940);
nand U8048 (N_8048,N_7604,N_7987);
nand U8049 (N_8049,N_7718,N_7770);
nand U8050 (N_8050,N_7935,N_7640);
and U8051 (N_8051,N_7620,N_7919);
or U8052 (N_8052,N_7853,N_7646);
nand U8053 (N_8053,N_7986,N_7866);
xnor U8054 (N_8054,N_7515,N_7643);
nor U8055 (N_8055,N_7995,N_7594);
or U8056 (N_8056,N_7621,N_7984);
or U8057 (N_8057,N_7512,N_7707);
or U8058 (N_8058,N_7930,N_7760);
nand U8059 (N_8059,N_7616,N_7795);
or U8060 (N_8060,N_7943,N_7553);
nor U8061 (N_8061,N_7904,N_7888);
or U8062 (N_8062,N_7818,N_7886);
and U8063 (N_8063,N_7780,N_7736);
nand U8064 (N_8064,N_7535,N_7916);
nor U8065 (N_8065,N_7806,N_7507);
nor U8066 (N_8066,N_7947,N_7650);
nand U8067 (N_8067,N_7653,N_7634);
or U8068 (N_8068,N_7563,N_7585);
nor U8069 (N_8069,N_7724,N_7740);
or U8070 (N_8070,N_7629,N_7520);
nand U8071 (N_8071,N_7598,N_7755);
or U8072 (N_8072,N_7979,N_7878);
and U8073 (N_8073,N_7654,N_7903);
nor U8074 (N_8074,N_7945,N_7989);
xor U8075 (N_8075,N_7656,N_7544);
nor U8076 (N_8076,N_7642,N_7698);
or U8077 (N_8077,N_7917,N_7799);
and U8078 (N_8078,N_7825,N_7958);
nor U8079 (N_8079,N_7664,N_7896);
and U8080 (N_8080,N_7934,N_7669);
or U8081 (N_8081,N_7722,N_7692);
nand U8082 (N_8082,N_7800,N_7745);
nor U8083 (N_8083,N_7677,N_7802);
and U8084 (N_8084,N_7767,N_7721);
nand U8085 (N_8085,N_7577,N_7578);
xor U8086 (N_8086,N_7710,N_7674);
nor U8087 (N_8087,N_7737,N_7505);
nand U8088 (N_8088,N_7881,N_7708);
or U8089 (N_8089,N_7949,N_7861);
xnor U8090 (N_8090,N_7757,N_7575);
nor U8091 (N_8091,N_7720,N_7699);
xor U8092 (N_8092,N_7822,N_7504);
nand U8093 (N_8093,N_7959,N_7637);
and U8094 (N_8094,N_7842,N_7953);
or U8095 (N_8095,N_7833,N_7717);
and U8096 (N_8096,N_7841,N_7936);
nor U8097 (N_8097,N_7774,N_7960);
nor U8098 (N_8098,N_7660,N_7676);
xnor U8099 (N_8099,N_7876,N_7541);
and U8100 (N_8100,N_7615,N_7996);
nor U8101 (N_8101,N_7764,N_7509);
nor U8102 (N_8102,N_7600,N_7791);
or U8103 (N_8103,N_7801,N_7521);
or U8104 (N_8104,N_7688,N_7680);
or U8105 (N_8105,N_7753,N_7735);
and U8106 (N_8106,N_7549,N_7689);
nor U8107 (N_8107,N_7531,N_7769);
and U8108 (N_8108,N_7611,N_7667);
xnor U8109 (N_8109,N_7994,N_7948);
xnor U8110 (N_8110,N_7734,N_7898);
nor U8111 (N_8111,N_7771,N_7567);
xnor U8112 (N_8112,N_7502,N_7762);
nand U8113 (N_8113,N_7829,N_7999);
nor U8114 (N_8114,N_7892,N_7514);
or U8115 (N_8115,N_7839,N_7652);
xor U8116 (N_8116,N_7713,N_7993);
nor U8117 (N_8117,N_7847,N_7906);
nor U8118 (N_8118,N_7895,N_7559);
and U8119 (N_8119,N_7912,N_7733);
xor U8120 (N_8120,N_7976,N_7648);
nand U8121 (N_8121,N_7666,N_7815);
and U8122 (N_8122,N_7665,N_7685);
nor U8123 (N_8123,N_7977,N_7978);
or U8124 (N_8124,N_7647,N_7662);
nor U8125 (N_8125,N_7682,N_7944);
xnor U8126 (N_8126,N_7796,N_7696);
and U8127 (N_8127,N_7523,N_7923);
nor U8128 (N_8128,N_7941,N_7982);
nor U8129 (N_8129,N_7614,N_7867);
nor U8130 (N_8130,N_7560,N_7612);
xnor U8131 (N_8131,N_7712,N_7673);
nand U8132 (N_8132,N_7985,N_7968);
xnor U8133 (N_8133,N_7910,N_7859);
nand U8134 (N_8134,N_7572,N_7623);
and U8135 (N_8135,N_7562,N_7950);
and U8136 (N_8136,N_7875,N_7715);
and U8137 (N_8137,N_7566,N_7599);
or U8138 (N_8138,N_7538,N_7814);
or U8139 (N_8139,N_7636,N_7628);
and U8140 (N_8140,N_7705,N_7659);
or U8141 (N_8141,N_7790,N_7877);
and U8142 (N_8142,N_7693,N_7850);
or U8143 (N_8143,N_7526,N_7775);
nand U8144 (N_8144,N_7823,N_7619);
nor U8145 (N_8145,N_7803,N_7668);
and U8146 (N_8146,N_7932,N_7826);
nor U8147 (N_8147,N_7794,N_7606);
nand U8148 (N_8148,N_7922,N_7601);
nor U8149 (N_8149,N_7732,N_7670);
or U8150 (N_8150,N_7820,N_7773);
nor U8151 (N_8151,N_7701,N_7638);
or U8152 (N_8152,N_7810,N_7962);
or U8153 (N_8153,N_7975,N_7914);
nor U8154 (N_8154,N_7807,N_7513);
nor U8155 (N_8155,N_7738,N_7849);
xnor U8156 (N_8156,N_7966,N_7990);
and U8157 (N_8157,N_7797,N_7542);
xor U8158 (N_8158,N_7843,N_7992);
or U8159 (N_8159,N_7725,N_7918);
and U8160 (N_8160,N_7776,N_7957);
xor U8161 (N_8161,N_7783,N_7519);
or U8162 (N_8162,N_7727,N_7649);
xnor U8163 (N_8163,N_7772,N_7729);
nand U8164 (N_8164,N_7907,N_7855);
or U8165 (N_8165,N_7954,N_7516);
or U8166 (N_8166,N_7586,N_7655);
nand U8167 (N_8167,N_7500,N_7813);
xor U8168 (N_8168,N_7763,N_7779);
or U8169 (N_8169,N_7857,N_7576);
and U8170 (N_8170,N_7851,N_7997);
nand U8171 (N_8171,N_7622,N_7645);
xor U8172 (N_8172,N_7778,N_7617);
and U8173 (N_8173,N_7931,N_7754);
or U8174 (N_8174,N_7874,N_7714);
xnor U8175 (N_8175,N_7536,N_7697);
and U8176 (N_8176,N_7927,N_7834);
xor U8177 (N_8177,N_7905,N_7746);
and U8178 (N_8178,N_7700,N_7980);
or U8179 (N_8179,N_7587,N_7681);
nand U8180 (N_8180,N_7821,N_7880);
nand U8181 (N_8181,N_7765,N_7835);
or U8182 (N_8182,N_7518,N_7706);
or U8183 (N_8183,N_7671,N_7630);
or U8184 (N_8184,N_7902,N_7747);
or U8185 (N_8185,N_7752,N_7804);
or U8186 (N_8186,N_7860,N_7879);
nand U8187 (N_8187,N_7926,N_7564);
xnor U8188 (N_8188,N_7675,N_7691);
or U8189 (N_8189,N_7686,N_7557);
nor U8190 (N_8190,N_7552,N_7952);
xnor U8191 (N_8191,N_7894,N_7723);
nand U8192 (N_8192,N_7704,N_7925);
and U8193 (N_8193,N_7683,N_7661);
and U8194 (N_8194,N_7836,N_7695);
xor U8195 (N_8195,N_7690,N_7595);
xor U8196 (N_8196,N_7759,N_7933);
and U8197 (N_8197,N_7593,N_7534);
xnor U8198 (N_8198,N_7969,N_7967);
or U8199 (N_8199,N_7973,N_7570);
xnor U8200 (N_8200,N_7726,N_7938);
nor U8201 (N_8201,N_7569,N_7506);
nand U8202 (N_8202,N_7583,N_7613);
xnor U8203 (N_8203,N_7786,N_7963);
nor U8204 (N_8204,N_7568,N_7525);
nand U8205 (N_8205,N_7766,N_7742);
and U8206 (N_8206,N_7588,N_7545);
nand U8207 (N_8207,N_7511,N_7580);
or U8208 (N_8208,N_7920,N_7921);
and U8209 (N_8209,N_7868,N_7731);
or U8210 (N_8210,N_7719,N_7663);
or U8211 (N_8211,N_7750,N_7543);
nand U8212 (N_8212,N_7618,N_7603);
nor U8213 (N_8213,N_7988,N_7956);
xor U8214 (N_8214,N_7573,N_7972);
or U8215 (N_8215,N_7609,N_7761);
xor U8216 (N_8216,N_7679,N_7749);
or U8217 (N_8217,N_7625,N_7558);
and U8218 (N_8218,N_7551,N_7651);
or U8219 (N_8219,N_7768,N_7784);
and U8220 (N_8220,N_7900,N_7711);
or U8221 (N_8221,N_7748,N_7631);
nor U8222 (N_8222,N_7811,N_7522);
xnor U8223 (N_8223,N_7632,N_7703);
or U8224 (N_8224,N_7831,N_7694);
or U8225 (N_8225,N_7658,N_7607);
and U8226 (N_8226,N_7524,N_7845);
nor U8227 (N_8227,N_7939,N_7971);
nor U8228 (N_8228,N_7862,N_7537);
nor U8229 (N_8229,N_7581,N_7882);
and U8230 (N_8230,N_7508,N_7589);
nand U8231 (N_8231,N_7858,N_7602);
and U8232 (N_8232,N_7870,N_7743);
or U8233 (N_8233,N_7574,N_7913);
nand U8234 (N_8234,N_7687,N_7756);
nor U8235 (N_8235,N_7816,N_7788);
and U8236 (N_8236,N_7530,N_7539);
or U8237 (N_8237,N_7911,N_7624);
nor U8238 (N_8238,N_7565,N_7639);
nor U8239 (N_8239,N_7873,N_7550);
xor U8240 (N_8240,N_7924,N_7838);
and U8241 (N_8241,N_7787,N_7517);
nor U8242 (N_8242,N_7608,N_7887);
or U8243 (N_8243,N_7627,N_7928);
or U8244 (N_8244,N_7546,N_7596);
and U8245 (N_8245,N_7792,N_7929);
nand U8246 (N_8246,N_7812,N_7716);
and U8247 (N_8247,N_7852,N_7597);
or U8248 (N_8248,N_7832,N_7869);
xor U8249 (N_8249,N_7501,N_7579);
nand U8250 (N_8250,N_7966,N_7572);
nor U8251 (N_8251,N_7745,N_7614);
and U8252 (N_8252,N_7581,N_7526);
nor U8253 (N_8253,N_7743,N_7664);
nand U8254 (N_8254,N_7712,N_7736);
xor U8255 (N_8255,N_7942,N_7946);
nand U8256 (N_8256,N_7860,N_7753);
and U8257 (N_8257,N_7946,N_7748);
nor U8258 (N_8258,N_7890,N_7834);
or U8259 (N_8259,N_7722,N_7663);
and U8260 (N_8260,N_7608,N_7737);
nor U8261 (N_8261,N_7692,N_7585);
xnor U8262 (N_8262,N_7821,N_7751);
xor U8263 (N_8263,N_7792,N_7631);
and U8264 (N_8264,N_7796,N_7519);
and U8265 (N_8265,N_7950,N_7729);
or U8266 (N_8266,N_7602,N_7730);
and U8267 (N_8267,N_7957,N_7718);
or U8268 (N_8268,N_7554,N_7545);
nor U8269 (N_8269,N_7608,N_7931);
or U8270 (N_8270,N_7782,N_7908);
xnor U8271 (N_8271,N_7936,N_7938);
xor U8272 (N_8272,N_7793,N_7795);
nor U8273 (N_8273,N_7510,N_7585);
xor U8274 (N_8274,N_7666,N_7516);
nor U8275 (N_8275,N_7580,N_7513);
xnor U8276 (N_8276,N_7761,N_7804);
or U8277 (N_8277,N_7630,N_7806);
nand U8278 (N_8278,N_7652,N_7608);
nor U8279 (N_8279,N_7549,N_7916);
or U8280 (N_8280,N_7974,N_7601);
nand U8281 (N_8281,N_7610,N_7671);
nor U8282 (N_8282,N_7804,N_7572);
xnor U8283 (N_8283,N_7575,N_7504);
nor U8284 (N_8284,N_7810,N_7508);
nand U8285 (N_8285,N_7816,N_7852);
xnor U8286 (N_8286,N_7601,N_7773);
nand U8287 (N_8287,N_7870,N_7648);
xor U8288 (N_8288,N_7601,N_7536);
and U8289 (N_8289,N_7752,N_7906);
nor U8290 (N_8290,N_7542,N_7587);
or U8291 (N_8291,N_7980,N_7612);
nand U8292 (N_8292,N_7602,N_7639);
xnor U8293 (N_8293,N_7558,N_7520);
and U8294 (N_8294,N_7716,N_7578);
and U8295 (N_8295,N_7918,N_7737);
nand U8296 (N_8296,N_7723,N_7764);
nor U8297 (N_8297,N_7521,N_7913);
nor U8298 (N_8298,N_7700,N_7569);
or U8299 (N_8299,N_7682,N_7879);
or U8300 (N_8300,N_7863,N_7735);
nor U8301 (N_8301,N_7898,N_7730);
nor U8302 (N_8302,N_7961,N_7963);
nand U8303 (N_8303,N_7773,N_7939);
nor U8304 (N_8304,N_7948,N_7700);
nand U8305 (N_8305,N_7647,N_7880);
or U8306 (N_8306,N_7882,N_7930);
nand U8307 (N_8307,N_7500,N_7638);
nor U8308 (N_8308,N_7939,N_7564);
nor U8309 (N_8309,N_7620,N_7899);
and U8310 (N_8310,N_7812,N_7631);
nor U8311 (N_8311,N_7652,N_7611);
nand U8312 (N_8312,N_7682,N_7713);
or U8313 (N_8313,N_7849,N_7766);
or U8314 (N_8314,N_7567,N_7643);
nand U8315 (N_8315,N_7941,N_7647);
nor U8316 (N_8316,N_7950,N_7829);
or U8317 (N_8317,N_7551,N_7623);
xor U8318 (N_8318,N_7947,N_7504);
or U8319 (N_8319,N_7653,N_7710);
nand U8320 (N_8320,N_7963,N_7992);
xor U8321 (N_8321,N_7874,N_7643);
and U8322 (N_8322,N_7911,N_7666);
and U8323 (N_8323,N_7873,N_7783);
nand U8324 (N_8324,N_7549,N_7706);
nor U8325 (N_8325,N_7672,N_7627);
or U8326 (N_8326,N_7844,N_7762);
and U8327 (N_8327,N_7890,N_7905);
nor U8328 (N_8328,N_7820,N_7530);
nor U8329 (N_8329,N_7954,N_7850);
nand U8330 (N_8330,N_7714,N_7620);
nor U8331 (N_8331,N_7747,N_7833);
nand U8332 (N_8332,N_7621,N_7552);
or U8333 (N_8333,N_7676,N_7932);
nor U8334 (N_8334,N_7986,N_7560);
nand U8335 (N_8335,N_7955,N_7956);
nand U8336 (N_8336,N_7924,N_7750);
and U8337 (N_8337,N_7867,N_7593);
xor U8338 (N_8338,N_7969,N_7958);
nor U8339 (N_8339,N_7573,N_7867);
nand U8340 (N_8340,N_7560,N_7617);
nand U8341 (N_8341,N_7868,N_7665);
xnor U8342 (N_8342,N_7953,N_7966);
or U8343 (N_8343,N_7694,N_7832);
nand U8344 (N_8344,N_7658,N_7641);
nor U8345 (N_8345,N_7647,N_7899);
xnor U8346 (N_8346,N_7740,N_7748);
nor U8347 (N_8347,N_7507,N_7926);
nand U8348 (N_8348,N_7667,N_7649);
and U8349 (N_8349,N_7651,N_7681);
and U8350 (N_8350,N_7813,N_7894);
xor U8351 (N_8351,N_7674,N_7576);
and U8352 (N_8352,N_7895,N_7977);
or U8353 (N_8353,N_7873,N_7506);
and U8354 (N_8354,N_7781,N_7847);
and U8355 (N_8355,N_7710,N_7546);
xor U8356 (N_8356,N_7918,N_7562);
and U8357 (N_8357,N_7555,N_7897);
xor U8358 (N_8358,N_7874,N_7914);
nor U8359 (N_8359,N_7998,N_7649);
nor U8360 (N_8360,N_7582,N_7961);
xor U8361 (N_8361,N_7631,N_7949);
nor U8362 (N_8362,N_7610,N_7755);
xnor U8363 (N_8363,N_7563,N_7646);
and U8364 (N_8364,N_7903,N_7772);
xor U8365 (N_8365,N_7931,N_7559);
xnor U8366 (N_8366,N_7694,N_7797);
xor U8367 (N_8367,N_7712,N_7665);
nand U8368 (N_8368,N_7993,N_7509);
xnor U8369 (N_8369,N_7997,N_7934);
xor U8370 (N_8370,N_7699,N_7709);
nand U8371 (N_8371,N_7761,N_7798);
nor U8372 (N_8372,N_7931,N_7766);
and U8373 (N_8373,N_7900,N_7811);
or U8374 (N_8374,N_7983,N_7720);
or U8375 (N_8375,N_7746,N_7725);
nor U8376 (N_8376,N_7778,N_7579);
nor U8377 (N_8377,N_7506,N_7604);
or U8378 (N_8378,N_7651,N_7925);
and U8379 (N_8379,N_7925,N_7674);
or U8380 (N_8380,N_7513,N_7572);
and U8381 (N_8381,N_7847,N_7628);
or U8382 (N_8382,N_7658,N_7614);
nand U8383 (N_8383,N_7775,N_7896);
nor U8384 (N_8384,N_7972,N_7890);
or U8385 (N_8385,N_7559,N_7800);
nand U8386 (N_8386,N_7739,N_7628);
nand U8387 (N_8387,N_7638,N_7611);
and U8388 (N_8388,N_7542,N_7586);
xnor U8389 (N_8389,N_7877,N_7661);
nand U8390 (N_8390,N_7540,N_7857);
or U8391 (N_8391,N_7956,N_7529);
or U8392 (N_8392,N_7734,N_7871);
nor U8393 (N_8393,N_7528,N_7851);
or U8394 (N_8394,N_7963,N_7551);
nor U8395 (N_8395,N_7887,N_7536);
nor U8396 (N_8396,N_7705,N_7773);
nor U8397 (N_8397,N_7675,N_7856);
nand U8398 (N_8398,N_7950,N_7551);
or U8399 (N_8399,N_7788,N_7560);
and U8400 (N_8400,N_7879,N_7788);
nor U8401 (N_8401,N_7691,N_7683);
or U8402 (N_8402,N_7633,N_7964);
nor U8403 (N_8403,N_7769,N_7577);
xnor U8404 (N_8404,N_7879,N_7671);
xor U8405 (N_8405,N_7955,N_7738);
nand U8406 (N_8406,N_7718,N_7727);
and U8407 (N_8407,N_7827,N_7502);
or U8408 (N_8408,N_7534,N_7664);
or U8409 (N_8409,N_7990,N_7650);
nand U8410 (N_8410,N_7651,N_7954);
nor U8411 (N_8411,N_7862,N_7564);
nor U8412 (N_8412,N_7607,N_7613);
nor U8413 (N_8413,N_7689,N_7952);
nor U8414 (N_8414,N_7528,N_7587);
nand U8415 (N_8415,N_7627,N_7613);
or U8416 (N_8416,N_7804,N_7936);
and U8417 (N_8417,N_7937,N_7713);
and U8418 (N_8418,N_7539,N_7717);
nand U8419 (N_8419,N_7599,N_7632);
nor U8420 (N_8420,N_7581,N_7929);
xnor U8421 (N_8421,N_7742,N_7928);
and U8422 (N_8422,N_7927,N_7770);
xnor U8423 (N_8423,N_7576,N_7810);
and U8424 (N_8424,N_7748,N_7772);
xor U8425 (N_8425,N_7595,N_7877);
or U8426 (N_8426,N_7567,N_7593);
and U8427 (N_8427,N_7655,N_7598);
or U8428 (N_8428,N_7579,N_7633);
nor U8429 (N_8429,N_7665,N_7705);
and U8430 (N_8430,N_7978,N_7971);
nor U8431 (N_8431,N_7516,N_7779);
nor U8432 (N_8432,N_7730,N_7837);
nor U8433 (N_8433,N_7961,N_7833);
or U8434 (N_8434,N_7769,N_7584);
xor U8435 (N_8435,N_7988,N_7523);
xnor U8436 (N_8436,N_7501,N_7519);
xnor U8437 (N_8437,N_7993,N_7809);
and U8438 (N_8438,N_7582,N_7747);
nand U8439 (N_8439,N_7573,N_7848);
nand U8440 (N_8440,N_7724,N_7817);
xnor U8441 (N_8441,N_7709,N_7623);
nor U8442 (N_8442,N_7520,N_7951);
nor U8443 (N_8443,N_7874,N_7710);
and U8444 (N_8444,N_7858,N_7826);
or U8445 (N_8445,N_7658,N_7639);
or U8446 (N_8446,N_7628,N_7714);
nand U8447 (N_8447,N_7539,N_7833);
nand U8448 (N_8448,N_7641,N_7842);
nor U8449 (N_8449,N_7905,N_7799);
or U8450 (N_8450,N_7661,N_7698);
and U8451 (N_8451,N_7546,N_7694);
xor U8452 (N_8452,N_7660,N_7701);
nor U8453 (N_8453,N_7782,N_7983);
or U8454 (N_8454,N_7868,N_7670);
or U8455 (N_8455,N_7561,N_7924);
and U8456 (N_8456,N_7630,N_7686);
xnor U8457 (N_8457,N_7821,N_7774);
and U8458 (N_8458,N_7637,N_7932);
or U8459 (N_8459,N_7805,N_7934);
or U8460 (N_8460,N_7819,N_7576);
xor U8461 (N_8461,N_7863,N_7544);
nand U8462 (N_8462,N_7975,N_7577);
nor U8463 (N_8463,N_7984,N_7551);
nand U8464 (N_8464,N_7954,N_7588);
nor U8465 (N_8465,N_7866,N_7946);
xor U8466 (N_8466,N_7950,N_7548);
xnor U8467 (N_8467,N_7874,N_7754);
nor U8468 (N_8468,N_7509,N_7555);
nor U8469 (N_8469,N_7823,N_7782);
xnor U8470 (N_8470,N_7718,N_7935);
and U8471 (N_8471,N_7772,N_7972);
and U8472 (N_8472,N_7641,N_7989);
xnor U8473 (N_8473,N_7968,N_7633);
xor U8474 (N_8474,N_7902,N_7544);
and U8475 (N_8475,N_7638,N_7976);
xnor U8476 (N_8476,N_7903,N_7784);
and U8477 (N_8477,N_7806,N_7941);
nand U8478 (N_8478,N_7728,N_7703);
xor U8479 (N_8479,N_7724,N_7676);
and U8480 (N_8480,N_7796,N_7981);
or U8481 (N_8481,N_7666,N_7594);
nor U8482 (N_8482,N_7763,N_7875);
or U8483 (N_8483,N_7818,N_7786);
nand U8484 (N_8484,N_7815,N_7622);
nand U8485 (N_8485,N_7832,N_7766);
or U8486 (N_8486,N_7503,N_7549);
xnor U8487 (N_8487,N_7724,N_7581);
nor U8488 (N_8488,N_7602,N_7933);
nand U8489 (N_8489,N_7792,N_7594);
nand U8490 (N_8490,N_7637,N_7751);
or U8491 (N_8491,N_7714,N_7824);
nand U8492 (N_8492,N_7729,N_7641);
nor U8493 (N_8493,N_7501,N_7671);
nand U8494 (N_8494,N_7814,N_7524);
nand U8495 (N_8495,N_7944,N_7643);
and U8496 (N_8496,N_7943,N_7744);
nand U8497 (N_8497,N_7530,N_7537);
xor U8498 (N_8498,N_7948,N_7733);
xnor U8499 (N_8499,N_7900,N_7862);
nor U8500 (N_8500,N_8095,N_8191);
nor U8501 (N_8501,N_8242,N_8247);
and U8502 (N_8502,N_8213,N_8328);
or U8503 (N_8503,N_8188,N_8063);
or U8504 (N_8504,N_8365,N_8319);
or U8505 (N_8505,N_8079,N_8433);
nor U8506 (N_8506,N_8019,N_8056);
or U8507 (N_8507,N_8012,N_8417);
nand U8508 (N_8508,N_8218,N_8399);
nor U8509 (N_8509,N_8129,N_8042);
xnor U8510 (N_8510,N_8131,N_8226);
or U8511 (N_8511,N_8179,N_8177);
xnor U8512 (N_8512,N_8461,N_8344);
and U8513 (N_8513,N_8041,N_8215);
xnor U8514 (N_8514,N_8371,N_8406);
nor U8515 (N_8515,N_8462,N_8094);
or U8516 (N_8516,N_8361,N_8064);
xor U8517 (N_8517,N_8102,N_8241);
or U8518 (N_8518,N_8111,N_8379);
xor U8519 (N_8519,N_8029,N_8481);
nand U8520 (N_8520,N_8071,N_8496);
xor U8521 (N_8521,N_8023,N_8137);
xor U8522 (N_8522,N_8125,N_8122);
xnor U8523 (N_8523,N_8415,N_8031);
nor U8524 (N_8524,N_8002,N_8336);
nor U8525 (N_8525,N_8374,N_8109);
nor U8526 (N_8526,N_8455,N_8157);
nor U8527 (N_8527,N_8495,N_8225);
and U8528 (N_8528,N_8259,N_8091);
and U8529 (N_8529,N_8083,N_8018);
xnor U8530 (N_8530,N_8103,N_8312);
nand U8531 (N_8531,N_8222,N_8076);
and U8532 (N_8532,N_8460,N_8234);
or U8533 (N_8533,N_8421,N_8150);
or U8534 (N_8534,N_8113,N_8420);
nand U8535 (N_8535,N_8273,N_8473);
nand U8536 (N_8536,N_8450,N_8178);
and U8537 (N_8537,N_8491,N_8090);
and U8538 (N_8538,N_8112,N_8405);
xnor U8539 (N_8539,N_8118,N_8401);
and U8540 (N_8540,N_8490,N_8077);
nand U8541 (N_8541,N_8132,N_8224);
nor U8542 (N_8542,N_8182,N_8258);
nand U8543 (N_8543,N_8343,N_8161);
and U8544 (N_8544,N_8313,N_8010);
xor U8545 (N_8545,N_8232,N_8159);
xor U8546 (N_8546,N_8096,N_8016);
nand U8547 (N_8547,N_8230,N_8398);
and U8548 (N_8548,N_8283,N_8423);
xnor U8549 (N_8549,N_8451,N_8410);
nand U8550 (N_8550,N_8291,N_8395);
xor U8551 (N_8551,N_8075,N_8456);
or U8552 (N_8552,N_8289,N_8204);
xnor U8553 (N_8553,N_8447,N_8219);
nand U8554 (N_8554,N_8381,N_8295);
and U8555 (N_8555,N_8358,N_8020);
xor U8556 (N_8556,N_8181,N_8373);
nor U8557 (N_8557,N_8439,N_8338);
and U8558 (N_8558,N_8209,N_8434);
or U8559 (N_8559,N_8354,N_8176);
xor U8560 (N_8560,N_8380,N_8144);
xnor U8561 (N_8561,N_8217,N_8248);
and U8562 (N_8562,N_8277,N_8081);
nand U8563 (N_8563,N_8123,N_8389);
or U8564 (N_8564,N_8087,N_8073);
or U8565 (N_8565,N_8337,N_8452);
nand U8566 (N_8566,N_8292,N_8257);
or U8567 (N_8567,N_8483,N_8326);
and U8568 (N_8568,N_8418,N_8133);
nand U8569 (N_8569,N_8160,N_8397);
nand U8570 (N_8570,N_8249,N_8093);
xor U8571 (N_8571,N_8287,N_8032);
nor U8572 (N_8572,N_8175,N_8408);
nor U8573 (N_8573,N_8026,N_8015);
nor U8574 (N_8574,N_8255,N_8383);
nand U8575 (N_8575,N_8364,N_8021);
nor U8576 (N_8576,N_8311,N_8169);
nand U8577 (N_8577,N_8477,N_8430);
nand U8578 (N_8578,N_8274,N_8005);
and U8579 (N_8579,N_8369,N_8282);
nor U8580 (N_8580,N_8432,N_8046);
and U8581 (N_8581,N_8186,N_8448);
or U8582 (N_8582,N_8356,N_8074);
nand U8583 (N_8583,N_8372,N_8411);
nor U8584 (N_8584,N_8139,N_8040);
xnor U8585 (N_8585,N_8302,N_8315);
or U8586 (N_8586,N_8285,N_8055);
xor U8587 (N_8587,N_8350,N_8107);
nor U8588 (N_8588,N_8396,N_8297);
nor U8589 (N_8589,N_8011,N_8489);
xor U8590 (N_8590,N_8252,N_8256);
nor U8591 (N_8591,N_8378,N_8000);
xor U8592 (N_8592,N_8281,N_8233);
or U8593 (N_8593,N_8286,N_8146);
nand U8594 (N_8594,N_8480,N_8054);
nor U8595 (N_8595,N_8322,N_8310);
xnor U8596 (N_8596,N_8008,N_8488);
nor U8597 (N_8597,N_8268,N_8001);
or U8598 (N_8598,N_8105,N_8009);
nor U8599 (N_8599,N_8275,N_8168);
nor U8600 (N_8600,N_8429,N_8470);
xnor U8601 (N_8601,N_8366,N_8299);
or U8602 (N_8602,N_8143,N_8030);
nor U8603 (N_8603,N_8185,N_8493);
xor U8604 (N_8604,N_8329,N_8393);
xor U8605 (N_8605,N_8476,N_8239);
nand U8606 (N_8606,N_8135,N_8266);
xor U8607 (N_8607,N_8084,N_8147);
or U8608 (N_8608,N_8116,N_8419);
or U8609 (N_8609,N_8082,N_8163);
nor U8610 (N_8610,N_8216,N_8196);
and U8611 (N_8611,N_8183,N_8067);
or U8612 (N_8612,N_8357,N_8246);
nand U8613 (N_8613,N_8442,N_8482);
and U8614 (N_8614,N_8335,N_8154);
and U8615 (N_8615,N_8101,N_8057);
nor U8616 (N_8616,N_8036,N_8052);
nor U8617 (N_8617,N_8492,N_8426);
xnor U8618 (N_8618,N_8245,N_8059);
nor U8619 (N_8619,N_8013,N_8263);
xor U8620 (N_8620,N_8099,N_8276);
or U8621 (N_8621,N_8068,N_8404);
nor U8622 (N_8622,N_8235,N_8307);
nand U8623 (N_8623,N_8321,N_8278);
and U8624 (N_8624,N_8047,N_8089);
or U8625 (N_8625,N_8317,N_8388);
nor U8626 (N_8626,N_8375,N_8466);
nand U8627 (N_8627,N_8170,N_8352);
or U8628 (N_8628,N_8022,N_8192);
or U8629 (N_8629,N_8413,N_8271);
nand U8630 (N_8630,N_8262,N_8114);
nand U8631 (N_8631,N_8035,N_8007);
and U8632 (N_8632,N_8376,N_8141);
and U8633 (N_8633,N_8444,N_8156);
nor U8634 (N_8634,N_8060,N_8117);
nor U8635 (N_8635,N_8211,N_8458);
nor U8636 (N_8636,N_8305,N_8304);
nand U8637 (N_8637,N_8202,N_8485);
nor U8638 (N_8638,N_8228,N_8284);
or U8639 (N_8639,N_8203,N_8260);
or U8640 (N_8640,N_8360,N_8049);
or U8641 (N_8641,N_8425,N_8334);
xor U8642 (N_8642,N_8479,N_8104);
or U8643 (N_8643,N_8330,N_8208);
xnor U8644 (N_8644,N_8180,N_8237);
and U8645 (N_8645,N_8377,N_8184);
nand U8646 (N_8646,N_8347,N_8390);
or U8647 (N_8647,N_8353,N_8153);
or U8648 (N_8648,N_8323,N_8409);
and U8649 (N_8649,N_8387,N_8086);
xor U8650 (N_8650,N_8223,N_8288);
nor U8651 (N_8651,N_8043,N_8497);
nor U8652 (N_8652,N_8454,N_8333);
nor U8653 (N_8653,N_8424,N_8440);
nand U8654 (N_8654,N_8342,N_8435);
and U8655 (N_8655,N_8126,N_8340);
nand U8656 (N_8656,N_8048,N_8200);
nand U8657 (N_8657,N_8092,N_8155);
nor U8658 (N_8658,N_8058,N_8412);
or U8659 (N_8659,N_8345,N_8051);
xnor U8660 (N_8660,N_8003,N_8494);
and U8661 (N_8661,N_8320,N_8151);
and U8662 (N_8662,N_8072,N_8128);
nand U8663 (N_8663,N_8484,N_8486);
nor U8664 (N_8664,N_8261,N_8270);
nor U8665 (N_8665,N_8088,N_8045);
and U8666 (N_8666,N_8199,N_8314);
nand U8667 (N_8667,N_8253,N_8348);
nand U8668 (N_8668,N_8301,N_8325);
xor U8669 (N_8669,N_8264,N_8148);
or U8670 (N_8670,N_8244,N_8171);
nand U8671 (N_8671,N_8472,N_8362);
or U8672 (N_8672,N_8351,N_8368);
or U8673 (N_8673,N_8308,N_8487);
and U8674 (N_8674,N_8229,N_8498);
nor U8675 (N_8675,N_8385,N_8392);
or U8676 (N_8676,N_8106,N_8053);
xor U8677 (N_8677,N_8173,N_8427);
xor U8678 (N_8678,N_8166,N_8227);
xnor U8679 (N_8679,N_8386,N_8316);
xor U8680 (N_8680,N_8197,N_8475);
xor U8681 (N_8681,N_8469,N_8459);
and U8682 (N_8682,N_8457,N_8165);
or U8683 (N_8683,N_8294,N_8303);
nor U8684 (N_8684,N_8212,N_8400);
xnor U8685 (N_8685,N_8471,N_8024);
or U8686 (N_8686,N_8130,N_8474);
nor U8687 (N_8687,N_8441,N_8231);
xor U8688 (N_8688,N_8422,N_8119);
and U8689 (N_8689,N_8044,N_8164);
and U8690 (N_8690,N_8414,N_8250);
nor U8691 (N_8691,N_8201,N_8463);
xor U8692 (N_8692,N_8428,N_8062);
nand U8693 (N_8693,N_8443,N_8341);
nand U8694 (N_8694,N_8193,N_8346);
or U8695 (N_8695,N_8145,N_8403);
and U8696 (N_8696,N_8134,N_8070);
nand U8697 (N_8697,N_8198,N_8167);
and U8698 (N_8698,N_8120,N_8267);
nand U8699 (N_8699,N_8391,N_8033);
xor U8700 (N_8700,N_8190,N_8355);
and U8701 (N_8701,N_8431,N_8124);
and U8702 (N_8702,N_8446,N_8115);
or U8703 (N_8703,N_8017,N_8014);
or U8704 (N_8704,N_8449,N_8367);
nor U8705 (N_8705,N_8382,N_8453);
xor U8706 (N_8706,N_8078,N_8006);
xnor U8707 (N_8707,N_8324,N_8331);
nand U8708 (N_8708,N_8272,N_8085);
nor U8709 (N_8709,N_8158,N_8437);
and U8710 (N_8710,N_8110,N_8066);
nand U8711 (N_8711,N_8384,N_8416);
xor U8712 (N_8712,N_8478,N_8306);
nor U8713 (N_8713,N_8243,N_8254);
nand U8714 (N_8714,N_8214,N_8300);
and U8715 (N_8715,N_8327,N_8298);
nor U8716 (N_8716,N_8332,N_8069);
xor U8717 (N_8717,N_8004,N_8136);
or U8718 (N_8718,N_8038,N_8318);
xor U8719 (N_8719,N_8065,N_8269);
xor U8720 (N_8720,N_8370,N_8050);
nand U8721 (N_8721,N_8034,N_8028);
nor U8722 (N_8722,N_8468,N_8207);
nand U8723 (N_8723,N_8363,N_8025);
nor U8724 (N_8724,N_8187,N_8174);
nor U8725 (N_8725,N_8100,N_8039);
nand U8726 (N_8726,N_8098,N_8499);
or U8727 (N_8727,N_8296,N_8359);
or U8728 (N_8728,N_8206,N_8097);
nand U8729 (N_8729,N_8265,N_8438);
xor U8730 (N_8730,N_8445,N_8279);
and U8731 (N_8731,N_8037,N_8339);
and U8732 (N_8732,N_8407,N_8220);
nor U8733 (N_8733,N_8189,N_8061);
xor U8734 (N_8734,N_8309,N_8402);
nor U8735 (N_8735,N_8108,N_8195);
or U8736 (N_8736,N_8027,N_8465);
xor U8737 (N_8737,N_8138,N_8194);
nor U8738 (N_8738,N_8236,N_8349);
nor U8739 (N_8739,N_8149,N_8221);
nor U8740 (N_8740,N_8290,N_8280);
or U8741 (N_8741,N_8205,N_8464);
nand U8742 (N_8742,N_8142,N_8162);
nor U8743 (N_8743,N_8080,N_8140);
and U8744 (N_8744,N_8293,N_8121);
nor U8745 (N_8745,N_8394,N_8251);
nor U8746 (N_8746,N_8467,N_8127);
and U8747 (N_8747,N_8436,N_8210);
or U8748 (N_8748,N_8172,N_8152);
xnor U8749 (N_8749,N_8238,N_8240);
xor U8750 (N_8750,N_8499,N_8431);
nand U8751 (N_8751,N_8035,N_8389);
nand U8752 (N_8752,N_8316,N_8130);
nor U8753 (N_8753,N_8051,N_8098);
and U8754 (N_8754,N_8101,N_8279);
xor U8755 (N_8755,N_8404,N_8073);
nand U8756 (N_8756,N_8472,N_8034);
or U8757 (N_8757,N_8096,N_8383);
or U8758 (N_8758,N_8425,N_8440);
nand U8759 (N_8759,N_8019,N_8313);
nand U8760 (N_8760,N_8271,N_8284);
or U8761 (N_8761,N_8242,N_8108);
xnor U8762 (N_8762,N_8078,N_8087);
or U8763 (N_8763,N_8450,N_8155);
or U8764 (N_8764,N_8348,N_8188);
and U8765 (N_8765,N_8179,N_8229);
nand U8766 (N_8766,N_8250,N_8324);
or U8767 (N_8767,N_8222,N_8127);
nor U8768 (N_8768,N_8202,N_8310);
or U8769 (N_8769,N_8105,N_8471);
nor U8770 (N_8770,N_8042,N_8223);
nand U8771 (N_8771,N_8311,N_8208);
xor U8772 (N_8772,N_8259,N_8331);
xor U8773 (N_8773,N_8041,N_8216);
nor U8774 (N_8774,N_8142,N_8490);
or U8775 (N_8775,N_8301,N_8167);
nand U8776 (N_8776,N_8127,N_8098);
nor U8777 (N_8777,N_8216,N_8191);
xnor U8778 (N_8778,N_8346,N_8460);
nor U8779 (N_8779,N_8187,N_8420);
or U8780 (N_8780,N_8282,N_8240);
xnor U8781 (N_8781,N_8292,N_8374);
or U8782 (N_8782,N_8466,N_8232);
nor U8783 (N_8783,N_8157,N_8045);
nand U8784 (N_8784,N_8485,N_8287);
xnor U8785 (N_8785,N_8241,N_8227);
xnor U8786 (N_8786,N_8477,N_8157);
and U8787 (N_8787,N_8458,N_8217);
and U8788 (N_8788,N_8093,N_8374);
xnor U8789 (N_8789,N_8068,N_8342);
or U8790 (N_8790,N_8132,N_8397);
nand U8791 (N_8791,N_8449,N_8028);
nand U8792 (N_8792,N_8294,N_8119);
nand U8793 (N_8793,N_8009,N_8413);
nor U8794 (N_8794,N_8336,N_8182);
nand U8795 (N_8795,N_8162,N_8377);
xor U8796 (N_8796,N_8187,N_8027);
nand U8797 (N_8797,N_8364,N_8298);
nor U8798 (N_8798,N_8090,N_8330);
or U8799 (N_8799,N_8310,N_8407);
nor U8800 (N_8800,N_8400,N_8476);
nor U8801 (N_8801,N_8462,N_8385);
nand U8802 (N_8802,N_8346,N_8366);
nor U8803 (N_8803,N_8003,N_8425);
or U8804 (N_8804,N_8478,N_8297);
or U8805 (N_8805,N_8444,N_8425);
or U8806 (N_8806,N_8162,N_8112);
nor U8807 (N_8807,N_8469,N_8209);
and U8808 (N_8808,N_8428,N_8453);
nand U8809 (N_8809,N_8021,N_8005);
and U8810 (N_8810,N_8173,N_8043);
or U8811 (N_8811,N_8020,N_8287);
nand U8812 (N_8812,N_8368,N_8213);
or U8813 (N_8813,N_8461,N_8140);
or U8814 (N_8814,N_8065,N_8203);
nand U8815 (N_8815,N_8155,N_8252);
nor U8816 (N_8816,N_8268,N_8047);
nand U8817 (N_8817,N_8029,N_8224);
nor U8818 (N_8818,N_8482,N_8451);
xor U8819 (N_8819,N_8403,N_8460);
xnor U8820 (N_8820,N_8126,N_8117);
nor U8821 (N_8821,N_8351,N_8029);
xor U8822 (N_8822,N_8197,N_8369);
and U8823 (N_8823,N_8332,N_8463);
and U8824 (N_8824,N_8185,N_8145);
nand U8825 (N_8825,N_8317,N_8140);
and U8826 (N_8826,N_8223,N_8246);
nor U8827 (N_8827,N_8189,N_8310);
nor U8828 (N_8828,N_8156,N_8288);
or U8829 (N_8829,N_8391,N_8232);
and U8830 (N_8830,N_8382,N_8035);
xor U8831 (N_8831,N_8078,N_8134);
nand U8832 (N_8832,N_8408,N_8144);
or U8833 (N_8833,N_8474,N_8486);
and U8834 (N_8834,N_8092,N_8451);
and U8835 (N_8835,N_8319,N_8405);
or U8836 (N_8836,N_8196,N_8198);
and U8837 (N_8837,N_8143,N_8015);
nand U8838 (N_8838,N_8314,N_8272);
nand U8839 (N_8839,N_8296,N_8363);
or U8840 (N_8840,N_8115,N_8374);
and U8841 (N_8841,N_8243,N_8489);
nor U8842 (N_8842,N_8145,N_8279);
xor U8843 (N_8843,N_8258,N_8015);
and U8844 (N_8844,N_8092,N_8452);
nor U8845 (N_8845,N_8384,N_8032);
or U8846 (N_8846,N_8131,N_8472);
or U8847 (N_8847,N_8128,N_8479);
and U8848 (N_8848,N_8355,N_8221);
or U8849 (N_8849,N_8362,N_8293);
xor U8850 (N_8850,N_8137,N_8260);
nor U8851 (N_8851,N_8038,N_8252);
nand U8852 (N_8852,N_8342,N_8362);
nor U8853 (N_8853,N_8491,N_8139);
or U8854 (N_8854,N_8407,N_8370);
and U8855 (N_8855,N_8004,N_8324);
nor U8856 (N_8856,N_8010,N_8135);
nor U8857 (N_8857,N_8484,N_8306);
and U8858 (N_8858,N_8302,N_8082);
and U8859 (N_8859,N_8023,N_8134);
nor U8860 (N_8860,N_8435,N_8074);
and U8861 (N_8861,N_8362,N_8416);
and U8862 (N_8862,N_8029,N_8080);
nor U8863 (N_8863,N_8476,N_8204);
or U8864 (N_8864,N_8421,N_8100);
nand U8865 (N_8865,N_8042,N_8173);
or U8866 (N_8866,N_8375,N_8417);
and U8867 (N_8867,N_8207,N_8292);
and U8868 (N_8868,N_8105,N_8347);
nor U8869 (N_8869,N_8355,N_8130);
or U8870 (N_8870,N_8198,N_8463);
nor U8871 (N_8871,N_8336,N_8017);
nand U8872 (N_8872,N_8234,N_8133);
nand U8873 (N_8873,N_8238,N_8392);
and U8874 (N_8874,N_8387,N_8280);
nor U8875 (N_8875,N_8150,N_8118);
nand U8876 (N_8876,N_8227,N_8127);
nor U8877 (N_8877,N_8021,N_8212);
xnor U8878 (N_8878,N_8428,N_8410);
xnor U8879 (N_8879,N_8209,N_8270);
nor U8880 (N_8880,N_8057,N_8013);
nand U8881 (N_8881,N_8428,N_8308);
nor U8882 (N_8882,N_8237,N_8125);
or U8883 (N_8883,N_8388,N_8032);
xor U8884 (N_8884,N_8144,N_8399);
xnor U8885 (N_8885,N_8141,N_8050);
xor U8886 (N_8886,N_8406,N_8353);
or U8887 (N_8887,N_8319,N_8358);
xor U8888 (N_8888,N_8440,N_8423);
nand U8889 (N_8889,N_8315,N_8244);
or U8890 (N_8890,N_8489,N_8387);
and U8891 (N_8891,N_8142,N_8445);
and U8892 (N_8892,N_8299,N_8173);
nand U8893 (N_8893,N_8300,N_8155);
nand U8894 (N_8894,N_8108,N_8323);
or U8895 (N_8895,N_8044,N_8473);
and U8896 (N_8896,N_8103,N_8301);
nor U8897 (N_8897,N_8168,N_8432);
nor U8898 (N_8898,N_8295,N_8200);
nand U8899 (N_8899,N_8177,N_8420);
nand U8900 (N_8900,N_8151,N_8160);
nor U8901 (N_8901,N_8396,N_8181);
nand U8902 (N_8902,N_8113,N_8487);
and U8903 (N_8903,N_8157,N_8178);
xor U8904 (N_8904,N_8348,N_8050);
and U8905 (N_8905,N_8395,N_8348);
xor U8906 (N_8906,N_8423,N_8184);
or U8907 (N_8907,N_8250,N_8496);
nand U8908 (N_8908,N_8031,N_8140);
nand U8909 (N_8909,N_8248,N_8034);
and U8910 (N_8910,N_8279,N_8414);
and U8911 (N_8911,N_8454,N_8064);
nand U8912 (N_8912,N_8051,N_8350);
or U8913 (N_8913,N_8143,N_8084);
xor U8914 (N_8914,N_8202,N_8399);
xor U8915 (N_8915,N_8399,N_8074);
and U8916 (N_8916,N_8222,N_8310);
and U8917 (N_8917,N_8081,N_8226);
nand U8918 (N_8918,N_8031,N_8477);
and U8919 (N_8919,N_8018,N_8030);
xnor U8920 (N_8920,N_8031,N_8272);
nor U8921 (N_8921,N_8138,N_8002);
or U8922 (N_8922,N_8189,N_8315);
nor U8923 (N_8923,N_8114,N_8191);
nand U8924 (N_8924,N_8054,N_8370);
nor U8925 (N_8925,N_8480,N_8237);
nand U8926 (N_8926,N_8100,N_8016);
xor U8927 (N_8927,N_8243,N_8323);
xor U8928 (N_8928,N_8006,N_8350);
nand U8929 (N_8929,N_8433,N_8475);
and U8930 (N_8930,N_8157,N_8275);
nor U8931 (N_8931,N_8212,N_8051);
and U8932 (N_8932,N_8418,N_8338);
nor U8933 (N_8933,N_8393,N_8029);
or U8934 (N_8934,N_8043,N_8013);
or U8935 (N_8935,N_8444,N_8084);
nand U8936 (N_8936,N_8084,N_8375);
nand U8937 (N_8937,N_8323,N_8221);
nor U8938 (N_8938,N_8431,N_8447);
xor U8939 (N_8939,N_8018,N_8438);
nand U8940 (N_8940,N_8136,N_8206);
and U8941 (N_8941,N_8083,N_8101);
nor U8942 (N_8942,N_8292,N_8038);
nand U8943 (N_8943,N_8066,N_8026);
nand U8944 (N_8944,N_8250,N_8073);
nand U8945 (N_8945,N_8370,N_8280);
and U8946 (N_8946,N_8042,N_8447);
or U8947 (N_8947,N_8153,N_8454);
or U8948 (N_8948,N_8156,N_8048);
xor U8949 (N_8949,N_8093,N_8172);
nand U8950 (N_8950,N_8100,N_8395);
nor U8951 (N_8951,N_8450,N_8463);
xor U8952 (N_8952,N_8289,N_8449);
or U8953 (N_8953,N_8198,N_8309);
nor U8954 (N_8954,N_8049,N_8171);
and U8955 (N_8955,N_8266,N_8260);
nor U8956 (N_8956,N_8409,N_8026);
nor U8957 (N_8957,N_8222,N_8106);
and U8958 (N_8958,N_8260,N_8114);
nor U8959 (N_8959,N_8365,N_8411);
or U8960 (N_8960,N_8251,N_8111);
nand U8961 (N_8961,N_8071,N_8056);
and U8962 (N_8962,N_8135,N_8019);
xor U8963 (N_8963,N_8386,N_8477);
or U8964 (N_8964,N_8184,N_8334);
and U8965 (N_8965,N_8381,N_8435);
xnor U8966 (N_8966,N_8404,N_8460);
or U8967 (N_8967,N_8211,N_8352);
or U8968 (N_8968,N_8198,N_8107);
or U8969 (N_8969,N_8133,N_8142);
and U8970 (N_8970,N_8433,N_8162);
nor U8971 (N_8971,N_8038,N_8235);
nor U8972 (N_8972,N_8171,N_8225);
xor U8973 (N_8973,N_8152,N_8224);
and U8974 (N_8974,N_8488,N_8322);
and U8975 (N_8975,N_8041,N_8188);
nand U8976 (N_8976,N_8037,N_8491);
or U8977 (N_8977,N_8140,N_8245);
or U8978 (N_8978,N_8112,N_8226);
xor U8979 (N_8979,N_8105,N_8412);
and U8980 (N_8980,N_8424,N_8198);
and U8981 (N_8981,N_8296,N_8124);
nor U8982 (N_8982,N_8494,N_8419);
or U8983 (N_8983,N_8152,N_8453);
nor U8984 (N_8984,N_8424,N_8027);
nand U8985 (N_8985,N_8311,N_8386);
or U8986 (N_8986,N_8224,N_8431);
xnor U8987 (N_8987,N_8331,N_8317);
xor U8988 (N_8988,N_8292,N_8046);
and U8989 (N_8989,N_8067,N_8263);
xnor U8990 (N_8990,N_8055,N_8208);
nor U8991 (N_8991,N_8024,N_8138);
and U8992 (N_8992,N_8235,N_8105);
and U8993 (N_8993,N_8197,N_8136);
nand U8994 (N_8994,N_8428,N_8089);
or U8995 (N_8995,N_8415,N_8052);
nor U8996 (N_8996,N_8432,N_8408);
nand U8997 (N_8997,N_8139,N_8326);
and U8998 (N_8998,N_8372,N_8498);
nand U8999 (N_8999,N_8289,N_8326);
xor U9000 (N_9000,N_8959,N_8580);
nand U9001 (N_9001,N_8935,N_8940);
or U9002 (N_9002,N_8833,N_8504);
nor U9003 (N_9003,N_8747,N_8626);
nand U9004 (N_9004,N_8948,N_8752);
xnor U9005 (N_9005,N_8583,N_8568);
nor U9006 (N_9006,N_8880,N_8772);
nor U9007 (N_9007,N_8901,N_8511);
xor U9008 (N_9008,N_8905,N_8814);
xnor U9009 (N_9009,N_8849,N_8910);
and U9010 (N_9010,N_8803,N_8933);
or U9011 (N_9011,N_8534,N_8947);
nand U9012 (N_9012,N_8770,N_8980);
nor U9013 (N_9013,N_8506,N_8544);
nand U9014 (N_9014,N_8919,N_8605);
nand U9015 (N_9015,N_8804,N_8885);
or U9016 (N_9016,N_8711,N_8657);
and U9017 (N_9017,N_8864,N_8682);
nand U9018 (N_9018,N_8547,N_8665);
or U9019 (N_9019,N_8956,N_8855);
xor U9020 (N_9020,N_8684,N_8923);
nor U9021 (N_9021,N_8955,N_8782);
or U9022 (N_9022,N_8694,N_8845);
nand U9023 (N_9023,N_8664,N_8687);
and U9024 (N_9024,N_8979,N_8899);
or U9025 (N_9025,N_8718,N_8915);
or U9026 (N_9026,N_8674,N_8517);
or U9027 (N_9027,N_8774,N_8525);
nor U9028 (N_9028,N_8603,N_8843);
nand U9029 (N_9029,N_8810,N_8714);
nor U9030 (N_9030,N_8937,N_8699);
or U9031 (N_9031,N_8667,N_8705);
nor U9032 (N_9032,N_8670,N_8668);
nor U9033 (N_9033,N_8823,N_8552);
xor U9034 (N_9034,N_8591,N_8872);
nor U9035 (N_9035,N_8912,N_8863);
nor U9036 (N_9036,N_8573,N_8817);
and U9037 (N_9037,N_8725,N_8613);
nand U9038 (N_9038,N_8615,N_8928);
xor U9039 (N_9039,N_8913,N_8777);
xor U9040 (N_9040,N_8637,N_8761);
xnor U9041 (N_9041,N_8743,N_8695);
xnor U9042 (N_9042,N_8530,N_8733);
and U9043 (N_9043,N_8622,N_8726);
or U9044 (N_9044,N_8543,N_8712);
or U9045 (N_9045,N_8867,N_8531);
and U9046 (N_9046,N_8852,N_8986);
nand U9047 (N_9047,N_8997,N_8848);
nand U9048 (N_9048,N_8798,N_8529);
or U9049 (N_9049,N_8588,N_8751);
nor U9050 (N_9050,N_8775,N_8697);
nand U9051 (N_9051,N_8945,N_8551);
xor U9052 (N_9052,N_8930,N_8505);
xnor U9053 (N_9053,N_8784,N_8541);
and U9054 (N_9054,N_8837,N_8688);
xnor U9055 (N_9055,N_8652,N_8851);
nand U9056 (N_9056,N_8510,N_8553);
nand U9057 (N_9057,N_8520,N_8918);
nor U9058 (N_9058,N_8644,N_8868);
and U9059 (N_9059,N_8710,N_8981);
nor U9060 (N_9060,N_8883,N_8974);
nand U9061 (N_9061,N_8653,N_8716);
or U9062 (N_9062,N_8819,N_8965);
nor U9063 (N_9063,N_8987,N_8985);
nand U9064 (N_9064,N_8528,N_8713);
nor U9065 (N_9065,N_8834,N_8917);
nor U9066 (N_9066,N_8691,N_8887);
and U9067 (N_9067,N_8602,N_8732);
nand U9068 (N_9068,N_8526,N_8572);
or U9069 (N_9069,N_8701,N_8642);
nor U9070 (N_9070,N_8686,N_8633);
and U9071 (N_9071,N_8621,N_8562);
or U9072 (N_9072,N_8557,N_8856);
nor U9073 (N_9073,N_8973,N_8595);
nor U9074 (N_9074,N_8574,N_8735);
xnor U9075 (N_9075,N_8627,N_8625);
xnor U9076 (N_9076,N_8631,N_8600);
or U9077 (N_9077,N_8961,N_8779);
and U9078 (N_9078,N_8767,N_8607);
nor U9079 (N_9079,N_8717,N_8599);
and U9080 (N_9080,N_8921,N_8828);
and U9081 (N_9081,N_8629,N_8820);
and U9082 (N_9082,N_8728,N_8939);
nor U9083 (N_9083,N_8748,N_8651);
xor U9084 (N_9084,N_8739,N_8976);
and U9085 (N_9085,N_8860,N_8857);
and U9086 (N_9086,N_8677,N_8821);
xnor U9087 (N_9087,N_8753,N_8720);
or U9088 (N_9088,N_8805,N_8620);
xor U9089 (N_9089,N_8755,N_8978);
nor U9090 (N_9090,N_8795,N_8922);
and U9091 (N_9091,N_8990,N_8598);
and U9092 (N_9092,N_8508,N_8892);
or U9093 (N_9093,N_8962,N_8842);
xnor U9094 (N_9094,N_8991,N_8877);
or U9095 (N_9095,N_8632,N_8781);
or U9096 (N_9096,N_8999,N_8865);
xnor U9097 (N_9097,N_8916,N_8659);
nor U9098 (N_9098,N_8731,N_8938);
xnor U9099 (N_9099,N_8623,N_8815);
nor U9100 (N_9100,N_8903,N_8610);
nor U9101 (N_9101,N_8749,N_8730);
nand U9102 (N_9102,N_8908,N_8567);
or U9103 (N_9103,N_8869,N_8709);
and U9104 (N_9104,N_8617,N_8523);
nor U9105 (N_9105,N_8967,N_8744);
or U9106 (N_9106,N_8931,N_8545);
nand U9107 (N_9107,N_8745,N_8977);
or U9108 (N_9108,N_8764,N_8746);
nand U9109 (N_9109,N_8886,N_8783);
xor U9110 (N_9110,N_8952,N_8638);
and U9111 (N_9111,N_8565,N_8540);
and U9112 (N_9112,N_8862,N_8584);
nor U9113 (N_9113,N_8577,N_8693);
nand U9114 (N_9114,N_8970,N_8509);
xor U9115 (N_9115,N_8757,N_8776);
or U9116 (N_9116,N_8640,N_8563);
nor U9117 (N_9117,N_8786,N_8972);
xor U9118 (N_9118,N_8942,N_8953);
xor U9119 (N_9119,N_8721,N_8888);
xnor U9120 (N_9120,N_8788,N_8966);
nand U9121 (N_9121,N_8984,N_8507);
nand U9122 (N_9122,N_8581,N_8809);
and U9123 (N_9123,N_8822,N_8616);
or U9124 (N_9124,N_8590,N_8554);
and U9125 (N_9125,N_8858,N_8654);
nand U9126 (N_9126,N_8597,N_8762);
and U9127 (N_9127,N_8946,N_8983);
xor U9128 (N_9128,N_8854,N_8927);
or U9129 (N_9129,N_8614,N_8649);
and U9130 (N_9130,N_8894,N_8904);
nor U9131 (N_9131,N_8555,N_8835);
and U9132 (N_9132,N_8518,N_8715);
xor U9133 (N_9133,N_8660,N_8673);
or U9134 (N_9134,N_8698,N_8811);
or U9135 (N_9135,N_8995,N_8870);
nand U9136 (N_9136,N_8890,N_8796);
xnor U9137 (N_9137,N_8592,N_8683);
or U9138 (N_9138,N_8909,N_8969);
and U9139 (N_9139,N_8502,N_8911);
or U9140 (N_9140,N_8832,N_8576);
or U9141 (N_9141,N_8550,N_8926);
xnor U9142 (N_9142,N_8586,N_8706);
or U9143 (N_9143,N_8643,N_8521);
nand U9144 (N_9144,N_8900,N_8645);
and U9145 (N_9145,N_8636,N_8839);
nor U9146 (N_9146,N_8561,N_8873);
and U9147 (N_9147,N_8758,N_8662);
and U9148 (N_9148,N_8516,N_8846);
or U9149 (N_9149,N_8532,N_8988);
or U9150 (N_9150,N_8612,N_8708);
xnor U9151 (N_9151,N_8794,N_8771);
nor U9152 (N_9152,N_8963,N_8558);
xor U9153 (N_9153,N_8537,N_8907);
xnor U9154 (N_9154,N_8703,N_8527);
and U9155 (N_9155,N_8524,N_8736);
and U9156 (N_9156,N_8679,N_8719);
and U9157 (N_9157,N_8941,N_8676);
or U9158 (N_9158,N_8853,N_8648);
nand U9159 (N_9159,N_8756,N_8785);
or U9160 (N_9160,N_8875,N_8797);
nand U9161 (N_9161,N_8964,N_8876);
nor U9162 (N_9162,N_8929,N_8608);
xnor U9163 (N_9163,N_8889,N_8696);
or U9164 (N_9164,N_8950,N_8704);
and U9165 (N_9165,N_8800,N_8601);
nand U9166 (N_9166,N_8639,N_8850);
or U9167 (N_9167,N_8951,N_8861);
xnor U9168 (N_9168,N_8968,N_8829);
and U9169 (N_9169,N_8564,N_8884);
and U9170 (N_9170,N_8570,N_8936);
xor U9171 (N_9171,N_8826,N_8738);
and U9172 (N_9172,N_8723,N_8944);
and U9173 (N_9173,N_8932,N_8878);
or U9174 (N_9174,N_8596,N_8998);
or U9175 (N_9175,N_8957,N_8992);
xor U9176 (N_9176,N_8994,N_8658);
xor U9177 (N_9177,N_8802,N_8535);
nand U9178 (N_9178,N_8896,N_8836);
xor U9179 (N_9179,N_8801,N_8678);
and U9180 (N_9180,N_8575,N_8647);
nor U9181 (N_9181,N_8840,N_8895);
nand U9182 (N_9182,N_8655,N_8898);
xnor U9183 (N_9183,N_8727,N_8816);
or U9184 (N_9184,N_8806,N_8750);
nor U9185 (N_9185,N_8827,N_8866);
or U9186 (N_9186,N_8996,N_8650);
or U9187 (N_9187,N_8793,N_8675);
nand U9188 (N_9188,N_8954,N_8663);
xnor U9189 (N_9189,N_8734,N_8538);
xnor U9190 (N_9190,N_8808,N_8635);
or U9191 (N_9191,N_8780,N_8807);
nor U9192 (N_9192,N_8702,N_8542);
xnor U9193 (N_9193,N_8812,N_8740);
nor U9194 (N_9194,N_8949,N_8766);
nand U9195 (N_9195,N_8585,N_8533);
or U9196 (N_9196,N_8566,N_8859);
nand U9197 (N_9197,N_8813,N_8559);
or U9198 (N_9198,N_8666,N_8539);
and U9199 (N_9199,N_8619,N_8501);
or U9200 (N_9200,N_8993,N_8789);
and U9201 (N_9201,N_8871,N_8790);
nand U9202 (N_9202,N_8891,N_8515);
or U9203 (N_9203,N_8519,N_8844);
nand U9204 (N_9204,N_8513,N_8881);
or U9205 (N_9205,N_8742,N_8556);
nand U9206 (N_9206,N_8924,N_8609);
and U9207 (N_9207,N_8594,N_8689);
xor U9208 (N_9208,N_8641,N_8611);
xor U9209 (N_9209,N_8989,N_8671);
or U9210 (N_9210,N_8646,N_8549);
nor U9211 (N_9211,N_8522,N_8824);
and U9212 (N_9212,N_8792,N_8536);
xor U9213 (N_9213,N_8773,N_8879);
xor U9214 (N_9214,N_8512,N_8765);
or U9215 (N_9215,N_8624,N_8690);
or U9216 (N_9216,N_8604,N_8759);
nor U9217 (N_9217,N_8825,N_8787);
nor U9218 (N_9218,N_8982,N_8634);
or U9219 (N_9219,N_8882,N_8724);
nor U9220 (N_9220,N_8778,N_8669);
nand U9221 (N_9221,N_8582,N_8831);
xnor U9222 (N_9222,N_8587,N_8958);
or U9223 (N_9223,N_8500,N_8578);
xnor U9224 (N_9224,N_8589,N_8548);
nor U9225 (N_9225,N_8681,N_8754);
and U9226 (N_9226,N_8707,N_8656);
nor U9227 (N_9227,N_8571,N_8902);
xor U9228 (N_9228,N_8769,N_8893);
and U9229 (N_9229,N_8685,N_8841);
nand U9230 (N_9230,N_8838,N_8503);
xor U9231 (N_9231,N_8763,N_8630);
nand U9232 (N_9232,N_8672,N_8741);
nand U9233 (N_9233,N_8628,N_8768);
xor U9234 (N_9234,N_8680,N_8943);
nor U9235 (N_9235,N_8818,N_8925);
and U9236 (N_9236,N_8593,N_8722);
nand U9237 (N_9237,N_8791,N_8569);
and U9238 (N_9238,N_8847,N_8546);
or U9239 (N_9239,N_8960,N_8700);
nand U9240 (N_9240,N_8737,N_8906);
nand U9241 (N_9241,N_8560,N_8920);
nand U9242 (N_9242,N_8514,N_8975);
nor U9243 (N_9243,N_8914,N_8830);
or U9244 (N_9244,N_8897,N_8874);
and U9245 (N_9245,N_8971,N_8799);
or U9246 (N_9246,N_8661,N_8729);
nor U9247 (N_9247,N_8692,N_8579);
nor U9248 (N_9248,N_8606,N_8934);
nand U9249 (N_9249,N_8618,N_8760);
and U9250 (N_9250,N_8678,N_8785);
and U9251 (N_9251,N_8596,N_8564);
and U9252 (N_9252,N_8533,N_8779);
nand U9253 (N_9253,N_8996,N_8711);
xnor U9254 (N_9254,N_8984,N_8645);
nor U9255 (N_9255,N_8517,N_8653);
nor U9256 (N_9256,N_8501,N_8535);
nor U9257 (N_9257,N_8506,N_8821);
and U9258 (N_9258,N_8700,N_8800);
or U9259 (N_9259,N_8955,N_8968);
xnor U9260 (N_9260,N_8953,N_8670);
nand U9261 (N_9261,N_8584,N_8713);
nor U9262 (N_9262,N_8743,N_8770);
nor U9263 (N_9263,N_8737,N_8793);
and U9264 (N_9264,N_8767,N_8731);
or U9265 (N_9265,N_8585,N_8638);
and U9266 (N_9266,N_8870,N_8592);
nand U9267 (N_9267,N_8544,N_8594);
xnor U9268 (N_9268,N_8725,N_8636);
xnor U9269 (N_9269,N_8944,N_8993);
or U9270 (N_9270,N_8788,N_8699);
nand U9271 (N_9271,N_8984,N_8732);
and U9272 (N_9272,N_8501,N_8945);
nand U9273 (N_9273,N_8924,N_8804);
nand U9274 (N_9274,N_8692,N_8724);
or U9275 (N_9275,N_8579,N_8814);
xnor U9276 (N_9276,N_8939,N_8708);
nor U9277 (N_9277,N_8598,N_8622);
or U9278 (N_9278,N_8550,N_8915);
nand U9279 (N_9279,N_8678,N_8550);
and U9280 (N_9280,N_8755,N_8802);
nor U9281 (N_9281,N_8741,N_8589);
nor U9282 (N_9282,N_8614,N_8929);
xnor U9283 (N_9283,N_8948,N_8919);
nor U9284 (N_9284,N_8817,N_8876);
nor U9285 (N_9285,N_8595,N_8969);
nand U9286 (N_9286,N_8520,N_8897);
xnor U9287 (N_9287,N_8878,N_8966);
nor U9288 (N_9288,N_8638,N_8621);
or U9289 (N_9289,N_8833,N_8961);
or U9290 (N_9290,N_8723,N_8777);
and U9291 (N_9291,N_8526,N_8589);
and U9292 (N_9292,N_8895,N_8971);
xor U9293 (N_9293,N_8751,N_8934);
and U9294 (N_9294,N_8545,N_8520);
nand U9295 (N_9295,N_8957,N_8731);
or U9296 (N_9296,N_8723,N_8593);
xor U9297 (N_9297,N_8628,N_8664);
and U9298 (N_9298,N_8971,N_8879);
xnor U9299 (N_9299,N_8508,N_8851);
nand U9300 (N_9300,N_8554,N_8581);
nand U9301 (N_9301,N_8622,N_8648);
nand U9302 (N_9302,N_8825,N_8684);
or U9303 (N_9303,N_8732,N_8841);
nand U9304 (N_9304,N_8779,N_8518);
nor U9305 (N_9305,N_8718,N_8500);
xnor U9306 (N_9306,N_8836,N_8823);
or U9307 (N_9307,N_8562,N_8940);
and U9308 (N_9308,N_8832,N_8677);
or U9309 (N_9309,N_8665,N_8663);
and U9310 (N_9310,N_8623,N_8924);
and U9311 (N_9311,N_8821,N_8518);
xor U9312 (N_9312,N_8749,N_8731);
and U9313 (N_9313,N_8826,N_8982);
xnor U9314 (N_9314,N_8579,N_8654);
or U9315 (N_9315,N_8865,N_8567);
xor U9316 (N_9316,N_8784,N_8525);
nor U9317 (N_9317,N_8910,N_8847);
nand U9318 (N_9318,N_8685,N_8574);
xnor U9319 (N_9319,N_8810,N_8727);
and U9320 (N_9320,N_8590,N_8696);
or U9321 (N_9321,N_8722,N_8573);
or U9322 (N_9322,N_8706,N_8544);
xnor U9323 (N_9323,N_8828,N_8833);
nand U9324 (N_9324,N_8610,N_8819);
nand U9325 (N_9325,N_8596,N_8715);
xnor U9326 (N_9326,N_8736,N_8690);
or U9327 (N_9327,N_8603,N_8943);
nand U9328 (N_9328,N_8647,N_8533);
nand U9329 (N_9329,N_8533,N_8783);
and U9330 (N_9330,N_8664,N_8643);
and U9331 (N_9331,N_8744,N_8913);
xnor U9332 (N_9332,N_8584,N_8976);
and U9333 (N_9333,N_8911,N_8804);
xor U9334 (N_9334,N_8923,N_8503);
nand U9335 (N_9335,N_8573,N_8690);
xnor U9336 (N_9336,N_8824,N_8581);
nor U9337 (N_9337,N_8781,N_8666);
nand U9338 (N_9338,N_8789,N_8604);
and U9339 (N_9339,N_8563,N_8524);
and U9340 (N_9340,N_8819,N_8781);
nand U9341 (N_9341,N_8855,N_8742);
and U9342 (N_9342,N_8627,N_8807);
nor U9343 (N_9343,N_8884,N_8574);
nand U9344 (N_9344,N_8962,N_8524);
or U9345 (N_9345,N_8869,N_8529);
or U9346 (N_9346,N_8552,N_8806);
xor U9347 (N_9347,N_8548,N_8662);
xor U9348 (N_9348,N_8707,N_8926);
nor U9349 (N_9349,N_8735,N_8583);
xor U9350 (N_9350,N_8557,N_8967);
and U9351 (N_9351,N_8935,N_8548);
and U9352 (N_9352,N_8899,N_8943);
nand U9353 (N_9353,N_8717,N_8876);
nand U9354 (N_9354,N_8743,N_8832);
and U9355 (N_9355,N_8730,N_8755);
nor U9356 (N_9356,N_8628,N_8945);
xor U9357 (N_9357,N_8752,N_8717);
and U9358 (N_9358,N_8562,N_8766);
xor U9359 (N_9359,N_8672,N_8594);
xor U9360 (N_9360,N_8896,N_8898);
xnor U9361 (N_9361,N_8554,N_8694);
nor U9362 (N_9362,N_8665,N_8693);
xnor U9363 (N_9363,N_8556,N_8544);
and U9364 (N_9364,N_8767,N_8818);
and U9365 (N_9365,N_8665,N_8977);
xnor U9366 (N_9366,N_8963,N_8687);
nand U9367 (N_9367,N_8812,N_8553);
or U9368 (N_9368,N_8544,N_8616);
nor U9369 (N_9369,N_8516,N_8557);
nand U9370 (N_9370,N_8882,N_8632);
xor U9371 (N_9371,N_8652,N_8817);
nand U9372 (N_9372,N_8804,N_8869);
nor U9373 (N_9373,N_8985,N_8602);
nor U9374 (N_9374,N_8536,N_8996);
nand U9375 (N_9375,N_8578,N_8664);
nor U9376 (N_9376,N_8754,N_8739);
xor U9377 (N_9377,N_8796,N_8665);
or U9378 (N_9378,N_8584,N_8606);
nand U9379 (N_9379,N_8850,N_8813);
nor U9380 (N_9380,N_8900,N_8647);
or U9381 (N_9381,N_8975,N_8520);
nor U9382 (N_9382,N_8533,N_8790);
or U9383 (N_9383,N_8822,N_8992);
nor U9384 (N_9384,N_8844,N_8997);
and U9385 (N_9385,N_8543,N_8953);
nor U9386 (N_9386,N_8879,N_8925);
xor U9387 (N_9387,N_8572,N_8919);
nor U9388 (N_9388,N_8750,N_8508);
nor U9389 (N_9389,N_8667,N_8584);
and U9390 (N_9390,N_8721,N_8720);
xor U9391 (N_9391,N_8715,N_8956);
and U9392 (N_9392,N_8518,N_8678);
and U9393 (N_9393,N_8736,N_8946);
nor U9394 (N_9394,N_8569,N_8980);
and U9395 (N_9395,N_8852,N_8906);
and U9396 (N_9396,N_8725,N_8956);
xnor U9397 (N_9397,N_8596,N_8912);
xor U9398 (N_9398,N_8765,N_8880);
xor U9399 (N_9399,N_8851,N_8816);
or U9400 (N_9400,N_8507,N_8539);
nor U9401 (N_9401,N_8983,N_8908);
or U9402 (N_9402,N_8640,N_8534);
xor U9403 (N_9403,N_8803,N_8769);
and U9404 (N_9404,N_8815,N_8755);
and U9405 (N_9405,N_8828,N_8883);
or U9406 (N_9406,N_8908,N_8997);
nand U9407 (N_9407,N_8558,N_8889);
xnor U9408 (N_9408,N_8539,N_8700);
or U9409 (N_9409,N_8805,N_8529);
and U9410 (N_9410,N_8743,N_8736);
or U9411 (N_9411,N_8795,N_8860);
xor U9412 (N_9412,N_8838,N_8887);
nand U9413 (N_9413,N_8654,N_8713);
or U9414 (N_9414,N_8675,N_8593);
and U9415 (N_9415,N_8706,N_8984);
nand U9416 (N_9416,N_8950,N_8614);
or U9417 (N_9417,N_8959,N_8684);
nand U9418 (N_9418,N_8879,N_8680);
or U9419 (N_9419,N_8876,N_8642);
nor U9420 (N_9420,N_8987,N_8825);
nor U9421 (N_9421,N_8623,N_8834);
nor U9422 (N_9422,N_8756,N_8549);
and U9423 (N_9423,N_8989,N_8911);
and U9424 (N_9424,N_8681,N_8756);
and U9425 (N_9425,N_8671,N_8938);
or U9426 (N_9426,N_8564,N_8995);
nand U9427 (N_9427,N_8933,N_8679);
nand U9428 (N_9428,N_8955,N_8904);
or U9429 (N_9429,N_8546,N_8833);
nand U9430 (N_9430,N_8898,N_8917);
nand U9431 (N_9431,N_8887,N_8956);
nand U9432 (N_9432,N_8981,N_8863);
xnor U9433 (N_9433,N_8913,N_8594);
nor U9434 (N_9434,N_8988,N_8806);
and U9435 (N_9435,N_8838,N_8693);
nand U9436 (N_9436,N_8942,N_8597);
or U9437 (N_9437,N_8727,N_8757);
or U9438 (N_9438,N_8950,N_8975);
or U9439 (N_9439,N_8833,N_8902);
and U9440 (N_9440,N_8673,N_8749);
and U9441 (N_9441,N_8768,N_8576);
xor U9442 (N_9442,N_8967,N_8521);
and U9443 (N_9443,N_8611,N_8888);
nand U9444 (N_9444,N_8995,N_8569);
nand U9445 (N_9445,N_8738,N_8667);
and U9446 (N_9446,N_8838,N_8927);
nor U9447 (N_9447,N_8557,N_8504);
and U9448 (N_9448,N_8948,N_8846);
xnor U9449 (N_9449,N_8960,N_8521);
and U9450 (N_9450,N_8936,N_8829);
nor U9451 (N_9451,N_8811,N_8771);
nand U9452 (N_9452,N_8565,N_8944);
and U9453 (N_9453,N_8692,N_8591);
xor U9454 (N_9454,N_8608,N_8872);
or U9455 (N_9455,N_8964,N_8614);
nand U9456 (N_9456,N_8537,N_8672);
and U9457 (N_9457,N_8605,N_8767);
and U9458 (N_9458,N_8995,N_8613);
nor U9459 (N_9459,N_8641,N_8766);
xor U9460 (N_9460,N_8794,N_8987);
or U9461 (N_9461,N_8675,N_8963);
nor U9462 (N_9462,N_8568,N_8821);
nand U9463 (N_9463,N_8721,N_8593);
xor U9464 (N_9464,N_8887,N_8931);
or U9465 (N_9465,N_8553,N_8828);
or U9466 (N_9466,N_8666,N_8963);
nand U9467 (N_9467,N_8584,N_8790);
and U9468 (N_9468,N_8804,N_8620);
and U9469 (N_9469,N_8674,N_8669);
xnor U9470 (N_9470,N_8967,N_8853);
xor U9471 (N_9471,N_8577,N_8590);
nor U9472 (N_9472,N_8586,N_8974);
and U9473 (N_9473,N_8546,N_8551);
nand U9474 (N_9474,N_8842,N_8843);
nor U9475 (N_9475,N_8620,N_8712);
nor U9476 (N_9476,N_8644,N_8837);
nand U9477 (N_9477,N_8587,N_8900);
xnor U9478 (N_9478,N_8658,N_8965);
nor U9479 (N_9479,N_8950,N_8773);
or U9480 (N_9480,N_8629,N_8716);
nor U9481 (N_9481,N_8772,N_8517);
xnor U9482 (N_9482,N_8708,N_8592);
nor U9483 (N_9483,N_8953,N_8824);
or U9484 (N_9484,N_8776,N_8604);
xor U9485 (N_9485,N_8650,N_8632);
or U9486 (N_9486,N_8745,N_8596);
and U9487 (N_9487,N_8741,N_8586);
or U9488 (N_9488,N_8861,N_8997);
nand U9489 (N_9489,N_8854,N_8902);
nor U9490 (N_9490,N_8876,N_8576);
and U9491 (N_9491,N_8750,N_8509);
and U9492 (N_9492,N_8650,N_8805);
and U9493 (N_9493,N_8944,N_8698);
and U9494 (N_9494,N_8583,N_8902);
nor U9495 (N_9495,N_8545,N_8875);
nand U9496 (N_9496,N_8678,N_8896);
and U9497 (N_9497,N_8720,N_8806);
and U9498 (N_9498,N_8645,N_8649);
nor U9499 (N_9499,N_8978,N_8503);
and U9500 (N_9500,N_9322,N_9453);
xor U9501 (N_9501,N_9475,N_9058);
nand U9502 (N_9502,N_9019,N_9366);
xor U9503 (N_9503,N_9422,N_9283);
or U9504 (N_9504,N_9444,N_9212);
xor U9505 (N_9505,N_9285,N_9015);
or U9506 (N_9506,N_9070,N_9384);
xor U9507 (N_9507,N_9011,N_9448);
and U9508 (N_9508,N_9498,N_9077);
and U9509 (N_9509,N_9093,N_9338);
nor U9510 (N_9510,N_9412,N_9080);
nor U9511 (N_9511,N_9378,N_9001);
xnor U9512 (N_9512,N_9220,N_9067);
xnor U9513 (N_9513,N_9097,N_9006);
or U9514 (N_9514,N_9348,N_9180);
nand U9515 (N_9515,N_9101,N_9364);
or U9516 (N_9516,N_9167,N_9007);
nand U9517 (N_9517,N_9330,N_9194);
or U9518 (N_9518,N_9091,N_9243);
nor U9519 (N_9519,N_9290,N_9172);
nand U9520 (N_9520,N_9173,N_9151);
and U9521 (N_9521,N_9240,N_9022);
xor U9522 (N_9522,N_9195,N_9009);
or U9523 (N_9523,N_9408,N_9121);
xnor U9524 (N_9524,N_9315,N_9153);
or U9525 (N_9525,N_9239,N_9265);
and U9526 (N_9526,N_9490,N_9462);
and U9527 (N_9527,N_9276,N_9032);
and U9528 (N_9528,N_9040,N_9424);
or U9529 (N_9529,N_9487,N_9386);
and U9530 (N_9530,N_9416,N_9423);
and U9531 (N_9531,N_9041,N_9132);
or U9532 (N_9532,N_9446,N_9339);
xor U9533 (N_9533,N_9392,N_9211);
nor U9534 (N_9534,N_9217,N_9419);
or U9535 (N_9535,N_9479,N_9391);
nor U9536 (N_9536,N_9088,N_9090);
nor U9537 (N_9537,N_9385,N_9267);
xor U9538 (N_9538,N_9174,N_9254);
nor U9539 (N_9539,N_9469,N_9038);
or U9540 (N_9540,N_9439,N_9472);
or U9541 (N_9541,N_9409,N_9034);
xor U9542 (N_9542,N_9299,N_9044);
or U9543 (N_9543,N_9209,N_9154);
xor U9544 (N_9544,N_9326,N_9109);
and U9545 (N_9545,N_9181,N_9431);
nor U9546 (N_9546,N_9450,N_9141);
nor U9547 (N_9547,N_9470,N_9221);
xor U9548 (N_9548,N_9486,N_9355);
or U9549 (N_9549,N_9455,N_9036);
or U9550 (N_9550,N_9107,N_9365);
xor U9551 (N_9551,N_9345,N_9065);
or U9552 (N_9552,N_9307,N_9202);
and U9553 (N_9553,N_9237,N_9316);
and U9554 (N_9554,N_9263,N_9166);
nor U9555 (N_9555,N_9112,N_9147);
and U9556 (N_9556,N_9137,N_9157);
and U9557 (N_9557,N_9397,N_9425);
nand U9558 (N_9558,N_9351,N_9359);
nor U9559 (N_9559,N_9328,N_9466);
or U9560 (N_9560,N_9260,N_9028);
nor U9561 (N_9561,N_9200,N_9272);
xor U9562 (N_9562,N_9060,N_9131);
or U9563 (N_9563,N_9155,N_9241);
and U9564 (N_9564,N_9027,N_9465);
nand U9565 (N_9565,N_9158,N_9052);
nand U9566 (N_9566,N_9456,N_9396);
xor U9567 (N_9567,N_9269,N_9336);
nand U9568 (N_9568,N_9246,N_9075);
or U9569 (N_9569,N_9005,N_9467);
nor U9570 (N_9570,N_9324,N_9230);
xor U9571 (N_9571,N_9440,N_9306);
xor U9572 (N_9572,N_9099,N_9297);
and U9573 (N_9573,N_9128,N_9226);
xnor U9574 (N_9574,N_9102,N_9414);
nand U9575 (N_9575,N_9135,N_9062);
xor U9576 (N_9576,N_9063,N_9333);
xor U9577 (N_9577,N_9370,N_9049);
nor U9578 (N_9578,N_9301,N_9257);
and U9579 (N_9579,N_9421,N_9096);
nand U9580 (N_9580,N_9059,N_9335);
and U9581 (N_9581,N_9012,N_9054);
nor U9582 (N_9582,N_9064,N_9341);
nor U9583 (N_9583,N_9304,N_9227);
and U9584 (N_9584,N_9332,N_9494);
xor U9585 (N_9585,N_9004,N_9213);
and U9586 (N_9586,N_9327,N_9176);
nor U9587 (N_9587,N_9250,N_9106);
nor U9588 (N_9588,N_9252,N_9152);
xnor U9589 (N_9589,N_9098,N_9436);
or U9590 (N_9590,N_9206,N_9480);
nor U9591 (N_9591,N_9356,N_9282);
xor U9592 (N_9592,N_9492,N_9406);
nor U9593 (N_9593,N_9248,N_9325);
xor U9594 (N_9594,N_9134,N_9317);
xnor U9595 (N_9595,N_9183,N_9369);
or U9596 (N_9596,N_9043,N_9177);
and U9597 (N_9597,N_9346,N_9274);
nand U9598 (N_9598,N_9048,N_9125);
nor U9599 (N_9599,N_9319,N_9484);
or U9600 (N_9600,N_9160,N_9394);
and U9601 (N_9601,N_9114,N_9280);
xnor U9602 (N_9602,N_9235,N_9066);
nand U9603 (N_9603,N_9197,N_9219);
or U9604 (N_9604,N_9300,N_9100);
and U9605 (N_9605,N_9375,N_9105);
and U9606 (N_9606,N_9461,N_9008);
nor U9607 (N_9607,N_9196,N_9372);
and U9608 (N_9608,N_9228,N_9076);
or U9609 (N_9609,N_9418,N_9122);
nor U9610 (N_9610,N_9310,N_9024);
xor U9611 (N_9611,N_9496,N_9203);
and U9612 (N_9612,N_9292,N_9129);
and U9613 (N_9613,N_9377,N_9308);
nor U9614 (N_9614,N_9287,N_9441);
xor U9615 (N_9615,N_9251,N_9312);
nand U9616 (N_9616,N_9092,N_9123);
or U9617 (N_9617,N_9030,N_9020);
xnor U9618 (N_9618,N_9434,N_9204);
nor U9619 (N_9619,N_9233,N_9124);
nand U9620 (N_9620,N_9078,N_9175);
xor U9621 (N_9621,N_9072,N_9050);
nand U9622 (N_9622,N_9103,N_9061);
and U9623 (N_9623,N_9231,N_9199);
nor U9624 (N_9624,N_9383,N_9451);
nand U9625 (N_9625,N_9382,N_9089);
xnor U9626 (N_9626,N_9142,N_9162);
and U9627 (N_9627,N_9120,N_9161);
and U9628 (N_9628,N_9293,N_9340);
or U9629 (N_9629,N_9046,N_9417);
xnor U9630 (N_9630,N_9457,N_9413);
or U9631 (N_9631,N_9415,N_9139);
or U9632 (N_9632,N_9182,N_9427);
nor U9633 (N_9633,N_9373,N_9399);
nand U9634 (N_9634,N_9420,N_9463);
nand U9635 (N_9635,N_9053,N_9296);
nor U9636 (N_9636,N_9018,N_9111);
and U9637 (N_9637,N_9321,N_9284);
nor U9638 (N_9638,N_9320,N_9309);
nand U9639 (N_9639,N_9187,N_9426);
xor U9640 (N_9640,N_9170,N_9016);
nor U9641 (N_9641,N_9026,N_9144);
or U9642 (N_9642,N_9395,N_9108);
and U9643 (N_9643,N_9095,N_9482);
or U9644 (N_9644,N_9238,N_9037);
nor U9645 (N_9645,N_9491,N_9488);
nand U9646 (N_9646,N_9331,N_9130);
nand U9647 (N_9647,N_9435,N_9270);
and U9648 (N_9648,N_9318,N_9113);
nand U9649 (N_9649,N_9236,N_9010);
nand U9650 (N_9650,N_9085,N_9208);
xor U9651 (N_9651,N_9249,N_9216);
or U9652 (N_9652,N_9305,N_9387);
xor U9653 (N_9653,N_9165,N_9334);
and U9654 (N_9654,N_9357,N_9192);
or U9655 (N_9655,N_9277,N_9218);
and U9656 (N_9656,N_9074,N_9262);
nor U9657 (N_9657,N_9255,N_9082);
or U9658 (N_9658,N_9352,N_9454);
or U9659 (N_9659,N_9118,N_9485);
nor U9660 (N_9660,N_9055,N_9266);
nand U9661 (N_9661,N_9073,N_9476);
and U9662 (N_9662,N_9468,N_9127);
xor U9663 (N_9663,N_9489,N_9003);
or U9664 (N_9664,N_9405,N_9354);
or U9665 (N_9665,N_9376,N_9311);
nand U9666 (N_9666,N_9258,N_9483);
and U9667 (N_9667,N_9458,N_9140);
xnor U9668 (N_9668,N_9256,N_9362);
xnor U9669 (N_9669,N_9402,N_9302);
xor U9670 (N_9670,N_9000,N_9344);
and U9671 (N_9671,N_9403,N_9207);
xor U9672 (N_9672,N_9150,N_9433);
or U9673 (N_9673,N_9401,N_9445);
and U9674 (N_9674,N_9298,N_9164);
and U9675 (N_9675,N_9343,N_9159);
and U9676 (N_9676,N_9286,N_9013);
nor U9677 (N_9677,N_9186,N_9389);
or U9678 (N_9678,N_9149,N_9138);
or U9679 (N_9679,N_9303,N_9407);
or U9680 (N_9680,N_9393,N_9342);
or U9681 (N_9681,N_9261,N_9184);
nand U9682 (N_9682,N_9232,N_9279);
nor U9683 (N_9683,N_9079,N_9294);
nor U9684 (N_9684,N_9247,N_9400);
or U9685 (N_9685,N_9117,N_9410);
and U9686 (N_9686,N_9363,N_9259);
nor U9687 (N_9687,N_9264,N_9495);
nor U9688 (N_9688,N_9143,N_9133);
or U9689 (N_9689,N_9314,N_9337);
xnor U9690 (N_9690,N_9481,N_9452);
xor U9691 (N_9691,N_9268,N_9210);
xor U9692 (N_9692,N_9021,N_9201);
xor U9693 (N_9693,N_9358,N_9214);
xor U9694 (N_9694,N_9094,N_9477);
or U9695 (N_9695,N_9350,N_9361);
or U9696 (N_9696,N_9411,N_9493);
or U9697 (N_9697,N_9388,N_9380);
xnor U9698 (N_9698,N_9025,N_9047);
nand U9699 (N_9699,N_9273,N_9045);
nand U9700 (N_9700,N_9179,N_9190);
nand U9701 (N_9701,N_9367,N_9404);
and U9702 (N_9702,N_9432,N_9460);
or U9703 (N_9703,N_9329,N_9459);
nand U9704 (N_9704,N_9083,N_9442);
xnor U9705 (N_9705,N_9313,N_9295);
and U9706 (N_9706,N_9443,N_9437);
nor U9707 (N_9707,N_9289,N_9081);
nand U9708 (N_9708,N_9398,N_9222);
xnor U9709 (N_9709,N_9163,N_9146);
and U9710 (N_9710,N_9430,N_9205);
or U9711 (N_9711,N_9223,N_9171);
and U9712 (N_9712,N_9115,N_9449);
nor U9713 (N_9713,N_9035,N_9168);
nor U9714 (N_9714,N_9271,N_9464);
nand U9715 (N_9715,N_9374,N_9002);
or U9716 (N_9716,N_9039,N_9225);
or U9717 (N_9717,N_9447,N_9428);
nor U9718 (N_9718,N_9017,N_9242);
and U9719 (N_9719,N_9349,N_9126);
nor U9720 (N_9720,N_9368,N_9288);
nand U9721 (N_9721,N_9069,N_9244);
and U9722 (N_9722,N_9478,N_9438);
xnor U9723 (N_9723,N_9145,N_9023);
nor U9724 (N_9724,N_9390,N_9178);
nand U9725 (N_9725,N_9169,N_9185);
or U9726 (N_9726,N_9278,N_9084);
nand U9727 (N_9727,N_9371,N_9473);
and U9728 (N_9728,N_9029,N_9360);
and U9729 (N_9729,N_9474,N_9347);
and U9730 (N_9730,N_9057,N_9379);
nand U9731 (N_9731,N_9245,N_9224);
nor U9732 (N_9732,N_9253,N_9188);
xnor U9733 (N_9733,N_9042,N_9056);
nor U9734 (N_9734,N_9381,N_9353);
and U9735 (N_9735,N_9215,N_9229);
nor U9736 (N_9736,N_9110,N_9136);
nor U9737 (N_9737,N_9191,N_9119);
nor U9738 (N_9738,N_9104,N_9281);
nand U9739 (N_9739,N_9156,N_9198);
xor U9740 (N_9740,N_9068,N_9116);
nor U9741 (N_9741,N_9033,N_9193);
nand U9742 (N_9742,N_9148,N_9291);
nand U9743 (N_9743,N_9497,N_9189);
and U9744 (N_9744,N_9031,N_9429);
xor U9745 (N_9745,N_9087,N_9086);
xor U9746 (N_9746,N_9071,N_9051);
xnor U9747 (N_9747,N_9471,N_9323);
and U9748 (N_9748,N_9275,N_9499);
nand U9749 (N_9749,N_9234,N_9014);
xor U9750 (N_9750,N_9281,N_9132);
and U9751 (N_9751,N_9305,N_9386);
nand U9752 (N_9752,N_9022,N_9436);
xnor U9753 (N_9753,N_9341,N_9009);
or U9754 (N_9754,N_9284,N_9374);
xor U9755 (N_9755,N_9194,N_9251);
nand U9756 (N_9756,N_9301,N_9373);
and U9757 (N_9757,N_9256,N_9180);
and U9758 (N_9758,N_9431,N_9116);
or U9759 (N_9759,N_9289,N_9025);
and U9760 (N_9760,N_9494,N_9105);
nand U9761 (N_9761,N_9064,N_9258);
and U9762 (N_9762,N_9469,N_9182);
nand U9763 (N_9763,N_9099,N_9126);
or U9764 (N_9764,N_9102,N_9266);
and U9765 (N_9765,N_9456,N_9328);
nand U9766 (N_9766,N_9399,N_9017);
and U9767 (N_9767,N_9315,N_9140);
xnor U9768 (N_9768,N_9241,N_9164);
nor U9769 (N_9769,N_9495,N_9067);
nand U9770 (N_9770,N_9237,N_9339);
or U9771 (N_9771,N_9280,N_9314);
xnor U9772 (N_9772,N_9373,N_9237);
xor U9773 (N_9773,N_9080,N_9128);
or U9774 (N_9774,N_9353,N_9435);
xnor U9775 (N_9775,N_9374,N_9352);
xnor U9776 (N_9776,N_9171,N_9074);
nor U9777 (N_9777,N_9228,N_9001);
or U9778 (N_9778,N_9282,N_9181);
nand U9779 (N_9779,N_9483,N_9404);
nor U9780 (N_9780,N_9199,N_9090);
or U9781 (N_9781,N_9338,N_9164);
nor U9782 (N_9782,N_9398,N_9362);
or U9783 (N_9783,N_9401,N_9248);
or U9784 (N_9784,N_9041,N_9428);
or U9785 (N_9785,N_9401,N_9375);
and U9786 (N_9786,N_9345,N_9049);
nor U9787 (N_9787,N_9016,N_9206);
xnor U9788 (N_9788,N_9336,N_9310);
and U9789 (N_9789,N_9094,N_9365);
and U9790 (N_9790,N_9137,N_9384);
xor U9791 (N_9791,N_9060,N_9348);
nand U9792 (N_9792,N_9230,N_9444);
xor U9793 (N_9793,N_9436,N_9326);
nand U9794 (N_9794,N_9080,N_9315);
nand U9795 (N_9795,N_9439,N_9096);
nor U9796 (N_9796,N_9138,N_9139);
nor U9797 (N_9797,N_9353,N_9042);
and U9798 (N_9798,N_9420,N_9345);
nor U9799 (N_9799,N_9043,N_9407);
or U9800 (N_9800,N_9144,N_9400);
or U9801 (N_9801,N_9345,N_9114);
nand U9802 (N_9802,N_9341,N_9492);
and U9803 (N_9803,N_9452,N_9093);
and U9804 (N_9804,N_9024,N_9073);
nor U9805 (N_9805,N_9440,N_9406);
nand U9806 (N_9806,N_9231,N_9339);
xor U9807 (N_9807,N_9498,N_9093);
or U9808 (N_9808,N_9044,N_9032);
nor U9809 (N_9809,N_9369,N_9338);
and U9810 (N_9810,N_9313,N_9393);
and U9811 (N_9811,N_9108,N_9412);
nand U9812 (N_9812,N_9494,N_9266);
and U9813 (N_9813,N_9179,N_9278);
nor U9814 (N_9814,N_9436,N_9417);
and U9815 (N_9815,N_9000,N_9454);
nor U9816 (N_9816,N_9454,N_9314);
or U9817 (N_9817,N_9496,N_9329);
or U9818 (N_9818,N_9180,N_9253);
nor U9819 (N_9819,N_9101,N_9089);
and U9820 (N_9820,N_9496,N_9388);
and U9821 (N_9821,N_9327,N_9100);
xnor U9822 (N_9822,N_9009,N_9178);
nand U9823 (N_9823,N_9396,N_9207);
and U9824 (N_9824,N_9249,N_9156);
xor U9825 (N_9825,N_9187,N_9123);
and U9826 (N_9826,N_9150,N_9469);
and U9827 (N_9827,N_9236,N_9430);
nand U9828 (N_9828,N_9206,N_9136);
nor U9829 (N_9829,N_9074,N_9256);
or U9830 (N_9830,N_9117,N_9138);
nand U9831 (N_9831,N_9250,N_9125);
and U9832 (N_9832,N_9233,N_9390);
nand U9833 (N_9833,N_9464,N_9062);
and U9834 (N_9834,N_9491,N_9080);
and U9835 (N_9835,N_9183,N_9011);
nor U9836 (N_9836,N_9056,N_9112);
xor U9837 (N_9837,N_9039,N_9479);
nor U9838 (N_9838,N_9303,N_9414);
nand U9839 (N_9839,N_9010,N_9133);
or U9840 (N_9840,N_9075,N_9443);
nor U9841 (N_9841,N_9170,N_9480);
nand U9842 (N_9842,N_9227,N_9119);
nor U9843 (N_9843,N_9361,N_9058);
xor U9844 (N_9844,N_9254,N_9485);
and U9845 (N_9845,N_9099,N_9177);
xnor U9846 (N_9846,N_9135,N_9416);
xor U9847 (N_9847,N_9262,N_9377);
xor U9848 (N_9848,N_9193,N_9228);
nor U9849 (N_9849,N_9288,N_9345);
nor U9850 (N_9850,N_9330,N_9306);
xor U9851 (N_9851,N_9338,N_9386);
xnor U9852 (N_9852,N_9465,N_9012);
nand U9853 (N_9853,N_9498,N_9063);
nand U9854 (N_9854,N_9477,N_9276);
or U9855 (N_9855,N_9072,N_9096);
nand U9856 (N_9856,N_9134,N_9345);
nor U9857 (N_9857,N_9008,N_9084);
and U9858 (N_9858,N_9339,N_9071);
nor U9859 (N_9859,N_9467,N_9044);
nor U9860 (N_9860,N_9078,N_9088);
or U9861 (N_9861,N_9457,N_9364);
nand U9862 (N_9862,N_9256,N_9305);
nor U9863 (N_9863,N_9000,N_9112);
nand U9864 (N_9864,N_9202,N_9231);
xnor U9865 (N_9865,N_9289,N_9398);
nor U9866 (N_9866,N_9418,N_9133);
nor U9867 (N_9867,N_9114,N_9336);
xnor U9868 (N_9868,N_9323,N_9026);
nand U9869 (N_9869,N_9419,N_9236);
and U9870 (N_9870,N_9443,N_9324);
nand U9871 (N_9871,N_9337,N_9245);
nor U9872 (N_9872,N_9381,N_9072);
and U9873 (N_9873,N_9180,N_9441);
and U9874 (N_9874,N_9430,N_9488);
and U9875 (N_9875,N_9471,N_9387);
and U9876 (N_9876,N_9329,N_9374);
or U9877 (N_9877,N_9448,N_9392);
and U9878 (N_9878,N_9135,N_9437);
nor U9879 (N_9879,N_9103,N_9083);
and U9880 (N_9880,N_9047,N_9323);
xor U9881 (N_9881,N_9155,N_9084);
or U9882 (N_9882,N_9421,N_9310);
nor U9883 (N_9883,N_9110,N_9417);
nand U9884 (N_9884,N_9088,N_9051);
and U9885 (N_9885,N_9366,N_9140);
and U9886 (N_9886,N_9369,N_9196);
xnor U9887 (N_9887,N_9455,N_9078);
or U9888 (N_9888,N_9159,N_9425);
or U9889 (N_9889,N_9020,N_9289);
or U9890 (N_9890,N_9461,N_9330);
or U9891 (N_9891,N_9104,N_9314);
or U9892 (N_9892,N_9486,N_9217);
xor U9893 (N_9893,N_9431,N_9247);
or U9894 (N_9894,N_9000,N_9083);
xnor U9895 (N_9895,N_9432,N_9182);
xor U9896 (N_9896,N_9037,N_9479);
xnor U9897 (N_9897,N_9225,N_9017);
or U9898 (N_9898,N_9054,N_9436);
nor U9899 (N_9899,N_9220,N_9345);
xnor U9900 (N_9900,N_9297,N_9101);
nand U9901 (N_9901,N_9441,N_9364);
or U9902 (N_9902,N_9162,N_9149);
xnor U9903 (N_9903,N_9392,N_9345);
and U9904 (N_9904,N_9099,N_9106);
or U9905 (N_9905,N_9319,N_9196);
or U9906 (N_9906,N_9371,N_9233);
nand U9907 (N_9907,N_9089,N_9384);
nor U9908 (N_9908,N_9267,N_9441);
xor U9909 (N_9909,N_9014,N_9263);
nor U9910 (N_9910,N_9463,N_9130);
and U9911 (N_9911,N_9202,N_9109);
nand U9912 (N_9912,N_9143,N_9083);
nor U9913 (N_9913,N_9138,N_9178);
or U9914 (N_9914,N_9475,N_9319);
or U9915 (N_9915,N_9179,N_9298);
nor U9916 (N_9916,N_9258,N_9150);
and U9917 (N_9917,N_9137,N_9420);
and U9918 (N_9918,N_9290,N_9109);
nand U9919 (N_9919,N_9149,N_9072);
and U9920 (N_9920,N_9294,N_9404);
nor U9921 (N_9921,N_9449,N_9055);
xor U9922 (N_9922,N_9319,N_9401);
nor U9923 (N_9923,N_9065,N_9293);
or U9924 (N_9924,N_9442,N_9401);
or U9925 (N_9925,N_9181,N_9033);
xnor U9926 (N_9926,N_9052,N_9334);
or U9927 (N_9927,N_9456,N_9163);
nor U9928 (N_9928,N_9139,N_9436);
and U9929 (N_9929,N_9461,N_9211);
xnor U9930 (N_9930,N_9284,N_9157);
nor U9931 (N_9931,N_9017,N_9295);
nor U9932 (N_9932,N_9096,N_9430);
nand U9933 (N_9933,N_9372,N_9189);
xnor U9934 (N_9934,N_9178,N_9185);
or U9935 (N_9935,N_9186,N_9069);
and U9936 (N_9936,N_9394,N_9343);
nor U9937 (N_9937,N_9263,N_9419);
nand U9938 (N_9938,N_9480,N_9228);
or U9939 (N_9939,N_9413,N_9212);
or U9940 (N_9940,N_9212,N_9477);
or U9941 (N_9941,N_9205,N_9066);
xnor U9942 (N_9942,N_9497,N_9411);
or U9943 (N_9943,N_9086,N_9458);
nand U9944 (N_9944,N_9404,N_9062);
or U9945 (N_9945,N_9272,N_9365);
xnor U9946 (N_9946,N_9316,N_9378);
and U9947 (N_9947,N_9272,N_9463);
nor U9948 (N_9948,N_9139,N_9431);
or U9949 (N_9949,N_9411,N_9442);
nand U9950 (N_9950,N_9480,N_9219);
xnor U9951 (N_9951,N_9497,N_9117);
or U9952 (N_9952,N_9161,N_9112);
nand U9953 (N_9953,N_9465,N_9075);
or U9954 (N_9954,N_9039,N_9483);
nand U9955 (N_9955,N_9479,N_9180);
xnor U9956 (N_9956,N_9122,N_9094);
nor U9957 (N_9957,N_9110,N_9022);
nor U9958 (N_9958,N_9073,N_9010);
nor U9959 (N_9959,N_9483,N_9378);
nand U9960 (N_9960,N_9006,N_9117);
or U9961 (N_9961,N_9413,N_9344);
xnor U9962 (N_9962,N_9075,N_9043);
and U9963 (N_9963,N_9044,N_9497);
and U9964 (N_9964,N_9420,N_9414);
and U9965 (N_9965,N_9435,N_9036);
or U9966 (N_9966,N_9036,N_9021);
nand U9967 (N_9967,N_9399,N_9037);
and U9968 (N_9968,N_9282,N_9384);
nand U9969 (N_9969,N_9334,N_9021);
xnor U9970 (N_9970,N_9102,N_9416);
and U9971 (N_9971,N_9442,N_9365);
or U9972 (N_9972,N_9323,N_9385);
nand U9973 (N_9973,N_9351,N_9428);
nand U9974 (N_9974,N_9096,N_9022);
and U9975 (N_9975,N_9084,N_9484);
nand U9976 (N_9976,N_9159,N_9432);
or U9977 (N_9977,N_9499,N_9143);
and U9978 (N_9978,N_9262,N_9029);
nor U9979 (N_9979,N_9335,N_9365);
and U9980 (N_9980,N_9049,N_9399);
and U9981 (N_9981,N_9314,N_9226);
nor U9982 (N_9982,N_9452,N_9101);
or U9983 (N_9983,N_9375,N_9384);
nor U9984 (N_9984,N_9060,N_9076);
and U9985 (N_9985,N_9211,N_9288);
nand U9986 (N_9986,N_9108,N_9046);
nor U9987 (N_9987,N_9317,N_9083);
nand U9988 (N_9988,N_9352,N_9449);
nand U9989 (N_9989,N_9185,N_9414);
and U9990 (N_9990,N_9234,N_9370);
nand U9991 (N_9991,N_9247,N_9049);
nor U9992 (N_9992,N_9063,N_9218);
nand U9993 (N_9993,N_9090,N_9063);
nor U9994 (N_9994,N_9393,N_9122);
or U9995 (N_9995,N_9177,N_9335);
xor U9996 (N_9996,N_9239,N_9308);
nand U9997 (N_9997,N_9221,N_9379);
or U9998 (N_9998,N_9273,N_9455);
or U9999 (N_9999,N_9085,N_9013);
nand UO_0 (O_0,N_9568,N_9893);
nand UO_1 (O_1,N_9789,N_9942);
or UO_2 (O_2,N_9565,N_9819);
nor UO_3 (O_3,N_9556,N_9929);
nor UO_4 (O_4,N_9595,N_9676);
nand UO_5 (O_5,N_9992,N_9754);
xor UO_6 (O_6,N_9817,N_9959);
and UO_7 (O_7,N_9701,N_9896);
or UO_8 (O_8,N_9784,N_9615);
nand UO_9 (O_9,N_9545,N_9830);
or UO_10 (O_10,N_9671,N_9862);
and UO_11 (O_11,N_9639,N_9648);
xnor UO_12 (O_12,N_9696,N_9823);
xnor UO_13 (O_13,N_9650,N_9704);
or UO_14 (O_14,N_9699,N_9961);
nor UO_15 (O_15,N_9557,N_9736);
nand UO_16 (O_16,N_9620,N_9617);
and UO_17 (O_17,N_9502,N_9969);
xnor UO_18 (O_18,N_9587,N_9955);
nand UO_19 (O_19,N_9713,N_9535);
nor UO_20 (O_20,N_9803,N_9850);
nor UO_21 (O_21,N_9665,N_9619);
and UO_22 (O_22,N_9579,N_9738);
or UO_23 (O_23,N_9740,N_9814);
and UO_24 (O_24,N_9834,N_9555);
or UO_25 (O_25,N_9581,N_9885);
and UO_26 (O_26,N_9626,N_9731);
nor UO_27 (O_27,N_9614,N_9625);
and UO_28 (O_28,N_9642,N_9933);
nand UO_29 (O_29,N_9739,N_9807);
or UO_30 (O_30,N_9745,N_9646);
xor UO_31 (O_31,N_9723,N_9781);
nand UO_32 (O_32,N_9543,N_9546);
nor UO_33 (O_33,N_9981,N_9735);
or UO_34 (O_34,N_9652,N_9831);
and UO_35 (O_35,N_9726,N_9971);
xor UO_36 (O_36,N_9668,N_9763);
xnor UO_37 (O_37,N_9965,N_9944);
and UO_38 (O_38,N_9703,N_9859);
nand UO_39 (O_39,N_9629,N_9846);
xor UO_40 (O_40,N_9570,N_9957);
nand UO_41 (O_41,N_9911,N_9536);
nor UO_42 (O_42,N_9698,N_9842);
xor UO_43 (O_43,N_9963,N_9953);
or UO_44 (O_44,N_9867,N_9621);
or UO_45 (O_45,N_9907,N_9688);
or UO_46 (O_46,N_9954,N_9769);
nand UO_47 (O_47,N_9573,N_9932);
nor UO_48 (O_48,N_9529,N_9750);
nand UO_49 (O_49,N_9623,N_9572);
nand UO_50 (O_50,N_9538,N_9810);
or UO_51 (O_51,N_9506,N_9835);
nor UO_52 (O_52,N_9993,N_9649);
and UO_53 (O_53,N_9583,N_9542);
or UO_54 (O_54,N_9684,N_9998);
xor UO_55 (O_55,N_9633,N_9719);
or UO_56 (O_56,N_9990,N_9563);
or UO_57 (O_57,N_9721,N_9946);
nor UO_58 (O_58,N_9507,N_9692);
nor UO_59 (O_59,N_9999,N_9931);
and UO_60 (O_60,N_9837,N_9559);
and UO_61 (O_61,N_9611,N_9589);
nand UO_62 (O_62,N_9891,N_9966);
and UO_63 (O_63,N_9744,N_9515);
and UO_64 (O_64,N_9791,N_9972);
and UO_65 (O_65,N_9586,N_9612);
nand UO_66 (O_66,N_9662,N_9730);
xor UO_67 (O_67,N_9964,N_9947);
nand UO_68 (O_68,N_9590,N_9548);
or UO_69 (O_69,N_9805,N_9577);
nand UO_70 (O_70,N_9751,N_9934);
nor UO_71 (O_71,N_9511,N_9773);
nand UO_72 (O_72,N_9551,N_9926);
nand UO_73 (O_73,N_9657,N_9682);
or UO_74 (O_74,N_9925,N_9549);
nor UO_75 (O_75,N_9779,N_9802);
nor UO_76 (O_76,N_9674,N_9984);
and UO_77 (O_77,N_9886,N_9743);
and UO_78 (O_78,N_9895,N_9876);
or UO_79 (O_79,N_9602,N_9637);
nor UO_80 (O_80,N_9500,N_9798);
nor UO_81 (O_81,N_9788,N_9737);
and UO_82 (O_82,N_9596,N_9787);
or UO_83 (O_83,N_9613,N_9764);
nand UO_84 (O_84,N_9540,N_9974);
and UO_85 (O_85,N_9707,N_9628);
and UO_86 (O_86,N_9574,N_9917);
nor UO_87 (O_87,N_9767,N_9973);
xnor UO_88 (O_88,N_9725,N_9785);
and UO_89 (O_89,N_9811,N_9909);
or UO_90 (O_90,N_9760,N_9683);
nor UO_91 (O_91,N_9761,N_9517);
or UO_92 (O_92,N_9967,N_9575);
nand UO_93 (O_93,N_9533,N_9681);
and UO_94 (O_94,N_9913,N_9792);
and UO_95 (O_95,N_9591,N_9938);
nor UO_96 (O_96,N_9976,N_9525);
or UO_97 (O_97,N_9845,N_9605);
and UO_98 (O_98,N_9706,N_9503);
or UO_99 (O_99,N_9618,N_9797);
and UO_100 (O_100,N_9833,N_9790);
xnor UO_101 (O_101,N_9588,N_9679);
and UO_102 (O_102,N_9501,N_9853);
or UO_103 (O_103,N_9627,N_9531);
or UO_104 (O_104,N_9635,N_9943);
nor UO_105 (O_105,N_9941,N_9770);
and UO_106 (O_106,N_9912,N_9937);
nand UO_107 (O_107,N_9970,N_9765);
and UO_108 (O_108,N_9766,N_9729);
or UO_109 (O_109,N_9958,N_9844);
xor UO_110 (O_110,N_9928,N_9513);
or UO_111 (O_111,N_9658,N_9894);
nor UO_112 (O_112,N_9560,N_9554);
and UO_113 (O_113,N_9951,N_9847);
nand UO_114 (O_114,N_9801,N_9804);
nand UO_115 (O_115,N_9600,N_9888);
nor UO_116 (O_116,N_9651,N_9717);
xor UO_117 (O_117,N_9901,N_9567);
nand UO_118 (O_118,N_9910,N_9996);
nor UO_119 (O_119,N_9728,N_9660);
nand UO_120 (O_120,N_9991,N_9783);
and UO_121 (O_121,N_9510,N_9950);
nor UO_122 (O_122,N_9832,N_9860);
or UO_123 (O_123,N_9647,N_9908);
nand UO_124 (O_124,N_9848,N_9762);
nor UO_125 (O_125,N_9983,N_9768);
nand UO_126 (O_126,N_9793,N_9582);
and UO_127 (O_127,N_9936,N_9865);
nor UO_128 (O_128,N_9914,N_9697);
and UO_129 (O_129,N_9806,N_9524);
nand UO_130 (O_130,N_9708,N_9836);
nor UO_131 (O_131,N_9732,N_9906);
or UO_132 (O_132,N_9816,N_9512);
xnor UO_133 (O_133,N_9838,N_9712);
nand UO_134 (O_134,N_9576,N_9622);
and UO_135 (O_135,N_9505,N_9884);
nor UO_136 (O_136,N_9889,N_9858);
xnor UO_137 (O_137,N_9564,N_9880);
xnor UO_138 (O_138,N_9922,N_9873);
and UO_139 (O_139,N_9700,N_9630);
and UO_140 (O_140,N_9869,N_9989);
or UO_141 (O_141,N_9852,N_9636);
nand UO_142 (O_142,N_9553,N_9753);
nand UO_143 (O_143,N_9987,N_9733);
or UO_144 (O_144,N_9872,N_9718);
or UO_145 (O_145,N_9691,N_9986);
nand UO_146 (O_146,N_9571,N_9879);
xnor UO_147 (O_147,N_9638,N_9558);
nand UO_148 (O_148,N_9742,N_9851);
nor UO_149 (O_149,N_9856,N_9849);
or UO_150 (O_150,N_9669,N_9948);
and UO_151 (O_151,N_9689,N_9666);
nor UO_152 (O_152,N_9685,N_9923);
and UO_153 (O_153,N_9727,N_9566);
and UO_154 (O_154,N_9822,N_9655);
and UO_155 (O_155,N_9874,N_9710);
xor UO_156 (O_156,N_9897,N_9772);
xnor UO_157 (O_157,N_9758,N_9799);
or UO_158 (O_158,N_9599,N_9661);
or UO_159 (O_159,N_9978,N_9795);
or UO_160 (O_160,N_9827,N_9526);
or UO_161 (O_161,N_9825,N_9747);
or UO_162 (O_162,N_9949,N_9645);
or UO_163 (O_163,N_9741,N_9824);
nand UO_164 (O_164,N_9716,N_9532);
or UO_165 (O_165,N_9794,N_9550);
nand UO_166 (O_166,N_9659,N_9530);
or UO_167 (O_167,N_9552,N_9678);
and UO_168 (O_168,N_9695,N_9868);
and UO_169 (O_169,N_9919,N_9641);
nor UO_170 (O_170,N_9521,N_9654);
xor UO_171 (O_171,N_9809,N_9663);
nor UO_172 (O_172,N_9749,N_9624);
or UO_173 (O_173,N_9643,N_9634);
nand UO_174 (O_174,N_9920,N_9709);
nor UO_175 (O_175,N_9640,N_9609);
nor UO_176 (O_176,N_9687,N_9539);
and UO_177 (O_177,N_9693,N_9956);
nor UO_178 (O_178,N_9927,N_9980);
xor UO_179 (O_179,N_9939,N_9905);
or UO_180 (O_180,N_9561,N_9598);
or UO_181 (O_181,N_9601,N_9610);
and UO_182 (O_182,N_9516,N_9813);
nor UO_183 (O_183,N_9569,N_9724);
or UO_184 (O_184,N_9673,N_9690);
or UO_185 (O_185,N_9680,N_9930);
nor UO_186 (O_186,N_9714,N_9829);
xnor UO_187 (O_187,N_9776,N_9607);
nor UO_188 (O_188,N_9916,N_9962);
or UO_189 (O_189,N_9854,N_9828);
nor UO_190 (O_190,N_9997,N_9593);
nand UO_191 (O_191,N_9523,N_9757);
nand UO_192 (O_192,N_9902,N_9584);
or UO_193 (O_193,N_9544,N_9870);
nor UO_194 (O_194,N_9782,N_9715);
and UO_195 (O_195,N_9778,N_9861);
nand UO_196 (O_196,N_9866,N_9898);
nand UO_197 (O_197,N_9720,N_9924);
nand UO_198 (O_198,N_9722,N_9578);
xor UO_199 (O_199,N_9541,N_9815);
xnor UO_200 (O_200,N_9877,N_9606);
nand UO_201 (O_201,N_9608,N_9771);
and UO_202 (O_202,N_9892,N_9903);
nand UO_203 (O_203,N_9871,N_9752);
nand UO_204 (O_204,N_9780,N_9887);
xnor UO_205 (O_205,N_9520,N_9777);
and UO_206 (O_206,N_9839,N_9644);
xnor UO_207 (O_207,N_9653,N_9857);
xor UO_208 (O_208,N_9734,N_9632);
or UO_209 (O_209,N_9975,N_9960);
nor UO_210 (O_210,N_9786,N_9952);
nand UO_211 (O_211,N_9812,N_9631);
nand UO_212 (O_212,N_9821,N_9694);
nor UO_213 (O_213,N_9918,N_9664);
nor UO_214 (O_214,N_9968,N_9616);
nor UO_215 (O_215,N_9882,N_9921);
xnor UO_216 (O_216,N_9899,N_9979);
and UO_217 (O_217,N_9528,N_9840);
and UO_218 (O_218,N_9875,N_9514);
and UO_219 (O_219,N_9534,N_9748);
and UO_220 (O_220,N_9580,N_9656);
nor UO_221 (O_221,N_9820,N_9826);
or UO_222 (O_222,N_9988,N_9800);
nand UO_223 (O_223,N_9675,N_9667);
xor UO_224 (O_224,N_9547,N_9755);
nand UO_225 (O_225,N_9686,N_9518);
and UO_226 (O_226,N_9808,N_9864);
or UO_227 (O_227,N_9841,N_9603);
or UO_228 (O_228,N_9711,N_9519);
or UO_229 (O_229,N_9672,N_9843);
and UO_230 (O_230,N_9855,N_9508);
nand UO_231 (O_231,N_9818,N_9604);
xnor UO_232 (O_232,N_9759,N_9982);
and UO_233 (O_233,N_9881,N_9985);
xnor UO_234 (O_234,N_9915,N_9883);
nand UO_235 (O_235,N_9585,N_9774);
nand UO_236 (O_236,N_9670,N_9994);
nor UO_237 (O_237,N_9878,N_9863);
nand UO_238 (O_238,N_9890,N_9527);
nand UO_239 (O_239,N_9995,N_9904);
and UO_240 (O_240,N_9900,N_9977);
xnor UO_241 (O_241,N_9935,N_9504);
xor UO_242 (O_242,N_9592,N_9746);
and UO_243 (O_243,N_9940,N_9522);
nand UO_244 (O_244,N_9702,N_9705);
nor UO_245 (O_245,N_9537,N_9796);
and UO_246 (O_246,N_9756,N_9775);
xnor UO_247 (O_247,N_9597,N_9677);
or UO_248 (O_248,N_9509,N_9945);
xor UO_249 (O_249,N_9562,N_9594);
nand UO_250 (O_250,N_9978,N_9692);
nor UO_251 (O_251,N_9974,N_9638);
and UO_252 (O_252,N_9690,N_9695);
and UO_253 (O_253,N_9584,N_9726);
and UO_254 (O_254,N_9837,N_9722);
and UO_255 (O_255,N_9553,N_9988);
xor UO_256 (O_256,N_9713,N_9660);
or UO_257 (O_257,N_9995,N_9743);
nand UO_258 (O_258,N_9824,N_9725);
nor UO_259 (O_259,N_9657,N_9913);
nand UO_260 (O_260,N_9824,N_9822);
and UO_261 (O_261,N_9990,N_9826);
and UO_262 (O_262,N_9622,N_9833);
nand UO_263 (O_263,N_9674,N_9812);
and UO_264 (O_264,N_9793,N_9524);
or UO_265 (O_265,N_9877,N_9672);
xor UO_266 (O_266,N_9895,N_9608);
nor UO_267 (O_267,N_9712,N_9827);
and UO_268 (O_268,N_9699,N_9926);
nor UO_269 (O_269,N_9764,N_9536);
nor UO_270 (O_270,N_9753,N_9562);
nor UO_271 (O_271,N_9881,N_9948);
or UO_272 (O_272,N_9889,N_9654);
xor UO_273 (O_273,N_9914,N_9948);
nor UO_274 (O_274,N_9737,N_9817);
and UO_275 (O_275,N_9978,N_9788);
or UO_276 (O_276,N_9639,N_9607);
and UO_277 (O_277,N_9501,N_9902);
or UO_278 (O_278,N_9654,N_9981);
or UO_279 (O_279,N_9647,N_9530);
nand UO_280 (O_280,N_9579,N_9833);
and UO_281 (O_281,N_9797,N_9679);
nor UO_282 (O_282,N_9713,N_9942);
nor UO_283 (O_283,N_9899,N_9620);
and UO_284 (O_284,N_9641,N_9875);
nor UO_285 (O_285,N_9743,N_9827);
nand UO_286 (O_286,N_9965,N_9617);
nor UO_287 (O_287,N_9513,N_9636);
nor UO_288 (O_288,N_9502,N_9538);
nor UO_289 (O_289,N_9523,N_9937);
nand UO_290 (O_290,N_9648,N_9544);
xnor UO_291 (O_291,N_9782,N_9913);
xnor UO_292 (O_292,N_9524,N_9910);
nand UO_293 (O_293,N_9848,N_9698);
and UO_294 (O_294,N_9875,N_9555);
and UO_295 (O_295,N_9595,N_9952);
nor UO_296 (O_296,N_9733,N_9919);
xnor UO_297 (O_297,N_9645,N_9546);
nor UO_298 (O_298,N_9665,N_9852);
nand UO_299 (O_299,N_9684,N_9547);
nor UO_300 (O_300,N_9554,N_9578);
nor UO_301 (O_301,N_9641,N_9512);
and UO_302 (O_302,N_9784,N_9834);
and UO_303 (O_303,N_9974,N_9908);
nor UO_304 (O_304,N_9839,N_9840);
or UO_305 (O_305,N_9774,N_9708);
nand UO_306 (O_306,N_9522,N_9511);
xor UO_307 (O_307,N_9989,N_9539);
or UO_308 (O_308,N_9741,N_9907);
and UO_309 (O_309,N_9880,N_9590);
nor UO_310 (O_310,N_9826,N_9866);
nand UO_311 (O_311,N_9562,N_9502);
xor UO_312 (O_312,N_9796,N_9763);
nand UO_313 (O_313,N_9613,N_9967);
or UO_314 (O_314,N_9831,N_9860);
nand UO_315 (O_315,N_9927,N_9713);
nand UO_316 (O_316,N_9748,N_9820);
nor UO_317 (O_317,N_9591,N_9714);
or UO_318 (O_318,N_9944,N_9978);
or UO_319 (O_319,N_9602,N_9845);
and UO_320 (O_320,N_9906,N_9836);
nor UO_321 (O_321,N_9927,N_9510);
xnor UO_322 (O_322,N_9711,N_9506);
and UO_323 (O_323,N_9868,N_9758);
nand UO_324 (O_324,N_9660,N_9927);
or UO_325 (O_325,N_9901,N_9515);
and UO_326 (O_326,N_9551,N_9817);
nand UO_327 (O_327,N_9808,N_9989);
xnor UO_328 (O_328,N_9549,N_9851);
or UO_329 (O_329,N_9557,N_9946);
xnor UO_330 (O_330,N_9939,N_9635);
or UO_331 (O_331,N_9949,N_9827);
xnor UO_332 (O_332,N_9556,N_9954);
and UO_333 (O_333,N_9627,N_9829);
nand UO_334 (O_334,N_9565,N_9986);
xnor UO_335 (O_335,N_9638,N_9675);
nor UO_336 (O_336,N_9789,N_9818);
nand UO_337 (O_337,N_9787,N_9642);
or UO_338 (O_338,N_9691,N_9733);
or UO_339 (O_339,N_9539,N_9985);
and UO_340 (O_340,N_9663,N_9872);
or UO_341 (O_341,N_9864,N_9953);
or UO_342 (O_342,N_9794,N_9765);
and UO_343 (O_343,N_9594,N_9528);
or UO_344 (O_344,N_9987,N_9883);
nor UO_345 (O_345,N_9757,N_9520);
and UO_346 (O_346,N_9748,N_9702);
and UO_347 (O_347,N_9537,N_9555);
nor UO_348 (O_348,N_9578,N_9627);
or UO_349 (O_349,N_9820,N_9589);
xnor UO_350 (O_350,N_9908,N_9936);
nand UO_351 (O_351,N_9899,N_9826);
nor UO_352 (O_352,N_9753,N_9736);
and UO_353 (O_353,N_9692,N_9665);
nand UO_354 (O_354,N_9982,N_9987);
nor UO_355 (O_355,N_9646,N_9643);
xor UO_356 (O_356,N_9679,N_9836);
xnor UO_357 (O_357,N_9873,N_9683);
or UO_358 (O_358,N_9667,N_9789);
or UO_359 (O_359,N_9526,N_9900);
nand UO_360 (O_360,N_9977,N_9815);
nor UO_361 (O_361,N_9938,N_9652);
nor UO_362 (O_362,N_9939,N_9602);
and UO_363 (O_363,N_9795,N_9764);
and UO_364 (O_364,N_9801,N_9633);
nand UO_365 (O_365,N_9987,N_9862);
nor UO_366 (O_366,N_9696,N_9882);
xor UO_367 (O_367,N_9813,N_9862);
or UO_368 (O_368,N_9618,N_9793);
xnor UO_369 (O_369,N_9558,N_9642);
and UO_370 (O_370,N_9911,N_9943);
nand UO_371 (O_371,N_9989,N_9638);
nor UO_372 (O_372,N_9513,N_9712);
and UO_373 (O_373,N_9761,N_9924);
nand UO_374 (O_374,N_9955,N_9753);
and UO_375 (O_375,N_9596,N_9929);
or UO_376 (O_376,N_9526,N_9808);
and UO_377 (O_377,N_9882,N_9936);
xor UO_378 (O_378,N_9882,N_9537);
nor UO_379 (O_379,N_9732,N_9765);
and UO_380 (O_380,N_9586,N_9812);
xnor UO_381 (O_381,N_9648,N_9955);
nand UO_382 (O_382,N_9580,N_9909);
or UO_383 (O_383,N_9762,N_9750);
nand UO_384 (O_384,N_9705,N_9769);
or UO_385 (O_385,N_9672,N_9951);
nand UO_386 (O_386,N_9707,N_9744);
nor UO_387 (O_387,N_9884,N_9841);
nand UO_388 (O_388,N_9973,N_9997);
nand UO_389 (O_389,N_9894,N_9608);
and UO_390 (O_390,N_9997,N_9569);
nand UO_391 (O_391,N_9618,N_9892);
xnor UO_392 (O_392,N_9537,N_9540);
or UO_393 (O_393,N_9800,N_9977);
nand UO_394 (O_394,N_9748,N_9838);
or UO_395 (O_395,N_9756,N_9543);
and UO_396 (O_396,N_9509,N_9790);
xnor UO_397 (O_397,N_9740,N_9853);
nor UO_398 (O_398,N_9841,N_9820);
nand UO_399 (O_399,N_9637,N_9734);
or UO_400 (O_400,N_9901,N_9984);
nor UO_401 (O_401,N_9777,N_9705);
and UO_402 (O_402,N_9532,N_9579);
xnor UO_403 (O_403,N_9818,N_9839);
nor UO_404 (O_404,N_9725,N_9536);
nand UO_405 (O_405,N_9599,N_9512);
and UO_406 (O_406,N_9957,N_9965);
or UO_407 (O_407,N_9982,N_9652);
nor UO_408 (O_408,N_9598,N_9845);
nand UO_409 (O_409,N_9621,N_9686);
xor UO_410 (O_410,N_9842,N_9707);
xor UO_411 (O_411,N_9695,N_9883);
or UO_412 (O_412,N_9595,N_9661);
nand UO_413 (O_413,N_9570,N_9853);
nand UO_414 (O_414,N_9924,N_9641);
nand UO_415 (O_415,N_9994,N_9687);
nor UO_416 (O_416,N_9583,N_9813);
or UO_417 (O_417,N_9739,N_9651);
or UO_418 (O_418,N_9816,N_9985);
nand UO_419 (O_419,N_9971,N_9731);
or UO_420 (O_420,N_9604,N_9521);
nand UO_421 (O_421,N_9505,N_9585);
and UO_422 (O_422,N_9546,N_9639);
and UO_423 (O_423,N_9807,N_9955);
nor UO_424 (O_424,N_9974,N_9736);
nand UO_425 (O_425,N_9658,N_9981);
nor UO_426 (O_426,N_9670,N_9578);
or UO_427 (O_427,N_9894,N_9588);
nand UO_428 (O_428,N_9543,N_9880);
xor UO_429 (O_429,N_9640,N_9902);
nand UO_430 (O_430,N_9912,N_9532);
xnor UO_431 (O_431,N_9708,N_9503);
xor UO_432 (O_432,N_9916,N_9541);
or UO_433 (O_433,N_9996,N_9750);
nor UO_434 (O_434,N_9669,N_9531);
xor UO_435 (O_435,N_9647,N_9717);
nand UO_436 (O_436,N_9739,N_9732);
xor UO_437 (O_437,N_9585,N_9560);
nor UO_438 (O_438,N_9520,N_9932);
xor UO_439 (O_439,N_9702,N_9799);
xor UO_440 (O_440,N_9965,N_9565);
and UO_441 (O_441,N_9900,N_9756);
xnor UO_442 (O_442,N_9791,N_9728);
xnor UO_443 (O_443,N_9790,N_9827);
or UO_444 (O_444,N_9794,N_9698);
nand UO_445 (O_445,N_9554,N_9544);
xor UO_446 (O_446,N_9713,N_9717);
or UO_447 (O_447,N_9891,N_9997);
or UO_448 (O_448,N_9604,N_9995);
nor UO_449 (O_449,N_9912,N_9985);
or UO_450 (O_450,N_9554,N_9816);
or UO_451 (O_451,N_9769,N_9896);
or UO_452 (O_452,N_9822,N_9669);
xnor UO_453 (O_453,N_9964,N_9732);
xor UO_454 (O_454,N_9752,N_9550);
and UO_455 (O_455,N_9945,N_9902);
nand UO_456 (O_456,N_9611,N_9536);
nor UO_457 (O_457,N_9896,N_9860);
and UO_458 (O_458,N_9819,N_9930);
nand UO_459 (O_459,N_9545,N_9826);
xnor UO_460 (O_460,N_9837,N_9669);
nand UO_461 (O_461,N_9850,N_9637);
and UO_462 (O_462,N_9687,N_9575);
or UO_463 (O_463,N_9589,N_9930);
nor UO_464 (O_464,N_9521,N_9529);
nor UO_465 (O_465,N_9967,N_9881);
xor UO_466 (O_466,N_9591,N_9980);
nand UO_467 (O_467,N_9629,N_9718);
nor UO_468 (O_468,N_9734,N_9733);
nor UO_469 (O_469,N_9707,N_9909);
xor UO_470 (O_470,N_9997,N_9964);
nand UO_471 (O_471,N_9647,N_9666);
xnor UO_472 (O_472,N_9651,N_9756);
nor UO_473 (O_473,N_9689,N_9577);
or UO_474 (O_474,N_9644,N_9647);
nor UO_475 (O_475,N_9919,N_9576);
and UO_476 (O_476,N_9701,N_9992);
xnor UO_477 (O_477,N_9946,N_9686);
and UO_478 (O_478,N_9750,N_9769);
nand UO_479 (O_479,N_9707,N_9615);
nor UO_480 (O_480,N_9995,N_9783);
nor UO_481 (O_481,N_9511,N_9860);
xor UO_482 (O_482,N_9720,N_9590);
and UO_483 (O_483,N_9544,N_9933);
nor UO_484 (O_484,N_9625,N_9542);
and UO_485 (O_485,N_9834,N_9607);
xor UO_486 (O_486,N_9823,N_9772);
nand UO_487 (O_487,N_9884,N_9798);
and UO_488 (O_488,N_9773,N_9902);
nand UO_489 (O_489,N_9558,N_9591);
and UO_490 (O_490,N_9563,N_9980);
and UO_491 (O_491,N_9643,N_9570);
or UO_492 (O_492,N_9700,N_9852);
nand UO_493 (O_493,N_9540,N_9626);
and UO_494 (O_494,N_9727,N_9810);
nor UO_495 (O_495,N_9774,N_9527);
and UO_496 (O_496,N_9514,N_9741);
xor UO_497 (O_497,N_9628,N_9625);
xor UO_498 (O_498,N_9576,N_9674);
xnor UO_499 (O_499,N_9813,N_9677);
nand UO_500 (O_500,N_9847,N_9758);
nor UO_501 (O_501,N_9715,N_9803);
nand UO_502 (O_502,N_9635,N_9743);
xnor UO_503 (O_503,N_9562,N_9782);
or UO_504 (O_504,N_9691,N_9993);
nand UO_505 (O_505,N_9743,N_9772);
nand UO_506 (O_506,N_9534,N_9947);
or UO_507 (O_507,N_9552,N_9887);
or UO_508 (O_508,N_9967,N_9840);
nor UO_509 (O_509,N_9847,N_9707);
nor UO_510 (O_510,N_9555,N_9972);
nor UO_511 (O_511,N_9806,N_9730);
xnor UO_512 (O_512,N_9865,N_9709);
or UO_513 (O_513,N_9910,N_9860);
xor UO_514 (O_514,N_9768,N_9577);
or UO_515 (O_515,N_9757,N_9553);
xnor UO_516 (O_516,N_9610,N_9535);
and UO_517 (O_517,N_9608,N_9604);
and UO_518 (O_518,N_9526,N_9892);
nand UO_519 (O_519,N_9544,N_9514);
nor UO_520 (O_520,N_9670,N_9713);
and UO_521 (O_521,N_9620,N_9948);
nand UO_522 (O_522,N_9947,N_9726);
nand UO_523 (O_523,N_9731,N_9614);
and UO_524 (O_524,N_9555,N_9914);
and UO_525 (O_525,N_9775,N_9629);
nand UO_526 (O_526,N_9608,N_9927);
nor UO_527 (O_527,N_9957,N_9909);
or UO_528 (O_528,N_9825,N_9646);
xnor UO_529 (O_529,N_9684,N_9930);
nor UO_530 (O_530,N_9814,N_9566);
and UO_531 (O_531,N_9674,N_9627);
nand UO_532 (O_532,N_9993,N_9581);
nor UO_533 (O_533,N_9793,N_9542);
nor UO_534 (O_534,N_9961,N_9954);
and UO_535 (O_535,N_9709,N_9926);
and UO_536 (O_536,N_9999,N_9743);
or UO_537 (O_537,N_9684,N_9643);
nand UO_538 (O_538,N_9965,N_9980);
nor UO_539 (O_539,N_9698,N_9695);
nand UO_540 (O_540,N_9682,N_9968);
nand UO_541 (O_541,N_9743,N_9965);
nor UO_542 (O_542,N_9854,N_9839);
or UO_543 (O_543,N_9580,N_9840);
nand UO_544 (O_544,N_9732,N_9945);
or UO_545 (O_545,N_9934,N_9868);
xnor UO_546 (O_546,N_9505,N_9571);
xor UO_547 (O_547,N_9843,N_9690);
xor UO_548 (O_548,N_9940,N_9590);
nand UO_549 (O_549,N_9825,N_9560);
xnor UO_550 (O_550,N_9817,N_9519);
or UO_551 (O_551,N_9997,N_9668);
xnor UO_552 (O_552,N_9539,N_9579);
and UO_553 (O_553,N_9702,N_9605);
xnor UO_554 (O_554,N_9833,N_9772);
or UO_555 (O_555,N_9748,N_9817);
nand UO_556 (O_556,N_9735,N_9826);
nand UO_557 (O_557,N_9577,N_9720);
and UO_558 (O_558,N_9660,N_9937);
and UO_559 (O_559,N_9560,N_9623);
xnor UO_560 (O_560,N_9835,N_9744);
or UO_561 (O_561,N_9981,N_9533);
nand UO_562 (O_562,N_9754,N_9618);
and UO_563 (O_563,N_9762,N_9682);
nand UO_564 (O_564,N_9940,N_9814);
or UO_565 (O_565,N_9881,N_9563);
and UO_566 (O_566,N_9832,N_9675);
and UO_567 (O_567,N_9970,N_9646);
nand UO_568 (O_568,N_9554,N_9624);
xor UO_569 (O_569,N_9926,N_9830);
or UO_570 (O_570,N_9919,N_9948);
nand UO_571 (O_571,N_9732,N_9756);
nand UO_572 (O_572,N_9923,N_9925);
xor UO_573 (O_573,N_9584,N_9871);
nor UO_574 (O_574,N_9732,N_9901);
nand UO_575 (O_575,N_9847,N_9502);
and UO_576 (O_576,N_9763,N_9874);
xor UO_577 (O_577,N_9802,N_9891);
or UO_578 (O_578,N_9804,N_9971);
nand UO_579 (O_579,N_9925,N_9949);
or UO_580 (O_580,N_9676,N_9885);
nand UO_581 (O_581,N_9760,N_9909);
nand UO_582 (O_582,N_9595,N_9792);
xnor UO_583 (O_583,N_9711,N_9732);
xor UO_584 (O_584,N_9843,N_9893);
or UO_585 (O_585,N_9847,N_9828);
nor UO_586 (O_586,N_9740,N_9599);
nand UO_587 (O_587,N_9606,N_9861);
and UO_588 (O_588,N_9733,N_9888);
or UO_589 (O_589,N_9798,N_9644);
nand UO_590 (O_590,N_9912,N_9885);
and UO_591 (O_591,N_9586,N_9848);
xor UO_592 (O_592,N_9984,N_9709);
and UO_593 (O_593,N_9614,N_9840);
nor UO_594 (O_594,N_9506,N_9562);
nand UO_595 (O_595,N_9995,N_9795);
nand UO_596 (O_596,N_9505,N_9657);
nand UO_597 (O_597,N_9609,N_9627);
or UO_598 (O_598,N_9773,N_9637);
nand UO_599 (O_599,N_9759,N_9969);
nor UO_600 (O_600,N_9818,N_9513);
nor UO_601 (O_601,N_9545,N_9627);
and UO_602 (O_602,N_9989,N_9731);
and UO_603 (O_603,N_9580,N_9874);
xnor UO_604 (O_604,N_9782,N_9989);
xor UO_605 (O_605,N_9572,N_9987);
or UO_606 (O_606,N_9761,N_9939);
nand UO_607 (O_607,N_9639,N_9541);
and UO_608 (O_608,N_9868,N_9504);
nor UO_609 (O_609,N_9745,N_9728);
and UO_610 (O_610,N_9909,N_9601);
and UO_611 (O_611,N_9850,N_9561);
nand UO_612 (O_612,N_9610,N_9545);
and UO_613 (O_613,N_9946,N_9520);
nor UO_614 (O_614,N_9541,N_9773);
or UO_615 (O_615,N_9621,N_9733);
or UO_616 (O_616,N_9872,N_9539);
and UO_617 (O_617,N_9912,N_9603);
xor UO_618 (O_618,N_9788,N_9779);
xor UO_619 (O_619,N_9852,N_9890);
nor UO_620 (O_620,N_9964,N_9642);
xnor UO_621 (O_621,N_9799,N_9668);
nor UO_622 (O_622,N_9655,N_9629);
or UO_623 (O_623,N_9682,N_9561);
or UO_624 (O_624,N_9787,N_9601);
nand UO_625 (O_625,N_9839,N_9745);
and UO_626 (O_626,N_9848,N_9945);
nand UO_627 (O_627,N_9599,N_9574);
and UO_628 (O_628,N_9802,N_9520);
xor UO_629 (O_629,N_9654,N_9793);
nand UO_630 (O_630,N_9756,N_9645);
or UO_631 (O_631,N_9875,N_9820);
xnor UO_632 (O_632,N_9899,N_9617);
xnor UO_633 (O_633,N_9961,N_9552);
or UO_634 (O_634,N_9942,N_9733);
nor UO_635 (O_635,N_9702,N_9938);
nor UO_636 (O_636,N_9970,N_9509);
xnor UO_637 (O_637,N_9772,N_9627);
nor UO_638 (O_638,N_9973,N_9881);
nor UO_639 (O_639,N_9755,N_9706);
nand UO_640 (O_640,N_9712,N_9509);
xnor UO_641 (O_641,N_9564,N_9574);
nand UO_642 (O_642,N_9574,N_9891);
and UO_643 (O_643,N_9894,N_9825);
nand UO_644 (O_644,N_9809,N_9774);
nand UO_645 (O_645,N_9661,N_9813);
nand UO_646 (O_646,N_9821,N_9723);
nand UO_647 (O_647,N_9522,N_9970);
xnor UO_648 (O_648,N_9978,N_9704);
nand UO_649 (O_649,N_9921,N_9586);
and UO_650 (O_650,N_9789,N_9613);
xnor UO_651 (O_651,N_9984,N_9778);
or UO_652 (O_652,N_9868,N_9832);
xor UO_653 (O_653,N_9537,N_9838);
and UO_654 (O_654,N_9854,N_9638);
nand UO_655 (O_655,N_9822,N_9881);
nand UO_656 (O_656,N_9833,N_9973);
or UO_657 (O_657,N_9632,N_9783);
nor UO_658 (O_658,N_9664,N_9503);
nor UO_659 (O_659,N_9932,N_9840);
xor UO_660 (O_660,N_9673,N_9919);
xnor UO_661 (O_661,N_9831,N_9857);
nor UO_662 (O_662,N_9827,N_9866);
nand UO_663 (O_663,N_9663,N_9708);
xnor UO_664 (O_664,N_9939,N_9653);
nor UO_665 (O_665,N_9942,N_9637);
nor UO_666 (O_666,N_9921,N_9927);
or UO_667 (O_667,N_9570,N_9929);
xnor UO_668 (O_668,N_9713,N_9861);
nor UO_669 (O_669,N_9515,N_9922);
nor UO_670 (O_670,N_9565,N_9633);
and UO_671 (O_671,N_9750,N_9674);
xnor UO_672 (O_672,N_9996,N_9759);
and UO_673 (O_673,N_9914,N_9989);
nor UO_674 (O_674,N_9827,N_9551);
nor UO_675 (O_675,N_9779,N_9914);
xor UO_676 (O_676,N_9521,N_9999);
nor UO_677 (O_677,N_9634,N_9871);
xor UO_678 (O_678,N_9714,N_9824);
nand UO_679 (O_679,N_9925,N_9575);
or UO_680 (O_680,N_9908,N_9845);
xnor UO_681 (O_681,N_9883,N_9519);
and UO_682 (O_682,N_9987,N_9906);
xnor UO_683 (O_683,N_9749,N_9796);
nor UO_684 (O_684,N_9913,N_9768);
or UO_685 (O_685,N_9714,N_9652);
or UO_686 (O_686,N_9727,N_9760);
or UO_687 (O_687,N_9732,N_9517);
nand UO_688 (O_688,N_9770,N_9867);
and UO_689 (O_689,N_9944,N_9661);
nor UO_690 (O_690,N_9731,N_9860);
or UO_691 (O_691,N_9912,N_9731);
nor UO_692 (O_692,N_9630,N_9547);
nand UO_693 (O_693,N_9977,N_9648);
nand UO_694 (O_694,N_9883,N_9673);
and UO_695 (O_695,N_9852,N_9933);
nor UO_696 (O_696,N_9620,N_9720);
and UO_697 (O_697,N_9880,N_9562);
and UO_698 (O_698,N_9892,N_9801);
nor UO_699 (O_699,N_9987,N_9595);
nand UO_700 (O_700,N_9561,N_9677);
nor UO_701 (O_701,N_9880,N_9966);
and UO_702 (O_702,N_9736,N_9692);
xor UO_703 (O_703,N_9800,N_9545);
or UO_704 (O_704,N_9971,N_9875);
or UO_705 (O_705,N_9601,N_9512);
and UO_706 (O_706,N_9892,N_9852);
or UO_707 (O_707,N_9622,N_9604);
nor UO_708 (O_708,N_9630,N_9635);
or UO_709 (O_709,N_9885,N_9598);
nor UO_710 (O_710,N_9758,N_9723);
nor UO_711 (O_711,N_9815,N_9889);
or UO_712 (O_712,N_9993,N_9990);
or UO_713 (O_713,N_9791,N_9956);
xnor UO_714 (O_714,N_9550,N_9508);
nor UO_715 (O_715,N_9854,N_9591);
and UO_716 (O_716,N_9815,N_9818);
and UO_717 (O_717,N_9576,N_9753);
and UO_718 (O_718,N_9618,N_9827);
nand UO_719 (O_719,N_9660,N_9924);
or UO_720 (O_720,N_9594,N_9999);
or UO_721 (O_721,N_9832,N_9679);
and UO_722 (O_722,N_9604,N_9522);
or UO_723 (O_723,N_9940,N_9986);
and UO_724 (O_724,N_9978,N_9593);
nor UO_725 (O_725,N_9501,N_9860);
nand UO_726 (O_726,N_9618,N_9999);
and UO_727 (O_727,N_9880,N_9932);
and UO_728 (O_728,N_9919,N_9621);
or UO_729 (O_729,N_9957,N_9873);
nor UO_730 (O_730,N_9639,N_9608);
and UO_731 (O_731,N_9602,N_9679);
and UO_732 (O_732,N_9758,N_9779);
and UO_733 (O_733,N_9718,N_9792);
nor UO_734 (O_734,N_9678,N_9922);
nor UO_735 (O_735,N_9997,N_9821);
or UO_736 (O_736,N_9782,N_9672);
and UO_737 (O_737,N_9979,N_9941);
and UO_738 (O_738,N_9891,N_9878);
nor UO_739 (O_739,N_9746,N_9594);
nand UO_740 (O_740,N_9938,N_9730);
xor UO_741 (O_741,N_9751,N_9787);
nor UO_742 (O_742,N_9678,N_9788);
nor UO_743 (O_743,N_9902,N_9956);
nor UO_744 (O_744,N_9902,N_9608);
or UO_745 (O_745,N_9575,N_9670);
or UO_746 (O_746,N_9978,N_9612);
xor UO_747 (O_747,N_9701,N_9565);
and UO_748 (O_748,N_9542,N_9806);
and UO_749 (O_749,N_9544,N_9890);
xor UO_750 (O_750,N_9775,N_9813);
xnor UO_751 (O_751,N_9873,N_9723);
or UO_752 (O_752,N_9616,N_9786);
nor UO_753 (O_753,N_9963,N_9537);
nor UO_754 (O_754,N_9951,N_9721);
nor UO_755 (O_755,N_9571,N_9892);
nor UO_756 (O_756,N_9992,N_9783);
nor UO_757 (O_757,N_9735,N_9709);
nor UO_758 (O_758,N_9545,N_9749);
or UO_759 (O_759,N_9733,N_9624);
nor UO_760 (O_760,N_9742,N_9946);
xor UO_761 (O_761,N_9740,N_9704);
and UO_762 (O_762,N_9976,N_9784);
xor UO_763 (O_763,N_9750,N_9508);
or UO_764 (O_764,N_9714,N_9813);
or UO_765 (O_765,N_9642,N_9673);
nor UO_766 (O_766,N_9792,N_9600);
nor UO_767 (O_767,N_9804,N_9521);
xnor UO_768 (O_768,N_9709,N_9703);
nor UO_769 (O_769,N_9960,N_9622);
nand UO_770 (O_770,N_9913,N_9901);
xnor UO_771 (O_771,N_9946,N_9749);
nand UO_772 (O_772,N_9777,N_9889);
nand UO_773 (O_773,N_9659,N_9936);
nor UO_774 (O_774,N_9912,N_9502);
nor UO_775 (O_775,N_9773,N_9864);
xor UO_776 (O_776,N_9560,N_9702);
xnor UO_777 (O_777,N_9575,N_9524);
or UO_778 (O_778,N_9657,N_9845);
nand UO_779 (O_779,N_9538,N_9925);
xor UO_780 (O_780,N_9606,N_9675);
nor UO_781 (O_781,N_9585,N_9599);
xnor UO_782 (O_782,N_9792,N_9844);
nand UO_783 (O_783,N_9826,N_9956);
nand UO_784 (O_784,N_9729,N_9829);
and UO_785 (O_785,N_9794,N_9568);
nor UO_786 (O_786,N_9999,N_9925);
and UO_787 (O_787,N_9785,N_9531);
xnor UO_788 (O_788,N_9743,N_9650);
and UO_789 (O_789,N_9778,N_9767);
or UO_790 (O_790,N_9846,N_9765);
xnor UO_791 (O_791,N_9877,N_9534);
xnor UO_792 (O_792,N_9961,N_9897);
nand UO_793 (O_793,N_9831,N_9637);
xor UO_794 (O_794,N_9773,N_9894);
nor UO_795 (O_795,N_9533,N_9576);
and UO_796 (O_796,N_9787,N_9501);
or UO_797 (O_797,N_9748,N_9821);
nor UO_798 (O_798,N_9800,N_9924);
nand UO_799 (O_799,N_9771,N_9803);
xor UO_800 (O_800,N_9873,N_9533);
or UO_801 (O_801,N_9641,N_9622);
xnor UO_802 (O_802,N_9849,N_9770);
nor UO_803 (O_803,N_9538,N_9554);
xnor UO_804 (O_804,N_9908,N_9916);
xnor UO_805 (O_805,N_9751,N_9769);
nor UO_806 (O_806,N_9623,N_9906);
or UO_807 (O_807,N_9657,N_9835);
xor UO_808 (O_808,N_9933,N_9849);
xor UO_809 (O_809,N_9736,N_9671);
nor UO_810 (O_810,N_9771,N_9764);
and UO_811 (O_811,N_9537,N_9904);
or UO_812 (O_812,N_9830,N_9707);
nand UO_813 (O_813,N_9505,N_9982);
and UO_814 (O_814,N_9583,N_9854);
xor UO_815 (O_815,N_9921,N_9831);
xnor UO_816 (O_816,N_9878,N_9681);
nor UO_817 (O_817,N_9690,N_9779);
nor UO_818 (O_818,N_9952,N_9891);
and UO_819 (O_819,N_9744,N_9713);
nor UO_820 (O_820,N_9924,N_9810);
xor UO_821 (O_821,N_9697,N_9594);
nand UO_822 (O_822,N_9727,N_9509);
or UO_823 (O_823,N_9907,N_9549);
nor UO_824 (O_824,N_9814,N_9663);
xor UO_825 (O_825,N_9693,N_9597);
or UO_826 (O_826,N_9552,N_9860);
nor UO_827 (O_827,N_9561,N_9876);
or UO_828 (O_828,N_9936,N_9551);
xnor UO_829 (O_829,N_9948,N_9557);
or UO_830 (O_830,N_9506,N_9654);
and UO_831 (O_831,N_9632,N_9976);
nor UO_832 (O_832,N_9579,N_9549);
and UO_833 (O_833,N_9778,N_9881);
nor UO_834 (O_834,N_9593,N_9559);
and UO_835 (O_835,N_9814,N_9521);
nand UO_836 (O_836,N_9888,N_9800);
nand UO_837 (O_837,N_9684,N_9678);
or UO_838 (O_838,N_9564,N_9532);
and UO_839 (O_839,N_9823,N_9837);
nor UO_840 (O_840,N_9579,N_9754);
or UO_841 (O_841,N_9564,N_9654);
or UO_842 (O_842,N_9624,N_9993);
xnor UO_843 (O_843,N_9603,N_9666);
nor UO_844 (O_844,N_9679,N_9702);
xnor UO_845 (O_845,N_9523,N_9758);
nand UO_846 (O_846,N_9750,N_9879);
or UO_847 (O_847,N_9573,N_9995);
xor UO_848 (O_848,N_9506,N_9734);
nor UO_849 (O_849,N_9699,N_9771);
xor UO_850 (O_850,N_9562,N_9761);
and UO_851 (O_851,N_9543,N_9714);
xor UO_852 (O_852,N_9701,N_9568);
and UO_853 (O_853,N_9555,N_9892);
nand UO_854 (O_854,N_9625,N_9606);
and UO_855 (O_855,N_9941,N_9774);
xnor UO_856 (O_856,N_9646,N_9978);
xnor UO_857 (O_857,N_9889,N_9604);
and UO_858 (O_858,N_9586,N_9846);
xor UO_859 (O_859,N_9898,N_9979);
nand UO_860 (O_860,N_9541,N_9938);
or UO_861 (O_861,N_9570,N_9962);
nand UO_862 (O_862,N_9878,N_9885);
nor UO_863 (O_863,N_9741,N_9588);
nor UO_864 (O_864,N_9605,N_9626);
nor UO_865 (O_865,N_9898,N_9920);
nor UO_866 (O_866,N_9774,N_9502);
and UO_867 (O_867,N_9598,N_9523);
xnor UO_868 (O_868,N_9611,N_9621);
and UO_869 (O_869,N_9669,N_9954);
xnor UO_870 (O_870,N_9819,N_9815);
and UO_871 (O_871,N_9698,N_9889);
xor UO_872 (O_872,N_9853,N_9875);
nand UO_873 (O_873,N_9675,N_9906);
or UO_874 (O_874,N_9766,N_9902);
and UO_875 (O_875,N_9676,N_9658);
and UO_876 (O_876,N_9814,N_9619);
xnor UO_877 (O_877,N_9605,N_9802);
nor UO_878 (O_878,N_9975,N_9625);
nor UO_879 (O_879,N_9919,N_9983);
nand UO_880 (O_880,N_9989,N_9856);
and UO_881 (O_881,N_9601,N_9808);
or UO_882 (O_882,N_9846,N_9912);
nand UO_883 (O_883,N_9718,N_9809);
or UO_884 (O_884,N_9705,N_9703);
nor UO_885 (O_885,N_9697,N_9763);
nor UO_886 (O_886,N_9711,N_9671);
or UO_887 (O_887,N_9667,N_9507);
nor UO_888 (O_888,N_9833,N_9731);
nor UO_889 (O_889,N_9550,N_9728);
nor UO_890 (O_890,N_9916,N_9841);
nand UO_891 (O_891,N_9552,N_9734);
nor UO_892 (O_892,N_9847,N_9974);
nor UO_893 (O_893,N_9964,N_9725);
nor UO_894 (O_894,N_9840,N_9657);
or UO_895 (O_895,N_9769,N_9681);
or UO_896 (O_896,N_9861,N_9770);
or UO_897 (O_897,N_9638,N_9623);
xor UO_898 (O_898,N_9571,N_9990);
nand UO_899 (O_899,N_9784,N_9891);
nand UO_900 (O_900,N_9544,N_9718);
nor UO_901 (O_901,N_9560,N_9614);
or UO_902 (O_902,N_9769,N_9931);
or UO_903 (O_903,N_9971,N_9805);
nor UO_904 (O_904,N_9562,N_9503);
nor UO_905 (O_905,N_9738,N_9567);
nand UO_906 (O_906,N_9602,N_9761);
nor UO_907 (O_907,N_9662,N_9591);
or UO_908 (O_908,N_9593,N_9916);
and UO_909 (O_909,N_9623,N_9863);
nand UO_910 (O_910,N_9515,N_9646);
xor UO_911 (O_911,N_9888,N_9646);
xnor UO_912 (O_912,N_9972,N_9930);
nor UO_913 (O_913,N_9793,N_9628);
nand UO_914 (O_914,N_9552,N_9854);
or UO_915 (O_915,N_9863,N_9900);
nand UO_916 (O_916,N_9993,N_9612);
nand UO_917 (O_917,N_9605,N_9504);
and UO_918 (O_918,N_9700,N_9582);
xor UO_919 (O_919,N_9889,N_9671);
nand UO_920 (O_920,N_9733,N_9618);
or UO_921 (O_921,N_9946,N_9941);
nand UO_922 (O_922,N_9561,N_9515);
xor UO_923 (O_923,N_9836,N_9986);
or UO_924 (O_924,N_9545,N_9969);
and UO_925 (O_925,N_9824,N_9739);
nor UO_926 (O_926,N_9648,N_9810);
xnor UO_927 (O_927,N_9754,N_9907);
xor UO_928 (O_928,N_9942,N_9976);
xnor UO_929 (O_929,N_9948,N_9746);
nand UO_930 (O_930,N_9976,N_9824);
nand UO_931 (O_931,N_9890,N_9602);
and UO_932 (O_932,N_9561,N_9745);
or UO_933 (O_933,N_9946,N_9896);
nor UO_934 (O_934,N_9871,N_9788);
nand UO_935 (O_935,N_9564,N_9972);
or UO_936 (O_936,N_9711,N_9600);
and UO_937 (O_937,N_9853,N_9612);
xnor UO_938 (O_938,N_9797,N_9817);
or UO_939 (O_939,N_9561,N_9605);
and UO_940 (O_940,N_9601,N_9738);
and UO_941 (O_941,N_9764,N_9830);
nor UO_942 (O_942,N_9705,N_9719);
nor UO_943 (O_943,N_9741,N_9627);
nand UO_944 (O_944,N_9789,N_9758);
or UO_945 (O_945,N_9517,N_9692);
nand UO_946 (O_946,N_9890,N_9970);
xor UO_947 (O_947,N_9952,N_9600);
or UO_948 (O_948,N_9980,N_9544);
nand UO_949 (O_949,N_9841,N_9850);
nor UO_950 (O_950,N_9781,N_9537);
or UO_951 (O_951,N_9932,N_9675);
xnor UO_952 (O_952,N_9797,N_9870);
nor UO_953 (O_953,N_9868,N_9636);
or UO_954 (O_954,N_9890,N_9867);
or UO_955 (O_955,N_9594,N_9645);
or UO_956 (O_956,N_9722,N_9850);
nor UO_957 (O_957,N_9845,N_9731);
and UO_958 (O_958,N_9847,N_9909);
nor UO_959 (O_959,N_9846,N_9549);
nand UO_960 (O_960,N_9870,N_9818);
or UO_961 (O_961,N_9671,N_9999);
nor UO_962 (O_962,N_9714,N_9800);
and UO_963 (O_963,N_9737,N_9814);
nor UO_964 (O_964,N_9944,N_9908);
nand UO_965 (O_965,N_9891,N_9535);
xor UO_966 (O_966,N_9909,N_9895);
nor UO_967 (O_967,N_9661,N_9716);
nor UO_968 (O_968,N_9526,N_9746);
and UO_969 (O_969,N_9586,N_9666);
nand UO_970 (O_970,N_9554,N_9541);
xor UO_971 (O_971,N_9954,N_9810);
xor UO_972 (O_972,N_9994,N_9590);
and UO_973 (O_973,N_9505,N_9661);
nor UO_974 (O_974,N_9628,N_9639);
nor UO_975 (O_975,N_9598,N_9672);
nor UO_976 (O_976,N_9500,N_9503);
xor UO_977 (O_977,N_9838,N_9778);
and UO_978 (O_978,N_9556,N_9545);
or UO_979 (O_979,N_9882,N_9956);
nand UO_980 (O_980,N_9781,N_9619);
or UO_981 (O_981,N_9786,N_9529);
and UO_982 (O_982,N_9718,N_9901);
nand UO_983 (O_983,N_9826,N_9728);
or UO_984 (O_984,N_9639,N_9903);
and UO_985 (O_985,N_9920,N_9581);
or UO_986 (O_986,N_9776,N_9755);
and UO_987 (O_987,N_9814,N_9685);
nand UO_988 (O_988,N_9707,N_9915);
nand UO_989 (O_989,N_9928,N_9983);
and UO_990 (O_990,N_9745,N_9641);
and UO_991 (O_991,N_9913,N_9793);
or UO_992 (O_992,N_9758,N_9853);
nor UO_993 (O_993,N_9923,N_9607);
or UO_994 (O_994,N_9893,N_9530);
nor UO_995 (O_995,N_9571,N_9527);
nor UO_996 (O_996,N_9526,N_9671);
and UO_997 (O_997,N_9599,N_9875);
xor UO_998 (O_998,N_9991,N_9560);
or UO_999 (O_999,N_9609,N_9809);
nand UO_1000 (O_1000,N_9958,N_9562);
xnor UO_1001 (O_1001,N_9786,N_9623);
nor UO_1002 (O_1002,N_9995,N_9787);
nor UO_1003 (O_1003,N_9983,N_9680);
and UO_1004 (O_1004,N_9799,N_9683);
xnor UO_1005 (O_1005,N_9901,N_9876);
xnor UO_1006 (O_1006,N_9868,N_9941);
and UO_1007 (O_1007,N_9834,N_9529);
or UO_1008 (O_1008,N_9718,N_9609);
nand UO_1009 (O_1009,N_9638,N_9580);
or UO_1010 (O_1010,N_9759,N_9908);
and UO_1011 (O_1011,N_9936,N_9866);
xnor UO_1012 (O_1012,N_9672,N_9611);
nor UO_1013 (O_1013,N_9736,N_9547);
xnor UO_1014 (O_1014,N_9739,N_9676);
or UO_1015 (O_1015,N_9508,N_9786);
or UO_1016 (O_1016,N_9541,N_9750);
nor UO_1017 (O_1017,N_9761,N_9600);
nor UO_1018 (O_1018,N_9757,N_9996);
nor UO_1019 (O_1019,N_9776,N_9632);
xnor UO_1020 (O_1020,N_9644,N_9796);
nand UO_1021 (O_1021,N_9591,N_9636);
nand UO_1022 (O_1022,N_9673,N_9537);
and UO_1023 (O_1023,N_9871,N_9720);
or UO_1024 (O_1024,N_9715,N_9562);
nor UO_1025 (O_1025,N_9695,N_9681);
nor UO_1026 (O_1026,N_9923,N_9550);
and UO_1027 (O_1027,N_9696,N_9677);
and UO_1028 (O_1028,N_9680,N_9781);
xnor UO_1029 (O_1029,N_9506,N_9832);
or UO_1030 (O_1030,N_9839,N_9870);
and UO_1031 (O_1031,N_9603,N_9685);
nor UO_1032 (O_1032,N_9781,N_9600);
nor UO_1033 (O_1033,N_9512,N_9858);
and UO_1034 (O_1034,N_9543,N_9772);
nand UO_1035 (O_1035,N_9916,N_9535);
nor UO_1036 (O_1036,N_9547,N_9503);
nor UO_1037 (O_1037,N_9774,N_9510);
xnor UO_1038 (O_1038,N_9905,N_9953);
xor UO_1039 (O_1039,N_9742,N_9693);
and UO_1040 (O_1040,N_9607,N_9951);
xnor UO_1041 (O_1041,N_9768,N_9759);
and UO_1042 (O_1042,N_9759,N_9647);
nor UO_1043 (O_1043,N_9576,N_9732);
or UO_1044 (O_1044,N_9967,N_9752);
and UO_1045 (O_1045,N_9902,N_9704);
nand UO_1046 (O_1046,N_9606,N_9846);
nand UO_1047 (O_1047,N_9788,N_9734);
nor UO_1048 (O_1048,N_9858,N_9577);
or UO_1049 (O_1049,N_9752,N_9983);
xor UO_1050 (O_1050,N_9762,N_9519);
and UO_1051 (O_1051,N_9507,N_9788);
and UO_1052 (O_1052,N_9964,N_9752);
nand UO_1053 (O_1053,N_9763,N_9739);
or UO_1054 (O_1054,N_9698,N_9598);
nor UO_1055 (O_1055,N_9835,N_9663);
nand UO_1056 (O_1056,N_9817,N_9648);
nand UO_1057 (O_1057,N_9716,N_9515);
xnor UO_1058 (O_1058,N_9664,N_9597);
xor UO_1059 (O_1059,N_9595,N_9861);
nand UO_1060 (O_1060,N_9549,N_9928);
xnor UO_1061 (O_1061,N_9987,N_9640);
xnor UO_1062 (O_1062,N_9694,N_9895);
xor UO_1063 (O_1063,N_9997,N_9676);
xnor UO_1064 (O_1064,N_9832,N_9559);
nand UO_1065 (O_1065,N_9780,N_9738);
and UO_1066 (O_1066,N_9914,N_9865);
xnor UO_1067 (O_1067,N_9905,N_9907);
nor UO_1068 (O_1068,N_9678,N_9832);
and UO_1069 (O_1069,N_9584,N_9577);
and UO_1070 (O_1070,N_9800,N_9676);
and UO_1071 (O_1071,N_9573,N_9826);
xnor UO_1072 (O_1072,N_9872,N_9841);
xor UO_1073 (O_1073,N_9894,N_9926);
xor UO_1074 (O_1074,N_9599,N_9506);
nand UO_1075 (O_1075,N_9608,N_9720);
xnor UO_1076 (O_1076,N_9506,N_9866);
or UO_1077 (O_1077,N_9943,N_9687);
nor UO_1078 (O_1078,N_9887,N_9768);
nand UO_1079 (O_1079,N_9754,N_9749);
nand UO_1080 (O_1080,N_9806,N_9891);
or UO_1081 (O_1081,N_9894,N_9882);
xor UO_1082 (O_1082,N_9965,N_9576);
xnor UO_1083 (O_1083,N_9742,N_9521);
nor UO_1084 (O_1084,N_9988,N_9544);
and UO_1085 (O_1085,N_9976,N_9905);
xnor UO_1086 (O_1086,N_9882,N_9633);
nor UO_1087 (O_1087,N_9546,N_9946);
nor UO_1088 (O_1088,N_9631,N_9814);
xnor UO_1089 (O_1089,N_9955,N_9970);
and UO_1090 (O_1090,N_9847,N_9590);
nand UO_1091 (O_1091,N_9754,N_9839);
and UO_1092 (O_1092,N_9913,N_9639);
xor UO_1093 (O_1093,N_9523,N_9867);
and UO_1094 (O_1094,N_9537,N_9657);
nor UO_1095 (O_1095,N_9880,N_9638);
nand UO_1096 (O_1096,N_9737,N_9575);
or UO_1097 (O_1097,N_9653,N_9640);
nor UO_1098 (O_1098,N_9570,N_9793);
nor UO_1099 (O_1099,N_9941,N_9844);
nand UO_1100 (O_1100,N_9708,N_9511);
or UO_1101 (O_1101,N_9663,N_9764);
and UO_1102 (O_1102,N_9682,N_9555);
nor UO_1103 (O_1103,N_9686,N_9813);
xor UO_1104 (O_1104,N_9655,N_9590);
nand UO_1105 (O_1105,N_9689,N_9866);
xor UO_1106 (O_1106,N_9817,N_9705);
or UO_1107 (O_1107,N_9517,N_9551);
or UO_1108 (O_1108,N_9555,N_9818);
nand UO_1109 (O_1109,N_9691,N_9820);
or UO_1110 (O_1110,N_9964,N_9829);
and UO_1111 (O_1111,N_9520,N_9837);
xnor UO_1112 (O_1112,N_9663,N_9619);
xnor UO_1113 (O_1113,N_9936,N_9857);
nor UO_1114 (O_1114,N_9965,N_9816);
or UO_1115 (O_1115,N_9736,N_9942);
and UO_1116 (O_1116,N_9914,N_9690);
nand UO_1117 (O_1117,N_9956,N_9755);
and UO_1118 (O_1118,N_9535,N_9528);
nor UO_1119 (O_1119,N_9577,N_9625);
or UO_1120 (O_1120,N_9621,N_9657);
and UO_1121 (O_1121,N_9763,N_9671);
or UO_1122 (O_1122,N_9551,N_9589);
and UO_1123 (O_1123,N_9848,N_9712);
nor UO_1124 (O_1124,N_9809,N_9550);
nand UO_1125 (O_1125,N_9828,N_9565);
nand UO_1126 (O_1126,N_9570,N_9700);
xnor UO_1127 (O_1127,N_9966,N_9892);
nand UO_1128 (O_1128,N_9805,N_9763);
xnor UO_1129 (O_1129,N_9933,N_9826);
nand UO_1130 (O_1130,N_9780,N_9825);
nand UO_1131 (O_1131,N_9991,N_9785);
nor UO_1132 (O_1132,N_9542,N_9635);
nand UO_1133 (O_1133,N_9858,N_9545);
or UO_1134 (O_1134,N_9517,N_9918);
and UO_1135 (O_1135,N_9628,N_9676);
or UO_1136 (O_1136,N_9956,N_9915);
and UO_1137 (O_1137,N_9549,N_9873);
nor UO_1138 (O_1138,N_9661,N_9567);
or UO_1139 (O_1139,N_9761,N_9926);
nand UO_1140 (O_1140,N_9656,N_9595);
or UO_1141 (O_1141,N_9735,N_9578);
and UO_1142 (O_1142,N_9854,N_9988);
nand UO_1143 (O_1143,N_9607,N_9717);
nand UO_1144 (O_1144,N_9925,N_9825);
nand UO_1145 (O_1145,N_9704,N_9529);
and UO_1146 (O_1146,N_9882,N_9690);
or UO_1147 (O_1147,N_9562,N_9811);
and UO_1148 (O_1148,N_9800,N_9792);
and UO_1149 (O_1149,N_9820,N_9866);
and UO_1150 (O_1150,N_9748,N_9950);
nor UO_1151 (O_1151,N_9887,N_9653);
xor UO_1152 (O_1152,N_9930,N_9714);
and UO_1153 (O_1153,N_9829,N_9647);
nor UO_1154 (O_1154,N_9666,N_9585);
xor UO_1155 (O_1155,N_9847,N_9788);
or UO_1156 (O_1156,N_9527,N_9792);
or UO_1157 (O_1157,N_9714,N_9593);
or UO_1158 (O_1158,N_9639,N_9684);
or UO_1159 (O_1159,N_9922,N_9532);
or UO_1160 (O_1160,N_9898,N_9601);
and UO_1161 (O_1161,N_9758,N_9935);
xnor UO_1162 (O_1162,N_9985,N_9926);
and UO_1163 (O_1163,N_9694,N_9716);
or UO_1164 (O_1164,N_9870,N_9549);
nand UO_1165 (O_1165,N_9977,N_9653);
nand UO_1166 (O_1166,N_9523,N_9831);
and UO_1167 (O_1167,N_9659,N_9963);
xor UO_1168 (O_1168,N_9839,N_9580);
nor UO_1169 (O_1169,N_9730,N_9838);
and UO_1170 (O_1170,N_9756,N_9781);
and UO_1171 (O_1171,N_9571,N_9759);
or UO_1172 (O_1172,N_9674,N_9679);
nand UO_1173 (O_1173,N_9838,N_9669);
xor UO_1174 (O_1174,N_9503,N_9924);
and UO_1175 (O_1175,N_9684,N_9569);
nand UO_1176 (O_1176,N_9978,N_9676);
nand UO_1177 (O_1177,N_9667,N_9811);
or UO_1178 (O_1178,N_9823,N_9939);
nand UO_1179 (O_1179,N_9521,N_9613);
xnor UO_1180 (O_1180,N_9835,N_9575);
nor UO_1181 (O_1181,N_9880,N_9550);
xor UO_1182 (O_1182,N_9876,N_9589);
or UO_1183 (O_1183,N_9676,N_9867);
and UO_1184 (O_1184,N_9627,N_9933);
nor UO_1185 (O_1185,N_9839,N_9582);
nand UO_1186 (O_1186,N_9720,N_9741);
nand UO_1187 (O_1187,N_9798,N_9719);
and UO_1188 (O_1188,N_9578,N_9816);
nand UO_1189 (O_1189,N_9527,N_9813);
nor UO_1190 (O_1190,N_9937,N_9983);
nor UO_1191 (O_1191,N_9648,N_9880);
xnor UO_1192 (O_1192,N_9531,N_9953);
xnor UO_1193 (O_1193,N_9887,N_9594);
and UO_1194 (O_1194,N_9811,N_9669);
and UO_1195 (O_1195,N_9749,N_9858);
and UO_1196 (O_1196,N_9801,N_9550);
or UO_1197 (O_1197,N_9500,N_9690);
nand UO_1198 (O_1198,N_9727,N_9807);
or UO_1199 (O_1199,N_9932,N_9541);
nor UO_1200 (O_1200,N_9892,N_9979);
nand UO_1201 (O_1201,N_9733,N_9511);
nand UO_1202 (O_1202,N_9792,N_9736);
and UO_1203 (O_1203,N_9501,N_9834);
nand UO_1204 (O_1204,N_9590,N_9633);
and UO_1205 (O_1205,N_9524,N_9750);
nor UO_1206 (O_1206,N_9561,N_9734);
nand UO_1207 (O_1207,N_9972,N_9768);
nand UO_1208 (O_1208,N_9852,N_9821);
nor UO_1209 (O_1209,N_9532,N_9979);
xnor UO_1210 (O_1210,N_9604,N_9901);
nand UO_1211 (O_1211,N_9704,N_9526);
nor UO_1212 (O_1212,N_9541,N_9842);
nor UO_1213 (O_1213,N_9695,N_9667);
xnor UO_1214 (O_1214,N_9512,N_9883);
and UO_1215 (O_1215,N_9877,N_9759);
xnor UO_1216 (O_1216,N_9860,N_9986);
nand UO_1217 (O_1217,N_9918,N_9628);
and UO_1218 (O_1218,N_9660,N_9678);
nor UO_1219 (O_1219,N_9946,N_9558);
xnor UO_1220 (O_1220,N_9743,N_9785);
nand UO_1221 (O_1221,N_9742,N_9779);
and UO_1222 (O_1222,N_9546,N_9694);
and UO_1223 (O_1223,N_9779,N_9698);
nand UO_1224 (O_1224,N_9863,N_9685);
nor UO_1225 (O_1225,N_9668,N_9907);
nor UO_1226 (O_1226,N_9637,N_9677);
and UO_1227 (O_1227,N_9832,N_9568);
nand UO_1228 (O_1228,N_9738,N_9669);
nand UO_1229 (O_1229,N_9598,N_9766);
nor UO_1230 (O_1230,N_9842,N_9710);
or UO_1231 (O_1231,N_9632,N_9801);
xnor UO_1232 (O_1232,N_9860,N_9962);
or UO_1233 (O_1233,N_9799,N_9894);
or UO_1234 (O_1234,N_9560,N_9514);
xnor UO_1235 (O_1235,N_9726,N_9725);
xnor UO_1236 (O_1236,N_9688,N_9779);
or UO_1237 (O_1237,N_9742,N_9765);
nand UO_1238 (O_1238,N_9605,N_9925);
xor UO_1239 (O_1239,N_9734,N_9652);
nand UO_1240 (O_1240,N_9853,N_9784);
nor UO_1241 (O_1241,N_9624,N_9668);
and UO_1242 (O_1242,N_9953,N_9964);
nand UO_1243 (O_1243,N_9598,N_9659);
xnor UO_1244 (O_1244,N_9523,N_9555);
nand UO_1245 (O_1245,N_9570,N_9725);
and UO_1246 (O_1246,N_9882,N_9657);
xor UO_1247 (O_1247,N_9650,N_9628);
nor UO_1248 (O_1248,N_9893,N_9697);
xor UO_1249 (O_1249,N_9818,N_9771);
nor UO_1250 (O_1250,N_9575,N_9614);
nor UO_1251 (O_1251,N_9651,N_9705);
nor UO_1252 (O_1252,N_9996,N_9870);
and UO_1253 (O_1253,N_9917,N_9612);
and UO_1254 (O_1254,N_9585,N_9629);
or UO_1255 (O_1255,N_9900,N_9568);
xor UO_1256 (O_1256,N_9667,N_9897);
or UO_1257 (O_1257,N_9698,N_9934);
nor UO_1258 (O_1258,N_9773,N_9912);
and UO_1259 (O_1259,N_9967,N_9779);
nor UO_1260 (O_1260,N_9584,N_9564);
nand UO_1261 (O_1261,N_9891,N_9664);
or UO_1262 (O_1262,N_9879,N_9547);
xor UO_1263 (O_1263,N_9578,N_9522);
nand UO_1264 (O_1264,N_9507,N_9693);
nand UO_1265 (O_1265,N_9693,N_9504);
or UO_1266 (O_1266,N_9935,N_9661);
and UO_1267 (O_1267,N_9551,N_9686);
and UO_1268 (O_1268,N_9737,N_9608);
and UO_1269 (O_1269,N_9787,N_9774);
nor UO_1270 (O_1270,N_9605,N_9785);
or UO_1271 (O_1271,N_9557,N_9937);
nand UO_1272 (O_1272,N_9866,N_9615);
and UO_1273 (O_1273,N_9521,N_9915);
or UO_1274 (O_1274,N_9941,N_9570);
nor UO_1275 (O_1275,N_9782,N_9970);
nand UO_1276 (O_1276,N_9820,N_9814);
and UO_1277 (O_1277,N_9656,N_9558);
or UO_1278 (O_1278,N_9937,N_9847);
nand UO_1279 (O_1279,N_9714,N_9844);
xor UO_1280 (O_1280,N_9617,N_9901);
xor UO_1281 (O_1281,N_9978,N_9754);
nor UO_1282 (O_1282,N_9745,N_9922);
xnor UO_1283 (O_1283,N_9624,N_9900);
xor UO_1284 (O_1284,N_9914,N_9571);
nor UO_1285 (O_1285,N_9595,N_9818);
and UO_1286 (O_1286,N_9925,N_9820);
nand UO_1287 (O_1287,N_9949,N_9636);
xor UO_1288 (O_1288,N_9705,N_9963);
or UO_1289 (O_1289,N_9838,N_9552);
nand UO_1290 (O_1290,N_9823,N_9687);
or UO_1291 (O_1291,N_9534,N_9692);
nor UO_1292 (O_1292,N_9850,N_9963);
nand UO_1293 (O_1293,N_9643,N_9561);
or UO_1294 (O_1294,N_9744,N_9689);
nand UO_1295 (O_1295,N_9625,N_9897);
and UO_1296 (O_1296,N_9668,N_9747);
and UO_1297 (O_1297,N_9776,N_9544);
and UO_1298 (O_1298,N_9597,N_9864);
and UO_1299 (O_1299,N_9779,N_9541);
nor UO_1300 (O_1300,N_9997,N_9557);
and UO_1301 (O_1301,N_9683,N_9907);
and UO_1302 (O_1302,N_9700,N_9808);
nor UO_1303 (O_1303,N_9606,N_9542);
xnor UO_1304 (O_1304,N_9787,N_9718);
nand UO_1305 (O_1305,N_9756,N_9888);
nand UO_1306 (O_1306,N_9780,N_9537);
and UO_1307 (O_1307,N_9603,N_9830);
xor UO_1308 (O_1308,N_9795,N_9724);
nand UO_1309 (O_1309,N_9661,N_9517);
or UO_1310 (O_1310,N_9568,N_9928);
nor UO_1311 (O_1311,N_9709,N_9625);
or UO_1312 (O_1312,N_9529,N_9623);
and UO_1313 (O_1313,N_9798,N_9710);
and UO_1314 (O_1314,N_9786,N_9900);
and UO_1315 (O_1315,N_9580,N_9670);
nor UO_1316 (O_1316,N_9742,N_9808);
and UO_1317 (O_1317,N_9801,N_9674);
and UO_1318 (O_1318,N_9607,N_9914);
and UO_1319 (O_1319,N_9903,N_9910);
xnor UO_1320 (O_1320,N_9509,N_9824);
and UO_1321 (O_1321,N_9629,N_9706);
or UO_1322 (O_1322,N_9809,N_9798);
nand UO_1323 (O_1323,N_9625,N_9626);
nor UO_1324 (O_1324,N_9564,N_9891);
or UO_1325 (O_1325,N_9753,N_9693);
nor UO_1326 (O_1326,N_9591,N_9976);
or UO_1327 (O_1327,N_9928,N_9639);
and UO_1328 (O_1328,N_9954,N_9994);
nand UO_1329 (O_1329,N_9797,N_9787);
nand UO_1330 (O_1330,N_9771,N_9576);
or UO_1331 (O_1331,N_9700,N_9705);
nor UO_1332 (O_1332,N_9904,N_9524);
nor UO_1333 (O_1333,N_9712,N_9556);
nand UO_1334 (O_1334,N_9512,N_9645);
nor UO_1335 (O_1335,N_9804,N_9579);
or UO_1336 (O_1336,N_9915,N_9535);
xor UO_1337 (O_1337,N_9535,N_9521);
nand UO_1338 (O_1338,N_9689,N_9782);
nand UO_1339 (O_1339,N_9825,N_9602);
and UO_1340 (O_1340,N_9763,N_9598);
or UO_1341 (O_1341,N_9834,N_9666);
and UO_1342 (O_1342,N_9513,N_9989);
and UO_1343 (O_1343,N_9586,N_9506);
or UO_1344 (O_1344,N_9736,N_9921);
or UO_1345 (O_1345,N_9608,N_9664);
and UO_1346 (O_1346,N_9854,N_9933);
xnor UO_1347 (O_1347,N_9951,N_9784);
or UO_1348 (O_1348,N_9666,N_9571);
and UO_1349 (O_1349,N_9544,N_9688);
nor UO_1350 (O_1350,N_9633,N_9761);
or UO_1351 (O_1351,N_9541,N_9678);
or UO_1352 (O_1352,N_9641,N_9964);
nor UO_1353 (O_1353,N_9592,N_9575);
nand UO_1354 (O_1354,N_9573,N_9769);
and UO_1355 (O_1355,N_9509,N_9904);
xor UO_1356 (O_1356,N_9721,N_9720);
and UO_1357 (O_1357,N_9830,N_9698);
xnor UO_1358 (O_1358,N_9509,N_9633);
and UO_1359 (O_1359,N_9826,N_9932);
nand UO_1360 (O_1360,N_9872,N_9903);
or UO_1361 (O_1361,N_9978,N_9991);
or UO_1362 (O_1362,N_9923,N_9527);
nor UO_1363 (O_1363,N_9958,N_9735);
nand UO_1364 (O_1364,N_9731,N_9862);
xor UO_1365 (O_1365,N_9820,N_9732);
or UO_1366 (O_1366,N_9520,N_9753);
nor UO_1367 (O_1367,N_9548,N_9514);
or UO_1368 (O_1368,N_9647,N_9735);
nand UO_1369 (O_1369,N_9534,N_9932);
or UO_1370 (O_1370,N_9787,N_9591);
nand UO_1371 (O_1371,N_9597,N_9512);
xnor UO_1372 (O_1372,N_9803,N_9553);
xor UO_1373 (O_1373,N_9944,N_9982);
nand UO_1374 (O_1374,N_9989,N_9628);
xor UO_1375 (O_1375,N_9611,N_9690);
nor UO_1376 (O_1376,N_9957,N_9779);
and UO_1377 (O_1377,N_9519,N_9695);
nand UO_1378 (O_1378,N_9509,N_9521);
xor UO_1379 (O_1379,N_9704,N_9826);
and UO_1380 (O_1380,N_9639,N_9617);
or UO_1381 (O_1381,N_9923,N_9880);
and UO_1382 (O_1382,N_9631,N_9752);
or UO_1383 (O_1383,N_9514,N_9554);
xnor UO_1384 (O_1384,N_9840,N_9675);
nor UO_1385 (O_1385,N_9542,N_9678);
nand UO_1386 (O_1386,N_9934,N_9617);
and UO_1387 (O_1387,N_9539,N_9536);
xor UO_1388 (O_1388,N_9694,N_9800);
and UO_1389 (O_1389,N_9849,N_9785);
and UO_1390 (O_1390,N_9932,N_9753);
xnor UO_1391 (O_1391,N_9669,N_9706);
nand UO_1392 (O_1392,N_9808,N_9790);
nor UO_1393 (O_1393,N_9746,N_9755);
xor UO_1394 (O_1394,N_9610,N_9626);
and UO_1395 (O_1395,N_9877,N_9950);
nand UO_1396 (O_1396,N_9588,N_9560);
and UO_1397 (O_1397,N_9762,N_9899);
and UO_1398 (O_1398,N_9833,N_9805);
xor UO_1399 (O_1399,N_9706,N_9765);
nand UO_1400 (O_1400,N_9955,N_9568);
xor UO_1401 (O_1401,N_9922,N_9516);
xor UO_1402 (O_1402,N_9568,N_9770);
or UO_1403 (O_1403,N_9666,N_9782);
nor UO_1404 (O_1404,N_9772,N_9685);
xnor UO_1405 (O_1405,N_9586,N_9830);
nor UO_1406 (O_1406,N_9947,N_9722);
nand UO_1407 (O_1407,N_9904,N_9902);
or UO_1408 (O_1408,N_9803,N_9867);
xnor UO_1409 (O_1409,N_9574,N_9554);
and UO_1410 (O_1410,N_9868,N_9667);
xnor UO_1411 (O_1411,N_9841,N_9614);
and UO_1412 (O_1412,N_9869,N_9808);
nand UO_1413 (O_1413,N_9843,N_9709);
or UO_1414 (O_1414,N_9997,N_9693);
nor UO_1415 (O_1415,N_9846,N_9696);
and UO_1416 (O_1416,N_9782,N_9968);
nand UO_1417 (O_1417,N_9709,N_9866);
nand UO_1418 (O_1418,N_9871,N_9632);
nand UO_1419 (O_1419,N_9508,N_9682);
xor UO_1420 (O_1420,N_9779,N_9909);
and UO_1421 (O_1421,N_9963,N_9649);
nor UO_1422 (O_1422,N_9873,N_9516);
and UO_1423 (O_1423,N_9722,N_9729);
or UO_1424 (O_1424,N_9997,N_9827);
xnor UO_1425 (O_1425,N_9690,N_9903);
xor UO_1426 (O_1426,N_9543,N_9697);
and UO_1427 (O_1427,N_9672,N_9871);
xor UO_1428 (O_1428,N_9508,N_9987);
nor UO_1429 (O_1429,N_9671,N_9970);
nor UO_1430 (O_1430,N_9510,N_9980);
nor UO_1431 (O_1431,N_9545,N_9856);
nand UO_1432 (O_1432,N_9521,N_9568);
nor UO_1433 (O_1433,N_9886,N_9918);
xor UO_1434 (O_1434,N_9907,N_9544);
nand UO_1435 (O_1435,N_9605,N_9552);
or UO_1436 (O_1436,N_9904,N_9597);
nor UO_1437 (O_1437,N_9693,N_9685);
nand UO_1438 (O_1438,N_9797,N_9783);
xnor UO_1439 (O_1439,N_9920,N_9938);
nand UO_1440 (O_1440,N_9957,N_9513);
and UO_1441 (O_1441,N_9901,N_9747);
nor UO_1442 (O_1442,N_9824,N_9761);
nor UO_1443 (O_1443,N_9783,N_9929);
or UO_1444 (O_1444,N_9995,N_9785);
or UO_1445 (O_1445,N_9861,N_9873);
or UO_1446 (O_1446,N_9959,N_9695);
nand UO_1447 (O_1447,N_9922,N_9916);
and UO_1448 (O_1448,N_9859,N_9961);
nor UO_1449 (O_1449,N_9895,N_9922);
nand UO_1450 (O_1450,N_9719,N_9858);
nand UO_1451 (O_1451,N_9583,N_9983);
nand UO_1452 (O_1452,N_9962,N_9536);
and UO_1453 (O_1453,N_9574,N_9749);
or UO_1454 (O_1454,N_9888,N_9637);
or UO_1455 (O_1455,N_9786,N_9609);
or UO_1456 (O_1456,N_9753,N_9709);
or UO_1457 (O_1457,N_9533,N_9575);
and UO_1458 (O_1458,N_9701,N_9934);
xor UO_1459 (O_1459,N_9582,N_9778);
and UO_1460 (O_1460,N_9862,N_9531);
xor UO_1461 (O_1461,N_9889,N_9748);
and UO_1462 (O_1462,N_9971,N_9538);
xor UO_1463 (O_1463,N_9998,N_9590);
nand UO_1464 (O_1464,N_9791,N_9836);
nor UO_1465 (O_1465,N_9805,N_9520);
xor UO_1466 (O_1466,N_9500,N_9532);
nand UO_1467 (O_1467,N_9840,N_9622);
nand UO_1468 (O_1468,N_9515,N_9577);
nand UO_1469 (O_1469,N_9672,N_9623);
or UO_1470 (O_1470,N_9557,N_9819);
xnor UO_1471 (O_1471,N_9637,N_9991);
nor UO_1472 (O_1472,N_9874,N_9792);
xor UO_1473 (O_1473,N_9760,N_9710);
xor UO_1474 (O_1474,N_9813,N_9704);
xnor UO_1475 (O_1475,N_9858,N_9554);
nor UO_1476 (O_1476,N_9664,N_9901);
or UO_1477 (O_1477,N_9553,N_9659);
or UO_1478 (O_1478,N_9535,N_9613);
or UO_1479 (O_1479,N_9649,N_9717);
nand UO_1480 (O_1480,N_9840,N_9736);
and UO_1481 (O_1481,N_9853,N_9556);
nor UO_1482 (O_1482,N_9751,N_9591);
xor UO_1483 (O_1483,N_9881,N_9909);
nand UO_1484 (O_1484,N_9564,N_9608);
nand UO_1485 (O_1485,N_9585,N_9661);
or UO_1486 (O_1486,N_9791,N_9714);
nor UO_1487 (O_1487,N_9919,N_9566);
nand UO_1488 (O_1488,N_9866,N_9851);
nor UO_1489 (O_1489,N_9742,N_9892);
or UO_1490 (O_1490,N_9698,N_9766);
xor UO_1491 (O_1491,N_9604,N_9772);
nand UO_1492 (O_1492,N_9765,N_9945);
xnor UO_1493 (O_1493,N_9688,N_9754);
or UO_1494 (O_1494,N_9899,N_9978);
and UO_1495 (O_1495,N_9565,N_9967);
or UO_1496 (O_1496,N_9856,N_9995);
xnor UO_1497 (O_1497,N_9505,N_9752);
nor UO_1498 (O_1498,N_9808,N_9586);
nand UO_1499 (O_1499,N_9841,N_9868);
endmodule