module basic_1000_10000_1500_20_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_296,In_176);
or U1 (N_1,In_792,In_286);
or U2 (N_2,In_518,In_449);
and U3 (N_3,In_23,In_260);
nor U4 (N_4,In_890,In_558);
and U5 (N_5,In_227,In_95);
or U6 (N_6,In_240,In_880);
nand U7 (N_7,In_212,In_363);
nor U8 (N_8,In_503,In_840);
or U9 (N_9,In_771,In_366);
and U10 (N_10,In_443,In_780);
nor U11 (N_11,In_610,In_859);
and U12 (N_12,In_330,In_837);
or U13 (N_13,In_469,In_399);
and U14 (N_14,In_949,In_321);
and U15 (N_15,In_101,In_854);
nor U16 (N_16,In_957,In_373);
xnor U17 (N_17,In_672,In_462);
nor U18 (N_18,In_965,In_257);
and U19 (N_19,In_579,In_109);
and U20 (N_20,In_812,In_842);
nand U21 (N_21,In_698,In_261);
or U22 (N_22,In_285,In_265);
nand U23 (N_23,In_552,In_828);
or U24 (N_24,In_487,In_270);
or U25 (N_25,In_216,In_700);
nor U26 (N_26,In_678,In_565);
nand U27 (N_27,In_543,In_488);
nand U28 (N_28,In_375,In_675);
nand U29 (N_29,In_279,In_703);
nand U30 (N_30,In_184,In_929);
or U31 (N_31,In_605,In_20);
and U32 (N_32,In_519,In_422);
and U33 (N_33,In_343,In_676);
nor U34 (N_34,In_102,In_355);
nand U35 (N_35,In_215,In_453);
nand U36 (N_36,In_458,In_909);
and U37 (N_37,In_657,In_421);
or U38 (N_38,In_968,In_262);
and U39 (N_39,In_960,In_747);
or U40 (N_40,In_434,In_540);
or U41 (N_41,In_685,In_522);
nand U42 (N_42,In_951,In_902);
nor U43 (N_43,In_602,In_74);
and U44 (N_44,In_199,In_819);
nand U45 (N_45,In_441,In_148);
and U46 (N_46,In_1,In_695);
and U47 (N_47,In_710,In_759);
nand U48 (N_48,In_614,In_752);
or U49 (N_49,In_903,In_244);
nand U50 (N_50,In_40,In_997);
or U51 (N_51,In_353,In_91);
nor U52 (N_52,In_895,In_418);
nand U53 (N_53,In_641,In_581);
nand U54 (N_54,In_745,In_735);
and U55 (N_55,In_674,In_495);
nand U56 (N_56,In_996,In_527);
nand U57 (N_57,In_654,In_222);
and U58 (N_58,In_966,In_106);
and U59 (N_59,In_599,In_410);
nor U60 (N_60,In_162,In_437);
nor U61 (N_61,In_19,In_165);
nand U62 (N_62,In_457,In_755);
nor U63 (N_63,In_790,In_801);
nand U64 (N_64,In_838,In_728);
or U65 (N_65,In_175,In_750);
nor U66 (N_66,In_653,In_535);
nor U67 (N_67,In_17,In_897);
nor U68 (N_68,In_389,In_390);
and U69 (N_69,In_636,In_200);
xor U70 (N_70,In_133,In_228);
nor U71 (N_71,In_100,In_513);
nand U72 (N_72,In_928,In_303);
and U73 (N_73,In_797,In_746);
nand U74 (N_74,In_911,In_971);
or U75 (N_75,In_907,In_651);
nand U76 (N_76,In_119,In_937);
and U77 (N_77,In_379,In_368);
and U78 (N_78,In_584,In_575);
and U79 (N_79,In_712,In_736);
or U80 (N_80,In_901,In_939);
or U81 (N_81,In_409,In_476);
nor U82 (N_82,In_888,In_22);
nand U83 (N_83,In_271,In_521);
nor U84 (N_84,In_510,In_11);
or U85 (N_85,In_655,In_740);
nand U86 (N_86,In_696,In_941);
and U87 (N_87,In_727,In_826);
or U88 (N_88,In_440,In_174);
nor U89 (N_89,In_258,In_652);
nor U90 (N_90,In_58,In_130);
or U91 (N_91,In_294,In_423);
and U92 (N_92,In_638,In_841);
nand U93 (N_93,In_961,In_977);
nor U94 (N_94,In_874,In_63);
or U95 (N_95,In_810,In_336);
or U96 (N_96,In_482,In_239);
and U97 (N_97,In_537,In_549);
or U98 (N_98,In_196,In_405);
and U99 (N_99,In_591,In_255);
nor U100 (N_100,In_640,In_96);
nand U101 (N_101,In_892,In_26);
and U102 (N_102,In_4,In_129);
and U103 (N_103,In_592,In_154);
and U104 (N_104,In_808,In_10);
nand U105 (N_105,In_626,In_8);
nor U106 (N_106,In_974,In_548);
nor U107 (N_107,In_427,In_145);
or U108 (N_108,In_166,In_182);
nor U109 (N_109,In_97,In_147);
xor U110 (N_110,In_112,In_406);
xnor U111 (N_111,In_172,In_71);
and U112 (N_112,In_304,In_217);
nor U113 (N_113,In_35,In_77);
nor U114 (N_114,In_231,In_501);
nand U115 (N_115,In_291,In_822);
and U116 (N_116,In_55,In_875);
or U117 (N_117,In_551,In_992);
nor U118 (N_118,In_480,In_531);
nand U119 (N_119,In_936,In_944);
or U120 (N_120,In_690,In_699);
or U121 (N_121,In_734,In_138);
nor U122 (N_122,In_542,In_791);
nor U123 (N_123,In_75,In_357);
or U124 (N_124,In_871,In_621);
nand U125 (N_125,In_319,In_65);
or U126 (N_126,In_673,In_436);
nand U127 (N_127,In_221,In_984);
xor U128 (N_128,In_191,In_397);
or U129 (N_129,In_724,In_39);
nor U130 (N_130,In_802,In_135);
nand U131 (N_131,In_149,In_416);
and U132 (N_132,In_985,In_297);
nor U133 (N_133,In_447,In_232);
and U134 (N_134,In_624,In_364);
and U135 (N_135,In_254,In_253);
or U136 (N_136,In_940,In_34);
or U137 (N_137,In_720,In_702);
nor U138 (N_138,In_391,In_594);
nand U139 (N_139,In_497,In_793);
nor U140 (N_140,In_205,In_387);
or U141 (N_141,In_586,In_511);
nand U142 (N_142,In_134,In_692);
nor U143 (N_143,In_386,In_408);
and U144 (N_144,In_33,In_276);
nor U145 (N_145,In_952,In_814);
nor U146 (N_146,In_224,In_546);
and U147 (N_147,In_648,In_123);
and U148 (N_148,In_632,In_889);
nor U149 (N_149,In_25,In_852);
and U150 (N_150,In_128,In_432);
and U151 (N_151,In_629,In_878);
or U152 (N_152,In_798,In_744);
and U153 (N_153,In_66,In_248);
and U154 (N_154,In_243,In_915);
and U155 (N_155,In_318,In_668);
and U156 (N_156,In_807,In_472);
xor U157 (N_157,In_464,In_47);
or U158 (N_158,In_588,In_721);
nor U159 (N_159,In_316,In_933);
nor U160 (N_160,In_836,In_557);
nor U161 (N_161,In_496,In_282);
nor U162 (N_162,In_99,In_956);
nand U163 (N_163,In_351,In_555);
or U164 (N_164,In_980,In_656);
and U165 (N_165,In_990,In_438);
nor U166 (N_166,In_796,In_385);
nor U167 (N_167,In_446,In_693);
or U168 (N_168,In_664,In_864);
nor U169 (N_169,In_863,In_562);
and U170 (N_170,In_86,In_43);
nor U171 (N_171,In_920,In_139);
nand U172 (N_172,In_765,In_927);
nand U173 (N_173,In_331,In_881);
nand U174 (N_174,In_954,In_839);
xor U175 (N_175,In_795,In_310);
or U176 (N_176,In_587,In_794);
nor U177 (N_177,In_328,In_981);
nor U178 (N_178,In_650,In_54);
or U179 (N_179,In_601,In_732);
and U180 (N_180,In_302,In_516);
or U181 (N_181,In_714,In_84);
nor U182 (N_182,In_783,In_748);
nand U183 (N_183,In_107,In_754);
or U184 (N_184,In_742,In_273);
and U185 (N_185,In_394,In_942);
nand U186 (N_186,In_862,In_250);
or U187 (N_187,In_959,In_547);
nor U188 (N_188,In_152,In_179);
nand U189 (N_189,In_603,In_799);
nand U190 (N_190,In_772,In_483);
and U191 (N_191,In_381,In_18);
nor U192 (N_192,In_681,In_931);
nor U193 (N_193,In_717,In_924);
nor U194 (N_194,In_877,In_701);
or U195 (N_195,In_781,In_885);
nand U196 (N_196,In_338,In_570);
nor U197 (N_197,In_670,In_383);
and U198 (N_198,In_972,In_813);
nand U199 (N_199,In_268,In_121);
nor U200 (N_200,In_61,In_341);
or U201 (N_201,In_269,In_994);
nor U202 (N_202,In_667,In_183);
nand U203 (N_203,In_13,In_362);
nand U204 (N_204,In_499,In_161);
or U205 (N_205,In_975,In_156);
nand U206 (N_206,In_999,In_644);
or U207 (N_207,In_485,In_206);
or U208 (N_208,In_709,In_876);
or U209 (N_209,In_62,In_83);
nand U210 (N_210,In_950,In_529);
nand U211 (N_211,In_263,In_884);
nor U212 (N_212,In_858,In_775);
nand U213 (N_213,In_913,In_860);
nand U214 (N_214,In_467,In_372);
nand U215 (N_215,In_855,In_350);
nand U216 (N_216,In_333,In_354);
nand U217 (N_217,In_169,In_204);
nor U218 (N_218,In_12,In_137);
nand U219 (N_219,In_31,In_825);
nor U220 (N_220,In_340,In_886);
or U221 (N_221,In_42,In_64);
nand U222 (N_222,In_92,In_502);
or U223 (N_223,In_226,In_274);
nor U224 (N_224,In_751,In_361);
nor U225 (N_225,In_607,In_523);
nor U226 (N_226,In_103,In_56);
or U227 (N_227,In_367,In_559);
or U228 (N_228,In_188,In_52);
nand U229 (N_229,In_705,In_157);
or U230 (N_230,In_213,In_317);
or U231 (N_231,In_713,In_823);
and U232 (N_232,In_207,In_512);
or U233 (N_233,In_509,In_113);
or U234 (N_234,In_891,In_583);
nor U235 (N_235,In_150,In_989);
nor U236 (N_236,In_556,In_633);
or U237 (N_237,In_893,In_337);
nand U238 (N_238,In_392,In_867);
and U239 (N_239,In_308,In_976);
and U240 (N_240,In_768,In_782);
and U241 (N_241,In_843,In_143);
and U242 (N_242,In_604,In_335);
nand U243 (N_243,In_197,In_490);
or U244 (N_244,In_926,In_370);
nand U245 (N_245,In_643,In_193);
and U246 (N_246,In_846,In_287);
and U247 (N_247,In_687,In_349);
or U248 (N_248,In_760,In_324);
nand U249 (N_249,In_73,In_766);
nand U250 (N_250,In_600,In_585);
or U251 (N_251,In_388,In_192);
nand U252 (N_252,In_275,In_79);
nor U253 (N_253,In_439,In_141);
or U254 (N_254,In_290,In_816);
nor U255 (N_255,In_117,In_778);
nor U256 (N_256,In_229,In_805);
nor U257 (N_257,In_342,In_115);
or U258 (N_258,In_380,In_5);
nand U259 (N_259,In_131,In_442);
nor U260 (N_260,In_233,In_534);
and U261 (N_261,In_646,In_120);
nor U262 (N_262,In_569,In_946);
nor U263 (N_263,In_395,In_108);
or U264 (N_264,In_627,In_571);
or U265 (N_265,In_195,In_76);
nor U266 (N_266,In_506,In_314);
nand U267 (N_267,In_568,In_983);
or U268 (N_268,In_329,In_616);
nor U269 (N_269,In_545,In_609);
and U270 (N_270,In_634,In_576);
or U271 (N_271,In_683,In_619);
nand U272 (N_272,In_853,In_16);
or U273 (N_273,In_708,In_628);
nand U274 (N_274,In_378,In_582);
and U275 (N_275,In_278,In_749);
and U276 (N_276,In_359,In_284);
and U277 (N_277,In_868,In_809);
nand U278 (N_278,In_67,In_637);
nor U279 (N_279,In_245,In_468);
xor U280 (N_280,In_639,In_567);
nor U281 (N_281,In_396,In_272);
and U282 (N_282,In_723,In_525);
nand U283 (N_283,In_234,In_160);
nor U284 (N_284,In_982,In_326);
xor U285 (N_285,In_831,In_861);
and U286 (N_286,In_671,In_190);
and U287 (N_287,In_185,In_763);
and U288 (N_288,In_598,In_649);
and U289 (N_289,In_382,In_371);
or U290 (N_290,In_666,In_277);
or U291 (N_291,In_677,In_315);
nand U292 (N_292,In_945,In_292);
nor U293 (N_293,In_753,In_856);
nor U294 (N_294,In_847,In_694);
and U295 (N_295,In_764,In_281);
nand U296 (N_296,In_922,In_544);
nor U297 (N_297,In_48,In_352);
and U298 (N_298,In_530,In_198);
and U299 (N_299,In_615,In_124);
nand U300 (N_300,In_729,In_832);
nor U301 (N_301,In_219,In_566);
or U302 (N_302,In_743,In_898);
nand U303 (N_303,In_536,In_631);
or U304 (N_304,In_256,In_948);
xor U305 (N_305,In_804,In_325);
nor U306 (N_306,In_470,In_322);
nand U307 (N_307,In_305,In_526);
and U308 (N_308,In_622,In_613);
nand U309 (N_309,In_144,In_460);
and U310 (N_310,In_953,In_905);
xnor U311 (N_311,In_384,In_704);
or U312 (N_312,In_578,In_815);
and U313 (N_313,In_98,In_327);
or U314 (N_314,In_663,In_851);
and U315 (N_315,In_21,In_970);
or U316 (N_316,In_360,In_938);
nand U317 (N_317,In_919,In_0);
nand U318 (N_318,In_741,In_90);
and U319 (N_319,In_455,In_312);
nor U320 (N_320,In_433,In_116);
and U321 (N_321,In_82,In_210);
and U322 (N_322,In_517,In_110);
or U323 (N_323,In_37,In_168);
nand U324 (N_324,In_923,In_554);
nor U325 (N_325,In_998,In_606);
nand U326 (N_326,In_718,In_311);
nor U327 (N_327,In_934,In_28);
or U328 (N_328,In_454,In_251);
or U329 (N_329,In_126,In_158);
or U330 (N_330,In_824,In_356);
nand U331 (N_331,In_682,In_969);
nand U332 (N_332,In_7,In_323);
and U333 (N_333,In_180,In_127);
and U334 (N_334,In_125,In_3);
nor U335 (N_335,In_964,In_142);
or U336 (N_336,In_403,In_461);
xnor U337 (N_337,In_561,In_45);
nand U338 (N_338,In_865,In_987);
and U339 (N_339,In_402,In_105);
nand U340 (N_340,In_550,In_298);
or U341 (N_341,In_833,In_612);
and U342 (N_342,In_164,In_220);
and U343 (N_343,In_111,In_829);
nand U344 (N_344,In_623,In_689);
nor U345 (N_345,In_289,In_658);
nand U346 (N_346,In_787,In_800);
nand U347 (N_347,In_15,In_266);
nor U348 (N_348,In_334,In_492);
and U349 (N_349,In_140,In_475);
and U350 (N_350,In_917,In_608);
nor U351 (N_351,In_466,In_153);
nand U352 (N_352,In_293,In_620);
nand U353 (N_353,In_882,In_507);
or U354 (N_354,In_456,In_280);
nor U355 (N_355,In_171,In_844);
xor U356 (N_356,In_887,In_553);
nor U357 (N_357,In_756,In_617);
and U358 (N_358,In_769,In_2);
and U359 (N_359,In_834,In_572);
nand U360 (N_360,In_779,In_786);
or U361 (N_361,In_784,In_412);
nor U362 (N_362,In_202,In_104);
nor U363 (N_363,In_738,In_267);
or U364 (N_364,In_424,In_203);
or U365 (N_365,In_733,In_417);
nor U366 (N_366,In_850,In_870);
nand U367 (N_367,In_635,In_912);
and U368 (N_368,In_306,In_679);
nand U369 (N_369,In_827,In_935);
or U370 (N_370,In_465,In_473);
xnor U371 (N_371,In_595,In_869);
xor U372 (N_372,In_358,In_925);
or U373 (N_373,In_50,In_246);
or U374 (N_374,In_159,In_347);
nand U375 (N_375,In_848,In_259);
nand U376 (N_376,In_504,In_533);
and U377 (N_377,In_967,In_430);
nor U378 (N_378,In_484,In_214);
or U379 (N_379,In_264,In_564);
and U380 (N_380,In_151,In_489);
nand U381 (N_381,In_563,In_908);
or U382 (N_382,In_514,In_818);
nand U383 (N_383,In_498,In_737);
or U384 (N_384,In_345,In_242);
and U385 (N_385,In_776,In_177);
nand U386 (N_386,In_774,In_398);
nor U387 (N_387,In_894,In_660);
nor U388 (N_388,In_872,In_46);
nand U389 (N_389,In_665,In_866);
and U390 (N_390,In_68,In_81);
and U391 (N_391,In_988,In_508);
nand U392 (N_392,In_400,In_524);
or U393 (N_393,In_155,In_597);
nor U394 (N_394,In_44,In_299);
nand U395 (N_395,In_170,In_659);
or U396 (N_396,In_916,In_580);
nand U397 (N_397,In_346,In_85);
and U398 (N_398,In_491,In_173);
nor U399 (N_399,In_577,In_72);
or U400 (N_400,In_943,In_914);
and U401 (N_401,In_896,In_87);
nand U402 (N_402,In_415,In_767);
nand U403 (N_403,In_288,In_761);
nor U404 (N_404,In_49,In_900);
nand U405 (N_405,In_930,In_731);
or U406 (N_406,In_820,In_520);
nor U407 (N_407,In_78,In_477);
or U408 (N_408,In_51,In_53);
and U409 (N_409,In_691,In_539);
nor U410 (N_410,In_132,In_38);
and U411 (N_411,In_835,In_236);
nand U412 (N_412,In_471,In_230);
nor U413 (N_413,In_611,In_830);
xnor U414 (N_414,In_986,In_500);
nand U415 (N_415,In_459,In_194);
nand U416 (N_416,In_332,In_590);
nand U417 (N_417,In_574,In_435);
nand U418 (N_418,In_348,In_6);
nor U419 (N_419,In_57,In_369);
nand U420 (N_420,In_377,In_344);
or U421 (N_421,In_426,In_873);
and U422 (N_422,In_494,In_947);
nand U423 (N_423,In_376,In_9);
nand U424 (N_424,In_69,In_313);
nand U425 (N_425,In_955,In_27);
nor U426 (N_426,In_589,In_680);
nand U427 (N_427,In_910,In_425);
or U428 (N_428,In_993,In_669);
and U429 (N_429,In_647,In_80);
or U430 (N_430,In_618,In_450);
or U431 (N_431,In_770,In_283);
or U432 (N_432,In_41,In_857);
or U433 (N_433,In_505,In_451);
nor U434 (N_434,In_295,In_904);
nand U435 (N_435,In_486,In_420);
and U436 (N_436,In_448,In_806);
or U437 (N_437,In_187,In_719);
nor U438 (N_438,In_235,In_252);
nand U439 (N_439,In_593,In_789);
nand U440 (N_440,In_625,In_411);
and U441 (N_441,In_979,In_684);
nor U442 (N_442,In_879,In_70);
or U443 (N_443,In_208,In_249);
xnor U444 (N_444,In_722,In_59);
and U445 (N_445,In_541,In_532);
nand U446 (N_446,In_716,In_991);
or U447 (N_447,In_444,In_181);
nand U448 (N_448,In_596,In_393);
nand U449 (N_449,In_60,In_247);
nor U450 (N_450,In_560,In_706);
nand U451 (N_451,In_29,In_146);
and U452 (N_452,In_413,In_32);
and U453 (N_453,In_89,In_538);
and U454 (N_454,In_688,In_479);
nand U455 (N_455,In_711,In_642);
nand U456 (N_456,In_201,In_209);
nand U457 (N_457,In_686,In_758);
or U458 (N_458,In_883,In_404);
nor U459 (N_459,In_24,In_118);
and U460 (N_460,In_463,In_762);
or U461 (N_461,In_899,In_995);
nand U462 (N_462,In_707,In_122);
nor U463 (N_463,In_493,In_973);
and U464 (N_464,In_211,In_645);
nand U465 (N_465,In_662,In_186);
nor U466 (N_466,In_93,In_401);
nor U467 (N_467,In_431,In_474);
or U468 (N_468,In_414,In_189);
or U469 (N_469,In_715,In_726);
and U470 (N_470,In_528,In_573);
nand U471 (N_471,In_374,In_163);
or U472 (N_472,In_773,In_307);
nor U473 (N_473,In_661,In_757);
and U474 (N_474,In_725,In_225);
and U475 (N_475,In_30,In_178);
nor U476 (N_476,In_739,In_429);
or U477 (N_477,In_481,In_320);
nand U478 (N_478,In_14,In_365);
or U479 (N_479,In_237,In_906);
or U480 (N_480,In_428,In_811);
or U481 (N_481,In_630,In_88);
nand U482 (N_482,In_136,In_407);
nand U483 (N_483,In_821,In_452);
nand U484 (N_484,In_803,In_36);
nand U485 (N_485,In_167,In_958);
and U486 (N_486,In_309,In_932);
and U487 (N_487,In_978,In_963);
and U488 (N_488,In_301,In_962);
nor U489 (N_489,In_817,In_114);
or U490 (N_490,In_339,In_241);
nand U491 (N_491,In_94,In_849);
nor U492 (N_492,In_777,In_785);
or U493 (N_493,In_515,In_697);
nand U494 (N_494,In_788,In_918);
nor U495 (N_495,In_730,In_419);
or U496 (N_496,In_445,In_238);
nand U497 (N_497,In_223,In_921);
nor U498 (N_498,In_300,In_478);
and U499 (N_499,In_218,In_845);
or U500 (N_500,N_165,N_239);
or U501 (N_501,N_243,N_58);
and U502 (N_502,N_322,N_261);
and U503 (N_503,N_182,N_190);
or U504 (N_504,N_480,N_153);
or U505 (N_505,N_24,N_309);
and U506 (N_506,N_85,N_276);
or U507 (N_507,N_47,N_352);
or U508 (N_508,N_180,N_465);
nand U509 (N_509,N_428,N_469);
or U510 (N_510,N_226,N_50);
or U511 (N_511,N_392,N_35);
nand U512 (N_512,N_211,N_23);
or U513 (N_513,N_415,N_136);
or U514 (N_514,N_474,N_235);
or U515 (N_515,N_269,N_342);
or U516 (N_516,N_257,N_44);
nor U517 (N_517,N_156,N_344);
nand U518 (N_518,N_464,N_424);
and U519 (N_519,N_193,N_305);
nand U520 (N_520,N_214,N_338);
or U521 (N_521,N_216,N_200);
and U522 (N_522,N_423,N_408);
and U523 (N_523,N_53,N_476);
or U524 (N_524,N_181,N_233);
and U525 (N_525,N_75,N_5);
nand U526 (N_526,N_270,N_337);
nand U527 (N_527,N_238,N_323);
nor U528 (N_528,N_391,N_160);
and U529 (N_529,N_348,N_314);
and U530 (N_530,N_185,N_63);
nand U531 (N_531,N_9,N_46);
and U532 (N_532,N_37,N_183);
nor U533 (N_533,N_264,N_496);
and U534 (N_534,N_402,N_378);
nand U535 (N_535,N_293,N_256);
or U536 (N_536,N_297,N_110);
and U537 (N_537,N_225,N_365);
or U538 (N_538,N_72,N_25);
nor U539 (N_539,N_466,N_401);
nand U540 (N_540,N_353,N_371);
or U541 (N_541,N_55,N_260);
or U542 (N_542,N_277,N_92);
nor U543 (N_543,N_358,N_141);
or U544 (N_544,N_333,N_86);
or U545 (N_545,N_355,N_307);
nor U546 (N_546,N_306,N_409);
nor U547 (N_547,N_76,N_390);
or U548 (N_548,N_395,N_335);
nand U549 (N_549,N_191,N_71);
nand U550 (N_550,N_117,N_280);
or U551 (N_551,N_123,N_278);
nand U552 (N_552,N_387,N_368);
nor U553 (N_553,N_328,N_351);
nand U554 (N_554,N_412,N_294);
or U555 (N_555,N_356,N_431);
or U556 (N_556,N_445,N_189);
nor U557 (N_557,N_32,N_155);
nand U558 (N_558,N_282,N_427);
or U559 (N_559,N_285,N_393);
nor U560 (N_560,N_206,N_299);
nor U561 (N_561,N_486,N_96);
or U562 (N_562,N_478,N_223);
and U563 (N_563,N_467,N_375);
nand U564 (N_564,N_18,N_34);
and U565 (N_565,N_12,N_458);
nand U566 (N_566,N_376,N_176);
and U567 (N_567,N_97,N_129);
nand U568 (N_568,N_184,N_361);
nand U569 (N_569,N_384,N_219);
xor U570 (N_570,N_255,N_324);
or U571 (N_571,N_103,N_405);
xnor U572 (N_572,N_51,N_265);
and U573 (N_573,N_281,N_48);
nand U574 (N_574,N_186,N_274);
nand U575 (N_575,N_263,N_144);
nor U576 (N_576,N_109,N_432);
nor U577 (N_577,N_454,N_380);
and U578 (N_578,N_388,N_490);
and U579 (N_579,N_435,N_119);
or U580 (N_580,N_493,N_317);
nand U581 (N_581,N_227,N_242);
or U582 (N_582,N_475,N_69);
nor U583 (N_583,N_203,N_481);
nand U584 (N_584,N_217,N_291);
and U585 (N_585,N_229,N_349);
nand U586 (N_586,N_171,N_89);
nor U587 (N_587,N_316,N_441);
xor U588 (N_588,N_52,N_379);
and U589 (N_589,N_443,N_252);
nand U590 (N_590,N_42,N_78);
nor U591 (N_591,N_472,N_138);
nand U592 (N_592,N_275,N_347);
nor U593 (N_593,N_396,N_421);
and U594 (N_594,N_450,N_383);
nor U595 (N_595,N_341,N_66);
or U596 (N_596,N_462,N_150);
and U597 (N_597,N_404,N_3);
nor U598 (N_598,N_363,N_204);
and U599 (N_599,N_177,N_403);
or U600 (N_600,N_115,N_374);
nor U601 (N_601,N_170,N_372);
or U602 (N_602,N_112,N_7);
or U603 (N_603,N_362,N_438);
or U604 (N_604,N_461,N_369);
nand U605 (N_605,N_471,N_311);
nor U606 (N_606,N_77,N_482);
nor U607 (N_607,N_198,N_143);
nor U608 (N_608,N_116,N_433);
or U609 (N_609,N_308,N_83);
nand U610 (N_610,N_303,N_498);
or U611 (N_611,N_179,N_407);
or U612 (N_612,N_253,N_329);
nand U613 (N_613,N_240,N_146);
and U614 (N_614,N_87,N_137);
nor U615 (N_615,N_298,N_377);
and U616 (N_616,N_343,N_487);
and U617 (N_617,N_367,N_221);
nor U618 (N_618,N_447,N_95);
and U619 (N_619,N_149,N_159);
nand U620 (N_620,N_381,N_151);
or U621 (N_621,N_147,N_82);
and U622 (N_622,N_398,N_222);
and U623 (N_623,N_187,N_249);
and U624 (N_624,N_301,N_33);
nor U625 (N_625,N_406,N_36);
or U626 (N_626,N_489,N_312);
xor U627 (N_627,N_266,N_73);
nor U628 (N_628,N_325,N_286);
or U629 (N_629,N_131,N_429);
xnor U630 (N_630,N_65,N_479);
or U631 (N_631,N_102,N_114);
nand U632 (N_632,N_470,N_172);
nor U633 (N_633,N_457,N_205);
nand U634 (N_634,N_339,N_14);
nor U635 (N_635,N_289,N_440);
and U636 (N_636,N_332,N_57);
or U637 (N_637,N_357,N_473);
nand U638 (N_638,N_28,N_494);
nand U639 (N_639,N_157,N_350);
nand U640 (N_640,N_212,N_60);
or U641 (N_641,N_439,N_340);
or U642 (N_642,N_290,N_459);
nand U643 (N_643,N_122,N_346);
or U644 (N_644,N_237,N_236);
and U645 (N_645,N_99,N_100);
nor U646 (N_646,N_118,N_126);
or U647 (N_647,N_16,N_254);
nor U648 (N_648,N_202,N_444);
nor U649 (N_649,N_484,N_313);
nand U650 (N_650,N_84,N_272);
xnor U651 (N_651,N_326,N_174);
nor U652 (N_652,N_283,N_245);
nor U653 (N_653,N_111,N_492);
or U654 (N_654,N_38,N_468);
or U655 (N_655,N_130,N_104);
and U656 (N_656,N_22,N_244);
nand U657 (N_657,N_15,N_19);
and U658 (N_658,N_246,N_108);
nand U659 (N_659,N_8,N_319);
nor U660 (N_660,N_224,N_2);
nor U661 (N_661,N_135,N_68);
nand U662 (N_662,N_477,N_91);
or U663 (N_663,N_70,N_56);
nor U664 (N_664,N_162,N_426);
and U665 (N_665,N_161,N_196);
and U666 (N_666,N_210,N_142);
and U667 (N_667,N_310,N_41);
or U668 (N_668,N_295,N_419);
nor U669 (N_669,N_241,N_359);
nor U670 (N_670,N_296,N_140);
or U671 (N_671,N_437,N_448);
nor U672 (N_672,N_321,N_148);
nand U673 (N_673,N_373,N_336);
or U674 (N_674,N_158,N_121);
or U675 (N_675,N_154,N_394);
nand U676 (N_676,N_389,N_132);
nand U677 (N_677,N_267,N_43);
and U678 (N_678,N_54,N_300);
nand U679 (N_679,N_345,N_13);
and U680 (N_680,N_334,N_133);
nor U681 (N_681,N_201,N_152);
nor U682 (N_682,N_456,N_287);
and U683 (N_683,N_168,N_215);
nor U684 (N_684,N_59,N_483);
or U685 (N_685,N_209,N_268);
xnor U686 (N_686,N_213,N_79);
xor U687 (N_687,N_400,N_385);
and U688 (N_688,N_232,N_134);
xor U689 (N_689,N_248,N_6);
or U690 (N_690,N_61,N_167);
or U691 (N_691,N_105,N_418);
nand U692 (N_692,N_382,N_29);
or U693 (N_693,N_208,N_113);
nor U694 (N_694,N_485,N_262);
or U695 (N_695,N_88,N_45);
nand U696 (N_696,N_26,N_331);
and U697 (N_697,N_31,N_320);
xnor U698 (N_698,N_315,N_218);
and U699 (N_699,N_64,N_284);
nor U700 (N_700,N_247,N_499);
and U701 (N_701,N_279,N_425);
or U702 (N_702,N_327,N_175);
nand U703 (N_703,N_0,N_98);
and U704 (N_704,N_139,N_292);
nor U705 (N_705,N_107,N_164);
and U706 (N_706,N_106,N_30);
or U707 (N_707,N_192,N_94);
or U708 (N_708,N_250,N_452);
nand U709 (N_709,N_360,N_39);
or U710 (N_710,N_497,N_195);
nand U711 (N_711,N_386,N_81);
and U712 (N_712,N_145,N_453);
and U713 (N_713,N_304,N_1);
nand U714 (N_714,N_10,N_128);
nand U715 (N_715,N_318,N_67);
nor U716 (N_716,N_194,N_488);
or U717 (N_717,N_163,N_220);
nor U718 (N_718,N_410,N_93);
xor U719 (N_719,N_491,N_302);
or U720 (N_720,N_188,N_27);
nor U721 (N_721,N_463,N_178);
or U722 (N_722,N_234,N_197);
nand U723 (N_723,N_330,N_228);
and U724 (N_724,N_173,N_166);
nor U725 (N_725,N_288,N_399);
and U726 (N_726,N_259,N_416);
nand U727 (N_727,N_460,N_370);
and U728 (N_728,N_62,N_420);
and U729 (N_729,N_446,N_169);
or U730 (N_730,N_124,N_11);
nor U731 (N_731,N_417,N_434);
and U732 (N_732,N_49,N_413);
or U733 (N_733,N_127,N_271);
and U734 (N_734,N_74,N_397);
nor U735 (N_735,N_251,N_125);
and U736 (N_736,N_90,N_354);
or U737 (N_737,N_414,N_273);
or U738 (N_738,N_20,N_258);
nor U739 (N_739,N_411,N_21);
nor U740 (N_740,N_40,N_4);
nor U741 (N_741,N_451,N_231);
or U742 (N_742,N_436,N_442);
and U743 (N_743,N_364,N_17);
and U744 (N_744,N_120,N_101);
and U745 (N_745,N_207,N_422);
nand U746 (N_746,N_449,N_455);
or U747 (N_747,N_495,N_366);
and U748 (N_748,N_80,N_230);
or U749 (N_749,N_430,N_199);
or U750 (N_750,N_338,N_18);
nand U751 (N_751,N_413,N_101);
nor U752 (N_752,N_440,N_203);
nor U753 (N_753,N_3,N_121);
nand U754 (N_754,N_302,N_317);
or U755 (N_755,N_215,N_276);
nor U756 (N_756,N_436,N_165);
and U757 (N_757,N_495,N_310);
nand U758 (N_758,N_389,N_216);
nand U759 (N_759,N_6,N_132);
nand U760 (N_760,N_82,N_35);
or U761 (N_761,N_238,N_147);
nor U762 (N_762,N_40,N_55);
and U763 (N_763,N_191,N_400);
nand U764 (N_764,N_415,N_445);
nor U765 (N_765,N_286,N_368);
nor U766 (N_766,N_218,N_328);
nand U767 (N_767,N_269,N_326);
nor U768 (N_768,N_85,N_359);
or U769 (N_769,N_85,N_467);
nand U770 (N_770,N_438,N_149);
nor U771 (N_771,N_397,N_38);
nand U772 (N_772,N_247,N_345);
nor U773 (N_773,N_128,N_92);
and U774 (N_774,N_425,N_155);
nand U775 (N_775,N_19,N_343);
or U776 (N_776,N_311,N_249);
and U777 (N_777,N_36,N_115);
nand U778 (N_778,N_368,N_487);
or U779 (N_779,N_196,N_216);
nor U780 (N_780,N_59,N_185);
and U781 (N_781,N_56,N_403);
nand U782 (N_782,N_126,N_300);
nor U783 (N_783,N_131,N_191);
nor U784 (N_784,N_41,N_394);
nor U785 (N_785,N_88,N_110);
nor U786 (N_786,N_43,N_108);
or U787 (N_787,N_320,N_303);
and U788 (N_788,N_118,N_363);
nor U789 (N_789,N_430,N_170);
and U790 (N_790,N_100,N_268);
and U791 (N_791,N_36,N_490);
nor U792 (N_792,N_389,N_283);
and U793 (N_793,N_62,N_224);
nor U794 (N_794,N_8,N_292);
and U795 (N_795,N_52,N_491);
or U796 (N_796,N_348,N_126);
or U797 (N_797,N_88,N_47);
nor U798 (N_798,N_70,N_145);
or U799 (N_799,N_31,N_147);
nor U800 (N_800,N_265,N_60);
nor U801 (N_801,N_282,N_252);
nand U802 (N_802,N_359,N_463);
nand U803 (N_803,N_280,N_484);
nor U804 (N_804,N_291,N_230);
nor U805 (N_805,N_59,N_369);
nand U806 (N_806,N_323,N_268);
and U807 (N_807,N_453,N_43);
and U808 (N_808,N_203,N_114);
and U809 (N_809,N_204,N_112);
and U810 (N_810,N_268,N_228);
nor U811 (N_811,N_386,N_9);
nand U812 (N_812,N_103,N_302);
or U813 (N_813,N_204,N_462);
nor U814 (N_814,N_485,N_7);
or U815 (N_815,N_71,N_371);
xor U816 (N_816,N_298,N_356);
nor U817 (N_817,N_298,N_133);
nand U818 (N_818,N_293,N_483);
and U819 (N_819,N_234,N_312);
nor U820 (N_820,N_317,N_385);
nor U821 (N_821,N_42,N_44);
nand U822 (N_822,N_225,N_413);
nor U823 (N_823,N_418,N_368);
nand U824 (N_824,N_328,N_185);
and U825 (N_825,N_29,N_181);
and U826 (N_826,N_476,N_194);
and U827 (N_827,N_210,N_432);
nor U828 (N_828,N_93,N_417);
and U829 (N_829,N_480,N_99);
or U830 (N_830,N_18,N_242);
nor U831 (N_831,N_233,N_441);
nand U832 (N_832,N_492,N_312);
or U833 (N_833,N_152,N_437);
nand U834 (N_834,N_276,N_45);
nand U835 (N_835,N_374,N_207);
nand U836 (N_836,N_427,N_144);
nand U837 (N_837,N_436,N_494);
nand U838 (N_838,N_441,N_412);
nor U839 (N_839,N_84,N_424);
nor U840 (N_840,N_415,N_306);
nand U841 (N_841,N_106,N_77);
nor U842 (N_842,N_118,N_71);
nand U843 (N_843,N_76,N_384);
and U844 (N_844,N_167,N_297);
and U845 (N_845,N_366,N_360);
and U846 (N_846,N_460,N_487);
nand U847 (N_847,N_320,N_146);
or U848 (N_848,N_292,N_48);
and U849 (N_849,N_12,N_17);
nand U850 (N_850,N_382,N_345);
or U851 (N_851,N_450,N_361);
nand U852 (N_852,N_234,N_434);
or U853 (N_853,N_441,N_280);
and U854 (N_854,N_289,N_207);
nor U855 (N_855,N_420,N_418);
and U856 (N_856,N_88,N_434);
and U857 (N_857,N_287,N_83);
and U858 (N_858,N_290,N_45);
or U859 (N_859,N_240,N_14);
xor U860 (N_860,N_297,N_248);
and U861 (N_861,N_402,N_450);
and U862 (N_862,N_372,N_305);
and U863 (N_863,N_408,N_313);
nand U864 (N_864,N_465,N_454);
nor U865 (N_865,N_190,N_98);
nand U866 (N_866,N_100,N_199);
nand U867 (N_867,N_257,N_400);
or U868 (N_868,N_104,N_487);
nor U869 (N_869,N_498,N_355);
nand U870 (N_870,N_247,N_64);
nand U871 (N_871,N_97,N_6);
nor U872 (N_872,N_153,N_138);
nand U873 (N_873,N_326,N_316);
nor U874 (N_874,N_220,N_93);
nor U875 (N_875,N_43,N_352);
nand U876 (N_876,N_28,N_238);
nand U877 (N_877,N_346,N_169);
or U878 (N_878,N_61,N_143);
nor U879 (N_879,N_59,N_265);
and U880 (N_880,N_253,N_494);
nor U881 (N_881,N_261,N_367);
nand U882 (N_882,N_5,N_372);
nand U883 (N_883,N_182,N_98);
nand U884 (N_884,N_416,N_218);
nor U885 (N_885,N_330,N_434);
xor U886 (N_886,N_204,N_263);
nor U887 (N_887,N_263,N_78);
nand U888 (N_888,N_79,N_153);
nand U889 (N_889,N_442,N_489);
nand U890 (N_890,N_22,N_407);
nand U891 (N_891,N_40,N_396);
nand U892 (N_892,N_452,N_65);
nor U893 (N_893,N_350,N_431);
and U894 (N_894,N_163,N_322);
nand U895 (N_895,N_191,N_62);
and U896 (N_896,N_123,N_36);
nor U897 (N_897,N_190,N_188);
nor U898 (N_898,N_277,N_409);
nor U899 (N_899,N_236,N_284);
xnor U900 (N_900,N_189,N_145);
and U901 (N_901,N_248,N_54);
nand U902 (N_902,N_104,N_287);
and U903 (N_903,N_344,N_244);
or U904 (N_904,N_66,N_166);
nor U905 (N_905,N_271,N_175);
or U906 (N_906,N_81,N_268);
and U907 (N_907,N_146,N_311);
nand U908 (N_908,N_92,N_112);
nand U909 (N_909,N_416,N_294);
nor U910 (N_910,N_333,N_222);
nand U911 (N_911,N_479,N_48);
and U912 (N_912,N_425,N_58);
or U913 (N_913,N_335,N_94);
nor U914 (N_914,N_213,N_332);
and U915 (N_915,N_322,N_304);
nand U916 (N_916,N_145,N_264);
or U917 (N_917,N_146,N_173);
and U918 (N_918,N_49,N_443);
or U919 (N_919,N_7,N_461);
nor U920 (N_920,N_16,N_126);
nor U921 (N_921,N_322,N_369);
nor U922 (N_922,N_120,N_65);
and U923 (N_923,N_40,N_349);
nor U924 (N_924,N_200,N_6);
and U925 (N_925,N_498,N_468);
nand U926 (N_926,N_92,N_119);
or U927 (N_927,N_175,N_82);
nand U928 (N_928,N_44,N_319);
xnor U929 (N_929,N_51,N_361);
nor U930 (N_930,N_206,N_4);
nor U931 (N_931,N_88,N_195);
and U932 (N_932,N_88,N_438);
or U933 (N_933,N_167,N_396);
or U934 (N_934,N_77,N_46);
and U935 (N_935,N_402,N_61);
nor U936 (N_936,N_269,N_31);
nand U937 (N_937,N_222,N_484);
nor U938 (N_938,N_237,N_369);
and U939 (N_939,N_122,N_404);
nor U940 (N_940,N_434,N_400);
and U941 (N_941,N_232,N_141);
nand U942 (N_942,N_53,N_277);
and U943 (N_943,N_119,N_359);
xor U944 (N_944,N_431,N_374);
nor U945 (N_945,N_301,N_164);
or U946 (N_946,N_432,N_289);
or U947 (N_947,N_94,N_313);
nor U948 (N_948,N_442,N_481);
and U949 (N_949,N_377,N_212);
nand U950 (N_950,N_425,N_169);
nand U951 (N_951,N_311,N_342);
or U952 (N_952,N_123,N_128);
nor U953 (N_953,N_370,N_451);
nand U954 (N_954,N_8,N_96);
and U955 (N_955,N_195,N_241);
or U956 (N_956,N_415,N_260);
and U957 (N_957,N_419,N_385);
and U958 (N_958,N_423,N_16);
or U959 (N_959,N_488,N_60);
or U960 (N_960,N_409,N_82);
and U961 (N_961,N_311,N_15);
nor U962 (N_962,N_221,N_128);
nand U963 (N_963,N_484,N_494);
nand U964 (N_964,N_125,N_359);
and U965 (N_965,N_360,N_200);
or U966 (N_966,N_144,N_138);
or U967 (N_967,N_159,N_206);
or U968 (N_968,N_377,N_333);
and U969 (N_969,N_173,N_259);
or U970 (N_970,N_326,N_21);
or U971 (N_971,N_290,N_207);
nand U972 (N_972,N_375,N_196);
or U973 (N_973,N_356,N_204);
nand U974 (N_974,N_404,N_198);
nand U975 (N_975,N_227,N_347);
or U976 (N_976,N_162,N_7);
or U977 (N_977,N_449,N_119);
nor U978 (N_978,N_438,N_296);
nand U979 (N_979,N_293,N_415);
or U980 (N_980,N_423,N_174);
and U981 (N_981,N_96,N_134);
nor U982 (N_982,N_198,N_334);
or U983 (N_983,N_311,N_250);
and U984 (N_984,N_249,N_72);
or U985 (N_985,N_216,N_112);
and U986 (N_986,N_410,N_59);
xnor U987 (N_987,N_313,N_196);
and U988 (N_988,N_233,N_409);
nand U989 (N_989,N_116,N_68);
and U990 (N_990,N_244,N_472);
or U991 (N_991,N_223,N_277);
nor U992 (N_992,N_123,N_438);
nor U993 (N_993,N_69,N_329);
or U994 (N_994,N_366,N_351);
nand U995 (N_995,N_108,N_70);
or U996 (N_996,N_296,N_485);
and U997 (N_997,N_339,N_350);
and U998 (N_998,N_117,N_148);
and U999 (N_999,N_359,N_377);
and U1000 (N_1000,N_866,N_731);
nand U1001 (N_1001,N_674,N_571);
or U1002 (N_1002,N_645,N_560);
or U1003 (N_1003,N_549,N_532);
nor U1004 (N_1004,N_935,N_543);
and U1005 (N_1005,N_874,N_569);
and U1006 (N_1006,N_746,N_816);
nand U1007 (N_1007,N_715,N_921);
or U1008 (N_1008,N_535,N_949);
or U1009 (N_1009,N_834,N_891);
nand U1010 (N_1010,N_855,N_859);
nand U1011 (N_1011,N_554,N_660);
nand U1012 (N_1012,N_649,N_975);
and U1013 (N_1013,N_599,N_735);
and U1014 (N_1014,N_681,N_594);
or U1015 (N_1015,N_888,N_576);
nor U1016 (N_1016,N_792,N_787);
and U1017 (N_1017,N_690,N_580);
nor U1018 (N_1018,N_887,N_820);
nor U1019 (N_1019,N_676,N_992);
nor U1020 (N_1020,N_971,N_752);
or U1021 (N_1021,N_770,N_922);
and U1022 (N_1022,N_913,N_893);
nor U1023 (N_1023,N_826,N_555);
and U1024 (N_1024,N_798,N_501);
nand U1025 (N_1025,N_698,N_617);
and U1026 (N_1026,N_979,N_999);
nand U1027 (N_1027,N_601,N_616);
nand U1028 (N_1028,N_765,N_609);
nand U1029 (N_1029,N_635,N_791);
or U1030 (N_1030,N_602,N_663);
nand U1031 (N_1031,N_824,N_961);
nor U1032 (N_1032,N_693,N_627);
and U1033 (N_1033,N_854,N_926);
nor U1034 (N_1034,N_694,N_908);
or U1035 (N_1035,N_699,N_907);
or U1036 (N_1036,N_520,N_568);
nand U1037 (N_1037,N_729,N_689);
or U1038 (N_1038,N_559,N_800);
xnor U1039 (N_1039,N_864,N_719);
nand U1040 (N_1040,N_574,N_714);
nor U1041 (N_1041,N_626,N_769);
nor U1042 (N_1042,N_942,N_563);
and U1043 (N_1043,N_784,N_598);
or U1044 (N_1044,N_890,N_675);
xnor U1045 (N_1045,N_723,N_783);
nand U1046 (N_1046,N_621,N_788);
and U1047 (N_1047,N_822,N_958);
or U1048 (N_1048,N_604,N_722);
or U1049 (N_1049,N_768,N_688);
nand U1050 (N_1050,N_696,N_998);
and U1051 (N_1051,N_780,N_751);
and U1052 (N_1052,N_940,N_686);
nor U1053 (N_1053,N_644,N_778);
nor U1054 (N_1054,N_502,N_705);
or U1055 (N_1055,N_795,N_753);
nor U1056 (N_1056,N_589,N_670);
nor U1057 (N_1057,N_880,N_703);
nand U1058 (N_1058,N_619,N_678);
and U1059 (N_1059,N_558,N_623);
nand U1060 (N_1060,N_588,N_881);
xnor U1061 (N_1061,N_804,N_643);
nand U1062 (N_1062,N_779,N_664);
nor U1063 (N_1063,N_527,N_572);
or U1064 (N_1064,N_716,N_831);
nand U1065 (N_1065,N_565,N_658);
and U1066 (N_1066,N_758,N_882);
nand U1067 (N_1067,N_823,N_615);
and U1068 (N_1068,N_692,N_657);
or U1069 (N_1069,N_785,N_513);
and U1070 (N_1070,N_550,N_841);
and U1071 (N_1071,N_772,N_595);
nor U1072 (N_1072,N_761,N_628);
and U1073 (N_1073,N_759,N_988);
or U1074 (N_1074,N_835,N_906);
nor U1075 (N_1075,N_957,N_512);
nor U1076 (N_1076,N_947,N_633);
nor U1077 (N_1077,N_687,N_585);
nand U1078 (N_1078,N_685,N_732);
or U1079 (N_1079,N_600,N_624);
and U1080 (N_1080,N_548,N_805);
nor U1081 (N_1081,N_630,N_954);
nor U1082 (N_1082,N_587,N_684);
nand U1083 (N_1083,N_724,N_525);
or U1084 (N_1084,N_782,N_544);
or U1085 (N_1085,N_611,N_781);
and U1086 (N_1086,N_567,N_905);
or U1087 (N_1087,N_755,N_523);
nand U1088 (N_1088,N_683,N_648);
or U1089 (N_1089,N_959,N_740);
and U1090 (N_1090,N_937,N_836);
and U1091 (N_1091,N_797,N_597);
or U1092 (N_1092,N_857,N_931);
or U1093 (N_1093,N_516,N_825);
nand U1094 (N_1094,N_744,N_873);
nand U1095 (N_1095,N_970,N_612);
and U1096 (N_1096,N_876,N_878);
nand U1097 (N_1097,N_528,N_861);
nand U1098 (N_1098,N_605,N_529);
and U1099 (N_1099,N_654,N_741);
nand U1100 (N_1100,N_712,N_511);
and U1101 (N_1101,N_659,N_933);
nor U1102 (N_1102,N_691,N_706);
nor U1103 (N_1103,N_538,N_897);
xnor U1104 (N_1104,N_849,N_673);
nor U1105 (N_1105,N_725,N_522);
nor U1106 (N_1106,N_738,N_540);
nor U1107 (N_1107,N_514,N_636);
nand U1108 (N_1108,N_943,N_914);
nor U1109 (N_1109,N_794,N_989);
nand U1110 (N_1110,N_556,N_868);
nand U1111 (N_1111,N_981,N_570);
nand U1112 (N_1112,N_754,N_742);
or U1113 (N_1113,N_777,N_813);
nor U1114 (N_1114,N_899,N_695);
or U1115 (N_1115,N_966,N_726);
nor U1116 (N_1116,N_721,N_996);
and U1117 (N_1117,N_542,N_507);
xor U1118 (N_1118,N_923,N_817);
nand U1119 (N_1119,N_832,N_713);
or U1120 (N_1120,N_924,N_620);
or U1121 (N_1121,N_750,N_521);
and U1122 (N_1122,N_736,N_904);
or U1123 (N_1123,N_504,N_919);
or U1124 (N_1124,N_969,N_747);
nor U1125 (N_1125,N_889,N_566);
and U1126 (N_1126,N_745,N_980);
nor U1127 (N_1127,N_925,N_991);
and U1128 (N_1128,N_707,N_710);
nand U1129 (N_1129,N_728,N_978);
or U1130 (N_1130,N_531,N_642);
or U1131 (N_1131,N_877,N_557);
or U1132 (N_1132,N_774,N_596);
nand U1133 (N_1133,N_972,N_709);
nor U1134 (N_1134,N_995,N_739);
nor U1135 (N_1135,N_500,N_900);
nor U1136 (N_1136,N_869,N_842);
nor U1137 (N_1137,N_871,N_551);
or U1138 (N_1138,N_679,N_677);
nor U1139 (N_1139,N_639,N_509);
nor U1140 (N_1140,N_879,N_593);
or U1141 (N_1141,N_718,N_662);
or U1142 (N_1142,N_524,N_872);
or U1143 (N_1143,N_833,N_505);
nor U1144 (N_1144,N_902,N_766);
or U1145 (N_1145,N_666,N_917);
nand U1146 (N_1146,N_837,N_641);
nor U1147 (N_1147,N_968,N_927);
and U1148 (N_1148,N_590,N_536);
nand U1149 (N_1149,N_821,N_618);
or U1150 (N_1150,N_843,N_840);
and U1151 (N_1151,N_591,N_844);
and U1152 (N_1152,N_862,N_976);
or U1153 (N_1153,N_898,N_748);
or U1154 (N_1154,N_870,N_682);
nor U1155 (N_1155,N_965,N_967);
and U1156 (N_1156,N_672,N_892);
and U1157 (N_1157,N_720,N_903);
nand U1158 (N_1158,N_951,N_809);
nor U1159 (N_1159,N_727,N_583);
nor U1160 (N_1160,N_952,N_910);
or U1161 (N_1161,N_646,N_582);
or U1162 (N_1162,N_749,N_883);
or U1163 (N_1163,N_786,N_652);
or U1164 (N_1164,N_547,N_743);
nand U1165 (N_1165,N_956,N_962);
and U1166 (N_1166,N_929,N_515);
or U1167 (N_1167,N_993,N_847);
nand U1168 (N_1168,N_896,N_796);
nor U1169 (N_1169,N_577,N_901);
and U1170 (N_1170,N_858,N_944);
and U1171 (N_1171,N_909,N_702);
or U1172 (N_1172,N_828,N_885);
nor U1173 (N_1173,N_517,N_762);
nor U1174 (N_1174,N_819,N_603);
nand U1175 (N_1175,N_848,N_632);
and U1176 (N_1176,N_669,N_985);
and U1177 (N_1177,N_799,N_553);
and U1178 (N_1178,N_997,N_561);
and U1179 (N_1179,N_983,N_650);
nand U1180 (N_1180,N_814,N_506);
xnor U1181 (N_1181,N_533,N_773);
nand U1182 (N_1182,N_928,N_578);
or U1183 (N_1183,N_775,N_960);
nor U1184 (N_1184,N_860,N_584);
nand U1185 (N_1185,N_579,N_990);
nor U1186 (N_1186,N_552,N_622);
or U1187 (N_1187,N_934,N_936);
nand U1188 (N_1188,N_946,N_808);
nor U1189 (N_1189,N_802,N_793);
nor U1190 (N_1190,N_733,N_939);
and U1191 (N_1191,N_845,N_730);
nor U1192 (N_1192,N_661,N_867);
nand U1193 (N_1193,N_994,N_656);
and U1194 (N_1194,N_575,N_987);
or U1195 (N_1195,N_941,N_704);
or U1196 (N_1196,N_625,N_853);
and U1197 (N_1197,N_518,N_838);
nand U1198 (N_1198,N_912,N_963);
nor U1199 (N_1199,N_886,N_767);
nor U1200 (N_1200,N_564,N_829);
nand U1201 (N_1201,N_607,N_915);
nor U1202 (N_1202,N_810,N_610);
or U1203 (N_1203,N_634,N_916);
nor U1204 (N_1204,N_647,N_667);
or U1205 (N_1205,N_760,N_606);
and U1206 (N_1206,N_790,N_545);
nand U1207 (N_1207,N_974,N_865);
or U1208 (N_1208,N_653,N_763);
and U1209 (N_1209,N_608,N_982);
or U1210 (N_1210,N_519,N_614);
nor U1211 (N_1211,N_592,N_894);
nand U1212 (N_1212,N_640,N_711);
nor U1213 (N_1213,N_953,N_530);
nand U1214 (N_1214,N_701,N_984);
nand U1215 (N_1215,N_700,N_771);
nand U1216 (N_1216,N_911,N_734);
nor U1217 (N_1217,N_977,N_586);
nor U1218 (N_1218,N_671,N_708);
nand U1219 (N_1219,N_930,N_546);
or U1220 (N_1220,N_812,N_537);
and U1221 (N_1221,N_955,N_613);
nor U1222 (N_1222,N_801,N_803);
nand U1223 (N_1223,N_932,N_717);
or U1224 (N_1224,N_851,N_839);
and U1225 (N_1225,N_806,N_697);
or U1226 (N_1226,N_850,N_918);
xor U1227 (N_1227,N_581,N_651);
and U1228 (N_1228,N_852,N_503);
nor U1229 (N_1229,N_973,N_562);
or U1230 (N_1230,N_920,N_508);
or U1231 (N_1231,N_573,N_526);
and U1232 (N_1232,N_541,N_510);
nand U1233 (N_1233,N_948,N_789);
and U1234 (N_1234,N_986,N_830);
or U1235 (N_1235,N_638,N_818);
nand U1236 (N_1236,N_539,N_856);
and U1237 (N_1237,N_875,N_665);
and U1238 (N_1238,N_764,N_631);
and U1239 (N_1239,N_950,N_668);
and U1240 (N_1240,N_807,N_964);
nand U1241 (N_1241,N_895,N_938);
nand U1242 (N_1242,N_846,N_680);
nor U1243 (N_1243,N_945,N_655);
nor U1244 (N_1244,N_629,N_815);
and U1245 (N_1245,N_811,N_637);
nand U1246 (N_1246,N_756,N_827);
and U1247 (N_1247,N_757,N_534);
xnor U1248 (N_1248,N_884,N_863);
nor U1249 (N_1249,N_737,N_776);
nor U1250 (N_1250,N_801,N_832);
nor U1251 (N_1251,N_838,N_644);
or U1252 (N_1252,N_571,N_577);
nand U1253 (N_1253,N_562,N_561);
or U1254 (N_1254,N_763,N_839);
nand U1255 (N_1255,N_778,N_693);
and U1256 (N_1256,N_692,N_809);
nor U1257 (N_1257,N_800,N_511);
or U1258 (N_1258,N_524,N_730);
or U1259 (N_1259,N_783,N_815);
or U1260 (N_1260,N_642,N_590);
and U1261 (N_1261,N_660,N_875);
or U1262 (N_1262,N_827,N_724);
nor U1263 (N_1263,N_721,N_709);
and U1264 (N_1264,N_842,N_887);
nand U1265 (N_1265,N_583,N_982);
nand U1266 (N_1266,N_504,N_848);
or U1267 (N_1267,N_864,N_736);
and U1268 (N_1268,N_714,N_813);
nand U1269 (N_1269,N_530,N_655);
or U1270 (N_1270,N_686,N_510);
and U1271 (N_1271,N_724,N_850);
xnor U1272 (N_1272,N_976,N_843);
nand U1273 (N_1273,N_691,N_821);
nor U1274 (N_1274,N_925,N_689);
or U1275 (N_1275,N_576,N_610);
nand U1276 (N_1276,N_747,N_765);
nor U1277 (N_1277,N_728,N_560);
nor U1278 (N_1278,N_699,N_928);
nand U1279 (N_1279,N_852,N_689);
nand U1280 (N_1280,N_597,N_603);
nor U1281 (N_1281,N_784,N_962);
or U1282 (N_1282,N_530,N_505);
nand U1283 (N_1283,N_922,N_616);
nand U1284 (N_1284,N_866,N_589);
or U1285 (N_1285,N_992,N_561);
nor U1286 (N_1286,N_953,N_637);
nand U1287 (N_1287,N_980,N_797);
and U1288 (N_1288,N_948,N_821);
nand U1289 (N_1289,N_766,N_593);
nand U1290 (N_1290,N_921,N_592);
and U1291 (N_1291,N_964,N_658);
and U1292 (N_1292,N_735,N_883);
and U1293 (N_1293,N_715,N_991);
nand U1294 (N_1294,N_775,N_856);
and U1295 (N_1295,N_515,N_638);
or U1296 (N_1296,N_534,N_628);
or U1297 (N_1297,N_800,N_542);
nand U1298 (N_1298,N_555,N_753);
and U1299 (N_1299,N_747,N_980);
nor U1300 (N_1300,N_715,N_624);
nor U1301 (N_1301,N_681,N_664);
or U1302 (N_1302,N_595,N_612);
and U1303 (N_1303,N_541,N_901);
nand U1304 (N_1304,N_661,N_686);
or U1305 (N_1305,N_802,N_986);
nor U1306 (N_1306,N_514,N_766);
or U1307 (N_1307,N_857,N_944);
and U1308 (N_1308,N_544,N_699);
nand U1309 (N_1309,N_675,N_575);
nand U1310 (N_1310,N_743,N_674);
nor U1311 (N_1311,N_828,N_920);
nand U1312 (N_1312,N_833,N_611);
nand U1313 (N_1313,N_700,N_755);
or U1314 (N_1314,N_930,N_970);
and U1315 (N_1315,N_963,N_594);
nor U1316 (N_1316,N_562,N_637);
nor U1317 (N_1317,N_889,N_950);
nor U1318 (N_1318,N_706,N_876);
nand U1319 (N_1319,N_605,N_641);
and U1320 (N_1320,N_736,N_771);
nor U1321 (N_1321,N_677,N_512);
and U1322 (N_1322,N_909,N_819);
nand U1323 (N_1323,N_867,N_681);
or U1324 (N_1324,N_559,N_849);
or U1325 (N_1325,N_792,N_815);
nand U1326 (N_1326,N_624,N_954);
and U1327 (N_1327,N_519,N_940);
nor U1328 (N_1328,N_793,N_764);
or U1329 (N_1329,N_936,N_649);
nand U1330 (N_1330,N_893,N_900);
nand U1331 (N_1331,N_635,N_901);
nand U1332 (N_1332,N_574,N_972);
or U1333 (N_1333,N_579,N_986);
nand U1334 (N_1334,N_700,N_846);
and U1335 (N_1335,N_699,N_640);
nand U1336 (N_1336,N_965,N_526);
or U1337 (N_1337,N_882,N_554);
nor U1338 (N_1338,N_673,N_527);
and U1339 (N_1339,N_813,N_655);
xnor U1340 (N_1340,N_737,N_730);
or U1341 (N_1341,N_798,N_634);
nor U1342 (N_1342,N_766,N_865);
nand U1343 (N_1343,N_718,N_533);
nor U1344 (N_1344,N_669,N_937);
or U1345 (N_1345,N_733,N_601);
and U1346 (N_1346,N_984,N_851);
and U1347 (N_1347,N_722,N_663);
and U1348 (N_1348,N_758,N_770);
or U1349 (N_1349,N_666,N_510);
and U1350 (N_1350,N_879,N_762);
nand U1351 (N_1351,N_517,N_942);
or U1352 (N_1352,N_909,N_820);
nand U1353 (N_1353,N_954,N_671);
xor U1354 (N_1354,N_596,N_503);
or U1355 (N_1355,N_671,N_806);
nor U1356 (N_1356,N_629,N_968);
or U1357 (N_1357,N_563,N_847);
and U1358 (N_1358,N_550,N_576);
and U1359 (N_1359,N_612,N_880);
nor U1360 (N_1360,N_554,N_540);
and U1361 (N_1361,N_626,N_863);
nand U1362 (N_1362,N_747,N_879);
nor U1363 (N_1363,N_507,N_587);
or U1364 (N_1364,N_706,N_789);
and U1365 (N_1365,N_987,N_939);
nand U1366 (N_1366,N_992,N_798);
nor U1367 (N_1367,N_794,N_862);
and U1368 (N_1368,N_946,N_627);
nand U1369 (N_1369,N_512,N_792);
or U1370 (N_1370,N_672,N_734);
nand U1371 (N_1371,N_862,N_825);
and U1372 (N_1372,N_736,N_651);
nor U1373 (N_1373,N_710,N_889);
nand U1374 (N_1374,N_675,N_940);
nand U1375 (N_1375,N_826,N_742);
or U1376 (N_1376,N_934,N_993);
and U1377 (N_1377,N_912,N_545);
and U1378 (N_1378,N_559,N_967);
nor U1379 (N_1379,N_604,N_602);
or U1380 (N_1380,N_931,N_893);
nor U1381 (N_1381,N_703,N_940);
or U1382 (N_1382,N_598,N_684);
and U1383 (N_1383,N_942,N_721);
or U1384 (N_1384,N_792,N_585);
or U1385 (N_1385,N_606,N_586);
and U1386 (N_1386,N_893,N_551);
or U1387 (N_1387,N_630,N_642);
nor U1388 (N_1388,N_945,N_826);
nor U1389 (N_1389,N_725,N_802);
or U1390 (N_1390,N_570,N_702);
nor U1391 (N_1391,N_795,N_632);
nor U1392 (N_1392,N_921,N_918);
and U1393 (N_1393,N_756,N_745);
nand U1394 (N_1394,N_836,N_578);
and U1395 (N_1395,N_997,N_725);
nand U1396 (N_1396,N_621,N_544);
nor U1397 (N_1397,N_550,N_962);
or U1398 (N_1398,N_912,N_524);
and U1399 (N_1399,N_943,N_606);
nand U1400 (N_1400,N_983,N_752);
and U1401 (N_1401,N_881,N_734);
or U1402 (N_1402,N_543,N_894);
nand U1403 (N_1403,N_623,N_929);
nand U1404 (N_1404,N_736,N_719);
nor U1405 (N_1405,N_808,N_714);
and U1406 (N_1406,N_809,N_787);
xor U1407 (N_1407,N_876,N_901);
nand U1408 (N_1408,N_722,N_528);
nand U1409 (N_1409,N_904,N_748);
and U1410 (N_1410,N_738,N_552);
nor U1411 (N_1411,N_951,N_716);
nand U1412 (N_1412,N_765,N_657);
or U1413 (N_1413,N_682,N_749);
or U1414 (N_1414,N_751,N_975);
and U1415 (N_1415,N_939,N_897);
xor U1416 (N_1416,N_647,N_980);
or U1417 (N_1417,N_735,N_527);
or U1418 (N_1418,N_992,N_838);
nor U1419 (N_1419,N_593,N_769);
nor U1420 (N_1420,N_532,N_676);
nand U1421 (N_1421,N_511,N_751);
xnor U1422 (N_1422,N_638,N_748);
or U1423 (N_1423,N_931,N_834);
and U1424 (N_1424,N_646,N_955);
or U1425 (N_1425,N_884,N_853);
nand U1426 (N_1426,N_805,N_891);
nand U1427 (N_1427,N_730,N_822);
and U1428 (N_1428,N_648,N_853);
or U1429 (N_1429,N_957,N_645);
nand U1430 (N_1430,N_891,N_506);
and U1431 (N_1431,N_852,N_805);
nand U1432 (N_1432,N_533,N_850);
nor U1433 (N_1433,N_793,N_913);
nand U1434 (N_1434,N_620,N_691);
nor U1435 (N_1435,N_833,N_668);
and U1436 (N_1436,N_506,N_901);
and U1437 (N_1437,N_941,N_992);
nand U1438 (N_1438,N_713,N_908);
and U1439 (N_1439,N_688,N_789);
and U1440 (N_1440,N_583,N_703);
xor U1441 (N_1441,N_916,N_502);
nand U1442 (N_1442,N_893,N_928);
nor U1443 (N_1443,N_970,N_884);
nand U1444 (N_1444,N_976,N_735);
or U1445 (N_1445,N_898,N_820);
nand U1446 (N_1446,N_589,N_746);
or U1447 (N_1447,N_511,N_748);
nor U1448 (N_1448,N_578,N_648);
nand U1449 (N_1449,N_951,N_548);
nor U1450 (N_1450,N_888,N_603);
nand U1451 (N_1451,N_938,N_522);
and U1452 (N_1452,N_890,N_651);
nor U1453 (N_1453,N_531,N_587);
and U1454 (N_1454,N_804,N_904);
nor U1455 (N_1455,N_648,N_985);
or U1456 (N_1456,N_836,N_556);
or U1457 (N_1457,N_615,N_957);
nor U1458 (N_1458,N_648,N_868);
nor U1459 (N_1459,N_977,N_820);
or U1460 (N_1460,N_959,N_846);
or U1461 (N_1461,N_709,N_584);
nor U1462 (N_1462,N_644,N_735);
nor U1463 (N_1463,N_902,N_767);
or U1464 (N_1464,N_683,N_815);
nand U1465 (N_1465,N_527,N_832);
or U1466 (N_1466,N_901,N_759);
nor U1467 (N_1467,N_560,N_912);
nor U1468 (N_1468,N_513,N_890);
nand U1469 (N_1469,N_893,N_967);
nor U1470 (N_1470,N_748,N_961);
or U1471 (N_1471,N_952,N_822);
nor U1472 (N_1472,N_914,N_848);
and U1473 (N_1473,N_603,N_784);
and U1474 (N_1474,N_892,N_600);
nand U1475 (N_1475,N_943,N_904);
nor U1476 (N_1476,N_802,N_537);
and U1477 (N_1477,N_990,N_790);
nor U1478 (N_1478,N_795,N_565);
or U1479 (N_1479,N_730,N_571);
nor U1480 (N_1480,N_711,N_934);
and U1481 (N_1481,N_646,N_978);
and U1482 (N_1482,N_509,N_773);
nand U1483 (N_1483,N_826,N_790);
nand U1484 (N_1484,N_818,N_867);
and U1485 (N_1485,N_801,N_930);
nor U1486 (N_1486,N_910,N_941);
nand U1487 (N_1487,N_963,N_914);
or U1488 (N_1488,N_912,N_634);
nor U1489 (N_1489,N_563,N_588);
nand U1490 (N_1490,N_759,N_810);
nor U1491 (N_1491,N_731,N_581);
and U1492 (N_1492,N_515,N_581);
and U1493 (N_1493,N_779,N_907);
nand U1494 (N_1494,N_989,N_504);
nor U1495 (N_1495,N_957,N_761);
and U1496 (N_1496,N_899,N_589);
or U1497 (N_1497,N_813,N_978);
and U1498 (N_1498,N_899,N_825);
nand U1499 (N_1499,N_951,N_928);
xnor U1500 (N_1500,N_1357,N_1128);
and U1501 (N_1501,N_1374,N_1102);
and U1502 (N_1502,N_1142,N_1344);
and U1503 (N_1503,N_1338,N_1148);
xor U1504 (N_1504,N_1440,N_1218);
nand U1505 (N_1505,N_1205,N_1144);
and U1506 (N_1506,N_1215,N_1348);
xnor U1507 (N_1507,N_1352,N_1345);
and U1508 (N_1508,N_1196,N_1353);
and U1509 (N_1509,N_1384,N_1254);
and U1510 (N_1510,N_1108,N_1233);
nand U1511 (N_1511,N_1434,N_1458);
or U1512 (N_1512,N_1069,N_1299);
nor U1513 (N_1513,N_1376,N_1214);
or U1514 (N_1514,N_1415,N_1267);
nand U1515 (N_1515,N_1258,N_1307);
nor U1516 (N_1516,N_1208,N_1221);
or U1517 (N_1517,N_1043,N_1400);
nor U1518 (N_1518,N_1492,N_1136);
or U1519 (N_1519,N_1485,N_1068);
nor U1520 (N_1520,N_1279,N_1422);
nand U1521 (N_1521,N_1073,N_1427);
nor U1522 (N_1522,N_1182,N_1217);
and U1523 (N_1523,N_1119,N_1240);
nor U1524 (N_1524,N_1096,N_1029);
nand U1525 (N_1525,N_1014,N_1364);
nand U1526 (N_1526,N_1482,N_1220);
or U1527 (N_1527,N_1253,N_1245);
and U1528 (N_1528,N_1388,N_1405);
and U1529 (N_1529,N_1126,N_1152);
or U1530 (N_1530,N_1235,N_1448);
nor U1531 (N_1531,N_1171,N_1329);
or U1532 (N_1532,N_1019,N_1351);
nand U1533 (N_1533,N_1391,N_1060);
nor U1534 (N_1534,N_1457,N_1012);
xor U1535 (N_1535,N_1410,N_1334);
nand U1536 (N_1536,N_1354,N_1179);
xnor U1537 (N_1537,N_1127,N_1450);
nand U1538 (N_1538,N_1264,N_1439);
and U1539 (N_1539,N_1383,N_1447);
nand U1540 (N_1540,N_1495,N_1487);
or U1541 (N_1541,N_1035,N_1170);
nand U1542 (N_1542,N_1370,N_1257);
and U1543 (N_1543,N_1079,N_1356);
nor U1544 (N_1544,N_1222,N_1067);
or U1545 (N_1545,N_1163,N_1046);
and U1546 (N_1546,N_1207,N_1135);
and U1547 (N_1547,N_1286,N_1032);
nor U1548 (N_1548,N_1187,N_1028);
or U1549 (N_1549,N_1022,N_1049);
nand U1550 (N_1550,N_1349,N_1494);
nand U1551 (N_1551,N_1411,N_1341);
or U1552 (N_1552,N_1275,N_1438);
nand U1553 (N_1553,N_1365,N_1030);
and U1554 (N_1554,N_1201,N_1191);
nor U1555 (N_1555,N_1092,N_1330);
or U1556 (N_1556,N_1038,N_1403);
or U1557 (N_1557,N_1333,N_1003);
or U1558 (N_1558,N_1317,N_1483);
and U1559 (N_1559,N_1442,N_1099);
nand U1560 (N_1560,N_1057,N_1313);
nand U1561 (N_1561,N_1204,N_1390);
nor U1562 (N_1562,N_1074,N_1355);
xnor U1563 (N_1563,N_1146,N_1117);
xor U1564 (N_1564,N_1430,N_1291);
nand U1565 (N_1565,N_1072,N_1282);
nor U1566 (N_1566,N_1089,N_1005);
nand U1567 (N_1567,N_1467,N_1015);
nand U1568 (N_1568,N_1292,N_1158);
nor U1569 (N_1569,N_1475,N_1017);
nand U1570 (N_1570,N_1001,N_1070);
nand U1571 (N_1571,N_1496,N_1386);
and U1572 (N_1572,N_1155,N_1219);
and U1573 (N_1573,N_1104,N_1431);
nand U1574 (N_1574,N_1284,N_1466);
nand U1575 (N_1575,N_1407,N_1036);
and U1576 (N_1576,N_1443,N_1369);
nand U1577 (N_1577,N_1472,N_1160);
and U1578 (N_1578,N_1133,N_1193);
nor U1579 (N_1579,N_1236,N_1167);
nor U1580 (N_1580,N_1200,N_1413);
nor U1581 (N_1581,N_1223,N_1209);
nand U1582 (N_1582,N_1414,N_1086);
nand U1583 (N_1583,N_1302,N_1326);
and U1584 (N_1584,N_1381,N_1016);
xor U1585 (N_1585,N_1285,N_1190);
and U1586 (N_1586,N_1259,N_1296);
nand U1587 (N_1587,N_1082,N_1412);
and U1588 (N_1588,N_1361,N_1094);
nand U1589 (N_1589,N_1402,N_1100);
and U1590 (N_1590,N_1062,N_1417);
nand U1591 (N_1591,N_1024,N_1168);
or U1592 (N_1592,N_1047,N_1262);
or U1593 (N_1593,N_1106,N_1123);
xor U1594 (N_1594,N_1175,N_1323);
and U1595 (N_1595,N_1396,N_1394);
nor U1596 (N_1596,N_1159,N_1452);
nor U1597 (N_1597,N_1366,N_1423);
or U1598 (N_1598,N_1425,N_1037);
nor U1599 (N_1599,N_1061,N_1229);
and U1600 (N_1600,N_1121,N_1371);
nand U1601 (N_1601,N_1143,N_1301);
nand U1602 (N_1602,N_1056,N_1116);
and U1603 (N_1603,N_1319,N_1164);
nand U1604 (N_1604,N_1419,N_1234);
nor U1605 (N_1605,N_1436,N_1137);
and U1606 (N_1606,N_1195,N_1304);
or U1607 (N_1607,N_1198,N_1033);
nor U1608 (N_1608,N_1004,N_1406);
xor U1609 (N_1609,N_1461,N_1125);
or U1610 (N_1610,N_1327,N_1449);
nor U1611 (N_1611,N_1109,N_1178);
nand U1612 (N_1612,N_1098,N_1080);
nand U1613 (N_1613,N_1031,N_1465);
and U1614 (N_1614,N_1263,N_1310);
or U1615 (N_1615,N_1150,N_1339);
nor U1616 (N_1616,N_1145,N_1273);
and U1617 (N_1617,N_1210,N_1122);
or U1618 (N_1618,N_1241,N_1071);
nand U1619 (N_1619,N_1020,N_1249);
and U1620 (N_1620,N_1295,N_1097);
and U1621 (N_1621,N_1387,N_1053);
nor U1622 (N_1622,N_1139,N_1078);
and U1623 (N_1623,N_1230,N_1045);
or U1624 (N_1624,N_1320,N_1260);
nand U1625 (N_1625,N_1256,N_1088);
and U1626 (N_1626,N_1293,N_1156);
nor U1627 (N_1627,N_1459,N_1130);
and U1628 (N_1628,N_1007,N_1213);
nor U1629 (N_1629,N_1373,N_1276);
nand U1630 (N_1630,N_1059,N_1114);
and U1631 (N_1631,N_1244,N_1120);
nor U1632 (N_1632,N_1397,N_1322);
nand U1633 (N_1633,N_1184,N_1473);
and U1634 (N_1634,N_1281,N_1277);
nor U1635 (N_1635,N_1469,N_1451);
nand U1636 (N_1636,N_1489,N_1006);
and U1637 (N_1637,N_1476,N_1034);
nor U1638 (N_1638,N_1392,N_1342);
nand U1639 (N_1639,N_1358,N_1134);
and U1640 (N_1640,N_1157,N_1497);
and U1641 (N_1641,N_1382,N_1379);
nor U1642 (N_1642,N_1328,N_1261);
nor U1643 (N_1643,N_1008,N_1308);
nand U1644 (N_1644,N_1471,N_1231);
or U1645 (N_1645,N_1010,N_1271);
nor U1646 (N_1646,N_1360,N_1445);
and U1647 (N_1647,N_1147,N_1112);
and U1648 (N_1648,N_1237,N_1181);
nor U1649 (N_1649,N_1018,N_1224);
nor U1650 (N_1650,N_1149,N_1162);
and U1651 (N_1651,N_1493,N_1435);
nand U1652 (N_1652,N_1305,N_1194);
nor U1653 (N_1653,N_1081,N_1336);
and U1654 (N_1654,N_1332,N_1199);
and U1655 (N_1655,N_1270,N_1300);
and U1656 (N_1656,N_1027,N_1474);
and U1657 (N_1657,N_1232,N_1380);
nor U1658 (N_1658,N_1206,N_1021);
or U1659 (N_1659,N_1189,N_1183);
nor U1660 (N_1660,N_1129,N_1166);
nor U1661 (N_1661,N_1077,N_1491);
and U1662 (N_1662,N_1470,N_1481);
and U1663 (N_1663,N_1176,N_1227);
or U1664 (N_1664,N_1343,N_1346);
nor U1665 (N_1665,N_1479,N_1453);
or U1666 (N_1666,N_1363,N_1103);
nor U1667 (N_1667,N_1278,N_1362);
nand U1668 (N_1668,N_1076,N_1314);
or U1669 (N_1669,N_1424,N_1052);
nor U1670 (N_1670,N_1367,N_1311);
nor U1671 (N_1671,N_1478,N_1454);
and U1672 (N_1672,N_1186,N_1289);
nor U1673 (N_1673,N_1177,N_1058);
or U1674 (N_1674,N_1420,N_1255);
nor U1675 (N_1675,N_1173,N_1226);
xnor U1676 (N_1676,N_1404,N_1246);
nand U1677 (N_1677,N_1401,N_1083);
or U1678 (N_1678,N_1228,N_1303);
and U1679 (N_1679,N_1013,N_1188);
xor U1680 (N_1680,N_1324,N_1375);
and U1681 (N_1681,N_1272,N_1131);
nand U1682 (N_1682,N_1238,N_1247);
nand U1683 (N_1683,N_1151,N_1274);
nand U1684 (N_1684,N_1460,N_1075);
or U1685 (N_1685,N_1115,N_1161);
and U1686 (N_1686,N_1216,N_1490);
nand U1687 (N_1687,N_1084,N_1153);
or U1688 (N_1688,N_1118,N_1321);
or U1689 (N_1689,N_1197,N_1368);
and U1690 (N_1690,N_1337,N_1040);
or U1691 (N_1691,N_1389,N_1185);
nand U1692 (N_1692,N_1064,N_1251);
nand U1693 (N_1693,N_1023,N_1347);
and U1694 (N_1694,N_1087,N_1093);
or U1695 (N_1695,N_1331,N_1002);
nand U1696 (N_1696,N_1372,N_1340);
nand U1697 (N_1697,N_1456,N_1312);
nor U1698 (N_1698,N_1265,N_1429);
and U1699 (N_1699,N_1172,N_1416);
nand U1700 (N_1700,N_1174,N_1066);
and U1701 (N_1701,N_1165,N_1000);
and U1702 (N_1702,N_1225,N_1306);
or U1703 (N_1703,N_1202,N_1441);
or U1704 (N_1704,N_1464,N_1192);
nor U1705 (N_1705,N_1433,N_1252);
nor U1706 (N_1706,N_1318,N_1107);
or U1707 (N_1707,N_1211,N_1280);
nand U1708 (N_1708,N_1063,N_1044);
nand U1709 (N_1709,N_1426,N_1283);
and U1710 (N_1710,N_1011,N_1385);
or U1711 (N_1711,N_1141,N_1042);
nor U1712 (N_1712,N_1051,N_1054);
and U1713 (N_1713,N_1085,N_1335);
nand U1714 (N_1714,N_1110,N_1239);
and U1715 (N_1715,N_1250,N_1203);
nand U1716 (N_1716,N_1446,N_1399);
nor U1717 (N_1717,N_1444,N_1325);
or U1718 (N_1718,N_1242,N_1294);
and U1719 (N_1719,N_1039,N_1359);
and U1720 (N_1720,N_1050,N_1169);
nor U1721 (N_1721,N_1154,N_1499);
and U1722 (N_1722,N_1398,N_1065);
and U1723 (N_1723,N_1418,N_1498);
and U1724 (N_1724,N_1428,N_1455);
and U1725 (N_1725,N_1288,N_1132);
and U1726 (N_1726,N_1350,N_1484);
nor U1727 (N_1727,N_1138,N_1048);
and U1728 (N_1728,N_1180,N_1316);
nand U1729 (N_1729,N_1268,N_1124);
nand U1730 (N_1730,N_1463,N_1243);
nor U1731 (N_1731,N_1290,N_1378);
or U1732 (N_1732,N_1377,N_1468);
or U1733 (N_1733,N_1432,N_1140);
and U1734 (N_1734,N_1009,N_1101);
and U1735 (N_1735,N_1409,N_1488);
and U1736 (N_1736,N_1025,N_1212);
nand U1737 (N_1737,N_1480,N_1041);
nor U1738 (N_1738,N_1269,N_1287);
nand U1739 (N_1739,N_1111,N_1297);
nor U1740 (N_1740,N_1090,N_1248);
nand U1741 (N_1741,N_1393,N_1105);
nand U1742 (N_1742,N_1315,N_1298);
or U1743 (N_1743,N_1437,N_1421);
and U1744 (N_1744,N_1309,N_1486);
nand U1745 (N_1745,N_1462,N_1091);
nor U1746 (N_1746,N_1408,N_1026);
and U1747 (N_1747,N_1095,N_1395);
nand U1748 (N_1748,N_1055,N_1113);
nand U1749 (N_1749,N_1266,N_1477);
nand U1750 (N_1750,N_1001,N_1484);
or U1751 (N_1751,N_1121,N_1321);
and U1752 (N_1752,N_1466,N_1268);
nand U1753 (N_1753,N_1491,N_1215);
nor U1754 (N_1754,N_1328,N_1349);
nor U1755 (N_1755,N_1276,N_1016);
nor U1756 (N_1756,N_1320,N_1293);
nand U1757 (N_1757,N_1093,N_1403);
xnor U1758 (N_1758,N_1117,N_1031);
or U1759 (N_1759,N_1223,N_1098);
nor U1760 (N_1760,N_1166,N_1275);
or U1761 (N_1761,N_1123,N_1171);
and U1762 (N_1762,N_1235,N_1383);
nand U1763 (N_1763,N_1390,N_1383);
nor U1764 (N_1764,N_1351,N_1185);
nor U1765 (N_1765,N_1381,N_1276);
or U1766 (N_1766,N_1229,N_1250);
nor U1767 (N_1767,N_1198,N_1015);
nor U1768 (N_1768,N_1446,N_1411);
or U1769 (N_1769,N_1296,N_1322);
nor U1770 (N_1770,N_1095,N_1109);
and U1771 (N_1771,N_1159,N_1064);
nand U1772 (N_1772,N_1254,N_1051);
nor U1773 (N_1773,N_1386,N_1405);
and U1774 (N_1774,N_1284,N_1495);
and U1775 (N_1775,N_1426,N_1083);
nor U1776 (N_1776,N_1092,N_1476);
and U1777 (N_1777,N_1250,N_1497);
nand U1778 (N_1778,N_1330,N_1271);
or U1779 (N_1779,N_1056,N_1389);
nor U1780 (N_1780,N_1293,N_1134);
nand U1781 (N_1781,N_1350,N_1394);
or U1782 (N_1782,N_1146,N_1462);
nand U1783 (N_1783,N_1043,N_1386);
nand U1784 (N_1784,N_1083,N_1453);
xor U1785 (N_1785,N_1172,N_1263);
nor U1786 (N_1786,N_1478,N_1331);
nand U1787 (N_1787,N_1041,N_1342);
nor U1788 (N_1788,N_1099,N_1002);
nand U1789 (N_1789,N_1047,N_1198);
or U1790 (N_1790,N_1208,N_1361);
nand U1791 (N_1791,N_1103,N_1155);
nand U1792 (N_1792,N_1127,N_1063);
or U1793 (N_1793,N_1084,N_1478);
or U1794 (N_1794,N_1059,N_1417);
nand U1795 (N_1795,N_1088,N_1435);
or U1796 (N_1796,N_1080,N_1318);
and U1797 (N_1797,N_1236,N_1393);
or U1798 (N_1798,N_1203,N_1128);
or U1799 (N_1799,N_1150,N_1391);
or U1800 (N_1800,N_1031,N_1021);
nor U1801 (N_1801,N_1210,N_1002);
nand U1802 (N_1802,N_1109,N_1368);
or U1803 (N_1803,N_1357,N_1115);
and U1804 (N_1804,N_1488,N_1293);
or U1805 (N_1805,N_1384,N_1238);
and U1806 (N_1806,N_1254,N_1180);
nand U1807 (N_1807,N_1396,N_1415);
nor U1808 (N_1808,N_1333,N_1454);
nand U1809 (N_1809,N_1172,N_1097);
nor U1810 (N_1810,N_1383,N_1250);
nor U1811 (N_1811,N_1000,N_1403);
or U1812 (N_1812,N_1010,N_1285);
nand U1813 (N_1813,N_1031,N_1048);
or U1814 (N_1814,N_1360,N_1160);
nor U1815 (N_1815,N_1183,N_1429);
or U1816 (N_1816,N_1042,N_1498);
or U1817 (N_1817,N_1439,N_1445);
nand U1818 (N_1818,N_1423,N_1122);
and U1819 (N_1819,N_1326,N_1184);
nor U1820 (N_1820,N_1465,N_1193);
nand U1821 (N_1821,N_1349,N_1330);
nor U1822 (N_1822,N_1473,N_1377);
or U1823 (N_1823,N_1194,N_1165);
nor U1824 (N_1824,N_1178,N_1056);
nor U1825 (N_1825,N_1469,N_1084);
nand U1826 (N_1826,N_1018,N_1465);
and U1827 (N_1827,N_1311,N_1094);
nand U1828 (N_1828,N_1433,N_1269);
nor U1829 (N_1829,N_1277,N_1090);
nor U1830 (N_1830,N_1136,N_1190);
nand U1831 (N_1831,N_1309,N_1187);
or U1832 (N_1832,N_1277,N_1206);
or U1833 (N_1833,N_1337,N_1235);
nor U1834 (N_1834,N_1253,N_1192);
and U1835 (N_1835,N_1397,N_1345);
nand U1836 (N_1836,N_1485,N_1060);
nor U1837 (N_1837,N_1186,N_1093);
nor U1838 (N_1838,N_1338,N_1119);
or U1839 (N_1839,N_1485,N_1131);
or U1840 (N_1840,N_1010,N_1398);
nand U1841 (N_1841,N_1147,N_1227);
xnor U1842 (N_1842,N_1207,N_1440);
nor U1843 (N_1843,N_1033,N_1357);
or U1844 (N_1844,N_1226,N_1460);
or U1845 (N_1845,N_1029,N_1411);
and U1846 (N_1846,N_1110,N_1184);
or U1847 (N_1847,N_1139,N_1484);
nor U1848 (N_1848,N_1252,N_1122);
nand U1849 (N_1849,N_1127,N_1186);
nor U1850 (N_1850,N_1022,N_1293);
nor U1851 (N_1851,N_1437,N_1101);
or U1852 (N_1852,N_1307,N_1361);
nor U1853 (N_1853,N_1001,N_1276);
nand U1854 (N_1854,N_1393,N_1489);
or U1855 (N_1855,N_1083,N_1434);
and U1856 (N_1856,N_1011,N_1071);
nor U1857 (N_1857,N_1380,N_1243);
nor U1858 (N_1858,N_1072,N_1082);
and U1859 (N_1859,N_1458,N_1476);
or U1860 (N_1860,N_1083,N_1021);
nand U1861 (N_1861,N_1033,N_1129);
or U1862 (N_1862,N_1050,N_1453);
nor U1863 (N_1863,N_1343,N_1192);
nand U1864 (N_1864,N_1213,N_1018);
nor U1865 (N_1865,N_1215,N_1043);
or U1866 (N_1866,N_1194,N_1268);
nand U1867 (N_1867,N_1040,N_1048);
nand U1868 (N_1868,N_1442,N_1473);
nor U1869 (N_1869,N_1421,N_1130);
nor U1870 (N_1870,N_1066,N_1275);
nand U1871 (N_1871,N_1091,N_1409);
or U1872 (N_1872,N_1443,N_1461);
or U1873 (N_1873,N_1092,N_1370);
nand U1874 (N_1874,N_1335,N_1450);
nand U1875 (N_1875,N_1316,N_1439);
nand U1876 (N_1876,N_1358,N_1299);
or U1877 (N_1877,N_1481,N_1106);
and U1878 (N_1878,N_1402,N_1371);
xnor U1879 (N_1879,N_1237,N_1063);
or U1880 (N_1880,N_1087,N_1086);
and U1881 (N_1881,N_1112,N_1398);
nor U1882 (N_1882,N_1122,N_1027);
nor U1883 (N_1883,N_1035,N_1231);
or U1884 (N_1884,N_1159,N_1320);
or U1885 (N_1885,N_1271,N_1156);
nand U1886 (N_1886,N_1467,N_1155);
nand U1887 (N_1887,N_1339,N_1037);
nand U1888 (N_1888,N_1277,N_1169);
nor U1889 (N_1889,N_1290,N_1266);
xnor U1890 (N_1890,N_1240,N_1421);
nor U1891 (N_1891,N_1043,N_1430);
and U1892 (N_1892,N_1272,N_1018);
nor U1893 (N_1893,N_1092,N_1002);
nand U1894 (N_1894,N_1078,N_1372);
or U1895 (N_1895,N_1167,N_1439);
nor U1896 (N_1896,N_1153,N_1276);
and U1897 (N_1897,N_1052,N_1247);
nor U1898 (N_1898,N_1386,N_1053);
xor U1899 (N_1899,N_1081,N_1019);
or U1900 (N_1900,N_1453,N_1060);
or U1901 (N_1901,N_1320,N_1220);
or U1902 (N_1902,N_1192,N_1013);
or U1903 (N_1903,N_1027,N_1041);
and U1904 (N_1904,N_1218,N_1153);
or U1905 (N_1905,N_1108,N_1009);
and U1906 (N_1906,N_1091,N_1208);
nor U1907 (N_1907,N_1396,N_1120);
or U1908 (N_1908,N_1191,N_1087);
nand U1909 (N_1909,N_1156,N_1261);
nand U1910 (N_1910,N_1231,N_1067);
xnor U1911 (N_1911,N_1170,N_1073);
or U1912 (N_1912,N_1180,N_1051);
and U1913 (N_1913,N_1493,N_1285);
nor U1914 (N_1914,N_1056,N_1101);
nand U1915 (N_1915,N_1330,N_1355);
nand U1916 (N_1916,N_1198,N_1494);
or U1917 (N_1917,N_1056,N_1421);
and U1918 (N_1918,N_1471,N_1016);
or U1919 (N_1919,N_1427,N_1418);
nor U1920 (N_1920,N_1186,N_1411);
or U1921 (N_1921,N_1459,N_1386);
or U1922 (N_1922,N_1080,N_1099);
and U1923 (N_1923,N_1019,N_1365);
and U1924 (N_1924,N_1141,N_1434);
nor U1925 (N_1925,N_1327,N_1026);
or U1926 (N_1926,N_1106,N_1389);
and U1927 (N_1927,N_1408,N_1238);
and U1928 (N_1928,N_1485,N_1061);
nand U1929 (N_1929,N_1336,N_1073);
nand U1930 (N_1930,N_1135,N_1453);
or U1931 (N_1931,N_1494,N_1034);
nand U1932 (N_1932,N_1216,N_1123);
or U1933 (N_1933,N_1064,N_1112);
xnor U1934 (N_1934,N_1122,N_1082);
and U1935 (N_1935,N_1143,N_1090);
and U1936 (N_1936,N_1128,N_1417);
and U1937 (N_1937,N_1134,N_1143);
nand U1938 (N_1938,N_1072,N_1256);
nor U1939 (N_1939,N_1057,N_1292);
nor U1940 (N_1940,N_1454,N_1073);
and U1941 (N_1941,N_1405,N_1403);
nand U1942 (N_1942,N_1368,N_1012);
nor U1943 (N_1943,N_1351,N_1006);
nor U1944 (N_1944,N_1082,N_1184);
and U1945 (N_1945,N_1179,N_1166);
nor U1946 (N_1946,N_1001,N_1128);
or U1947 (N_1947,N_1115,N_1226);
nand U1948 (N_1948,N_1411,N_1464);
and U1949 (N_1949,N_1363,N_1256);
or U1950 (N_1950,N_1120,N_1207);
nand U1951 (N_1951,N_1310,N_1021);
and U1952 (N_1952,N_1149,N_1134);
or U1953 (N_1953,N_1437,N_1322);
or U1954 (N_1954,N_1115,N_1401);
nor U1955 (N_1955,N_1464,N_1306);
nor U1956 (N_1956,N_1181,N_1156);
and U1957 (N_1957,N_1205,N_1441);
nor U1958 (N_1958,N_1159,N_1325);
or U1959 (N_1959,N_1440,N_1090);
and U1960 (N_1960,N_1155,N_1133);
and U1961 (N_1961,N_1306,N_1494);
nand U1962 (N_1962,N_1408,N_1315);
or U1963 (N_1963,N_1176,N_1381);
nand U1964 (N_1964,N_1497,N_1094);
and U1965 (N_1965,N_1396,N_1469);
or U1966 (N_1966,N_1126,N_1161);
nand U1967 (N_1967,N_1196,N_1221);
nor U1968 (N_1968,N_1260,N_1173);
nor U1969 (N_1969,N_1229,N_1107);
nor U1970 (N_1970,N_1215,N_1478);
nor U1971 (N_1971,N_1008,N_1371);
nand U1972 (N_1972,N_1129,N_1189);
or U1973 (N_1973,N_1473,N_1472);
nor U1974 (N_1974,N_1234,N_1201);
and U1975 (N_1975,N_1352,N_1047);
and U1976 (N_1976,N_1352,N_1480);
nor U1977 (N_1977,N_1230,N_1023);
nand U1978 (N_1978,N_1282,N_1243);
nand U1979 (N_1979,N_1350,N_1235);
nand U1980 (N_1980,N_1279,N_1433);
or U1981 (N_1981,N_1161,N_1038);
nand U1982 (N_1982,N_1185,N_1440);
nor U1983 (N_1983,N_1139,N_1420);
and U1984 (N_1984,N_1171,N_1246);
and U1985 (N_1985,N_1347,N_1327);
nand U1986 (N_1986,N_1390,N_1361);
and U1987 (N_1987,N_1290,N_1377);
nor U1988 (N_1988,N_1453,N_1216);
and U1989 (N_1989,N_1395,N_1196);
nand U1990 (N_1990,N_1227,N_1168);
nor U1991 (N_1991,N_1369,N_1088);
nand U1992 (N_1992,N_1369,N_1026);
and U1993 (N_1993,N_1466,N_1137);
xnor U1994 (N_1994,N_1045,N_1007);
nand U1995 (N_1995,N_1392,N_1380);
nand U1996 (N_1996,N_1190,N_1206);
and U1997 (N_1997,N_1082,N_1069);
and U1998 (N_1998,N_1113,N_1237);
xnor U1999 (N_1999,N_1086,N_1490);
or U2000 (N_2000,N_1671,N_1979);
nand U2001 (N_2001,N_1756,N_1903);
nor U2002 (N_2002,N_1964,N_1775);
and U2003 (N_2003,N_1922,N_1956);
nor U2004 (N_2004,N_1622,N_1628);
xnor U2005 (N_2005,N_1914,N_1777);
and U2006 (N_2006,N_1550,N_1716);
or U2007 (N_2007,N_1978,N_1860);
nand U2008 (N_2008,N_1508,N_1613);
nand U2009 (N_2009,N_1990,N_1534);
nor U2010 (N_2010,N_1941,N_1778);
or U2011 (N_2011,N_1981,N_1538);
nor U2012 (N_2012,N_1806,N_1863);
or U2013 (N_2013,N_1760,N_1834);
and U2014 (N_2014,N_1604,N_1839);
or U2015 (N_2015,N_1676,N_1629);
nand U2016 (N_2016,N_1901,N_1561);
nor U2017 (N_2017,N_1967,N_1663);
and U2018 (N_2018,N_1747,N_1723);
nor U2019 (N_2019,N_1845,N_1898);
nand U2020 (N_2020,N_1578,N_1678);
nor U2021 (N_2021,N_1969,N_1951);
nor U2022 (N_2022,N_1531,N_1603);
or U2023 (N_2023,N_1579,N_1892);
xnor U2024 (N_2024,N_1985,N_1942);
or U2025 (N_2025,N_1817,N_1692);
or U2026 (N_2026,N_1635,N_1795);
or U2027 (N_2027,N_1709,N_1543);
or U2028 (N_2028,N_1615,N_1877);
or U2029 (N_2029,N_1848,N_1913);
and U2030 (N_2030,N_1606,N_1896);
nor U2031 (N_2031,N_1961,N_1626);
and U2032 (N_2032,N_1646,N_1642);
or U2033 (N_2033,N_1900,N_1734);
and U2034 (N_2034,N_1955,N_1510);
nor U2035 (N_2035,N_1544,N_1590);
xnor U2036 (N_2036,N_1746,N_1878);
or U2037 (N_2037,N_1682,N_1876);
or U2038 (N_2038,N_1827,N_1562);
or U2039 (N_2039,N_1673,N_1593);
nand U2040 (N_2040,N_1844,N_1623);
nor U2041 (N_2041,N_1809,N_1702);
and U2042 (N_2042,N_1779,N_1825);
nand U2043 (N_2043,N_1584,N_1596);
nand U2044 (N_2044,N_1754,N_1840);
nand U2045 (N_2045,N_1588,N_1713);
and U2046 (N_2046,N_1767,N_1652);
or U2047 (N_2047,N_1665,N_1826);
nand U2048 (N_2048,N_1897,N_1935);
nor U2049 (N_2049,N_1759,N_1998);
nor U2050 (N_2050,N_1851,N_1977);
or U2051 (N_2051,N_1614,N_1943);
xnor U2052 (N_2052,N_1973,N_1949);
nor U2053 (N_2053,N_1743,N_1572);
nand U2054 (N_2054,N_1835,N_1636);
nor U2055 (N_2055,N_1703,N_1776);
and U2056 (N_2056,N_1651,N_1980);
and U2057 (N_2057,N_1810,N_1733);
nor U2058 (N_2058,N_1624,N_1755);
and U2059 (N_2059,N_1854,N_1698);
or U2060 (N_2060,N_1947,N_1830);
nor U2061 (N_2061,N_1822,N_1905);
nor U2062 (N_2062,N_1974,N_1871);
nor U2063 (N_2063,N_1783,N_1660);
or U2064 (N_2064,N_1563,N_1730);
nand U2065 (N_2065,N_1565,N_1855);
and U2066 (N_2066,N_1946,N_1766);
nor U2067 (N_2067,N_1794,N_1714);
nor U2068 (N_2068,N_1558,N_1971);
nor U2069 (N_2069,N_1894,N_1881);
and U2070 (N_2070,N_1735,N_1966);
nor U2071 (N_2071,N_1654,N_1753);
and U2072 (N_2072,N_1884,N_1571);
nor U2073 (N_2073,N_1551,N_1939);
nor U2074 (N_2074,N_1643,N_1736);
or U2075 (N_2075,N_1828,N_1582);
nand U2076 (N_2076,N_1886,N_1532);
nand U2077 (N_2077,N_1731,N_1518);
nor U2078 (N_2078,N_1683,N_1972);
nand U2079 (N_2079,N_1690,N_1514);
or U2080 (N_2080,N_1920,N_1983);
or U2081 (N_2081,N_1540,N_1772);
and U2082 (N_2082,N_1539,N_1798);
and U2083 (N_2083,N_1704,N_1616);
nor U2084 (N_2084,N_1824,N_1658);
or U2085 (N_2085,N_1793,N_1918);
nand U2086 (N_2086,N_1960,N_1814);
nor U2087 (N_2087,N_1899,N_1668);
and U2088 (N_2088,N_1869,N_1748);
nand U2089 (N_2089,N_1675,N_1750);
and U2090 (N_2090,N_1792,N_1988);
nand U2091 (N_2091,N_1823,N_1535);
nor U2092 (N_2092,N_1502,N_1577);
or U2093 (N_2093,N_1653,N_1926);
nand U2094 (N_2094,N_1936,N_1799);
xor U2095 (N_2095,N_1545,N_1929);
xor U2096 (N_2096,N_1583,N_1568);
and U2097 (N_2097,N_1890,N_1986);
or U2098 (N_2098,N_1501,N_1873);
nor U2099 (N_2099,N_1962,N_1993);
xnor U2100 (N_2100,N_1933,N_1711);
xor U2101 (N_2101,N_1728,N_1803);
or U2102 (N_2102,N_1987,N_1959);
nand U2103 (N_2103,N_1630,N_1696);
nor U2104 (N_2104,N_1589,N_1891);
or U2105 (N_2105,N_1925,N_1526);
or U2106 (N_2106,N_1618,N_1576);
nor U2107 (N_2107,N_1764,N_1557);
and U2108 (N_2108,N_1677,N_1507);
and U2109 (N_2109,N_1601,N_1849);
or U2110 (N_2110,N_1525,N_1564);
or U2111 (N_2111,N_1742,N_1740);
and U2112 (N_2112,N_1994,N_1511);
and U2113 (N_2113,N_1811,N_1715);
and U2114 (N_2114,N_1529,N_1607);
or U2115 (N_2115,N_1989,N_1634);
and U2116 (N_2116,N_1857,N_1627);
nand U2117 (N_2117,N_1852,N_1732);
or U2118 (N_2118,N_1608,N_1940);
xor U2119 (N_2119,N_1705,N_1841);
nor U2120 (N_2120,N_1695,N_1672);
and U2121 (N_2121,N_1975,N_1659);
nand U2122 (N_2122,N_1808,N_1575);
and U2123 (N_2123,N_1552,N_1952);
or U2124 (N_2124,N_1739,N_1587);
or U2125 (N_2125,N_1512,N_1697);
nand U2126 (N_2126,N_1681,N_1684);
or U2127 (N_2127,N_1997,N_1694);
nand U2128 (N_2128,N_1815,N_1519);
nor U2129 (N_2129,N_1717,N_1667);
or U2130 (N_2130,N_1887,N_1641);
or U2131 (N_2131,N_1982,N_1797);
xnor U2132 (N_2132,N_1829,N_1882);
nand U2133 (N_2133,N_1872,N_1609);
nand U2134 (N_2134,N_1533,N_1586);
and U2135 (N_2135,N_1765,N_1595);
nand U2136 (N_2136,N_1515,N_1761);
nor U2137 (N_2137,N_1948,N_1687);
and U2138 (N_2138,N_1693,N_1908);
xor U2139 (N_2139,N_1738,N_1996);
nor U2140 (N_2140,N_1724,N_1885);
or U2141 (N_2141,N_1784,N_1640);
and U2142 (N_2142,N_1812,N_1611);
or U2143 (N_2143,N_1859,N_1954);
nand U2144 (N_2144,N_1927,N_1720);
or U2145 (N_2145,N_1602,N_1883);
xor U2146 (N_2146,N_1820,N_1520);
and U2147 (N_2147,N_1867,N_1560);
nand U2148 (N_2148,N_1866,N_1836);
nor U2149 (N_2149,N_1553,N_1712);
and U2150 (N_2150,N_1580,N_1895);
and U2151 (N_2151,N_1774,N_1707);
nor U2152 (N_2152,N_1699,N_1548);
xor U2153 (N_2153,N_1649,N_1541);
nand U2154 (N_2154,N_1605,N_1727);
nand U2155 (N_2155,N_1581,N_1843);
nand U2156 (N_2156,N_1556,N_1637);
and U2157 (N_2157,N_1600,N_1610);
or U2158 (N_2158,N_1680,N_1633);
nand U2159 (N_2159,N_1970,N_1864);
nor U2160 (N_2160,N_1710,N_1865);
or U2161 (N_2161,N_1786,N_1912);
and U2162 (N_2162,N_1632,N_1800);
nor U2163 (N_2163,N_1757,N_1638);
and U2164 (N_2164,N_1500,N_1957);
and U2165 (N_2165,N_1991,N_1995);
or U2166 (N_2166,N_1874,N_1932);
nand U2167 (N_2167,N_1612,N_1506);
and U2168 (N_2168,N_1685,N_1968);
nor U2169 (N_2169,N_1549,N_1537);
nor U2170 (N_2170,N_1770,N_1700);
and U2171 (N_2171,N_1833,N_1505);
nor U2172 (N_2172,N_1664,N_1819);
or U2173 (N_2173,N_1782,N_1617);
or U2174 (N_2174,N_1984,N_1679);
and U2175 (N_2175,N_1796,N_1513);
and U2176 (N_2176,N_1842,N_1689);
nand U2177 (N_2177,N_1846,N_1911);
or U2178 (N_2178,N_1893,N_1861);
nand U2179 (N_2179,N_1928,N_1751);
nand U2180 (N_2180,N_1701,N_1858);
nand U2181 (N_2181,N_1801,N_1523);
and U2182 (N_2182,N_1522,N_1921);
nand U2183 (N_2183,N_1787,N_1771);
and U2184 (N_2184,N_1818,N_1645);
nand U2185 (N_2185,N_1773,N_1569);
or U2186 (N_2186,N_1938,N_1945);
and U2187 (N_2187,N_1503,N_1788);
or U2188 (N_2188,N_1524,N_1752);
and U2189 (N_2189,N_1530,N_1850);
nor U2190 (N_2190,N_1737,N_1889);
nand U2191 (N_2191,N_1729,N_1910);
and U2192 (N_2192,N_1528,N_1907);
and U2193 (N_2193,N_1726,N_1669);
and U2194 (N_2194,N_1923,N_1516);
nor U2195 (N_2195,N_1655,N_1647);
or U2196 (N_2196,N_1999,N_1762);
and U2197 (N_2197,N_1597,N_1619);
nand U2198 (N_2198,N_1725,N_1944);
or U2199 (N_2199,N_1813,N_1598);
nor U2200 (N_2200,N_1706,N_1666);
nor U2201 (N_2201,N_1749,N_1585);
nand U2202 (N_2202,N_1708,N_1790);
or U2203 (N_2203,N_1536,N_1662);
and U2204 (N_2204,N_1934,N_1574);
nor U2205 (N_2205,N_1592,N_1566);
and U2206 (N_2206,N_1650,N_1821);
or U2207 (N_2207,N_1718,N_1856);
or U2208 (N_2208,N_1924,N_1879);
nor U2209 (N_2209,N_1909,N_1527);
nor U2210 (N_2210,N_1763,N_1904);
or U2211 (N_2211,N_1930,N_1768);
and U2212 (N_2212,N_1521,N_1554);
or U2213 (N_2213,N_1902,N_1570);
nand U2214 (N_2214,N_1745,N_1517);
nand U2215 (N_2215,N_1657,N_1831);
or U2216 (N_2216,N_1621,N_1917);
nand U2217 (N_2217,N_1573,N_1789);
and U2218 (N_2218,N_1915,N_1802);
nor U2219 (N_2219,N_1837,N_1555);
and U2220 (N_2220,N_1744,N_1916);
or U2221 (N_2221,N_1870,N_1880);
nand U2222 (N_2222,N_1931,N_1547);
xor U2223 (N_2223,N_1937,N_1965);
nor U2224 (N_2224,N_1791,N_1816);
and U2225 (N_2225,N_1976,N_1781);
or U2226 (N_2226,N_1688,N_1691);
nand U2227 (N_2227,N_1906,N_1591);
nor U2228 (N_2228,N_1992,N_1639);
nor U2229 (N_2229,N_1559,N_1719);
nand U2230 (N_2230,N_1804,N_1805);
or U2231 (N_2231,N_1888,N_1875);
or U2232 (N_2232,N_1661,N_1832);
and U2233 (N_2233,N_1862,N_1741);
nor U2234 (N_2234,N_1599,N_1620);
nand U2235 (N_2235,N_1807,N_1780);
and U2236 (N_2236,N_1674,N_1958);
nor U2237 (N_2237,N_1504,N_1567);
and U2238 (N_2238,N_1721,N_1625);
or U2239 (N_2239,N_1963,N_1631);
nor U2240 (N_2240,N_1686,N_1769);
nor U2241 (N_2241,N_1509,N_1644);
nor U2242 (N_2242,N_1648,N_1950);
nor U2243 (N_2243,N_1853,N_1868);
nor U2244 (N_2244,N_1722,N_1953);
nand U2245 (N_2245,N_1919,N_1785);
nand U2246 (N_2246,N_1670,N_1758);
or U2247 (N_2247,N_1838,N_1542);
nand U2248 (N_2248,N_1546,N_1594);
or U2249 (N_2249,N_1847,N_1656);
nor U2250 (N_2250,N_1895,N_1969);
and U2251 (N_2251,N_1679,N_1597);
xor U2252 (N_2252,N_1805,N_1920);
and U2253 (N_2253,N_1560,N_1999);
or U2254 (N_2254,N_1695,N_1891);
or U2255 (N_2255,N_1793,N_1565);
and U2256 (N_2256,N_1788,N_1774);
and U2257 (N_2257,N_1786,N_1766);
nand U2258 (N_2258,N_1948,N_1828);
nand U2259 (N_2259,N_1989,N_1834);
and U2260 (N_2260,N_1737,N_1892);
or U2261 (N_2261,N_1654,N_1874);
or U2262 (N_2262,N_1983,N_1825);
nor U2263 (N_2263,N_1690,N_1644);
or U2264 (N_2264,N_1667,N_1589);
nor U2265 (N_2265,N_1538,N_1743);
or U2266 (N_2266,N_1546,N_1977);
nand U2267 (N_2267,N_1698,N_1773);
nand U2268 (N_2268,N_1716,N_1539);
and U2269 (N_2269,N_1885,N_1936);
nand U2270 (N_2270,N_1851,N_1886);
or U2271 (N_2271,N_1769,N_1665);
nor U2272 (N_2272,N_1614,N_1535);
nor U2273 (N_2273,N_1808,N_1525);
and U2274 (N_2274,N_1885,N_1595);
and U2275 (N_2275,N_1530,N_1675);
nor U2276 (N_2276,N_1849,N_1923);
nand U2277 (N_2277,N_1978,N_1787);
nand U2278 (N_2278,N_1743,N_1777);
nor U2279 (N_2279,N_1624,N_1521);
nand U2280 (N_2280,N_1550,N_1763);
or U2281 (N_2281,N_1761,N_1520);
or U2282 (N_2282,N_1577,N_1620);
or U2283 (N_2283,N_1905,N_1850);
nor U2284 (N_2284,N_1685,N_1747);
nand U2285 (N_2285,N_1699,N_1759);
and U2286 (N_2286,N_1652,N_1982);
nand U2287 (N_2287,N_1537,N_1903);
nand U2288 (N_2288,N_1555,N_1719);
nand U2289 (N_2289,N_1922,N_1963);
nor U2290 (N_2290,N_1750,N_1967);
and U2291 (N_2291,N_1649,N_1861);
xnor U2292 (N_2292,N_1852,N_1648);
nand U2293 (N_2293,N_1588,N_1561);
and U2294 (N_2294,N_1849,N_1540);
or U2295 (N_2295,N_1599,N_1559);
or U2296 (N_2296,N_1776,N_1750);
nor U2297 (N_2297,N_1863,N_1893);
nor U2298 (N_2298,N_1513,N_1877);
and U2299 (N_2299,N_1672,N_1794);
nor U2300 (N_2300,N_1732,N_1560);
nand U2301 (N_2301,N_1806,N_1529);
and U2302 (N_2302,N_1969,N_1598);
nand U2303 (N_2303,N_1559,N_1644);
nor U2304 (N_2304,N_1974,N_1889);
and U2305 (N_2305,N_1920,N_1652);
and U2306 (N_2306,N_1515,N_1706);
nor U2307 (N_2307,N_1921,N_1514);
nand U2308 (N_2308,N_1637,N_1690);
nor U2309 (N_2309,N_1905,N_1514);
nand U2310 (N_2310,N_1670,N_1971);
nand U2311 (N_2311,N_1810,N_1756);
nor U2312 (N_2312,N_1536,N_1845);
and U2313 (N_2313,N_1796,N_1978);
and U2314 (N_2314,N_1979,N_1595);
or U2315 (N_2315,N_1954,N_1782);
or U2316 (N_2316,N_1889,N_1887);
and U2317 (N_2317,N_1792,N_1719);
or U2318 (N_2318,N_1980,N_1639);
or U2319 (N_2319,N_1840,N_1772);
nor U2320 (N_2320,N_1722,N_1931);
nor U2321 (N_2321,N_1791,N_1951);
nand U2322 (N_2322,N_1603,N_1614);
or U2323 (N_2323,N_1957,N_1715);
nor U2324 (N_2324,N_1815,N_1614);
or U2325 (N_2325,N_1841,N_1837);
nor U2326 (N_2326,N_1533,N_1977);
and U2327 (N_2327,N_1962,N_1959);
nand U2328 (N_2328,N_1968,N_1928);
nand U2329 (N_2329,N_1689,N_1577);
nand U2330 (N_2330,N_1501,N_1979);
nor U2331 (N_2331,N_1899,N_1812);
or U2332 (N_2332,N_1767,N_1570);
nand U2333 (N_2333,N_1988,N_1932);
nor U2334 (N_2334,N_1846,N_1741);
nor U2335 (N_2335,N_1679,N_1595);
nor U2336 (N_2336,N_1850,N_1535);
and U2337 (N_2337,N_1532,N_1564);
xor U2338 (N_2338,N_1712,N_1514);
nor U2339 (N_2339,N_1550,N_1847);
nor U2340 (N_2340,N_1572,N_1963);
or U2341 (N_2341,N_1892,N_1945);
or U2342 (N_2342,N_1703,N_1970);
or U2343 (N_2343,N_1965,N_1860);
nand U2344 (N_2344,N_1558,N_1783);
or U2345 (N_2345,N_1710,N_1937);
nor U2346 (N_2346,N_1964,N_1654);
nor U2347 (N_2347,N_1524,N_1610);
xor U2348 (N_2348,N_1529,N_1594);
or U2349 (N_2349,N_1577,N_1666);
or U2350 (N_2350,N_1544,N_1799);
nor U2351 (N_2351,N_1909,N_1815);
nor U2352 (N_2352,N_1582,N_1604);
or U2353 (N_2353,N_1793,N_1656);
or U2354 (N_2354,N_1923,N_1626);
and U2355 (N_2355,N_1585,N_1640);
nor U2356 (N_2356,N_1626,N_1503);
nor U2357 (N_2357,N_1673,N_1993);
or U2358 (N_2358,N_1600,N_1691);
or U2359 (N_2359,N_1976,N_1576);
nand U2360 (N_2360,N_1662,N_1806);
or U2361 (N_2361,N_1656,N_1538);
or U2362 (N_2362,N_1617,N_1954);
or U2363 (N_2363,N_1532,N_1720);
and U2364 (N_2364,N_1833,N_1834);
and U2365 (N_2365,N_1609,N_1636);
nand U2366 (N_2366,N_1812,N_1586);
nand U2367 (N_2367,N_1767,N_1721);
or U2368 (N_2368,N_1959,N_1752);
nor U2369 (N_2369,N_1749,N_1634);
or U2370 (N_2370,N_1866,N_1592);
nand U2371 (N_2371,N_1542,N_1968);
and U2372 (N_2372,N_1643,N_1557);
and U2373 (N_2373,N_1654,N_1928);
nand U2374 (N_2374,N_1514,N_1653);
nor U2375 (N_2375,N_1506,N_1797);
nand U2376 (N_2376,N_1957,N_1633);
and U2377 (N_2377,N_1953,N_1873);
or U2378 (N_2378,N_1773,N_1643);
and U2379 (N_2379,N_1523,N_1596);
and U2380 (N_2380,N_1898,N_1893);
nor U2381 (N_2381,N_1660,N_1523);
xnor U2382 (N_2382,N_1636,N_1850);
nand U2383 (N_2383,N_1880,N_1500);
nor U2384 (N_2384,N_1776,N_1854);
and U2385 (N_2385,N_1784,N_1920);
nand U2386 (N_2386,N_1864,N_1801);
or U2387 (N_2387,N_1647,N_1796);
and U2388 (N_2388,N_1881,N_1726);
nor U2389 (N_2389,N_1803,N_1799);
and U2390 (N_2390,N_1646,N_1941);
or U2391 (N_2391,N_1606,N_1625);
xor U2392 (N_2392,N_1658,N_1616);
or U2393 (N_2393,N_1702,N_1834);
or U2394 (N_2394,N_1602,N_1549);
xor U2395 (N_2395,N_1854,N_1868);
nor U2396 (N_2396,N_1556,N_1744);
or U2397 (N_2397,N_1770,N_1779);
and U2398 (N_2398,N_1797,N_1932);
nor U2399 (N_2399,N_1578,N_1674);
and U2400 (N_2400,N_1587,N_1723);
or U2401 (N_2401,N_1981,N_1755);
or U2402 (N_2402,N_1802,N_1794);
and U2403 (N_2403,N_1536,N_1560);
and U2404 (N_2404,N_1640,N_1907);
nand U2405 (N_2405,N_1592,N_1546);
nor U2406 (N_2406,N_1690,N_1618);
nor U2407 (N_2407,N_1837,N_1709);
nor U2408 (N_2408,N_1729,N_1603);
and U2409 (N_2409,N_1814,N_1768);
and U2410 (N_2410,N_1519,N_1926);
nand U2411 (N_2411,N_1926,N_1916);
or U2412 (N_2412,N_1776,N_1506);
or U2413 (N_2413,N_1661,N_1567);
or U2414 (N_2414,N_1804,N_1795);
nand U2415 (N_2415,N_1547,N_1992);
nand U2416 (N_2416,N_1552,N_1503);
nor U2417 (N_2417,N_1544,N_1701);
nand U2418 (N_2418,N_1935,N_1595);
or U2419 (N_2419,N_1779,N_1650);
and U2420 (N_2420,N_1549,N_1891);
or U2421 (N_2421,N_1681,N_1869);
or U2422 (N_2422,N_1942,N_1990);
nand U2423 (N_2423,N_1899,N_1852);
or U2424 (N_2424,N_1853,N_1967);
nand U2425 (N_2425,N_1584,N_1669);
or U2426 (N_2426,N_1669,N_1870);
and U2427 (N_2427,N_1973,N_1926);
nor U2428 (N_2428,N_1691,N_1668);
nand U2429 (N_2429,N_1884,N_1837);
xor U2430 (N_2430,N_1716,N_1564);
and U2431 (N_2431,N_1959,N_1965);
and U2432 (N_2432,N_1903,N_1774);
and U2433 (N_2433,N_1774,N_1616);
nand U2434 (N_2434,N_1646,N_1731);
nand U2435 (N_2435,N_1687,N_1732);
and U2436 (N_2436,N_1507,N_1509);
and U2437 (N_2437,N_1915,N_1596);
or U2438 (N_2438,N_1545,N_1792);
and U2439 (N_2439,N_1513,N_1856);
or U2440 (N_2440,N_1941,N_1543);
nand U2441 (N_2441,N_1815,N_1703);
nor U2442 (N_2442,N_1526,N_1521);
nor U2443 (N_2443,N_1669,N_1874);
and U2444 (N_2444,N_1611,N_1727);
nand U2445 (N_2445,N_1906,N_1613);
nor U2446 (N_2446,N_1855,N_1998);
and U2447 (N_2447,N_1960,N_1640);
nand U2448 (N_2448,N_1795,N_1808);
nand U2449 (N_2449,N_1941,N_1782);
nand U2450 (N_2450,N_1822,N_1584);
nand U2451 (N_2451,N_1507,N_1830);
and U2452 (N_2452,N_1793,N_1895);
and U2453 (N_2453,N_1500,N_1929);
nand U2454 (N_2454,N_1922,N_1548);
nor U2455 (N_2455,N_1974,N_1635);
nand U2456 (N_2456,N_1952,N_1795);
nor U2457 (N_2457,N_1526,N_1810);
or U2458 (N_2458,N_1570,N_1634);
and U2459 (N_2459,N_1512,N_1861);
nand U2460 (N_2460,N_1871,N_1959);
and U2461 (N_2461,N_1535,N_1731);
nand U2462 (N_2462,N_1731,N_1577);
or U2463 (N_2463,N_1543,N_1626);
nor U2464 (N_2464,N_1687,N_1558);
and U2465 (N_2465,N_1828,N_1748);
nand U2466 (N_2466,N_1960,N_1949);
xnor U2467 (N_2467,N_1816,N_1905);
or U2468 (N_2468,N_1847,N_1994);
and U2469 (N_2469,N_1957,N_1837);
nor U2470 (N_2470,N_1756,N_1666);
and U2471 (N_2471,N_1880,N_1633);
or U2472 (N_2472,N_1823,N_1972);
and U2473 (N_2473,N_1952,N_1671);
nand U2474 (N_2474,N_1844,N_1905);
nand U2475 (N_2475,N_1881,N_1816);
nand U2476 (N_2476,N_1863,N_1787);
and U2477 (N_2477,N_1790,N_1593);
or U2478 (N_2478,N_1564,N_1773);
nand U2479 (N_2479,N_1731,N_1848);
nand U2480 (N_2480,N_1561,N_1644);
nand U2481 (N_2481,N_1867,N_1724);
and U2482 (N_2482,N_1709,N_1581);
or U2483 (N_2483,N_1724,N_1668);
xnor U2484 (N_2484,N_1631,N_1527);
or U2485 (N_2485,N_1869,N_1745);
nand U2486 (N_2486,N_1826,N_1635);
nor U2487 (N_2487,N_1729,N_1829);
nand U2488 (N_2488,N_1920,N_1786);
and U2489 (N_2489,N_1935,N_1597);
nand U2490 (N_2490,N_1612,N_1682);
nand U2491 (N_2491,N_1944,N_1994);
and U2492 (N_2492,N_1961,N_1627);
nor U2493 (N_2493,N_1695,N_1875);
or U2494 (N_2494,N_1980,N_1534);
and U2495 (N_2495,N_1525,N_1745);
nand U2496 (N_2496,N_1760,N_1526);
or U2497 (N_2497,N_1919,N_1690);
nand U2498 (N_2498,N_1672,N_1642);
and U2499 (N_2499,N_1739,N_1737);
nand U2500 (N_2500,N_2247,N_2057);
or U2501 (N_2501,N_2426,N_2234);
and U2502 (N_2502,N_2094,N_2015);
or U2503 (N_2503,N_2091,N_2150);
nor U2504 (N_2504,N_2290,N_2005);
nand U2505 (N_2505,N_2085,N_2284);
nand U2506 (N_2506,N_2497,N_2035);
nand U2507 (N_2507,N_2288,N_2257);
nor U2508 (N_2508,N_2326,N_2049);
and U2509 (N_2509,N_2180,N_2066);
and U2510 (N_2510,N_2296,N_2036);
or U2511 (N_2511,N_2480,N_2068);
nand U2512 (N_2512,N_2424,N_2281);
or U2513 (N_2513,N_2221,N_2215);
and U2514 (N_2514,N_2159,N_2210);
or U2515 (N_2515,N_2414,N_2071);
or U2516 (N_2516,N_2367,N_2208);
nand U2517 (N_2517,N_2047,N_2053);
and U2518 (N_2518,N_2170,N_2302);
or U2519 (N_2519,N_2492,N_2463);
nor U2520 (N_2520,N_2113,N_2146);
nor U2521 (N_2521,N_2255,N_2218);
xor U2522 (N_2522,N_2327,N_2173);
and U2523 (N_2523,N_2483,N_2306);
nor U2524 (N_2524,N_2007,N_2259);
nor U2525 (N_2525,N_2486,N_2298);
nand U2526 (N_2526,N_2462,N_2217);
nor U2527 (N_2527,N_2164,N_2148);
nor U2528 (N_2528,N_2158,N_2044);
nand U2529 (N_2529,N_2446,N_2373);
nor U2530 (N_2530,N_2376,N_2229);
nor U2531 (N_2531,N_2398,N_2470);
and U2532 (N_2532,N_2484,N_2351);
nand U2533 (N_2533,N_2467,N_2419);
and U2534 (N_2534,N_2272,N_2030);
and U2535 (N_2535,N_2372,N_2293);
or U2536 (N_2536,N_2109,N_2136);
or U2537 (N_2537,N_2198,N_2421);
and U2538 (N_2538,N_2065,N_2400);
nand U2539 (N_2539,N_2292,N_2494);
nor U2540 (N_2540,N_2123,N_2453);
and U2541 (N_2541,N_2029,N_2072);
or U2542 (N_2542,N_2097,N_2360);
or U2543 (N_2543,N_2416,N_2037);
or U2544 (N_2544,N_2407,N_2013);
nor U2545 (N_2545,N_2375,N_2267);
and U2546 (N_2546,N_2336,N_2429);
and U2547 (N_2547,N_2063,N_2058);
nor U2548 (N_2548,N_2264,N_2382);
or U2549 (N_2549,N_2498,N_2124);
nor U2550 (N_2550,N_2265,N_2458);
or U2551 (N_2551,N_2112,N_2415);
and U2552 (N_2552,N_2239,N_2411);
or U2553 (N_2553,N_2254,N_2399);
and U2554 (N_2554,N_2041,N_2337);
or U2555 (N_2555,N_2020,N_2342);
or U2556 (N_2556,N_2045,N_2008);
and U2557 (N_2557,N_2280,N_2493);
nor U2558 (N_2558,N_2316,N_2196);
and U2559 (N_2559,N_2006,N_2475);
or U2560 (N_2560,N_2413,N_2385);
nand U2561 (N_2561,N_2182,N_2436);
nand U2562 (N_2562,N_2115,N_2330);
nor U2563 (N_2563,N_2389,N_2219);
and U2564 (N_2564,N_2025,N_2346);
and U2565 (N_2565,N_2171,N_2294);
and U2566 (N_2566,N_2111,N_2250);
nand U2567 (N_2567,N_2197,N_2354);
nand U2568 (N_2568,N_2039,N_2489);
nand U2569 (N_2569,N_2323,N_2224);
nor U2570 (N_2570,N_2417,N_2258);
or U2571 (N_2571,N_2279,N_2391);
or U2572 (N_2572,N_2418,N_2018);
nand U2573 (N_2573,N_2050,N_2321);
nand U2574 (N_2574,N_2477,N_2232);
nand U2575 (N_2575,N_2108,N_2012);
and U2576 (N_2576,N_2178,N_2393);
nand U2577 (N_2577,N_2460,N_2226);
and U2578 (N_2578,N_2153,N_2349);
or U2579 (N_2579,N_2437,N_2185);
nand U2580 (N_2580,N_2093,N_2353);
xnor U2581 (N_2581,N_2128,N_2248);
nor U2582 (N_2582,N_2485,N_2131);
and U2583 (N_2583,N_2089,N_2069);
and U2584 (N_2584,N_2273,N_2021);
and U2585 (N_2585,N_2023,N_2166);
nor U2586 (N_2586,N_2076,N_2121);
xnor U2587 (N_2587,N_2320,N_2114);
nand U2588 (N_2588,N_2103,N_2003);
nor U2589 (N_2589,N_2220,N_2362);
and U2590 (N_2590,N_2433,N_2435);
nor U2591 (N_2591,N_2213,N_2242);
or U2592 (N_2592,N_2117,N_2074);
and U2593 (N_2593,N_2409,N_2397);
nand U2594 (N_2594,N_2380,N_2371);
and U2595 (N_2595,N_2363,N_2423);
nand U2596 (N_2596,N_2252,N_2135);
or U2597 (N_2597,N_2245,N_2238);
nor U2598 (N_2598,N_2461,N_2473);
xor U2599 (N_2599,N_2187,N_2471);
and U2600 (N_2600,N_2268,N_2033);
nor U2601 (N_2601,N_2341,N_2105);
or U2602 (N_2602,N_2042,N_2356);
xor U2603 (N_2603,N_2443,N_2163);
or U2604 (N_2604,N_2143,N_2445);
and U2605 (N_2605,N_2328,N_2133);
nor U2606 (N_2606,N_2455,N_2396);
and U2607 (N_2607,N_2086,N_2343);
nand U2608 (N_2608,N_2274,N_2102);
xor U2609 (N_2609,N_2137,N_2392);
and U2610 (N_2610,N_2191,N_2287);
and U2611 (N_2611,N_2054,N_2243);
or U2612 (N_2612,N_2456,N_2043);
and U2613 (N_2613,N_2237,N_2016);
and U2614 (N_2614,N_2308,N_2231);
and U2615 (N_2615,N_2165,N_2395);
nand U2616 (N_2616,N_2212,N_2203);
nor U2617 (N_2617,N_2099,N_2096);
and U2618 (N_2618,N_2017,N_2228);
or U2619 (N_2619,N_2001,N_2495);
or U2620 (N_2620,N_2200,N_2004);
nor U2621 (N_2621,N_2269,N_2055);
nand U2622 (N_2622,N_2022,N_2240);
and U2623 (N_2623,N_2476,N_2034);
and U2624 (N_2624,N_2390,N_2009);
or U2625 (N_2625,N_2438,N_2449);
nand U2626 (N_2626,N_2087,N_2184);
nor U2627 (N_2627,N_2233,N_2019);
nor U2628 (N_2628,N_2079,N_2011);
nand U2629 (N_2629,N_2078,N_2144);
or U2630 (N_2630,N_2469,N_2075);
or U2631 (N_2631,N_2046,N_2127);
and U2632 (N_2632,N_2277,N_2080);
nand U2633 (N_2633,N_2186,N_2451);
or U2634 (N_2634,N_2325,N_2090);
and U2635 (N_2635,N_2310,N_2285);
and U2636 (N_2636,N_2410,N_2106);
nor U2637 (N_2637,N_2262,N_2324);
xnor U2638 (N_2638,N_2434,N_2309);
and U2639 (N_2639,N_2010,N_2125);
or U2640 (N_2640,N_2002,N_2110);
nand U2641 (N_2641,N_2152,N_2139);
nand U2642 (N_2642,N_2312,N_2408);
nand U2643 (N_2643,N_2179,N_2073);
and U2644 (N_2644,N_2358,N_2251);
or U2645 (N_2645,N_2126,N_2100);
and U2646 (N_2646,N_2420,N_2332);
or U2647 (N_2647,N_2168,N_2369);
and U2648 (N_2648,N_2056,N_2261);
and U2649 (N_2649,N_2194,N_2081);
nand U2650 (N_2650,N_2027,N_2468);
and U2651 (N_2651,N_2295,N_2404);
nand U2652 (N_2652,N_2064,N_2490);
and U2653 (N_2653,N_2300,N_2307);
or U2654 (N_2654,N_2236,N_2028);
nor U2655 (N_2655,N_2402,N_2225);
or U2656 (N_2656,N_2394,N_2347);
or U2657 (N_2657,N_2192,N_2052);
or U2658 (N_2658,N_2183,N_2365);
nor U2659 (N_2659,N_2283,N_2403);
nand U2660 (N_2660,N_2452,N_2361);
nand U2661 (N_2661,N_2157,N_2059);
and U2662 (N_2662,N_2024,N_2088);
nor U2663 (N_2663,N_2289,N_2303);
nand U2664 (N_2664,N_2211,N_2377);
and U2665 (N_2665,N_2286,N_2340);
nor U2666 (N_2666,N_2301,N_2266);
nor U2667 (N_2667,N_2026,N_2032);
or U2668 (N_2668,N_2175,N_2318);
nor U2669 (N_2669,N_2161,N_2061);
nor U2670 (N_2670,N_2313,N_2107);
or U2671 (N_2671,N_2195,N_2174);
or U2672 (N_2672,N_2223,N_2297);
nand U2673 (N_2673,N_2275,N_2122);
or U2674 (N_2674,N_2140,N_2207);
or U2675 (N_2675,N_2199,N_2241);
or U2676 (N_2676,N_2104,N_2422);
nor U2677 (N_2677,N_2487,N_2364);
nand U2678 (N_2678,N_2482,N_2401);
and U2679 (N_2679,N_2335,N_2314);
and U2680 (N_2680,N_2141,N_2383);
nor U2681 (N_2681,N_2244,N_2441);
nand U2682 (N_2682,N_2176,N_2406);
or U2683 (N_2683,N_2132,N_2428);
and U2684 (N_2684,N_2048,N_2142);
or U2685 (N_2685,N_2189,N_2038);
or U2686 (N_2686,N_2387,N_2384);
nor U2687 (N_2687,N_2350,N_2160);
or U2688 (N_2688,N_2379,N_2051);
nand U2689 (N_2689,N_2442,N_2425);
and U2690 (N_2690,N_2319,N_2271);
nor U2691 (N_2691,N_2134,N_2120);
nor U2692 (N_2692,N_2167,N_2444);
and U2693 (N_2693,N_2172,N_2070);
and U2694 (N_2694,N_2188,N_2499);
or U2695 (N_2695,N_2249,N_2431);
or U2696 (N_2696,N_2260,N_2177);
nand U2697 (N_2697,N_2270,N_2317);
xor U2698 (N_2698,N_2077,N_2031);
nand U2699 (N_2699,N_2204,N_2227);
and U2700 (N_2700,N_2465,N_2405);
or U2701 (N_2701,N_2216,N_2155);
nor U2702 (N_2702,N_2092,N_2095);
nand U2703 (N_2703,N_2479,N_2378);
and U2704 (N_2704,N_2206,N_2448);
or U2705 (N_2705,N_2256,N_2491);
and U2706 (N_2706,N_2119,N_2230);
and U2707 (N_2707,N_2374,N_2331);
or U2708 (N_2708,N_2083,N_2334);
or U2709 (N_2709,N_2282,N_2149);
nor U2710 (N_2710,N_2322,N_2381);
nand U2711 (N_2711,N_2368,N_2014);
or U2712 (N_2712,N_2000,N_2062);
nand U2713 (N_2713,N_2412,N_2386);
nand U2714 (N_2714,N_2067,N_2235);
and U2715 (N_2715,N_2344,N_2246);
nor U2716 (N_2716,N_2478,N_2457);
or U2717 (N_2717,N_2357,N_2299);
xor U2718 (N_2718,N_2116,N_2339);
nor U2719 (N_2719,N_2366,N_2447);
and U2720 (N_2720,N_2129,N_2345);
nor U2721 (N_2721,N_2329,N_2388);
nand U2722 (N_2722,N_2201,N_2202);
nand U2723 (N_2723,N_2278,N_2181);
and U2724 (N_2724,N_2145,N_2305);
nor U2725 (N_2725,N_2370,N_2466);
or U2726 (N_2726,N_2439,N_2162);
xnor U2727 (N_2727,N_2459,N_2333);
or U2728 (N_2728,N_2464,N_2084);
and U2729 (N_2729,N_2474,N_2138);
or U2730 (N_2730,N_2130,N_2205);
and U2731 (N_2731,N_2263,N_2082);
nand U2732 (N_2732,N_2315,N_2151);
and U2733 (N_2733,N_2118,N_2481);
and U2734 (N_2734,N_2156,N_2454);
or U2735 (N_2735,N_2432,N_2472);
or U2736 (N_2736,N_2304,N_2311);
xor U2737 (N_2737,N_2276,N_2190);
or U2738 (N_2738,N_2214,N_2169);
nor U2739 (N_2739,N_2427,N_2488);
nor U2740 (N_2740,N_2222,N_2450);
or U2741 (N_2741,N_2101,N_2209);
xor U2742 (N_2742,N_2060,N_2430);
nand U2743 (N_2743,N_2098,N_2440);
and U2744 (N_2744,N_2040,N_2154);
or U2745 (N_2745,N_2291,N_2359);
and U2746 (N_2746,N_2348,N_2496);
or U2747 (N_2747,N_2338,N_2253);
and U2748 (N_2748,N_2193,N_2147);
nand U2749 (N_2749,N_2355,N_2352);
nand U2750 (N_2750,N_2018,N_2229);
xor U2751 (N_2751,N_2118,N_2491);
nand U2752 (N_2752,N_2162,N_2469);
or U2753 (N_2753,N_2064,N_2311);
nor U2754 (N_2754,N_2021,N_2177);
nor U2755 (N_2755,N_2186,N_2460);
nand U2756 (N_2756,N_2444,N_2300);
or U2757 (N_2757,N_2173,N_2435);
xor U2758 (N_2758,N_2287,N_2248);
or U2759 (N_2759,N_2420,N_2313);
and U2760 (N_2760,N_2386,N_2498);
or U2761 (N_2761,N_2114,N_2112);
nand U2762 (N_2762,N_2313,N_2308);
nand U2763 (N_2763,N_2048,N_2024);
and U2764 (N_2764,N_2082,N_2315);
and U2765 (N_2765,N_2181,N_2117);
nand U2766 (N_2766,N_2296,N_2194);
or U2767 (N_2767,N_2204,N_2141);
nand U2768 (N_2768,N_2068,N_2106);
or U2769 (N_2769,N_2424,N_2035);
or U2770 (N_2770,N_2391,N_2341);
nand U2771 (N_2771,N_2024,N_2239);
xnor U2772 (N_2772,N_2333,N_2190);
and U2773 (N_2773,N_2232,N_2145);
nand U2774 (N_2774,N_2159,N_2205);
and U2775 (N_2775,N_2389,N_2409);
nand U2776 (N_2776,N_2075,N_2123);
or U2777 (N_2777,N_2091,N_2131);
nor U2778 (N_2778,N_2012,N_2424);
and U2779 (N_2779,N_2154,N_2213);
and U2780 (N_2780,N_2340,N_2396);
and U2781 (N_2781,N_2417,N_2493);
xor U2782 (N_2782,N_2410,N_2370);
nor U2783 (N_2783,N_2172,N_2184);
nor U2784 (N_2784,N_2313,N_2239);
nand U2785 (N_2785,N_2423,N_2186);
and U2786 (N_2786,N_2258,N_2486);
nor U2787 (N_2787,N_2415,N_2094);
and U2788 (N_2788,N_2401,N_2477);
and U2789 (N_2789,N_2231,N_2123);
and U2790 (N_2790,N_2039,N_2373);
nand U2791 (N_2791,N_2404,N_2494);
and U2792 (N_2792,N_2376,N_2001);
nor U2793 (N_2793,N_2008,N_2339);
nor U2794 (N_2794,N_2272,N_2380);
or U2795 (N_2795,N_2056,N_2355);
nand U2796 (N_2796,N_2404,N_2210);
and U2797 (N_2797,N_2172,N_2099);
and U2798 (N_2798,N_2267,N_2056);
nor U2799 (N_2799,N_2097,N_2042);
and U2800 (N_2800,N_2071,N_2053);
nor U2801 (N_2801,N_2040,N_2384);
and U2802 (N_2802,N_2150,N_2251);
nand U2803 (N_2803,N_2376,N_2490);
nand U2804 (N_2804,N_2218,N_2248);
and U2805 (N_2805,N_2064,N_2076);
or U2806 (N_2806,N_2076,N_2062);
or U2807 (N_2807,N_2078,N_2071);
xor U2808 (N_2808,N_2011,N_2033);
and U2809 (N_2809,N_2149,N_2057);
nor U2810 (N_2810,N_2110,N_2324);
nand U2811 (N_2811,N_2007,N_2002);
or U2812 (N_2812,N_2405,N_2081);
nand U2813 (N_2813,N_2451,N_2355);
nand U2814 (N_2814,N_2425,N_2458);
and U2815 (N_2815,N_2050,N_2293);
nor U2816 (N_2816,N_2257,N_2178);
nor U2817 (N_2817,N_2364,N_2290);
nand U2818 (N_2818,N_2338,N_2487);
nor U2819 (N_2819,N_2453,N_2167);
and U2820 (N_2820,N_2100,N_2024);
xnor U2821 (N_2821,N_2063,N_2423);
nor U2822 (N_2822,N_2228,N_2350);
nand U2823 (N_2823,N_2068,N_2035);
and U2824 (N_2824,N_2157,N_2291);
and U2825 (N_2825,N_2470,N_2164);
nor U2826 (N_2826,N_2191,N_2116);
nor U2827 (N_2827,N_2327,N_2428);
nor U2828 (N_2828,N_2075,N_2408);
nand U2829 (N_2829,N_2037,N_2153);
and U2830 (N_2830,N_2217,N_2417);
and U2831 (N_2831,N_2406,N_2327);
or U2832 (N_2832,N_2467,N_2240);
and U2833 (N_2833,N_2089,N_2075);
nor U2834 (N_2834,N_2064,N_2332);
nor U2835 (N_2835,N_2254,N_2303);
nor U2836 (N_2836,N_2272,N_2295);
and U2837 (N_2837,N_2029,N_2479);
and U2838 (N_2838,N_2224,N_2428);
nand U2839 (N_2839,N_2077,N_2356);
nand U2840 (N_2840,N_2343,N_2406);
and U2841 (N_2841,N_2195,N_2438);
or U2842 (N_2842,N_2171,N_2113);
nor U2843 (N_2843,N_2299,N_2173);
nor U2844 (N_2844,N_2105,N_2403);
nor U2845 (N_2845,N_2056,N_2348);
nand U2846 (N_2846,N_2104,N_2047);
or U2847 (N_2847,N_2153,N_2163);
or U2848 (N_2848,N_2385,N_2466);
nor U2849 (N_2849,N_2244,N_2382);
or U2850 (N_2850,N_2261,N_2297);
and U2851 (N_2851,N_2446,N_2480);
nor U2852 (N_2852,N_2233,N_2370);
or U2853 (N_2853,N_2222,N_2239);
or U2854 (N_2854,N_2293,N_2180);
nor U2855 (N_2855,N_2406,N_2171);
nor U2856 (N_2856,N_2429,N_2044);
nor U2857 (N_2857,N_2238,N_2452);
or U2858 (N_2858,N_2080,N_2102);
nand U2859 (N_2859,N_2026,N_2147);
nand U2860 (N_2860,N_2117,N_2007);
xnor U2861 (N_2861,N_2230,N_2437);
nor U2862 (N_2862,N_2250,N_2333);
nand U2863 (N_2863,N_2398,N_2097);
nor U2864 (N_2864,N_2408,N_2486);
xor U2865 (N_2865,N_2486,N_2242);
nor U2866 (N_2866,N_2072,N_2438);
nor U2867 (N_2867,N_2101,N_2055);
or U2868 (N_2868,N_2292,N_2228);
and U2869 (N_2869,N_2266,N_2265);
nor U2870 (N_2870,N_2065,N_2090);
xnor U2871 (N_2871,N_2196,N_2338);
and U2872 (N_2872,N_2306,N_2393);
nor U2873 (N_2873,N_2167,N_2390);
or U2874 (N_2874,N_2065,N_2182);
or U2875 (N_2875,N_2043,N_2002);
and U2876 (N_2876,N_2490,N_2346);
and U2877 (N_2877,N_2185,N_2007);
and U2878 (N_2878,N_2196,N_2434);
nand U2879 (N_2879,N_2016,N_2195);
and U2880 (N_2880,N_2078,N_2072);
xnor U2881 (N_2881,N_2418,N_2118);
nand U2882 (N_2882,N_2240,N_2153);
and U2883 (N_2883,N_2325,N_2066);
and U2884 (N_2884,N_2145,N_2447);
or U2885 (N_2885,N_2413,N_2400);
xor U2886 (N_2886,N_2154,N_2237);
and U2887 (N_2887,N_2241,N_2109);
or U2888 (N_2888,N_2389,N_2447);
or U2889 (N_2889,N_2094,N_2209);
nor U2890 (N_2890,N_2459,N_2153);
and U2891 (N_2891,N_2498,N_2038);
or U2892 (N_2892,N_2446,N_2476);
nor U2893 (N_2893,N_2423,N_2079);
nor U2894 (N_2894,N_2098,N_2197);
xnor U2895 (N_2895,N_2100,N_2253);
and U2896 (N_2896,N_2216,N_2339);
and U2897 (N_2897,N_2044,N_2108);
nor U2898 (N_2898,N_2060,N_2302);
nand U2899 (N_2899,N_2444,N_2313);
and U2900 (N_2900,N_2013,N_2231);
nor U2901 (N_2901,N_2218,N_2179);
and U2902 (N_2902,N_2037,N_2455);
xnor U2903 (N_2903,N_2317,N_2264);
or U2904 (N_2904,N_2164,N_2250);
and U2905 (N_2905,N_2383,N_2342);
or U2906 (N_2906,N_2432,N_2254);
or U2907 (N_2907,N_2493,N_2440);
or U2908 (N_2908,N_2456,N_2470);
nand U2909 (N_2909,N_2217,N_2327);
nand U2910 (N_2910,N_2374,N_2029);
nor U2911 (N_2911,N_2025,N_2162);
nand U2912 (N_2912,N_2186,N_2224);
nand U2913 (N_2913,N_2207,N_2240);
nor U2914 (N_2914,N_2146,N_2192);
nor U2915 (N_2915,N_2457,N_2001);
and U2916 (N_2916,N_2095,N_2184);
and U2917 (N_2917,N_2492,N_2310);
nand U2918 (N_2918,N_2499,N_2266);
nor U2919 (N_2919,N_2236,N_2425);
nand U2920 (N_2920,N_2284,N_2228);
nor U2921 (N_2921,N_2262,N_2194);
nor U2922 (N_2922,N_2070,N_2093);
nand U2923 (N_2923,N_2233,N_2148);
and U2924 (N_2924,N_2370,N_2465);
nor U2925 (N_2925,N_2273,N_2318);
nor U2926 (N_2926,N_2383,N_2072);
or U2927 (N_2927,N_2131,N_2472);
nand U2928 (N_2928,N_2428,N_2048);
nand U2929 (N_2929,N_2482,N_2070);
or U2930 (N_2930,N_2152,N_2213);
xnor U2931 (N_2931,N_2318,N_2081);
nor U2932 (N_2932,N_2389,N_2037);
and U2933 (N_2933,N_2463,N_2060);
and U2934 (N_2934,N_2349,N_2249);
and U2935 (N_2935,N_2259,N_2299);
nand U2936 (N_2936,N_2429,N_2034);
nand U2937 (N_2937,N_2192,N_2306);
nor U2938 (N_2938,N_2497,N_2065);
nand U2939 (N_2939,N_2244,N_2197);
nor U2940 (N_2940,N_2117,N_2318);
and U2941 (N_2941,N_2322,N_2202);
nor U2942 (N_2942,N_2414,N_2423);
nor U2943 (N_2943,N_2111,N_2311);
and U2944 (N_2944,N_2194,N_2138);
or U2945 (N_2945,N_2323,N_2459);
or U2946 (N_2946,N_2055,N_2459);
or U2947 (N_2947,N_2124,N_2368);
nor U2948 (N_2948,N_2139,N_2116);
or U2949 (N_2949,N_2158,N_2480);
and U2950 (N_2950,N_2474,N_2270);
and U2951 (N_2951,N_2035,N_2488);
nand U2952 (N_2952,N_2492,N_2117);
nand U2953 (N_2953,N_2348,N_2288);
and U2954 (N_2954,N_2177,N_2093);
and U2955 (N_2955,N_2348,N_2430);
nand U2956 (N_2956,N_2343,N_2233);
or U2957 (N_2957,N_2392,N_2189);
nor U2958 (N_2958,N_2094,N_2202);
and U2959 (N_2959,N_2460,N_2224);
nor U2960 (N_2960,N_2488,N_2274);
and U2961 (N_2961,N_2020,N_2165);
nand U2962 (N_2962,N_2465,N_2236);
nand U2963 (N_2963,N_2126,N_2207);
nor U2964 (N_2964,N_2487,N_2348);
and U2965 (N_2965,N_2472,N_2231);
or U2966 (N_2966,N_2365,N_2117);
and U2967 (N_2967,N_2103,N_2281);
xor U2968 (N_2968,N_2347,N_2085);
or U2969 (N_2969,N_2027,N_2383);
or U2970 (N_2970,N_2144,N_2377);
and U2971 (N_2971,N_2095,N_2015);
nand U2972 (N_2972,N_2459,N_2322);
or U2973 (N_2973,N_2081,N_2267);
and U2974 (N_2974,N_2344,N_2038);
or U2975 (N_2975,N_2082,N_2060);
and U2976 (N_2976,N_2025,N_2418);
nor U2977 (N_2977,N_2339,N_2174);
and U2978 (N_2978,N_2154,N_2098);
nor U2979 (N_2979,N_2255,N_2499);
nor U2980 (N_2980,N_2455,N_2331);
or U2981 (N_2981,N_2220,N_2466);
nor U2982 (N_2982,N_2203,N_2330);
or U2983 (N_2983,N_2288,N_2020);
or U2984 (N_2984,N_2302,N_2327);
and U2985 (N_2985,N_2333,N_2243);
or U2986 (N_2986,N_2235,N_2377);
and U2987 (N_2987,N_2283,N_2454);
or U2988 (N_2988,N_2397,N_2065);
nor U2989 (N_2989,N_2328,N_2058);
nor U2990 (N_2990,N_2278,N_2277);
nor U2991 (N_2991,N_2339,N_2132);
or U2992 (N_2992,N_2014,N_2186);
nand U2993 (N_2993,N_2155,N_2091);
nand U2994 (N_2994,N_2384,N_2405);
nor U2995 (N_2995,N_2034,N_2045);
nand U2996 (N_2996,N_2104,N_2405);
or U2997 (N_2997,N_2134,N_2207);
nor U2998 (N_2998,N_2278,N_2132);
and U2999 (N_2999,N_2114,N_2405);
nor U3000 (N_3000,N_2673,N_2827);
and U3001 (N_3001,N_2637,N_2764);
nor U3002 (N_3002,N_2661,N_2842);
nand U3003 (N_3003,N_2856,N_2976);
or U3004 (N_3004,N_2912,N_2687);
or U3005 (N_3005,N_2895,N_2735);
and U3006 (N_3006,N_2678,N_2745);
nand U3007 (N_3007,N_2890,N_2664);
or U3008 (N_3008,N_2520,N_2791);
nor U3009 (N_3009,N_2925,N_2830);
nand U3010 (N_3010,N_2961,N_2505);
nand U3011 (N_3011,N_2816,N_2647);
nand U3012 (N_3012,N_2972,N_2589);
nand U3013 (N_3013,N_2758,N_2694);
or U3014 (N_3014,N_2815,N_2723);
and U3015 (N_3015,N_2851,N_2573);
nand U3016 (N_3016,N_2992,N_2556);
or U3017 (N_3017,N_2787,N_2886);
and U3018 (N_3018,N_2594,N_2737);
and U3019 (N_3019,N_2662,N_2833);
nor U3020 (N_3020,N_2575,N_2826);
nand U3021 (N_3021,N_2755,N_2742);
and U3022 (N_3022,N_2808,N_2654);
and U3023 (N_3023,N_2528,N_2638);
nor U3024 (N_3024,N_2635,N_2521);
xor U3025 (N_3025,N_2538,N_2853);
and U3026 (N_3026,N_2574,N_2820);
nor U3027 (N_3027,N_2885,N_2844);
or U3028 (N_3028,N_2968,N_2536);
or U3029 (N_3029,N_2843,N_2867);
and U3030 (N_3030,N_2922,N_2719);
and U3031 (N_3031,N_2718,N_2571);
nand U3032 (N_3032,N_2683,N_2974);
nor U3033 (N_3033,N_2532,N_2730);
nor U3034 (N_3034,N_2558,N_2898);
nand U3035 (N_3035,N_2552,N_2775);
and U3036 (N_3036,N_2956,N_2850);
and U3037 (N_3037,N_2762,N_2915);
xor U3038 (N_3038,N_2653,N_2734);
and U3039 (N_3039,N_2636,N_2513);
nor U3040 (N_3040,N_2917,N_2965);
nand U3041 (N_3041,N_2811,N_2875);
xnor U3042 (N_3042,N_2582,N_2697);
nor U3043 (N_3043,N_2523,N_2907);
and U3044 (N_3044,N_2616,N_2861);
or U3045 (N_3045,N_2768,N_2911);
nor U3046 (N_3046,N_2519,N_2620);
nor U3047 (N_3047,N_2892,N_2685);
or U3048 (N_3048,N_2793,N_2502);
nand U3049 (N_3049,N_2522,N_2702);
xor U3050 (N_3050,N_2899,N_2964);
or U3051 (N_3051,N_2786,N_2810);
and U3052 (N_3052,N_2684,N_2946);
or U3053 (N_3053,N_2645,N_2507);
and U3054 (N_3054,N_2710,N_2708);
or U3055 (N_3055,N_2557,N_2749);
or U3056 (N_3056,N_2887,N_2691);
nand U3057 (N_3057,N_2568,N_2999);
and U3058 (N_3058,N_2948,N_2772);
or U3059 (N_3059,N_2966,N_2872);
nor U3060 (N_3060,N_2865,N_2659);
nand U3061 (N_3061,N_2585,N_2931);
and U3062 (N_3062,N_2801,N_2997);
or U3063 (N_3063,N_2590,N_2562);
nor U3064 (N_3064,N_2705,N_2839);
nand U3065 (N_3065,N_2790,N_2676);
and U3066 (N_3066,N_2696,N_2858);
and U3067 (N_3067,N_2903,N_2543);
nor U3068 (N_3068,N_2733,N_2615);
and U3069 (N_3069,N_2567,N_2945);
and U3070 (N_3070,N_2717,N_2955);
nor U3071 (N_3071,N_2648,N_2747);
nor U3072 (N_3072,N_2546,N_2909);
or U3073 (N_3073,N_2792,N_2751);
and U3074 (N_3074,N_2501,N_2977);
or U3075 (N_3075,N_2566,N_2927);
or U3076 (N_3076,N_2725,N_2930);
nor U3077 (N_3077,N_2517,N_2681);
nor U3078 (N_3078,N_2619,N_2918);
nor U3079 (N_3079,N_2914,N_2668);
and U3080 (N_3080,N_2770,N_2729);
and U3081 (N_3081,N_2525,N_2537);
nand U3082 (N_3082,N_2560,N_2539);
nor U3083 (N_3083,N_2510,N_2672);
nand U3084 (N_3084,N_2554,N_2923);
and U3085 (N_3085,N_2941,N_2877);
or U3086 (N_3086,N_2712,N_2595);
nor U3087 (N_3087,N_2626,N_2933);
nor U3088 (N_3088,N_2863,N_2613);
or U3089 (N_3089,N_2722,N_2879);
and U3090 (N_3090,N_2800,N_2766);
and U3091 (N_3091,N_2689,N_2643);
nor U3092 (N_3092,N_2876,N_2852);
nor U3093 (N_3093,N_2860,N_2646);
or U3094 (N_3094,N_2604,N_2511);
or U3095 (N_3095,N_2658,N_2698);
or U3096 (N_3096,N_2541,N_2782);
or U3097 (N_3097,N_2623,N_2514);
or U3098 (N_3098,N_2627,N_2802);
and U3099 (N_3099,N_2576,N_2906);
and U3100 (N_3100,N_2910,N_2748);
and U3101 (N_3101,N_2551,N_2893);
nor U3102 (N_3102,N_2971,N_2845);
nand U3103 (N_3103,N_2550,N_2908);
nand U3104 (N_3104,N_2726,N_2670);
nand U3105 (N_3105,N_2859,N_2652);
or U3106 (N_3106,N_2980,N_2944);
nand U3107 (N_3107,N_2690,N_2570);
and U3108 (N_3108,N_2937,N_2709);
nor U3109 (N_3109,N_2655,N_2625);
or U3110 (N_3110,N_2967,N_2740);
or U3111 (N_3111,N_2544,N_2897);
or U3112 (N_3112,N_2817,N_2932);
and U3113 (N_3113,N_2862,N_2555);
nand U3114 (N_3114,N_2883,N_2973);
or U3115 (N_3115,N_2515,N_2996);
nor U3116 (N_3116,N_2916,N_2644);
or U3117 (N_3117,N_2744,N_2991);
and U3118 (N_3118,N_2987,N_2783);
or U3119 (N_3119,N_2854,N_2963);
nand U3120 (N_3120,N_2754,N_2591);
and U3121 (N_3121,N_2531,N_2796);
nor U3122 (N_3122,N_2848,N_2641);
and U3123 (N_3123,N_2617,N_2821);
nand U3124 (N_3124,N_2612,N_2732);
or U3125 (N_3125,N_2957,N_2855);
or U3126 (N_3126,N_2773,N_2518);
or U3127 (N_3127,N_2985,N_2524);
or U3128 (N_3128,N_2958,N_2632);
xor U3129 (N_3129,N_2765,N_2981);
nor U3130 (N_3130,N_2936,N_2679);
xor U3131 (N_3131,N_2831,N_2716);
or U3132 (N_3132,N_2504,N_2778);
and U3133 (N_3133,N_2559,N_2888);
nor U3134 (N_3134,N_2516,N_2864);
nor U3135 (N_3135,N_2509,N_2953);
or U3136 (N_3136,N_2547,N_2540);
and U3137 (N_3137,N_2869,N_2603);
nand U3138 (N_3138,N_2902,N_2707);
and U3139 (N_3139,N_2846,N_2878);
nand U3140 (N_3140,N_2789,N_2759);
or U3141 (N_3141,N_2753,N_2938);
or U3142 (N_3142,N_2610,N_2534);
or U3143 (N_3143,N_2774,N_2621);
nand U3144 (N_3144,N_2714,N_2896);
xor U3145 (N_3145,N_2785,N_2609);
nand U3146 (N_3146,N_2564,N_2695);
nor U3147 (N_3147,N_2978,N_2935);
xor U3148 (N_3148,N_2784,N_2738);
or U3149 (N_3149,N_2840,N_2951);
nand U3150 (N_3150,N_2703,N_2553);
nand U3151 (N_3151,N_2812,N_2822);
nand U3152 (N_3152,N_2950,N_2736);
nor U3153 (N_3153,N_2666,N_2970);
and U3154 (N_3154,N_2624,N_2807);
nand U3155 (N_3155,N_2577,N_2934);
or U3156 (N_3156,N_2767,N_2752);
and U3157 (N_3157,N_2629,N_2686);
or U3158 (N_3158,N_2640,N_2769);
and U3159 (N_3159,N_2593,N_2866);
and U3160 (N_3160,N_2823,N_2706);
nand U3161 (N_3161,N_2874,N_2870);
or U3162 (N_3162,N_2871,N_2746);
and U3163 (N_3163,N_2873,N_2512);
nor U3164 (N_3164,N_2693,N_2959);
or U3165 (N_3165,N_2928,N_2545);
nor U3166 (N_3166,N_2803,N_2835);
and U3167 (N_3167,N_2634,N_2587);
nor U3168 (N_3168,N_2924,N_2583);
nor U3169 (N_3169,N_2838,N_2663);
nand U3170 (N_3170,N_2776,N_2715);
or U3171 (N_3171,N_2671,N_2614);
or U3172 (N_3172,N_2799,N_2565);
or U3173 (N_3173,N_2984,N_2704);
or U3174 (N_3174,N_2677,N_2527);
xor U3175 (N_3175,N_2795,N_2969);
xnor U3176 (N_3176,N_2542,N_2628);
nand U3177 (N_3177,N_2600,N_2599);
or U3178 (N_3178,N_2572,N_2584);
nor U3179 (N_3179,N_2529,N_2757);
nand U3180 (N_3180,N_2761,N_2642);
nand U3181 (N_3181,N_2756,N_2829);
or U3182 (N_3182,N_2805,N_2889);
nand U3183 (N_3183,N_2926,N_2580);
or U3184 (N_3184,N_2739,N_2727);
nand U3185 (N_3185,N_2804,N_2994);
nor U3186 (N_3186,N_2506,N_2500);
xnor U3187 (N_3187,N_2763,N_2880);
or U3188 (N_3188,N_2962,N_2633);
or U3189 (N_3189,N_2868,N_2650);
and U3190 (N_3190,N_2998,N_2503);
and U3191 (N_3191,N_2891,N_2901);
xor U3192 (N_3192,N_2597,N_2586);
or U3193 (N_3193,N_2780,N_2699);
nand U3194 (N_3194,N_2779,N_2882);
nor U3195 (N_3195,N_2549,N_2667);
or U3196 (N_3196,N_2884,N_2724);
or U3197 (N_3197,N_2605,N_2982);
nor U3198 (N_3198,N_2601,N_2988);
nor U3199 (N_3199,N_2608,N_2949);
nand U3200 (N_3200,N_2760,N_2788);
and U3201 (N_3201,N_2692,N_2657);
nor U3202 (N_3202,N_2824,N_2849);
nor U3203 (N_3203,N_2943,N_2607);
nor U3204 (N_3204,N_2618,N_2904);
nor U3205 (N_3205,N_2993,N_2797);
nand U3206 (N_3206,N_2952,N_2665);
nor U3207 (N_3207,N_2596,N_2622);
and U3208 (N_3208,N_2526,N_2819);
xor U3209 (N_3209,N_2905,N_2913);
xor U3210 (N_3210,N_2535,N_2781);
and U3211 (N_3211,N_2929,N_2674);
nand U3212 (N_3212,N_2611,N_2809);
nor U3213 (N_3213,N_2832,N_2741);
and U3214 (N_3214,N_2979,N_2688);
nand U3215 (N_3215,N_2794,N_2900);
nor U3216 (N_3216,N_2682,N_2533);
or U3217 (N_3217,N_2806,N_2940);
and U3218 (N_3218,N_2881,N_2639);
or U3219 (N_3219,N_2798,N_2530);
or U3220 (N_3220,N_2649,N_2508);
or U3221 (N_3221,N_2602,N_2569);
and U3222 (N_3222,N_2836,N_2983);
and U3223 (N_3223,N_2701,N_2651);
and U3224 (N_3224,N_2548,N_2975);
or U3225 (N_3225,N_2921,N_2606);
nand U3226 (N_3226,N_2954,N_2731);
or U3227 (N_3227,N_2563,N_2680);
nor U3228 (N_3228,N_2894,N_2743);
nand U3229 (N_3229,N_2592,N_2598);
or U3230 (N_3230,N_2828,N_2675);
and U3231 (N_3231,N_2818,N_2777);
nor U3232 (N_3232,N_2920,N_2995);
nor U3233 (N_3233,N_2630,N_2579);
nor U3234 (N_3234,N_2561,N_2578);
or U3235 (N_3235,N_2631,N_2947);
or U3236 (N_3236,N_2660,N_2942);
and U3237 (N_3237,N_2721,N_2939);
nand U3238 (N_3238,N_2713,N_2814);
nor U3239 (N_3239,N_2986,N_2750);
nand U3240 (N_3240,N_2588,N_2834);
and U3241 (N_3241,N_2825,N_2847);
and U3242 (N_3242,N_2919,N_2837);
or U3243 (N_3243,N_2700,N_2728);
nand U3244 (N_3244,N_2711,N_2813);
nand U3245 (N_3245,N_2841,N_2720);
and U3246 (N_3246,N_2989,N_2960);
nand U3247 (N_3247,N_2581,N_2990);
or U3248 (N_3248,N_2669,N_2771);
nand U3249 (N_3249,N_2656,N_2857);
or U3250 (N_3250,N_2973,N_2674);
xnor U3251 (N_3251,N_2715,N_2692);
or U3252 (N_3252,N_2850,N_2695);
nor U3253 (N_3253,N_2639,N_2810);
nand U3254 (N_3254,N_2847,N_2741);
and U3255 (N_3255,N_2861,N_2794);
xor U3256 (N_3256,N_2804,N_2581);
nor U3257 (N_3257,N_2998,N_2965);
or U3258 (N_3258,N_2842,N_2973);
nand U3259 (N_3259,N_2645,N_2924);
nand U3260 (N_3260,N_2981,N_2812);
and U3261 (N_3261,N_2845,N_2777);
nand U3262 (N_3262,N_2717,N_2545);
and U3263 (N_3263,N_2535,N_2600);
or U3264 (N_3264,N_2593,N_2863);
or U3265 (N_3265,N_2507,N_2860);
nand U3266 (N_3266,N_2759,N_2773);
xor U3267 (N_3267,N_2990,N_2991);
nor U3268 (N_3268,N_2741,N_2785);
nand U3269 (N_3269,N_2608,N_2571);
and U3270 (N_3270,N_2579,N_2760);
or U3271 (N_3271,N_2563,N_2654);
nor U3272 (N_3272,N_2912,N_2672);
and U3273 (N_3273,N_2670,N_2573);
and U3274 (N_3274,N_2771,N_2549);
nand U3275 (N_3275,N_2934,N_2889);
nand U3276 (N_3276,N_2629,N_2657);
xor U3277 (N_3277,N_2690,N_2703);
nand U3278 (N_3278,N_2652,N_2811);
nor U3279 (N_3279,N_2622,N_2885);
nand U3280 (N_3280,N_2800,N_2816);
nand U3281 (N_3281,N_2650,N_2822);
nor U3282 (N_3282,N_2850,N_2845);
nand U3283 (N_3283,N_2660,N_2984);
nor U3284 (N_3284,N_2778,N_2937);
nor U3285 (N_3285,N_2572,N_2992);
and U3286 (N_3286,N_2503,N_2816);
nand U3287 (N_3287,N_2694,N_2848);
and U3288 (N_3288,N_2520,N_2962);
or U3289 (N_3289,N_2583,N_2624);
nand U3290 (N_3290,N_2934,N_2875);
and U3291 (N_3291,N_2625,N_2721);
or U3292 (N_3292,N_2782,N_2844);
and U3293 (N_3293,N_2709,N_2964);
or U3294 (N_3294,N_2748,N_2554);
nand U3295 (N_3295,N_2755,N_2526);
and U3296 (N_3296,N_2564,N_2797);
nor U3297 (N_3297,N_2508,N_2877);
nand U3298 (N_3298,N_2572,N_2823);
nor U3299 (N_3299,N_2640,N_2688);
and U3300 (N_3300,N_2550,N_2847);
nor U3301 (N_3301,N_2969,N_2860);
nand U3302 (N_3302,N_2942,N_2766);
and U3303 (N_3303,N_2844,N_2831);
and U3304 (N_3304,N_2981,N_2656);
or U3305 (N_3305,N_2521,N_2621);
and U3306 (N_3306,N_2885,N_2809);
nand U3307 (N_3307,N_2646,N_2761);
nand U3308 (N_3308,N_2868,N_2823);
nand U3309 (N_3309,N_2812,N_2577);
nand U3310 (N_3310,N_2678,N_2860);
or U3311 (N_3311,N_2991,N_2596);
or U3312 (N_3312,N_2774,N_2877);
nor U3313 (N_3313,N_2670,N_2885);
and U3314 (N_3314,N_2761,N_2868);
nor U3315 (N_3315,N_2645,N_2516);
or U3316 (N_3316,N_2575,N_2521);
nor U3317 (N_3317,N_2539,N_2655);
nor U3318 (N_3318,N_2565,N_2643);
or U3319 (N_3319,N_2704,N_2647);
and U3320 (N_3320,N_2798,N_2731);
nor U3321 (N_3321,N_2758,N_2891);
or U3322 (N_3322,N_2854,N_2522);
and U3323 (N_3323,N_2678,N_2912);
and U3324 (N_3324,N_2564,N_2756);
and U3325 (N_3325,N_2721,N_2903);
nand U3326 (N_3326,N_2671,N_2965);
and U3327 (N_3327,N_2636,N_2806);
and U3328 (N_3328,N_2886,N_2965);
nor U3329 (N_3329,N_2871,N_2901);
or U3330 (N_3330,N_2789,N_2609);
nor U3331 (N_3331,N_2642,N_2861);
or U3332 (N_3332,N_2814,N_2926);
nor U3333 (N_3333,N_2508,N_2911);
and U3334 (N_3334,N_2908,N_2846);
nand U3335 (N_3335,N_2572,N_2510);
nor U3336 (N_3336,N_2977,N_2773);
and U3337 (N_3337,N_2773,N_2569);
or U3338 (N_3338,N_2894,N_2593);
nand U3339 (N_3339,N_2803,N_2772);
and U3340 (N_3340,N_2905,N_2934);
or U3341 (N_3341,N_2676,N_2763);
nand U3342 (N_3342,N_2919,N_2956);
nor U3343 (N_3343,N_2782,N_2596);
or U3344 (N_3344,N_2510,N_2690);
or U3345 (N_3345,N_2939,N_2515);
and U3346 (N_3346,N_2700,N_2736);
nand U3347 (N_3347,N_2519,N_2955);
or U3348 (N_3348,N_2716,N_2747);
and U3349 (N_3349,N_2999,N_2932);
nor U3350 (N_3350,N_2641,N_2946);
nand U3351 (N_3351,N_2696,N_2567);
nor U3352 (N_3352,N_2820,N_2698);
and U3353 (N_3353,N_2500,N_2654);
and U3354 (N_3354,N_2662,N_2522);
nor U3355 (N_3355,N_2503,N_2806);
nor U3356 (N_3356,N_2850,N_2551);
nand U3357 (N_3357,N_2697,N_2758);
and U3358 (N_3358,N_2783,N_2805);
or U3359 (N_3359,N_2601,N_2932);
nor U3360 (N_3360,N_2545,N_2812);
nand U3361 (N_3361,N_2668,N_2883);
or U3362 (N_3362,N_2640,N_2503);
nor U3363 (N_3363,N_2570,N_2860);
nand U3364 (N_3364,N_2794,N_2739);
nand U3365 (N_3365,N_2599,N_2619);
nand U3366 (N_3366,N_2799,N_2635);
and U3367 (N_3367,N_2913,N_2567);
and U3368 (N_3368,N_2754,N_2973);
xor U3369 (N_3369,N_2659,N_2533);
nand U3370 (N_3370,N_2665,N_2662);
or U3371 (N_3371,N_2865,N_2711);
or U3372 (N_3372,N_2797,N_2934);
nand U3373 (N_3373,N_2670,N_2649);
nand U3374 (N_3374,N_2704,N_2905);
nor U3375 (N_3375,N_2924,N_2834);
nor U3376 (N_3376,N_2691,N_2935);
nand U3377 (N_3377,N_2556,N_2790);
or U3378 (N_3378,N_2865,N_2718);
or U3379 (N_3379,N_2824,N_2968);
or U3380 (N_3380,N_2783,N_2632);
nand U3381 (N_3381,N_2597,N_2882);
and U3382 (N_3382,N_2949,N_2707);
nor U3383 (N_3383,N_2625,N_2818);
and U3384 (N_3384,N_2597,N_2725);
nor U3385 (N_3385,N_2979,N_2763);
and U3386 (N_3386,N_2994,N_2891);
nor U3387 (N_3387,N_2968,N_2562);
nand U3388 (N_3388,N_2593,N_2709);
nor U3389 (N_3389,N_2675,N_2767);
nor U3390 (N_3390,N_2659,N_2751);
and U3391 (N_3391,N_2688,N_2572);
or U3392 (N_3392,N_2705,N_2915);
nor U3393 (N_3393,N_2991,N_2670);
and U3394 (N_3394,N_2680,N_2978);
nor U3395 (N_3395,N_2913,N_2698);
and U3396 (N_3396,N_2868,N_2891);
and U3397 (N_3397,N_2787,N_2975);
nand U3398 (N_3398,N_2918,N_2788);
or U3399 (N_3399,N_2532,N_2630);
nand U3400 (N_3400,N_2524,N_2870);
and U3401 (N_3401,N_2707,N_2676);
and U3402 (N_3402,N_2500,N_2729);
or U3403 (N_3403,N_2897,N_2572);
nor U3404 (N_3404,N_2651,N_2525);
nor U3405 (N_3405,N_2778,N_2519);
and U3406 (N_3406,N_2610,N_2590);
nand U3407 (N_3407,N_2858,N_2533);
nor U3408 (N_3408,N_2888,N_2767);
and U3409 (N_3409,N_2882,N_2671);
and U3410 (N_3410,N_2986,N_2513);
or U3411 (N_3411,N_2611,N_2690);
and U3412 (N_3412,N_2878,N_2901);
nor U3413 (N_3413,N_2614,N_2823);
and U3414 (N_3414,N_2604,N_2568);
or U3415 (N_3415,N_2807,N_2544);
or U3416 (N_3416,N_2569,N_2672);
nor U3417 (N_3417,N_2845,N_2871);
xnor U3418 (N_3418,N_2778,N_2901);
nor U3419 (N_3419,N_2889,N_2815);
nand U3420 (N_3420,N_2852,N_2648);
or U3421 (N_3421,N_2750,N_2654);
or U3422 (N_3422,N_2546,N_2569);
nor U3423 (N_3423,N_2925,N_2833);
nor U3424 (N_3424,N_2587,N_2872);
or U3425 (N_3425,N_2755,N_2877);
nand U3426 (N_3426,N_2728,N_2606);
nor U3427 (N_3427,N_2635,N_2645);
and U3428 (N_3428,N_2720,N_2832);
or U3429 (N_3429,N_2749,N_2877);
and U3430 (N_3430,N_2618,N_2719);
or U3431 (N_3431,N_2834,N_2519);
nor U3432 (N_3432,N_2850,N_2940);
and U3433 (N_3433,N_2523,N_2810);
or U3434 (N_3434,N_2966,N_2614);
nor U3435 (N_3435,N_2942,N_2861);
nor U3436 (N_3436,N_2799,N_2674);
nor U3437 (N_3437,N_2989,N_2702);
and U3438 (N_3438,N_2873,N_2642);
nand U3439 (N_3439,N_2993,N_2827);
and U3440 (N_3440,N_2688,N_2756);
nor U3441 (N_3441,N_2849,N_2959);
nand U3442 (N_3442,N_2884,N_2727);
and U3443 (N_3443,N_2618,N_2718);
or U3444 (N_3444,N_2790,N_2887);
nand U3445 (N_3445,N_2819,N_2719);
or U3446 (N_3446,N_2774,N_2696);
nor U3447 (N_3447,N_2532,N_2774);
nor U3448 (N_3448,N_2752,N_2645);
and U3449 (N_3449,N_2993,N_2590);
and U3450 (N_3450,N_2560,N_2696);
nor U3451 (N_3451,N_2817,N_2517);
nor U3452 (N_3452,N_2685,N_2955);
nor U3453 (N_3453,N_2538,N_2840);
nor U3454 (N_3454,N_2997,N_2909);
nor U3455 (N_3455,N_2588,N_2803);
or U3456 (N_3456,N_2974,N_2843);
nor U3457 (N_3457,N_2617,N_2999);
and U3458 (N_3458,N_2891,N_2789);
or U3459 (N_3459,N_2976,N_2930);
and U3460 (N_3460,N_2969,N_2889);
or U3461 (N_3461,N_2591,N_2839);
or U3462 (N_3462,N_2703,N_2715);
or U3463 (N_3463,N_2750,N_2824);
nor U3464 (N_3464,N_2893,N_2669);
nor U3465 (N_3465,N_2734,N_2764);
or U3466 (N_3466,N_2802,N_2601);
or U3467 (N_3467,N_2638,N_2701);
nor U3468 (N_3468,N_2783,N_2652);
or U3469 (N_3469,N_2675,N_2964);
nor U3470 (N_3470,N_2837,N_2586);
and U3471 (N_3471,N_2995,N_2698);
or U3472 (N_3472,N_2976,N_2631);
or U3473 (N_3473,N_2750,N_2893);
or U3474 (N_3474,N_2589,N_2645);
nor U3475 (N_3475,N_2821,N_2887);
nand U3476 (N_3476,N_2646,N_2743);
nand U3477 (N_3477,N_2846,N_2723);
or U3478 (N_3478,N_2940,N_2594);
nor U3479 (N_3479,N_2921,N_2934);
nor U3480 (N_3480,N_2604,N_2932);
nand U3481 (N_3481,N_2593,N_2797);
nand U3482 (N_3482,N_2849,N_2904);
or U3483 (N_3483,N_2617,N_2720);
or U3484 (N_3484,N_2547,N_2627);
nand U3485 (N_3485,N_2788,N_2656);
xor U3486 (N_3486,N_2742,N_2916);
nor U3487 (N_3487,N_2743,N_2865);
nor U3488 (N_3488,N_2521,N_2592);
and U3489 (N_3489,N_2784,N_2709);
xor U3490 (N_3490,N_2965,N_2713);
nand U3491 (N_3491,N_2613,N_2765);
nand U3492 (N_3492,N_2519,N_2682);
nand U3493 (N_3493,N_2841,N_2687);
nand U3494 (N_3494,N_2610,N_2614);
nand U3495 (N_3495,N_2597,N_2692);
nand U3496 (N_3496,N_2767,N_2592);
nand U3497 (N_3497,N_2609,N_2562);
and U3498 (N_3498,N_2784,N_2681);
and U3499 (N_3499,N_2904,N_2812);
nor U3500 (N_3500,N_3474,N_3000);
nor U3501 (N_3501,N_3336,N_3137);
nand U3502 (N_3502,N_3182,N_3268);
or U3503 (N_3503,N_3105,N_3296);
nand U3504 (N_3504,N_3347,N_3155);
and U3505 (N_3505,N_3381,N_3353);
or U3506 (N_3506,N_3255,N_3305);
and U3507 (N_3507,N_3470,N_3188);
nor U3508 (N_3508,N_3042,N_3205);
nor U3509 (N_3509,N_3372,N_3186);
and U3510 (N_3510,N_3266,N_3049);
or U3511 (N_3511,N_3242,N_3120);
nor U3512 (N_3512,N_3425,N_3262);
nand U3513 (N_3513,N_3030,N_3265);
nor U3514 (N_3514,N_3085,N_3253);
or U3515 (N_3515,N_3061,N_3244);
nor U3516 (N_3516,N_3204,N_3481);
nand U3517 (N_3517,N_3286,N_3412);
and U3518 (N_3518,N_3064,N_3306);
or U3519 (N_3519,N_3135,N_3366);
nand U3520 (N_3520,N_3029,N_3348);
xnor U3521 (N_3521,N_3373,N_3415);
nand U3522 (N_3522,N_3399,N_3054);
nor U3523 (N_3523,N_3050,N_3014);
nor U3524 (N_3524,N_3375,N_3156);
nor U3525 (N_3525,N_3220,N_3334);
nor U3526 (N_3526,N_3411,N_3307);
nand U3527 (N_3527,N_3312,N_3012);
or U3528 (N_3528,N_3211,N_3047);
nor U3529 (N_3529,N_3421,N_3221);
nor U3530 (N_3530,N_3429,N_3100);
nand U3531 (N_3531,N_3232,N_3361);
or U3532 (N_3532,N_3489,N_3403);
nand U3533 (N_3533,N_3027,N_3450);
and U3534 (N_3534,N_3349,N_3033);
or U3535 (N_3535,N_3330,N_3274);
and U3536 (N_3536,N_3081,N_3059);
and U3537 (N_3537,N_3010,N_3031);
nand U3538 (N_3538,N_3230,N_3319);
nand U3539 (N_3539,N_3432,N_3393);
nor U3540 (N_3540,N_3289,N_3037);
and U3541 (N_3541,N_3413,N_3351);
nor U3542 (N_3542,N_3368,N_3103);
and U3543 (N_3543,N_3091,N_3370);
nor U3544 (N_3544,N_3102,N_3422);
or U3545 (N_3545,N_3486,N_3391);
nor U3546 (N_3546,N_3028,N_3377);
nor U3547 (N_3547,N_3068,N_3036);
nor U3548 (N_3548,N_3109,N_3325);
and U3549 (N_3549,N_3404,N_3076);
nor U3550 (N_3550,N_3476,N_3473);
or U3551 (N_3551,N_3389,N_3339);
nand U3552 (N_3552,N_3275,N_3408);
or U3553 (N_3553,N_3157,N_3176);
and U3554 (N_3554,N_3199,N_3226);
nor U3555 (N_3555,N_3446,N_3099);
or U3556 (N_3556,N_3097,N_3075);
nand U3557 (N_3557,N_3024,N_3066);
nor U3558 (N_3558,N_3082,N_3487);
and U3559 (N_3559,N_3189,N_3171);
nor U3560 (N_3560,N_3235,N_3332);
and U3561 (N_3561,N_3417,N_3467);
nor U3562 (N_3562,N_3313,N_3290);
nand U3563 (N_3563,N_3113,N_3087);
or U3564 (N_3564,N_3447,N_3115);
or U3565 (N_3565,N_3406,N_3227);
nor U3566 (N_3566,N_3214,N_3045);
nor U3567 (N_3567,N_3496,N_3371);
or U3568 (N_3568,N_3111,N_3299);
nand U3569 (N_3569,N_3346,N_3472);
or U3570 (N_3570,N_3090,N_3453);
or U3571 (N_3571,N_3207,N_3302);
or U3572 (N_3572,N_3252,N_3094);
or U3573 (N_3573,N_3023,N_3224);
nor U3574 (N_3574,N_3292,N_3471);
nand U3575 (N_3575,N_3291,N_3271);
nor U3576 (N_3576,N_3151,N_3078);
or U3577 (N_3577,N_3365,N_3132);
nor U3578 (N_3578,N_3177,N_3048);
nor U3579 (N_3579,N_3465,N_3044);
or U3580 (N_3580,N_3294,N_3492);
or U3581 (N_3581,N_3498,N_3152);
and U3582 (N_3582,N_3164,N_3469);
or U3583 (N_3583,N_3251,N_3070);
nor U3584 (N_3584,N_3246,N_3195);
and U3585 (N_3585,N_3213,N_3180);
or U3586 (N_3586,N_3034,N_3279);
or U3587 (N_3587,N_3172,N_3258);
nand U3588 (N_3588,N_3146,N_3394);
nand U3589 (N_3589,N_3430,N_3245);
and U3590 (N_3590,N_3276,N_3494);
and U3591 (N_3591,N_3369,N_3285);
xor U3592 (N_3592,N_3114,N_3280);
nand U3593 (N_3593,N_3136,N_3468);
nand U3594 (N_3594,N_3269,N_3239);
nor U3595 (N_3595,N_3362,N_3181);
or U3596 (N_3596,N_3005,N_3298);
or U3597 (N_3597,N_3052,N_3456);
and U3598 (N_3598,N_3193,N_3317);
nand U3599 (N_3599,N_3236,N_3179);
and U3600 (N_3600,N_3122,N_3021);
and U3601 (N_3601,N_3046,N_3287);
and U3602 (N_3602,N_3163,N_3282);
or U3603 (N_3603,N_3215,N_3378);
nor U3604 (N_3604,N_3022,N_3327);
and U3605 (N_3605,N_3457,N_3088);
or U3606 (N_3606,N_3444,N_3400);
nor U3607 (N_3607,N_3416,N_3101);
or U3608 (N_3608,N_3301,N_3475);
xor U3609 (N_3609,N_3315,N_3055);
or U3610 (N_3610,N_3324,N_3187);
nand U3611 (N_3611,N_3360,N_3013);
or U3612 (N_3612,N_3223,N_3126);
nand U3613 (N_3613,N_3154,N_3060);
nand U3614 (N_3614,N_3237,N_3462);
nor U3615 (N_3615,N_3284,N_3147);
or U3616 (N_3616,N_3428,N_3380);
nand U3617 (N_3617,N_3019,N_3201);
or U3618 (N_3618,N_3383,N_3166);
or U3619 (N_3619,N_3278,N_3104);
and U3620 (N_3620,N_3004,N_3162);
nand U3621 (N_3621,N_3263,N_3144);
nand U3622 (N_3622,N_3148,N_3451);
nor U3623 (N_3623,N_3058,N_3238);
nand U3624 (N_3624,N_3379,N_3077);
nor U3625 (N_3625,N_3455,N_3397);
or U3626 (N_3626,N_3420,N_3130);
nand U3627 (N_3627,N_3338,N_3234);
and U3628 (N_3628,N_3056,N_3020);
or U3629 (N_3629,N_3203,N_3198);
nand U3630 (N_3630,N_3478,N_3174);
and U3631 (N_3631,N_3441,N_3001);
nand U3632 (N_3632,N_3337,N_3431);
nor U3633 (N_3633,N_3304,N_3288);
and U3634 (N_3634,N_3173,N_3384);
nand U3635 (N_3635,N_3386,N_3131);
xnor U3636 (N_3636,N_3159,N_3150);
nor U3637 (N_3637,N_3231,N_3364);
or U3638 (N_3638,N_3409,N_3035);
nand U3639 (N_3639,N_3065,N_3062);
nor U3640 (N_3640,N_3356,N_3320);
nor U3641 (N_3641,N_3488,N_3323);
nand U3642 (N_3642,N_3321,N_3141);
nor U3643 (N_3643,N_3350,N_3390);
nor U3644 (N_3644,N_3424,N_3032);
and U3645 (N_3645,N_3281,N_3098);
nor U3646 (N_3646,N_3250,N_3210);
xnor U3647 (N_3647,N_3463,N_3359);
and U3648 (N_3648,N_3303,N_3329);
nor U3649 (N_3649,N_3084,N_3459);
nand U3650 (N_3650,N_3343,N_3477);
nand U3651 (N_3651,N_3039,N_3086);
nand U3652 (N_3652,N_3015,N_3192);
nand U3653 (N_3653,N_3106,N_3016);
nand U3654 (N_3654,N_3092,N_3200);
or U3655 (N_3655,N_3143,N_3074);
and U3656 (N_3656,N_3376,N_3121);
xnor U3657 (N_3657,N_3443,N_3483);
nor U3658 (N_3658,N_3308,N_3485);
or U3659 (N_3659,N_3040,N_3057);
nand U3660 (N_3660,N_3388,N_3335);
or U3661 (N_3661,N_3112,N_3125);
and U3662 (N_3662,N_3003,N_3093);
nor U3663 (N_3663,N_3160,N_3426);
nand U3664 (N_3664,N_3352,N_3316);
and U3665 (N_3665,N_3161,N_3017);
nor U3666 (N_3666,N_3196,N_3079);
or U3667 (N_3667,N_3018,N_3354);
or U3668 (N_3668,N_3295,N_3318);
or U3669 (N_3669,N_3395,N_3293);
and U3670 (N_3670,N_3405,N_3260);
or U3671 (N_3671,N_3493,N_3026);
or U3672 (N_3672,N_3149,N_3460);
and U3673 (N_3673,N_3217,N_3466);
nand U3674 (N_3674,N_3449,N_3358);
or U3675 (N_3675,N_3256,N_3249);
or U3676 (N_3676,N_3414,N_3464);
nand U3677 (N_3677,N_3233,N_3490);
nor U3678 (N_3678,N_3385,N_3438);
nor U3679 (N_3679,N_3427,N_3208);
nor U3680 (N_3680,N_3401,N_3259);
and U3681 (N_3681,N_3297,N_3300);
nor U3682 (N_3682,N_3439,N_3340);
nor U3683 (N_3683,N_3442,N_3071);
or U3684 (N_3684,N_3202,N_3218);
or U3685 (N_3685,N_3219,N_3479);
nand U3686 (N_3686,N_3452,N_3168);
nor U3687 (N_3687,N_3435,N_3491);
nor U3688 (N_3688,N_3434,N_3326);
or U3689 (N_3689,N_3261,N_3053);
or U3690 (N_3690,N_3212,N_3345);
or U3691 (N_3691,N_3341,N_3433);
nand U3692 (N_3692,N_3423,N_3095);
nand U3693 (N_3693,N_3096,N_3191);
or U3694 (N_3694,N_3264,N_3480);
and U3695 (N_3695,N_3225,N_3119);
and U3696 (N_3696,N_3254,N_3407);
or U3697 (N_3697,N_3272,N_3138);
nor U3698 (N_3698,N_3170,N_3002);
nor U3699 (N_3699,N_3140,N_3216);
and U3700 (N_3700,N_3185,N_3398);
and U3701 (N_3701,N_3041,N_3310);
nand U3702 (N_3702,N_3243,N_3038);
or U3703 (N_3703,N_3153,N_3314);
nand U3704 (N_3704,N_3367,N_3197);
and U3705 (N_3705,N_3117,N_3437);
or U3706 (N_3706,N_3333,N_3178);
nor U3707 (N_3707,N_3374,N_3110);
nor U3708 (N_3708,N_3145,N_3241);
or U3709 (N_3709,N_3089,N_3183);
and U3710 (N_3710,N_3497,N_3248);
and U3711 (N_3711,N_3129,N_3134);
and U3712 (N_3712,N_3283,N_3402);
and U3713 (N_3713,N_3167,N_3495);
xnor U3714 (N_3714,N_3116,N_3229);
and U3715 (N_3715,N_3277,N_3382);
nor U3716 (N_3716,N_3007,N_3273);
or U3717 (N_3717,N_3107,N_3328);
or U3718 (N_3718,N_3133,N_3169);
and U3719 (N_3719,N_3387,N_3436);
nor U3720 (N_3720,N_3458,N_3445);
nor U3721 (N_3721,N_3194,N_3461);
nand U3722 (N_3722,N_3396,N_3222);
or U3723 (N_3723,N_3051,N_3175);
or U3724 (N_3724,N_3331,N_3209);
nand U3725 (N_3725,N_3009,N_3228);
nand U3726 (N_3726,N_3083,N_3484);
and U3727 (N_3727,N_3190,N_3184);
nand U3728 (N_3728,N_3069,N_3322);
nor U3729 (N_3729,N_3142,N_3499);
and U3730 (N_3730,N_3355,N_3342);
or U3731 (N_3731,N_3008,N_3309);
or U3732 (N_3732,N_3206,N_3419);
or U3733 (N_3733,N_3344,N_3454);
nor U3734 (N_3734,N_3043,N_3357);
xor U3735 (N_3735,N_3108,N_3418);
nand U3736 (N_3736,N_3247,N_3128);
and U3737 (N_3737,N_3073,N_3311);
nor U3738 (N_3738,N_3006,N_3139);
or U3739 (N_3739,N_3482,N_3158);
nor U3740 (N_3740,N_3363,N_3011);
and U3741 (N_3741,N_3165,N_3267);
or U3742 (N_3742,N_3025,N_3410);
and U3743 (N_3743,N_3063,N_3270);
nand U3744 (N_3744,N_3072,N_3440);
and U3745 (N_3745,N_3240,N_3448);
nor U3746 (N_3746,N_3067,N_3127);
nor U3747 (N_3747,N_3118,N_3257);
nand U3748 (N_3748,N_3080,N_3124);
or U3749 (N_3749,N_3123,N_3392);
nor U3750 (N_3750,N_3000,N_3419);
nor U3751 (N_3751,N_3397,N_3327);
nand U3752 (N_3752,N_3047,N_3221);
nand U3753 (N_3753,N_3380,N_3196);
and U3754 (N_3754,N_3440,N_3368);
nand U3755 (N_3755,N_3249,N_3020);
and U3756 (N_3756,N_3475,N_3002);
and U3757 (N_3757,N_3168,N_3435);
nand U3758 (N_3758,N_3002,N_3205);
or U3759 (N_3759,N_3202,N_3344);
and U3760 (N_3760,N_3465,N_3113);
nand U3761 (N_3761,N_3123,N_3075);
or U3762 (N_3762,N_3133,N_3019);
or U3763 (N_3763,N_3333,N_3486);
nor U3764 (N_3764,N_3377,N_3078);
or U3765 (N_3765,N_3093,N_3253);
nand U3766 (N_3766,N_3184,N_3087);
and U3767 (N_3767,N_3202,N_3057);
nor U3768 (N_3768,N_3341,N_3268);
nand U3769 (N_3769,N_3151,N_3107);
or U3770 (N_3770,N_3286,N_3225);
nand U3771 (N_3771,N_3097,N_3021);
and U3772 (N_3772,N_3285,N_3426);
and U3773 (N_3773,N_3079,N_3418);
or U3774 (N_3774,N_3266,N_3279);
nor U3775 (N_3775,N_3356,N_3020);
nand U3776 (N_3776,N_3105,N_3214);
and U3777 (N_3777,N_3024,N_3128);
and U3778 (N_3778,N_3152,N_3001);
nor U3779 (N_3779,N_3131,N_3037);
or U3780 (N_3780,N_3013,N_3383);
and U3781 (N_3781,N_3216,N_3267);
nor U3782 (N_3782,N_3007,N_3204);
and U3783 (N_3783,N_3111,N_3391);
or U3784 (N_3784,N_3244,N_3423);
and U3785 (N_3785,N_3437,N_3045);
nor U3786 (N_3786,N_3345,N_3170);
or U3787 (N_3787,N_3017,N_3495);
nor U3788 (N_3788,N_3117,N_3251);
or U3789 (N_3789,N_3360,N_3129);
and U3790 (N_3790,N_3201,N_3458);
and U3791 (N_3791,N_3267,N_3353);
nand U3792 (N_3792,N_3413,N_3068);
nor U3793 (N_3793,N_3412,N_3113);
nor U3794 (N_3794,N_3219,N_3083);
and U3795 (N_3795,N_3352,N_3208);
and U3796 (N_3796,N_3344,N_3292);
and U3797 (N_3797,N_3091,N_3037);
or U3798 (N_3798,N_3464,N_3412);
nand U3799 (N_3799,N_3216,N_3291);
and U3800 (N_3800,N_3094,N_3073);
or U3801 (N_3801,N_3011,N_3030);
and U3802 (N_3802,N_3340,N_3266);
and U3803 (N_3803,N_3052,N_3419);
or U3804 (N_3804,N_3362,N_3357);
or U3805 (N_3805,N_3390,N_3464);
or U3806 (N_3806,N_3350,N_3273);
xnor U3807 (N_3807,N_3120,N_3262);
nand U3808 (N_3808,N_3244,N_3222);
or U3809 (N_3809,N_3338,N_3068);
nor U3810 (N_3810,N_3135,N_3430);
nand U3811 (N_3811,N_3007,N_3406);
or U3812 (N_3812,N_3138,N_3337);
nand U3813 (N_3813,N_3023,N_3282);
and U3814 (N_3814,N_3417,N_3466);
nand U3815 (N_3815,N_3327,N_3412);
and U3816 (N_3816,N_3449,N_3243);
and U3817 (N_3817,N_3438,N_3284);
xnor U3818 (N_3818,N_3169,N_3002);
or U3819 (N_3819,N_3278,N_3006);
nand U3820 (N_3820,N_3051,N_3413);
nand U3821 (N_3821,N_3017,N_3197);
or U3822 (N_3822,N_3045,N_3268);
nor U3823 (N_3823,N_3116,N_3309);
and U3824 (N_3824,N_3434,N_3486);
or U3825 (N_3825,N_3071,N_3019);
nor U3826 (N_3826,N_3477,N_3313);
nor U3827 (N_3827,N_3141,N_3332);
or U3828 (N_3828,N_3208,N_3369);
nand U3829 (N_3829,N_3492,N_3081);
nand U3830 (N_3830,N_3162,N_3213);
nand U3831 (N_3831,N_3404,N_3016);
nand U3832 (N_3832,N_3372,N_3101);
nor U3833 (N_3833,N_3286,N_3436);
nand U3834 (N_3834,N_3265,N_3003);
or U3835 (N_3835,N_3175,N_3075);
or U3836 (N_3836,N_3160,N_3095);
nand U3837 (N_3837,N_3114,N_3271);
and U3838 (N_3838,N_3454,N_3238);
and U3839 (N_3839,N_3141,N_3252);
nand U3840 (N_3840,N_3284,N_3420);
nand U3841 (N_3841,N_3395,N_3282);
nor U3842 (N_3842,N_3042,N_3097);
nand U3843 (N_3843,N_3092,N_3368);
or U3844 (N_3844,N_3066,N_3209);
nor U3845 (N_3845,N_3113,N_3225);
nor U3846 (N_3846,N_3457,N_3135);
nor U3847 (N_3847,N_3105,N_3409);
and U3848 (N_3848,N_3196,N_3401);
nand U3849 (N_3849,N_3167,N_3369);
or U3850 (N_3850,N_3300,N_3309);
nand U3851 (N_3851,N_3333,N_3257);
and U3852 (N_3852,N_3384,N_3439);
nand U3853 (N_3853,N_3399,N_3039);
and U3854 (N_3854,N_3317,N_3380);
or U3855 (N_3855,N_3020,N_3491);
nor U3856 (N_3856,N_3457,N_3378);
or U3857 (N_3857,N_3139,N_3257);
nand U3858 (N_3858,N_3033,N_3470);
and U3859 (N_3859,N_3234,N_3147);
or U3860 (N_3860,N_3474,N_3370);
and U3861 (N_3861,N_3335,N_3363);
and U3862 (N_3862,N_3244,N_3015);
nand U3863 (N_3863,N_3497,N_3017);
nor U3864 (N_3864,N_3191,N_3062);
nand U3865 (N_3865,N_3231,N_3337);
nor U3866 (N_3866,N_3455,N_3207);
nor U3867 (N_3867,N_3486,N_3281);
nand U3868 (N_3868,N_3375,N_3356);
nor U3869 (N_3869,N_3366,N_3237);
nor U3870 (N_3870,N_3484,N_3467);
or U3871 (N_3871,N_3180,N_3444);
nor U3872 (N_3872,N_3396,N_3047);
and U3873 (N_3873,N_3166,N_3424);
nand U3874 (N_3874,N_3223,N_3271);
and U3875 (N_3875,N_3395,N_3193);
nand U3876 (N_3876,N_3482,N_3072);
nand U3877 (N_3877,N_3495,N_3440);
nor U3878 (N_3878,N_3129,N_3000);
nor U3879 (N_3879,N_3214,N_3288);
nor U3880 (N_3880,N_3005,N_3183);
or U3881 (N_3881,N_3311,N_3366);
nor U3882 (N_3882,N_3044,N_3384);
or U3883 (N_3883,N_3401,N_3283);
nor U3884 (N_3884,N_3014,N_3260);
nor U3885 (N_3885,N_3160,N_3269);
nor U3886 (N_3886,N_3461,N_3212);
nand U3887 (N_3887,N_3351,N_3027);
or U3888 (N_3888,N_3113,N_3413);
nand U3889 (N_3889,N_3107,N_3339);
nor U3890 (N_3890,N_3079,N_3021);
or U3891 (N_3891,N_3128,N_3048);
or U3892 (N_3892,N_3340,N_3198);
nor U3893 (N_3893,N_3223,N_3491);
and U3894 (N_3894,N_3369,N_3049);
nand U3895 (N_3895,N_3198,N_3249);
nand U3896 (N_3896,N_3418,N_3461);
or U3897 (N_3897,N_3003,N_3419);
nand U3898 (N_3898,N_3373,N_3234);
and U3899 (N_3899,N_3424,N_3357);
or U3900 (N_3900,N_3338,N_3064);
and U3901 (N_3901,N_3033,N_3178);
or U3902 (N_3902,N_3015,N_3079);
nor U3903 (N_3903,N_3337,N_3145);
nor U3904 (N_3904,N_3257,N_3115);
nand U3905 (N_3905,N_3142,N_3167);
and U3906 (N_3906,N_3287,N_3446);
nand U3907 (N_3907,N_3315,N_3073);
nor U3908 (N_3908,N_3481,N_3099);
nand U3909 (N_3909,N_3283,N_3265);
nor U3910 (N_3910,N_3337,N_3232);
and U3911 (N_3911,N_3047,N_3253);
nand U3912 (N_3912,N_3099,N_3167);
nor U3913 (N_3913,N_3303,N_3388);
or U3914 (N_3914,N_3024,N_3440);
and U3915 (N_3915,N_3001,N_3291);
or U3916 (N_3916,N_3182,N_3437);
or U3917 (N_3917,N_3421,N_3414);
nand U3918 (N_3918,N_3216,N_3480);
or U3919 (N_3919,N_3334,N_3052);
nand U3920 (N_3920,N_3092,N_3018);
nor U3921 (N_3921,N_3071,N_3353);
nor U3922 (N_3922,N_3157,N_3489);
nand U3923 (N_3923,N_3254,N_3398);
or U3924 (N_3924,N_3061,N_3167);
or U3925 (N_3925,N_3071,N_3179);
nor U3926 (N_3926,N_3351,N_3174);
nand U3927 (N_3927,N_3046,N_3030);
and U3928 (N_3928,N_3228,N_3091);
nor U3929 (N_3929,N_3055,N_3242);
or U3930 (N_3930,N_3265,N_3339);
nand U3931 (N_3931,N_3044,N_3283);
nand U3932 (N_3932,N_3382,N_3290);
xor U3933 (N_3933,N_3086,N_3415);
or U3934 (N_3934,N_3326,N_3152);
or U3935 (N_3935,N_3189,N_3489);
nand U3936 (N_3936,N_3368,N_3191);
or U3937 (N_3937,N_3119,N_3257);
nand U3938 (N_3938,N_3165,N_3026);
nand U3939 (N_3939,N_3449,N_3273);
or U3940 (N_3940,N_3250,N_3272);
or U3941 (N_3941,N_3280,N_3382);
nand U3942 (N_3942,N_3339,N_3118);
and U3943 (N_3943,N_3041,N_3009);
nand U3944 (N_3944,N_3494,N_3158);
nand U3945 (N_3945,N_3248,N_3436);
and U3946 (N_3946,N_3437,N_3268);
nor U3947 (N_3947,N_3154,N_3163);
or U3948 (N_3948,N_3238,N_3448);
and U3949 (N_3949,N_3014,N_3261);
or U3950 (N_3950,N_3003,N_3440);
nor U3951 (N_3951,N_3054,N_3037);
nor U3952 (N_3952,N_3207,N_3411);
nand U3953 (N_3953,N_3086,N_3186);
nand U3954 (N_3954,N_3025,N_3226);
or U3955 (N_3955,N_3359,N_3325);
nor U3956 (N_3956,N_3079,N_3202);
and U3957 (N_3957,N_3374,N_3066);
or U3958 (N_3958,N_3143,N_3408);
nor U3959 (N_3959,N_3328,N_3348);
nor U3960 (N_3960,N_3136,N_3014);
and U3961 (N_3961,N_3493,N_3043);
or U3962 (N_3962,N_3400,N_3387);
and U3963 (N_3963,N_3387,N_3234);
nor U3964 (N_3964,N_3053,N_3243);
or U3965 (N_3965,N_3219,N_3478);
or U3966 (N_3966,N_3371,N_3312);
nand U3967 (N_3967,N_3087,N_3010);
and U3968 (N_3968,N_3054,N_3113);
or U3969 (N_3969,N_3202,N_3001);
nand U3970 (N_3970,N_3108,N_3367);
and U3971 (N_3971,N_3182,N_3271);
nand U3972 (N_3972,N_3034,N_3035);
or U3973 (N_3973,N_3481,N_3154);
nand U3974 (N_3974,N_3118,N_3427);
or U3975 (N_3975,N_3185,N_3405);
and U3976 (N_3976,N_3288,N_3071);
or U3977 (N_3977,N_3021,N_3082);
nand U3978 (N_3978,N_3328,N_3273);
and U3979 (N_3979,N_3026,N_3006);
nor U3980 (N_3980,N_3312,N_3131);
nand U3981 (N_3981,N_3068,N_3370);
or U3982 (N_3982,N_3330,N_3062);
nor U3983 (N_3983,N_3179,N_3095);
and U3984 (N_3984,N_3194,N_3354);
xnor U3985 (N_3985,N_3241,N_3069);
and U3986 (N_3986,N_3155,N_3278);
nor U3987 (N_3987,N_3307,N_3285);
and U3988 (N_3988,N_3440,N_3164);
nand U3989 (N_3989,N_3411,N_3449);
or U3990 (N_3990,N_3412,N_3305);
and U3991 (N_3991,N_3425,N_3304);
or U3992 (N_3992,N_3091,N_3011);
nand U3993 (N_3993,N_3311,N_3255);
nor U3994 (N_3994,N_3364,N_3253);
and U3995 (N_3995,N_3370,N_3318);
nor U3996 (N_3996,N_3377,N_3480);
and U3997 (N_3997,N_3425,N_3396);
and U3998 (N_3998,N_3395,N_3353);
nor U3999 (N_3999,N_3287,N_3355);
nand U4000 (N_4000,N_3985,N_3912);
or U4001 (N_4001,N_3965,N_3510);
nor U4002 (N_4002,N_3562,N_3831);
xnor U4003 (N_4003,N_3757,N_3668);
xnor U4004 (N_4004,N_3826,N_3778);
and U4005 (N_4005,N_3901,N_3825);
or U4006 (N_4006,N_3730,N_3807);
nand U4007 (N_4007,N_3517,N_3950);
nand U4008 (N_4008,N_3819,N_3586);
nor U4009 (N_4009,N_3526,N_3560);
or U4010 (N_4010,N_3905,N_3556);
or U4011 (N_4011,N_3536,N_3899);
nor U4012 (N_4012,N_3610,N_3764);
and U4013 (N_4013,N_3916,N_3760);
and U4014 (N_4014,N_3928,N_3933);
and U4015 (N_4015,N_3902,N_3742);
and U4016 (N_4016,N_3660,N_3973);
or U4017 (N_4017,N_3789,N_3733);
and U4018 (N_4018,N_3615,N_3593);
nand U4019 (N_4019,N_3518,N_3587);
nand U4020 (N_4020,N_3860,N_3881);
nor U4021 (N_4021,N_3590,N_3867);
and U4022 (N_4022,N_3983,N_3704);
or U4023 (N_4023,N_3635,N_3670);
nand U4024 (N_4024,N_3618,N_3966);
and U4025 (N_4025,N_3833,N_3997);
nand U4026 (N_4026,N_3600,N_3781);
nor U4027 (N_4027,N_3845,N_3580);
nand U4028 (N_4028,N_3688,N_3666);
and U4029 (N_4029,N_3525,N_3565);
or U4030 (N_4030,N_3543,N_3793);
nor U4031 (N_4031,N_3754,N_3715);
nand U4032 (N_4032,N_3628,N_3703);
nor U4033 (N_4033,N_3541,N_3568);
and U4034 (N_4034,N_3577,N_3913);
nand U4035 (N_4035,N_3918,N_3980);
nand U4036 (N_4036,N_3741,N_3623);
nor U4037 (N_4037,N_3563,N_3995);
nand U4038 (N_4038,N_3837,N_3561);
or U4039 (N_4039,N_3520,N_3603);
nor U4040 (N_4040,N_3522,N_3751);
and U4041 (N_4041,N_3964,N_3683);
or U4042 (N_4042,N_3582,N_3842);
nor U4043 (N_4043,N_3524,N_3863);
or U4044 (N_4044,N_3967,N_3699);
or U4045 (N_4045,N_3925,N_3709);
nand U4046 (N_4046,N_3680,N_3874);
or U4047 (N_4047,N_3725,N_3803);
nand U4048 (N_4048,N_3970,N_3854);
and U4049 (N_4049,N_3707,N_3776);
xor U4050 (N_4050,N_3551,N_3639);
nor U4051 (N_4051,N_3534,N_3987);
nor U4052 (N_4052,N_3914,N_3936);
nor U4053 (N_4053,N_3975,N_3828);
nor U4054 (N_4054,N_3808,N_3662);
and U4055 (N_4055,N_3920,N_3927);
or U4056 (N_4056,N_3996,N_3578);
and U4057 (N_4057,N_3636,N_3546);
nand U4058 (N_4058,N_3759,N_3686);
nor U4059 (N_4059,N_3718,N_3992);
nand U4060 (N_4060,N_3511,N_3872);
and U4061 (N_4061,N_3566,N_3542);
or U4062 (N_4062,N_3609,N_3513);
and U4063 (N_4063,N_3711,N_3604);
or U4064 (N_4064,N_3951,N_3756);
nand U4065 (N_4065,N_3772,N_3801);
or U4066 (N_4066,N_3592,N_3583);
or U4067 (N_4067,N_3716,N_3829);
nand U4068 (N_4068,N_3953,N_3588);
or U4069 (N_4069,N_3750,N_3871);
nand U4070 (N_4070,N_3972,N_3572);
nand U4071 (N_4071,N_3642,N_3647);
nand U4072 (N_4072,N_3521,N_3601);
or U4073 (N_4073,N_3891,N_3653);
or U4074 (N_4074,N_3782,N_3728);
nor U4075 (N_4075,N_3768,N_3752);
nand U4076 (N_4076,N_3974,N_3700);
or U4077 (N_4077,N_3597,N_3625);
xnor U4078 (N_4078,N_3640,N_3948);
and U4079 (N_4079,N_3523,N_3570);
or U4080 (N_4080,N_3947,N_3806);
nor U4081 (N_4081,N_3573,N_3619);
or U4082 (N_4082,N_3994,N_3721);
or U4083 (N_4083,N_3851,N_3911);
or U4084 (N_4084,N_3797,N_3514);
nor U4085 (N_4085,N_3540,N_3701);
and U4086 (N_4086,N_3740,N_3931);
nor U4087 (N_4087,N_3836,N_3726);
or U4088 (N_4088,N_3919,N_3645);
and U4089 (N_4089,N_3755,N_3855);
nor U4090 (N_4090,N_3873,N_3922);
or U4091 (N_4091,N_3841,N_3569);
nand U4092 (N_4092,N_3900,N_3736);
nor U4093 (N_4093,N_3917,N_3866);
nor U4094 (N_4094,N_3702,N_3823);
xnor U4095 (N_4095,N_3611,N_3631);
or U4096 (N_4096,N_3676,N_3976);
nand U4097 (N_4097,N_3554,N_3839);
and U4098 (N_4098,N_3945,N_3719);
nor U4099 (N_4099,N_3545,N_3780);
nor U4100 (N_4100,N_3656,N_3870);
nand U4101 (N_4101,N_3838,N_3691);
nor U4102 (N_4102,N_3713,N_3658);
nand U4103 (N_4103,N_3633,N_3681);
or U4104 (N_4104,N_3811,N_3937);
and U4105 (N_4105,N_3977,N_3963);
nor U4106 (N_4106,N_3978,N_3739);
nor U4107 (N_4107,N_3960,N_3903);
nor U4108 (N_4108,N_3930,N_3706);
and U4109 (N_4109,N_3584,N_3575);
nand U4110 (N_4110,N_3850,N_3761);
or U4111 (N_4111,N_3880,N_3651);
and U4112 (N_4112,N_3904,N_3548);
nand U4113 (N_4113,N_3817,N_3506);
nand U4114 (N_4114,N_3895,N_3596);
and U4115 (N_4115,N_3832,N_3792);
nor U4116 (N_4116,N_3650,N_3763);
and U4117 (N_4117,N_3813,N_3652);
nand U4118 (N_4118,N_3884,N_3678);
nand U4119 (N_4119,N_3932,N_3737);
nor U4120 (N_4120,N_3939,N_3847);
and U4121 (N_4121,N_3698,N_3693);
or U4122 (N_4122,N_3538,N_3717);
nor U4123 (N_4123,N_3613,N_3815);
and U4124 (N_4124,N_3798,N_3720);
nand U4125 (N_4125,N_3910,N_3685);
and U4126 (N_4126,N_3794,N_3775);
nor U4127 (N_4127,N_3629,N_3557);
nand U4128 (N_4128,N_3766,N_3504);
nand U4129 (N_4129,N_3508,N_3677);
nor U4130 (N_4130,N_3800,N_3500);
and U4131 (N_4131,N_3567,N_3893);
nor U4132 (N_4132,N_3791,N_3859);
and U4133 (N_4133,N_3762,N_3649);
and U4134 (N_4134,N_3787,N_3594);
nand U4135 (N_4135,N_3991,N_3669);
nand U4136 (N_4136,N_3690,N_3888);
nor U4137 (N_4137,N_3559,N_3501);
nor U4138 (N_4138,N_3942,N_3537);
and U4139 (N_4139,N_3956,N_3887);
and U4140 (N_4140,N_3687,N_3955);
nand U4141 (N_4141,N_3984,N_3773);
and U4142 (N_4142,N_3555,N_3843);
and U4143 (N_4143,N_3796,N_3877);
or U4144 (N_4144,N_3878,N_3857);
and U4145 (N_4145,N_3862,N_3799);
and U4146 (N_4146,N_3599,N_3765);
or U4147 (N_4147,N_3824,N_3814);
or U4148 (N_4148,N_3503,N_3864);
nor U4149 (N_4149,N_3868,N_3509);
nor U4150 (N_4150,N_3858,N_3571);
and U4151 (N_4151,N_3889,N_3682);
and U4152 (N_4152,N_3705,N_3758);
or U4153 (N_4153,N_3883,N_3783);
and U4154 (N_4154,N_3897,N_3608);
and U4155 (N_4155,N_3969,N_3812);
nor U4156 (N_4156,N_3738,N_3602);
nor U4157 (N_4157,N_3989,N_3530);
nor U4158 (N_4158,N_3856,N_3674);
nand U4159 (N_4159,N_3830,N_3879);
nand U4160 (N_4160,N_3767,N_3809);
and U4161 (N_4161,N_3723,N_3923);
nand U4162 (N_4162,N_3753,N_3971);
nand U4163 (N_4163,N_3502,N_3954);
or U4164 (N_4164,N_3747,N_3938);
or U4165 (N_4165,N_3790,N_3531);
and U4166 (N_4166,N_3581,N_3894);
and U4167 (N_4167,N_3549,N_3654);
nand U4168 (N_4168,N_3946,N_3779);
xnor U4169 (N_4169,N_3614,N_3802);
nand U4170 (N_4170,N_3574,N_3885);
nand U4171 (N_4171,N_3852,N_3915);
and U4172 (N_4172,N_3550,N_3990);
nor U4173 (N_4173,N_3632,N_3708);
and U4174 (N_4174,N_3617,N_3528);
and U4175 (N_4175,N_3516,N_3999);
or U4176 (N_4176,N_3641,N_3710);
and U4177 (N_4177,N_3929,N_3553);
nand U4178 (N_4178,N_3876,N_3846);
and U4179 (N_4179,N_3646,N_3539);
or U4180 (N_4180,N_3732,N_3844);
nand U4181 (N_4181,N_3935,N_3890);
nor U4182 (N_4182,N_3770,N_3659);
and U4183 (N_4183,N_3907,N_3591);
nor U4184 (N_4184,N_3959,N_3952);
and U4185 (N_4185,N_3748,N_3626);
nand U4186 (N_4186,N_3692,N_3865);
nor U4187 (N_4187,N_3558,N_3598);
and U4188 (N_4188,N_3810,N_3684);
nand U4189 (N_4189,N_3667,N_3712);
or U4190 (N_4190,N_3777,N_3875);
nand U4191 (N_4191,N_3547,N_3630);
and U4192 (N_4192,N_3958,N_3786);
and U4193 (N_4193,N_3924,N_3949);
or U4194 (N_4194,N_3771,N_3535);
nand U4195 (N_4195,N_3697,N_3512);
or U4196 (N_4196,N_3507,N_3622);
nand U4197 (N_4197,N_3898,N_3605);
nand U4198 (N_4198,N_3993,N_3634);
nand U4199 (N_4199,N_3769,N_3818);
or U4200 (N_4200,N_3886,N_3988);
or U4201 (N_4201,N_3744,N_3627);
xnor U4202 (N_4202,N_3616,N_3784);
nor U4203 (N_4203,N_3962,N_3848);
xor U4204 (N_4204,N_3552,N_3944);
nor U4205 (N_4205,N_3743,N_3820);
nand U4206 (N_4206,N_3979,N_3735);
nor U4207 (N_4207,N_3729,N_3696);
or U4208 (N_4208,N_3657,N_3673);
nand U4209 (N_4209,N_3606,N_3816);
or U4210 (N_4210,N_3644,N_3861);
or U4211 (N_4211,N_3745,N_3595);
nand U4212 (N_4212,N_3638,N_3505);
and U4213 (N_4213,N_3795,N_3869);
nand U4214 (N_4214,N_3986,N_3805);
nand U4215 (N_4215,N_3661,N_3998);
nand U4216 (N_4216,N_3564,N_3694);
or U4217 (N_4217,N_3648,N_3620);
nand U4218 (N_4218,N_3957,N_3934);
nand U4219 (N_4219,N_3746,N_3940);
xor U4220 (N_4220,N_3822,N_3532);
nor U4221 (N_4221,N_3908,N_3679);
nor U4222 (N_4222,N_3734,N_3714);
nor U4223 (N_4223,N_3892,N_3621);
nor U4224 (N_4224,N_3827,N_3821);
nand U4225 (N_4225,N_3906,N_3788);
and U4226 (N_4226,N_3909,N_3941);
nand U4227 (N_4227,N_3982,N_3749);
nor U4228 (N_4228,N_3774,N_3664);
nand U4229 (N_4229,N_3675,N_3579);
nor U4230 (N_4230,N_3968,N_3724);
nor U4231 (N_4231,N_3943,N_3624);
and U4232 (N_4232,N_3527,N_3835);
nor U4233 (N_4233,N_3515,N_3544);
and U4234 (N_4234,N_3849,N_3607);
nor U4235 (N_4235,N_3804,N_3576);
and U4236 (N_4236,N_3882,N_3961);
nand U4237 (N_4237,N_3921,N_3529);
and U4238 (N_4238,N_3785,N_3533);
nor U4239 (N_4239,N_3637,N_3981);
nand U4240 (N_4240,N_3643,N_3519);
nand U4241 (N_4241,N_3689,N_3853);
and U4242 (N_4242,N_3672,N_3589);
nor U4243 (N_4243,N_3896,N_3727);
nand U4244 (N_4244,N_3671,N_3840);
nor U4245 (N_4245,N_3665,N_3612);
or U4246 (N_4246,N_3655,N_3731);
and U4247 (N_4247,N_3585,N_3663);
nand U4248 (N_4248,N_3695,N_3722);
or U4249 (N_4249,N_3834,N_3926);
or U4250 (N_4250,N_3970,N_3908);
nand U4251 (N_4251,N_3792,N_3991);
and U4252 (N_4252,N_3942,N_3548);
xor U4253 (N_4253,N_3849,N_3964);
or U4254 (N_4254,N_3581,N_3824);
nor U4255 (N_4255,N_3976,N_3782);
nor U4256 (N_4256,N_3539,N_3682);
and U4257 (N_4257,N_3928,N_3532);
nand U4258 (N_4258,N_3828,N_3863);
or U4259 (N_4259,N_3813,N_3920);
nor U4260 (N_4260,N_3873,N_3851);
or U4261 (N_4261,N_3659,N_3771);
nor U4262 (N_4262,N_3940,N_3617);
nor U4263 (N_4263,N_3834,N_3892);
or U4264 (N_4264,N_3776,N_3780);
or U4265 (N_4265,N_3673,N_3997);
nand U4266 (N_4266,N_3965,N_3977);
and U4267 (N_4267,N_3872,N_3533);
nor U4268 (N_4268,N_3731,N_3685);
nand U4269 (N_4269,N_3621,N_3628);
or U4270 (N_4270,N_3596,N_3771);
nor U4271 (N_4271,N_3994,N_3711);
or U4272 (N_4272,N_3811,N_3846);
or U4273 (N_4273,N_3956,N_3799);
nand U4274 (N_4274,N_3728,N_3564);
or U4275 (N_4275,N_3893,N_3569);
or U4276 (N_4276,N_3834,N_3605);
nand U4277 (N_4277,N_3544,N_3738);
or U4278 (N_4278,N_3863,N_3899);
or U4279 (N_4279,N_3515,N_3894);
nand U4280 (N_4280,N_3571,N_3880);
xor U4281 (N_4281,N_3981,N_3629);
nor U4282 (N_4282,N_3890,N_3507);
nand U4283 (N_4283,N_3833,N_3771);
nand U4284 (N_4284,N_3560,N_3651);
xnor U4285 (N_4285,N_3660,N_3956);
nand U4286 (N_4286,N_3806,N_3572);
nor U4287 (N_4287,N_3712,N_3561);
or U4288 (N_4288,N_3853,N_3901);
or U4289 (N_4289,N_3879,N_3623);
or U4290 (N_4290,N_3791,N_3763);
and U4291 (N_4291,N_3910,N_3735);
nor U4292 (N_4292,N_3633,N_3527);
or U4293 (N_4293,N_3546,N_3648);
nand U4294 (N_4294,N_3999,N_3938);
and U4295 (N_4295,N_3790,N_3544);
or U4296 (N_4296,N_3710,N_3779);
and U4297 (N_4297,N_3936,N_3988);
and U4298 (N_4298,N_3927,N_3898);
nand U4299 (N_4299,N_3935,N_3882);
or U4300 (N_4300,N_3784,N_3814);
or U4301 (N_4301,N_3846,N_3707);
nand U4302 (N_4302,N_3603,N_3645);
and U4303 (N_4303,N_3555,N_3867);
nor U4304 (N_4304,N_3904,N_3870);
and U4305 (N_4305,N_3755,N_3712);
nor U4306 (N_4306,N_3501,N_3954);
nor U4307 (N_4307,N_3758,N_3570);
nand U4308 (N_4308,N_3889,N_3567);
and U4309 (N_4309,N_3767,N_3664);
nand U4310 (N_4310,N_3907,N_3833);
xor U4311 (N_4311,N_3672,N_3922);
or U4312 (N_4312,N_3562,N_3575);
nor U4313 (N_4313,N_3680,N_3648);
nor U4314 (N_4314,N_3681,N_3716);
or U4315 (N_4315,N_3622,N_3781);
nand U4316 (N_4316,N_3775,N_3949);
nor U4317 (N_4317,N_3893,N_3543);
nor U4318 (N_4318,N_3522,N_3579);
nor U4319 (N_4319,N_3735,N_3798);
nand U4320 (N_4320,N_3980,N_3714);
nand U4321 (N_4321,N_3604,N_3856);
nand U4322 (N_4322,N_3906,N_3770);
or U4323 (N_4323,N_3845,N_3575);
and U4324 (N_4324,N_3649,N_3836);
and U4325 (N_4325,N_3649,N_3589);
and U4326 (N_4326,N_3938,N_3794);
nand U4327 (N_4327,N_3550,N_3749);
or U4328 (N_4328,N_3830,N_3510);
or U4329 (N_4329,N_3519,N_3979);
xnor U4330 (N_4330,N_3924,N_3569);
nand U4331 (N_4331,N_3928,N_3800);
and U4332 (N_4332,N_3941,N_3647);
and U4333 (N_4333,N_3825,N_3767);
and U4334 (N_4334,N_3949,N_3943);
nor U4335 (N_4335,N_3997,N_3722);
nand U4336 (N_4336,N_3597,N_3793);
or U4337 (N_4337,N_3700,N_3706);
and U4338 (N_4338,N_3640,N_3893);
and U4339 (N_4339,N_3670,N_3506);
nand U4340 (N_4340,N_3531,N_3984);
or U4341 (N_4341,N_3725,N_3750);
and U4342 (N_4342,N_3877,N_3750);
xnor U4343 (N_4343,N_3682,N_3866);
or U4344 (N_4344,N_3646,N_3939);
nor U4345 (N_4345,N_3641,N_3565);
nand U4346 (N_4346,N_3608,N_3772);
and U4347 (N_4347,N_3714,N_3764);
and U4348 (N_4348,N_3782,N_3894);
nor U4349 (N_4349,N_3702,N_3887);
and U4350 (N_4350,N_3514,N_3547);
nor U4351 (N_4351,N_3803,N_3812);
nor U4352 (N_4352,N_3696,N_3700);
and U4353 (N_4353,N_3801,N_3881);
or U4354 (N_4354,N_3938,N_3565);
nand U4355 (N_4355,N_3916,N_3910);
and U4356 (N_4356,N_3712,N_3751);
and U4357 (N_4357,N_3606,N_3862);
or U4358 (N_4358,N_3880,N_3601);
nor U4359 (N_4359,N_3818,N_3540);
nor U4360 (N_4360,N_3574,N_3725);
nand U4361 (N_4361,N_3909,N_3632);
nand U4362 (N_4362,N_3631,N_3511);
or U4363 (N_4363,N_3951,N_3932);
nor U4364 (N_4364,N_3532,N_3716);
nor U4365 (N_4365,N_3561,N_3729);
nand U4366 (N_4366,N_3826,N_3624);
nor U4367 (N_4367,N_3918,N_3648);
nor U4368 (N_4368,N_3711,N_3550);
and U4369 (N_4369,N_3530,N_3836);
or U4370 (N_4370,N_3655,N_3719);
and U4371 (N_4371,N_3611,N_3806);
nand U4372 (N_4372,N_3985,N_3560);
or U4373 (N_4373,N_3522,N_3628);
and U4374 (N_4374,N_3845,N_3592);
and U4375 (N_4375,N_3904,N_3816);
nor U4376 (N_4376,N_3948,N_3967);
nand U4377 (N_4377,N_3846,N_3722);
nand U4378 (N_4378,N_3787,N_3795);
nand U4379 (N_4379,N_3951,N_3720);
xnor U4380 (N_4380,N_3813,N_3873);
or U4381 (N_4381,N_3812,N_3800);
nand U4382 (N_4382,N_3924,N_3685);
and U4383 (N_4383,N_3602,N_3949);
nor U4384 (N_4384,N_3509,N_3689);
and U4385 (N_4385,N_3646,N_3798);
nand U4386 (N_4386,N_3638,N_3912);
and U4387 (N_4387,N_3772,N_3747);
nand U4388 (N_4388,N_3563,N_3628);
nor U4389 (N_4389,N_3960,N_3638);
nor U4390 (N_4390,N_3850,N_3953);
or U4391 (N_4391,N_3719,N_3677);
or U4392 (N_4392,N_3898,N_3616);
and U4393 (N_4393,N_3887,N_3695);
nor U4394 (N_4394,N_3771,N_3866);
xnor U4395 (N_4395,N_3946,N_3994);
or U4396 (N_4396,N_3741,N_3656);
nand U4397 (N_4397,N_3543,N_3833);
or U4398 (N_4398,N_3930,N_3874);
or U4399 (N_4399,N_3865,N_3564);
nor U4400 (N_4400,N_3677,N_3976);
or U4401 (N_4401,N_3566,N_3778);
nand U4402 (N_4402,N_3827,N_3839);
and U4403 (N_4403,N_3739,N_3932);
nor U4404 (N_4404,N_3821,N_3730);
nand U4405 (N_4405,N_3706,N_3515);
nor U4406 (N_4406,N_3595,N_3541);
nor U4407 (N_4407,N_3587,N_3502);
or U4408 (N_4408,N_3740,N_3981);
xnor U4409 (N_4409,N_3791,N_3747);
and U4410 (N_4410,N_3644,N_3716);
nand U4411 (N_4411,N_3546,N_3561);
or U4412 (N_4412,N_3700,N_3982);
nand U4413 (N_4413,N_3617,N_3856);
or U4414 (N_4414,N_3868,N_3702);
or U4415 (N_4415,N_3735,N_3616);
and U4416 (N_4416,N_3839,N_3928);
xor U4417 (N_4417,N_3815,N_3541);
xnor U4418 (N_4418,N_3770,N_3752);
or U4419 (N_4419,N_3592,N_3813);
and U4420 (N_4420,N_3558,N_3536);
and U4421 (N_4421,N_3792,N_3723);
and U4422 (N_4422,N_3933,N_3565);
nand U4423 (N_4423,N_3715,N_3546);
nand U4424 (N_4424,N_3656,N_3719);
xnor U4425 (N_4425,N_3543,N_3875);
or U4426 (N_4426,N_3753,N_3916);
or U4427 (N_4427,N_3708,N_3792);
nand U4428 (N_4428,N_3825,N_3596);
nand U4429 (N_4429,N_3843,N_3788);
and U4430 (N_4430,N_3646,N_3685);
or U4431 (N_4431,N_3672,N_3556);
xor U4432 (N_4432,N_3925,N_3544);
and U4433 (N_4433,N_3511,N_3738);
and U4434 (N_4434,N_3750,N_3879);
nor U4435 (N_4435,N_3842,N_3586);
and U4436 (N_4436,N_3567,N_3928);
or U4437 (N_4437,N_3859,N_3872);
nand U4438 (N_4438,N_3581,N_3813);
xor U4439 (N_4439,N_3558,N_3774);
and U4440 (N_4440,N_3638,N_3796);
and U4441 (N_4441,N_3647,N_3917);
and U4442 (N_4442,N_3544,N_3521);
and U4443 (N_4443,N_3871,N_3623);
nand U4444 (N_4444,N_3590,N_3743);
nor U4445 (N_4445,N_3606,N_3899);
nand U4446 (N_4446,N_3530,N_3562);
nor U4447 (N_4447,N_3747,N_3560);
or U4448 (N_4448,N_3911,N_3529);
nor U4449 (N_4449,N_3583,N_3545);
nand U4450 (N_4450,N_3662,N_3657);
or U4451 (N_4451,N_3884,N_3931);
nand U4452 (N_4452,N_3545,N_3697);
or U4453 (N_4453,N_3965,N_3787);
nor U4454 (N_4454,N_3674,N_3662);
nor U4455 (N_4455,N_3525,N_3833);
and U4456 (N_4456,N_3750,N_3739);
and U4457 (N_4457,N_3999,N_3576);
and U4458 (N_4458,N_3613,N_3757);
and U4459 (N_4459,N_3661,N_3718);
nor U4460 (N_4460,N_3923,N_3801);
or U4461 (N_4461,N_3830,N_3766);
and U4462 (N_4462,N_3508,N_3860);
nor U4463 (N_4463,N_3545,N_3678);
nand U4464 (N_4464,N_3589,N_3560);
or U4465 (N_4465,N_3749,N_3909);
and U4466 (N_4466,N_3851,N_3668);
xnor U4467 (N_4467,N_3677,N_3901);
or U4468 (N_4468,N_3955,N_3707);
nand U4469 (N_4469,N_3857,N_3622);
or U4470 (N_4470,N_3673,N_3915);
nor U4471 (N_4471,N_3932,N_3599);
nor U4472 (N_4472,N_3802,N_3965);
and U4473 (N_4473,N_3551,N_3918);
nor U4474 (N_4474,N_3996,N_3816);
nor U4475 (N_4475,N_3538,N_3888);
nor U4476 (N_4476,N_3529,N_3526);
or U4477 (N_4477,N_3714,N_3968);
nor U4478 (N_4478,N_3773,N_3581);
or U4479 (N_4479,N_3518,N_3805);
or U4480 (N_4480,N_3698,N_3758);
and U4481 (N_4481,N_3728,N_3998);
and U4482 (N_4482,N_3811,N_3865);
nand U4483 (N_4483,N_3562,N_3664);
and U4484 (N_4484,N_3643,N_3631);
nor U4485 (N_4485,N_3935,N_3650);
or U4486 (N_4486,N_3505,N_3839);
nor U4487 (N_4487,N_3568,N_3622);
or U4488 (N_4488,N_3917,N_3907);
and U4489 (N_4489,N_3602,N_3849);
xnor U4490 (N_4490,N_3677,N_3857);
nor U4491 (N_4491,N_3758,N_3704);
and U4492 (N_4492,N_3674,N_3624);
nand U4493 (N_4493,N_3854,N_3670);
or U4494 (N_4494,N_3676,N_3943);
or U4495 (N_4495,N_3894,N_3540);
nor U4496 (N_4496,N_3888,N_3875);
or U4497 (N_4497,N_3515,N_3956);
and U4498 (N_4498,N_3752,N_3819);
nor U4499 (N_4499,N_3889,N_3734);
or U4500 (N_4500,N_4352,N_4328);
and U4501 (N_4501,N_4499,N_4423);
or U4502 (N_4502,N_4173,N_4120);
or U4503 (N_4503,N_4222,N_4064);
nand U4504 (N_4504,N_4250,N_4284);
and U4505 (N_4505,N_4267,N_4391);
nor U4506 (N_4506,N_4124,N_4459);
nand U4507 (N_4507,N_4096,N_4119);
nor U4508 (N_4508,N_4287,N_4341);
xnor U4509 (N_4509,N_4445,N_4439);
and U4510 (N_4510,N_4159,N_4342);
or U4511 (N_4511,N_4481,N_4355);
nand U4512 (N_4512,N_4377,N_4407);
nor U4513 (N_4513,N_4312,N_4310);
nand U4514 (N_4514,N_4288,N_4317);
and U4515 (N_4515,N_4474,N_4118);
or U4516 (N_4516,N_4327,N_4145);
nor U4517 (N_4517,N_4150,N_4030);
nor U4518 (N_4518,N_4031,N_4464);
nor U4519 (N_4519,N_4191,N_4373);
and U4520 (N_4520,N_4236,N_4498);
nor U4521 (N_4521,N_4356,N_4285);
or U4522 (N_4522,N_4162,N_4005);
nor U4523 (N_4523,N_4131,N_4240);
nand U4524 (N_4524,N_4244,N_4335);
or U4525 (N_4525,N_4234,N_4345);
and U4526 (N_4526,N_4478,N_4416);
and U4527 (N_4527,N_4062,N_4289);
or U4528 (N_4528,N_4020,N_4007);
nand U4529 (N_4529,N_4209,N_4252);
or U4530 (N_4530,N_4227,N_4013);
nor U4531 (N_4531,N_4494,N_4475);
nand U4532 (N_4532,N_4155,N_4491);
or U4533 (N_4533,N_4186,N_4054);
nand U4534 (N_4534,N_4023,N_4309);
and U4535 (N_4535,N_4410,N_4071);
and U4536 (N_4536,N_4477,N_4146);
or U4537 (N_4537,N_4219,N_4393);
nor U4538 (N_4538,N_4261,N_4292);
nand U4539 (N_4539,N_4266,N_4347);
and U4540 (N_4540,N_4090,N_4431);
or U4541 (N_4541,N_4121,N_4138);
xnor U4542 (N_4542,N_4251,N_4259);
or U4543 (N_4543,N_4094,N_4056);
or U4544 (N_4544,N_4081,N_4390);
and U4545 (N_4545,N_4116,N_4492);
nor U4546 (N_4546,N_4334,N_4230);
nand U4547 (N_4547,N_4369,N_4111);
nand U4548 (N_4548,N_4398,N_4165);
nand U4549 (N_4549,N_4067,N_4057);
and U4550 (N_4550,N_4238,N_4144);
and U4551 (N_4551,N_4098,N_4350);
and U4552 (N_4552,N_4281,N_4467);
and U4553 (N_4553,N_4348,N_4117);
nand U4554 (N_4554,N_4060,N_4280);
nand U4555 (N_4555,N_4426,N_4212);
nand U4556 (N_4556,N_4106,N_4156);
nand U4557 (N_4557,N_4091,N_4453);
and U4558 (N_4558,N_4041,N_4093);
nor U4559 (N_4559,N_4151,N_4465);
nor U4560 (N_4560,N_4260,N_4339);
nor U4561 (N_4561,N_4170,N_4493);
or U4562 (N_4562,N_4387,N_4318);
or U4563 (N_4563,N_4421,N_4322);
nand U4564 (N_4564,N_4455,N_4040);
or U4565 (N_4565,N_4346,N_4193);
and U4566 (N_4566,N_4277,N_4010);
and U4567 (N_4567,N_4485,N_4408);
nor U4568 (N_4568,N_4226,N_4296);
nand U4569 (N_4569,N_4384,N_4022);
nand U4570 (N_4570,N_4396,N_4206);
nand U4571 (N_4571,N_4179,N_4037);
and U4572 (N_4572,N_4458,N_4133);
nor U4573 (N_4573,N_4305,N_4050);
nand U4574 (N_4574,N_4202,N_4084);
or U4575 (N_4575,N_4297,N_4363);
nand U4576 (N_4576,N_4269,N_4129);
nand U4577 (N_4577,N_4332,N_4446);
nor U4578 (N_4578,N_4300,N_4441);
nand U4579 (N_4579,N_4204,N_4365);
nand U4580 (N_4580,N_4069,N_4205);
nor U4581 (N_4581,N_4070,N_4237);
and U4582 (N_4582,N_4157,N_4075);
nand U4583 (N_4583,N_4409,N_4419);
and U4584 (N_4584,N_4315,N_4198);
nor U4585 (N_4585,N_4476,N_4126);
and U4586 (N_4586,N_4325,N_4239);
and U4587 (N_4587,N_4141,N_4123);
nand U4588 (N_4588,N_4233,N_4397);
nand U4589 (N_4589,N_4270,N_4189);
nand U4590 (N_4590,N_4381,N_4053);
and U4591 (N_4591,N_4473,N_4038);
nor U4592 (N_4592,N_4436,N_4044);
or U4593 (N_4593,N_4258,N_4132);
and U4594 (N_4594,N_4001,N_4454);
nor U4595 (N_4595,N_4437,N_4282);
nand U4596 (N_4596,N_4032,N_4462);
and U4597 (N_4597,N_4021,N_4364);
or U4598 (N_4598,N_4203,N_4488);
and U4599 (N_4599,N_4243,N_4166);
or U4600 (N_4600,N_4307,N_4142);
and U4601 (N_4601,N_4367,N_4174);
and U4602 (N_4602,N_4154,N_4003);
or U4603 (N_4603,N_4447,N_4048);
and U4604 (N_4604,N_4401,N_4324);
and U4605 (N_4605,N_4424,N_4482);
nor U4606 (N_4606,N_4224,N_4479);
nand U4607 (N_4607,N_4158,N_4089);
or U4608 (N_4608,N_4366,N_4480);
and U4609 (N_4609,N_4185,N_4264);
or U4610 (N_4610,N_4027,N_4374);
and U4611 (N_4611,N_4283,N_4077);
nor U4612 (N_4612,N_4086,N_4128);
and U4613 (N_4613,N_4109,N_4354);
nand U4614 (N_4614,N_4450,N_4405);
and U4615 (N_4615,N_4055,N_4026);
or U4616 (N_4616,N_4182,N_4201);
or U4617 (N_4617,N_4135,N_4388);
nand U4618 (N_4618,N_4351,N_4248);
or U4619 (N_4619,N_4349,N_4427);
nor U4620 (N_4620,N_4471,N_4034);
or U4621 (N_4621,N_4180,N_4035);
or U4622 (N_4622,N_4058,N_4461);
nand U4623 (N_4623,N_4432,N_4291);
nand U4624 (N_4624,N_4100,N_4358);
xor U4625 (N_4625,N_4370,N_4196);
nor U4626 (N_4626,N_4379,N_4148);
nand U4627 (N_4627,N_4273,N_4457);
and U4628 (N_4628,N_4046,N_4460);
and U4629 (N_4629,N_4199,N_4192);
nand U4630 (N_4630,N_4127,N_4306);
and U4631 (N_4631,N_4340,N_4456);
and U4632 (N_4632,N_4028,N_4357);
nand U4633 (N_4633,N_4006,N_4143);
or U4634 (N_4634,N_4415,N_4149);
and U4635 (N_4635,N_4112,N_4045);
xor U4636 (N_4636,N_4249,N_4009);
or U4637 (N_4637,N_4105,N_4442);
nand U4638 (N_4638,N_4378,N_4042);
nand U4639 (N_4639,N_4400,N_4072);
and U4640 (N_4640,N_4019,N_4164);
and U4641 (N_4641,N_4108,N_4463);
nand U4642 (N_4642,N_4392,N_4211);
nand U4643 (N_4643,N_4451,N_4286);
nor U4644 (N_4644,N_4320,N_4301);
or U4645 (N_4645,N_4223,N_4311);
nand U4646 (N_4646,N_4043,N_4438);
nor U4647 (N_4647,N_4484,N_4080);
nand U4648 (N_4648,N_4331,N_4122);
and U4649 (N_4649,N_4015,N_4329);
nor U4650 (N_4650,N_4172,N_4101);
nand U4651 (N_4651,N_4215,N_4294);
and U4652 (N_4652,N_4229,N_4114);
nor U4653 (N_4653,N_4130,N_4353);
and U4654 (N_4654,N_4195,N_4073);
and U4655 (N_4655,N_4420,N_4171);
or U4656 (N_4656,N_4385,N_4319);
or U4657 (N_4657,N_4496,N_4274);
nor U4658 (N_4658,N_4107,N_4217);
nor U4659 (N_4659,N_4246,N_4413);
nor U4660 (N_4660,N_4276,N_4359);
nand U4661 (N_4661,N_4220,N_4207);
or U4662 (N_4662,N_4371,N_4448);
nand U4663 (N_4663,N_4403,N_4399);
nor U4664 (N_4664,N_4472,N_4061);
or U4665 (N_4665,N_4242,N_4414);
or U4666 (N_4666,N_4103,N_4085);
nand U4667 (N_4667,N_4383,N_4235);
and U4668 (N_4668,N_4422,N_4362);
or U4669 (N_4669,N_4025,N_4299);
nand U4670 (N_4670,N_4161,N_4290);
nand U4671 (N_4671,N_4360,N_4303);
or U4672 (N_4672,N_4308,N_4167);
nor U4673 (N_4673,N_4429,N_4298);
nand U4674 (N_4674,N_4102,N_4218);
and U4675 (N_4675,N_4083,N_4160);
or U4676 (N_4676,N_4097,N_4406);
nand U4677 (N_4677,N_4068,N_4033);
and U4678 (N_4678,N_4434,N_4036);
and U4679 (N_4679,N_4216,N_4425);
and U4680 (N_4680,N_4483,N_4095);
nand U4681 (N_4681,N_4184,N_4361);
or U4682 (N_4682,N_4268,N_4272);
nor U4683 (N_4683,N_4368,N_4486);
nand U4684 (N_4684,N_4049,N_4210);
or U4685 (N_4685,N_4163,N_4323);
nand U4686 (N_4686,N_4402,N_4190);
nor U4687 (N_4687,N_4326,N_4452);
nand U4688 (N_4688,N_4417,N_4411);
xor U4689 (N_4689,N_4330,N_4262);
xnor U4690 (N_4690,N_4278,N_4440);
nand U4691 (N_4691,N_4002,N_4197);
and U4692 (N_4692,N_4016,N_4168);
and U4693 (N_4693,N_4079,N_4245);
or U4694 (N_4694,N_4257,N_4395);
xnor U4695 (N_4695,N_4372,N_4232);
or U4696 (N_4696,N_4344,N_4018);
and U4697 (N_4697,N_4275,N_4466);
and U4698 (N_4698,N_4304,N_4169);
nand U4699 (N_4699,N_4052,N_4134);
or U4700 (N_4700,N_4113,N_4208);
or U4701 (N_4701,N_4078,N_4074);
or U4702 (N_4702,N_4468,N_4221);
and U4703 (N_4703,N_4039,N_4313);
nand U4704 (N_4704,N_4213,N_4147);
or U4705 (N_4705,N_4316,N_4293);
nor U4706 (N_4706,N_4029,N_4337);
or U4707 (N_4707,N_4265,N_4183);
or U4708 (N_4708,N_4256,N_4125);
or U4709 (N_4709,N_4066,N_4051);
and U4710 (N_4710,N_4225,N_4487);
and U4711 (N_4711,N_4087,N_4469);
nor U4712 (N_4712,N_4376,N_4497);
or U4713 (N_4713,N_4333,N_4389);
and U4714 (N_4714,N_4382,N_4011);
or U4715 (N_4715,N_4014,N_4443);
nor U4716 (N_4716,N_4177,N_4489);
and U4717 (N_4717,N_4253,N_4375);
or U4718 (N_4718,N_4271,N_4490);
and U4719 (N_4719,N_4115,N_4012);
or U4720 (N_4720,N_4088,N_4152);
nand U4721 (N_4721,N_4231,N_4444);
and U4722 (N_4722,N_4140,N_4433);
or U4723 (N_4723,N_4047,N_4241);
nand U4724 (N_4724,N_4024,N_4279);
or U4725 (N_4725,N_4187,N_4470);
nor U4726 (N_4726,N_4228,N_4428);
or U4727 (N_4727,N_4386,N_4200);
and U4728 (N_4728,N_4314,N_4065);
or U4729 (N_4729,N_4247,N_4136);
or U4730 (N_4730,N_4255,N_4194);
nand U4731 (N_4731,N_4254,N_4188);
or U4732 (N_4732,N_4435,N_4495);
nand U4733 (N_4733,N_4263,N_4181);
nand U4734 (N_4734,N_4092,N_4295);
nor U4735 (N_4735,N_4076,N_4404);
and U4736 (N_4736,N_4176,N_4104);
and U4737 (N_4737,N_4412,N_4343);
nor U4738 (N_4738,N_4137,N_4008);
or U4739 (N_4739,N_4017,N_4430);
and U4740 (N_4740,N_4178,N_4336);
nand U4741 (N_4741,N_4059,N_4000);
or U4742 (N_4742,N_4338,N_4214);
nand U4743 (N_4743,N_4082,N_4449);
nor U4744 (N_4744,N_4063,N_4139);
nor U4745 (N_4745,N_4394,N_4110);
nor U4746 (N_4746,N_4175,N_4321);
nor U4747 (N_4747,N_4418,N_4004);
nor U4748 (N_4748,N_4380,N_4302);
or U4749 (N_4749,N_4099,N_4153);
nand U4750 (N_4750,N_4416,N_4193);
and U4751 (N_4751,N_4349,N_4282);
and U4752 (N_4752,N_4354,N_4108);
nand U4753 (N_4753,N_4217,N_4480);
nor U4754 (N_4754,N_4185,N_4179);
nand U4755 (N_4755,N_4205,N_4058);
or U4756 (N_4756,N_4277,N_4468);
nor U4757 (N_4757,N_4079,N_4247);
or U4758 (N_4758,N_4329,N_4448);
nand U4759 (N_4759,N_4075,N_4357);
nand U4760 (N_4760,N_4260,N_4192);
nand U4761 (N_4761,N_4309,N_4027);
nand U4762 (N_4762,N_4260,N_4217);
and U4763 (N_4763,N_4136,N_4222);
or U4764 (N_4764,N_4090,N_4168);
or U4765 (N_4765,N_4212,N_4177);
nor U4766 (N_4766,N_4339,N_4011);
nand U4767 (N_4767,N_4227,N_4170);
and U4768 (N_4768,N_4300,N_4283);
nor U4769 (N_4769,N_4428,N_4004);
nor U4770 (N_4770,N_4083,N_4062);
nor U4771 (N_4771,N_4373,N_4389);
nor U4772 (N_4772,N_4071,N_4259);
nor U4773 (N_4773,N_4436,N_4221);
nor U4774 (N_4774,N_4362,N_4084);
nor U4775 (N_4775,N_4372,N_4261);
nand U4776 (N_4776,N_4288,N_4085);
and U4777 (N_4777,N_4281,N_4452);
nand U4778 (N_4778,N_4441,N_4392);
nor U4779 (N_4779,N_4176,N_4288);
nor U4780 (N_4780,N_4328,N_4367);
or U4781 (N_4781,N_4340,N_4499);
or U4782 (N_4782,N_4062,N_4363);
nor U4783 (N_4783,N_4230,N_4364);
nor U4784 (N_4784,N_4472,N_4300);
or U4785 (N_4785,N_4014,N_4467);
and U4786 (N_4786,N_4289,N_4005);
or U4787 (N_4787,N_4390,N_4158);
nand U4788 (N_4788,N_4023,N_4077);
nand U4789 (N_4789,N_4250,N_4433);
nor U4790 (N_4790,N_4481,N_4448);
or U4791 (N_4791,N_4168,N_4178);
or U4792 (N_4792,N_4309,N_4318);
nand U4793 (N_4793,N_4043,N_4056);
or U4794 (N_4794,N_4069,N_4427);
or U4795 (N_4795,N_4089,N_4215);
nor U4796 (N_4796,N_4013,N_4298);
nor U4797 (N_4797,N_4008,N_4028);
nor U4798 (N_4798,N_4258,N_4358);
nor U4799 (N_4799,N_4012,N_4223);
nand U4800 (N_4800,N_4305,N_4240);
and U4801 (N_4801,N_4438,N_4452);
or U4802 (N_4802,N_4171,N_4270);
and U4803 (N_4803,N_4133,N_4359);
nand U4804 (N_4804,N_4454,N_4205);
nand U4805 (N_4805,N_4365,N_4463);
and U4806 (N_4806,N_4315,N_4448);
or U4807 (N_4807,N_4188,N_4056);
nand U4808 (N_4808,N_4218,N_4129);
and U4809 (N_4809,N_4107,N_4475);
and U4810 (N_4810,N_4144,N_4194);
or U4811 (N_4811,N_4223,N_4264);
or U4812 (N_4812,N_4396,N_4398);
or U4813 (N_4813,N_4073,N_4042);
or U4814 (N_4814,N_4340,N_4394);
or U4815 (N_4815,N_4280,N_4255);
xnor U4816 (N_4816,N_4035,N_4428);
or U4817 (N_4817,N_4296,N_4004);
nand U4818 (N_4818,N_4332,N_4282);
and U4819 (N_4819,N_4453,N_4141);
and U4820 (N_4820,N_4316,N_4173);
nor U4821 (N_4821,N_4220,N_4250);
and U4822 (N_4822,N_4015,N_4469);
nand U4823 (N_4823,N_4289,N_4348);
or U4824 (N_4824,N_4168,N_4325);
nor U4825 (N_4825,N_4313,N_4261);
or U4826 (N_4826,N_4446,N_4142);
nor U4827 (N_4827,N_4209,N_4148);
nand U4828 (N_4828,N_4174,N_4342);
and U4829 (N_4829,N_4413,N_4245);
or U4830 (N_4830,N_4409,N_4323);
and U4831 (N_4831,N_4074,N_4214);
and U4832 (N_4832,N_4076,N_4420);
and U4833 (N_4833,N_4221,N_4335);
nand U4834 (N_4834,N_4336,N_4452);
and U4835 (N_4835,N_4463,N_4499);
or U4836 (N_4836,N_4465,N_4453);
nand U4837 (N_4837,N_4101,N_4047);
xnor U4838 (N_4838,N_4400,N_4208);
nand U4839 (N_4839,N_4428,N_4010);
nor U4840 (N_4840,N_4450,N_4031);
nor U4841 (N_4841,N_4412,N_4128);
nand U4842 (N_4842,N_4320,N_4116);
nor U4843 (N_4843,N_4399,N_4209);
nand U4844 (N_4844,N_4057,N_4321);
nand U4845 (N_4845,N_4342,N_4134);
nand U4846 (N_4846,N_4455,N_4491);
nor U4847 (N_4847,N_4340,N_4259);
and U4848 (N_4848,N_4270,N_4095);
xor U4849 (N_4849,N_4354,N_4480);
nor U4850 (N_4850,N_4320,N_4239);
or U4851 (N_4851,N_4018,N_4140);
nand U4852 (N_4852,N_4162,N_4279);
nor U4853 (N_4853,N_4239,N_4279);
and U4854 (N_4854,N_4475,N_4496);
nor U4855 (N_4855,N_4220,N_4371);
or U4856 (N_4856,N_4431,N_4181);
and U4857 (N_4857,N_4336,N_4208);
and U4858 (N_4858,N_4186,N_4334);
nor U4859 (N_4859,N_4491,N_4310);
or U4860 (N_4860,N_4377,N_4341);
nand U4861 (N_4861,N_4039,N_4016);
nand U4862 (N_4862,N_4204,N_4074);
nand U4863 (N_4863,N_4071,N_4380);
and U4864 (N_4864,N_4378,N_4389);
nand U4865 (N_4865,N_4411,N_4192);
nor U4866 (N_4866,N_4341,N_4006);
and U4867 (N_4867,N_4278,N_4469);
and U4868 (N_4868,N_4248,N_4047);
nor U4869 (N_4869,N_4323,N_4245);
and U4870 (N_4870,N_4229,N_4293);
nor U4871 (N_4871,N_4287,N_4294);
or U4872 (N_4872,N_4467,N_4356);
and U4873 (N_4873,N_4116,N_4045);
nand U4874 (N_4874,N_4247,N_4494);
or U4875 (N_4875,N_4391,N_4306);
and U4876 (N_4876,N_4272,N_4002);
nand U4877 (N_4877,N_4465,N_4468);
nor U4878 (N_4878,N_4349,N_4398);
and U4879 (N_4879,N_4492,N_4044);
and U4880 (N_4880,N_4188,N_4360);
nor U4881 (N_4881,N_4106,N_4232);
nand U4882 (N_4882,N_4037,N_4122);
nand U4883 (N_4883,N_4170,N_4179);
nor U4884 (N_4884,N_4218,N_4317);
nand U4885 (N_4885,N_4110,N_4091);
nand U4886 (N_4886,N_4425,N_4438);
and U4887 (N_4887,N_4067,N_4189);
nand U4888 (N_4888,N_4274,N_4116);
or U4889 (N_4889,N_4324,N_4267);
nor U4890 (N_4890,N_4164,N_4163);
nor U4891 (N_4891,N_4022,N_4399);
nor U4892 (N_4892,N_4355,N_4332);
nand U4893 (N_4893,N_4004,N_4005);
nor U4894 (N_4894,N_4367,N_4289);
or U4895 (N_4895,N_4289,N_4293);
nor U4896 (N_4896,N_4216,N_4292);
nand U4897 (N_4897,N_4004,N_4446);
or U4898 (N_4898,N_4420,N_4086);
and U4899 (N_4899,N_4306,N_4080);
nor U4900 (N_4900,N_4463,N_4219);
or U4901 (N_4901,N_4200,N_4402);
and U4902 (N_4902,N_4414,N_4185);
and U4903 (N_4903,N_4474,N_4081);
nor U4904 (N_4904,N_4479,N_4447);
or U4905 (N_4905,N_4495,N_4341);
or U4906 (N_4906,N_4013,N_4041);
nor U4907 (N_4907,N_4124,N_4399);
or U4908 (N_4908,N_4088,N_4351);
or U4909 (N_4909,N_4239,N_4445);
nand U4910 (N_4910,N_4459,N_4416);
and U4911 (N_4911,N_4362,N_4312);
or U4912 (N_4912,N_4055,N_4030);
or U4913 (N_4913,N_4330,N_4212);
nor U4914 (N_4914,N_4337,N_4122);
nand U4915 (N_4915,N_4385,N_4052);
nand U4916 (N_4916,N_4480,N_4267);
and U4917 (N_4917,N_4258,N_4137);
or U4918 (N_4918,N_4384,N_4465);
and U4919 (N_4919,N_4470,N_4337);
nand U4920 (N_4920,N_4293,N_4113);
nor U4921 (N_4921,N_4023,N_4131);
nand U4922 (N_4922,N_4285,N_4074);
nor U4923 (N_4923,N_4349,N_4317);
nand U4924 (N_4924,N_4274,N_4337);
nand U4925 (N_4925,N_4195,N_4233);
or U4926 (N_4926,N_4161,N_4495);
nor U4927 (N_4927,N_4307,N_4371);
nand U4928 (N_4928,N_4395,N_4306);
and U4929 (N_4929,N_4000,N_4168);
nor U4930 (N_4930,N_4451,N_4147);
xnor U4931 (N_4931,N_4196,N_4080);
nor U4932 (N_4932,N_4283,N_4159);
or U4933 (N_4933,N_4005,N_4452);
nand U4934 (N_4934,N_4288,N_4324);
nor U4935 (N_4935,N_4429,N_4234);
xnor U4936 (N_4936,N_4057,N_4011);
nand U4937 (N_4937,N_4022,N_4018);
nand U4938 (N_4938,N_4130,N_4424);
and U4939 (N_4939,N_4481,N_4089);
nand U4940 (N_4940,N_4019,N_4139);
nand U4941 (N_4941,N_4022,N_4336);
and U4942 (N_4942,N_4287,N_4141);
and U4943 (N_4943,N_4329,N_4395);
or U4944 (N_4944,N_4369,N_4064);
or U4945 (N_4945,N_4484,N_4183);
nand U4946 (N_4946,N_4028,N_4390);
and U4947 (N_4947,N_4432,N_4256);
nand U4948 (N_4948,N_4129,N_4261);
and U4949 (N_4949,N_4070,N_4368);
nor U4950 (N_4950,N_4152,N_4465);
and U4951 (N_4951,N_4401,N_4109);
nor U4952 (N_4952,N_4390,N_4217);
xnor U4953 (N_4953,N_4225,N_4331);
nor U4954 (N_4954,N_4414,N_4234);
nand U4955 (N_4955,N_4267,N_4175);
nand U4956 (N_4956,N_4173,N_4412);
nor U4957 (N_4957,N_4325,N_4191);
nor U4958 (N_4958,N_4496,N_4399);
nand U4959 (N_4959,N_4494,N_4034);
nor U4960 (N_4960,N_4058,N_4113);
nand U4961 (N_4961,N_4307,N_4298);
or U4962 (N_4962,N_4197,N_4059);
nor U4963 (N_4963,N_4270,N_4435);
or U4964 (N_4964,N_4269,N_4367);
nand U4965 (N_4965,N_4463,N_4024);
nand U4966 (N_4966,N_4265,N_4031);
xor U4967 (N_4967,N_4068,N_4453);
nand U4968 (N_4968,N_4090,N_4372);
nand U4969 (N_4969,N_4313,N_4027);
nand U4970 (N_4970,N_4008,N_4471);
nand U4971 (N_4971,N_4277,N_4086);
nand U4972 (N_4972,N_4291,N_4475);
and U4973 (N_4973,N_4466,N_4127);
and U4974 (N_4974,N_4257,N_4466);
and U4975 (N_4975,N_4017,N_4233);
nand U4976 (N_4976,N_4142,N_4250);
nand U4977 (N_4977,N_4283,N_4169);
nor U4978 (N_4978,N_4212,N_4197);
nor U4979 (N_4979,N_4399,N_4081);
and U4980 (N_4980,N_4043,N_4009);
nand U4981 (N_4981,N_4284,N_4317);
or U4982 (N_4982,N_4474,N_4146);
nor U4983 (N_4983,N_4061,N_4412);
nand U4984 (N_4984,N_4419,N_4007);
nor U4985 (N_4985,N_4168,N_4329);
or U4986 (N_4986,N_4392,N_4413);
or U4987 (N_4987,N_4194,N_4152);
nor U4988 (N_4988,N_4072,N_4301);
or U4989 (N_4989,N_4291,N_4292);
nor U4990 (N_4990,N_4039,N_4203);
or U4991 (N_4991,N_4302,N_4386);
and U4992 (N_4992,N_4431,N_4019);
nor U4993 (N_4993,N_4329,N_4301);
or U4994 (N_4994,N_4210,N_4372);
or U4995 (N_4995,N_4450,N_4442);
nor U4996 (N_4996,N_4295,N_4249);
and U4997 (N_4997,N_4252,N_4463);
or U4998 (N_4998,N_4268,N_4285);
nand U4999 (N_4999,N_4494,N_4022);
or U5000 (N_5000,N_4781,N_4703);
and U5001 (N_5001,N_4675,N_4667);
nor U5002 (N_5002,N_4830,N_4638);
and U5003 (N_5003,N_4714,N_4681);
nor U5004 (N_5004,N_4945,N_4741);
nor U5005 (N_5005,N_4580,N_4615);
and U5006 (N_5006,N_4548,N_4785);
or U5007 (N_5007,N_4616,N_4712);
nor U5008 (N_5008,N_4822,N_4550);
and U5009 (N_5009,N_4860,N_4735);
nor U5010 (N_5010,N_4931,N_4811);
and U5011 (N_5011,N_4632,N_4976);
xnor U5012 (N_5012,N_4956,N_4977);
nand U5013 (N_5013,N_4801,N_4889);
and U5014 (N_5014,N_4769,N_4588);
nor U5015 (N_5015,N_4509,N_4697);
nor U5016 (N_5016,N_4579,N_4888);
nor U5017 (N_5017,N_4549,N_4890);
nor U5018 (N_5018,N_4951,N_4870);
nand U5019 (N_5019,N_4850,N_4963);
nor U5020 (N_5020,N_4983,N_4605);
and U5021 (N_5021,N_4794,N_4671);
and U5022 (N_5022,N_4940,N_4919);
nand U5023 (N_5023,N_4784,N_4522);
or U5024 (N_5024,N_4751,N_4920);
nand U5025 (N_5025,N_4943,N_4901);
or U5026 (N_5026,N_4770,N_4904);
nand U5027 (N_5027,N_4907,N_4746);
nand U5028 (N_5028,N_4601,N_4718);
nand U5029 (N_5029,N_4578,N_4937);
and U5030 (N_5030,N_4866,N_4762);
nor U5031 (N_5031,N_4629,N_4849);
nor U5032 (N_5032,N_4600,N_4665);
nor U5033 (N_5033,N_4627,N_4926);
and U5034 (N_5034,N_4955,N_4704);
and U5035 (N_5035,N_4753,N_4898);
or U5036 (N_5036,N_4755,N_4599);
or U5037 (N_5037,N_4587,N_4541);
nand U5038 (N_5038,N_4612,N_4530);
or U5039 (N_5039,N_4613,N_4899);
and U5040 (N_5040,N_4756,N_4607);
and U5041 (N_5041,N_4654,N_4879);
nor U5042 (N_5042,N_4859,N_4772);
and U5043 (N_5043,N_4992,N_4805);
xor U5044 (N_5044,N_4643,N_4909);
nor U5045 (N_5045,N_4817,N_4854);
xor U5046 (N_5046,N_4614,N_4572);
and U5047 (N_5047,N_4574,N_4930);
and U5048 (N_5048,N_4964,N_4668);
nor U5049 (N_5049,N_4651,N_4840);
and U5050 (N_5050,N_4711,N_4551);
or U5051 (N_5051,N_4846,N_4820);
and U5052 (N_5052,N_4745,N_4744);
or U5053 (N_5053,N_4984,N_4799);
nor U5054 (N_5054,N_4670,N_4981);
nor U5055 (N_5055,N_4793,N_4912);
nor U5056 (N_5056,N_4944,N_4825);
and U5057 (N_5057,N_4748,N_4506);
nand U5058 (N_5058,N_4764,N_4637);
xor U5059 (N_5059,N_4639,N_4502);
or U5060 (N_5060,N_4826,N_4812);
nand U5061 (N_5061,N_4916,N_4832);
nor U5062 (N_5062,N_4966,N_4887);
nor U5063 (N_5063,N_4842,N_4581);
or U5064 (N_5064,N_4729,N_4526);
or U5065 (N_5065,N_4570,N_4975);
nand U5066 (N_5066,N_4518,N_4710);
nand U5067 (N_5067,N_4921,N_4693);
nand U5068 (N_5068,N_4686,N_4852);
or U5069 (N_5069,N_4653,N_4941);
and U5070 (N_5070,N_4758,N_4611);
nand U5071 (N_5071,N_4517,N_4935);
nand U5072 (N_5072,N_4939,N_4732);
or U5073 (N_5073,N_4584,N_4824);
and U5074 (N_5074,N_4942,N_4938);
nand U5075 (N_5075,N_4573,N_4989);
and U5076 (N_5076,N_4750,N_4682);
nor U5077 (N_5077,N_4836,N_4819);
or U5078 (N_5078,N_4680,N_4695);
and U5079 (N_5079,N_4647,N_4903);
or U5080 (N_5080,N_4765,N_4521);
and U5081 (N_5081,N_4527,N_4532);
or U5082 (N_5082,N_4576,N_4594);
or U5083 (N_5083,N_4933,N_4771);
nor U5084 (N_5084,N_4757,N_4617);
nand U5085 (N_5085,N_4848,N_4782);
and U5086 (N_5086,N_4650,N_4915);
and U5087 (N_5087,N_4731,N_4910);
nand U5088 (N_5088,N_4661,N_4664);
or U5089 (N_5089,N_4813,N_4561);
or U5090 (N_5090,N_4577,N_4766);
nor U5091 (N_5091,N_4698,N_4768);
nand U5092 (N_5092,N_4923,N_4918);
or U5093 (N_5093,N_4878,N_4928);
nand U5094 (N_5094,N_4986,N_4980);
or U5095 (N_5095,N_4531,N_4917);
nand U5096 (N_5096,N_4761,N_4990);
nor U5097 (N_5097,N_4666,N_4863);
nor U5098 (N_5098,N_4971,N_4677);
nor U5099 (N_5099,N_4688,N_4564);
and U5100 (N_5100,N_4857,N_4610);
nand U5101 (N_5101,N_4702,N_4511);
nand U5102 (N_5102,N_4501,N_4586);
and U5103 (N_5103,N_4893,N_4875);
and U5104 (N_5104,N_4823,N_4707);
nand U5105 (N_5105,N_4960,N_4592);
nand U5106 (N_5106,N_4700,N_4998);
nor U5107 (N_5107,N_4519,N_4958);
nand U5108 (N_5108,N_4692,N_4589);
nand U5109 (N_5109,N_4829,N_4914);
and U5110 (N_5110,N_4649,N_4835);
nor U5111 (N_5111,N_4721,N_4690);
xor U5112 (N_5112,N_4776,N_4885);
or U5113 (N_5113,N_4747,N_4795);
or U5114 (N_5114,N_4591,N_4708);
nand U5115 (N_5115,N_4683,N_4804);
nor U5116 (N_5116,N_4808,N_4728);
or U5117 (N_5117,N_4540,N_4725);
nand U5118 (N_5118,N_4537,N_4634);
or U5119 (N_5119,N_4557,N_4678);
nor U5120 (N_5120,N_4618,N_4694);
nor U5121 (N_5121,N_4554,N_4622);
nor U5122 (N_5122,N_4839,N_4743);
nor U5123 (N_5123,N_4844,N_4886);
nor U5124 (N_5124,N_4936,N_4633);
nor U5125 (N_5125,N_4630,N_4779);
or U5126 (N_5126,N_4985,N_4544);
nand U5127 (N_5127,N_4927,N_4696);
or U5128 (N_5128,N_4512,N_4645);
nand U5129 (N_5129,N_4833,N_4775);
and U5130 (N_5130,N_4628,N_4952);
or U5131 (N_5131,N_4996,N_4626);
or U5132 (N_5132,N_4507,N_4736);
and U5133 (N_5133,N_4896,N_4891);
or U5134 (N_5134,N_4814,N_4773);
nor U5135 (N_5135,N_4837,N_4834);
nor U5136 (N_5136,N_4767,N_4528);
nand U5137 (N_5137,N_4954,N_4566);
nand U5138 (N_5138,N_4991,N_4596);
nand U5139 (N_5139,N_4536,N_4913);
xor U5140 (N_5140,N_4806,N_4500);
and U5141 (N_5141,N_4624,N_4724);
nor U5142 (N_5142,N_4979,N_4906);
nor U5143 (N_5143,N_4734,N_4783);
and U5144 (N_5144,N_4908,N_4778);
nand U5145 (N_5145,N_4974,N_4603);
nand U5146 (N_5146,N_4663,N_4529);
and U5147 (N_5147,N_4791,N_4961);
nand U5148 (N_5148,N_4669,N_4740);
nor U5149 (N_5149,N_4546,N_4925);
and U5150 (N_5150,N_4993,N_4625);
nand U5151 (N_5151,N_4789,N_4569);
and U5152 (N_5152,N_4623,N_4602);
nor U5153 (N_5153,N_4988,N_4777);
nor U5154 (N_5154,N_4872,N_4962);
nor U5155 (N_5155,N_4585,N_4797);
nand U5156 (N_5156,N_4520,N_4523);
nor U5157 (N_5157,N_4553,N_4534);
and U5158 (N_5158,N_4709,N_4982);
or U5159 (N_5159,N_4796,N_4994);
or U5160 (N_5160,N_4722,N_4843);
and U5161 (N_5161,N_4723,N_4867);
and U5162 (N_5162,N_4593,N_4987);
nand U5163 (N_5163,N_4621,N_4868);
nor U5164 (N_5164,N_4881,N_4567);
nand U5165 (N_5165,N_4552,N_4590);
and U5166 (N_5166,N_4788,N_4905);
and U5167 (N_5167,N_4516,N_4687);
and U5168 (N_5168,N_4774,N_4949);
nand U5169 (N_5169,N_4539,N_4815);
and U5170 (N_5170,N_4871,N_4877);
nand U5171 (N_5171,N_4582,N_4884);
nand U5172 (N_5172,N_4543,N_4749);
or U5173 (N_5173,N_4575,N_4809);
and U5174 (N_5174,N_4672,N_4947);
nor U5175 (N_5175,N_4970,N_4929);
nor U5176 (N_5176,N_4999,N_4831);
nor U5177 (N_5177,N_4882,N_4739);
nor U5178 (N_5178,N_4715,N_4642);
or U5179 (N_5179,N_4864,N_4513);
or U5180 (N_5180,N_4595,N_4571);
nand U5181 (N_5181,N_4760,N_4763);
and U5182 (N_5182,N_4851,N_4644);
nand U5183 (N_5183,N_4894,N_4604);
nor U5184 (N_5184,N_4897,N_4717);
nor U5185 (N_5185,N_4946,N_4685);
nand U5186 (N_5186,N_4953,N_4560);
nor U5187 (N_5187,N_4895,N_4619);
nand U5188 (N_5188,N_4883,N_4847);
nor U5189 (N_5189,N_4597,N_4656);
nand U5190 (N_5190,N_4995,N_4738);
and U5191 (N_5191,N_4856,N_4606);
nand U5192 (N_5192,N_4706,N_4841);
or U5193 (N_5193,N_4558,N_4759);
nand U5194 (N_5194,N_4900,N_4807);
or U5195 (N_5195,N_4800,N_4858);
or U5196 (N_5196,N_4620,N_4533);
nor U5197 (N_5197,N_4640,N_4701);
nor U5198 (N_5198,N_4655,N_4828);
nor U5199 (N_5199,N_4659,N_4810);
and U5200 (N_5200,N_4737,N_4978);
and U5201 (N_5201,N_4934,N_4865);
nor U5202 (N_5202,N_4657,N_4818);
and U5203 (N_5203,N_4730,N_4827);
xnor U5204 (N_5204,N_4733,N_4727);
and U5205 (N_5205,N_4515,N_4699);
nor U5206 (N_5206,N_4631,N_4679);
nor U5207 (N_5207,N_4816,N_4742);
nor U5208 (N_5208,N_4514,N_4563);
and U5209 (N_5209,N_4562,N_4922);
and U5210 (N_5210,N_4924,N_4950);
and U5211 (N_5211,N_4689,N_4713);
nand U5212 (N_5212,N_4787,N_4691);
or U5213 (N_5213,N_4880,N_4948);
or U5214 (N_5214,N_4786,N_4973);
or U5215 (N_5215,N_4646,N_4969);
nor U5216 (N_5216,N_4608,N_4684);
nor U5217 (N_5217,N_4803,N_4641);
or U5218 (N_5218,N_4853,N_4568);
or U5219 (N_5219,N_4892,N_4673);
nor U5220 (N_5220,N_4676,N_4821);
and U5221 (N_5221,N_4932,N_4648);
or U5222 (N_5222,N_4752,N_4780);
or U5223 (N_5223,N_4662,N_4911);
or U5224 (N_5224,N_4583,N_4705);
nand U5225 (N_5225,N_4635,N_4720);
nor U5226 (N_5226,N_4542,N_4674);
or U5227 (N_5227,N_4658,N_4802);
xnor U5228 (N_5228,N_4598,N_4510);
nand U5229 (N_5229,N_4556,N_4545);
and U5230 (N_5230,N_4790,N_4716);
nor U5231 (N_5231,N_4524,N_4869);
nand U5232 (N_5232,N_4959,N_4874);
or U5233 (N_5233,N_4862,N_4972);
and U5234 (N_5234,N_4876,N_4547);
nor U5235 (N_5235,N_4968,N_4838);
or U5236 (N_5236,N_4535,N_4861);
or U5237 (N_5237,N_4726,N_4902);
and U5238 (N_5238,N_4525,N_4505);
nor U5239 (N_5239,N_4855,N_4660);
or U5240 (N_5240,N_4965,N_4538);
nor U5241 (N_5241,N_4957,N_4845);
nand U5242 (N_5242,N_4967,N_4559);
and U5243 (N_5243,N_4555,N_4719);
nor U5244 (N_5244,N_4565,N_4504);
nor U5245 (N_5245,N_4798,N_4503);
nand U5246 (N_5246,N_4792,N_4997);
or U5247 (N_5247,N_4873,N_4508);
and U5248 (N_5248,N_4609,N_4636);
or U5249 (N_5249,N_4754,N_4652);
and U5250 (N_5250,N_4875,N_4559);
and U5251 (N_5251,N_4513,N_4598);
and U5252 (N_5252,N_4501,N_4905);
or U5253 (N_5253,N_4564,N_4660);
nor U5254 (N_5254,N_4839,N_4602);
nand U5255 (N_5255,N_4529,N_4933);
nor U5256 (N_5256,N_4536,N_4789);
and U5257 (N_5257,N_4531,N_4568);
nor U5258 (N_5258,N_4753,N_4940);
or U5259 (N_5259,N_4599,N_4584);
and U5260 (N_5260,N_4828,N_4917);
or U5261 (N_5261,N_4501,N_4530);
nand U5262 (N_5262,N_4655,N_4561);
nand U5263 (N_5263,N_4619,N_4965);
or U5264 (N_5264,N_4840,N_4919);
nand U5265 (N_5265,N_4958,N_4798);
or U5266 (N_5266,N_4825,N_4981);
and U5267 (N_5267,N_4825,N_4632);
or U5268 (N_5268,N_4516,N_4848);
and U5269 (N_5269,N_4535,N_4594);
nor U5270 (N_5270,N_4672,N_4700);
nor U5271 (N_5271,N_4663,N_4949);
nand U5272 (N_5272,N_4521,N_4592);
or U5273 (N_5273,N_4594,N_4541);
nand U5274 (N_5274,N_4551,N_4540);
and U5275 (N_5275,N_4841,N_4835);
and U5276 (N_5276,N_4570,N_4923);
and U5277 (N_5277,N_4788,N_4965);
nand U5278 (N_5278,N_4631,N_4725);
nor U5279 (N_5279,N_4942,N_4882);
and U5280 (N_5280,N_4795,N_4529);
and U5281 (N_5281,N_4675,N_4833);
or U5282 (N_5282,N_4711,N_4619);
and U5283 (N_5283,N_4909,N_4732);
nand U5284 (N_5284,N_4620,N_4896);
nor U5285 (N_5285,N_4904,N_4817);
nand U5286 (N_5286,N_4785,N_4992);
or U5287 (N_5287,N_4587,N_4969);
and U5288 (N_5288,N_4944,N_4990);
or U5289 (N_5289,N_4674,N_4565);
nand U5290 (N_5290,N_4963,N_4739);
nor U5291 (N_5291,N_4817,N_4881);
nor U5292 (N_5292,N_4776,N_4832);
and U5293 (N_5293,N_4550,N_4959);
or U5294 (N_5294,N_4916,N_4953);
nand U5295 (N_5295,N_4726,N_4528);
nor U5296 (N_5296,N_4551,N_4741);
and U5297 (N_5297,N_4917,N_4856);
nor U5298 (N_5298,N_4543,N_4776);
and U5299 (N_5299,N_4829,N_4639);
and U5300 (N_5300,N_4609,N_4785);
nand U5301 (N_5301,N_4970,N_4723);
nor U5302 (N_5302,N_4972,N_4671);
or U5303 (N_5303,N_4957,N_4532);
nand U5304 (N_5304,N_4773,N_4647);
or U5305 (N_5305,N_4821,N_4707);
nand U5306 (N_5306,N_4944,N_4646);
or U5307 (N_5307,N_4628,N_4709);
nand U5308 (N_5308,N_4896,N_4503);
and U5309 (N_5309,N_4772,N_4700);
or U5310 (N_5310,N_4603,N_4923);
and U5311 (N_5311,N_4934,N_4668);
and U5312 (N_5312,N_4861,N_4772);
nor U5313 (N_5313,N_4793,N_4635);
nand U5314 (N_5314,N_4969,N_4655);
or U5315 (N_5315,N_4657,N_4794);
and U5316 (N_5316,N_4540,N_4522);
xnor U5317 (N_5317,N_4973,N_4891);
nand U5318 (N_5318,N_4718,N_4912);
nand U5319 (N_5319,N_4703,N_4884);
and U5320 (N_5320,N_4994,N_4583);
and U5321 (N_5321,N_4755,N_4533);
nand U5322 (N_5322,N_4697,N_4600);
and U5323 (N_5323,N_4609,N_4835);
nor U5324 (N_5324,N_4981,N_4563);
nand U5325 (N_5325,N_4915,N_4884);
or U5326 (N_5326,N_4662,N_4626);
nand U5327 (N_5327,N_4924,N_4942);
nand U5328 (N_5328,N_4578,N_4579);
nand U5329 (N_5329,N_4803,N_4584);
xor U5330 (N_5330,N_4988,N_4706);
nor U5331 (N_5331,N_4798,N_4764);
nand U5332 (N_5332,N_4716,N_4855);
nand U5333 (N_5333,N_4665,N_4953);
nand U5334 (N_5334,N_4798,N_4846);
and U5335 (N_5335,N_4542,N_4950);
nand U5336 (N_5336,N_4564,N_4664);
nor U5337 (N_5337,N_4940,N_4774);
nor U5338 (N_5338,N_4579,N_4939);
and U5339 (N_5339,N_4633,N_4850);
nand U5340 (N_5340,N_4703,N_4911);
nor U5341 (N_5341,N_4511,N_4943);
nor U5342 (N_5342,N_4710,N_4926);
nand U5343 (N_5343,N_4770,N_4660);
and U5344 (N_5344,N_4556,N_4535);
and U5345 (N_5345,N_4957,N_4808);
and U5346 (N_5346,N_4528,N_4837);
or U5347 (N_5347,N_4787,N_4920);
and U5348 (N_5348,N_4780,N_4647);
nor U5349 (N_5349,N_4916,N_4962);
and U5350 (N_5350,N_4851,N_4836);
xnor U5351 (N_5351,N_4796,N_4728);
or U5352 (N_5352,N_4890,N_4956);
or U5353 (N_5353,N_4520,N_4857);
nor U5354 (N_5354,N_4731,N_4939);
nand U5355 (N_5355,N_4672,N_4655);
nand U5356 (N_5356,N_4665,N_4685);
nor U5357 (N_5357,N_4573,N_4859);
nor U5358 (N_5358,N_4814,N_4792);
nand U5359 (N_5359,N_4702,N_4816);
and U5360 (N_5360,N_4730,N_4879);
nand U5361 (N_5361,N_4539,N_4564);
and U5362 (N_5362,N_4653,N_4800);
nand U5363 (N_5363,N_4734,N_4916);
nand U5364 (N_5364,N_4647,N_4931);
nor U5365 (N_5365,N_4500,N_4856);
nand U5366 (N_5366,N_4589,N_4964);
or U5367 (N_5367,N_4768,N_4839);
and U5368 (N_5368,N_4727,N_4865);
xnor U5369 (N_5369,N_4610,N_4939);
nor U5370 (N_5370,N_4964,N_4735);
or U5371 (N_5371,N_4575,N_4981);
nand U5372 (N_5372,N_4630,N_4647);
nor U5373 (N_5373,N_4610,N_4816);
nor U5374 (N_5374,N_4691,N_4879);
xnor U5375 (N_5375,N_4892,N_4879);
or U5376 (N_5376,N_4969,N_4840);
nand U5377 (N_5377,N_4718,N_4898);
and U5378 (N_5378,N_4789,N_4509);
or U5379 (N_5379,N_4871,N_4905);
nor U5380 (N_5380,N_4865,N_4660);
nand U5381 (N_5381,N_4899,N_4837);
nor U5382 (N_5382,N_4777,N_4549);
nand U5383 (N_5383,N_4722,N_4829);
nor U5384 (N_5384,N_4844,N_4900);
nand U5385 (N_5385,N_4706,N_4945);
or U5386 (N_5386,N_4949,N_4976);
nand U5387 (N_5387,N_4565,N_4677);
and U5388 (N_5388,N_4684,N_4744);
nor U5389 (N_5389,N_4619,N_4613);
and U5390 (N_5390,N_4610,N_4593);
nand U5391 (N_5391,N_4528,N_4576);
nand U5392 (N_5392,N_4790,N_4769);
and U5393 (N_5393,N_4661,N_4762);
and U5394 (N_5394,N_4948,N_4647);
and U5395 (N_5395,N_4743,N_4577);
or U5396 (N_5396,N_4524,N_4823);
and U5397 (N_5397,N_4793,N_4751);
nand U5398 (N_5398,N_4732,N_4828);
nand U5399 (N_5399,N_4887,N_4794);
or U5400 (N_5400,N_4643,N_4670);
nand U5401 (N_5401,N_4733,N_4618);
or U5402 (N_5402,N_4569,N_4549);
nand U5403 (N_5403,N_4986,N_4535);
nor U5404 (N_5404,N_4717,N_4957);
nor U5405 (N_5405,N_4660,N_4609);
and U5406 (N_5406,N_4690,N_4545);
nand U5407 (N_5407,N_4820,N_4758);
and U5408 (N_5408,N_4666,N_4707);
xnor U5409 (N_5409,N_4758,N_4789);
and U5410 (N_5410,N_4787,N_4813);
or U5411 (N_5411,N_4596,N_4912);
nor U5412 (N_5412,N_4746,N_4648);
nor U5413 (N_5413,N_4635,N_4554);
nor U5414 (N_5414,N_4959,N_4793);
and U5415 (N_5415,N_4764,N_4742);
and U5416 (N_5416,N_4540,N_4817);
and U5417 (N_5417,N_4750,N_4690);
nand U5418 (N_5418,N_4740,N_4606);
nor U5419 (N_5419,N_4602,N_4857);
nand U5420 (N_5420,N_4883,N_4653);
nand U5421 (N_5421,N_4663,N_4756);
and U5422 (N_5422,N_4895,N_4788);
nand U5423 (N_5423,N_4978,N_4816);
xor U5424 (N_5424,N_4841,N_4845);
nor U5425 (N_5425,N_4653,N_4989);
and U5426 (N_5426,N_4614,N_4503);
and U5427 (N_5427,N_4789,N_4801);
nand U5428 (N_5428,N_4532,N_4969);
and U5429 (N_5429,N_4723,N_4562);
or U5430 (N_5430,N_4866,N_4505);
and U5431 (N_5431,N_4606,N_4761);
or U5432 (N_5432,N_4891,N_4924);
nor U5433 (N_5433,N_4926,N_4633);
or U5434 (N_5434,N_4615,N_4572);
nor U5435 (N_5435,N_4594,N_4880);
and U5436 (N_5436,N_4972,N_4760);
nor U5437 (N_5437,N_4569,N_4522);
nor U5438 (N_5438,N_4843,N_4697);
and U5439 (N_5439,N_4542,N_4993);
or U5440 (N_5440,N_4892,N_4987);
or U5441 (N_5441,N_4500,N_4758);
and U5442 (N_5442,N_4616,N_4564);
or U5443 (N_5443,N_4943,N_4716);
or U5444 (N_5444,N_4537,N_4585);
nand U5445 (N_5445,N_4815,N_4728);
nor U5446 (N_5446,N_4691,N_4535);
nand U5447 (N_5447,N_4996,N_4654);
xor U5448 (N_5448,N_4639,N_4987);
or U5449 (N_5449,N_4675,N_4565);
or U5450 (N_5450,N_4579,N_4897);
xor U5451 (N_5451,N_4998,N_4900);
or U5452 (N_5452,N_4785,N_4789);
or U5453 (N_5453,N_4675,N_4772);
nand U5454 (N_5454,N_4877,N_4506);
nor U5455 (N_5455,N_4678,N_4649);
xnor U5456 (N_5456,N_4733,N_4689);
and U5457 (N_5457,N_4884,N_4726);
nor U5458 (N_5458,N_4783,N_4665);
or U5459 (N_5459,N_4797,N_4629);
nand U5460 (N_5460,N_4638,N_4588);
nand U5461 (N_5461,N_4869,N_4550);
nor U5462 (N_5462,N_4829,N_4526);
nor U5463 (N_5463,N_4844,N_4550);
and U5464 (N_5464,N_4889,N_4623);
and U5465 (N_5465,N_4631,N_4954);
and U5466 (N_5466,N_4965,N_4903);
or U5467 (N_5467,N_4718,N_4738);
nor U5468 (N_5468,N_4743,N_4993);
nand U5469 (N_5469,N_4838,N_4952);
nand U5470 (N_5470,N_4515,N_4967);
nand U5471 (N_5471,N_4647,N_4853);
or U5472 (N_5472,N_4695,N_4640);
nor U5473 (N_5473,N_4859,N_4568);
or U5474 (N_5474,N_4811,N_4585);
nor U5475 (N_5475,N_4979,N_4529);
and U5476 (N_5476,N_4790,N_4973);
or U5477 (N_5477,N_4583,N_4501);
nand U5478 (N_5478,N_4512,N_4960);
and U5479 (N_5479,N_4941,N_4600);
nand U5480 (N_5480,N_4976,N_4757);
xnor U5481 (N_5481,N_4815,N_4994);
nand U5482 (N_5482,N_4608,N_4923);
or U5483 (N_5483,N_4919,N_4538);
nor U5484 (N_5484,N_4942,N_4937);
nand U5485 (N_5485,N_4851,N_4991);
nand U5486 (N_5486,N_4685,N_4812);
nor U5487 (N_5487,N_4950,N_4815);
nor U5488 (N_5488,N_4672,N_4527);
nand U5489 (N_5489,N_4699,N_4620);
nor U5490 (N_5490,N_4506,N_4935);
nor U5491 (N_5491,N_4621,N_4641);
nor U5492 (N_5492,N_4952,N_4650);
nand U5493 (N_5493,N_4518,N_4920);
xor U5494 (N_5494,N_4579,N_4925);
and U5495 (N_5495,N_4810,N_4980);
and U5496 (N_5496,N_4584,N_4973);
and U5497 (N_5497,N_4655,N_4596);
and U5498 (N_5498,N_4981,N_4763);
and U5499 (N_5499,N_4783,N_4884);
nand U5500 (N_5500,N_5008,N_5270);
nand U5501 (N_5501,N_5108,N_5486);
or U5502 (N_5502,N_5407,N_5284);
nand U5503 (N_5503,N_5152,N_5352);
nor U5504 (N_5504,N_5368,N_5230);
and U5505 (N_5505,N_5034,N_5366);
or U5506 (N_5506,N_5421,N_5318);
nand U5507 (N_5507,N_5112,N_5350);
nor U5508 (N_5508,N_5335,N_5315);
and U5509 (N_5509,N_5290,N_5195);
or U5510 (N_5510,N_5193,N_5356);
nor U5511 (N_5511,N_5236,N_5477);
and U5512 (N_5512,N_5492,N_5169);
nor U5513 (N_5513,N_5093,N_5484);
nor U5514 (N_5514,N_5226,N_5158);
nor U5515 (N_5515,N_5105,N_5104);
nor U5516 (N_5516,N_5050,N_5085);
or U5517 (N_5517,N_5190,N_5205);
nor U5518 (N_5518,N_5417,N_5045);
nor U5519 (N_5519,N_5041,N_5082);
or U5520 (N_5520,N_5182,N_5410);
nor U5521 (N_5521,N_5124,N_5151);
or U5522 (N_5522,N_5208,N_5072);
and U5523 (N_5523,N_5483,N_5365);
or U5524 (N_5524,N_5061,N_5478);
and U5525 (N_5525,N_5038,N_5126);
and U5526 (N_5526,N_5420,N_5273);
and U5527 (N_5527,N_5428,N_5456);
and U5528 (N_5528,N_5431,N_5363);
and U5529 (N_5529,N_5166,N_5458);
or U5530 (N_5530,N_5001,N_5187);
nand U5531 (N_5531,N_5327,N_5445);
nand U5532 (N_5532,N_5090,N_5324);
nand U5533 (N_5533,N_5340,N_5252);
nor U5534 (N_5534,N_5444,N_5238);
or U5535 (N_5535,N_5092,N_5348);
or U5536 (N_5536,N_5218,N_5170);
or U5537 (N_5537,N_5387,N_5223);
or U5538 (N_5538,N_5308,N_5261);
or U5539 (N_5539,N_5217,N_5455);
or U5540 (N_5540,N_5286,N_5495);
or U5541 (N_5541,N_5010,N_5224);
or U5542 (N_5542,N_5147,N_5254);
nor U5543 (N_5543,N_5059,N_5405);
nand U5544 (N_5544,N_5314,N_5459);
nor U5545 (N_5545,N_5438,N_5080);
nand U5546 (N_5546,N_5115,N_5349);
or U5547 (N_5547,N_5296,N_5198);
nor U5548 (N_5548,N_5457,N_5344);
nand U5549 (N_5549,N_5269,N_5194);
nor U5550 (N_5550,N_5278,N_5109);
xor U5551 (N_5551,N_5019,N_5003);
or U5552 (N_5552,N_5282,N_5036);
nor U5553 (N_5553,N_5196,N_5075);
nor U5554 (N_5554,N_5331,N_5334);
nand U5555 (N_5555,N_5339,N_5107);
nand U5556 (N_5556,N_5361,N_5087);
nor U5557 (N_5557,N_5135,N_5371);
nor U5558 (N_5558,N_5227,N_5362);
nand U5559 (N_5559,N_5077,N_5121);
nor U5560 (N_5560,N_5244,N_5174);
and U5561 (N_5561,N_5228,N_5251);
or U5562 (N_5562,N_5162,N_5346);
or U5563 (N_5563,N_5088,N_5225);
nand U5564 (N_5564,N_5246,N_5298);
and U5565 (N_5565,N_5118,N_5436);
nor U5566 (N_5566,N_5289,N_5337);
and U5567 (N_5567,N_5063,N_5475);
nor U5568 (N_5568,N_5330,N_5117);
or U5569 (N_5569,N_5027,N_5023);
nand U5570 (N_5570,N_5233,N_5111);
nand U5571 (N_5571,N_5497,N_5287);
or U5572 (N_5572,N_5207,N_5048);
nor U5573 (N_5573,N_5219,N_5091);
and U5574 (N_5574,N_5496,N_5142);
nor U5575 (N_5575,N_5398,N_5262);
nor U5576 (N_5576,N_5221,N_5370);
nand U5577 (N_5577,N_5018,N_5393);
nor U5578 (N_5578,N_5402,N_5099);
nor U5579 (N_5579,N_5442,N_5447);
nor U5580 (N_5580,N_5413,N_5345);
nor U5581 (N_5581,N_5053,N_5357);
or U5582 (N_5582,N_5411,N_5000);
nand U5583 (N_5583,N_5199,N_5317);
nor U5584 (N_5584,N_5248,N_5129);
or U5585 (N_5585,N_5429,N_5030);
nand U5586 (N_5586,N_5240,N_5395);
or U5587 (N_5587,N_5209,N_5028);
nand U5588 (N_5588,N_5245,N_5042);
nand U5589 (N_5589,N_5434,N_5202);
nor U5590 (N_5590,N_5016,N_5277);
nor U5591 (N_5591,N_5263,N_5266);
nand U5592 (N_5592,N_5376,N_5412);
nor U5593 (N_5593,N_5253,N_5372);
and U5594 (N_5594,N_5177,N_5322);
and U5595 (N_5595,N_5103,N_5106);
and U5596 (N_5596,N_5178,N_5168);
nand U5597 (N_5597,N_5403,N_5157);
nor U5598 (N_5598,N_5443,N_5423);
nand U5599 (N_5599,N_5267,N_5414);
or U5600 (N_5600,N_5123,N_5154);
nor U5601 (N_5601,N_5052,N_5250);
or U5602 (N_5602,N_5096,N_5100);
nand U5603 (N_5603,N_5389,N_5325);
nand U5604 (N_5604,N_5037,N_5153);
nor U5605 (N_5605,N_5453,N_5229);
and U5606 (N_5606,N_5408,N_5285);
nand U5607 (N_5607,N_5264,N_5144);
and U5608 (N_5608,N_5451,N_5448);
nor U5609 (N_5609,N_5125,N_5441);
nand U5610 (N_5610,N_5243,N_5119);
nand U5611 (N_5611,N_5164,N_5313);
nand U5612 (N_5612,N_5300,N_5424);
and U5613 (N_5613,N_5463,N_5399);
nor U5614 (N_5614,N_5382,N_5247);
and U5615 (N_5615,N_5347,N_5396);
xor U5616 (N_5616,N_5401,N_5294);
and U5617 (N_5617,N_5473,N_5392);
and U5618 (N_5618,N_5148,N_5131);
nor U5619 (N_5619,N_5046,N_5328);
or U5620 (N_5620,N_5304,N_5481);
or U5621 (N_5621,N_5415,N_5005);
xnor U5622 (N_5622,N_5241,N_5498);
nor U5623 (N_5623,N_5472,N_5394);
or U5624 (N_5624,N_5275,N_5406);
nor U5625 (N_5625,N_5029,N_5427);
nand U5626 (N_5626,N_5215,N_5189);
nand U5627 (N_5627,N_5409,N_5114);
nor U5628 (N_5628,N_5465,N_5332);
or U5629 (N_5629,N_5200,N_5291);
nand U5630 (N_5630,N_5310,N_5171);
and U5631 (N_5631,N_5102,N_5165);
or U5632 (N_5632,N_5012,N_5388);
nor U5633 (N_5633,N_5487,N_5064);
nand U5634 (N_5634,N_5272,N_5184);
and U5635 (N_5635,N_5358,N_5482);
nor U5636 (N_5636,N_5035,N_5074);
and U5637 (N_5637,N_5128,N_5307);
or U5638 (N_5638,N_5049,N_5137);
nand U5639 (N_5639,N_5302,N_5316);
and U5640 (N_5640,N_5133,N_5094);
nor U5641 (N_5641,N_5450,N_5078);
nand U5642 (N_5642,N_5303,N_5425);
and U5643 (N_5643,N_5089,N_5116);
nor U5644 (N_5644,N_5130,N_5391);
and U5645 (N_5645,N_5081,N_5161);
nor U5646 (N_5646,N_5020,N_5257);
nand U5647 (N_5647,N_5134,N_5343);
or U5648 (N_5648,N_5186,N_5295);
or U5649 (N_5649,N_5281,N_5222);
nor U5650 (N_5650,N_5462,N_5390);
nor U5651 (N_5651,N_5176,N_5268);
or U5652 (N_5652,N_5360,N_5172);
nor U5653 (N_5653,N_5426,N_5054);
nor U5654 (N_5654,N_5369,N_5470);
nand U5655 (N_5655,N_5329,N_5017);
nand U5656 (N_5656,N_5466,N_5159);
and U5657 (N_5657,N_5309,N_5355);
nor U5658 (N_5658,N_5364,N_5386);
nand U5659 (N_5659,N_5323,N_5488);
nor U5660 (N_5660,N_5280,N_5211);
and U5661 (N_5661,N_5039,N_5060);
nor U5662 (N_5662,N_5336,N_5065);
or U5663 (N_5663,N_5397,N_5305);
nand U5664 (N_5664,N_5101,N_5004);
nand U5665 (N_5665,N_5367,N_5480);
and U5666 (N_5666,N_5373,N_5212);
nand U5667 (N_5667,N_5062,N_5288);
or U5668 (N_5668,N_5051,N_5432);
nor U5669 (N_5669,N_5474,N_5249);
nor U5670 (N_5670,N_5351,N_5311);
and U5671 (N_5671,N_5146,N_5083);
or U5672 (N_5672,N_5086,N_5140);
nor U5673 (N_5673,N_5179,N_5097);
or U5674 (N_5674,N_5057,N_5419);
nand U5675 (N_5675,N_5321,N_5239);
nand U5676 (N_5676,N_5132,N_5026);
nor U5677 (N_5677,N_5213,N_5485);
nor U5678 (N_5678,N_5489,N_5242);
and U5679 (N_5679,N_5237,N_5418);
nor U5680 (N_5680,N_5214,N_5299);
or U5681 (N_5681,N_5256,N_5491);
and U5682 (N_5682,N_5071,N_5452);
xnor U5683 (N_5683,N_5044,N_5067);
or U5684 (N_5684,N_5150,N_5192);
or U5685 (N_5685,N_5155,N_5191);
and U5686 (N_5686,N_5319,N_5306);
and U5687 (N_5687,N_5201,N_5359);
and U5688 (N_5688,N_5469,N_5110);
and U5689 (N_5689,N_5449,N_5255);
and U5690 (N_5690,N_5460,N_5031);
or U5691 (N_5691,N_5430,N_5467);
nand U5692 (N_5692,N_5033,N_5301);
nand U5693 (N_5693,N_5210,N_5279);
and U5694 (N_5694,N_5073,N_5464);
and U5695 (N_5695,N_5180,N_5095);
and U5696 (N_5696,N_5232,N_5032);
nor U5697 (N_5697,N_5378,N_5127);
nand U5698 (N_5698,N_5098,N_5056);
nand U5699 (N_5699,N_5468,N_5333);
nor U5700 (N_5700,N_5206,N_5040);
nor U5701 (N_5701,N_5231,N_5066);
nand U5702 (N_5702,N_5021,N_5374);
and U5703 (N_5703,N_5384,N_5381);
nor U5704 (N_5704,N_5007,N_5235);
nand U5705 (N_5705,N_5293,N_5258);
or U5706 (N_5706,N_5494,N_5197);
or U5707 (N_5707,N_5024,N_5175);
and U5708 (N_5708,N_5143,N_5341);
nand U5709 (N_5709,N_5493,N_5076);
nor U5710 (N_5710,N_5375,N_5377);
nand U5711 (N_5711,N_5312,N_5439);
xnor U5712 (N_5712,N_5120,N_5283);
or U5713 (N_5713,N_5043,N_5416);
or U5714 (N_5714,N_5446,N_5181);
nand U5715 (N_5715,N_5342,N_5167);
and U5716 (N_5716,N_5476,N_5499);
and U5717 (N_5717,N_5011,N_5013);
nand U5718 (N_5718,N_5383,N_5422);
and U5719 (N_5719,N_5025,N_5002);
and U5720 (N_5720,N_5379,N_5014);
nor U5721 (N_5721,N_5058,N_5353);
nand U5722 (N_5722,N_5163,N_5047);
and U5723 (N_5723,N_5138,N_5404);
nor U5724 (N_5724,N_5338,N_5055);
or U5725 (N_5725,N_5216,N_5006);
nand U5726 (N_5726,N_5260,N_5015);
nand U5727 (N_5727,N_5454,N_5259);
nor U5728 (N_5728,N_5079,N_5490);
and U5729 (N_5729,N_5204,N_5141);
xor U5730 (N_5730,N_5271,N_5084);
and U5731 (N_5731,N_5009,N_5149);
nor U5732 (N_5732,N_5068,N_5274);
or U5733 (N_5733,N_5185,N_5022);
nand U5734 (N_5734,N_5276,N_5069);
nor U5735 (N_5735,N_5136,N_5265);
nor U5736 (N_5736,N_5471,N_5173);
nor U5737 (N_5737,N_5461,N_5188);
or U5738 (N_5738,N_5435,N_5203);
or U5739 (N_5739,N_5326,N_5292);
and U5740 (N_5740,N_5122,N_5220);
and U5741 (N_5741,N_5320,N_5440);
nand U5742 (N_5742,N_5070,N_5479);
nand U5743 (N_5743,N_5113,N_5437);
and U5744 (N_5744,N_5380,N_5354);
or U5745 (N_5745,N_5160,N_5234);
or U5746 (N_5746,N_5385,N_5400);
and U5747 (N_5747,N_5183,N_5139);
nand U5748 (N_5748,N_5156,N_5433);
nand U5749 (N_5749,N_5297,N_5145);
or U5750 (N_5750,N_5310,N_5111);
or U5751 (N_5751,N_5303,N_5026);
and U5752 (N_5752,N_5469,N_5023);
and U5753 (N_5753,N_5368,N_5393);
nor U5754 (N_5754,N_5178,N_5315);
and U5755 (N_5755,N_5340,N_5483);
xor U5756 (N_5756,N_5286,N_5026);
or U5757 (N_5757,N_5442,N_5484);
or U5758 (N_5758,N_5155,N_5148);
xnor U5759 (N_5759,N_5473,N_5233);
nand U5760 (N_5760,N_5088,N_5189);
nor U5761 (N_5761,N_5395,N_5001);
or U5762 (N_5762,N_5346,N_5243);
nor U5763 (N_5763,N_5365,N_5165);
nand U5764 (N_5764,N_5497,N_5232);
nor U5765 (N_5765,N_5458,N_5481);
and U5766 (N_5766,N_5215,N_5030);
and U5767 (N_5767,N_5497,N_5108);
or U5768 (N_5768,N_5009,N_5224);
nand U5769 (N_5769,N_5188,N_5351);
and U5770 (N_5770,N_5207,N_5109);
and U5771 (N_5771,N_5499,N_5445);
and U5772 (N_5772,N_5474,N_5453);
nor U5773 (N_5773,N_5390,N_5257);
or U5774 (N_5774,N_5131,N_5461);
and U5775 (N_5775,N_5389,N_5482);
or U5776 (N_5776,N_5418,N_5295);
and U5777 (N_5777,N_5088,N_5466);
nand U5778 (N_5778,N_5449,N_5403);
or U5779 (N_5779,N_5099,N_5222);
and U5780 (N_5780,N_5281,N_5107);
and U5781 (N_5781,N_5367,N_5020);
nand U5782 (N_5782,N_5272,N_5321);
nor U5783 (N_5783,N_5111,N_5494);
or U5784 (N_5784,N_5164,N_5083);
or U5785 (N_5785,N_5010,N_5256);
or U5786 (N_5786,N_5013,N_5217);
nor U5787 (N_5787,N_5220,N_5409);
nand U5788 (N_5788,N_5047,N_5276);
nand U5789 (N_5789,N_5242,N_5119);
nand U5790 (N_5790,N_5467,N_5253);
or U5791 (N_5791,N_5177,N_5000);
nor U5792 (N_5792,N_5336,N_5410);
nor U5793 (N_5793,N_5112,N_5258);
nand U5794 (N_5794,N_5484,N_5134);
nor U5795 (N_5795,N_5256,N_5378);
nand U5796 (N_5796,N_5375,N_5482);
nor U5797 (N_5797,N_5168,N_5189);
and U5798 (N_5798,N_5263,N_5348);
and U5799 (N_5799,N_5470,N_5123);
and U5800 (N_5800,N_5274,N_5477);
nor U5801 (N_5801,N_5001,N_5003);
nor U5802 (N_5802,N_5360,N_5232);
nand U5803 (N_5803,N_5245,N_5424);
nand U5804 (N_5804,N_5331,N_5452);
and U5805 (N_5805,N_5415,N_5269);
and U5806 (N_5806,N_5137,N_5355);
and U5807 (N_5807,N_5254,N_5251);
nand U5808 (N_5808,N_5152,N_5025);
nor U5809 (N_5809,N_5455,N_5251);
nor U5810 (N_5810,N_5025,N_5247);
and U5811 (N_5811,N_5276,N_5306);
or U5812 (N_5812,N_5433,N_5126);
nand U5813 (N_5813,N_5344,N_5069);
nor U5814 (N_5814,N_5294,N_5267);
nor U5815 (N_5815,N_5283,N_5027);
nand U5816 (N_5816,N_5460,N_5006);
xor U5817 (N_5817,N_5023,N_5076);
and U5818 (N_5818,N_5288,N_5246);
xnor U5819 (N_5819,N_5476,N_5137);
or U5820 (N_5820,N_5326,N_5278);
nor U5821 (N_5821,N_5300,N_5116);
and U5822 (N_5822,N_5233,N_5304);
xor U5823 (N_5823,N_5214,N_5200);
nand U5824 (N_5824,N_5344,N_5400);
and U5825 (N_5825,N_5226,N_5275);
nand U5826 (N_5826,N_5352,N_5219);
nand U5827 (N_5827,N_5268,N_5379);
nand U5828 (N_5828,N_5257,N_5405);
and U5829 (N_5829,N_5352,N_5455);
and U5830 (N_5830,N_5334,N_5491);
nand U5831 (N_5831,N_5286,N_5176);
or U5832 (N_5832,N_5216,N_5296);
or U5833 (N_5833,N_5355,N_5068);
and U5834 (N_5834,N_5129,N_5367);
nor U5835 (N_5835,N_5243,N_5447);
nor U5836 (N_5836,N_5378,N_5343);
nor U5837 (N_5837,N_5171,N_5266);
or U5838 (N_5838,N_5081,N_5294);
or U5839 (N_5839,N_5402,N_5220);
nand U5840 (N_5840,N_5408,N_5353);
or U5841 (N_5841,N_5112,N_5271);
nand U5842 (N_5842,N_5045,N_5002);
and U5843 (N_5843,N_5233,N_5341);
nand U5844 (N_5844,N_5154,N_5397);
and U5845 (N_5845,N_5097,N_5053);
nor U5846 (N_5846,N_5095,N_5355);
and U5847 (N_5847,N_5288,N_5269);
and U5848 (N_5848,N_5472,N_5438);
nor U5849 (N_5849,N_5252,N_5088);
and U5850 (N_5850,N_5229,N_5459);
nand U5851 (N_5851,N_5304,N_5438);
nor U5852 (N_5852,N_5378,N_5025);
and U5853 (N_5853,N_5064,N_5357);
or U5854 (N_5854,N_5465,N_5373);
or U5855 (N_5855,N_5423,N_5391);
nor U5856 (N_5856,N_5387,N_5142);
nand U5857 (N_5857,N_5253,N_5280);
nor U5858 (N_5858,N_5488,N_5284);
or U5859 (N_5859,N_5485,N_5246);
nor U5860 (N_5860,N_5005,N_5011);
nand U5861 (N_5861,N_5329,N_5049);
nand U5862 (N_5862,N_5448,N_5394);
and U5863 (N_5863,N_5189,N_5110);
or U5864 (N_5864,N_5286,N_5134);
and U5865 (N_5865,N_5202,N_5078);
nand U5866 (N_5866,N_5290,N_5382);
and U5867 (N_5867,N_5340,N_5425);
xor U5868 (N_5868,N_5317,N_5136);
nand U5869 (N_5869,N_5383,N_5455);
or U5870 (N_5870,N_5472,N_5453);
nand U5871 (N_5871,N_5379,N_5316);
nand U5872 (N_5872,N_5116,N_5428);
and U5873 (N_5873,N_5170,N_5127);
xor U5874 (N_5874,N_5478,N_5104);
or U5875 (N_5875,N_5408,N_5481);
nor U5876 (N_5876,N_5307,N_5234);
and U5877 (N_5877,N_5341,N_5142);
nand U5878 (N_5878,N_5405,N_5345);
and U5879 (N_5879,N_5218,N_5264);
and U5880 (N_5880,N_5262,N_5069);
nor U5881 (N_5881,N_5018,N_5078);
nor U5882 (N_5882,N_5133,N_5264);
and U5883 (N_5883,N_5436,N_5147);
xor U5884 (N_5884,N_5460,N_5160);
nor U5885 (N_5885,N_5253,N_5465);
nand U5886 (N_5886,N_5107,N_5261);
nor U5887 (N_5887,N_5249,N_5307);
or U5888 (N_5888,N_5267,N_5197);
nor U5889 (N_5889,N_5256,N_5327);
nand U5890 (N_5890,N_5102,N_5111);
nor U5891 (N_5891,N_5135,N_5247);
or U5892 (N_5892,N_5296,N_5220);
and U5893 (N_5893,N_5273,N_5270);
nand U5894 (N_5894,N_5283,N_5389);
nand U5895 (N_5895,N_5268,N_5071);
nand U5896 (N_5896,N_5163,N_5022);
or U5897 (N_5897,N_5119,N_5334);
nand U5898 (N_5898,N_5486,N_5393);
nand U5899 (N_5899,N_5009,N_5054);
or U5900 (N_5900,N_5486,N_5233);
or U5901 (N_5901,N_5132,N_5161);
or U5902 (N_5902,N_5316,N_5180);
nand U5903 (N_5903,N_5269,N_5203);
nor U5904 (N_5904,N_5159,N_5076);
and U5905 (N_5905,N_5038,N_5343);
and U5906 (N_5906,N_5221,N_5312);
and U5907 (N_5907,N_5447,N_5478);
nand U5908 (N_5908,N_5273,N_5264);
nor U5909 (N_5909,N_5035,N_5243);
and U5910 (N_5910,N_5204,N_5136);
nand U5911 (N_5911,N_5436,N_5037);
nor U5912 (N_5912,N_5437,N_5183);
and U5913 (N_5913,N_5056,N_5078);
nand U5914 (N_5914,N_5117,N_5253);
or U5915 (N_5915,N_5041,N_5485);
and U5916 (N_5916,N_5415,N_5472);
and U5917 (N_5917,N_5478,N_5242);
nand U5918 (N_5918,N_5020,N_5171);
and U5919 (N_5919,N_5316,N_5148);
or U5920 (N_5920,N_5359,N_5164);
or U5921 (N_5921,N_5464,N_5427);
nor U5922 (N_5922,N_5278,N_5321);
nand U5923 (N_5923,N_5065,N_5418);
and U5924 (N_5924,N_5160,N_5366);
nand U5925 (N_5925,N_5306,N_5028);
and U5926 (N_5926,N_5051,N_5297);
or U5927 (N_5927,N_5298,N_5135);
nand U5928 (N_5928,N_5341,N_5120);
nor U5929 (N_5929,N_5322,N_5197);
nor U5930 (N_5930,N_5192,N_5113);
nor U5931 (N_5931,N_5137,N_5021);
nor U5932 (N_5932,N_5271,N_5445);
and U5933 (N_5933,N_5371,N_5249);
or U5934 (N_5934,N_5258,N_5139);
and U5935 (N_5935,N_5484,N_5282);
and U5936 (N_5936,N_5420,N_5426);
nor U5937 (N_5937,N_5155,N_5130);
or U5938 (N_5938,N_5064,N_5079);
nor U5939 (N_5939,N_5152,N_5367);
xnor U5940 (N_5940,N_5413,N_5369);
or U5941 (N_5941,N_5341,N_5073);
or U5942 (N_5942,N_5298,N_5466);
nor U5943 (N_5943,N_5126,N_5070);
and U5944 (N_5944,N_5008,N_5051);
or U5945 (N_5945,N_5235,N_5355);
nor U5946 (N_5946,N_5418,N_5160);
nand U5947 (N_5947,N_5150,N_5247);
or U5948 (N_5948,N_5360,N_5419);
and U5949 (N_5949,N_5126,N_5376);
or U5950 (N_5950,N_5409,N_5108);
and U5951 (N_5951,N_5141,N_5254);
and U5952 (N_5952,N_5035,N_5215);
nand U5953 (N_5953,N_5042,N_5461);
nor U5954 (N_5954,N_5498,N_5018);
and U5955 (N_5955,N_5414,N_5261);
nand U5956 (N_5956,N_5093,N_5067);
or U5957 (N_5957,N_5290,N_5412);
and U5958 (N_5958,N_5024,N_5027);
and U5959 (N_5959,N_5067,N_5495);
xnor U5960 (N_5960,N_5363,N_5327);
and U5961 (N_5961,N_5264,N_5084);
nor U5962 (N_5962,N_5484,N_5087);
and U5963 (N_5963,N_5095,N_5484);
nand U5964 (N_5964,N_5369,N_5208);
nand U5965 (N_5965,N_5251,N_5062);
nor U5966 (N_5966,N_5107,N_5197);
or U5967 (N_5967,N_5320,N_5256);
nor U5968 (N_5968,N_5138,N_5270);
or U5969 (N_5969,N_5306,N_5385);
or U5970 (N_5970,N_5449,N_5288);
nor U5971 (N_5971,N_5203,N_5241);
nor U5972 (N_5972,N_5095,N_5194);
or U5973 (N_5973,N_5196,N_5031);
nand U5974 (N_5974,N_5230,N_5098);
nand U5975 (N_5975,N_5492,N_5185);
nor U5976 (N_5976,N_5306,N_5377);
or U5977 (N_5977,N_5302,N_5034);
or U5978 (N_5978,N_5497,N_5014);
xor U5979 (N_5979,N_5446,N_5183);
nand U5980 (N_5980,N_5228,N_5370);
and U5981 (N_5981,N_5421,N_5006);
nor U5982 (N_5982,N_5101,N_5057);
and U5983 (N_5983,N_5383,N_5484);
or U5984 (N_5984,N_5077,N_5291);
or U5985 (N_5985,N_5034,N_5018);
or U5986 (N_5986,N_5427,N_5311);
or U5987 (N_5987,N_5450,N_5477);
nor U5988 (N_5988,N_5393,N_5376);
nand U5989 (N_5989,N_5255,N_5459);
or U5990 (N_5990,N_5300,N_5037);
or U5991 (N_5991,N_5016,N_5310);
nand U5992 (N_5992,N_5001,N_5263);
nor U5993 (N_5993,N_5367,N_5346);
nand U5994 (N_5994,N_5149,N_5100);
nor U5995 (N_5995,N_5217,N_5463);
nor U5996 (N_5996,N_5460,N_5474);
nor U5997 (N_5997,N_5147,N_5292);
xor U5998 (N_5998,N_5270,N_5133);
nand U5999 (N_5999,N_5084,N_5348);
and U6000 (N_6000,N_5903,N_5642);
nor U6001 (N_6001,N_5788,N_5835);
nand U6002 (N_6002,N_5750,N_5791);
nand U6003 (N_6003,N_5610,N_5851);
nand U6004 (N_6004,N_5776,N_5550);
nand U6005 (N_6005,N_5652,N_5937);
xor U6006 (N_6006,N_5969,N_5618);
xnor U6007 (N_6007,N_5962,N_5692);
nand U6008 (N_6008,N_5898,N_5760);
nor U6009 (N_6009,N_5648,N_5814);
nand U6010 (N_6010,N_5649,N_5868);
and U6011 (N_6011,N_5737,N_5772);
and U6012 (N_6012,N_5529,N_5906);
nor U6013 (N_6013,N_5634,N_5650);
and U6014 (N_6014,N_5712,N_5540);
and U6015 (N_6015,N_5894,N_5576);
nand U6016 (N_6016,N_5724,N_5735);
or U6017 (N_6017,N_5913,N_5646);
nand U6018 (N_6018,N_5543,N_5731);
nor U6019 (N_6019,N_5780,N_5720);
and U6020 (N_6020,N_5516,N_5966);
and U6021 (N_6021,N_5883,N_5619);
nor U6022 (N_6022,N_5802,N_5804);
nand U6023 (N_6023,N_5664,N_5899);
and U6024 (N_6024,N_5869,N_5683);
nor U6025 (N_6025,N_5567,N_5909);
nor U6026 (N_6026,N_5663,N_5528);
or U6027 (N_6027,N_5577,N_5555);
nand U6028 (N_6028,N_5614,N_5721);
or U6029 (N_6029,N_5603,N_5758);
nor U6030 (N_6030,N_5511,N_5671);
nand U6031 (N_6031,N_5942,N_5792);
nor U6032 (N_6032,N_5584,N_5531);
xnor U6033 (N_6033,N_5732,N_5609);
or U6034 (N_6034,N_5669,N_5964);
or U6035 (N_6035,N_5939,N_5515);
nand U6036 (N_6036,N_5554,N_5960);
or U6037 (N_6037,N_5711,N_5800);
or U6038 (N_6038,N_5926,N_5774);
nand U6039 (N_6039,N_5687,N_5977);
and U6040 (N_6040,N_5775,N_5752);
and U6041 (N_6041,N_5840,N_5636);
nand U6042 (N_6042,N_5521,N_5885);
nor U6043 (N_6043,N_5963,N_5902);
nor U6044 (N_6044,N_5863,N_5625);
nor U6045 (N_6045,N_5900,N_5799);
nor U6046 (N_6046,N_5917,N_5631);
and U6047 (N_6047,N_5936,N_5651);
or U6048 (N_6048,N_5698,N_5510);
and U6049 (N_6049,N_5604,N_5542);
nand U6050 (N_6050,N_5596,N_5701);
or U6051 (N_6051,N_5598,N_5973);
nand U6052 (N_6052,N_5988,N_5884);
or U6053 (N_6053,N_5507,N_5993);
nor U6054 (N_6054,N_5946,N_5867);
xnor U6055 (N_6055,N_5512,N_5877);
nor U6056 (N_6056,N_5809,N_5585);
nand U6057 (N_6057,N_5933,N_5762);
nor U6058 (N_6058,N_5726,N_5880);
nor U6059 (N_6059,N_5864,N_5624);
nand U6060 (N_6060,N_5819,N_5722);
nand U6061 (N_6061,N_5976,N_5647);
or U6062 (N_6062,N_5565,N_5532);
and U6063 (N_6063,N_5754,N_5539);
nor U6064 (N_6064,N_5680,N_5954);
xor U6065 (N_6065,N_5667,N_5556);
or U6066 (N_6066,N_5872,N_5911);
nor U6067 (N_6067,N_5925,N_5615);
and U6068 (N_6068,N_5738,N_5620);
and U6069 (N_6069,N_5771,N_5816);
or U6070 (N_6070,N_5560,N_5796);
nor U6071 (N_6071,N_5574,N_5718);
nand U6072 (N_6072,N_5617,N_5928);
or U6073 (N_6073,N_5578,N_5996);
or U6074 (N_6074,N_5546,N_5725);
or U6075 (N_6075,N_5744,N_5825);
nand U6076 (N_6076,N_5790,N_5641);
and U6077 (N_6077,N_5789,N_5590);
nand U6078 (N_6078,N_5901,N_5811);
or U6079 (N_6079,N_5570,N_5950);
nand U6080 (N_6080,N_5681,N_5686);
nor U6081 (N_6081,N_5706,N_5713);
nor U6082 (N_6082,N_5871,N_5748);
nand U6083 (N_6083,N_5632,N_5889);
and U6084 (N_6084,N_5621,N_5935);
or U6085 (N_6085,N_5568,N_5806);
nor U6086 (N_6086,N_5945,N_5653);
and U6087 (N_6087,N_5786,N_5708);
nand U6088 (N_6088,N_5929,N_5612);
or U6089 (N_6089,N_5690,N_5968);
and U6090 (N_6090,N_5691,N_5918);
and U6091 (N_6091,N_5888,N_5530);
or U6092 (N_6092,N_5998,N_5583);
and U6093 (N_6093,N_5832,N_5672);
nand U6094 (N_6094,N_5795,N_5756);
and U6095 (N_6095,N_5639,N_5729);
nor U6096 (N_6096,N_5992,N_5716);
nor U6097 (N_6097,N_5658,N_5745);
and U6098 (N_6098,N_5734,N_5654);
or U6099 (N_6099,N_5882,N_5915);
nor U6100 (N_6100,N_5893,N_5534);
xor U6101 (N_6101,N_5581,N_5812);
nand U6102 (N_6102,N_5769,N_5949);
and U6103 (N_6103,N_5566,N_5857);
and U6104 (N_6104,N_5628,N_5839);
nand U6105 (N_6105,N_5519,N_5695);
or U6106 (N_6106,N_5740,N_5940);
nand U6107 (N_6107,N_5573,N_5517);
or U6108 (N_6108,N_5861,N_5859);
or U6109 (N_6109,N_5958,N_5891);
and U6110 (N_6110,N_5873,N_5502);
nand U6111 (N_6111,N_5699,N_5862);
and U6112 (N_6112,N_5808,N_5593);
nor U6113 (N_6113,N_5506,N_5645);
and U6114 (N_6114,N_5674,N_5741);
nor U6115 (N_6115,N_5616,N_5999);
or U6116 (N_6116,N_5675,N_5829);
or U6117 (N_6117,N_5904,N_5678);
nand U6118 (N_6118,N_5848,N_5895);
nor U6119 (N_6119,N_5728,N_5665);
and U6120 (N_6120,N_5520,N_5697);
nor U6121 (N_6121,N_5548,N_5633);
and U6122 (N_6122,N_5710,N_5948);
nand U6123 (N_6123,N_5854,N_5777);
nor U6124 (N_6124,N_5919,N_5597);
and U6125 (N_6125,N_5827,N_5858);
nand U6126 (N_6126,N_5500,N_5533);
nand U6127 (N_6127,N_5525,N_5707);
xnor U6128 (N_6128,N_5763,N_5773);
nor U6129 (N_6129,N_5875,N_5905);
nand U6130 (N_6130,N_5561,N_5552);
or U6131 (N_6131,N_5892,N_5673);
and U6132 (N_6132,N_5759,N_5580);
nand U6133 (N_6133,N_5965,N_5696);
nor U6134 (N_6134,N_5944,N_5717);
nor U6135 (N_6135,N_5957,N_5833);
nor U6136 (N_6136,N_5881,N_5817);
and U6137 (N_6137,N_5821,N_5914);
nor U6138 (N_6138,N_5970,N_5504);
nor U6139 (N_6139,N_5505,N_5587);
nand U6140 (N_6140,N_5783,N_5844);
and U6141 (N_6141,N_5828,N_5757);
nor U6142 (N_6142,N_5770,N_5635);
and U6143 (N_6143,N_5779,N_5622);
nand U6144 (N_6144,N_5694,N_5997);
nor U6145 (N_6145,N_5630,N_5700);
or U6146 (N_6146,N_5599,N_5600);
nor U6147 (N_6147,N_5953,N_5685);
nand U6148 (N_6148,N_5736,N_5805);
or U6149 (N_6149,N_5987,N_5594);
and U6150 (N_6150,N_5842,N_5638);
and U6151 (N_6151,N_5715,N_5606);
or U6152 (N_6152,N_5764,N_5979);
nor U6153 (N_6153,N_5535,N_5781);
and U6154 (N_6154,N_5656,N_5569);
and U6155 (N_6155,N_5518,N_5865);
or U6156 (N_6156,N_5661,N_5676);
or U6157 (N_6157,N_5660,N_5723);
and U6158 (N_6158,N_5719,N_5682);
or U6159 (N_6159,N_5765,N_5582);
or U6160 (N_6160,N_5541,N_5579);
and U6161 (N_6161,N_5818,N_5916);
and U6162 (N_6162,N_5956,N_5834);
and U6163 (N_6163,N_5934,N_5659);
nand U6164 (N_6164,N_5984,N_5586);
xnor U6165 (N_6165,N_5727,N_5886);
nor U6166 (N_6166,N_5749,N_5513);
nand U6167 (N_6167,N_5855,N_5524);
nand U6168 (N_6168,N_5709,N_5822);
nor U6169 (N_6169,N_5559,N_5830);
or U6170 (N_6170,N_5766,N_5921);
or U6171 (N_6171,N_5689,N_5994);
and U6172 (N_6172,N_5755,N_5608);
nand U6173 (N_6173,N_5547,N_5688);
nor U6174 (N_6174,N_5611,N_5975);
or U6175 (N_6175,N_5982,N_5938);
or U6176 (N_6176,N_5924,N_5971);
and U6177 (N_6177,N_5959,N_5767);
xor U6178 (N_6178,N_5508,N_5787);
or U6179 (N_6179,N_5846,N_5501);
nand U6180 (N_6180,N_5536,N_5589);
and U6181 (N_6181,N_5784,N_5558);
and U6182 (N_6182,N_5952,N_5705);
or U6183 (N_6183,N_5850,N_5714);
and U6184 (N_6184,N_5836,N_5551);
nor U6185 (N_6185,N_5537,N_5843);
and U6186 (N_6186,N_5592,N_5803);
nor U6187 (N_6187,N_5793,N_5657);
nor U6188 (N_6188,N_5961,N_5887);
nor U6189 (N_6189,N_5640,N_5602);
or U6190 (N_6190,N_5986,N_5798);
nor U6191 (N_6191,N_5637,N_5831);
and U6192 (N_6192,N_5522,N_5991);
nand U6193 (N_6193,N_5878,N_5753);
or U6194 (N_6194,N_5820,N_5703);
and U6195 (N_6195,N_5983,N_5823);
or U6196 (N_6196,N_5778,N_5739);
and U6197 (N_6197,N_5605,N_5702);
or U6198 (N_6198,N_5747,N_5563);
nand U6199 (N_6199,N_5562,N_5751);
nand U6200 (N_6200,N_5845,N_5538);
nand U6201 (N_6201,N_5866,N_5662);
nor U6202 (N_6202,N_5981,N_5761);
nor U6203 (N_6203,N_5523,N_5613);
or U6204 (N_6204,N_5841,N_5932);
or U6205 (N_6205,N_5879,N_5572);
nand U6206 (N_6206,N_5927,N_5967);
or U6207 (N_6207,N_5972,N_5627);
nor U6208 (N_6208,N_5782,N_5852);
nand U6209 (N_6209,N_5943,N_5629);
and U6210 (N_6210,N_5838,N_5601);
nor U6211 (N_6211,N_5549,N_5930);
or U6212 (N_6212,N_5826,N_5923);
nand U6213 (N_6213,N_5874,N_5666);
and U6214 (N_6214,N_5890,N_5668);
or U6215 (N_6215,N_5704,N_5797);
or U6216 (N_6216,N_5974,N_5509);
or U6217 (N_6217,N_5643,N_5553);
or U6218 (N_6218,N_5557,N_5514);
and U6219 (N_6219,N_5837,N_5545);
and U6220 (N_6220,N_5985,N_5860);
nor U6221 (N_6221,N_5670,N_5807);
or U6222 (N_6222,N_5995,N_5876);
nand U6223 (N_6223,N_5743,N_5677);
nor U6224 (N_6224,N_5785,N_5746);
or U6225 (N_6225,N_5655,N_5626);
nand U6226 (N_6226,N_5941,N_5931);
nand U6227 (N_6227,N_5730,N_5742);
nand U6228 (N_6228,N_5813,N_5768);
nor U6229 (N_6229,N_5955,N_5824);
or U6230 (N_6230,N_5908,N_5693);
and U6231 (N_6231,N_5623,N_5951);
or U6232 (N_6232,N_5920,N_5980);
or U6233 (N_6233,N_5801,N_5527);
nand U6234 (N_6234,N_5595,N_5849);
nand U6235 (N_6235,N_5912,N_5910);
nor U6236 (N_6236,N_5544,N_5571);
nor U6237 (N_6237,N_5644,N_5853);
and U6238 (N_6238,N_5870,N_5607);
nand U6239 (N_6239,N_5503,N_5856);
or U6240 (N_6240,N_5564,N_5896);
or U6241 (N_6241,N_5575,N_5815);
nand U6242 (N_6242,N_5684,N_5591);
and U6243 (N_6243,N_5978,N_5794);
nand U6244 (N_6244,N_5947,N_5922);
nand U6245 (N_6245,N_5990,N_5810);
or U6246 (N_6246,N_5679,N_5897);
or U6247 (N_6247,N_5907,N_5588);
or U6248 (N_6248,N_5847,N_5733);
and U6249 (N_6249,N_5526,N_5989);
or U6250 (N_6250,N_5854,N_5882);
or U6251 (N_6251,N_5631,N_5618);
or U6252 (N_6252,N_5621,N_5975);
and U6253 (N_6253,N_5640,N_5627);
nor U6254 (N_6254,N_5970,N_5674);
or U6255 (N_6255,N_5812,N_5831);
or U6256 (N_6256,N_5703,N_5595);
nand U6257 (N_6257,N_5634,N_5866);
nor U6258 (N_6258,N_5966,N_5849);
or U6259 (N_6259,N_5919,N_5912);
or U6260 (N_6260,N_5645,N_5634);
xnor U6261 (N_6261,N_5622,N_5686);
or U6262 (N_6262,N_5956,N_5755);
nor U6263 (N_6263,N_5540,N_5806);
nand U6264 (N_6264,N_5951,N_5699);
and U6265 (N_6265,N_5700,N_5624);
nand U6266 (N_6266,N_5641,N_5976);
and U6267 (N_6267,N_5870,N_5970);
or U6268 (N_6268,N_5507,N_5934);
nor U6269 (N_6269,N_5964,N_5688);
nor U6270 (N_6270,N_5642,N_5896);
or U6271 (N_6271,N_5614,N_5960);
nor U6272 (N_6272,N_5921,N_5923);
nand U6273 (N_6273,N_5563,N_5722);
and U6274 (N_6274,N_5980,N_5946);
xor U6275 (N_6275,N_5860,N_5651);
nor U6276 (N_6276,N_5954,N_5924);
and U6277 (N_6277,N_5812,N_5714);
or U6278 (N_6278,N_5812,N_5991);
nor U6279 (N_6279,N_5822,N_5737);
or U6280 (N_6280,N_5529,N_5763);
nor U6281 (N_6281,N_5563,N_5657);
nor U6282 (N_6282,N_5687,N_5996);
nand U6283 (N_6283,N_5628,N_5932);
and U6284 (N_6284,N_5555,N_5811);
or U6285 (N_6285,N_5706,N_5773);
nand U6286 (N_6286,N_5922,N_5984);
or U6287 (N_6287,N_5944,N_5748);
nand U6288 (N_6288,N_5897,N_5712);
nor U6289 (N_6289,N_5710,N_5994);
nor U6290 (N_6290,N_5776,N_5694);
nor U6291 (N_6291,N_5953,N_5687);
and U6292 (N_6292,N_5796,N_5958);
or U6293 (N_6293,N_5640,N_5705);
nor U6294 (N_6294,N_5738,N_5740);
nor U6295 (N_6295,N_5736,N_5872);
nor U6296 (N_6296,N_5853,N_5536);
nor U6297 (N_6297,N_5587,N_5576);
and U6298 (N_6298,N_5942,N_5950);
nand U6299 (N_6299,N_5590,N_5968);
nand U6300 (N_6300,N_5619,N_5846);
and U6301 (N_6301,N_5978,N_5681);
nor U6302 (N_6302,N_5933,N_5681);
nand U6303 (N_6303,N_5953,N_5973);
or U6304 (N_6304,N_5954,N_5691);
and U6305 (N_6305,N_5966,N_5896);
nor U6306 (N_6306,N_5691,N_5501);
or U6307 (N_6307,N_5758,N_5672);
nor U6308 (N_6308,N_5836,N_5687);
and U6309 (N_6309,N_5756,N_5577);
and U6310 (N_6310,N_5552,N_5688);
or U6311 (N_6311,N_5954,N_5846);
nor U6312 (N_6312,N_5572,N_5966);
or U6313 (N_6313,N_5716,N_5771);
xnor U6314 (N_6314,N_5901,N_5833);
or U6315 (N_6315,N_5542,N_5794);
nor U6316 (N_6316,N_5838,N_5680);
and U6317 (N_6317,N_5563,N_5888);
and U6318 (N_6318,N_5895,N_5718);
nor U6319 (N_6319,N_5780,N_5756);
nor U6320 (N_6320,N_5999,N_5533);
and U6321 (N_6321,N_5608,N_5853);
nor U6322 (N_6322,N_5540,N_5618);
or U6323 (N_6323,N_5939,N_5820);
and U6324 (N_6324,N_5637,N_5995);
or U6325 (N_6325,N_5790,N_5637);
and U6326 (N_6326,N_5708,N_5621);
nand U6327 (N_6327,N_5868,N_5861);
or U6328 (N_6328,N_5876,N_5923);
nand U6329 (N_6329,N_5803,N_5978);
xnor U6330 (N_6330,N_5573,N_5528);
nand U6331 (N_6331,N_5861,N_5984);
nand U6332 (N_6332,N_5728,N_5533);
nor U6333 (N_6333,N_5581,N_5529);
and U6334 (N_6334,N_5819,N_5857);
nand U6335 (N_6335,N_5913,N_5817);
nor U6336 (N_6336,N_5750,N_5730);
or U6337 (N_6337,N_5915,N_5609);
or U6338 (N_6338,N_5761,N_5757);
or U6339 (N_6339,N_5986,N_5775);
nor U6340 (N_6340,N_5814,N_5863);
or U6341 (N_6341,N_5966,N_5702);
nor U6342 (N_6342,N_5920,N_5837);
and U6343 (N_6343,N_5653,N_5565);
nand U6344 (N_6344,N_5714,N_5575);
and U6345 (N_6345,N_5825,N_5546);
nand U6346 (N_6346,N_5636,N_5895);
nand U6347 (N_6347,N_5778,N_5937);
nand U6348 (N_6348,N_5941,N_5869);
nand U6349 (N_6349,N_5867,N_5667);
and U6350 (N_6350,N_5973,N_5551);
nand U6351 (N_6351,N_5902,N_5847);
or U6352 (N_6352,N_5783,N_5800);
and U6353 (N_6353,N_5548,N_5586);
or U6354 (N_6354,N_5724,N_5855);
nor U6355 (N_6355,N_5858,N_5880);
nor U6356 (N_6356,N_5779,N_5948);
or U6357 (N_6357,N_5613,N_5527);
nor U6358 (N_6358,N_5908,N_5856);
and U6359 (N_6359,N_5840,N_5851);
or U6360 (N_6360,N_5612,N_5624);
and U6361 (N_6361,N_5614,N_5749);
nor U6362 (N_6362,N_5844,N_5584);
nand U6363 (N_6363,N_5904,N_5547);
nor U6364 (N_6364,N_5901,N_5705);
nand U6365 (N_6365,N_5676,N_5752);
nor U6366 (N_6366,N_5709,N_5899);
nor U6367 (N_6367,N_5744,N_5995);
and U6368 (N_6368,N_5733,N_5627);
or U6369 (N_6369,N_5718,N_5504);
and U6370 (N_6370,N_5614,N_5951);
or U6371 (N_6371,N_5623,N_5900);
nand U6372 (N_6372,N_5531,N_5917);
nand U6373 (N_6373,N_5543,N_5507);
and U6374 (N_6374,N_5923,N_5742);
and U6375 (N_6375,N_5618,N_5509);
nor U6376 (N_6376,N_5656,N_5505);
nand U6377 (N_6377,N_5741,N_5749);
or U6378 (N_6378,N_5654,N_5911);
nand U6379 (N_6379,N_5882,N_5920);
nand U6380 (N_6380,N_5534,N_5655);
nand U6381 (N_6381,N_5632,N_5746);
nand U6382 (N_6382,N_5781,N_5621);
nor U6383 (N_6383,N_5802,N_5688);
nand U6384 (N_6384,N_5690,N_5691);
nand U6385 (N_6385,N_5671,N_5621);
and U6386 (N_6386,N_5579,N_5703);
nand U6387 (N_6387,N_5520,N_5932);
nor U6388 (N_6388,N_5729,N_5564);
or U6389 (N_6389,N_5566,N_5897);
xnor U6390 (N_6390,N_5934,N_5853);
or U6391 (N_6391,N_5518,N_5517);
or U6392 (N_6392,N_5526,N_5636);
or U6393 (N_6393,N_5975,N_5971);
or U6394 (N_6394,N_5931,N_5809);
and U6395 (N_6395,N_5760,N_5986);
nor U6396 (N_6396,N_5745,N_5627);
nand U6397 (N_6397,N_5609,N_5816);
nand U6398 (N_6398,N_5794,N_5706);
xor U6399 (N_6399,N_5699,N_5505);
nor U6400 (N_6400,N_5728,N_5536);
or U6401 (N_6401,N_5542,N_5765);
nor U6402 (N_6402,N_5893,N_5701);
or U6403 (N_6403,N_5537,N_5846);
or U6404 (N_6404,N_5751,N_5594);
and U6405 (N_6405,N_5507,N_5937);
nor U6406 (N_6406,N_5737,N_5798);
or U6407 (N_6407,N_5702,N_5872);
and U6408 (N_6408,N_5711,N_5843);
nor U6409 (N_6409,N_5550,N_5609);
nor U6410 (N_6410,N_5761,N_5583);
nor U6411 (N_6411,N_5836,N_5868);
xor U6412 (N_6412,N_5506,N_5589);
nand U6413 (N_6413,N_5892,N_5532);
nor U6414 (N_6414,N_5599,N_5533);
or U6415 (N_6415,N_5900,N_5969);
nor U6416 (N_6416,N_5926,N_5982);
and U6417 (N_6417,N_5719,N_5990);
or U6418 (N_6418,N_5525,N_5743);
and U6419 (N_6419,N_5799,N_5907);
nand U6420 (N_6420,N_5902,N_5820);
nand U6421 (N_6421,N_5749,N_5793);
nand U6422 (N_6422,N_5723,N_5999);
or U6423 (N_6423,N_5873,N_5952);
nor U6424 (N_6424,N_5976,N_5835);
and U6425 (N_6425,N_5926,N_5642);
nor U6426 (N_6426,N_5810,N_5515);
or U6427 (N_6427,N_5531,N_5512);
nor U6428 (N_6428,N_5881,N_5762);
nand U6429 (N_6429,N_5947,N_5581);
or U6430 (N_6430,N_5735,N_5539);
or U6431 (N_6431,N_5557,N_5763);
nand U6432 (N_6432,N_5793,N_5947);
nor U6433 (N_6433,N_5796,N_5616);
nor U6434 (N_6434,N_5930,N_5672);
nand U6435 (N_6435,N_5891,N_5872);
nand U6436 (N_6436,N_5780,N_5786);
nor U6437 (N_6437,N_5772,N_5872);
nand U6438 (N_6438,N_5793,N_5909);
nand U6439 (N_6439,N_5813,N_5726);
or U6440 (N_6440,N_5618,N_5537);
nor U6441 (N_6441,N_5759,N_5695);
or U6442 (N_6442,N_5979,N_5770);
nor U6443 (N_6443,N_5773,N_5934);
nand U6444 (N_6444,N_5723,N_5591);
nor U6445 (N_6445,N_5654,N_5516);
and U6446 (N_6446,N_5973,N_5659);
or U6447 (N_6447,N_5763,N_5619);
and U6448 (N_6448,N_5639,N_5676);
and U6449 (N_6449,N_5728,N_5903);
or U6450 (N_6450,N_5641,N_5826);
nand U6451 (N_6451,N_5587,N_5943);
or U6452 (N_6452,N_5944,N_5765);
and U6453 (N_6453,N_5962,N_5761);
nand U6454 (N_6454,N_5736,N_5930);
or U6455 (N_6455,N_5960,N_5818);
nor U6456 (N_6456,N_5759,N_5786);
nand U6457 (N_6457,N_5668,N_5633);
or U6458 (N_6458,N_5721,N_5956);
nand U6459 (N_6459,N_5876,N_5998);
or U6460 (N_6460,N_5509,N_5862);
nand U6461 (N_6461,N_5850,N_5511);
and U6462 (N_6462,N_5956,N_5743);
nand U6463 (N_6463,N_5577,N_5786);
nor U6464 (N_6464,N_5794,N_5647);
or U6465 (N_6465,N_5504,N_5530);
nor U6466 (N_6466,N_5758,N_5518);
nor U6467 (N_6467,N_5933,N_5903);
nor U6468 (N_6468,N_5974,N_5695);
nand U6469 (N_6469,N_5780,N_5636);
nor U6470 (N_6470,N_5751,N_5557);
or U6471 (N_6471,N_5776,N_5927);
nand U6472 (N_6472,N_5777,N_5936);
nand U6473 (N_6473,N_5713,N_5774);
or U6474 (N_6474,N_5914,N_5622);
nand U6475 (N_6475,N_5786,N_5958);
nand U6476 (N_6476,N_5631,N_5769);
nand U6477 (N_6477,N_5768,N_5948);
nand U6478 (N_6478,N_5809,N_5973);
and U6479 (N_6479,N_5549,N_5792);
or U6480 (N_6480,N_5504,N_5562);
nor U6481 (N_6481,N_5654,N_5503);
nor U6482 (N_6482,N_5896,N_5733);
or U6483 (N_6483,N_5837,N_5878);
nand U6484 (N_6484,N_5924,N_5631);
and U6485 (N_6485,N_5671,N_5921);
nand U6486 (N_6486,N_5622,N_5908);
nor U6487 (N_6487,N_5569,N_5996);
nand U6488 (N_6488,N_5634,N_5976);
nor U6489 (N_6489,N_5826,N_5751);
nor U6490 (N_6490,N_5622,N_5630);
or U6491 (N_6491,N_5711,N_5515);
nand U6492 (N_6492,N_5638,N_5614);
or U6493 (N_6493,N_5906,N_5506);
and U6494 (N_6494,N_5749,N_5521);
nor U6495 (N_6495,N_5885,N_5602);
nor U6496 (N_6496,N_5623,N_5646);
and U6497 (N_6497,N_5662,N_5925);
nand U6498 (N_6498,N_5829,N_5930);
or U6499 (N_6499,N_5707,N_5797);
and U6500 (N_6500,N_6015,N_6022);
and U6501 (N_6501,N_6318,N_6054);
or U6502 (N_6502,N_6096,N_6228);
nand U6503 (N_6503,N_6176,N_6001);
nor U6504 (N_6504,N_6213,N_6295);
nand U6505 (N_6505,N_6175,N_6117);
nor U6506 (N_6506,N_6358,N_6134);
nor U6507 (N_6507,N_6385,N_6173);
and U6508 (N_6508,N_6281,N_6434);
nor U6509 (N_6509,N_6480,N_6126);
nor U6510 (N_6510,N_6441,N_6377);
and U6511 (N_6511,N_6296,N_6216);
nand U6512 (N_6512,N_6143,N_6429);
and U6513 (N_6513,N_6060,N_6129);
nor U6514 (N_6514,N_6475,N_6118);
nor U6515 (N_6515,N_6158,N_6155);
nor U6516 (N_6516,N_6005,N_6468);
or U6517 (N_6517,N_6045,N_6363);
nor U6518 (N_6518,N_6386,N_6380);
nor U6519 (N_6519,N_6451,N_6472);
or U6520 (N_6520,N_6407,N_6337);
or U6521 (N_6521,N_6471,N_6348);
nand U6522 (N_6522,N_6113,N_6368);
nand U6523 (N_6523,N_6024,N_6391);
nand U6524 (N_6524,N_6362,N_6378);
nor U6525 (N_6525,N_6376,N_6254);
or U6526 (N_6526,N_6414,N_6319);
or U6527 (N_6527,N_6456,N_6427);
nand U6528 (N_6528,N_6112,N_6425);
or U6529 (N_6529,N_6459,N_6011);
nor U6530 (N_6530,N_6102,N_6068);
and U6531 (N_6531,N_6186,N_6342);
nor U6532 (N_6532,N_6244,N_6327);
nand U6533 (N_6533,N_6273,N_6283);
and U6534 (N_6534,N_6465,N_6181);
nand U6535 (N_6535,N_6087,N_6182);
and U6536 (N_6536,N_6360,N_6394);
or U6537 (N_6537,N_6245,N_6161);
nor U6538 (N_6538,N_6390,N_6311);
nand U6539 (N_6539,N_6092,N_6497);
or U6540 (N_6540,N_6089,N_6232);
or U6541 (N_6541,N_6168,N_6339);
or U6542 (N_6542,N_6462,N_6200);
or U6543 (N_6543,N_6028,N_6114);
nand U6544 (N_6544,N_6374,N_6490);
nand U6545 (N_6545,N_6449,N_6413);
nor U6546 (N_6546,N_6300,N_6235);
nor U6547 (N_6547,N_6344,N_6016);
nand U6548 (N_6548,N_6473,N_6333);
or U6549 (N_6549,N_6077,N_6306);
nor U6550 (N_6550,N_6018,N_6201);
nand U6551 (N_6551,N_6185,N_6119);
and U6552 (N_6552,N_6217,N_6152);
nor U6553 (N_6553,N_6046,N_6225);
and U6554 (N_6554,N_6088,N_6049);
nor U6555 (N_6555,N_6417,N_6169);
nand U6556 (N_6556,N_6063,N_6259);
nand U6557 (N_6557,N_6224,N_6345);
nand U6558 (N_6558,N_6062,N_6261);
nand U6559 (N_6559,N_6220,N_6108);
nand U6560 (N_6560,N_6234,N_6369);
and U6561 (N_6561,N_6267,N_6236);
or U6562 (N_6562,N_6122,N_6214);
or U6563 (N_6563,N_6042,N_6384);
nor U6564 (N_6564,N_6106,N_6304);
and U6565 (N_6565,N_6411,N_6227);
nor U6566 (N_6566,N_6041,N_6325);
and U6567 (N_6567,N_6021,N_6193);
and U6568 (N_6568,N_6257,N_6359);
and U6569 (N_6569,N_6381,N_6095);
or U6570 (N_6570,N_6316,N_6310);
and U6571 (N_6571,N_6166,N_6388);
or U6572 (N_6572,N_6489,N_6432);
and U6573 (N_6573,N_6293,N_6299);
or U6574 (N_6574,N_6066,N_6131);
and U6575 (N_6575,N_6171,N_6396);
nand U6576 (N_6576,N_6419,N_6150);
or U6577 (N_6577,N_6099,N_6104);
or U6578 (N_6578,N_6308,N_6035);
or U6579 (N_6579,N_6057,N_6382);
and U6580 (N_6580,N_6079,N_6167);
and U6581 (N_6581,N_6073,N_6215);
or U6582 (N_6582,N_6032,N_6205);
or U6583 (N_6583,N_6094,N_6233);
nor U6584 (N_6584,N_6443,N_6324);
nand U6585 (N_6585,N_6485,N_6460);
nand U6586 (N_6586,N_6002,N_6086);
nand U6587 (N_6587,N_6253,N_6255);
and U6588 (N_6588,N_6379,N_6195);
and U6589 (N_6589,N_6477,N_6194);
or U6590 (N_6590,N_6162,N_6137);
nand U6591 (N_6591,N_6353,N_6469);
nor U6592 (N_6592,N_6450,N_6053);
nor U6593 (N_6593,N_6499,N_6493);
nand U6594 (N_6594,N_6444,N_6492);
nor U6595 (N_6595,N_6078,N_6019);
nand U6596 (N_6596,N_6211,N_6426);
and U6597 (N_6597,N_6398,N_6340);
nor U6598 (N_6598,N_6415,N_6470);
or U6599 (N_6599,N_6303,N_6111);
nand U6600 (N_6600,N_6305,N_6356);
nor U6601 (N_6601,N_6481,N_6222);
or U6602 (N_6602,N_6457,N_6133);
nor U6603 (N_6603,N_6070,N_6190);
and U6604 (N_6604,N_6128,N_6071);
or U6605 (N_6605,N_6424,N_6284);
nand U6606 (N_6606,N_6445,N_6315);
nor U6607 (N_6607,N_6036,N_6055);
and U6608 (N_6608,N_6297,N_6031);
or U6609 (N_6609,N_6160,N_6349);
xnor U6610 (N_6610,N_6007,N_6229);
or U6611 (N_6611,N_6482,N_6240);
xor U6612 (N_6612,N_6314,N_6188);
or U6613 (N_6613,N_6332,N_6393);
or U6614 (N_6614,N_6208,N_6266);
nor U6615 (N_6615,N_6263,N_6288);
nor U6616 (N_6616,N_6474,N_6455);
nor U6617 (N_6617,N_6110,N_6335);
nand U6618 (N_6618,N_6370,N_6187);
nand U6619 (N_6619,N_6237,N_6392);
nand U6620 (N_6620,N_6412,N_6203);
nor U6621 (N_6621,N_6221,N_6000);
nor U6622 (N_6622,N_6366,N_6135);
nand U6623 (N_6623,N_6159,N_6009);
or U6624 (N_6624,N_6218,N_6163);
or U6625 (N_6625,N_6248,N_6256);
nand U6626 (N_6626,N_6210,N_6403);
nor U6627 (N_6627,N_6483,N_6436);
nand U6628 (N_6628,N_6453,N_6180);
or U6629 (N_6629,N_6437,N_6438);
and U6630 (N_6630,N_6479,N_6280);
nand U6631 (N_6631,N_6268,N_6097);
nor U6632 (N_6632,N_6389,N_6278);
nor U6633 (N_6633,N_6361,N_6383);
nor U6634 (N_6634,N_6026,N_6416);
or U6635 (N_6635,N_6476,N_6399);
and U6636 (N_6636,N_6090,N_6048);
nor U6637 (N_6637,N_6323,N_6302);
and U6638 (N_6638,N_6085,N_6331);
nand U6639 (N_6639,N_6226,N_6209);
nor U6640 (N_6640,N_6025,N_6013);
and U6641 (N_6641,N_6027,N_6294);
or U6642 (N_6642,N_6329,N_6404);
nor U6643 (N_6643,N_6290,N_6276);
or U6644 (N_6644,N_6487,N_6047);
nor U6645 (N_6645,N_6017,N_6375);
xnor U6646 (N_6646,N_6165,N_6080);
nor U6647 (N_6647,N_6145,N_6153);
or U6648 (N_6648,N_6367,N_6037);
and U6649 (N_6649,N_6464,N_6291);
or U6650 (N_6650,N_6498,N_6183);
and U6651 (N_6651,N_6322,N_6207);
nand U6652 (N_6652,N_6372,N_6198);
nor U6653 (N_6653,N_6156,N_6346);
nand U6654 (N_6654,N_6287,N_6116);
and U6655 (N_6655,N_6204,N_6402);
or U6656 (N_6656,N_6272,N_6478);
and U6657 (N_6657,N_6357,N_6251);
nand U6658 (N_6658,N_6400,N_6439);
nand U6659 (N_6659,N_6127,N_6039);
nand U6660 (N_6660,N_6149,N_6242);
nand U6661 (N_6661,N_6336,N_6285);
or U6662 (N_6662,N_6050,N_6270);
nand U6663 (N_6663,N_6212,N_6466);
or U6664 (N_6664,N_6279,N_6141);
or U6665 (N_6665,N_6130,N_6120);
or U6666 (N_6666,N_6387,N_6275);
nand U6667 (N_6667,N_6023,N_6132);
nor U6668 (N_6668,N_6355,N_6334);
or U6669 (N_6669,N_6052,N_6282);
nand U6670 (N_6670,N_6328,N_6494);
and U6671 (N_6671,N_6365,N_6074);
nor U6672 (N_6672,N_6431,N_6231);
nand U6673 (N_6673,N_6406,N_6286);
nand U6674 (N_6674,N_6184,N_6313);
and U6675 (N_6675,N_6421,N_6059);
or U6676 (N_6676,N_6298,N_6004);
nor U6677 (N_6677,N_6030,N_6252);
nand U6678 (N_6678,N_6418,N_6056);
or U6679 (N_6679,N_6238,N_6069);
nor U6680 (N_6680,N_6202,N_6189);
or U6681 (N_6681,N_6246,N_6148);
and U6682 (N_6682,N_6264,N_6100);
nor U6683 (N_6683,N_6409,N_6223);
and U6684 (N_6684,N_6309,N_6467);
or U6685 (N_6685,N_6241,N_6098);
or U6686 (N_6686,N_6250,N_6410);
or U6687 (N_6687,N_6491,N_6174);
xor U6688 (N_6688,N_6373,N_6012);
nor U6689 (N_6689,N_6454,N_6420);
and U6690 (N_6690,N_6197,N_6307);
nor U6691 (N_6691,N_6142,N_6051);
and U6692 (N_6692,N_6364,N_6486);
and U6693 (N_6693,N_6247,N_6458);
xor U6694 (N_6694,N_6433,N_6044);
nor U6695 (N_6695,N_6343,N_6371);
nor U6696 (N_6696,N_6067,N_6338);
or U6697 (N_6697,N_6351,N_6125);
or U6698 (N_6698,N_6292,N_6179);
nor U6699 (N_6699,N_6230,N_6447);
nor U6700 (N_6700,N_6265,N_6043);
or U6701 (N_6701,N_6347,N_6330);
nand U6702 (N_6702,N_6107,N_6350);
nor U6703 (N_6703,N_6239,N_6423);
nand U6704 (N_6704,N_6082,N_6010);
nand U6705 (N_6705,N_6003,N_6196);
and U6706 (N_6706,N_6014,N_6191);
and U6707 (N_6707,N_6260,N_6147);
or U6708 (N_6708,N_6146,N_6061);
or U6709 (N_6709,N_6033,N_6405);
nor U6710 (N_6710,N_6139,N_6154);
nand U6711 (N_6711,N_6326,N_6081);
nand U6712 (N_6712,N_6354,N_6271);
nor U6713 (N_6713,N_6177,N_6395);
nor U6714 (N_6714,N_6262,N_6124);
nand U6715 (N_6715,N_6463,N_6093);
nor U6716 (N_6716,N_6164,N_6064);
nand U6717 (N_6717,N_6408,N_6199);
xor U6718 (N_6718,N_6422,N_6452);
and U6719 (N_6719,N_6496,N_6115);
nor U6720 (N_6720,N_6428,N_6034);
nor U6721 (N_6721,N_6072,N_6101);
xnor U6722 (N_6722,N_6435,N_6430);
nor U6723 (N_6723,N_6312,N_6488);
and U6724 (N_6724,N_6065,N_6192);
nor U6725 (N_6725,N_6446,N_6144);
nand U6726 (N_6726,N_6206,N_6151);
nand U6727 (N_6727,N_6140,N_6301);
nor U6728 (N_6728,N_6121,N_6084);
and U6729 (N_6729,N_6076,N_6495);
or U6730 (N_6730,N_6440,N_6109);
or U6731 (N_6731,N_6277,N_6289);
nand U6732 (N_6732,N_6352,N_6058);
nand U6733 (N_6733,N_6038,N_6448);
nor U6734 (N_6734,N_6170,N_6178);
or U6735 (N_6735,N_6442,N_6249);
nand U6736 (N_6736,N_6123,N_6103);
or U6737 (N_6737,N_6172,N_6040);
nor U6738 (N_6738,N_6274,N_6008);
and U6739 (N_6739,N_6138,N_6461);
or U6740 (N_6740,N_6219,N_6029);
and U6741 (N_6741,N_6157,N_6321);
nor U6742 (N_6742,N_6243,N_6397);
or U6743 (N_6743,N_6317,N_6136);
and U6744 (N_6744,N_6341,N_6401);
and U6745 (N_6745,N_6105,N_6269);
or U6746 (N_6746,N_6258,N_6006);
nor U6747 (N_6747,N_6083,N_6091);
or U6748 (N_6748,N_6020,N_6320);
or U6749 (N_6749,N_6075,N_6484);
nand U6750 (N_6750,N_6328,N_6134);
nor U6751 (N_6751,N_6455,N_6380);
and U6752 (N_6752,N_6395,N_6169);
nand U6753 (N_6753,N_6209,N_6357);
and U6754 (N_6754,N_6422,N_6151);
or U6755 (N_6755,N_6446,N_6343);
nand U6756 (N_6756,N_6420,N_6244);
nand U6757 (N_6757,N_6091,N_6184);
and U6758 (N_6758,N_6412,N_6040);
xor U6759 (N_6759,N_6330,N_6255);
nand U6760 (N_6760,N_6428,N_6055);
nor U6761 (N_6761,N_6422,N_6015);
and U6762 (N_6762,N_6471,N_6314);
or U6763 (N_6763,N_6266,N_6271);
xor U6764 (N_6764,N_6438,N_6016);
and U6765 (N_6765,N_6244,N_6455);
nor U6766 (N_6766,N_6040,N_6487);
or U6767 (N_6767,N_6142,N_6067);
and U6768 (N_6768,N_6018,N_6336);
or U6769 (N_6769,N_6425,N_6066);
nand U6770 (N_6770,N_6152,N_6340);
nor U6771 (N_6771,N_6338,N_6195);
nand U6772 (N_6772,N_6396,N_6114);
nor U6773 (N_6773,N_6119,N_6458);
nor U6774 (N_6774,N_6249,N_6416);
and U6775 (N_6775,N_6100,N_6154);
or U6776 (N_6776,N_6015,N_6303);
and U6777 (N_6777,N_6209,N_6428);
nand U6778 (N_6778,N_6275,N_6224);
nand U6779 (N_6779,N_6425,N_6390);
nand U6780 (N_6780,N_6033,N_6168);
nor U6781 (N_6781,N_6067,N_6475);
nor U6782 (N_6782,N_6044,N_6226);
or U6783 (N_6783,N_6447,N_6284);
xnor U6784 (N_6784,N_6117,N_6356);
and U6785 (N_6785,N_6224,N_6240);
and U6786 (N_6786,N_6260,N_6083);
nor U6787 (N_6787,N_6072,N_6492);
nor U6788 (N_6788,N_6232,N_6135);
nand U6789 (N_6789,N_6208,N_6342);
nand U6790 (N_6790,N_6042,N_6292);
xnor U6791 (N_6791,N_6103,N_6073);
and U6792 (N_6792,N_6157,N_6220);
or U6793 (N_6793,N_6233,N_6190);
nand U6794 (N_6794,N_6250,N_6344);
nand U6795 (N_6795,N_6119,N_6005);
or U6796 (N_6796,N_6178,N_6483);
nor U6797 (N_6797,N_6321,N_6147);
nand U6798 (N_6798,N_6314,N_6202);
or U6799 (N_6799,N_6427,N_6136);
xnor U6800 (N_6800,N_6177,N_6446);
nor U6801 (N_6801,N_6247,N_6456);
xnor U6802 (N_6802,N_6139,N_6204);
or U6803 (N_6803,N_6424,N_6026);
or U6804 (N_6804,N_6006,N_6293);
nor U6805 (N_6805,N_6084,N_6352);
and U6806 (N_6806,N_6416,N_6289);
nor U6807 (N_6807,N_6387,N_6439);
or U6808 (N_6808,N_6467,N_6448);
and U6809 (N_6809,N_6447,N_6285);
and U6810 (N_6810,N_6287,N_6324);
nand U6811 (N_6811,N_6210,N_6142);
and U6812 (N_6812,N_6281,N_6118);
or U6813 (N_6813,N_6348,N_6386);
or U6814 (N_6814,N_6225,N_6409);
nor U6815 (N_6815,N_6248,N_6404);
or U6816 (N_6816,N_6004,N_6095);
and U6817 (N_6817,N_6127,N_6477);
or U6818 (N_6818,N_6326,N_6298);
nand U6819 (N_6819,N_6077,N_6273);
nand U6820 (N_6820,N_6054,N_6482);
nor U6821 (N_6821,N_6081,N_6027);
xnor U6822 (N_6822,N_6181,N_6225);
and U6823 (N_6823,N_6129,N_6428);
and U6824 (N_6824,N_6177,N_6094);
or U6825 (N_6825,N_6212,N_6021);
nand U6826 (N_6826,N_6117,N_6352);
and U6827 (N_6827,N_6288,N_6162);
nand U6828 (N_6828,N_6046,N_6297);
or U6829 (N_6829,N_6434,N_6275);
nor U6830 (N_6830,N_6370,N_6377);
or U6831 (N_6831,N_6196,N_6252);
or U6832 (N_6832,N_6398,N_6048);
and U6833 (N_6833,N_6092,N_6422);
or U6834 (N_6834,N_6215,N_6316);
or U6835 (N_6835,N_6486,N_6342);
and U6836 (N_6836,N_6452,N_6461);
nand U6837 (N_6837,N_6018,N_6132);
nand U6838 (N_6838,N_6376,N_6098);
and U6839 (N_6839,N_6370,N_6072);
and U6840 (N_6840,N_6089,N_6386);
xnor U6841 (N_6841,N_6251,N_6377);
nand U6842 (N_6842,N_6039,N_6147);
and U6843 (N_6843,N_6126,N_6159);
nand U6844 (N_6844,N_6478,N_6086);
nor U6845 (N_6845,N_6340,N_6266);
and U6846 (N_6846,N_6403,N_6448);
or U6847 (N_6847,N_6235,N_6226);
nand U6848 (N_6848,N_6367,N_6157);
nor U6849 (N_6849,N_6144,N_6132);
and U6850 (N_6850,N_6224,N_6439);
nor U6851 (N_6851,N_6194,N_6378);
and U6852 (N_6852,N_6009,N_6265);
and U6853 (N_6853,N_6456,N_6081);
or U6854 (N_6854,N_6090,N_6459);
or U6855 (N_6855,N_6114,N_6458);
nor U6856 (N_6856,N_6420,N_6424);
and U6857 (N_6857,N_6182,N_6106);
or U6858 (N_6858,N_6418,N_6283);
nand U6859 (N_6859,N_6279,N_6467);
nor U6860 (N_6860,N_6259,N_6415);
or U6861 (N_6861,N_6290,N_6330);
nand U6862 (N_6862,N_6319,N_6167);
and U6863 (N_6863,N_6448,N_6312);
nor U6864 (N_6864,N_6109,N_6284);
nand U6865 (N_6865,N_6300,N_6052);
nor U6866 (N_6866,N_6112,N_6127);
or U6867 (N_6867,N_6211,N_6098);
or U6868 (N_6868,N_6478,N_6321);
and U6869 (N_6869,N_6358,N_6330);
nor U6870 (N_6870,N_6277,N_6242);
and U6871 (N_6871,N_6481,N_6227);
nand U6872 (N_6872,N_6295,N_6033);
nor U6873 (N_6873,N_6427,N_6045);
nand U6874 (N_6874,N_6421,N_6467);
nand U6875 (N_6875,N_6231,N_6261);
nor U6876 (N_6876,N_6375,N_6213);
nor U6877 (N_6877,N_6381,N_6450);
nand U6878 (N_6878,N_6476,N_6404);
nor U6879 (N_6879,N_6099,N_6293);
or U6880 (N_6880,N_6164,N_6065);
nor U6881 (N_6881,N_6081,N_6115);
or U6882 (N_6882,N_6151,N_6407);
and U6883 (N_6883,N_6368,N_6458);
or U6884 (N_6884,N_6401,N_6180);
nand U6885 (N_6885,N_6266,N_6455);
nor U6886 (N_6886,N_6483,N_6489);
and U6887 (N_6887,N_6126,N_6083);
nand U6888 (N_6888,N_6040,N_6430);
or U6889 (N_6889,N_6149,N_6155);
nor U6890 (N_6890,N_6288,N_6181);
and U6891 (N_6891,N_6433,N_6174);
nand U6892 (N_6892,N_6087,N_6021);
and U6893 (N_6893,N_6016,N_6172);
and U6894 (N_6894,N_6288,N_6447);
nand U6895 (N_6895,N_6023,N_6241);
nand U6896 (N_6896,N_6412,N_6028);
nand U6897 (N_6897,N_6094,N_6040);
nand U6898 (N_6898,N_6354,N_6269);
nor U6899 (N_6899,N_6329,N_6004);
nand U6900 (N_6900,N_6063,N_6489);
nand U6901 (N_6901,N_6069,N_6106);
or U6902 (N_6902,N_6047,N_6304);
and U6903 (N_6903,N_6082,N_6043);
nand U6904 (N_6904,N_6205,N_6226);
and U6905 (N_6905,N_6271,N_6395);
and U6906 (N_6906,N_6420,N_6181);
or U6907 (N_6907,N_6480,N_6437);
and U6908 (N_6908,N_6228,N_6173);
nand U6909 (N_6909,N_6057,N_6313);
or U6910 (N_6910,N_6005,N_6381);
and U6911 (N_6911,N_6374,N_6479);
nor U6912 (N_6912,N_6356,N_6225);
nor U6913 (N_6913,N_6277,N_6456);
nor U6914 (N_6914,N_6498,N_6452);
or U6915 (N_6915,N_6043,N_6404);
and U6916 (N_6916,N_6455,N_6104);
nand U6917 (N_6917,N_6404,N_6255);
or U6918 (N_6918,N_6346,N_6024);
xnor U6919 (N_6919,N_6348,N_6476);
nand U6920 (N_6920,N_6058,N_6051);
or U6921 (N_6921,N_6401,N_6361);
nand U6922 (N_6922,N_6003,N_6008);
and U6923 (N_6923,N_6315,N_6133);
or U6924 (N_6924,N_6449,N_6493);
or U6925 (N_6925,N_6016,N_6073);
or U6926 (N_6926,N_6211,N_6150);
nor U6927 (N_6927,N_6255,N_6270);
and U6928 (N_6928,N_6347,N_6284);
nor U6929 (N_6929,N_6250,N_6254);
nand U6930 (N_6930,N_6492,N_6374);
nor U6931 (N_6931,N_6225,N_6379);
nor U6932 (N_6932,N_6427,N_6017);
and U6933 (N_6933,N_6015,N_6411);
or U6934 (N_6934,N_6245,N_6105);
and U6935 (N_6935,N_6165,N_6382);
nor U6936 (N_6936,N_6363,N_6020);
nand U6937 (N_6937,N_6127,N_6393);
or U6938 (N_6938,N_6360,N_6331);
or U6939 (N_6939,N_6240,N_6423);
or U6940 (N_6940,N_6353,N_6383);
nor U6941 (N_6941,N_6319,N_6195);
nor U6942 (N_6942,N_6433,N_6066);
or U6943 (N_6943,N_6393,N_6475);
or U6944 (N_6944,N_6304,N_6456);
or U6945 (N_6945,N_6036,N_6171);
and U6946 (N_6946,N_6392,N_6498);
or U6947 (N_6947,N_6276,N_6463);
and U6948 (N_6948,N_6326,N_6006);
or U6949 (N_6949,N_6406,N_6362);
and U6950 (N_6950,N_6338,N_6125);
and U6951 (N_6951,N_6374,N_6071);
nand U6952 (N_6952,N_6389,N_6248);
or U6953 (N_6953,N_6427,N_6012);
or U6954 (N_6954,N_6366,N_6226);
nand U6955 (N_6955,N_6221,N_6398);
or U6956 (N_6956,N_6360,N_6196);
nor U6957 (N_6957,N_6305,N_6133);
nor U6958 (N_6958,N_6030,N_6188);
nor U6959 (N_6959,N_6319,N_6267);
nor U6960 (N_6960,N_6290,N_6075);
nor U6961 (N_6961,N_6027,N_6413);
and U6962 (N_6962,N_6209,N_6309);
nand U6963 (N_6963,N_6482,N_6081);
nor U6964 (N_6964,N_6384,N_6478);
or U6965 (N_6965,N_6039,N_6019);
nor U6966 (N_6966,N_6280,N_6153);
or U6967 (N_6967,N_6334,N_6096);
nand U6968 (N_6968,N_6049,N_6449);
nand U6969 (N_6969,N_6404,N_6100);
and U6970 (N_6970,N_6112,N_6167);
and U6971 (N_6971,N_6283,N_6298);
nor U6972 (N_6972,N_6180,N_6492);
and U6973 (N_6973,N_6316,N_6074);
nor U6974 (N_6974,N_6039,N_6276);
or U6975 (N_6975,N_6455,N_6130);
nor U6976 (N_6976,N_6486,N_6427);
nand U6977 (N_6977,N_6416,N_6323);
or U6978 (N_6978,N_6312,N_6349);
or U6979 (N_6979,N_6380,N_6279);
or U6980 (N_6980,N_6315,N_6121);
or U6981 (N_6981,N_6127,N_6470);
and U6982 (N_6982,N_6125,N_6071);
nand U6983 (N_6983,N_6210,N_6094);
or U6984 (N_6984,N_6324,N_6260);
and U6985 (N_6985,N_6464,N_6143);
or U6986 (N_6986,N_6304,N_6406);
xor U6987 (N_6987,N_6351,N_6465);
and U6988 (N_6988,N_6049,N_6431);
or U6989 (N_6989,N_6329,N_6041);
or U6990 (N_6990,N_6495,N_6100);
or U6991 (N_6991,N_6427,N_6470);
nor U6992 (N_6992,N_6489,N_6391);
and U6993 (N_6993,N_6416,N_6457);
and U6994 (N_6994,N_6271,N_6127);
nand U6995 (N_6995,N_6042,N_6492);
and U6996 (N_6996,N_6079,N_6480);
nor U6997 (N_6997,N_6490,N_6200);
nand U6998 (N_6998,N_6483,N_6139);
nor U6999 (N_6999,N_6231,N_6433);
nor U7000 (N_7000,N_6783,N_6767);
or U7001 (N_7001,N_6661,N_6785);
nand U7002 (N_7002,N_6800,N_6920);
nor U7003 (N_7003,N_6521,N_6636);
nand U7004 (N_7004,N_6778,N_6958);
nand U7005 (N_7005,N_6674,N_6982);
or U7006 (N_7006,N_6504,N_6930);
nand U7007 (N_7007,N_6516,N_6538);
or U7008 (N_7008,N_6536,N_6608);
or U7009 (N_7009,N_6730,N_6720);
nand U7010 (N_7010,N_6946,N_6860);
and U7011 (N_7011,N_6959,N_6562);
xor U7012 (N_7012,N_6534,N_6977);
nor U7013 (N_7013,N_6786,N_6653);
nor U7014 (N_7014,N_6518,N_6769);
nand U7015 (N_7015,N_6847,N_6671);
and U7016 (N_7016,N_6500,N_6856);
nor U7017 (N_7017,N_6693,N_6704);
nor U7018 (N_7018,N_6590,N_6810);
nor U7019 (N_7019,N_6918,N_6954);
nand U7020 (N_7020,N_6923,N_6502);
and U7021 (N_7021,N_6995,N_6528);
xor U7022 (N_7022,N_6570,N_6972);
and U7023 (N_7023,N_6573,N_6666);
nor U7024 (N_7024,N_6823,N_6551);
nor U7025 (N_7025,N_6875,N_6939);
nor U7026 (N_7026,N_6619,N_6578);
xnor U7027 (N_7027,N_6659,N_6780);
and U7028 (N_7028,N_6895,N_6808);
or U7029 (N_7029,N_6522,N_6899);
and U7030 (N_7030,N_6701,N_6511);
or U7031 (N_7031,N_6848,N_6526);
and U7032 (N_7032,N_6634,N_6821);
or U7033 (N_7033,N_6706,N_6533);
nand U7034 (N_7034,N_6503,N_6906);
or U7035 (N_7035,N_6621,N_6952);
and U7036 (N_7036,N_6664,N_6736);
nand U7037 (N_7037,N_6603,N_6809);
nor U7038 (N_7038,N_6685,N_6622);
nand U7039 (N_7039,N_6903,N_6631);
or U7040 (N_7040,N_6639,N_6794);
or U7041 (N_7041,N_6609,N_6645);
or U7042 (N_7042,N_6680,N_6650);
or U7043 (N_7043,N_6566,N_6612);
and U7044 (N_7044,N_6712,N_6556);
nor U7045 (N_7045,N_6512,N_6589);
nand U7046 (N_7046,N_6579,N_6826);
nand U7047 (N_7047,N_6961,N_6886);
nor U7048 (N_7048,N_6818,N_6527);
or U7049 (N_7049,N_6673,N_6668);
nor U7050 (N_7050,N_6655,N_6694);
nand U7051 (N_7051,N_6925,N_6561);
nand U7052 (N_7052,N_6625,N_6870);
nor U7053 (N_7053,N_6738,N_6864);
or U7054 (N_7054,N_6565,N_6648);
nor U7055 (N_7055,N_6907,N_6599);
or U7056 (N_7056,N_6586,N_6803);
or U7057 (N_7057,N_6568,N_6768);
nand U7058 (N_7058,N_6862,N_6820);
or U7059 (N_7059,N_6732,N_6756);
nor U7060 (N_7060,N_6688,N_6937);
and U7061 (N_7061,N_6797,N_6830);
or U7062 (N_7062,N_6684,N_6601);
and U7063 (N_7063,N_6900,N_6980);
or U7064 (N_7064,N_6658,N_6515);
nor U7065 (N_7065,N_6764,N_6564);
nor U7066 (N_7066,N_6971,N_6981);
nor U7067 (N_7067,N_6838,N_6577);
nor U7068 (N_7068,N_6944,N_6874);
nor U7069 (N_7069,N_6908,N_6513);
nor U7070 (N_7070,N_6540,N_6716);
nor U7071 (N_7071,N_6752,N_6993);
and U7072 (N_7072,N_6611,N_6950);
nand U7073 (N_7073,N_6921,N_6559);
nor U7074 (N_7074,N_6751,N_6596);
or U7075 (N_7075,N_6530,N_6727);
or U7076 (N_7076,N_6916,N_6824);
nand U7077 (N_7077,N_6678,N_6731);
and U7078 (N_7078,N_6772,N_6807);
nor U7079 (N_7079,N_6748,N_6990);
or U7080 (N_7080,N_6884,N_6994);
nand U7081 (N_7081,N_6850,N_6805);
nand U7082 (N_7082,N_6859,N_6949);
nand U7083 (N_7083,N_6537,N_6894);
nand U7084 (N_7084,N_6877,N_6633);
nand U7085 (N_7085,N_6798,N_6852);
nor U7086 (N_7086,N_6630,N_6888);
nand U7087 (N_7087,N_6962,N_6983);
or U7088 (N_7088,N_6729,N_6989);
or U7089 (N_7089,N_6933,N_6984);
or U7090 (N_7090,N_6531,N_6607);
nand U7091 (N_7091,N_6876,N_6617);
or U7092 (N_7092,N_6893,N_6539);
nand U7093 (N_7093,N_6686,N_6905);
and U7094 (N_7094,N_6588,N_6721);
and U7095 (N_7095,N_6594,N_6996);
and U7096 (N_7096,N_6979,N_6763);
or U7097 (N_7097,N_6861,N_6765);
nor U7098 (N_7098,N_6691,N_6822);
or U7099 (N_7099,N_6714,N_6718);
and U7100 (N_7100,N_6828,N_6835);
or U7101 (N_7101,N_6928,N_6687);
or U7102 (N_7102,N_6887,N_6911);
and U7103 (N_7103,N_6670,N_6932);
nor U7104 (N_7104,N_6519,N_6508);
nor U7105 (N_7105,N_6739,N_6827);
nor U7106 (N_7106,N_6642,N_6753);
or U7107 (N_7107,N_6967,N_6717);
nand U7108 (N_7108,N_6935,N_6806);
nor U7109 (N_7109,N_6700,N_6858);
or U7110 (N_7110,N_6855,N_6947);
nor U7111 (N_7111,N_6627,N_6974);
nand U7112 (N_7112,N_6628,N_6544);
or U7113 (N_7113,N_6705,N_6616);
or U7114 (N_7114,N_6572,N_6575);
nand U7115 (N_7115,N_6698,N_6624);
nor U7116 (N_7116,N_6968,N_6535);
nand U7117 (N_7117,N_6901,N_6523);
and U7118 (N_7118,N_6784,N_6652);
nand U7119 (N_7119,N_6943,N_6604);
nor U7120 (N_7120,N_6872,N_6941);
or U7121 (N_7121,N_6675,N_6690);
or U7122 (N_7122,N_6992,N_6591);
nor U7123 (N_7123,N_6615,N_6597);
or U7124 (N_7124,N_6574,N_6743);
or U7125 (N_7125,N_6987,N_6999);
nor U7126 (N_7126,N_6646,N_6940);
or U7127 (N_7127,N_6529,N_6600);
and U7128 (N_7128,N_6563,N_6744);
nor U7129 (N_7129,N_6737,N_6867);
nor U7130 (N_7130,N_6879,N_6790);
and U7131 (N_7131,N_6724,N_6632);
or U7132 (N_7132,N_6558,N_6834);
and U7133 (N_7133,N_6567,N_6524);
nand U7134 (N_7134,N_6929,N_6878);
nor U7135 (N_7135,N_6552,N_6931);
or U7136 (N_7136,N_6733,N_6587);
nand U7137 (N_7137,N_6773,N_6750);
and U7138 (N_7138,N_6913,N_6505);
nand U7139 (N_7139,N_6814,N_6985);
nand U7140 (N_7140,N_6761,N_6677);
xnor U7141 (N_7141,N_6865,N_6917);
nand U7142 (N_7142,N_6897,N_6719);
nor U7143 (N_7143,N_6676,N_6910);
and U7144 (N_7144,N_6667,N_6965);
and U7145 (N_7145,N_6902,N_6734);
nor U7146 (N_7146,N_6606,N_6635);
nor U7147 (N_7147,N_6991,N_6507);
or U7148 (N_7148,N_6963,N_6747);
or U7149 (N_7149,N_6699,N_6833);
or U7150 (N_7150,N_6610,N_6711);
nand U7151 (N_7151,N_6919,N_6640);
nand U7152 (N_7152,N_6846,N_6843);
and U7153 (N_7153,N_6546,N_6509);
or U7154 (N_7154,N_6592,N_6759);
and U7155 (N_7155,N_6757,N_6754);
nor U7156 (N_7156,N_6945,N_6726);
and U7157 (N_7157,N_6569,N_6789);
and U7158 (N_7158,N_6660,N_6804);
or U7159 (N_7159,N_6857,N_6626);
nand U7160 (N_7160,N_6681,N_6922);
nand U7161 (N_7161,N_6960,N_6829);
or U7162 (N_7162,N_6793,N_6755);
and U7163 (N_7163,N_6880,N_6514);
and U7164 (N_7164,N_6543,N_6882);
nand U7165 (N_7165,N_6782,N_6863);
or U7166 (N_7166,N_6851,N_6555);
nand U7167 (N_7167,N_6813,N_6695);
nand U7168 (N_7168,N_6742,N_6657);
or U7169 (N_7169,N_6844,N_6836);
and U7170 (N_7170,N_6970,N_6973);
and U7171 (N_7171,N_6576,N_6598);
nor U7172 (N_7172,N_6868,N_6614);
or U7173 (N_7173,N_6741,N_6898);
nor U7174 (N_7174,N_6595,N_6715);
or U7175 (N_7175,N_6934,N_6663);
and U7176 (N_7176,N_6689,N_6891);
nand U7177 (N_7177,N_6506,N_6795);
nand U7178 (N_7178,N_6618,N_6998);
nand U7179 (N_7179,N_6771,N_6722);
and U7180 (N_7180,N_6707,N_6871);
and U7181 (N_7181,N_6777,N_6550);
or U7182 (N_7182,N_6584,N_6745);
nor U7183 (N_7183,N_6957,N_6560);
nand U7184 (N_7184,N_6866,N_6580);
nor U7185 (N_7185,N_6669,N_6740);
nor U7186 (N_7186,N_6787,N_6762);
or U7187 (N_7187,N_6926,N_6581);
nand U7188 (N_7188,N_6812,N_6881);
nand U7189 (N_7189,N_6770,N_6904);
and U7190 (N_7190,N_6637,N_6620);
nand U7191 (N_7191,N_6953,N_6702);
nand U7192 (N_7192,N_6924,N_6840);
and U7193 (N_7193,N_6725,N_6710);
or U7194 (N_7194,N_6713,N_6890);
nor U7195 (N_7195,N_6746,N_6542);
and U7196 (N_7196,N_6912,N_6679);
nand U7197 (N_7197,N_6966,N_6938);
or U7198 (N_7198,N_6708,N_6760);
and U7199 (N_7199,N_6656,N_6779);
or U7200 (N_7200,N_6697,N_6885);
nand U7201 (N_7201,N_6819,N_6781);
and U7202 (N_7202,N_6796,N_6582);
or U7203 (N_7203,N_6969,N_6896);
or U7204 (N_7204,N_6571,N_6816);
nor U7205 (N_7205,N_6703,N_6849);
or U7206 (N_7206,N_6692,N_6914);
and U7207 (N_7207,N_6585,N_6892);
or U7208 (N_7208,N_6986,N_6510);
or U7209 (N_7209,N_6825,N_6915);
xor U7210 (N_7210,N_6869,N_6651);
and U7211 (N_7211,N_6682,N_6517);
nor U7212 (N_7212,N_6665,N_6853);
and U7213 (N_7213,N_6520,N_6776);
nand U7214 (N_7214,N_6647,N_6775);
and U7215 (N_7215,N_6815,N_6709);
xor U7216 (N_7216,N_6811,N_6501);
xor U7217 (N_7217,N_6723,N_6641);
or U7218 (N_7218,N_6801,N_6735);
and U7219 (N_7219,N_6791,N_6774);
or U7220 (N_7220,N_6758,N_6942);
nand U7221 (N_7221,N_6605,N_6654);
and U7222 (N_7222,N_6978,N_6553);
and U7223 (N_7223,N_6644,N_6557);
and U7224 (N_7224,N_6927,N_6951);
nand U7225 (N_7225,N_6831,N_6788);
nand U7226 (N_7226,N_6547,N_6841);
or U7227 (N_7227,N_6873,N_6976);
xor U7228 (N_7228,N_6975,N_6948);
nor U7229 (N_7229,N_6593,N_6548);
and U7230 (N_7230,N_6988,N_6955);
nor U7231 (N_7231,N_6792,N_6638);
or U7232 (N_7232,N_6683,N_6696);
nand U7233 (N_7233,N_6845,N_6997);
nand U7234 (N_7234,N_6909,N_6649);
nor U7235 (N_7235,N_6549,N_6541);
or U7236 (N_7236,N_6956,N_6936);
or U7237 (N_7237,N_6629,N_6532);
or U7238 (N_7238,N_6525,N_6766);
nand U7239 (N_7239,N_6623,N_6545);
nor U7240 (N_7240,N_6643,N_6554);
nand U7241 (N_7241,N_6662,N_6839);
and U7242 (N_7242,N_6602,N_6749);
nor U7243 (N_7243,N_6583,N_6802);
or U7244 (N_7244,N_6964,N_6728);
or U7245 (N_7245,N_6842,N_6817);
nand U7246 (N_7246,N_6837,N_6883);
or U7247 (N_7247,N_6799,N_6832);
and U7248 (N_7248,N_6889,N_6613);
xor U7249 (N_7249,N_6672,N_6854);
or U7250 (N_7250,N_6752,N_6664);
or U7251 (N_7251,N_6608,N_6712);
nor U7252 (N_7252,N_6883,N_6699);
nand U7253 (N_7253,N_6732,N_6770);
nand U7254 (N_7254,N_6845,N_6996);
and U7255 (N_7255,N_6996,N_6840);
or U7256 (N_7256,N_6886,N_6766);
or U7257 (N_7257,N_6865,N_6847);
or U7258 (N_7258,N_6518,N_6893);
nor U7259 (N_7259,N_6586,N_6544);
or U7260 (N_7260,N_6522,N_6610);
or U7261 (N_7261,N_6715,N_6681);
nor U7262 (N_7262,N_6893,N_6788);
nand U7263 (N_7263,N_6799,N_6642);
or U7264 (N_7264,N_6948,N_6605);
and U7265 (N_7265,N_6909,N_6818);
and U7266 (N_7266,N_6635,N_6579);
nand U7267 (N_7267,N_6990,N_6926);
and U7268 (N_7268,N_6710,N_6778);
xor U7269 (N_7269,N_6956,N_6972);
or U7270 (N_7270,N_6973,N_6753);
and U7271 (N_7271,N_6852,N_6598);
nand U7272 (N_7272,N_6773,N_6617);
and U7273 (N_7273,N_6888,N_6884);
nor U7274 (N_7274,N_6737,N_6967);
nand U7275 (N_7275,N_6717,N_6718);
nor U7276 (N_7276,N_6900,N_6783);
and U7277 (N_7277,N_6736,N_6713);
nand U7278 (N_7278,N_6731,N_6540);
nand U7279 (N_7279,N_6958,N_6980);
or U7280 (N_7280,N_6866,N_6520);
and U7281 (N_7281,N_6774,N_6969);
and U7282 (N_7282,N_6989,N_6623);
nor U7283 (N_7283,N_6908,N_6763);
and U7284 (N_7284,N_6992,N_6514);
and U7285 (N_7285,N_6688,N_6716);
nor U7286 (N_7286,N_6784,N_6785);
nor U7287 (N_7287,N_6798,N_6867);
nand U7288 (N_7288,N_6546,N_6575);
nor U7289 (N_7289,N_6912,N_6837);
or U7290 (N_7290,N_6928,N_6607);
and U7291 (N_7291,N_6753,N_6541);
nor U7292 (N_7292,N_6535,N_6869);
and U7293 (N_7293,N_6520,N_6743);
or U7294 (N_7294,N_6549,N_6698);
and U7295 (N_7295,N_6828,N_6750);
nand U7296 (N_7296,N_6807,N_6538);
nor U7297 (N_7297,N_6714,N_6793);
nand U7298 (N_7298,N_6738,N_6566);
and U7299 (N_7299,N_6802,N_6629);
or U7300 (N_7300,N_6840,N_6630);
nor U7301 (N_7301,N_6857,N_6605);
or U7302 (N_7302,N_6759,N_6819);
and U7303 (N_7303,N_6756,N_6714);
xor U7304 (N_7304,N_6706,N_6914);
and U7305 (N_7305,N_6659,N_6586);
nand U7306 (N_7306,N_6929,N_6980);
or U7307 (N_7307,N_6649,N_6762);
or U7308 (N_7308,N_6871,N_6954);
or U7309 (N_7309,N_6673,N_6754);
nand U7310 (N_7310,N_6501,N_6833);
nor U7311 (N_7311,N_6951,N_6556);
and U7312 (N_7312,N_6527,N_6613);
or U7313 (N_7313,N_6724,N_6703);
nor U7314 (N_7314,N_6759,N_6556);
and U7315 (N_7315,N_6571,N_6681);
nand U7316 (N_7316,N_6571,N_6848);
nand U7317 (N_7317,N_6586,N_6796);
nor U7318 (N_7318,N_6624,N_6709);
nand U7319 (N_7319,N_6654,N_6556);
nor U7320 (N_7320,N_6511,N_6564);
and U7321 (N_7321,N_6537,N_6548);
nor U7322 (N_7322,N_6992,N_6596);
and U7323 (N_7323,N_6849,N_6890);
and U7324 (N_7324,N_6739,N_6747);
and U7325 (N_7325,N_6688,N_6546);
nor U7326 (N_7326,N_6766,N_6573);
and U7327 (N_7327,N_6650,N_6559);
or U7328 (N_7328,N_6901,N_6938);
nand U7329 (N_7329,N_6905,N_6910);
and U7330 (N_7330,N_6842,N_6500);
or U7331 (N_7331,N_6536,N_6617);
nor U7332 (N_7332,N_6813,N_6660);
nand U7333 (N_7333,N_6789,N_6872);
nand U7334 (N_7334,N_6865,N_6715);
nor U7335 (N_7335,N_6669,N_6653);
nand U7336 (N_7336,N_6524,N_6955);
or U7337 (N_7337,N_6646,N_6820);
and U7338 (N_7338,N_6622,N_6654);
or U7339 (N_7339,N_6641,N_6867);
nand U7340 (N_7340,N_6966,N_6723);
or U7341 (N_7341,N_6818,N_6843);
or U7342 (N_7342,N_6619,N_6710);
nor U7343 (N_7343,N_6697,N_6898);
and U7344 (N_7344,N_6654,N_6779);
or U7345 (N_7345,N_6727,N_6793);
nand U7346 (N_7346,N_6989,N_6526);
nor U7347 (N_7347,N_6995,N_6843);
or U7348 (N_7348,N_6662,N_6933);
or U7349 (N_7349,N_6531,N_6881);
and U7350 (N_7350,N_6746,N_6769);
nand U7351 (N_7351,N_6758,N_6999);
nor U7352 (N_7352,N_6675,N_6930);
and U7353 (N_7353,N_6902,N_6855);
or U7354 (N_7354,N_6557,N_6545);
or U7355 (N_7355,N_6863,N_6661);
nor U7356 (N_7356,N_6959,N_6609);
nor U7357 (N_7357,N_6661,N_6749);
nand U7358 (N_7358,N_6861,N_6615);
nor U7359 (N_7359,N_6750,N_6786);
nor U7360 (N_7360,N_6835,N_6879);
nor U7361 (N_7361,N_6831,N_6791);
nor U7362 (N_7362,N_6532,N_6577);
or U7363 (N_7363,N_6784,N_6978);
nor U7364 (N_7364,N_6937,N_6857);
nand U7365 (N_7365,N_6893,N_6723);
or U7366 (N_7366,N_6567,N_6919);
or U7367 (N_7367,N_6676,N_6909);
nand U7368 (N_7368,N_6849,N_6671);
nor U7369 (N_7369,N_6604,N_6618);
nor U7370 (N_7370,N_6875,N_6836);
nor U7371 (N_7371,N_6576,N_6790);
nor U7372 (N_7372,N_6609,N_6723);
and U7373 (N_7373,N_6821,N_6791);
nor U7374 (N_7374,N_6545,N_6692);
and U7375 (N_7375,N_6859,N_6602);
nor U7376 (N_7376,N_6726,N_6716);
and U7377 (N_7377,N_6779,N_6722);
nand U7378 (N_7378,N_6972,N_6807);
nand U7379 (N_7379,N_6680,N_6544);
nand U7380 (N_7380,N_6704,N_6641);
and U7381 (N_7381,N_6524,N_6678);
nor U7382 (N_7382,N_6814,N_6766);
nand U7383 (N_7383,N_6579,N_6521);
nand U7384 (N_7384,N_6694,N_6519);
nor U7385 (N_7385,N_6807,N_6784);
and U7386 (N_7386,N_6645,N_6814);
and U7387 (N_7387,N_6938,N_6624);
nand U7388 (N_7388,N_6914,N_6788);
or U7389 (N_7389,N_6563,N_6990);
nand U7390 (N_7390,N_6551,N_6610);
or U7391 (N_7391,N_6786,N_6979);
nor U7392 (N_7392,N_6941,N_6822);
and U7393 (N_7393,N_6694,N_6960);
or U7394 (N_7394,N_6974,N_6980);
nor U7395 (N_7395,N_6934,N_6839);
nor U7396 (N_7396,N_6538,N_6737);
and U7397 (N_7397,N_6543,N_6787);
nor U7398 (N_7398,N_6696,N_6998);
xnor U7399 (N_7399,N_6852,N_6941);
nor U7400 (N_7400,N_6536,N_6589);
or U7401 (N_7401,N_6747,N_6814);
nand U7402 (N_7402,N_6990,N_6968);
xor U7403 (N_7403,N_6794,N_6916);
nor U7404 (N_7404,N_6918,N_6881);
nand U7405 (N_7405,N_6836,N_6508);
or U7406 (N_7406,N_6559,N_6826);
or U7407 (N_7407,N_6633,N_6661);
and U7408 (N_7408,N_6874,N_6922);
nand U7409 (N_7409,N_6917,N_6881);
or U7410 (N_7410,N_6575,N_6930);
and U7411 (N_7411,N_6775,N_6619);
or U7412 (N_7412,N_6896,N_6794);
or U7413 (N_7413,N_6973,N_6962);
or U7414 (N_7414,N_6807,N_6557);
nand U7415 (N_7415,N_6902,N_6762);
nand U7416 (N_7416,N_6974,N_6554);
and U7417 (N_7417,N_6967,N_6977);
or U7418 (N_7418,N_6538,N_6596);
or U7419 (N_7419,N_6700,N_6795);
nand U7420 (N_7420,N_6828,N_6909);
or U7421 (N_7421,N_6873,N_6981);
or U7422 (N_7422,N_6632,N_6676);
nand U7423 (N_7423,N_6961,N_6887);
nor U7424 (N_7424,N_6732,N_6584);
nand U7425 (N_7425,N_6643,N_6966);
nor U7426 (N_7426,N_6631,N_6766);
nor U7427 (N_7427,N_6507,N_6949);
nand U7428 (N_7428,N_6883,N_6919);
nor U7429 (N_7429,N_6957,N_6826);
xor U7430 (N_7430,N_6919,N_6774);
xnor U7431 (N_7431,N_6838,N_6762);
and U7432 (N_7432,N_6507,N_6966);
nor U7433 (N_7433,N_6930,N_6800);
nand U7434 (N_7434,N_6860,N_6552);
nand U7435 (N_7435,N_6988,N_6922);
nor U7436 (N_7436,N_6697,N_6979);
xnor U7437 (N_7437,N_6702,N_6921);
nand U7438 (N_7438,N_6763,N_6910);
and U7439 (N_7439,N_6847,N_6537);
and U7440 (N_7440,N_6760,N_6983);
xor U7441 (N_7441,N_6731,N_6641);
and U7442 (N_7442,N_6961,N_6761);
nand U7443 (N_7443,N_6970,N_6637);
nand U7444 (N_7444,N_6824,N_6874);
nor U7445 (N_7445,N_6746,N_6975);
or U7446 (N_7446,N_6644,N_6684);
nand U7447 (N_7447,N_6500,N_6501);
nor U7448 (N_7448,N_6969,N_6636);
nand U7449 (N_7449,N_6953,N_6740);
and U7450 (N_7450,N_6693,N_6954);
or U7451 (N_7451,N_6512,N_6877);
nor U7452 (N_7452,N_6535,N_6698);
and U7453 (N_7453,N_6749,N_6897);
nand U7454 (N_7454,N_6905,N_6901);
or U7455 (N_7455,N_6840,N_6613);
nor U7456 (N_7456,N_6869,N_6679);
or U7457 (N_7457,N_6518,N_6666);
nor U7458 (N_7458,N_6914,N_6665);
and U7459 (N_7459,N_6671,N_6631);
nand U7460 (N_7460,N_6681,N_6669);
nor U7461 (N_7461,N_6787,N_6720);
nand U7462 (N_7462,N_6509,N_6724);
or U7463 (N_7463,N_6872,N_6969);
or U7464 (N_7464,N_6994,N_6629);
nor U7465 (N_7465,N_6636,N_6613);
or U7466 (N_7466,N_6560,N_6726);
and U7467 (N_7467,N_6876,N_6910);
nand U7468 (N_7468,N_6710,N_6868);
nor U7469 (N_7469,N_6703,N_6825);
nor U7470 (N_7470,N_6593,N_6873);
nor U7471 (N_7471,N_6751,N_6817);
nand U7472 (N_7472,N_6845,N_6802);
nand U7473 (N_7473,N_6772,N_6680);
and U7474 (N_7474,N_6846,N_6848);
and U7475 (N_7475,N_6813,N_6996);
nand U7476 (N_7476,N_6778,N_6782);
and U7477 (N_7477,N_6808,N_6856);
or U7478 (N_7478,N_6872,N_6834);
nor U7479 (N_7479,N_6758,N_6523);
or U7480 (N_7480,N_6810,N_6762);
or U7481 (N_7481,N_6763,N_6983);
or U7482 (N_7482,N_6691,N_6510);
nor U7483 (N_7483,N_6511,N_6957);
nor U7484 (N_7484,N_6597,N_6927);
or U7485 (N_7485,N_6906,N_6598);
nand U7486 (N_7486,N_6940,N_6848);
nand U7487 (N_7487,N_6768,N_6742);
nand U7488 (N_7488,N_6956,N_6670);
nand U7489 (N_7489,N_6828,N_6855);
xor U7490 (N_7490,N_6673,N_6519);
nor U7491 (N_7491,N_6897,N_6698);
nand U7492 (N_7492,N_6954,N_6605);
nor U7493 (N_7493,N_6800,N_6632);
nand U7494 (N_7494,N_6969,N_6638);
nand U7495 (N_7495,N_6956,N_6807);
and U7496 (N_7496,N_6660,N_6674);
nand U7497 (N_7497,N_6896,N_6997);
nor U7498 (N_7498,N_6648,N_6593);
nand U7499 (N_7499,N_6704,N_6646);
and U7500 (N_7500,N_7499,N_7004);
or U7501 (N_7501,N_7204,N_7296);
nor U7502 (N_7502,N_7130,N_7227);
and U7503 (N_7503,N_7370,N_7025);
or U7504 (N_7504,N_7372,N_7440);
nand U7505 (N_7505,N_7171,N_7097);
or U7506 (N_7506,N_7143,N_7389);
or U7507 (N_7507,N_7154,N_7173);
and U7508 (N_7508,N_7123,N_7045);
xnor U7509 (N_7509,N_7148,N_7387);
nand U7510 (N_7510,N_7246,N_7139);
or U7511 (N_7511,N_7495,N_7304);
nor U7512 (N_7512,N_7210,N_7396);
or U7513 (N_7513,N_7144,N_7053);
or U7514 (N_7514,N_7132,N_7454);
and U7515 (N_7515,N_7366,N_7032);
nand U7516 (N_7516,N_7422,N_7429);
nand U7517 (N_7517,N_7490,N_7088);
nor U7518 (N_7518,N_7466,N_7287);
nor U7519 (N_7519,N_7080,N_7207);
and U7520 (N_7520,N_7340,N_7375);
and U7521 (N_7521,N_7437,N_7086);
or U7522 (N_7522,N_7243,N_7250);
and U7523 (N_7523,N_7193,N_7410);
nor U7524 (N_7524,N_7234,N_7024);
or U7525 (N_7525,N_7232,N_7344);
and U7526 (N_7526,N_7455,N_7463);
nand U7527 (N_7527,N_7464,N_7073);
and U7528 (N_7528,N_7049,N_7009);
and U7529 (N_7529,N_7050,N_7117);
or U7530 (N_7530,N_7245,N_7394);
or U7531 (N_7531,N_7493,N_7260);
nor U7532 (N_7532,N_7069,N_7488);
nor U7533 (N_7533,N_7472,N_7252);
nand U7534 (N_7534,N_7022,N_7128);
nand U7535 (N_7535,N_7044,N_7236);
nand U7536 (N_7536,N_7182,N_7155);
nor U7537 (N_7537,N_7431,N_7308);
or U7538 (N_7538,N_7156,N_7424);
nand U7539 (N_7539,N_7197,N_7332);
or U7540 (N_7540,N_7483,N_7160);
nor U7541 (N_7541,N_7191,N_7075);
and U7542 (N_7542,N_7180,N_7238);
or U7543 (N_7543,N_7200,N_7166);
xnor U7544 (N_7544,N_7247,N_7381);
nand U7545 (N_7545,N_7237,N_7406);
nor U7546 (N_7546,N_7041,N_7063);
nor U7547 (N_7547,N_7167,N_7138);
xor U7548 (N_7548,N_7275,N_7416);
nand U7549 (N_7549,N_7333,N_7081);
nand U7550 (N_7550,N_7470,N_7468);
nand U7551 (N_7551,N_7496,N_7494);
nand U7552 (N_7552,N_7293,N_7030);
nor U7553 (N_7553,N_7355,N_7071);
and U7554 (N_7554,N_7048,N_7265);
nor U7555 (N_7555,N_7159,N_7354);
or U7556 (N_7556,N_7165,N_7388);
or U7557 (N_7557,N_7125,N_7395);
nor U7558 (N_7558,N_7404,N_7039);
nor U7559 (N_7559,N_7017,N_7435);
or U7560 (N_7560,N_7486,N_7013);
nand U7561 (N_7561,N_7262,N_7445);
nor U7562 (N_7562,N_7432,N_7299);
nor U7563 (N_7563,N_7038,N_7145);
nor U7564 (N_7564,N_7335,N_7297);
or U7565 (N_7565,N_7442,N_7391);
and U7566 (N_7566,N_7402,N_7096);
or U7567 (N_7567,N_7283,N_7256);
nand U7568 (N_7568,N_7428,N_7359);
or U7569 (N_7569,N_7360,N_7220);
and U7570 (N_7570,N_7228,N_7035);
nor U7571 (N_7571,N_7398,N_7356);
nand U7572 (N_7572,N_7303,N_7415);
or U7573 (N_7573,N_7007,N_7336);
or U7574 (N_7574,N_7380,N_7112);
nor U7575 (N_7575,N_7010,N_7043);
and U7576 (N_7576,N_7040,N_7068);
nor U7577 (N_7577,N_7272,N_7461);
nand U7578 (N_7578,N_7240,N_7401);
or U7579 (N_7579,N_7327,N_7076);
or U7580 (N_7580,N_7438,N_7479);
nor U7581 (N_7581,N_7326,N_7474);
nor U7582 (N_7582,N_7294,N_7364);
or U7583 (N_7583,N_7177,N_7201);
or U7584 (N_7584,N_7309,N_7315);
nand U7585 (N_7585,N_7295,N_7104);
nor U7586 (N_7586,N_7456,N_7184);
and U7587 (N_7587,N_7292,N_7186);
and U7588 (N_7588,N_7267,N_7343);
nand U7589 (N_7589,N_7122,N_7083);
and U7590 (N_7590,N_7168,N_7115);
and U7591 (N_7591,N_7286,N_7060);
nor U7592 (N_7592,N_7259,N_7172);
and U7593 (N_7593,N_7430,N_7385);
nand U7594 (N_7594,N_7106,N_7378);
nand U7595 (N_7595,N_7093,N_7280);
or U7596 (N_7596,N_7005,N_7042);
nand U7597 (N_7597,N_7188,N_7176);
or U7598 (N_7598,N_7189,N_7379);
nor U7599 (N_7599,N_7199,N_7498);
nand U7600 (N_7600,N_7313,N_7065);
nor U7601 (N_7601,N_7091,N_7345);
nand U7602 (N_7602,N_7175,N_7214);
or U7603 (N_7603,N_7151,N_7229);
nor U7604 (N_7604,N_7119,N_7383);
nor U7605 (N_7605,N_7459,N_7405);
or U7606 (N_7606,N_7001,N_7181);
and U7607 (N_7607,N_7449,N_7021);
nor U7608 (N_7608,N_7301,N_7027);
nand U7609 (N_7609,N_7031,N_7157);
or U7610 (N_7610,N_7342,N_7258);
nor U7611 (N_7611,N_7377,N_7161);
nor U7612 (N_7612,N_7358,N_7061);
and U7613 (N_7613,N_7028,N_7105);
xnor U7614 (N_7614,N_7290,N_7318);
nand U7615 (N_7615,N_7098,N_7215);
nor U7616 (N_7616,N_7339,N_7357);
or U7617 (N_7617,N_7298,N_7158);
nand U7618 (N_7618,N_7121,N_7102);
or U7619 (N_7619,N_7368,N_7000);
nor U7620 (N_7620,N_7420,N_7090);
and U7621 (N_7621,N_7037,N_7099);
and U7622 (N_7622,N_7064,N_7338);
and U7623 (N_7623,N_7433,N_7450);
nand U7624 (N_7624,N_7150,N_7101);
or U7625 (N_7625,N_7153,N_7311);
nor U7626 (N_7626,N_7020,N_7059);
or U7627 (N_7627,N_7261,N_7427);
nand U7628 (N_7628,N_7140,N_7439);
and U7629 (N_7629,N_7403,N_7003);
nor U7630 (N_7630,N_7334,N_7120);
or U7631 (N_7631,N_7070,N_7414);
nor U7632 (N_7632,N_7263,N_7255);
nor U7633 (N_7633,N_7163,N_7118);
or U7634 (N_7634,N_7284,N_7419);
nand U7635 (N_7635,N_7230,N_7477);
or U7636 (N_7636,N_7219,N_7094);
and U7637 (N_7637,N_7058,N_7471);
and U7638 (N_7638,N_7397,N_7476);
nor U7639 (N_7639,N_7282,N_7462);
and U7640 (N_7640,N_7131,N_7408);
nor U7641 (N_7641,N_7480,N_7187);
and U7642 (N_7642,N_7264,N_7085);
or U7643 (N_7643,N_7142,N_7051);
or U7644 (N_7644,N_7217,N_7253);
and U7645 (N_7645,N_7487,N_7390);
nor U7646 (N_7646,N_7162,N_7257);
or U7647 (N_7647,N_7341,N_7347);
nor U7648 (N_7648,N_7209,N_7235);
nor U7649 (N_7649,N_7135,N_7089);
or U7650 (N_7650,N_7337,N_7015);
nand U7651 (N_7651,N_7178,N_7224);
or U7652 (N_7652,N_7108,N_7113);
and U7653 (N_7653,N_7475,N_7393);
nand U7654 (N_7654,N_7348,N_7221);
or U7655 (N_7655,N_7465,N_7497);
nor U7656 (N_7656,N_7374,N_7399);
and U7657 (N_7657,N_7023,N_7268);
nor U7658 (N_7658,N_7141,N_7029);
or U7659 (N_7659,N_7183,N_7062);
nor U7660 (N_7660,N_7026,N_7376);
or U7661 (N_7661,N_7249,N_7254);
nor U7662 (N_7662,N_7458,N_7452);
nand U7663 (N_7663,N_7006,N_7129);
nand U7664 (N_7664,N_7231,N_7034);
nand U7665 (N_7665,N_7473,N_7111);
or U7666 (N_7666,N_7285,N_7306);
nand U7667 (N_7667,N_7077,N_7169);
or U7668 (N_7668,N_7087,N_7136);
or U7669 (N_7669,N_7434,N_7446);
and U7670 (N_7670,N_7222,N_7242);
nand U7671 (N_7671,N_7484,N_7353);
xor U7672 (N_7672,N_7164,N_7351);
nor U7673 (N_7673,N_7444,N_7382);
or U7674 (N_7674,N_7016,N_7270);
or U7675 (N_7675,N_7008,N_7448);
nor U7676 (N_7676,N_7365,N_7481);
and U7677 (N_7677,N_7320,N_7216);
and U7678 (N_7678,N_7205,N_7198);
or U7679 (N_7679,N_7491,N_7057);
nand U7680 (N_7680,N_7319,N_7047);
or U7681 (N_7681,N_7269,N_7443);
nand U7682 (N_7682,N_7072,N_7248);
nor U7683 (N_7683,N_7328,N_7478);
xor U7684 (N_7684,N_7469,N_7302);
and U7685 (N_7685,N_7194,N_7190);
and U7686 (N_7686,N_7244,N_7185);
or U7687 (N_7687,N_7307,N_7114);
or U7688 (N_7688,N_7067,N_7084);
or U7689 (N_7689,N_7300,N_7352);
or U7690 (N_7690,N_7100,N_7124);
nand U7691 (N_7691,N_7133,N_7195);
nand U7692 (N_7692,N_7134,N_7149);
nand U7693 (N_7693,N_7288,N_7281);
nor U7694 (N_7694,N_7251,N_7409);
nand U7695 (N_7695,N_7271,N_7453);
nor U7696 (N_7696,N_7277,N_7426);
or U7697 (N_7697,N_7324,N_7485);
or U7698 (N_7698,N_7384,N_7109);
nand U7699 (N_7699,N_7279,N_7202);
or U7700 (N_7700,N_7137,N_7146);
and U7701 (N_7701,N_7233,N_7460);
xnor U7702 (N_7702,N_7012,N_7386);
and U7703 (N_7703,N_7033,N_7436);
and U7704 (N_7704,N_7110,N_7467);
and U7705 (N_7705,N_7011,N_7482);
or U7706 (N_7706,N_7095,N_7126);
nor U7707 (N_7707,N_7441,N_7349);
and U7708 (N_7708,N_7014,N_7079);
nor U7709 (N_7709,N_7329,N_7363);
and U7710 (N_7710,N_7451,N_7196);
and U7711 (N_7711,N_7425,N_7066);
nand U7712 (N_7712,N_7211,N_7489);
nand U7713 (N_7713,N_7417,N_7322);
or U7714 (N_7714,N_7179,N_7019);
or U7715 (N_7715,N_7413,N_7103);
or U7716 (N_7716,N_7170,N_7316);
nor U7717 (N_7717,N_7423,N_7331);
nor U7718 (N_7718,N_7407,N_7447);
nand U7719 (N_7719,N_7321,N_7362);
and U7720 (N_7720,N_7213,N_7457);
or U7721 (N_7721,N_7367,N_7078);
and U7722 (N_7722,N_7092,N_7412);
nor U7723 (N_7723,N_7056,N_7036);
xnor U7724 (N_7724,N_7274,N_7273);
nor U7725 (N_7725,N_7174,N_7371);
nand U7726 (N_7726,N_7074,N_7203);
nand U7727 (N_7727,N_7278,N_7223);
or U7728 (N_7728,N_7369,N_7107);
nor U7729 (N_7729,N_7373,N_7310);
nand U7730 (N_7730,N_7400,N_7392);
nand U7731 (N_7731,N_7225,N_7239);
nor U7732 (N_7732,N_7218,N_7192);
nand U7733 (N_7733,N_7325,N_7346);
and U7734 (N_7734,N_7266,N_7116);
nand U7735 (N_7735,N_7147,N_7330);
nand U7736 (N_7736,N_7082,N_7350);
xor U7737 (N_7737,N_7276,N_7127);
or U7738 (N_7738,N_7055,N_7411);
or U7739 (N_7739,N_7054,N_7241);
and U7740 (N_7740,N_7291,N_7212);
nand U7741 (N_7741,N_7018,N_7312);
and U7742 (N_7742,N_7206,N_7152);
or U7743 (N_7743,N_7046,N_7492);
and U7744 (N_7744,N_7314,N_7289);
nor U7745 (N_7745,N_7421,N_7323);
nand U7746 (N_7746,N_7052,N_7418);
nand U7747 (N_7747,N_7002,N_7208);
nor U7748 (N_7748,N_7317,N_7226);
or U7749 (N_7749,N_7305,N_7361);
nor U7750 (N_7750,N_7482,N_7094);
nor U7751 (N_7751,N_7079,N_7004);
and U7752 (N_7752,N_7067,N_7344);
and U7753 (N_7753,N_7106,N_7050);
or U7754 (N_7754,N_7266,N_7185);
and U7755 (N_7755,N_7423,N_7270);
nor U7756 (N_7756,N_7348,N_7403);
nand U7757 (N_7757,N_7399,N_7427);
or U7758 (N_7758,N_7007,N_7385);
nor U7759 (N_7759,N_7004,N_7194);
or U7760 (N_7760,N_7170,N_7346);
nor U7761 (N_7761,N_7402,N_7039);
nand U7762 (N_7762,N_7352,N_7138);
nand U7763 (N_7763,N_7129,N_7355);
and U7764 (N_7764,N_7250,N_7120);
nor U7765 (N_7765,N_7084,N_7322);
nand U7766 (N_7766,N_7229,N_7160);
and U7767 (N_7767,N_7390,N_7090);
nor U7768 (N_7768,N_7386,N_7414);
nor U7769 (N_7769,N_7172,N_7342);
nor U7770 (N_7770,N_7476,N_7289);
nor U7771 (N_7771,N_7086,N_7104);
nand U7772 (N_7772,N_7216,N_7120);
nor U7773 (N_7773,N_7134,N_7083);
nor U7774 (N_7774,N_7174,N_7343);
or U7775 (N_7775,N_7498,N_7230);
nand U7776 (N_7776,N_7007,N_7004);
xor U7777 (N_7777,N_7301,N_7297);
and U7778 (N_7778,N_7032,N_7080);
nand U7779 (N_7779,N_7466,N_7481);
nand U7780 (N_7780,N_7061,N_7144);
or U7781 (N_7781,N_7249,N_7043);
and U7782 (N_7782,N_7462,N_7148);
xor U7783 (N_7783,N_7034,N_7234);
or U7784 (N_7784,N_7110,N_7388);
nor U7785 (N_7785,N_7325,N_7363);
or U7786 (N_7786,N_7187,N_7483);
and U7787 (N_7787,N_7429,N_7327);
nor U7788 (N_7788,N_7342,N_7430);
and U7789 (N_7789,N_7116,N_7083);
and U7790 (N_7790,N_7107,N_7153);
and U7791 (N_7791,N_7114,N_7065);
or U7792 (N_7792,N_7466,N_7096);
nand U7793 (N_7793,N_7405,N_7155);
or U7794 (N_7794,N_7061,N_7492);
nor U7795 (N_7795,N_7194,N_7075);
or U7796 (N_7796,N_7481,N_7002);
and U7797 (N_7797,N_7437,N_7029);
nand U7798 (N_7798,N_7385,N_7480);
or U7799 (N_7799,N_7244,N_7183);
nor U7800 (N_7800,N_7277,N_7030);
nand U7801 (N_7801,N_7388,N_7407);
nand U7802 (N_7802,N_7016,N_7039);
and U7803 (N_7803,N_7375,N_7035);
xnor U7804 (N_7804,N_7035,N_7219);
or U7805 (N_7805,N_7383,N_7406);
and U7806 (N_7806,N_7127,N_7204);
nor U7807 (N_7807,N_7119,N_7484);
and U7808 (N_7808,N_7405,N_7343);
xnor U7809 (N_7809,N_7033,N_7081);
nand U7810 (N_7810,N_7224,N_7196);
and U7811 (N_7811,N_7218,N_7012);
and U7812 (N_7812,N_7352,N_7485);
nor U7813 (N_7813,N_7172,N_7272);
or U7814 (N_7814,N_7435,N_7306);
xor U7815 (N_7815,N_7365,N_7115);
or U7816 (N_7816,N_7111,N_7125);
nor U7817 (N_7817,N_7457,N_7368);
and U7818 (N_7818,N_7146,N_7288);
and U7819 (N_7819,N_7144,N_7151);
or U7820 (N_7820,N_7371,N_7057);
and U7821 (N_7821,N_7195,N_7429);
nor U7822 (N_7822,N_7290,N_7282);
nor U7823 (N_7823,N_7119,N_7303);
nor U7824 (N_7824,N_7268,N_7294);
and U7825 (N_7825,N_7183,N_7102);
or U7826 (N_7826,N_7155,N_7252);
or U7827 (N_7827,N_7376,N_7269);
nand U7828 (N_7828,N_7173,N_7013);
or U7829 (N_7829,N_7391,N_7256);
or U7830 (N_7830,N_7103,N_7312);
and U7831 (N_7831,N_7050,N_7127);
and U7832 (N_7832,N_7419,N_7268);
and U7833 (N_7833,N_7354,N_7257);
nor U7834 (N_7834,N_7286,N_7434);
nor U7835 (N_7835,N_7182,N_7129);
and U7836 (N_7836,N_7404,N_7119);
or U7837 (N_7837,N_7383,N_7386);
and U7838 (N_7838,N_7492,N_7248);
nand U7839 (N_7839,N_7084,N_7047);
and U7840 (N_7840,N_7466,N_7315);
or U7841 (N_7841,N_7210,N_7358);
or U7842 (N_7842,N_7280,N_7216);
and U7843 (N_7843,N_7482,N_7091);
nand U7844 (N_7844,N_7034,N_7495);
or U7845 (N_7845,N_7163,N_7498);
or U7846 (N_7846,N_7365,N_7394);
and U7847 (N_7847,N_7216,N_7195);
and U7848 (N_7848,N_7356,N_7336);
or U7849 (N_7849,N_7049,N_7439);
or U7850 (N_7850,N_7177,N_7078);
nand U7851 (N_7851,N_7298,N_7165);
nor U7852 (N_7852,N_7333,N_7238);
nor U7853 (N_7853,N_7162,N_7347);
nor U7854 (N_7854,N_7280,N_7361);
or U7855 (N_7855,N_7110,N_7412);
or U7856 (N_7856,N_7257,N_7366);
or U7857 (N_7857,N_7043,N_7374);
nand U7858 (N_7858,N_7436,N_7410);
or U7859 (N_7859,N_7354,N_7274);
nand U7860 (N_7860,N_7119,N_7485);
nand U7861 (N_7861,N_7152,N_7174);
nand U7862 (N_7862,N_7017,N_7474);
or U7863 (N_7863,N_7276,N_7390);
and U7864 (N_7864,N_7322,N_7213);
nor U7865 (N_7865,N_7226,N_7095);
or U7866 (N_7866,N_7130,N_7421);
or U7867 (N_7867,N_7082,N_7447);
nand U7868 (N_7868,N_7155,N_7415);
nor U7869 (N_7869,N_7110,N_7332);
nor U7870 (N_7870,N_7448,N_7005);
and U7871 (N_7871,N_7266,N_7383);
or U7872 (N_7872,N_7127,N_7196);
and U7873 (N_7873,N_7231,N_7428);
or U7874 (N_7874,N_7003,N_7181);
nand U7875 (N_7875,N_7246,N_7429);
and U7876 (N_7876,N_7042,N_7279);
nand U7877 (N_7877,N_7148,N_7433);
and U7878 (N_7878,N_7379,N_7322);
and U7879 (N_7879,N_7293,N_7237);
nor U7880 (N_7880,N_7046,N_7429);
and U7881 (N_7881,N_7221,N_7134);
nand U7882 (N_7882,N_7456,N_7219);
nor U7883 (N_7883,N_7163,N_7253);
and U7884 (N_7884,N_7308,N_7456);
and U7885 (N_7885,N_7259,N_7295);
and U7886 (N_7886,N_7456,N_7268);
nand U7887 (N_7887,N_7382,N_7411);
nand U7888 (N_7888,N_7444,N_7352);
or U7889 (N_7889,N_7240,N_7197);
nand U7890 (N_7890,N_7308,N_7131);
nand U7891 (N_7891,N_7389,N_7163);
nand U7892 (N_7892,N_7021,N_7314);
or U7893 (N_7893,N_7388,N_7397);
and U7894 (N_7894,N_7209,N_7103);
nor U7895 (N_7895,N_7137,N_7049);
nor U7896 (N_7896,N_7335,N_7334);
and U7897 (N_7897,N_7156,N_7140);
nand U7898 (N_7898,N_7363,N_7164);
nand U7899 (N_7899,N_7452,N_7023);
or U7900 (N_7900,N_7089,N_7308);
and U7901 (N_7901,N_7304,N_7312);
nand U7902 (N_7902,N_7439,N_7114);
nor U7903 (N_7903,N_7396,N_7194);
and U7904 (N_7904,N_7283,N_7320);
nand U7905 (N_7905,N_7421,N_7194);
nor U7906 (N_7906,N_7031,N_7400);
nor U7907 (N_7907,N_7477,N_7381);
and U7908 (N_7908,N_7395,N_7258);
or U7909 (N_7909,N_7306,N_7413);
nand U7910 (N_7910,N_7099,N_7026);
or U7911 (N_7911,N_7221,N_7409);
and U7912 (N_7912,N_7116,N_7171);
or U7913 (N_7913,N_7421,N_7398);
nand U7914 (N_7914,N_7133,N_7176);
and U7915 (N_7915,N_7429,N_7347);
nor U7916 (N_7916,N_7225,N_7028);
nand U7917 (N_7917,N_7448,N_7055);
nand U7918 (N_7918,N_7381,N_7228);
nor U7919 (N_7919,N_7209,N_7202);
nor U7920 (N_7920,N_7022,N_7463);
nor U7921 (N_7921,N_7146,N_7083);
and U7922 (N_7922,N_7001,N_7352);
or U7923 (N_7923,N_7259,N_7049);
nor U7924 (N_7924,N_7091,N_7318);
and U7925 (N_7925,N_7369,N_7404);
nand U7926 (N_7926,N_7448,N_7175);
nand U7927 (N_7927,N_7388,N_7157);
and U7928 (N_7928,N_7152,N_7267);
nand U7929 (N_7929,N_7011,N_7154);
and U7930 (N_7930,N_7346,N_7185);
or U7931 (N_7931,N_7428,N_7170);
or U7932 (N_7932,N_7237,N_7093);
nor U7933 (N_7933,N_7022,N_7263);
nor U7934 (N_7934,N_7343,N_7076);
or U7935 (N_7935,N_7193,N_7021);
and U7936 (N_7936,N_7458,N_7202);
nor U7937 (N_7937,N_7345,N_7030);
nand U7938 (N_7938,N_7016,N_7346);
and U7939 (N_7939,N_7323,N_7257);
nor U7940 (N_7940,N_7200,N_7486);
nand U7941 (N_7941,N_7243,N_7418);
and U7942 (N_7942,N_7234,N_7009);
or U7943 (N_7943,N_7425,N_7207);
nor U7944 (N_7944,N_7405,N_7189);
and U7945 (N_7945,N_7034,N_7325);
nor U7946 (N_7946,N_7460,N_7324);
or U7947 (N_7947,N_7136,N_7282);
and U7948 (N_7948,N_7120,N_7111);
nand U7949 (N_7949,N_7151,N_7426);
nand U7950 (N_7950,N_7482,N_7361);
nand U7951 (N_7951,N_7205,N_7162);
or U7952 (N_7952,N_7430,N_7003);
nand U7953 (N_7953,N_7144,N_7098);
nor U7954 (N_7954,N_7348,N_7274);
or U7955 (N_7955,N_7428,N_7382);
nor U7956 (N_7956,N_7098,N_7119);
nand U7957 (N_7957,N_7488,N_7018);
nand U7958 (N_7958,N_7413,N_7029);
and U7959 (N_7959,N_7213,N_7374);
nand U7960 (N_7960,N_7344,N_7147);
nand U7961 (N_7961,N_7448,N_7491);
nand U7962 (N_7962,N_7426,N_7043);
nor U7963 (N_7963,N_7366,N_7220);
and U7964 (N_7964,N_7130,N_7100);
and U7965 (N_7965,N_7076,N_7016);
nor U7966 (N_7966,N_7377,N_7395);
nand U7967 (N_7967,N_7159,N_7449);
nor U7968 (N_7968,N_7234,N_7426);
nor U7969 (N_7969,N_7110,N_7009);
nor U7970 (N_7970,N_7364,N_7457);
nand U7971 (N_7971,N_7295,N_7147);
or U7972 (N_7972,N_7394,N_7170);
nand U7973 (N_7973,N_7057,N_7186);
or U7974 (N_7974,N_7316,N_7273);
nor U7975 (N_7975,N_7497,N_7001);
and U7976 (N_7976,N_7040,N_7193);
or U7977 (N_7977,N_7324,N_7101);
nand U7978 (N_7978,N_7084,N_7412);
nor U7979 (N_7979,N_7336,N_7460);
nand U7980 (N_7980,N_7169,N_7061);
or U7981 (N_7981,N_7205,N_7334);
nand U7982 (N_7982,N_7433,N_7029);
nor U7983 (N_7983,N_7358,N_7064);
and U7984 (N_7984,N_7130,N_7064);
xnor U7985 (N_7985,N_7163,N_7151);
nand U7986 (N_7986,N_7205,N_7020);
nor U7987 (N_7987,N_7075,N_7447);
nand U7988 (N_7988,N_7194,N_7384);
and U7989 (N_7989,N_7328,N_7139);
nand U7990 (N_7990,N_7424,N_7361);
nor U7991 (N_7991,N_7099,N_7357);
nor U7992 (N_7992,N_7437,N_7054);
nor U7993 (N_7993,N_7478,N_7435);
nand U7994 (N_7994,N_7216,N_7292);
nand U7995 (N_7995,N_7345,N_7471);
nand U7996 (N_7996,N_7121,N_7078);
and U7997 (N_7997,N_7419,N_7239);
and U7998 (N_7998,N_7242,N_7023);
nor U7999 (N_7999,N_7194,N_7207);
and U8000 (N_8000,N_7713,N_7873);
nor U8001 (N_8001,N_7678,N_7703);
nand U8002 (N_8002,N_7983,N_7972);
and U8003 (N_8003,N_7854,N_7715);
or U8004 (N_8004,N_7980,N_7749);
nand U8005 (N_8005,N_7765,N_7672);
and U8006 (N_8006,N_7926,N_7824);
or U8007 (N_8007,N_7805,N_7698);
or U8008 (N_8008,N_7619,N_7843);
nor U8009 (N_8009,N_7901,N_7754);
or U8010 (N_8010,N_7668,N_7652);
xnor U8011 (N_8011,N_7740,N_7595);
nand U8012 (N_8012,N_7530,N_7918);
nand U8013 (N_8013,N_7578,N_7964);
nor U8014 (N_8014,N_7823,N_7669);
and U8015 (N_8015,N_7724,N_7945);
nor U8016 (N_8016,N_7597,N_7676);
nand U8017 (N_8017,N_7653,N_7838);
nand U8018 (N_8018,N_7666,N_7558);
nor U8019 (N_8019,N_7999,N_7991);
and U8020 (N_8020,N_7542,N_7527);
and U8021 (N_8021,N_7910,N_7984);
and U8022 (N_8022,N_7665,N_7704);
nand U8023 (N_8023,N_7756,N_7543);
nand U8024 (N_8024,N_7744,N_7536);
or U8025 (N_8025,N_7528,N_7580);
or U8026 (N_8026,N_7747,N_7859);
and U8027 (N_8027,N_7917,N_7898);
and U8028 (N_8028,N_7872,N_7952);
xor U8029 (N_8029,N_7990,N_7947);
nand U8030 (N_8030,N_7525,N_7708);
nand U8031 (N_8031,N_7658,N_7520);
nand U8032 (N_8032,N_7936,N_7940);
and U8033 (N_8033,N_7569,N_7887);
nand U8034 (N_8034,N_7988,N_7884);
nor U8035 (N_8035,N_7941,N_7553);
or U8036 (N_8036,N_7590,N_7966);
and U8037 (N_8037,N_7723,N_7976);
nor U8038 (N_8038,N_7701,N_7870);
and U8039 (N_8039,N_7899,N_7538);
or U8040 (N_8040,N_7506,N_7924);
nand U8041 (N_8041,N_7853,N_7637);
and U8042 (N_8042,N_7997,N_7505);
nand U8043 (N_8043,N_7565,N_7531);
nor U8044 (N_8044,N_7800,N_7829);
or U8045 (N_8045,N_7741,N_7803);
nor U8046 (N_8046,N_7864,N_7816);
or U8047 (N_8047,N_7627,N_7721);
or U8048 (N_8048,N_7534,N_7822);
nand U8049 (N_8049,N_7512,N_7532);
and U8050 (N_8050,N_7552,N_7742);
nand U8051 (N_8051,N_7697,N_7944);
and U8052 (N_8052,N_7635,N_7570);
xnor U8053 (N_8053,N_7612,N_7562);
or U8054 (N_8054,N_7850,N_7857);
nor U8055 (N_8055,N_7762,N_7959);
xnor U8056 (N_8056,N_7557,N_7774);
nor U8057 (N_8057,N_7559,N_7719);
xnor U8058 (N_8058,N_7641,N_7663);
or U8059 (N_8059,N_7705,N_7793);
nor U8060 (N_8060,N_7912,N_7833);
or U8061 (N_8061,N_7847,N_7700);
and U8062 (N_8062,N_7636,N_7706);
and U8063 (N_8063,N_7720,N_7819);
nand U8064 (N_8064,N_7882,N_7521);
and U8065 (N_8065,N_7778,N_7848);
nor U8066 (N_8066,N_7757,N_7596);
nor U8067 (N_8067,N_7993,N_7573);
and U8068 (N_8068,N_7875,N_7913);
or U8069 (N_8069,N_7759,N_7807);
nor U8070 (N_8070,N_7893,N_7503);
and U8071 (N_8071,N_7630,N_7651);
and U8072 (N_8072,N_7517,N_7809);
and U8073 (N_8073,N_7812,N_7709);
and U8074 (N_8074,N_7982,N_7548);
and U8075 (N_8075,N_7830,N_7588);
nand U8076 (N_8076,N_7968,N_7922);
nand U8077 (N_8077,N_7662,N_7902);
nor U8078 (N_8078,N_7608,N_7726);
or U8079 (N_8079,N_7603,N_7518);
and U8080 (N_8080,N_7842,N_7963);
nand U8081 (N_8081,N_7745,N_7656);
nand U8082 (N_8082,N_7804,N_7828);
nor U8083 (N_8083,N_7681,N_7802);
nor U8084 (N_8084,N_7736,N_7643);
or U8085 (N_8085,N_7632,N_7622);
and U8086 (N_8086,N_7634,N_7675);
nand U8087 (N_8087,N_7956,N_7693);
nand U8088 (N_8088,N_7743,N_7592);
and U8089 (N_8089,N_7863,N_7561);
xnor U8090 (N_8090,N_7826,N_7815);
and U8091 (N_8091,N_7871,N_7738);
nor U8092 (N_8092,N_7647,N_7722);
or U8093 (N_8093,N_7795,N_7714);
nor U8094 (N_8094,N_7585,N_7576);
or U8095 (N_8095,N_7909,N_7667);
nor U8096 (N_8096,N_7954,N_7685);
nor U8097 (N_8097,N_7609,N_7925);
nand U8098 (N_8098,N_7877,N_7549);
and U8099 (N_8099,N_7867,N_7849);
and U8100 (N_8100,N_7735,N_7514);
and U8101 (N_8101,N_7564,N_7885);
and U8102 (N_8102,N_7568,N_7914);
nor U8103 (N_8103,N_7511,N_7616);
nand U8104 (N_8104,N_7975,N_7832);
nand U8105 (N_8105,N_7670,N_7648);
and U8106 (N_8106,N_7510,N_7507);
nor U8107 (N_8107,N_7814,N_7679);
and U8108 (N_8108,N_7671,N_7661);
or U8109 (N_8109,N_7604,N_7868);
nor U8110 (N_8110,N_7862,N_7907);
nor U8111 (N_8111,N_7890,N_7911);
or U8112 (N_8112,N_7792,N_7973);
nor U8113 (N_8113,N_7813,N_7811);
nand U8114 (N_8114,N_7626,N_7979);
nor U8115 (N_8115,N_7948,N_7563);
nand U8116 (N_8116,N_7739,N_7801);
nand U8117 (N_8117,N_7889,N_7628);
or U8118 (N_8118,N_7779,N_7737);
and U8119 (N_8119,N_7657,N_7555);
nor U8120 (N_8120,N_7974,N_7645);
and U8121 (N_8121,N_7845,N_7965);
xnor U8122 (N_8122,N_7821,N_7934);
and U8123 (N_8123,N_7888,N_7606);
nor U8124 (N_8124,N_7664,N_7996);
nor U8125 (N_8125,N_7776,N_7760);
and U8126 (N_8126,N_7906,N_7961);
and U8127 (N_8127,N_7969,N_7770);
and U8128 (N_8128,N_7900,N_7939);
nor U8129 (N_8129,N_7998,N_7572);
and U8130 (N_8130,N_7921,N_7855);
nand U8131 (N_8131,N_7836,N_7683);
nand U8132 (N_8132,N_7994,N_7541);
and U8133 (N_8133,N_7691,N_7650);
and U8134 (N_8134,N_7610,N_7930);
nand U8135 (N_8135,N_7699,N_7727);
nor U8136 (N_8136,N_7688,N_7718);
nor U8137 (N_8137,N_7995,N_7958);
xor U8138 (N_8138,N_7625,N_7615);
nand U8139 (N_8139,N_7690,N_7971);
nor U8140 (N_8140,N_7858,N_7710);
xnor U8141 (N_8141,N_7547,N_7808);
nor U8142 (N_8142,N_7659,N_7750);
and U8143 (N_8143,N_7689,N_7574);
or U8144 (N_8144,N_7866,N_7611);
and U8145 (N_8145,N_7748,N_7755);
and U8146 (N_8146,N_7878,N_7831);
or U8147 (N_8147,N_7560,N_7687);
and U8148 (N_8148,N_7602,N_7777);
or U8149 (N_8149,N_7545,N_7860);
xnor U8150 (N_8150,N_7856,N_7927);
or U8151 (N_8151,N_7733,N_7942);
and U8152 (N_8152,N_7929,N_7501);
nand U8153 (N_8153,N_7519,N_7571);
nor U8154 (N_8154,N_7782,N_7682);
or U8155 (N_8155,N_7938,N_7876);
or U8156 (N_8156,N_7614,N_7624);
or U8157 (N_8157,N_7932,N_7581);
nand U8158 (N_8158,N_7618,N_7783);
or U8159 (N_8159,N_7977,N_7582);
nand U8160 (N_8160,N_7768,N_7992);
nand U8161 (N_8161,N_7785,N_7950);
and U8162 (N_8162,N_7605,N_7791);
or U8163 (N_8163,N_7607,N_7796);
or U8164 (N_8164,N_7551,N_7753);
nor U8165 (N_8165,N_7660,N_7915);
nor U8166 (N_8166,N_7920,N_7953);
or U8167 (N_8167,N_7673,N_7535);
and U8168 (N_8168,N_7970,N_7655);
and U8169 (N_8169,N_7707,N_7623);
and U8170 (N_8170,N_7841,N_7732);
nor U8171 (N_8171,N_7613,N_7781);
nor U8172 (N_8172,N_7931,N_7820);
nor U8173 (N_8173,N_7790,N_7654);
nor U8174 (N_8174,N_7515,N_7540);
and U8175 (N_8175,N_7787,N_7839);
nor U8176 (N_8176,N_7644,N_7799);
nor U8177 (N_8177,N_7694,N_7734);
or U8178 (N_8178,N_7784,N_7810);
or U8179 (N_8179,N_7594,N_7874);
and U8180 (N_8180,N_7702,N_7638);
nor U8181 (N_8181,N_7529,N_7758);
or U8182 (N_8182,N_7817,N_7646);
nor U8183 (N_8183,N_7516,N_7806);
or U8184 (N_8184,N_7794,N_7567);
and U8185 (N_8185,N_7579,N_7502);
nand U8186 (N_8186,N_7599,N_7846);
nand U8187 (N_8187,N_7881,N_7896);
and U8188 (N_8188,N_7513,N_7894);
nand U8189 (N_8189,N_7978,N_7851);
nor U8190 (N_8190,N_7767,N_7680);
xor U8191 (N_8191,N_7633,N_7771);
nor U8192 (N_8192,N_7526,N_7923);
or U8193 (N_8193,N_7711,N_7844);
and U8194 (N_8194,N_7798,N_7827);
or U8195 (N_8195,N_7903,N_7761);
nor U8196 (N_8196,N_7712,N_7835);
nor U8197 (N_8197,N_7642,N_7967);
or U8198 (N_8198,N_7601,N_7617);
nor U8199 (N_8199,N_7880,N_7600);
or U8200 (N_8200,N_7575,N_7752);
and U8201 (N_8201,N_7869,N_7746);
nand U8202 (N_8202,N_7897,N_7591);
and U8203 (N_8203,N_7508,N_7772);
nand U8204 (N_8204,N_7677,N_7621);
or U8205 (N_8205,N_7937,N_7554);
nand U8206 (N_8206,N_7905,N_7587);
nor U8207 (N_8207,N_7577,N_7593);
or U8208 (N_8208,N_7696,N_7861);
and U8209 (N_8209,N_7586,N_7537);
nand U8210 (N_8210,N_7686,N_7955);
and U8211 (N_8211,N_7523,N_7786);
nor U8212 (N_8212,N_7935,N_7544);
or U8213 (N_8213,N_7933,N_7522);
nor U8214 (N_8214,N_7943,N_7556);
nor U8215 (N_8215,N_7730,N_7631);
and U8216 (N_8216,N_7639,N_7766);
or U8217 (N_8217,N_7589,N_7957);
and U8218 (N_8218,N_7865,N_7960);
and U8219 (N_8219,N_7928,N_7629);
nor U8220 (N_8220,N_7725,N_7904);
or U8221 (N_8221,N_7729,N_7751);
or U8222 (N_8222,N_7916,N_7788);
or U8223 (N_8223,N_7852,N_7763);
xnor U8224 (N_8224,N_7775,N_7583);
or U8225 (N_8225,N_7598,N_7986);
and U8226 (N_8226,N_7908,N_7500);
nor U8227 (N_8227,N_7818,N_7731);
or U8228 (N_8228,N_7533,N_7692);
nand U8229 (N_8229,N_7509,N_7550);
nand U8230 (N_8230,N_7892,N_7883);
nand U8231 (N_8231,N_7797,N_7837);
xor U8232 (N_8232,N_7649,N_7769);
and U8233 (N_8233,N_7695,N_7891);
nor U8234 (N_8234,N_7620,N_7728);
and U8235 (N_8235,N_7780,N_7640);
and U8236 (N_8236,N_7895,N_7539);
and U8237 (N_8237,N_7716,N_7684);
or U8238 (N_8238,N_7825,N_7919);
nor U8239 (N_8239,N_7566,N_7951);
or U8240 (N_8240,N_7764,N_7879);
and U8241 (N_8241,N_7789,N_7840);
nand U8242 (N_8242,N_7834,N_7886);
or U8243 (N_8243,N_7962,N_7674);
nand U8244 (N_8244,N_7717,N_7985);
and U8245 (N_8245,N_7989,N_7546);
or U8246 (N_8246,N_7773,N_7946);
nand U8247 (N_8247,N_7524,N_7949);
or U8248 (N_8248,N_7504,N_7584);
nand U8249 (N_8249,N_7981,N_7987);
nand U8250 (N_8250,N_7640,N_7704);
or U8251 (N_8251,N_7811,N_7860);
xnor U8252 (N_8252,N_7665,N_7713);
and U8253 (N_8253,N_7805,N_7808);
nand U8254 (N_8254,N_7914,N_7533);
nor U8255 (N_8255,N_7759,N_7854);
or U8256 (N_8256,N_7597,N_7839);
and U8257 (N_8257,N_7907,N_7949);
and U8258 (N_8258,N_7566,N_7994);
and U8259 (N_8259,N_7660,N_7790);
xnor U8260 (N_8260,N_7845,N_7923);
nand U8261 (N_8261,N_7720,N_7860);
nand U8262 (N_8262,N_7830,N_7638);
nand U8263 (N_8263,N_7740,N_7801);
and U8264 (N_8264,N_7951,N_7523);
nor U8265 (N_8265,N_7906,N_7792);
or U8266 (N_8266,N_7979,N_7550);
xor U8267 (N_8267,N_7514,N_7651);
nand U8268 (N_8268,N_7930,N_7761);
nand U8269 (N_8269,N_7903,N_7608);
nor U8270 (N_8270,N_7504,N_7680);
nand U8271 (N_8271,N_7788,N_7693);
or U8272 (N_8272,N_7793,N_7660);
nand U8273 (N_8273,N_7992,N_7623);
nand U8274 (N_8274,N_7680,N_7812);
nand U8275 (N_8275,N_7996,N_7758);
nand U8276 (N_8276,N_7899,N_7529);
nor U8277 (N_8277,N_7973,N_7994);
nand U8278 (N_8278,N_7980,N_7934);
and U8279 (N_8279,N_7577,N_7862);
nor U8280 (N_8280,N_7554,N_7920);
nor U8281 (N_8281,N_7907,N_7977);
xor U8282 (N_8282,N_7508,N_7649);
nand U8283 (N_8283,N_7755,N_7574);
and U8284 (N_8284,N_7970,N_7966);
or U8285 (N_8285,N_7598,N_7713);
nand U8286 (N_8286,N_7759,N_7645);
and U8287 (N_8287,N_7818,N_7796);
nor U8288 (N_8288,N_7593,N_7679);
nand U8289 (N_8289,N_7913,N_7666);
nor U8290 (N_8290,N_7801,N_7946);
and U8291 (N_8291,N_7916,N_7691);
and U8292 (N_8292,N_7907,N_7844);
or U8293 (N_8293,N_7522,N_7824);
nor U8294 (N_8294,N_7771,N_7631);
and U8295 (N_8295,N_7658,N_7638);
nand U8296 (N_8296,N_7519,N_7767);
nand U8297 (N_8297,N_7569,N_7600);
and U8298 (N_8298,N_7806,N_7771);
or U8299 (N_8299,N_7955,N_7532);
or U8300 (N_8300,N_7580,N_7829);
or U8301 (N_8301,N_7572,N_7660);
or U8302 (N_8302,N_7531,N_7705);
nand U8303 (N_8303,N_7511,N_7850);
nand U8304 (N_8304,N_7768,N_7997);
or U8305 (N_8305,N_7784,N_7801);
nand U8306 (N_8306,N_7599,N_7682);
nor U8307 (N_8307,N_7759,N_7646);
and U8308 (N_8308,N_7967,N_7751);
nand U8309 (N_8309,N_7659,N_7901);
and U8310 (N_8310,N_7634,N_7583);
and U8311 (N_8311,N_7700,N_7623);
nand U8312 (N_8312,N_7537,N_7741);
or U8313 (N_8313,N_7968,N_7870);
and U8314 (N_8314,N_7687,N_7999);
and U8315 (N_8315,N_7723,N_7811);
or U8316 (N_8316,N_7508,N_7699);
nand U8317 (N_8317,N_7898,N_7861);
nand U8318 (N_8318,N_7998,N_7905);
or U8319 (N_8319,N_7831,N_7611);
nor U8320 (N_8320,N_7529,N_7520);
nor U8321 (N_8321,N_7769,N_7765);
and U8322 (N_8322,N_7688,N_7894);
or U8323 (N_8323,N_7632,N_7641);
and U8324 (N_8324,N_7604,N_7622);
nor U8325 (N_8325,N_7824,N_7516);
or U8326 (N_8326,N_7965,N_7663);
or U8327 (N_8327,N_7575,N_7642);
or U8328 (N_8328,N_7734,N_7569);
nand U8329 (N_8329,N_7914,N_7907);
nand U8330 (N_8330,N_7883,N_7915);
and U8331 (N_8331,N_7867,N_7814);
nand U8332 (N_8332,N_7843,N_7894);
and U8333 (N_8333,N_7750,N_7527);
or U8334 (N_8334,N_7746,N_7515);
and U8335 (N_8335,N_7925,N_7847);
and U8336 (N_8336,N_7918,N_7680);
and U8337 (N_8337,N_7974,N_7721);
or U8338 (N_8338,N_7507,N_7752);
nor U8339 (N_8339,N_7822,N_7725);
or U8340 (N_8340,N_7954,N_7836);
nand U8341 (N_8341,N_7625,N_7573);
or U8342 (N_8342,N_7882,N_7907);
nor U8343 (N_8343,N_7925,N_7905);
nor U8344 (N_8344,N_7937,N_7841);
or U8345 (N_8345,N_7652,N_7687);
and U8346 (N_8346,N_7936,N_7660);
or U8347 (N_8347,N_7673,N_7881);
and U8348 (N_8348,N_7699,N_7674);
nor U8349 (N_8349,N_7509,N_7895);
or U8350 (N_8350,N_7849,N_7823);
and U8351 (N_8351,N_7674,N_7597);
xnor U8352 (N_8352,N_7912,N_7940);
nor U8353 (N_8353,N_7744,N_7922);
nand U8354 (N_8354,N_7610,N_7541);
or U8355 (N_8355,N_7634,N_7978);
and U8356 (N_8356,N_7548,N_7555);
nand U8357 (N_8357,N_7906,N_7970);
and U8358 (N_8358,N_7510,N_7561);
and U8359 (N_8359,N_7932,N_7588);
or U8360 (N_8360,N_7520,N_7642);
nor U8361 (N_8361,N_7600,N_7649);
or U8362 (N_8362,N_7972,N_7657);
nor U8363 (N_8363,N_7761,N_7574);
nor U8364 (N_8364,N_7941,N_7661);
nand U8365 (N_8365,N_7802,N_7744);
or U8366 (N_8366,N_7979,N_7632);
and U8367 (N_8367,N_7625,N_7798);
and U8368 (N_8368,N_7715,N_7866);
nand U8369 (N_8369,N_7566,N_7749);
nand U8370 (N_8370,N_7661,N_7647);
and U8371 (N_8371,N_7581,N_7988);
and U8372 (N_8372,N_7640,N_7963);
nand U8373 (N_8373,N_7795,N_7542);
nor U8374 (N_8374,N_7959,N_7830);
and U8375 (N_8375,N_7651,N_7863);
or U8376 (N_8376,N_7795,N_7970);
nor U8377 (N_8377,N_7831,N_7702);
nand U8378 (N_8378,N_7762,N_7739);
nand U8379 (N_8379,N_7606,N_7590);
nor U8380 (N_8380,N_7827,N_7986);
nor U8381 (N_8381,N_7873,N_7600);
nor U8382 (N_8382,N_7723,N_7515);
and U8383 (N_8383,N_7579,N_7636);
nand U8384 (N_8384,N_7736,N_7569);
nor U8385 (N_8385,N_7790,N_7574);
nand U8386 (N_8386,N_7869,N_7909);
or U8387 (N_8387,N_7949,N_7811);
nor U8388 (N_8388,N_7954,N_7853);
or U8389 (N_8389,N_7976,N_7602);
nand U8390 (N_8390,N_7800,N_7562);
and U8391 (N_8391,N_7795,N_7685);
nand U8392 (N_8392,N_7851,N_7926);
and U8393 (N_8393,N_7768,N_7500);
nand U8394 (N_8394,N_7666,N_7774);
nand U8395 (N_8395,N_7790,N_7855);
and U8396 (N_8396,N_7887,N_7813);
nand U8397 (N_8397,N_7650,N_7811);
or U8398 (N_8398,N_7693,N_7856);
or U8399 (N_8399,N_7521,N_7848);
nand U8400 (N_8400,N_7853,N_7953);
and U8401 (N_8401,N_7682,N_7735);
nor U8402 (N_8402,N_7823,N_7798);
nand U8403 (N_8403,N_7746,N_7707);
or U8404 (N_8404,N_7741,N_7966);
or U8405 (N_8405,N_7902,N_7959);
xnor U8406 (N_8406,N_7565,N_7890);
nor U8407 (N_8407,N_7814,N_7747);
xor U8408 (N_8408,N_7805,N_7650);
nand U8409 (N_8409,N_7713,N_7699);
nand U8410 (N_8410,N_7811,N_7529);
or U8411 (N_8411,N_7777,N_7893);
and U8412 (N_8412,N_7660,N_7808);
nor U8413 (N_8413,N_7516,N_7801);
nor U8414 (N_8414,N_7923,N_7898);
and U8415 (N_8415,N_7764,N_7636);
nand U8416 (N_8416,N_7691,N_7757);
and U8417 (N_8417,N_7991,N_7736);
nor U8418 (N_8418,N_7682,N_7602);
and U8419 (N_8419,N_7819,N_7563);
and U8420 (N_8420,N_7797,N_7700);
nor U8421 (N_8421,N_7585,N_7778);
nand U8422 (N_8422,N_7819,N_7964);
nor U8423 (N_8423,N_7965,N_7702);
nand U8424 (N_8424,N_7803,N_7674);
xor U8425 (N_8425,N_7637,N_7721);
nor U8426 (N_8426,N_7834,N_7645);
nor U8427 (N_8427,N_7756,N_7779);
and U8428 (N_8428,N_7530,N_7602);
nand U8429 (N_8429,N_7776,N_7949);
or U8430 (N_8430,N_7856,N_7917);
and U8431 (N_8431,N_7626,N_7698);
or U8432 (N_8432,N_7532,N_7558);
or U8433 (N_8433,N_7613,N_7690);
or U8434 (N_8434,N_7501,N_7882);
nand U8435 (N_8435,N_7570,N_7991);
nor U8436 (N_8436,N_7668,N_7624);
or U8437 (N_8437,N_7632,N_7671);
or U8438 (N_8438,N_7779,N_7677);
nor U8439 (N_8439,N_7969,N_7565);
or U8440 (N_8440,N_7777,N_7650);
nor U8441 (N_8441,N_7762,N_7675);
and U8442 (N_8442,N_7597,N_7812);
and U8443 (N_8443,N_7891,N_7749);
nand U8444 (N_8444,N_7907,N_7571);
and U8445 (N_8445,N_7731,N_7611);
or U8446 (N_8446,N_7909,N_7815);
xor U8447 (N_8447,N_7733,N_7823);
nor U8448 (N_8448,N_7998,N_7961);
nand U8449 (N_8449,N_7826,N_7808);
nor U8450 (N_8450,N_7698,N_7942);
xnor U8451 (N_8451,N_7512,N_7867);
nand U8452 (N_8452,N_7997,N_7977);
or U8453 (N_8453,N_7567,N_7686);
and U8454 (N_8454,N_7954,N_7577);
and U8455 (N_8455,N_7712,N_7831);
and U8456 (N_8456,N_7932,N_7760);
and U8457 (N_8457,N_7609,N_7973);
and U8458 (N_8458,N_7638,N_7721);
and U8459 (N_8459,N_7919,N_7526);
nor U8460 (N_8460,N_7983,N_7562);
and U8461 (N_8461,N_7863,N_7915);
nor U8462 (N_8462,N_7717,N_7521);
and U8463 (N_8463,N_7741,N_7718);
xnor U8464 (N_8464,N_7759,N_7822);
nand U8465 (N_8465,N_7610,N_7890);
and U8466 (N_8466,N_7720,N_7799);
nor U8467 (N_8467,N_7613,N_7711);
nor U8468 (N_8468,N_7512,N_7658);
or U8469 (N_8469,N_7748,N_7997);
nor U8470 (N_8470,N_7900,N_7794);
nand U8471 (N_8471,N_7997,N_7585);
xor U8472 (N_8472,N_7835,N_7801);
or U8473 (N_8473,N_7828,N_7941);
and U8474 (N_8474,N_7589,N_7633);
nor U8475 (N_8475,N_7858,N_7800);
nor U8476 (N_8476,N_7661,N_7526);
or U8477 (N_8477,N_7562,N_7699);
and U8478 (N_8478,N_7908,N_7669);
and U8479 (N_8479,N_7856,N_7637);
or U8480 (N_8480,N_7891,N_7871);
or U8481 (N_8481,N_7871,N_7573);
or U8482 (N_8482,N_7995,N_7847);
xor U8483 (N_8483,N_7511,N_7984);
nor U8484 (N_8484,N_7524,N_7624);
nand U8485 (N_8485,N_7955,N_7937);
nand U8486 (N_8486,N_7538,N_7673);
nor U8487 (N_8487,N_7830,N_7821);
or U8488 (N_8488,N_7573,N_7775);
or U8489 (N_8489,N_7513,N_7591);
or U8490 (N_8490,N_7590,N_7581);
and U8491 (N_8491,N_7735,N_7535);
nand U8492 (N_8492,N_7598,N_7504);
nor U8493 (N_8493,N_7791,N_7509);
or U8494 (N_8494,N_7652,N_7534);
or U8495 (N_8495,N_7748,N_7536);
nor U8496 (N_8496,N_7738,N_7889);
xnor U8497 (N_8497,N_7730,N_7740);
nand U8498 (N_8498,N_7541,N_7638);
xnor U8499 (N_8499,N_7942,N_7579);
and U8500 (N_8500,N_8308,N_8413);
and U8501 (N_8501,N_8179,N_8039);
or U8502 (N_8502,N_8303,N_8176);
xor U8503 (N_8503,N_8460,N_8040);
nand U8504 (N_8504,N_8276,N_8360);
and U8505 (N_8505,N_8107,N_8328);
nand U8506 (N_8506,N_8305,N_8028);
nor U8507 (N_8507,N_8472,N_8223);
nand U8508 (N_8508,N_8285,N_8012);
or U8509 (N_8509,N_8169,N_8064);
and U8510 (N_8510,N_8387,N_8250);
nand U8511 (N_8511,N_8093,N_8479);
and U8512 (N_8512,N_8022,N_8206);
nor U8513 (N_8513,N_8031,N_8484);
or U8514 (N_8514,N_8408,N_8162);
and U8515 (N_8515,N_8459,N_8197);
nor U8516 (N_8516,N_8378,N_8120);
nand U8517 (N_8517,N_8189,N_8058);
nand U8518 (N_8518,N_8001,N_8420);
and U8519 (N_8519,N_8428,N_8006);
nand U8520 (N_8520,N_8211,N_8152);
nand U8521 (N_8521,N_8256,N_8457);
nor U8522 (N_8522,N_8345,N_8016);
and U8523 (N_8523,N_8042,N_8079);
nand U8524 (N_8524,N_8337,N_8365);
nor U8525 (N_8525,N_8299,N_8074);
xnor U8526 (N_8526,N_8000,N_8359);
nor U8527 (N_8527,N_8220,N_8161);
or U8528 (N_8528,N_8214,N_8199);
and U8529 (N_8529,N_8190,N_8008);
and U8530 (N_8530,N_8030,N_8136);
nand U8531 (N_8531,N_8224,N_8132);
and U8532 (N_8532,N_8036,N_8174);
or U8533 (N_8533,N_8246,N_8080);
or U8534 (N_8534,N_8316,N_8057);
nor U8535 (N_8535,N_8452,N_8394);
or U8536 (N_8536,N_8264,N_8053);
and U8537 (N_8537,N_8118,N_8478);
nor U8538 (N_8538,N_8468,N_8320);
nor U8539 (N_8539,N_8386,N_8421);
nand U8540 (N_8540,N_8082,N_8068);
nand U8541 (N_8541,N_8336,N_8150);
and U8542 (N_8542,N_8350,N_8486);
nand U8543 (N_8543,N_8329,N_8495);
nand U8544 (N_8544,N_8153,N_8186);
nand U8545 (N_8545,N_8444,N_8464);
or U8546 (N_8546,N_8181,N_8352);
nand U8547 (N_8547,N_8281,N_8018);
or U8548 (N_8548,N_8419,N_8052);
nor U8549 (N_8549,N_8251,N_8023);
and U8550 (N_8550,N_8406,N_8157);
and U8551 (N_8551,N_8314,N_8088);
or U8552 (N_8552,N_8343,N_8496);
and U8553 (N_8553,N_8092,N_8182);
nand U8554 (N_8554,N_8498,N_8194);
or U8555 (N_8555,N_8395,N_8284);
and U8556 (N_8556,N_8255,N_8433);
or U8557 (N_8557,N_8405,N_8196);
and U8558 (N_8558,N_8095,N_8497);
nor U8559 (N_8559,N_8142,N_8207);
and U8560 (N_8560,N_8400,N_8200);
or U8561 (N_8561,N_8091,N_8245);
nor U8562 (N_8562,N_8191,N_8210);
nor U8563 (N_8563,N_8312,N_8193);
nor U8564 (N_8564,N_8442,N_8051);
nand U8565 (N_8565,N_8077,N_8121);
nand U8566 (N_8566,N_8310,N_8253);
nand U8567 (N_8567,N_8274,N_8380);
and U8568 (N_8568,N_8086,N_8168);
and U8569 (N_8569,N_8443,N_8104);
nand U8570 (N_8570,N_8390,N_8029);
nor U8571 (N_8571,N_8358,N_8249);
nand U8572 (N_8572,N_8205,N_8171);
nand U8573 (N_8573,N_8105,N_8278);
and U8574 (N_8574,N_8158,N_8002);
nor U8575 (N_8575,N_8146,N_8026);
or U8576 (N_8576,N_8247,N_8041);
nor U8577 (N_8577,N_8494,N_8014);
or U8578 (N_8578,N_8015,N_8208);
xor U8579 (N_8579,N_8163,N_8412);
or U8580 (N_8580,N_8111,N_8403);
nor U8581 (N_8581,N_8155,N_8259);
and U8582 (N_8582,N_8135,N_8137);
and U8583 (N_8583,N_8364,N_8034);
and U8584 (N_8584,N_8499,N_8315);
nand U8585 (N_8585,N_8177,N_8376);
and U8586 (N_8586,N_8455,N_8180);
or U8587 (N_8587,N_8017,N_8450);
or U8588 (N_8588,N_8235,N_8431);
nor U8589 (N_8589,N_8423,N_8090);
and U8590 (N_8590,N_8293,N_8125);
nor U8591 (N_8591,N_8324,N_8382);
xor U8592 (N_8592,N_8124,N_8279);
and U8593 (N_8593,N_8123,N_8144);
nand U8594 (N_8594,N_8258,N_8254);
and U8595 (N_8595,N_8415,N_8465);
and U8596 (N_8596,N_8165,N_8290);
nor U8597 (N_8597,N_8325,N_8113);
and U8598 (N_8598,N_8055,N_8096);
nand U8599 (N_8599,N_8449,N_8466);
and U8600 (N_8600,N_8139,N_8148);
nor U8601 (N_8601,N_8188,N_8453);
and U8602 (N_8602,N_8263,N_8213);
nor U8603 (N_8603,N_8348,N_8222);
nand U8604 (N_8604,N_8084,N_8291);
nand U8605 (N_8605,N_8354,N_8417);
nand U8606 (N_8606,N_8447,N_8047);
and U8607 (N_8607,N_8356,N_8363);
or U8608 (N_8608,N_8236,N_8393);
nand U8609 (N_8609,N_8005,N_8073);
nand U8610 (N_8610,N_8221,N_8045);
or U8611 (N_8611,N_8108,N_8302);
nor U8612 (N_8612,N_8319,N_8192);
and U8613 (N_8613,N_8019,N_8141);
nand U8614 (N_8614,N_8432,N_8094);
and U8615 (N_8615,N_8438,N_8409);
or U8616 (N_8616,N_8078,N_8402);
nor U8617 (N_8617,N_8437,N_8272);
nor U8618 (N_8618,N_8270,N_8178);
or U8619 (N_8619,N_8020,N_8355);
nor U8620 (N_8620,N_8441,N_8140);
nand U8621 (N_8621,N_8410,N_8375);
nand U8622 (N_8622,N_8071,N_8366);
or U8623 (N_8623,N_8240,N_8267);
nand U8624 (N_8624,N_8166,N_8377);
nor U8625 (N_8625,N_8327,N_8338);
or U8626 (N_8626,N_8225,N_8492);
or U8627 (N_8627,N_8145,N_8297);
nand U8628 (N_8628,N_8318,N_8330);
nand U8629 (N_8629,N_8167,N_8089);
or U8630 (N_8630,N_8404,N_8143);
and U8631 (N_8631,N_8147,N_8228);
and U8632 (N_8632,N_8226,N_8069);
nor U8633 (N_8633,N_8454,N_8361);
and U8634 (N_8634,N_8009,N_8011);
nand U8635 (N_8635,N_8097,N_8487);
or U8636 (N_8636,N_8271,N_8280);
and U8637 (N_8637,N_8480,N_8231);
nor U8638 (N_8638,N_8244,N_8151);
nand U8639 (N_8639,N_8066,N_8087);
or U8640 (N_8640,N_8204,N_8217);
nor U8641 (N_8641,N_8202,N_8372);
nor U8642 (N_8642,N_8288,N_8296);
and U8643 (N_8643,N_8416,N_8184);
or U8644 (N_8644,N_8368,N_8289);
or U8645 (N_8645,N_8203,N_8128);
nor U8646 (N_8646,N_8007,N_8075);
nor U8647 (N_8647,N_8379,N_8490);
or U8648 (N_8648,N_8122,N_8227);
or U8649 (N_8649,N_8114,N_8043);
nand U8650 (N_8650,N_8083,N_8391);
nor U8651 (N_8651,N_8138,N_8451);
and U8652 (N_8652,N_8357,N_8229);
nand U8653 (N_8653,N_8397,N_8277);
nor U8654 (N_8654,N_8238,N_8102);
or U8655 (N_8655,N_8369,N_8130);
nor U8656 (N_8656,N_8474,N_8230);
nand U8657 (N_8657,N_8212,N_8109);
nand U8658 (N_8658,N_8414,N_8117);
nor U8659 (N_8659,N_8347,N_8126);
nand U8660 (N_8660,N_8334,N_8021);
nand U8661 (N_8661,N_8475,N_8424);
and U8662 (N_8662,N_8301,N_8209);
nor U8663 (N_8663,N_8300,N_8063);
or U8664 (N_8664,N_8313,N_8339);
nor U8665 (N_8665,N_8046,N_8426);
nor U8666 (N_8666,N_8381,N_8187);
nor U8667 (N_8667,N_8072,N_8027);
or U8668 (N_8668,N_8103,N_8219);
or U8669 (N_8669,N_8004,N_8099);
or U8670 (N_8670,N_8399,N_8216);
and U8671 (N_8671,N_8389,N_8116);
or U8672 (N_8672,N_8434,N_8172);
and U8673 (N_8673,N_8341,N_8242);
xor U8674 (N_8674,N_8445,N_8134);
and U8675 (N_8675,N_8392,N_8489);
nor U8676 (N_8676,N_8233,N_8456);
nand U8677 (N_8677,N_8458,N_8234);
or U8678 (N_8678,N_8243,N_8110);
or U8679 (N_8679,N_8033,N_8218);
and U8680 (N_8680,N_8062,N_8059);
nor U8681 (N_8681,N_8311,N_8050);
or U8682 (N_8682,N_8085,N_8037);
nand U8683 (N_8683,N_8127,N_8248);
or U8684 (N_8684,N_8129,N_8101);
and U8685 (N_8685,N_8237,N_8385);
nor U8686 (N_8686,N_8032,N_8353);
nor U8687 (N_8687,N_8396,N_8439);
nand U8688 (N_8688,N_8383,N_8374);
and U8689 (N_8689,N_8373,N_8232);
or U8690 (N_8690,N_8106,N_8435);
nand U8691 (N_8691,N_8422,N_8349);
or U8692 (N_8692,N_8401,N_8481);
and U8693 (N_8693,N_8119,N_8309);
or U8694 (N_8694,N_8056,N_8160);
nand U8695 (N_8695,N_8010,N_8418);
nand U8696 (N_8696,N_8266,N_8195);
and U8697 (N_8697,N_8470,N_8265);
or U8698 (N_8698,N_8239,N_8269);
or U8699 (N_8699,N_8287,N_8185);
or U8700 (N_8700,N_8462,N_8013);
nor U8701 (N_8701,N_8425,N_8159);
or U8702 (N_8702,N_8154,N_8164);
xnor U8703 (N_8703,N_8215,N_8038);
or U8704 (N_8704,N_8483,N_8260);
and U8705 (N_8705,N_8183,N_8070);
and U8706 (N_8706,N_8471,N_8307);
nand U8707 (N_8707,N_8362,N_8411);
and U8708 (N_8708,N_8286,N_8252);
and U8709 (N_8709,N_8304,N_8398);
or U8710 (N_8710,N_8275,N_8346);
or U8711 (N_8711,N_8323,N_8384);
nor U8712 (N_8712,N_8351,N_8131);
or U8713 (N_8713,N_8461,N_8340);
nor U8714 (N_8714,N_8388,N_8333);
nor U8715 (N_8715,N_8035,N_8049);
and U8716 (N_8716,N_8261,N_8257);
nand U8717 (N_8717,N_8332,N_8156);
or U8718 (N_8718,N_8448,N_8048);
nand U8719 (N_8719,N_8317,N_8344);
and U8720 (N_8720,N_8133,N_8370);
nor U8721 (N_8721,N_8467,N_8322);
or U8722 (N_8722,N_8491,N_8469);
nor U8723 (N_8723,N_8273,N_8061);
and U8724 (N_8724,N_8482,N_8065);
and U8725 (N_8725,N_8098,N_8493);
and U8726 (N_8726,N_8367,N_8024);
nor U8727 (N_8727,N_8149,N_8060);
and U8728 (N_8728,N_8407,N_8335);
nand U8729 (N_8729,N_8298,N_8331);
nor U8730 (N_8730,N_8429,N_8463);
nor U8731 (N_8731,N_8115,N_8430);
nand U8732 (N_8732,N_8100,N_8025);
or U8733 (N_8733,N_8295,N_8067);
or U8734 (N_8734,N_8342,N_8446);
xor U8735 (N_8735,N_8282,N_8440);
or U8736 (N_8736,N_8198,N_8076);
or U8737 (N_8737,N_8473,N_8427);
xnor U8738 (N_8738,N_8175,N_8262);
and U8739 (N_8739,N_8294,N_8112);
or U8740 (N_8740,N_8477,N_8283);
or U8741 (N_8741,N_8321,N_8054);
or U8742 (N_8742,N_8292,N_8436);
nor U8743 (N_8743,N_8081,N_8003);
nand U8744 (N_8744,N_8371,N_8268);
or U8745 (N_8745,N_8306,N_8170);
nor U8746 (N_8746,N_8476,N_8044);
nand U8747 (N_8747,N_8326,N_8173);
or U8748 (N_8748,N_8201,N_8488);
nand U8749 (N_8749,N_8485,N_8241);
or U8750 (N_8750,N_8210,N_8498);
or U8751 (N_8751,N_8211,N_8179);
nor U8752 (N_8752,N_8198,N_8149);
or U8753 (N_8753,N_8097,N_8348);
or U8754 (N_8754,N_8112,N_8040);
and U8755 (N_8755,N_8125,N_8243);
nand U8756 (N_8756,N_8177,N_8422);
nand U8757 (N_8757,N_8359,N_8067);
nor U8758 (N_8758,N_8241,N_8356);
or U8759 (N_8759,N_8360,N_8155);
xnor U8760 (N_8760,N_8370,N_8410);
or U8761 (N_8761,N_8072,N_8498);
nand U8762 (N_8762,N_8220,N_8244);
nand U8763 (N_8763,N_8087,N_8215);
xor U8764 (N_8764,N_8428,N_8425);
or U8765 (N_8765,N_8279,N_8369);
or U8766 (N_8766,N_8314,N_8344);
or U8767 (N_8767,N_8075,N_8363);
and U8768 (N_8768,N_8168,N_8244);
nor U8769 (N_8769,N_8142,N_8182);
nor U8770 (N_8770,N_8039,N_8285);
nand U8771 (N_8771,N_8406,N_8160);
or U8772 (N_8772,N_8300,N_8126);
nand U8773 (N_8773,N_8380,N_8212);
nand U8774 (N_8774,N_8406,N_8479);
nand U8775 (N_8775,N_8010,N_8003);
or U8776 (N_8776,N_8262,N_8156);
nand U8777 (N_8777,N_8256,N_8369);
nand U8778 (N_8778,N_8487,N_8304);
nand U8779 (N_8779,N_8103,N_8182);
nor U8780 (N_8780,N_8368,N_8487);
and U8781 (N_8781,N_8208,N_8467);
or U8782 (N_8782,N_8133,N_8019);
or U8783 (N_8783,N_8079,N_8405);
and U8784 (N_8784,N_8224,N_8410);
and U8785 (N_8785,N_8197,N_8030);
nand U8786 (N_8786,N_8277,N_8338);
nor U8787 (N_8787,N_8215,N_8440);
or U8788 (N_8788,N_8237,N_8413);
and U8789 (N_8789,N_8438,N_8441);
and U8790 (N_8790,N_8220,N_8424);
nor U8791 (N_8791,N_8288,N_8294);
and U8792 (N_8792,N_8425,N_8411);
or U8793 (N_8793,N_8128,N_8376);
and U8794 (N_8794,N_8013,N_8235);
nand U8795 (N_8795,N_8392,N_8416);
and U8796 (N_8796,N_8169,N_8233);
nand U8797 (N_8797,N_8306,N_8310);
or U8798 (N_8798,N_8233,N_8277);
and U8799 (N_8799,N_8142,N_8300);
nor U8800 (N_8800,N_8098,N_8038);
nand U8801 (N_8801,N_8176,N_8098);
nor U8802 (N_8802,N_8055,N_8443);
xor U8803 (N_8803,N_8450,N_8132);
or U8804 (N_8804,N_8147,N_8161);
or U8805 (N_8805,N_8268,N_8427);
nand U8806 (N_8806,N_8059,N_8076);
nor U8807 (N_8807,N_8125,N_8300);
nand U8808 (N_8808,N_8247,N_8052);
or U8809 (N_8809,N_8311,N_8006);
nor U8810 (N_8810,N_8067,N_8036);
nand U8811 (N_8811,N_8110,N_8223);
or U8812 (N_8812,N_8169,N_8159);
or U8813 (N_8813,N_8189,N_8324);
nor U8814 (N_8814,N_8086,N_8496);
nor U8815 (N_8815,N_8499,N_8269);
and U8816 (N_8816,N_8377,N_8357);
or U8817 (N_8817,N_8356,N_8112);
nand U8818 (N_8818,N_8405,N_8037);
nand U8819 (N_8819,N_8139,N_8401);
or U8820 (N_8820,N_8287,N_8247);
and U8821 (N_8821,N_8009,N_8182);
and U8822 (N_8822,N_8061,N_8328);
nor U8823 (N_8823,N_8262,N_8065);
or U8824 (N_8824,N_8420,N_8307);
or U8825 (N_8825,N_8359,N_8291);
or U8826 (N_8826,N_8407,N_8329);
and U8827 (N_8827,N_8388,N_8487);
nor U8828 (N_8828,N_8339,N_8082);
nor U8829 (N_8829,N_8219,N_8323);
and U8830 (N_8830,N_8188,N_8243);
nand U8831 (N_8831,N_8491,N_8338);
nor U8832 (N_8832,N_8040,N_8029);
and U8833 (N_8833,N_8140,N_8457);
and U8834 (N_8834,N_8343,N_8371);
and U8835 (N_8835,N_8317,N_8066);
or U8836 (N_8836,N_8479,N_8083);
nand U8837 (N_8837,N_8073,N_8449);
or U8838 (N_8838,N_8007,N_8235);
or U8839 (N_8839,N_8276,N_8016);
and U8840 (N_8840,N_8473,N_8080);
nor U8841 (N_8841,N_8034,N_8104);
or U8842 (N_8842,N_8442,N_8103);
and U8843 (N_8843,N_8069,N_8098);
nor U8844 (N_8844,N_8076,N_8278);
nor U8845 (N_8845,N_8254,N_8490);
or U8846 (N_8846,N_8105,N_8233);
nand U8847 (N_8847,N_8487,N_8400);
and U8848 (N_8848,N_8140,N_8232);
or U8849 (N_8849,N_8342,N_8188);
nand U8850 (N_8850,N_8226,N_8379);
and U8851 (N_8851,N_8265,N_8438);
and U8852 (N_8852,N_8204,N_8154);
and U8853 (N_8853,N_8372,N_8464);
or U8854 (N_8854,N_8055,N_8031);
nand U8855 (N_8855,N_8137,N_8184);
or U8856 (N_8856,N_8331,N_8176);
or U8857 (N_8857,N_8001,N_8400);
and U8858 (N_8858,N_8387,N_8455);
nand U8859 (N_8859,N_8450,N_8193);
nand U8860 (N_8860,N_8353,N_8388);
nor U8861 (N_8861,N_8404,N_8047);
nor U8862 (N_8862,N_8030,N_8252);
nand U8863 (N_8863,N_8337,N_8425);
or U8864 (N_8864,N_8266,N_8477);
nand U8865 (N_8865,N_8201,N_8108);
nor U8866 (N_8866,N_8091,N_8039);
and U8867 (N_8867,N_8290,N_8138);
or U8868 (N_8868,N_8268,N_8031);
nand U8869 (N_8869,N_8134,N_8008);
nor U8870 (N_8870,N_8226,N_8203);
nand U8871 (N_8871,N_8043,N_8409);
or U8872 (N_8872,N_8066,N_8465);
and U8873 (N_8873,N_8073,N_8175);
and U8874 (N_8874,N_8105,N_8100);
or U8875 (N_8875,N_8004,N_8342);
nand U8876 (N_8876,N_8280,N_8028);
nand U8877 (N_8877,N_8431,N_8352);
nand U8878 (N_8878,N_8014,N_8348);
and U8879 (N_8879,N_8343,N_8083);
nor U8880 (N_8880,N_8103,N_8268);
and U8881 (N_8881,N_8303,N_8155);
nor U8882 (N_8882,N_8454,N_8084);
xnor U8883 (N_8883,N_8190,N_8199);
or U8884 (N_8884,N_8347,N_8249);
nor U8885 (N_8885,N_8046,N_8451);
nand U8886 (N_8886,N_8383,N_8019);
or U8887 (N_8887,N_8244,N_8481);
nand U8888 (N_8888,N_8293,N_8214);
and U8889 (N_8889,N_8472,N_8304);
and U8890 (N_8890,N_8497,N_8025);
nand U8891 (N_8891,N_8499,N_8290);
and U8892 (N_8892,N_8308,N_8454);
and U8893 (N_8893,N_8390,N_8277);
nor U8894 (N_8894,N_8426,N_8099);
or U8895 (N_8895,N_8452,N_8148);
nor U8896 (N_8896,N_8441,N_8113);
nand U8897 (N_8897,N_8043,N_8196);
or U8898 (N_8898,N_8098,N_8280);
nand U8899 (N_8899,N_8055,N_8272);
nand U8900 (N_8900,N_8285,N_8214);
nand U8901 (N_8901,N_8240,N_8473);
and U8902 (N_8902,N_8398,N_8481);
and U8903 (N_8903,N_8292,N_8406);
or U8904 (N_8904,N_8190,N_8064);
and U8905 (N_8905,N_8203,N_8249);
or U8906 (N_8906,N_8052,N_8264);
or U8907 (N_8907,N_8188,N_8352);
nor U8908 (N_8908,N_8183,N_8205);
and U8909 (N_8909,N_8151,N_8270);
nand U8910 (N_8910,N_8281,N_8349);
and U8911 (N_8911,N_8208,N_8420);
nor U8912 (N_8912,N_8453,N_8486);
nor U8913 (N_8913,N_8317,N_8254);
and U8914 (N_8914,N_8000,N_8002);
and U8915 (N_8915,N_8273,N_8039);
nand U8916 (N_8916,N_8085,N_8386);
and U8917 (N_8917,N_8318,N_8091);
or U8918 (N_8918,N_8478,N_8281);
or U8919 (N_8919,N_8013,N_8077);
nor U8920 (N_8920,N_8338,N_8115);
nor U8921 (N_8921,N_8070,N_8061);
and U8922 (N_8922,N_8125,N_8433);
nand U8923 (N_8923,N_8479,N_8122);
and U8924 (N_8924,N_8282,N_8418);
and U8925 (N_8925,N_8236,N_8295);
nand U8926 (N_8926,N_8295,N_8245);
nand U8927 (N_8927,N_8039,N_8469);
nand U8928 (N_8928,N_8207,N_8385);
nand U8929 (N_8929,N_8447,N_8289);
nand U8930 (N_8930,N_8480,N_8040);
nor U8931 (N_8931,N_8424,N_8017);
and U8932 (N_8932,N_8165,N_8486);
or U8933 (N_8933,N_8008,N_8340);
and U8934 (N_8934,N_8354,N_8101);
nor U8935 (N_8935,N_8398,N_8416);
or U8936 (N_8936,N_8335,N_8124);
nand U8937 (N_8937,N_8196,N_8218);
and U8938 (N_8938,N_8097,N_8061);
nand U8939 (N_8939,N_8212,N_8325);
and U8940 (N_8940,N_8259,N_8369);
nor U8941 (N_8941,N_8165,N_8274);
or U8942 (N_8942,N_8078,N_8375);
nor U8943 (N_8943,N_8303,N_8025);
or U8944 (N_8944,N_8118,N_8364);
and U8945 (N_8945,N_8137,N_8297);
and U8946 (N_8946,N_8204,N_8284);
nand U8947 (N_8947,N_8458,N_8178);
nor U8948 (N_8948,N_8261,N_8451);
and U8949 (N_8949,N_8366,N_8057);
or U8950 (N_8950,N_8154,N_8158);
or U8951 (N_8951,N_8165,N_8394);
and U8952 (N_8952,N_8187,N_8349);
and U8953 (N_8953,N_8443,N_8053);
nor U8954 (N_8954,N_8284,N_8126);
or U8955 (N_8955,N_8103,N_8165);
and U8956 (N_8956,N_8490,N_8451);
nor U8957 (N_8957,N_8243,N_8322);
xnor U8958 (N_8958,N_8267,N_8206);
or U8959 (N_8959,N_8134,N_8224);
or U8960 (N_8960,N_8181,N_8472);
nor U8961 (N_8961,N_8379,N_8311);
nor U8962 (N_8962,N_8066,N_8494);
or U8963 (N_8963,N_8396,N_8095);
and U8964 (N_8964,N_8220,N_8241);
nand U8965 (N_8965,N_8022,N_8381);
nand U8966 (N_8966,N_8292,N_8391);
nand U8967 (N_8967,N_8079,N_8040);
nor U8968 (N_8968,N_8284,N_8117);
nand U8969 (N_8969,N_8299,N_8447);
and U8970 (N_8970,N_8150,N_8416);
nand U8971 (N_8971,N_8218,N_8328);
nand U8972 (N_8972,N_8135,N_8045);
nand U8973 (N_8973,N_8019,N_8474);
nand U8974 (N_8974,N_8139,N_8355);
nand U8975 (N_8975,N_8419,N_8475);
and U8976 (N_8976,N_8184,N_8124);
and U8977 (N_8977,N_8329,N_8125);
nand U8978 (N_8978,N_8276,N_8248);
nand U8979 (N_8979,N_8485,N_8363);
and U8980 (N_8980,N_8164,N_8354);
and U8981 (N_8981,N_8405,N_8153);
nor U8982 (N_8982,N_8155,N_8254);
nor U8983 (N_8983,N_8480,N_8392);
nor U8984 (N_8984,N_8180,N_8458);
or U8985 (N_8985,N_8219,N_8305);
or U8986 (N_8986,N_8044,N_8073);
nor U8987 (N_8987,N_8356,N_8088);
nor U8988 (N_8988,N_8038,N_8334);
nor U8989 (N_8989,N_8254,N_8311);
nand U8990 (N_8990,N_8054,N_8389);
xnor U8991 (N_8991,N_8120,N_8088);
and U8992 (N_8992,N_8156,N_8031);
nor U8993 (N_8993,N_8270,N_8049);
nand U8994 (N_8994,N_8302,N_8018);
nand U8995 (N_8995,N_8154,N_8237);
and U8996 (N_8996,N_8431,N_8010);
and U8997 (N_8997,N_8280,N_8174);
nor U8998 (N_8998,N_8199,N_8176);
and U8999 (N_8999,N_8478,N_8226);
nand U9000 (N_9000,N_8698,N_8544);
or U9001 (N_9001,N_8896,N_8739);
or U9002 (N_9002,N_8561,N_8586);
nand U9003 (N_9003,N_8861,N_8898);
or U9004 (N_9004,N_8514,N_8902);
or U9005 (N_9005,N_8917,N_8505);
or U9006 (N_9006,N_8768,N_8655);
or U9007 (N_9007,N_8809,N_8527);
and U9008 (N_9008,N_8961,N_8747);
or U9009 (N_9009,N_8609,N_8873);
or U9010 (N_9010,N_8963,N_8745);
or U9011 (N_9011,N_8740,N_8910);
nand U9012 (N_9012,N_8560,N_8770);
and U9013 (N_9013,N_8969,N_8901);
and U9014 (N_9014,N_8869,N_8676);
or U9015 (N_9015,N_8881,N_8858);
nor U9016 (N_9016,N_8663,N_8801);
or U9017 (N_9017,N_8987,N_8593);
nor U9018 (N_9018,N_8570,N_8746);
or U9019 (N_9019,N_8839,N_8882);
nand U9020 (N_9020,N_8808,N_8693);
nand U9021 (N_9021,N_8893,N_8639);
and U9022 (N_9022,N_8712,N_8729);
nand U9023 (N_9023,N_8500,N_8918);
and U9024 (N_9024,N_8925,N_8989);
and U9025 (N_9025,N_8798,N_8767);
nor U9026 (N_9026,N_8684,N_8603);
or U9027 (N_9027,N_8580,N_8583);
nor U9028 (N_9028,N_8588,N_8935);
nand U9029 (N_9029,N_8678,N_8512);
nand U9030 (N_9030,N_8926,N_8995);
or U9031 (N_9031,N_8730,N_8535);
or U9032 (N_9032,N_8824,N_8792);
xor U9033 (N_9033,N_8857,N_8681);
or U9034 (N_9034,N_8673,N_8735);
or U9035 (N_9035,N_8933,N_8652);
nand U9036 (N_9036,N_8548,N_8744);
nor U9037 (N_9037,N_8725,N_8601);
nand U9038 (N_9038,N_8709,N_8870);
or U9039 (N_9039,N_8836,N_8728);
nor U9040 (N_9040,N_8856,N_8934);
nand U9041 (N_9041,N_8518,N_8618);
nand U9042 (N_9042,N_8617,N_8972);
nand U9043 (N_9043,N_8790,N_8846);
nand U9044 (N_9044,N_8531,N_8721);
nor U9045 (N_9045,N_8762,N_8960);
nor U9046 (N_9046,N_8868,N_8677);
or U9047 (N_9047,N_8822,N_8785);
or U9048 (N_9048,N_8853,N_8540);
nor U9049 (N_9049,N_8837,N_8890);
nor U9050 (N_9050,N_8754,N_8708);
or U9051 (N_9051,N_8920,N_8722);
nor U9052 (N_9052,N_8965,N_8766);
nand U9053 (N_9053,N_8862,N_8841);
xnor U9054 (N_9054,N_8664,N_8880);
or U9055 (N_9055,N_8973,N_8884);
nor U9056 (N_9056,N_8971,N_8760);
xnor U9057 (N_9057,N_8621,N_8634);
nor U9058 (N_9058,N_8707,N_8932);
nor U9059 (N_9059,N_8993,N_8945);
xnor U9060 (N_9060,N_8679,N_8631);
nor U9061 (N_9061,N_8930,N_8510);
and U9062 (N_9062,N_8562,N_8877);
nand U9063 (N_9063,N_8906,N_8619);
nand U9064 (N_9064,N_8661,N_8615);
nor U9065 (N_9065,N_8814,N_8635);
and U9066 (N_9066,N_8797,N_8694);
or U9067 (N_9067,N_8670,N_8688);
nor U9068 (N_9068,N_8795,N_8914);
nand U9069 (N_9069,N_8913,N_8602);
and U9070 (N_9070,N_8690,N_8563);
and U9071 (N_9071,N_8878,N_8522);
and U9072 (N_9072,N_8689,N_8867);
or U9073 (N_9073,N_8794,N_8992);
nand U9074 (N_9074,N_8549,N_8813);
nor U9075 (N_9075,N_8607,N_8843);
and U9076 (N_9076,N_8959,N_8592);
nand U9077 (N_9077,N_8953,N_8929);
or U9078 (N_9078,N_8581,N_8695);
or U9079 (N_9079,N_8682,N_8741);
nand U9080 (N_9080,N_8612,N_8598);
nand U9081 (N_9081,N_8590,N_8939);
nor U9082 (N_9082,N_8521,N_8657);
or U9083 (N_9083,N_8800,N_8916);
or U9084 (N_9084,N_8951,N_8622);
nor U9085 (N_9085,N_8530,N_8895);
nor U9086 (N_9086,N_8555,N_8523);
and U9087 (N_9087,N_8984,N_8541);
or U9088 (N_9088,N_8687,N_8921);
nor U9089 (N_9089,N_8724,N_8700);
nand U9090 (N_9090,N_8537,N_8937);
xor U9091 (N_9091,N_8966,N_8900);
or U9092 (N_9092,N_8641,N_8647);
or U9093 (N_9093,N_8737,N_8553);
nand U9094 (N_9094,N_8756,N_8557);
nand U9095 (N_9095,N_8646,N_8958);
or U9096 (N_9096,N_8576,N_8669);
or U9097 (N_9097,N_8788,N_8885);
nand U9098 (N_9098,N_8650,N_8651);
and U9099 (N_9099,N_8938,N_8772);
nand U9100 (N_9100,N_8823,N_8803);
nor U9101 (N_9101,N_8763,N_8587);
xnor U9102 (N_9102,N_8831,N_8940);
nand U9103 (N_9103,N_8571,N_8931);
nor U9104 (N_9104,N_8946,N_8671);
nand U9105 (N_9105,N_8637,N_8743);
nand U9106 (N_9106,N_8962,N_8977);
nand U9107 (N_9107,N_8828,N_8714);
nand U9108 (N_9108,N_8524,N_8628);
and U9109 (N_9109,N_8680,N_8723);
nand U9110 (N_9110,N_8738,N_8594);
nor U9111 (N_9111,N_8978,N_8720);
nor U9112 (N_9112,N_8791,N_8875);
and U9113 (N_9113,N_8928,N_8665);
nor U9114 (N_9114,N_8572,N_8950);
nor U9115 (N_9115,N_8852,N_8964);
and U9116 (N_9116,N_8784,N_8787);
nand U9117 (N_9117,N_8666,N_8886);
nor U9118 (N_9118,N_8879,N_8550);
nand U9119 (N_9119,N_8954,N_8513);
and U9120 (N_9120,N_8833,N_8713);
nand U9121 (N_9121,N_8585,N_8919);
nor U9122 (N_9122,N_8829,N_8630);
nor U9123 (N_9123,N_8614,N_8911);
and U9124 (N_9124,N_8776,N_8656);
nand U9125 (N_9125,N_8811,N_8591);
nand U9126 (N_9126,N_8922,N_8764);
or U9127 (N_9127,N_8696,N_8956);
and U9128 (N_9128,N_8558,N_8582);
or U9129 (N_9129,N_8819,N_8998);
and U9130 (N_9130,N_8575,N_8623);
nand U9131 (N_9131,N_8704,N_8699);
and U9132 (N_9132,N_8542,N_8817);
and U9133 (N_9133,N_8826,N_8711);
and U9134 (N_9134,N_8830,N_8848);
or U9135 (N_9135,N_8545,N_8662);
and U9136 (N_9136,N_8789,N_8955);
or U9137 (N_9137,N_8847,N_8683);
or U9138 (N_9138,N_8777,N_8812);
and U9139 (N_9139,N_8584,N_8927);
or U9140 (N_9140,N_8624,N_8838);
nor U9141 (N_9141,N_8627,N_8595);
and U9142 (N_9142,N_8717,N_8810);
nand U9143 (N_9143,N_8604,N_8804);
nor U9144 (N_9144,N_8509,N_8520);
nor U9145 (N_9145,N_8632,N_8556);
nor U9146 (N_9146,N_8779,N_8643);
or U9147 (N_9147,N_8716,N_8508);
nor U9148 (N_9148,N_8765,N_8775);
and U9149 (N_9149,N_8908,N_8807);
nor U9150 (N_9150,N_8999,N_8654);
or U9151 (N_9151,N_8517,N_8719);
and U9152 (N_9152,N_8751,N_8674);
or U9153 (N_9153,N_8596,N_8749);
nand U9154 (N_9154,N_8757,N_8949);
nor U9155 (N_9155,N_8990,N_8552);
nor U9156 (N_9156,N_8872,N_8706);
nand U9157 (N_9157,N_8793,N_8667);
and U9158 (N_9158,N_8608,N_8904);
or U9159 (N_9159,N_8988,N_8525);
and U9160 (N_9160,N_8539,N_8705);
and U9161 (N_9161,N_8806,N_8564);
or U9162 (N_9162,N_8726,N_8529);
nand U9163 (N_9163,N_8864,N_8502);
nand U9164 (N_9164,N_8907,N_8891);
or U9165 (N_9165,N_8805,N_8566);
and U9166 (N_9166,N_8511,N_8915);
or U9167 (N_9167,N_8503,N_8942);
nand U9168 (N_9168,N_8968,N_8547);
and U9169 (N_9169,N_8675,N_8578);
or U9170 (N_9170,N_8519,N_8597);
or U9171 (N_9171,N_8799,N_8515);
or U9172 (N_9172,N_8967,N_8644);
and U9173 (N_9173,N_8702,N_8626);
nand U9174 (N_9174,N_8753,N_8686);
and U9175 (N_9175,N_8820,N_8859);
and U9176 (N_9176,N_8783,N_8504);
and U9177 (N_9177,N_8874,N_8685);
nor U9178 (N_9178,N_8997,N_8835);
or U9179 (N_9179,N_8983,N_8701);
and U9180 (N_9180,N_8638,N_8815);
nand U9181 (N_9181,N_8780,N_8672);
nand U9182 (N_9182,N_8616,N_8970);
nand U9183 (N_9183,N_8589,N_8710);
nor U9184 (N_9184,N_8844,N_8736);
or U9185 (N_9185,N_8986,N_8568);
and U9186 (N_9186,N_8516,N_8936);
or U9187 (N_9187,N_8850,N_8645);
nor U9188 (N_9188,N_8871,N_8849);
nor U9189 (N_9189,N_8912,N_8827);
or U9190 (N_9190,N_8979,N_8957);
nor U9191 (N_9191,N_8565,N_8909);
nor U9192 (N_9192,N_8577,N_8818);
nor U9193 (N_9193,N_8976,N_8506);
and U9194 (N_9194,N_8752,N_8642);
or U9195 (N_9195,N_8854,N_8742);
nor U9196 (N_9196,N_8620,N_8629);
nor U9197 (N_9197,N_8842,N_8821);
nor U9198 (N_9198,N_8755,N_8733);
or U9199 (N_9199,N_8985,N_8692);
nor U9200 (N_9200,N_8802,N_8761);
nor U9201 (N_9201,N_8625,N_8579);
or U9202 (N_9202,N_8649,N_8982);
nand U9203 (N_9203,N_8528,N_8551);
nor U9204 (N_9204,N_8691,N_8860);
or U9205 (N_9205,N_8610,N_8981);
nand U9206 (N_9206,N_8507,N_8948);
and U9207 (N_9207,N_8892,N_8748);
nand U9208 (N_9208,N_8660,N_8974);
and U9209 (N_9209,N_8855,N_8703);
and U9210 (N_9210,N_8781,N_8786);
nor U9211 (N_9211,N_8559,N_8774);
nand U9212 (N_9212,N_8865,N_8866);
and U9213 (N_9213,N_8501,N_8876);
or U9214 (N_9214,N_8567,N_8889);
or U9215 (N_9215,N_8943,N_8554);
nor U9216 (N_9216,N_8863,N_8605);
and U9217 (N_9217,N_8536,N_8923);
or U9218 (N_9218,N_8758,N_8894);
and U9219 (N_9219,N_8825,N_8546);
or U9220 (N_9220,N_8599,N_8883);
or U9221 (N_9221,N_8727,N_8648);
or U9222 (N_9222,N_8796,N_8574);
nand U9223 (N_9223,N_8640,N_8947);
or U9224 (N_9224,N_8734,N_8653);
or U9225 (N_9225,N_8569,N_8975);
or U9226 (N_9226,N_8613,N_8899);
nand U9227 (N_9227,N_8538,N_8759);
nand U9228 (N_9228,N_8715,N_8534);
nor U9229 (N_9229,N_8816,N_8573);
and U9230 (N_9230,N_8903,N_8532);
and U9231 (N_9231,N_8851,N_8773);
nand U9232 (N_9232,N_8941,N_8887);
or U9233 (N_9233,N_8952,N_8533);
nor U9234 (N_9234,N_8905,N_8845);
xnor U9235 (N_9235,N_8731,N_8778);
or U9236 (N_9236,N_8718,N_8888);
nand U9237 (N_9237,N_8633,N_8980);
nor U9238 (N_9238,N_8658,N_8769);
xnor U9239 (N_9239,N_8600,N_8606);
nand U9240 (N_9240,N_8732,N_8668);
nor U9241 (N_9241,N_8832,N_8897);
nor U9242 (N_9242,N_8611,N_8924);
and U9243 (N_9243,N_8636,N_8659);
and U9244 (N_9244,N_8771,N_8543);
and U9245 (N_9245,N_8996,N_8697);
nand U9246 (N_9246,N_8526,N_8994);
and U9247 (N_9247,N_8782,N_8991);
nand U9248 (N_9248,N_8834,N_8840);
or U9249 (N_9249,N_8944,N_8750);
nand U9250 (N_9250,N_8865,N_8975);
nor U9251 (N_9251,N_8995,N_8572);
and U9252 (N_9252,N_8776,N_8531);
nand U9253 (N_9253,N_8655,N_8508);
nor U9254 (N_9254,N_8710,N_8911);
or U9255 (N_9255,N_8889,N_8790);
nand U9256 (N_9256,N_8987,N_8612);
nor U9257 (N_9257,N_8687,N_8901);
or U9258 (N_9258,N_8948,N_8668);
nand U9259 (N_9259,N_8520,N_8710);
or U9260 (N_9260,N_8572,N_8859);
and U9261 (N_9261,N_8557,N_8505);
or U9262 (N_9262,N_8728,N_8518);
nor U9263 (N_9263,N_8895,N_8817);
nand U9264 (N_9264,N_8661,N_8781);
or U9265 (N_9265,N_8712,N_8520);
xnor U9266 (N_9266,N_8547,N_8928);
nor U9267 (N_9267,N_8983,N_8896);
nand U9268 (N_9268,N_8723,N_8963);
nor U9269 (N_9269,N_8904,N_8585);
or U9270 (N_9270,N_8989,N_8949);
or U9271 (N_9271,N_8852,N_8578);
xnor U9272 (N_9272,N_8623,N_8528);
nor U9273 (N_9273,N_8816,N_8985);
or U9274 (N_9274,N_8884,N_8657);
and U9275 (N_9275,N_8858,N_8792);
nand U9276 (N_9276,N_8869,N_8731);
or U9277 (N_9277,N_8767,N_8667);
or U9278 (N_9278,N_8870,N_8927);
nor U9279 (N_9279,N_8729,N_8669);
nor U9280 (N_9280,N_8822,N_8686);
or U9281 (N_9281,N_8675,N_8534);
and U9282 (N_9282,N_8548,N_8934);
nor U9283 (N_9283,N_8832,N_8655);
and U9284 (N_9284,N_8547,N_8750);
and U9285 (N_9285,N_8666,N_8872);
and U9286 (N_9286,N_8966,N_8558);
or U9287 (N_9287,N_8813,N_8890);
or U9288 (N_9288,N_8753,N_8696);
nand U9289 (N_9289,N_8776,N_8827);
and U9290 (N_9290,N_8926,N_8510);
or U9291 (N_9291,N_8911,N_8864);
nand U9292 (N_9292,N_8644,N_8804);
and U9293 (N_9293,N_8533,N_8890);
and U9294 (N_9294,N_8785,N_8855);
xor U9295 (N_9295,N_8962,N_8664);
and U9296 (N_9296,N_8744,N_8939);
nor U9297 (N_9297,N_8551,N_8523);
or U9298 (N_9298,N_8936,N_8711);
or U9299 (N_9299,N_8801,N_8846);
or U9300 (N_9300,N_8670,N_8994);
or U9301 (N_9301,N_8864,N_8603);
and U9302 (N_9302,N_8580,N_8649);
nand U9303 (N_9303,N_8951,N_8722);
nor U9304 (N_9304,N_8506,N_8840);
or U9305 (N_9305,N_8947,N_8743);
or U9306 (N_9306,N_8821,N_8551);
and U9307 (N_9307,N_8536,N_8528);
nand U9308 (N_9308,N_8718,N_8622);
nor U9309 (N_9309,N_8998,N_8504);
nand U9310 (N_9310,N_8950,N_8795);
nor U9311 (N_9311,N_8747,N_8876);
and U9312 (N_9312,N_8752,N_8861);
nand U9313 (N_9313,N_8810,N_8770);
nor U9314 (N_9314,N_8915,N_8891);
nor U9315 (N_9315,N_8706,N_8683);
nand U9316 (N_9316,N_8751,N_8804);
nor U9317 (N_9317,N_8767,N_8546);
and U9318 (N_9318,N_8930,N_8894);
or U9319 (N_9319,N_8997,N_8930);
or U9320 (N_9320,N_8548,N_8637);
and U9321 (N_9321,N_8743,N_8649);
and U9322 (N_9322,N_8958,N_8884);
nor U9323 (N_9323,N_8676,N_8659);
nand U9324 (N_9324,N_8782,N_8756);
or U9325 (N_9325,N_8842,N_8802);
and U9326 (N_9326,N_8909,N_8865);
or U9327 (N_9327,N_8714,N_8992);
nor U9328 (N_9328,N_8997,N_8604);
nor U9329 (N_9329,N_8656,N_8633);
nand U9330 (N_9330,N_8648,N_8965);
nor U9331 (N_9331,N_8855,N_8682);
nand U9332 (N_9332,N_8503,N_8914);
nand U9333 (N_9333,N_8642,N_8760);
nor U9334 (N_9334,N_8849,N_8721);
nand U9335 (N_9335,N_8903,N_8577);
or U9336 (N_9336,N_8815,N_8681);
nor U9337 (N_9337,N_8788,N_8670);
nor U9338 (N_9338,N_8931,N_8669);
nand U9339 (N_9339,N_8577,N_8633);
nor U9340 (N_9340,N_8940,N_8681);
and U9341 (N_9341,N_8799,N_8598);
and U9342 (N_9342,N_8896,N_8528);
nor U9343 (N_9343,N_8766,N_8857);
or U9344 (N_9344,N_8779,N_8810);
or U9345 (N_9345,N_8667,N_8842);
or U9346 (N_9346,N_8878,N_8824);
or U9347 (N_9347,N_8886,N_8919);
nand U9348 (N_9348,N_8690,N_8583);
nor U9349 (N_9349,N_8915,N_8694);
nor U9350 (N_9350,N_8718,N_8877);
nor U9351 (N_9351,N_8733,N_8763);
nand U9352 (N_9352,N_8732,N_8752);
nand U9353 (N_9353,N_8925,N_8751);
and U9354 (N_9354,N_8721,N_8976);
or U9355 (N_9355,N_8696,N_8502);
and U9356 (N_9356,N_8957,N_8819);
nand U9357 (N_9357,N_8602,N_8667);
and U9358 (N_9358,N_8653,N_8882);
nand U9359 (N_9359,N_8574,N_8505);
xor U9360 (N_9360,N_8851,N_8658);
and U9361 (N_9361,N_8690,N_8785);
or U9362 (N_9362,N_8541,N_8656);
nand U9363 (N_9363,N_8921,N_8972);
or U9364 (N_9364,N_8737,N_8646);
and U9365 (N_9365,N_8792,N_8937);
and U9366 (N_9366,N_8657,N_8753);
or U9367 (N_9367,N_8730,N_8790);
and U9368 (N_9368,N_8797,N_8653);
nand U9369 (N_9369,N_8554,N_8682);
nor U9370 (N_9370,N_8559,N_8549);
and U9371 (N_9371,N_8925,N_8698);
or U9372 (N_9372,N_8526,N_8936);
and U9373 (N_9373,N_8875,N_8673);
nand U9374 (N_9374,N_8699,N_8920);
or U9375 (N_9375,N_8981,N_8641);
or U9376 (N_9376,N_8904,N_8725);
nand U9377 (N_9377,N_8670,N_8913);
or U9378 (N_9378,N_8542,N_8784);
or U9379 (N_9379,N_8666,N_8633);
nand U9380 (N_9380,N_8744,N_8958);
or U9381 (N_9381,N_8652,N_8641);
nand U9382 (N_9382,N_8613,N_8688);
and U9383 (N_9383,N_8661,N_8692);
nor U9384 (N_9384,N_8629,N_8782);
or U9385 (N_9385,N_8860,N_8698);
or U9386 (N_9386,N_8995,N_8841);
xor U9387 (N_9387,N_8658,N_8635);
nor U9388 (N_9388,N_8927,N_8894);
and U9389 (N_9389,N_8963,N_8760);
and U9390 (N_9390,N_8895,N_8600);
and U9391 (N_9391,N_8800,N_8920);
and U9392 (N_9392,N_8986,N_8881);
nand U9393 (N_9393,N_8772,N_8525);
and U9394 (N_9394,N_8670,N_8781);
and U9395 (N_9395,N_8712,N_8608);
nand U9396 (N_9396,N_8765,N_8675);
nand U9397 (N_9397,N_8959,N_8761);
nand U9398 (N_9398,N_8757,N_8625);
nand U9399 (N_9399,N_8779,N_8978);
or U9400 (N_9400,N_8548,N_8602);
nor U9401 (N_9401,N_8819,N_8996);
and U9402 (N_9402,N_8687,N_8746);
nand U9403 (N_9403,N_8996,N_8802);
and U9404 (N_9404,N_8757,N_8928);
nor U9405 (N_9405,N_8844,N_8777);
nor U9406 (N_9406,N_8770,N_8728);
nor U9407 (N_9407,N_8792,N_8784);
nor U9408 (N_9408,N_8825,N_8510);
nor U9409 (N_9409,N_8823,N_8525);
and U9410 (N_9410,N_8789,N_8646);
or U9411 (N_9411,N_8532,N_8988);
nand U9412 (N_9412,N_8706,N_8984);
and U9413 (N_9413,N_8771,N_8584);
or U9414 (N_9414,N_8980,N_8948);
nor U9415 (N_9415,N_8902,N_8958);
nor U9416 (N_9416,N_8690,N_8599);
xnor U9417 (N_9417,N_8605,N_8760);
nand U9418 (N_9418,N_8979,N_8898);
xnor U9419 (N_9419,N_8698,N_8737);
nor U9420 (N_9420,N_8666,N_8655);
and U9421 (N_9421,N_8600,N_8616);
or U9422 (N_9422,N_8861,N_8700);
nand U9423 (N_9423,N_8816,N_8612);
and U9424 (N_9424,N_8566,N_8870);
nand U9425 (N_9425,N_8893,N_8698);
or U9426 (N_9426,N_8514,N_8839);
or U9427 (N_9427,N_8773,N_8980);
nor U9428 (N_9428,N_8660,N_8528);
and U9429 (N_9429,N_8872,N_8772);
xnor U9430 (N_9430,N_8506,N_8969);
nor U9431 (N_9431,N_8708,N_8944);
or U9432 (N_9432,N_8586,N_8860);
or U9433 (N_9433,N_8776,N_8788);
nand U9434 (N_9434,N_8637,N_8792);
nor U9435 (N_9435,N_8559,N_8769);
nor U9436 (N_9436,N_8567,N_8911);
nand U9437 (N_9437,N_8663,N_8673);
nand U9438 (N_9438,N_8526,N_8548);
and U9439 (N_9439,N_8700,N_8782);
or U9440 (N_9440,N_8700,N_8622);
nand U9441 (N_9441,N_8635,N_8629);
nand U9442 (N_9442,N_8801,N_8700);
and U9443 (N_9443,N_8968,N_8639);
nand U9444 (N_9444,N_8815,N_8709);
nor U9445 (N_9445,N_8871,N_8834);
and U9446 (N_9446,N_8721,N_8540);
nor U9447 (N_9447,N_8603,N_8759);
nor U9448 (N_9448,N_8553,N_8733);
and U9449 (N_9449,N_8765,N_8936);
nor U9450 (N_9450,N_8969,N_8940);
and U9451 (N_9451,N_8539,N_8599);
or U9452 (N_9452,N_8865,N_8830);
nand U9453 (N_9453,N_8792,N_8541);
or U9454 (N_9454,N_8704,N_8700);
nand U9455 (N_9455,N_8935,N_8562);
or U9456 (N_9456,N_8508,N_8912);
nand U9457 (N_9457,N_8582,N_8969);
or U9458 (N_9458,N_8936,N_8856);
or U9459 (N_9459,N_8868,N_8834);
nor U9460 (N_9460,N_8795,N_8600);
or U9461 (N_9461,N_8513,N_8922);
nor U9462 (N_9462,N_8975,N_8866);
or U9463 (N_9463,N_8857,N_8859);
or U9464 (N_9464,N_8542,N_8722);
or U9465 (N_9465,N_8727,N_8812);
nor U9466 (N_9466,N_8603,N_8995);
nand U9467 (N_9467,N_8976,N_8980);
nor U9468 (N_9468,N_8741,N_8552);
nand U9469 (N_9469,N_8783,N_8803);
nor U9470 (N_9470,N_8748,N_8672);
nor U9471 (N_9471,N_8921,N_8708);
and U9472 (N_9472,N_8685,N_8675);
nand U9473 (N_9473,N_8553,N_8508);
nand U9474 (N_9474,N_8954,N_8521);
nor U9475 (N_9475,N_8803,N_8734);
and U9476 (N_9476,N_8750,N_8523);
and U9477 (N_9477,N_8634,N_8955);
nand U9478 (N_9478,N_8989,N_8887);
and U9479 (N_9479,N_8540,N_8808);
nor U9480 (N_9480,N_8673,N_8741);
or U9481 (N_9481,N_8537,N_8838);
and U9482 (N_9482,N_8710,N_8987);
or U9483 (N_9483,N_8609,N_8625);
nand U9484 (N_9484,N_8773,N_8698);
or U9485 (N_9485,N_8958,N_8914);
and U9486 (N_9486,N_8696,N_8651);
nor U9487 (N_9487,N_8556,N_8937);
or U9488 (N_9488,N_8740,N_8913);
nor U9489 (N_9489,N_8896,N_8780);
or U9490 (N_9490,N_8532,N_8767);
or U9491 (N_9491,N_8652,N_8562);
nor U9492 (N_9492,N_8605,N_8971);
or U9493 (N_9493,N_8795,N_8837);
nand U9494 (N_9494,N_8707,N_8865);
or U9495 (N_9495,N_8770,N_8753);
and U9496 (N_9496,N_8969,N_8674);
nor U9497 (N_9497,N_8650,N_8527);
nor U9498 (N_9498,N_8533,N_8711);
and U9499 (N_9499,N_8505,N_8641);
and U9500 (N_9500,N_9292,N_9468);
nor U9501 (N_9501,N_9391,N_9210);
and U9502 (N_9502,N_9484,N_9382);
or U9503 (N_9503,N_9365,N_9067);
and U9504 (N_9504,N_9122,N_9386);
nand U9505 (N_9505,N_9147,N_9070);
and U9506 (N_9506,N_9061,N_9306);
and U9507 (N_9507,N_9201,N_9102);
and U9508 (N_9508,N_9499,N_9463);
nand U9509 (N_9509,N_9334,N_9166);
and U9510 (N_9510,N_9310,N_9174);
nor U9511 (N_9511,N_9389,N_9221);
or U9512 (N_9512,N_9280,N_9426);
and U9513 (N_9513,N_9349,N_9316);
or U9514 (N_9514,N_9400,N_9282);
and U9515 (N_9515,N_9408,N_9084);
or U9516 (N_9516,N_9062,N_9225);
nor U9517 (N_9517,N_9248,N_9134);
or U9518 (N_9518,N_9112,N_9305);
nand U9519 (N_9519,N_9214,N_9233);
nor U9520 (N_9520,N_9157,N_9039);
nand U9521 (N_9521,N_9051,N_9080);
nand U9522 (N_9522,N_9317,N_9371);
and U9523 (N_9523,N_9375,N_9286);
or U9524 (N_9524,N_9268,N_9454);
nor U9525 (N_9525,N_9000,N_9381);
or U9526 (N_9526,N_9186,N_9226);
nand U9527 (N_9527,N_9362,N_9396);
nand U9528 (N_9528,N_9260,N_9239);
nor U9529 (N_9529,N_9103,N_9151);
nand U9530 (N_9530,N_9066,N_9133);
xnor U9531 (N_9531,N_9496,N_9483);
nand U9532 (N_9532,N_9207,N_9485);
nor U9533 (N_9533,N_9262,N_9372);
nor U9534 (N_9534,N_9418,N_9155);
or U9535 (N_9535,N_9290,N_9064);
nor U9536 (N_9536,N_9115,N_9342);
nor U9537 (N_9537,N_9321,N_9318);
or U9538 (N_9538,N_9407,N_9406);
and U9539 (N_9539,N_9459,N_9030);
and U9540 (N_9540,N_9356,N_9377);
or U9541 (N_9541,N_9093,N_9337);
or U9542 (N_9542,N_9163,N_9470);
nand U9543 (N_9543,N_9419,N_9118);
nand U9544 (N_9544,N_9440,N_9191);
nor U9545 (N_9545,N_9096,N_9224);
or U9546 (N_9546,N_9312,N_9117);
nor U9547 (N_9547,N_9417,N_9143);
or U9548 (N_9548,N_9244,N_9465);
nor U9549 (N_9549,N_9263,N_9431);
xor U9550 (N_9550,N_9104,N_9462);
nand U9551 (N_9551,N_9355,N_9179);
or U9552 (N_9552,N_9299,N_9083);
nor U9553 (N_9553,N_9475,N_9363);
nand U9554 (N_9554,N_9241,N_9235);
xnor U9555 (N_9555,N_9467,N_9351);
nand U9556 (N_9556,N_9136,N_9002);
or U9557 (N_9557,N_9183,N_9343);
and U9558 (N_9558,N_9314,N_9124);
or U9559 (N_9559,N_9116,N_9199);
nand U9560 (N_9560,N_9437,N_9211);
nand U9561 (N_9561,N_9283,N_9111);
and U9562 (N_9562,N_9326,N_9411);
and U9563 (N_9563,N_9410,N_9079);
nand U9564 (N_9564,N_9482,N_9088);
and U9565 (N_9565,N_9204,N_9229);
and U9566 (N_9566,N_9228,N_9378);
and U9567 (N_9567,N_9161,N_9087);
or U9568 (N_9568,N_9255,N_9453);
nand U9569 (N_9569,N_9150,N_9421);
nand U9570 (N_9570,N_9187,N_9276);
nand U9571 (N_9571,N_9497,N_9340);
nand U9572 (N_9572,N_9059,N_9285);
and U9573 (N_9573,N_9189,N_9309);
nor U9574 (N_9574,N_9298,N_9450);
or U9575 (N_9575,N_9395,N_9455);
or U9576 (N_9576,N_9113,N_9250);
nor U9577 (N_9577,N_9234,N_9322);
and U9578 (N_9578,N_9106,N_9324);
nor U9579 (N_9579,N_9137,N_9142);
or U9580 (N_9580,N_9020,N_9486);
nor U9581 (N_9581,N_9361,N_9054);
and U9582 (N_9582,N_9416,N_9045);
nor U9583 (N_9583,N_9456,N_9008);
nand U9584 (N_9584,N_9085,N_9293);
or U9585 (N_9585,N_9141,N_9279);
nand U9586 (N_9586,N_9217,N_9493);
and U9587 (N_9587,N_9458,N_9041);
nand U9588 (N_9588,N_9368,N_9056);
and U9589 (N_9589,N_9238,N_9190);
nand U9590 (N_9590,N_9320,N_9350);
xor U9591 (N_9591,N_9315,N_9009);
xnor U9592 (N_9592,N_9101,N_9025);
nor U9593 (N_9593,N_9478,N_9197);
and U9594 (N_9594,N_9153,N_9266);
nand U9595 (N_9595,N_9188,N_9307);
or U9596 (N_9596,N_9348,N_9127);
and U9597 (N_9597,N_9384,N_9077);
nor U9598 (N_9598,N_9376,N_9432);
and U9599 (N_9599,N_9247,N_9004);
nand U9600 (N_9600,N_9215,N_9222);
and U9601 (N_9601,N_9075,N_9249);
and U9602 (N_9602,N_9434,N_9379);
nor U9603 (N_9603,N_9178,N_9231);
and U9604 (N_9604,N_9369,N_9325);
nand U9605 (N_9605,N_9028,N_9130);
nor U9606 (N_9606,N_9071,N_9423);
and U9607 (N_9607,N_9167,N_9273);
nor U9608 (N_9608,N_9438,N_9010);
and U9609 (N_9609,N_9086,N_9100);
or U9610 (N_9610,N_9278,N_9095);
or U9611 (N_9611,N_9200,N_9339);
xnor U9612 (N_9612,N_9311,N_9257);
nor U9613 (N_9613,N_9464,N_9401);
and U9614 (N_9614,N_9441,N_9335);
and U9615 (N_9615,N_9284,N_9412);
nor U9616 (N_9616,N_9413,N_9073);
nand U9617 (N_9617,N_9494,N_9352);
nand U9618 (N_9618,N_9404,N_9331);
or U9619 (N_9619,N_9380,N_9182);
nand U9620 (N_9620,N_9001,N_9390);
or U9621 (N_9621,N_9345,N_9338);
and U9622 (N_9622,N_9265,N_9259);
nand U9623 (N_9623,N_9258,N_9146);
or U9624 (N_9624,N_9037,N_9357);
and U9625 (N_9625,N_9366,N_9439);
and U9626 (N_9626,N_9203,N_9367);
nor U9627 (N_9627,N_9253,N_9281);
nand U9628 (N_9628,N_9295,N_9415);
nor U9629 (N_9629,N_9358,N_9135);
nand U9630 (N_9630,N_9081,N_9303);
and U9631 (N_9631,N_9333,N_9196);
nor U9632 (N_9632,N_9192,N_9202);
nand U9633 (N_9633,N_9168,N_9240);
or U9634 (N_9634,N_9060,N_9429);
nand U9635 (N_9635,N_9033,N_9125);
nand U9636 (N_9636,N_9430,N_9492);
nor U9637 (N_9637,N_9016,N_9294);
xor U9638 (N_9638,N_9193,N_9383);
or U9639 (N_9639,N_9435,N_9107);
xnor U9640 (N_9640,N_9344,N_9402);
and U9641 (N_9641,N_9154,N_9021);
or U9642 (N_9642,N_9302,N_9047);
or U9643 (N_9643,N_9121,N_9422);
or U9644 (N_9644,N_9232,N_9110);
nor U9645 (N_9645,N_9068,N_9313);
nor U9646 (N_9646,N_9144,N_9319);
or U9647 (N_9647,N_9145,N_9223);
nor U9648 (N_9648,N_9354,N_9252);
nand U9649 (N_9649,N_9291,N_9181);
and U9650 (N_9650,N_9105,N_9148);
nand U9651 (N_9651,N_9092,N_9267);
and U9652 (N_9652,N_9022,N_9172);
nand U9653 (N_9653,N_9013,N_9444);
or U9654 (N_9654,N_9449,N_9393);
nand U9655 (N_9655,N_9029,N_9392);
and U9656 (N_9656,N_9304,N_9397);
or U9657 (N_9657,N_9387,N_9328);
and U9658 (N_9658,N_9332,N_9409);
nand U9659 (N_9659,N_9140,N_9341);
nor U9660 (N_9660,N_9212,N_9473);
and U9661 (N_9661,N_9198,N_9176);
and U9662 (N_9662,N_9003,N_9152);
nand U9663 (N_9663,N_9058,N_9452);
nand U9664 (N_9664,N_9461,N_9065);
nor U9665 (N_9665,N_9156,N_9094);
nor U9666 (N_9666,N_9180,N_9035);
nand U9667 (N_9667,N_9126,N_9169);
and U9668 (N_9668,N_9477,N_9006);
nor U9669 (N_9669,N_9300,N_9398);
and U9670 (N_9670,N_9194,N_9012);
nor U9671 (N_9671,N_9242,N_9296);
xor U9672 (N_9672,N_9011,N_9427);
or U9673 (N_9673,N_9405,N_9472);
nor U9674 (N_9674,N_9287,N_9443);
and U9675 (N_9675,N_9275,N_9120);
nand U9676 (N_9676,N_9347,N_9005);
and U9677 (N_9677,N_9481,N_9097);
nor U9678 (N_9678,N_9019,N_9032);
and U9679 (N_9679,N_9165,N_9460);
and U9680 (N_9680,N_9479,N_9251);
or U9681 (N_9681,N_9446,N_9206);
nor U9682 (N_9682,N_9098,N_9270);
and U9683 (N_9683,N_9243,N_9129);
nor U9684 (N_9684,N_9036,N_9254);
or U9685 (N_9685,N_9170,N_9445);
nand U9686 (N_9686,N_9425,N_9327);
or U9687 (N_9687,N_9399,N_9288);
nor U9688 (N_9688,N_9131,N_9216);
or U9689 (N_9689,N_9428,N_9164);
nor U9690 (N_9690,N_9230,N_9218);
xnor U9691 (N_9691,N_9301,N_9271);
or U9692 (N_9692,N_9274,N_9074);
and U9693 (N_9693,N_9323,N_9031);
or U9694 (N_9694,N_9027,N_9414);
nand U9695 (N_9695,N_9420,N_9034);
nor U9696 (N_9696,N_9160,N_9237);
or U9697 (N_9697,N_9448,N_9123);
and U9698 (N_9698,N_9469,N_9490);
and U9699 (N_9699,N_9272,N_9289);
nand U9700 (N_9700,N_9044,N_9388);
and U9701 (N_9701,N_9132,N_9208);
nor U9702 (N_9702,N_9209,N_9374);
and U9703 (N_9703,N_9043,N_9076);
or U9704 (N_9704,N_9480,N_9119);
nand U9705 (N_9705,N_9040,N_9474);
nand U9706 (N_9706,N_9042,N_9346);
or U9707 (N_9707,N_9336,N_9488);
and U9708 (N_9708,N_9359,N_9205);
nor U9709 (N_9709,N_9353,N_9329);
nand U9710 (N_9710,N_9017,N_9023);
nand U9711 (N_9711,N_9385,N_9063);
or U9712 (N_9712,N_9466,N_9246);
nor U9713 (N_9713,N_9007,N_9403);
or U9714 (N_9714,N_9308,N_9269);
or U9715 (N_9715,N_9495,N_9370);
and U9716 (N_9716,N_9360,N_9089);
nand U9717 (N_9717,N_9139,N_9213);
nand U9718 (N_9718,N_9261,N_9159);
nand U9719 (N_9719,N_9436,N_9114);
or U9720 (N_9720,N_9069,N_9277);
and U9721 (N_9721,N_9072,N_9082);
nor U9722 (N_9722,N_9018,N_9149);
and U9723 (N_9723,N_9108,N_9055);
nor U9724 (N_9724,N_9185,N_9220);
or U9725 (N_9725,N_9219,N_9498);
and U9726 (N_9726,N_9256,N_9038);
and U9727 (N_9727,N_9173,N_9090);
xnor U9728 (N_9728,N_9447,N_9091);
and U9729 (N_9729,N_9373,N_9109);
and U9730 (N_9730,N_9158,N_9184);
or U9731 (N_9731,N_9433,N_9491);
nand U9732 (N_9732,N_9424,N_9195);
and U9733 (N_9733,N_9364,N_9245);
nand U9734 (N_9734,N_9177,N_9046);
nor U9735 (N_9735,N_9471,N_9024);
or U9736 (N_9736,N_9476,N_9138);
nor U9737 (N_9737,N_9171,N_9099);
nand U9738 (N_9738,N_9264,N_9227);
nor U9739 (N_9739,N_9052,N_9451);
or U9740 (N_9740,N_9050,N_9297);
or U9741 (N_9741,N_9057,N_9489);
and U9742 (N_9742,N_9078,N_9330);
or U9743 (N_9743,N_9394,N_9162);
and U9744 (N_9744,N_9457,N_9014);
or U9745 (N_9745,N_9442,N_9053);
nor U9746 (N_9746,N_9015,N_9026);
nor U9747 (N_9747,N_9048,N_9049);
nor U9748 (N_9748,N_9175,N_9487);
or U9749 (N_9749,N_9128,N_9236);
nor U9750 (N_9750,N_9392,N_9389);
and U9751 (N_9751,N_9270,N_9453);
or U9752 (N_9752,N_9464,N_9023);
nor U9753 (N_9753,N_9291,N_9423);
and U9754 (N_9754,N_9123,N_9409);
nand U9755 (N_9755,N_9256,N_9320);
or U9756 (N_9756,N_9197,N_9255);
nor U9757 (N_9757,N_9047,N_9223);
nand U9758 (N_9758,N_9027,N_9332);
xnor U9759 (N_9759,N_9019,N_9480);
and U9760 (N_9760,N_9446,N_9472);
nor U9761 (N_9761,N_9060,N_9226);
or U9762 (N_9762,N_9351,N_9427);
nor U9763 (N_9763,N_9117,N_9345);
or U9764 (N_9764,N_9460,N_9243);
nor U9765 (N_9765,N_9110,N_9195);
nand U9766 (N_9766,N_9244,N_9212);
nor U9767 (N_9767,N_9364,N_9084);
and U9768 (N_9768,N_9392,N_9485);
nor U9769 (N_9769,N_9161,N_9386);
nor U9770 (N_9770,N_9211,N_9442);
nand U9771 (N_9771,N_9455,N_9042);
nand U9772 (N_9772,N_9496,N_9355);
or U9773 (N_9773,N_9098,N_9353);
and U9774 (N_9774,N_9339,N_9288);
or U9775 (N_9775,N_9391,N_9113);
and U9776 (N_9776,N_9245,N_9194);
and U9777 (N_9777,N_9158,N_9105);
or U9778 (N_9778,N_9050,N_9408);
nor U9779 (N_9779,N_9356,N_9195);
nor U9780 (N_9780,N_9019,N_9466);
nor U9781 (N_9781,N_9420,N_9405);
or U9782 (N_9782,N_9185,N_9138);
or U9783 (N_9783,N_9470,N_9422);
nor U9784 (N_9784,N_9018,N_9261);
or U9785 (N_9785,N_9030,N_9352);
nand U9786 (N_9786,N_9085,N_9452);
or U9787 (N_9787,N_9159,N_9027);
or U9788 (N_9788,N_9002,N_9067);
or U9789 (N_9789,N_9390,N_9443);
and U9790 (N_9790,N_9146,N_9164);
or U9791 (N_9791,N_9138,N_9469);
nor U9792 (N_9792,N_9415,N_9090);
or U9793 (N_9793,N_9103,N_9257);
nor U9794 (N_9794,N_9225,N_9396);
nor U9795 (N_9795,N_9277,N_9480);
nor U9796 (N_9796,N_9183,N_9260);
nand U9797 (N_9797,N_9139,N_9245);
or U9798 (N_9798,N_9160,N_9490);
and U9799 (N_9799,N_9044,N_9145);
or U9800 (N_9800,N_9194,N_9321);
nand U9801 (N_9801,N_9078,N_9280);
and U9802 (N_9802,N_9259,N_9116);
xor U9803 (N_9803,N_9107,N_9347);
or U9804 (N_9804,N_9258,N_9055);
or U9805 (N_9805,N_9016,N_9363);
nor U9806 (N_9806,N_9336,N_9478);
nand U9807 (N_9807,N_9096,N_9001);
or U9808 (N_9808,N_9363,N_9464);
and U9809 (N_9809,N_9477,N_9157);
nand U9810 (N_9810,N_9264,N_9297);
nor U9811 (N_9811,N_9370,N_9081);
or U9812 (N_9812,N_9100,N_9247);
and U9813 (N_9813,N_9046,N_9182);
and U9814 (N_9814,N_9226,N_9110);
and U9815 (N_9815,N_9067,N_9215);
nand U9816 (N_9816,N_9360,N_9291);
and U9817 (N_9817,N_9156,N_9358);
or U9818 (N_9818,N_9004,N_9246);
nand U9819 (N_9819,N_9361,N_9464);
or U9820 (N_9820,N_9259,N_9088);
and U9821 (N_9821,N_9204,N_9218);
and U9822 (N_9822,N_9165,N_9472);
xnor U9823 (N_9823,N_9175,N_9348);
nor U9824 (N_9824,N_9242,N_9357);
nor U9825 (N_9825,N_9176,N_9059);
and U9826 (N_9826,N_9041,N_9111);
nand U9827 (N_9827,N_9108,N_9244);
nand U9828 (N_9828,N_9196,N_9036);
nor U9829 (N_9829,N_9003,N_9466);
and U9830 (N_9830,N_9017,N_9106);
xor U9831 (N_9831,N_9180,N_9154);
nor U9832 (N_9832,N_9123,N_9273);
and U9833 (N_9833,N_9154,N_9129);
nor U9834 (N_9834,N_9409,N_9349);
and U9835 (N_9835,N_9115,N_9046);
or U9836 (N_9836,N_9349,N_9024);
nor U9837 (N_9837,N_9212,N_9000);
or U9838 (N_9838,N_9047,N_9039);
or U9839 (N_9839,N_9278,N_9447);
nor U9840 (N_9840,N_9019,N_9418);
nor U9841 (N_9841,N_9016,N_9329);
nand U9842 (N_9842,N_9259,N_9330);
nand U9843 (N_9843,N_9466,N_9125);
nor U9844 (N_9844,N_9467,N_9212);
nand U9845 (N_9845,N_9119,N_9127);
and U9846 (N_9846,N_9116,N_9366);
and U9847 (N_9847,N_9343,N_9040);
or U9848 (N_9848,N_9394,N_9181);
or U9849 (N_9849,N_9362,N_9199);
nor U9850 (N_9850,N_9208,N_9162);
or U9851 (N_9851,N_9313,N_9060);
nor U9852 (N_9852,N_9448,N_9137);
and U9853 (N_9853,N_9156,N_9169);
xor U9854 (N_9854,N_9118,N_9354);
nand U9855 (N_9855,N_9078,N_9193);
or U9856 (N_9856,N_9338,N_9334);
nor U9857 (N_9857,N_9078,N_9255);
and U9858 (N_9858,N_9093,N_9356);
nand U9859 (N_9859,N_9016,N_9105);
or U9860 (N_9860,N_9330,N_9004);
or U9861 (N_9861,N_9090,N_9283);
nand U9862 (N_9862,N_9233,N_9035);
or U9863 (N_9863,N_9063,N_9206);
or U9864 (N_9864,N_9380,N_9344);
nand U9865 (N_9865,N_9194,N_9401);
nor U9866 (N_9866,N_9335,N_9381);
and U9867 (N_9867,N_9378,N_9190);
and U9868 (N_9868,N_9149,N_9098);
nor U9869 (N_9869,N_9351,N_9456);
or U9870 (N_9870,N_9206,N_9046);
xnor U9871 (N_9871,N_9364,N_9305);
and U9872 (N_9872,N_9357,N_9341);
nor U9873 (N_9873,N_9209,N_9076);
or U9874 (N_9874,N_9443,N_9349);
nor U9875 (N_9875,N_9385,N_9119);
or U9876 (N_9876,N_9440,N_9240);
nand U9877 (N_9877,N_9088,N_9461);
nand U9878 (N_9878,N_9225,N_9091);
nor U9879 (N_9879,N_9139,N_9495);
nand U9880 (N_9880,N_9204,N_9375);
nor U9881 (N_9881,N_9439,N_9155);
or U9882 (N_9882,N_9076,N_9482);
nand U9883 (N_9883,N_9313,N_9363);
nand U9884 (N_9884,N_9079,N_9418);
or U9885 (N_9885,N_9228,N_9453);
nor U9886 (N_9886,N_9127,N_9269);
nor U9887 (N_9887,N_9050,N_9038);
or U9888 (N_9888,N_9154,N_9472);
nor U9889 (N_9889,N_9166,N_9061);
nand U9890 (N_9890,N_9114,N_9200);
nor U9891 (N_9891,N_9022,N_9448);
and U9892 (N_9892,N_9140,N_9488);
nor U9893 (N_9893,N_9209,N_9206);
nand U9894 (N_9894,N_9111,N_9472);
or U9895 (N_9895,N_9493,N_9059);
or U9896 (N_9896,N_9440,N_9145);
or U9897 (N_9897,N_9179,N_9302);
nor U9898 (N_9898,N_9448,N_9277);
nand U9899 (N_9899,N_9327,N_9397);
and U9900 (N_9900,N_9342,N_9425);
or U9901 (N_9901,N_9275,N_9136);
nand U9902 (N_9902,N_9325,N_9326);
or U9903 (N_9903,N_9476,N_9150);
and U9904 (N_9904,N_9133,N_9411);
nand U9905 (N_9905,N_9204,N_9339);
or U9906 (N_9906,N_9485,N_9294);
or U9907 (N_9907,N_9286,N_9006);
nand U9908 (N_9908,N_9356,N_9447);
and U9909 (N_9909,N_9447,N_9436);
nor U9910 (N_9910,N_9482,N_9052);
and U9911 (N_9911,N_9373,N_9216);
or U9912 (N_9912,N_9264,N_9018);
and U9913 (N_9913,N_9296,N_9294);
nand U9914 (N_9914,N_9085,N_9188);
nor U9915 (N_9915,N_9211,N_9015);
nor U9916 (N_9916,N_9376,N_9139);
or U9917 (N_9917,N_9396,N_9435);
xnor U9918 (N_9918,N_9322,N_9267);
nand U9919 (N_9919,N_9071,N_9421);
nand U9920 (N_9920,N_9238,N_9428);
nand U9921 (N_9921,N_9257,N_9084);
nor U9922 (N_9922,N_9343,N_9241);
nor U9923 (N_9923,N_9301,N_9247);
and U9924 (N_9924,N_9499,N_9144);
nor U9925 (N_9925,N_9347,N_9474);
nor U9926 (N_9926,N_9449,N_9082);
nor U9927 (N_9927,N_9018,N_9389);
or U9928 (N_9928,N_9044,N_9426);
nor U9929 (N_9929,N_9032,N_9474);
nand U9930 (N_9930,N_9136,N_9381);
and U9931 (N_9931,N_9119,N_9424);
or U9932 (N_9932,N_9392,N_9062);
nand U9933 (N_9933,N_9392,N_9171);
and U9934 (N_9934,N_9256,N_9185);
nor U9935 (N_9935,N_9241,N_9356);
nand U9936 (N_9936,N_9262,N_9156);
and U9937 (N_9937,N_9104,N_9321);
nor U9938 (N_9938,N_9156,N_9457);
nor U9939 (N_9939,N_9102,N_9361);
nand U9940 (N_9940,N_9374,N_9219);
or U9941 (N_9941,N_9293,N_9031);
nor U9942 (N_9942,N_9097,N_9124);
or U9943 (N_9943,N_9035,N_9317);
nand U9944 (N_9944,N_9473,N_9129);
or U9945 (N_9945,N_9165,N_9267);
and U9946 (N_9946,N_9424,N_9144);
or U9947 (N_9947,N_9180,N_9026);
or U9948 (N_9948,N_9061,N_9375);
or U9949 (N_9949,N_9111,N_9212);
and U9950 (N_9950,N_9272,N_9048);
nor U9951 (N_9951,N_9310,N_9429);
or U9952 (N_9952,N_9118,N_9156);
or U9953 (N_9953,N_9467,N_9162);
or U9954 (N_9954,N_9382,N_9043);
xor U9955 (N_9955,N_9461,N_9307);
nand U9956 (N_9956,N_9347,N_9153);
nor U9957 (N_9957,N_9059,N_9319);
and U9958 (N_9958,N_9051,N_9282);
nand U9959 (N_9959,N_9198,N_9330);
nand U9960 (N_9960,N_9266,N_9381);
and U9961 (N_9961,N_9489,N_9100);
nand U9962 (N_9962,N_9444,N_9348);
nand U9963 (N_9963,N_9363,N_9012);
nor U9964 (N_9964,N_9430,N_9024);
nor U9965 (N_9965,N_9440,N_9438);
nand U9966 (N_9966,N_9083,N_9448);
and U9967 (N_9967,N_9124,N_9235);
and U9968 (N_9968,N_9034,N_9078);
nand U9969 (N_9969,N_9339,N_9135);
and U9970 (N_9970,N_9051,N_9191);
or U9971 (N_9971,N_9117,N_9285);
nor U9972 (N_9972,N_9114,N_9265);
nand U9973 (N_9973,N_9049,N_9353);
xnor U9974 (N_9974,N_9349,N_9262);
and U9975 (N_9975,N_9374,N_9141);
nand U9976 (N_9976,N_9054,N_9276);
and U9977 (N_9977,N_9251,N_9056);
nand U9978 (N_9978,N_9065,N_9199);
and U9979 (N_9979,N_9302,N_9488);
nand U9980 (N_9980,N_9327,N_9261);
nand U9981 (N_9981,N_9368,N_9150);
and U9982 (N_9982,N_9487,N_9352);
nor U9983 (N_9983,N_9342,N_9363);
nor U9984 (N_9984,N_9175,N_9172);
and U9985 (N_9985,N_9283,N_9174);
and U9986 (N_9986,N_9425,N_9219);
nor U9987 (N_9987,N_9417,N_9088);
or U9988 (N_9988,N_9365,N_9004);
nand U9989 (N_9989,N_9191,N_9039);
and U9990 (N_9990,N_9001,N_9292);
and U9991 (N_9991,N_9169,N_9212);
and U9992 (N_9992,N_9085,N_9454);
or U9993 (N_9993,N_9233,N_9042);
nor U9994 (N_9994,N_9368,N_9137);
or U9995 (N_9995,N_9095,N_9346);
or U9996 (N_9996,N_9378,N_9172);
nor U9997 (N_9997,N_9183,N_9141);
and U9998 (N_9998,N_9090,N_9011);
nor U9999 (N_9999,N_9078,N_9220);
or UO_0 (O_0,N_9759,N_9975);
or UO_1 (O_1,N_9680,N_9754);
and UO_2 (O_2,N_9540,N_9512);
xor UO_3 (O_3,N_9600,N_9871);
and UO_4 (O_4,N_9623,N_9552);
or UO_5 (O_5,N_9706,N_9633);
and UO_6 (O_6,N_9542,N_9947);
and UO_7 (O_7,N_9539,N_9650);
nand UO_8 (O_8,N_9939,N_9955);
nor UO_9 (O_9,N_9849,N_9764);
and UO_10 (O_10,N_9991,N_9701);
nor UO_11 (O_11,N_9642,N_9836);
nor UO_12 (O_12,N_9956,N_9762);
and UO_13 (O_13,N_9570,N_9506);
nor UO_14 (O_14,N_9658,N_9949);
nor UO_15 (O_15,N_9758,N_9832);
and UO_16 (O_16,N_9692,N_9704);
nor UO_17 (O_17,N_9630,N_9860);
or UO_18 (O_18,N_9880,N_9757);
xnor UO_19 (O_19,N_9514,N_9798);
nand UO_20 (O_20,N_9502,N_9935);
and UO_21 (O_21,N_9550,N_9793);
nor UO_22 (O_22,N_9903,N_9715);
nor UO_23 (O_23,N_9978,N_9727);
nand UO_24 (O_24,N_9588,N_9675);
nor UO_25 (O_25,N_9568,N_9792);
nand UO_26 (O_26,N_9594,N_9719);
nand UO_27 (O_27,N_9609,N_9928);
or UO_28 (O_28,N_9918,N_9932);
nand UO_29 (O_29,N_9638,N_9868);
nand UO_30 (O_30,N_9522,N_9584);
nor UO_31 (O_31,N_9778,N_9553);
nand UO_32 (O_32,N_9547,N_9566);
xnor UO_33 (O_33,N_9894,N_9543);
nand UO_34 (O_34,N_9743,N_9571);
nor UO_35 (O_35,N_9614,N_9765);
nor UO_36 (O_36,N_9527,N_9523);
and UO_37 (O_37,N_9933,N_9659);
nand UO_38 (O_38,N_9740,N_9672);
and UO_39 (O_39,N_9677,N_9687);
nor UO_40 (O_40,N_9822,N_9653);
nand UO_41 (O_41,N_9603,N_9818);
or UO_42 (O_42,N_9965,N_9856);
nand UO_43 (O_43,N_9580,N_9852);
nor UO_44 (O_44,N_9707,N_9745);
nand UO_45 (O_45,N_9744,N_9877);
nor UO_46 (O_46,N_9927,N_9845);
nor UO_47 (O_47,N_9731,N_9769);
or UO_48 (O_48,N_9721,N_9673);
nor UO_49 (O_49,N_9859,N_9773);
nand UO_50 (O_50,N_9708,N_9940);
nor UO_51 (O_51,N_9901,N_9620);
xor UO_52 (O_52,N_9733,N_9801);
nor UO_53 (O_53,N_9662,N_9957);
and UO_54 (O_54,N_9914,N_9632);
nand UO_55 (O_55,N_9851,N_9612);
nor UO_56 (O_56,N_9747,N_9709);
or UO_57 (O_57,N_9627,N_9908);
and UO_58 (O_58,N_9923,N_9645);
and UO_59 (O_59,N_9775,N_9587);
nor UO_60 (O_60,N_9693,N_9924);
nor UO_61 (O_61,N_9828,N_9861);
or UO_62 (O_62,N_9814,N_9700);
nor UO_63 (O_63,N_9639,N_9511);
nor UO_64 (O_64,N_9999,N_9799);
and UO_65 (O_65,N_9628,N_9590);
nand UO_66 (O_66,N_9878,N_9994);
and UO_67 (O_67,N_9724,N_9920);
and UO_68 (O_68,N_9907,N_9886);
nand UO_69 (O_69,N_9810,N_9837);
and UO_70 (O_70,N_9870,N_9624);
or UO_71 (O_71,N_9839,N_9997);
nor UO_72 (O_72,N_9718,N_9591);
nand UO_73 (O_73,N_9616,N_9763);
nand UO_74 (O_74,N_9881,N_9528);
and UO_75 (O_75,N_9898,N_9643);
nand UO_76 (O_76,N_9986,N_9637);
or UO_77 (O_77,N_9842,N_9572);
or UO_78 (O_78,N_9711,N_9501);
or UO_79 (O_79,N_9667,N_9931);
and UO_80 (O_80,N_9507,N_9685);
or UO_81 (O_81,N_9794,N_9846);
nand UO_82 (O_82,N_9848,N_9926);
or UO_83 (O_83,N_9728,N_9951);
nor UO_84 (O_84,N_9695,N_9873);
and UO_85 (O_85,N_9517,N_9738);
and UO_86 (O_86,N_9909,N_9983);
and UO_87 (O_87,N_9649,N_9875);
or UO_88 (O_88,N_9670,N_9592);
nand UO_89 (O_89,N_9608,N_9817);
or UO_90 (O_90,N_9500,N_9884);
or UO_91 (O_91,N_9936,N_9698);
nor UO_92 (O_92,N_9644,N_9676);
and UO_93 (O_93,N_9751,N_9660);
and UO_94 (O_94,N_9558,N_9897);
or UO_95 (O_95,N_9525,N_9551);
nand UO_96 (O_96,N_9583,N_9858);
nor UO_97 (O_97,N_9554,N_9979);
and UO_98 (O_98,N_9888,N_9833);
nand UO_99 (O_99,N_9508,N_9838);
or UO_100 (O_100,N_9546,N_9705);
or UO_101 (O_101,N_9647,N_9518);
or UO_102 (O_102,N_9988,N_9651);
and UO_103 (O_103,N_9944,N_9567);
or UO_104 (O_104,N_9736,N_9879);
nand UO_105 (O_105,N_9857,N_9816);
nand UO_106 (O_106,N_9797,N_9937);
nand UO_107 (O_107,N_9661,N_9841);
and UO_108 (O_108,N_9824,N_9656);
and UO_109 (O_109,N_9786,N_9560);
or UO_110 (O_110,N_9510,N_9804);
and UO_111 (O_111,N_9809,N_9772);
or UO_112 (O_112,N_9948,N_9867);
nor UO_113 (O_113,N_9844,N_9569);
nand UO_114 (O_114,N_9722,N_9617);
and UO_115 (O_115,N_9900,N_9976);
nor UO_116 (O_116,N_9820,N_9771);
and UO_117 (O_117,N_9813,N_9941);
xnor UO_118 (O_118,N_9782,N_9938);
or UO_119 (O_119,N_9713,N_9912);
or UO_120 (O_120,N_9834,N_9779);
nor UO_121 (O_121,N_9829,N_9974);
nor UO_122 (O_122,N_9819,N_9674);
nor UO_123 (O_123,N_9619,N_9597);
nand UO_124 (O_124,N_9734,N_9712);
nand UO_125 (O_125,N_9635,N_9987);
or UO_126 (O_126,N_9812,N_9526);
nand UO_127 (O_127,N_9582,N_9530);
nand UO_128 (O_128,N_9995,N_9989);
or UO_129 (O_129,N_9690,N_9545);
nand UO_130 (O_130,N_9885,N_9827);
or UO_131 (O_131,N_9521,N_9902);
and UO_132 (O_132,N_9889,N_9689);
or UO_133 (O_133,N_9919,N_9843);
nand UO_134 (O_134,N_9893,N_9958);
and UO_135 (O_135,N_9595,N_9679);
nand UO_136 (O_136,N_9952,N_9883);
and UO_137 (O_137,N_9629,N_9576);
nand UO_138 (O_138,N_9646,N_9726);
nand UO_139 (O_139,N_9904,N_9513);
nand UO_140 (O_140,N_9921,N_9815);
nor UO_141 (O_141,N_9790,N_9648);
nor UO_142 (O_142,N_9657,N_9821);
nor UO_143 (O_143,N_9892,N_9741);
nor UO_144 (O_144,N_9548,N_9925);
nand UO_145 (O_145,N_9756,N_9800);
and UO_146 (O_146,N_9516,N_9699);
and UO_147 (O_147,N_9766,N_9618);
and UO_148 (O_148,N_9641,N_9714);
or UO_149 (O_149,N_9780,N_9961);
nand UO_150 (O_150,N_9515,N_9805);
nand UO_151 (O_151,N_9625,N_9746);
nor UO_152 (O_152,N_9929,N_9943);
nand UO_153 (O_153,N_9696,N_9795);
nand UO_154 (O_154,N_9564,N_9752);
or UO_155 (O_155,N_9990,N_9874);
nor UO_156 (O_156,N_9524,N_9964);
nand UO_157 (O_157,N_9730,N_9755);
nand UO_158 (O_158,N_9942,N_9697);
nor UO_159 (O_159,N_9579,N_9748);
nand UO_160 (O_160,N_9922,N_9787);
and UO_161 (O_161,N_9847,N_9984);
and UO_162 (O_162,N_9774,N_9574);
nor UO_163 (O_163,N_9504,N_9509);
nor UO_164 (O_164,N_9606,N_9982);
and UO_165 (O_165,N_9681,N_9575);
and UO_166 (O_166,N_9654,N_9854);
nand UO_167 (O_167,N_9945,N_9960);
nand UO_168 (O_168,N_9998,N_9622);
or UO_169 (O_169,N_9586,N_9725);
nor UO_170 (O_170,N_9864,N_9710);
or UO_171 (O_171,N_9981,N_9573);
or UO_172 (O_172,N_9593,N_9615);
and UO_173 (O_173,N_9634,N_9910);
or UO_174 (O_174,N_9581,N_9631);
or UO_175 (O_175,N_9749,N_9520);
and UO_176 (O_176,N_9876,N_9640);
nor UO_177 (O_177,N_9605,N_9808);
nor UO_178 (O_178,N_9716,N_9531);
nand UO_179 (O_179,N_9613,N_9503);
and UO_180 (O_180,N_9980,N_9544);
and UO_181 (O_181,N_9789,N_9720);
or UO_182 (O_182,N_9831,N_9535);
nand UO_183 (O_183,N_9563,N_9823);
or UO_184 (O_184,N_9686,N_9768);
or UO_185 (O_185,N_9556,N_9962);
and UO_186 (O_186,N_9652,N_9869);
and UO_187 (O_187,N_9655,N_9826);
or UO_188 (O_188,N_9565,N_9985);
or UO_189 (O_189,N_9555,N_9917);
nand UO_190 (O_190,N_9536,N_9682);
or UO_191 (O_191,N_9611,N_9862);
and UO_192 (O_192,N_9750,N_9684);
or UO_193 (O_193,N_9895,N_9806);
nand UO_194 (O_194,N_9777,N_9934);
nor UO_195 (O_195,N_9959,N_9865);
or UO_196 (O_196,N_9866,N_9664);
nand UO_197 (O_197,N_9596,N_9791);
nand UO_198 (O_198,N_9578,N_9770);
or UO_199 (O_199,N_9967,N_9850);
and UO_200 (O_200,N_9825,N_9916);
and UO_201 (O_201,N_9977,N_9992);
nand UO_202 (O_202,N_9604,N_9911);
nor UO_203 (O_203,N_9946,N_9784);
and UO_204 (O_204,N_9802,N_9970);
nor UO_205 (O_205,N_9549,N_9971);
nor UO_206 (O_206,N_9599,N_9803);
nor UO_207 (O_207,N_9783,N_9561);
or UO_208 (O_208,N_9863,N_9688);
nor UO_209 (O_209,N_9621,N_9703);
nand UO_210 (O_210,N_9723,N_9585);
nor UO_211 (O_211,N_9969,N_9830);
nor UO_212 (O_212,N_9872,N_9760);
and UO_213 (O_213,N_9598,N_9915);
nor UO_214 (O_214,N_9966,N_9529);
or UO_215 (O_215,N_9737,N_9669);
xnor UO_216 (O_216,N_9683,N_9717);
nand UO_217 (O_217,N_9538,N_9905);
nand UO_218 (O_218,N_9950,N_9557);
nor UO_219 (O_219,N_9519,N_9739);
and UO_220 (O_220,N_9887,N_9732);
nor UO_221 (O_221,N_9855,N_9899);
nor UO_222 (O_222,N_9835,N_9742);
nor UO_223 (O_223,N_9776,N_9626);
and UO_224 (O_224,N_9577,N_9890);
and UO_225 (O_225,N_9559,N_9807);
nor UO_226 (O_226,N_9678,N_9666);
and UO_227 (O_227,N_9505,N_9663);
and UO_228 (O_228,N_9811,N_9996);
nand UO_229 (O_229,N_9691,N_9973);
and UO_230 (O_230,N_9785,N_9930);
nor UO_231 (O_231,N_9533,N_9913);
nor UO_232 (O_232,N_9882,N_9702);
and UO_233 (O_233,N_9694,N_9602);
or UO_234 (O_234,N_9953,N_9753);
nor UO_235 (O_235,N_9610,N_9963);
or UO_236 (O_236,N_9993,N_9729);
nor UO_237 (O_237,N_9853,N_9636);
nor UO_238 (O_238,N_9671,N_9735);
or UO_239 (O_239,N_9840,N_9668);
nand UO_240 (O_240,N_9589,N_9781);
or UO_241 (O_241,N_9761,N_9954);
nor UO_242 (O_242,N_9534,N_9968);
or UO_243 (O_243,N_9607,N_9665);
and UO_244 (O_244,N_9767,N_9796);
nand UO_245 (O_245,N_9601,N_9896);
nand UO_246 (O_246,N_9788,N_9532);
or UO_247 (O_247,N_9537,N_9906);
nand UO_248 (O_248,N_9972,N_9562);
and UO_249 (O_249,N_9891,N_9541);
nor UO_250 (O_250,N_9640,N_9745);
or UO_251 (O_251,N_9672,N_9626);
nand UO_252 (O_252,N_9733,N_9643);
nor UO_253 (O_253,N_9507,N_9813);
nand UO_254 (O_254,N_9705,N_9776);
nor UO_255 (O_255,N_9731,N_9900);
or UO_256 (O_256,N_9595,N_9889);
and UO_257 (O_257,N_9968,N_9951);
nor UO_258 (O_258,N_9718,N_9642);
or UO_259 (O_259,N_9835,N_9893);
nor UO_260 (O_260,N_9920,N_9540);
or UO_261 (O_261,N_9877,N_9908);
and UO_262 (O_262,N_9664,N_9783);
nor UO_263 (O_263,N_9990,N_9885);
or UO_264 (O_264,N_9643,N_9750);
nor UO_265 (O_265,N_9610,N_9942);
and UO_266 (O_266,N_9708,N_9721);
and UO_267 (O_267,N_9538,N_9958);
and UO_268 (O_268,N_9558,N_9972);
nor UO_269 (O_269,N_9953,N_9980);
nand UO_270 (O_270,N_9912,N_9589);
nand UO_271 (O_271,N_9554,N_9731);
or UO_272 (O_272,N_9572,N_9751);
or UO_273 (O_273,N_9511,N_9627);
or UO_274 (O_274,N_9773,N_9986);
and UO_275 (O_275,N_9589,N_9694);
or UO_276 (O_276,N_9530,N_9781);
and UO_277 (O_277,N_9635,N_9649);
xor UO_278 (O_278,N_9591,N_9798);
and UO_279 (O_279,N_9739,N_9530);
nand UO_280 (O_280,N_9568,N_9941);
nor UO_281 (O_281,N_9663,N_9530);
and UO_282 (O_282,N_9689,N_9858);
or UO_283 (O_283,N_9938,N_9538);
and UO_284 (O_284,N_9607,N_9572);
or UO_285 (O_285,N_9633,N_9696);
or UO_286 (O_286,N_9753,N_9657);
nor UO_287 (O_287,N_9708,N_9563);
and UO_288 (O_288,N_9515,N_9686);
and UO_289 (O_289,N_9873,N_9704);
and UO_290 (O_290,N_9586,N_9904);
nor UO_291 (O_291,N_9961,N_9618);
or UO_292 (O_292,N_9714,N_9726);
or UO_293 (O_293,N_9977,N_9966);
and UO_294 (O_294,N_9958,N_9509);
nand UO_295 (O_295,N_9925,N_9566);
and UO_296 (O_296,N_9998,N_9992);
nor UO_297 (O_297,N_9739,N_9915);
nand UO_298 (O_298,N_9965,N_9731);
or UO_299 (O_299,N_9695,N_9744);
nor UO_300 (O_300,N_9517,N_9586);
nor UO_301 (O_301,N_9973,N_9767);
or UO_302 (O_302,N_9976,N_9881);
nand UO_303 (O_303,N_9587,N_9892);
or UO_304 (O_304,N_9993,N_9857);
or UO_305 (O_305,N_9881,N_9622);
nand UO_306 (O_306,N_9999,N_9729);
and UO_307 (O_307,N_9852,N_9956);
nand UO_308 (O_308,N_9999,N_9833);
and UO_309 (O_309,N_9727,N_9757);
nand UO_310 (O_310,N_9594,N_9813);
nor UO_311 (O_311,N_9818,N_9519);
nor UO_312 (O_312,N_9994,N_9922);
and UO_313 (O_313,N_9653,N_9647);
nor UO_314 (O_314,N_9774,N_9939);
nor UO_315 (O_315,N_9720,N_9673);
and UO_316 (O_316,N_9591,N_9736);
and UO_317 (O_317,N_9984,N_9788);
nor UO_318 (O_318,N_9551,N_9655);
and UO_319 (O_319,N_9544,N_9908);
or UO_320 (O_320,N_9598,N_9726);
nand UO_321 (O_321,N_9531,N_9755);
nor UO_322 (O_322,N_9900,N_9788);
or UO_323 (O_323,N_9872,N_9818);
and UO_324 (O_324,N_9816,N_9690);
nand UO_325 (O_325,N_9792,N_9899);
nor UO_326 (O_326,N_9802,N_9680);
and UO_327 (O_327,N_9711,N_9789);
nand UO_328 (O_328,N_9944,N_9613);
xnor UO_329 (O_329,N_9678,N_9849);
and UO_330 (O_330,N_9958,N_9790);
nand UO_331 (O_331,N_9764,N_9875);
or UO_332 (O_332,N_9546,N_9813);
or UO_333 (O_333,N_9910,N_9907);
or UO_334 (O_334,N_9782,N_9645);
and UO_335 (O_335,N_9754,N_9975);
or UO_336 (O_336,N_9685,N_9901);
or UO_337 (O_337,N_9710,N_9896);
and UO_338 (O_338,N_9515,N_9529);
or UO_339 (O_339,N_9881,N_9725);
or UO_340 (O_340,N_9613,N_9577);
nand UO_341 (O_341,N_9953,N_9943);
nand UO_342 (O_342,N_9636,N_9577);
nor UO_343 (O_343,N_9998,N_9831);
and UO_344 (O_344,N_9563,N_9870);
or UO_345 (O_345,N_9727,N_9825);
or UO_346 (O_346,N_9603,N_9793);
nor UO_347 (O_347,N_9759,N_9869);
nor UO_348 (O_348,N_9654,N_9856);
or UO_349 (O_349,N_9731,N_9891);
nor UO_350 (O_350,N_9739,N_9612);
nand UO_351 (O_351,N_9569,N_9901);
nor UO_352 (O_352,N_9565,N_9935);
xor UO_353 (O_353,N_9759,N_9606);
nand UO_354 (O_354,N_9623,N_9888);
or UO_355 (O_355,N_9625,N_9867);
and UO_356 (O_356,N_9691,N_9536);
or UO_357 (O_357,N_9856,N_9604);
and UO_358 (O_358,N_9999,N_9519);
nand UO_359 (O_359,N_9962,N_9786);
and UO_360 (O_360,N_9979,N_9769);
or UO_361 (O_361,N_9906,N_9640);
or UO_362 (O_362,N_9631,N_9730);
nor UO_363 (O_363,N_9701,N_9577);
nand UO_364 (O_364,N_9599,N_9697);
nor UO_365 (O_365,N_9539,N_9526);
nor UO_366 (O_366,N_9576,N_9658);
nor UO_367 (O_367,N_9551,N_9634);
nor UO_368 (O_368,N_9616,N_9553);
and UO_369 (O_369,N_9700,N_9606);
and UO_370 (O_370,N_9565,N_9525);
and UO_371 (O_371,N_9670,N_9752);
or UO_372 (O_372,N_9872,N_9531);
nor UO_373 (O_373,N_9602,N_9662);
and UO_374 (O_374,N_9536,N_9582);
nor UO_375 (O_375,N_9882,N_9693);
or UO_376 (O_376,N_9620,N_9618);
and UO_377 (O_377,N_9725,N_9686);
and UO_378 (O_378,N_9793,N_9619);
or UO_379 (O_379,N_9927,N_9978);
or UO_380 (O_380,N_9766,N_9711);
or UO_381 (O_381,N_9902,N_9913);
and UO_382 (O_382,N_9703,N_9685);
nand UO_383 (O_383,N_9943,N_9690);
and UO_384 (O_384,N_9709,N_9626);
and UO_385 (O_385,N_9559,N_9769);
nor UO_386 (O_386,N_9820,N_9934);
or UO_387 (O_387,N_9508,N_9973);
or UO_388 (O_388,N_9963,N_9827);
and UO_389 (O_389,N_9978,N_9932);
and UO_390 (O_390,N_9865,N_9512);
or UO_391 (O_391,N_9605,N_9952);
nand UO_392 (O_392,N_9919,N_9693);
nor UO_393 (O_393,N_9501,N_9961);
or UO_394 (O_394,N_9878,N_9848);
and UO_395 (O_395,N_9858,N_9962);
nand UO_396 (O_396,N_9957,N_9985);
xnor UO_397 (O_397,N_9537,N_9931);
or UO_398 (O_398,N_9593,N_9813);
nand UO_399 (O_399,N_9739,N_9575);
and UO_400 (O_400,N_9509,N_9678);
or UO_401 (O_401,N_9597,N_9607);
or UO_402 (O_402,N_9973,N_9776);
nand UO_403 (O_403,N_9734,N_9745);
nand UO_404 (O_404,N_9845,N_9602);
nand UO_405 (O_405,N_9508,N_9596);
or UO_406 (O_406,N_9925,N_9609);
nand UO_407 (O_407,N_9868,N_9782);
nand UO_408 (O_408,N_9763,N_9742);
nand UO_409 (O_409,N_9918,N_9626);
nor UO_410 (O_410,N_9673,N_9899);
nand UO_411 (O_411,N_9867,N_9830);
or UO_412 (O_412,N_9871,N_9818);
or UO_413 (O_413,N_9714,N_9729);
nor UO_414 (O_414,N_9640,N_9648);
or UO_415 (O_415,N_9725,N_9527);
nand UO_416 (O_416,N_9988,N_9879);
and UO_417 (O_417,N_9519,N_9939);
nand UO_418 (O_418,N_9747,N_9951);
nor UO_419 (O_419,N_9637,N_9946);
nand UO_420 (O_420,N_9693,N_9679);
and UO_421 (O_421,N_9687,N_9980);
or UO_422 (O_422,N_9890,N_9893);
or UO_423 (O_423,N_9684,N_9599);
nor UO_424 (O_424,N_9602,N_9706);
nand UO_425 (O_425,N_9646,N_9849);
or UO_426 (O_426,N_9782,N_9834);
nand UO_427 (O_427,N_9536,N_9718);
or UO_428 (O_428,N_9642,N_9772);
nand UO_429 (O_429,N_9841,N_9598);
or UO_430 (O_430,N_9917,N_9690);
nor UO_431 (O_431,N_9870,N_9617);
nand UO_432 (O_432,N_9788,N_9637);
nand UO_433 (O_433,N_9944,N_9648);
nor UO_434 (O_434,N_9875,N_9820);
nor UO_435 (O_435,N_9562,N_9544);
or UO_436 (O_436,N_9660,N_9563);
or UO_437 (O_437,N_9755,N_9800);
or UO_438 (O_438,N_9581,N_9841);
nor UO_439 (O_439,N_9786,N_9934);
or UO_440 (O_440,N_9878,N_9822);
nor UO_441 (O_441,N_9917,N_9515);
nand UO_442 (O_442,N_9933,N_9905);
nor UO_443 (O_443,N_9556,N_9626);
nor UO_444 (O_444,N_9856,N_9630);
nand UO_445 (O_445,N_9508,N_9777);
or UO_446 (O_446,N_9537,N_9589);
nor UO_447 (O_447,N_9529,N_9740);
nor UO_448 (O_448,N_9665,N_9851);
and UO_449 (O_449,N_9998,N_9954);
nand UO_450 (O_450,N_9779,N_9708);
nand UO_451 (O_451,N_9524,N_9815);
nand UO_452 (O_452,N_9994,N_9864);
or UO_453 (O_453,N_9726,N_9515);
nand UO_454 (O_454,N_9802,N_9985);
xor UO_455 (O_455,N_9977,N_9687);
nand UO_456 (O_456,N_9507,N_9766);
nor UO_457 (O_457,N_9876,N_9898);
nor UO_458 (O_458,N_9796,N_9659);
and UO_459 (O_459,N_9955,N_9950);
or UO_460 (O_460,N_9800,N_9604);
nand UO_461 (O_461,N_9569,N_9929);
or UO_462 (O_462,N_9998,N_9625);
and UO_463 (O_463,N_9550,N_9839);
nand UO_464 (O_464,N_9854,N_9771);
and UO_465 (O_465,N_9572,N_9623);
nand UO_466 (O_466,N_9693,N_9891);
or UO_467 (O_467,N_9811,N_9679);
or UO_468 (O_468,N_9930,N_9560);
or UO_469 (O_469,N_9736,N_9756);
or UO_470 (O_470,N_9597,N_9605);
and UO_471 (O_471,N_9680,N_9535);
and UO_472 (O_472,N_9903,N_9956);
or UO_473 (O_473,N_9530,N_9960);
or UO_474 (O_474,N_9808,N_9667);
or UO_475 (O_475,N_9810,N_9889);
nor UO_476 (O_476,N_9914,N_9916);
nor UO_477 (O_477,N_9626,N_9899);
nor UO_478 (O_478,N_9976,N_9733);
nand UO_479 (O_479,N_9644,N_9684);
and UO_480 (O_480,N_9952,N_9771);
nor UO_481 (O_481,N_9983,N_9605);
and UO_482 (O_482,N_9611,N_9943);
or UO_483 (O_483,N_9877,N_9814);
and UO_484 (O_484,N_9629,N_9539);
nor UO_485 (O_485,N_9568,N_9887);
nor UO_486 (O_486,N_9668,N_9751);
nor UO_487 (O_487,N_9822,N_9663);
nand UO_488 (O_488,N_9548,N_9716);
nor UO_489 (O_489,N_9803,N_9926);
or UO_490 (O_490,N_9995,N_9942);
xnor UO_491 (O_491,N_9850,N_9707);
or UO_492 (O_492,N_9858,N_9901);
and UO_493 (O_493,N_9943,N_9683);
and UO_494 (O_494,N_9698,N_9580);
nor UO_495 (O_495,N_9512,N_9728);
and UO_496 (O_496,N_9691,N_9777);
xnor UO_497 (O_497,N_9848,N_9801);
and UO_498 (O_498,N_9955,N_9974);
nor UO_499 (O_499,N_9971,N_9662);
nand UO_500 (O_500,N_9936,N_9939);
nand UO_501 (O_501,N_9671,N_9722);
nand UO_502 (O_502,N_9966,N_9762);
and UO_503 (O_503,N_9732,N_9623);
nor UO_504 (O_504,N_9740,N_9550);
and UO_505 (O_505,N_9884,N_9873);
nand UO_506 (O_506,N_9582,N_9610);
nand UO_507 (O_507,N_9571,N_9835);
and UO_508 (O_508,N_9971,N_9754);
nand UO_509 (O_509,N_9770,N_9581);
nand UO_510 (O_510,N_9866,N_9989);
nor UO_511 (O_511,N_9971,N_9584);
nand UO_512 (O_512,N_9749,N_9887);
and UO_513 (O_513,N_9606,N_9910);
nor UO_514 (O_514,N_9960,N_9884);
nor UO_515 (O_515,N_9529,N_9545);
nand UO_516 (O_516,N_9904,N_9892);
or UO_517 (O_517,N_9895,N_9737);
and UO_518 (O_518,N_9844,N_9953);
or UO_519 (O_519,N_9913,N_9963);
and UO_520 (O_520,N_9909,N_9768);
and UO_521 (O_521,N_9675,N_9748);
or UO_522 (O_522,N_9707,N_9998);
nand UO_523 (O_523,N_9870,N_9584);
nor UO_524 (O_524,N_9859,N_9967);
and UO_525 (O_525,N_9939,N_9947);
nand UO_526 (O_526,N_9657,N_9532);
nand UO_527 (O_527,N_9745,N_9740);
and UO_528 (O_528,N_9865,N_9919);
or UO_529 (O_529,N_9638,N_9540);
nand UO_530 (O_530,N_9980,N_9972);
or UO_531 (O_531,N_9513,N_9763);
nor UO_532 (O_532,N_9625,N_9618);
nand UO_533 (O_533,N_9664,N_9786);
or UO_534 (O_534,N_9786,N_9854);
nand UO_535 (O_535,N_9608,N_9996);
or UO_536 (O_536,N_9811,N_9672);
nor UO_537 (O_537,N_9501,N_9735);
nand UO_538 (O_538,N_9954,N_9801);
or UO_539 (O_539,N_9790,N_9672);
and UO_540 (O_540,N_9654,N_9631);
and UO_541 (O_541,N_9609,N_9836);
or UO_542 (O_542,N_9849,N_9584);
nand UO_543 (O_543,N_9823,N_9587);
nor UO_544 (O_544,N_9815,N_9946);
nand UO_545 (O_545,N_9800,N_9666);
nor UO_546 (O_546,N_9940,N_9636);
or UO_547 (O_547,N_9636,N_9730);
nor UO_548 (O_548,N_9796,N_9730);
or UO_549 (O_549,N_9962,N_9619);
and UO_550 (O_550,N_9644,N_9719);
nor UO_551 (O_551,N_9662,N_9964);
and UO_552 (O_552,N_9970,N_9902);
and UO_553 (O_553,N_9549,N_9568);
nand UO_554 (O_554,N_9896,N_9988);
and UO_555 (O_555,N_9562,N_9893);
and UO_556 (O_556,N_9530,N_9738);
and UO_557 (O_557,N_9620,N_9556);
and UO_558 (O_558,N_9806,N_9964);
nor UO_559 (O_559,N_9774,N_9602);
and UO_560 (O_560,N_9800,N_9891);
and UO_561 (O_561,N_9697,N_9944);
nand UO_562 (O_562,N_9916,N_9684);
and UO_563 (O_563,N_9996,N_9891);
and UO_564 (O_564,N_9545,N_9920);
nand UO_565 (O_565,N_9758,N_9547);
nor UO_566 (O_566,N_9635,N_9537);
and UO_567 (O_567,N_9999,N_9551);
xor UO_568 (O_568,N_9656,N_9959);
or UO_569 (O_569,N_9890,N_9556);
nand UO_570 (O_570,N_9982,N_9877);
and UO_571 (O_571,N_9898,N_9600);
nor UO_572 (O_572,N_9770,N_9648);
and UO_573 (O_573,N_9627,N_9589);
nand UO_574 (O_574,N_9889,N_9839);
and UO_575 (O_575,N_9590,N_9802);
nor UO_576 (O_576,N_9857,N_9583);
and UO_577 (O_577,N_9957,N_9922);
nor UO_578 (O_578,N_9706,N_9548);
nor UO_579 (O_579,N_9507,N_9546);
nand UO_580 (O_580,N_9970,N_9851);
nand UO_581 (O_581,N_9544,N_9673);
and UO_582 (O_582,N_9968,N_9795);
and UO_583 (O_583,N_9611,N_9945);
nor UO_584 (O_584,N_9540,N_9780);
and UO_585 (O_585,N_9685,N_9526);
nor UO_586 (O_586,N_9722,N_9872);
nand UO_587 (O_587,N_9859,N_9881);
or UO_588 (O_588,N_9833,N_9733);
or UO_589 (O_589,N_9540,N_9575);
nand UO_590 (O_590,N_9867,N_9582);
and UO_591 (O_591,N_9739,N_9547);
nand UO_592 (O_592,N_9974,N_9603);
nor UO_593 (O_593,N_9540,N_9987);
or UO_594 (O_594,N_9609,N_9996);
nand UO_595 (O_595,N_9977,N_9849);
nor UO_596 (O_596,N_9534,N_9874);
nand UO_597 (O_597,N_9937,N_9934);
nand UO_598 (O_598,N_9774,N_9531);
and UO_599 (O_599,N_9811,N_9539);
nand UO_600 (O_600,N_9678,N_9788);
nand UO_601 (O_601,N_9834,N_9875);
nand UO_602 (O_602,N_9696,N_9932);
or UO_603 (O_603,N_9937,N_9723);
nand UO_604 (O_604,N_9862,N_9912);
nor UO_605 (O_605,N_9521,N_9870);
nand UO_606 (O_606,N_9787,N_9585);
nand UO_607 (O_607,N_9507,N_9967);
xor UO_608 (O_608,N_9654,N_9934);
and UO_609 (O_609,N_9538,N_9572);
or UO_610 (O_610,N_9954,N_9557);
and UO_611 (O_611,N_9794,N_9798);
or UO_612 (O_612,N_9602,N_9836);
nand UO_613 (O_613,N_9772,N_9817);
or UO_614 (O_614,N_9748,N_9640);
nor UO_615 (O_615,N_9823,N_9882);
nor UO_616 (O_616,N_9543,N_9646);
and UO_617 (O_617,N_9915,N_9620);
nand UO_618 (O_618,N_9618,N_9978);
nand UO_619 (O_619,N_9717,N_9757);
nand UO_620 (O_620,N_9597,N_9806);
or UO_621 (O_621,N_9516,N_9557);
and UO_622 (O_622,N_9853,N_9642);
nand UO_623 (O_623,N_9750,N_9867);
nand UO_624 (O_624,N_9829,N_9677);
nor UO_625 (O_625,N_9575,N_9729);
and UO_626 (O_626,N_9542,N_9818);
and UO_627 (O_627,N_9513,N_9779);
or UO_628 (O_628,N_9742,N_9883);
nand UO_629 (O_629,N_9676,N_9787);
and UO_630 (O_630,N_9913,N_9614);
and UO_631 (O_631,N_9687,N_9748);
nand UO_632 (O_632,N_9847,N_9725);
nand UO_633 (O_633,N_9737,N_9641);
nand UO_634 (O_634,N_9755,N_9996);
xor UO_635 (O_635,N_9853,N_9962);
and UO_636 (O_636,N_9817,N_9504);
and UO_637 (O_637,N_9813,N_9859);
or UO_638 (O_638,N_9789,N_9955);
nor UO_639 (O_639,N_9892,N_9865);
or UO_640 (O_640,N_9615,N_9987);
and UO_641 (O_641,N_9793,N_9577);
nor UO_642 (O_642,N_9509,N_9596);
nor UO_643 (O_643,N_9896,N_9913);
or UO_644 (O_644,N_9771,N_9973);
or UO_645 (O_645,N_9977,N_9733);
nor UO_646 (O_646,N_9830,N_9533);
or UO_647 (O_647,N_9773,N_9718);
and UO_648 (O_648,N_9652,N_9560);
nand UO_649 (O_649,N_9923,N_9749);
nand UO_650 (O_650,N_9692,N_9639);
nor UO_651 (O_651,N_9554,N_9601);
nand UO_652 (O_652,N_9928,N_9700);
nor UO_653 (O_653,N_9615,N_9740);
nand UO_654 (O_654,N_9970,N_9652);
nand UO_655 (O_655,N_9948,N_9967);
or UO_656 (O_656,N_9788,N_9849);
and UO_657 (O_657,N_9673,N_9835);
nor UO_658 (O_658,N_9679,N_9933);
nor UO_659 (O_659,N_9632,N_9633);
and UO_660 (O_660,N_9638,N_9853);
nand UO_661 (O_661,N_9982,N_9974);
and UO_662 (O_662,N_9883,N_9758);
nand UO_663 (O_663,N_9509,N_9983);
and UO_664 (O_664,N_9777,N_9901);
or UO_665 (O_665,N_9724,N_9591);
and UO_666 (O_666,N_9885,N_9880);
nor UO_667 (O_667,N_9567,N_9571);
or UO_668 (O_668,N_9532,N_9650);
or UO_669 (O_669,N_9516,N_9940);
nor UO_670 (O_670,N_9726,N_9674);
nand UO_671 (O_671,N_9819,N_9880);
nor UO_672 (O_672,N_9650,N_9559);
nand UO_673 (O_673,N_9787,N_9785);
or UO_674 (O_674,N_9513,N_9575);
or UO_675 (O_675,N_9654,N_9884);
and UO_676 (O_676,N_9811,N_9662);
or UO_677 (O_677,N_9751,N_9603);
and UO_678 (O_678,N_9769,N_9682);
and UO_679 (O_679,N_9620,N_9591);
nor UO_680 (O_680,N_9745,N_9604);
nor UO_681 (O_681,N_9720,N_9836);
and UO_682 (O_682,N_9838,N_9869);
nand UO_683 (O_683,N_9929,N_9671);
nand UO_684 (O_684,N_9752,N_9730);
nor UO_685 (O_685,N_9761,N_9891);
and UO_686 (O_686,N_9805,N_9534);
nor UO_687 (O_687,N_9572,N_9677);
nor UO_688 (O_688,N_9990,N_9652);
xor UO_689 (O_689,N_9936,N_9752);
nand UO_690 (O_690,N_9678,N_9689);
nand UO_691 (O_691,N_9865,N_9953);
and UO_692 (O_692,N_9772,N_9806);
nand UO_693 (O_693,N_9845,N_9597);
nor UO_694 (O_694,N_9951,N_9799);
nand UO_695 (O_695,N_9663,N_9781);
or UO_696 (O_696,N_9718,N_9616);
nor UO_697 (O_697,N_9522,N_9575);
nand UO_698 (O_698,N_9789,N_9614);
and UO_699 (O_699,N_9716,N_9595);
or UO_700 (O_700,N_9501,N_9715);
xnor UO_701 (O_701,N_9540,N_9985);
nand UO_702 (O_702,N_9967,N_9511);
nor UO_703 (O_703,N_9978,N_9993);
nor UO_704 (O_704,N_9635,N_9654);
nor UO_705 (O_705,N_9503,N_9830);
and UO_706 (O_706,N_9701,N_9581);
or UO_707 (O_707,N_9625,N_9623);
nor UO_708 (O_708,N_9730,N_9995);
or UO_709 (O_709,N_9667,N_9854);
and UO_710 (O_710,N_9681,N_9831);
nor UO_711 (O_711,N_9551,N_9878);
or UO_712 (O_712,N_9870,N_9565);
nand UO_713 (O_713,N_9679,N_9986);
nand UO_714 (O_714,N_9559,N_9982);
nand UO_715 (O_715,N_9515,N_9612);
nand UO_716 (O_716,N_9705,N_9524);
and UO_717 (O_717,N_9630,N_9987);
nor UO_718 (O_718,N_9906,N_9524);
nor UO_719 (O_719,N_9984,N_9851);
and UO_720 (O_720,N_9926,N_9882);
and UO_721 (O_721,N_9614,N_9944);
or UO_722 (O_722,N_9815,N_9713);
or UO_723 (O_723,N_9890,N_9772);
and UO_724 (O_724,N_9856,N_9859);
and UO_725 (O_725,N_9508,N_9604);
or UO_726 (O_726,N_9946,N_9525);
nand UO_727 (O_727,N_9550,N_9636);
nand UO_728 (O_728,N_9962,N_9633);
nand UO_729 (O_729,N_9634,N_9538);
or UO_730 (O_730,N_9782,N_9758);
nand UO_731 (O_731,N_9600,N_9583);
and UO_732 (O_732,N_9530,N_9902);
nor UO_733 (O_733,N_9709,N_9545);
or UO_734 (O_734,N_9950,N_9765);
and UO_735 (O_735,N_9770,N_9607);
and UO_736 (O_736,N_9822,N_9910);
nor UO_737 (O_737,N_9626,N_9545);
and UO_738 (O_738,N_9866,N_9717);
xnor UO_739 (O_739,N_9625,N_9843);
nand UO_740 (O_740,N_9848,N_9514);
nor UO_741 (O_741,N_9697,N_9865);
xnor UO_742 (O_742,N_9908,N_9619);
nor UO_743 (O_743,N_9547,N_9619);
and UO_744 (O_744,N_9581,N_9585);
and UO_745 (O_745,N_9839,N_9794);
nand UO_746 (O_746,N_9549,N_9694);
nand UO_747 (O_747,N_9666,N_9951);
or UO_748 (O_748,N_9788,N_9761);
nor UO_749 (O_749,N_9920,N_9744);
or UO_750 (O_750,N_9532,N_9851);
nand UO_751 (O_751,N_9551,N_9602);
nor UO_752 (O_752,N_9536,N_9717);
or UO_753 (O_753,N_9827,N_9797);
nor UO_754 (O_754,N_9813,N_9523);
or UO_755 (O_755,N_9535,N_9911);
nand UO_756 (O_756,N_9741,N_9659);
nand UO_757 (O_757,N_9577,N_9814);
and UO_758 (O_758,N_9951,N_9636);
and UO_759 (O_759,N_9674,N_9841);
and UO_760 (O_760,N_9573,N_9986);
nor UO_761 (O_761,N_9817,N_9577);
and UO_762 (O_762,N_9546,N_9592);
nor UO_763 (O_763,N_9600,N_9602);
or UO_764 (O_764,N_9961,N_9802);
nor UO_765 (O_765,N_9660,N_9852);
and UO_766 (O_766,N_9850,N_9734);
nor UO_767 (O_767,N_9592,N_9551);
and UO_768 (O_768,N_9786,N_9568);
and UO_769 (O_769,N_9968,N_9917);
and UO_770 (O_770,N_9806,N_9750);
nor UO_771 (O_771,N_9963,N_9743);
and UO_772 (O_772,N_9938,N_9508);
and UO_773 (O_773,N_9928,N_9797);
nand UO_774 (O_774,N_9507,N_9748);
or UO_775 (O_775,N_9634,N_9673);
nand UO_776 (O_776,N_9548,N_9524);
nand UO_777 (O_777,N_9533,N_9887);
nand UO_778 (O_778,N_9552,N_9814);
nand UO_779 (O_779,N_9886,N_9987);
nand UO_780 (O_780,N_9604,N_9723);
nand UO_781 (O_781,N_9902,N_9641);
and UO_782 (O_782,N_9907,N_9947);
and UO_783 (O_783,N_9865,N_9912);
or UO_784 (O_784,N_9959,N_9586);
and UO_785 (O_785,N_9856,N_9841);
or UO_786 (O_786,N_9891,N_9524);
or UO_787 (O_787,N_9628,N_9874);
or UO_788 (O_788,N_9517,N_9601);
nor UO_789 (O_789,N_9891,N_9758);
or UO_790 (O_790,N_9514,N_9809);
nor UO_791 (O_791,N_9665,N_9774);
nand UO_792 (O_792,N_9931,N_9612);
nor UO_793 (O_793,N_9795,N_9595);
nand UO_794 (O_794,N_9501,N_9608);
nand UO_795 (O_795,N_9743,N_9741);
and UO_796 (O_796,N_9607,N_9982);
and UO_797 (O_797,N_9541,N_9803);
nor UO_798 (O_798,N_9961,N_9786);
nand UO_799 (O_799,N_9943,N_9978);
nand UO_800 (O_800,N_9599,N_9911);
xnor UO_801 (O_801,N_9575,N_9911);
nor UO_802 (O_802,N_9533,N_9806);
and UO_803 (O_803,N_9694,N_9862);
and UO_804 (O_804,N_9960,N_9893);
nor UO_805 (O_805,N_9648,N_9661);
and UO_806 (O_806,N_9554,N_9736);
nand UO_807 (O_807,N_9895,N_9928);
and UO_808 (O_808,N_9877,N_9714);
and UO_809 (O_809,N_9560,N_9936);
or UO_810 (O_810,N_9975,N_9863);
and UO_811 (O_811,N_9512,N_9923);
nand UO_812 (O_812,N_9547,N_9986);
nor UO_813 (O_813,N_9762,N_9699);
nor UO_814 (O_814,N_9871,N_9905);
and UO_815 (O_815,N_9946,N_9719);
or UO_816 (O_816,N_9789,N_9551);
nor UO_817 (O_817,N_9869,N_9875);
or UO_818 (O_818,N_9641,N_9768);
or UO_819 (O_819,N_9551,N_9617);
and UO_820 (O_820,N_9681,N_9716);
and UO_821 (O_821,N_9954,N_9535);
nor UO_822 (O_822,N_9832,N_9931);
or UO_823 (O_823,N_9640,N_9717);
nand UO_824 (O_824,N_9624,N_9863);
or UO_825 (O_825,N_9832,N_9546);
and UO_826 (O_826,N_9876,N_9878);
xor UO_827 (O_827,N_9989,N_9712);
or UO_828 (O_828,N_9653,N_9517);
nor UO_829 (O_829,N_9572,N_9883);
or UO_830 (O_830,N_9839,N_9505);
nand UO_831 (O_831,N_9949,N_9639);
nor UO_832 (O_832,N_9889,N_9966);
or UO_833 (O_833,N_9853,N_9874);
nand UO_834 (O_834,N_9770,N_9673);
nand UO_835 (O_835,N_9575,N_9712);
and UO_836 (O_836,N_9620,N_9582);
and UO_837 (O_837,N_9546,N_9825);
nor UO_838 (O_838,N_9576,N_9692);
or UO_839 (O_839,N_9707,N_9551);
nand UO_840 (O_840,N_9536,N_9899);
nor UO_841 (O_841,N_9860,N_9792);
and UO_842 (O_842,N_9609,N_9863);
or UO_843 (O_843,N_9684,N_9520);
or UO_844 (O_844,N_9513,N_9927);
nand UO_845 (O_845,N_9952,N_9897);
nor UO_846 (O_846,N_9889,N_9678);
nor UO_847 (O_847,N_9647,N_9750);
or UO_848 (O_848,N_9814,N_9840);
nand UO_849 (O_849,N_9765,N_9974);
and UO_850 (O_850,N_9653,N_9592);
nor UO_851 (O_851,N_9710,N_9889);
or UO_852 (O_852,N_9664,N_9758);
nand UO_853 (O_853,N_9871,N_9834);
xor UO_854 (O_854,N_9565,N_9602);
or UO_855 (O_855,N_9779,N_9536);
xnor UO_856 (O_856,N_9630,N_9910);
nor UO_857 (O_857,N_9780,N_9960);
nand UO_858 (O_858,N_9838,N_9923);
nand UO_859 (O_859,N_9888,N_9684);
or UO_860 (O_860,N_9550,N_9676);
or UO_861 (O_861,N_9794,N_9955);
or UO_862 (O_862,N_9564,N_9618);
or UO_863 (O_863,N_9858,N_9805);
or UO_864 (O_864,N_9990,N_9594);
or UO_865 (O_865,N_9621,N_9997);
and UO_866 (O_866,N_9565,N_9661);
nor UO_867 (O_867,N_9994,N_9911);
nor UO_868 (O_868,N_9775,N_9584);
nor UO_869 (O_869,N_9653,N_9587);
and UO_870 (O_870,N_9819,N_9969);
nor UO_871 (O_871,N_9638,N_9598);
or UO_872 (O_872,N_9935,N_9678);
nand UO_873 (O_873,N_9761,N_9547);
and UO_874 (O_874,N_9597,N_9506);
nand UO_875 (O_875,N_9580,N_9516);
nand UO_876 (O_876,N_9517,N_9788);
and UO_877 (O_877,N_9602,N_9539);
or UO_878 (O_878,N_9967,N_9510);
nand UO_879 (O_879,N_9790,N_9526);
and UO_880 (O_880,N_9647,N_9545);
nand UO_881 (O_881,N_9951,N_9632);
nand UO_882 (O_882,N_9866,N_9776);
nand UO_883 (O_883,N_9929,N_9861);
or UO_884 (O_884,N_9825,N_9809);
nor UO_885 (O_885,N_9584,N_9751);
nor UO_886 (O_886,N_9719,N_9816);
nand UO_887 (O_887,N_9894,N_9606);
nor UO_888 (O_888,N_9696,N_9837);
nor UO_889 (O_889,N_9901,N_9637);
nor UO_890 (O_890,N_9520,N_9903);
or UO_891 (O_891,N_9865,N_9544);
nor UO_892 (O_892,N_9998,N_9848);
and UO_893 (O_893,N_9844,N_9881);
nand UO_894 (O_894,N_9757,N_9808);
or UO_895 (O_895,N_9920,N_9846);
nor UO_896 (O_896,N_9813,N_9954);
or UO_897 (O_897,N_9701,N_9754);
nand UO_898 (O_898,N_9675,N_9690);
nand UO_899 (O_899,N_9705,N_9951);
nor UO_900 (O_900,N_9823,N_9532);
and UO_901 (O_901,N_9545,N_9640);
xnor UO_902 (O_902,N_9615,N_9878);
xor UO_903 (O_903,N_9644,N_9619);
nand UO_904 (O_904,N_9582,N_9785);
or UO_905 (O_905,N_9583,N_9848);
nand UO_906 (O_906,N_9726,N_9524);
and UO_907 (O_907,N_9959,N_9939);
or UO_908 (O_908,N_9820,N_9710);
or UO_909 (O_909,N_9745,N_9694);
and UO_910 (O_910,N_9799,N_9913);
or UO_911 (O_911,N_9762,N_9779);
or UO_912 (O_912,N_9843,N_9821);
nand UO_913 (O_913,N_9954,N_9540);
and UO_914 (O_914,N_9944,N_9533);
nand UO_915 (O_915,N_9968,N_9807);
nor UO_916 (O_916,N_9618,N_9697);
or UO_917 (O_917,N_9691,N_9692);
and UO_918 (O_918,N_9652,N_9758);
nor UO_919 (O_919,N_9700,N_9990);
and UO_920 (O_920,N_9534,N_9902);
or UO_921 (O_921,N_9510,N_9942);
or UO_922 (O_922,N_9527,N_9786);
nand UO_923 (O_923,N_9580,N_9907);
nor UO_924 (O_924,N_9889,N_9814);
and UO_925 (O_925,N_9632,N_9933);
nand UO_926 (O_926,N_9781,N_9656);
nor UO_927 (O_927,N_9742,N_9950);
or UO_928 (O_928,N_9539,N_9618);
or UO_929 (O_929,N_9990,N_9507);
and UO_930 (O_930,N_9665,N_9937);
and UO_931 (O_931,N_9718,N_9639);
nor UO_932 (O_932,N_9795,N_9649);
and UO_933 (O_933,N_9862,N_9774);
nand UO_934 (O_934,N_9921,N_9635);
and UO_935 (O_935,N_9740,N_9781);
or UO_936 (O_936,N_9930,N_9914);
or UO_937 (O_937,N_9595,N_9823);
nor UO_938 (O_938,N_9785,N_9736);
or UO_939 (O_939,N_9787,N_9893);
nand UO_940 (O_940,N_9693,N_9544);
nor UO_941 (O_941,N_9838,N_9611);
or UO_942 (O_942,N_9651,N_9949);
and UO_943 (O_943,N_9778,N_9961);
nor UO_944 (O_944,N_9952,N_9566);
or UO_945 (O_945,N_9720,N_9795);
and UO_946 (O_946,N_9960,N_9636);
nand UO_947 (O_947,N_9511,N_9617);
and UO_948 (O_948,N_9515,N_9913);
or UO_949 (O_949,N_9819,N_9889);
nand UO_950 (O_950,N_9525,N_9860);
xnor UO_951 (O_951,N_9638,N_9707);
nor UO_952 (O_952,N_9997,N_9814);
and UO_953 (O_953,N_9886,N_9613);
nor UO_954 (O_954,N_9930,N_9965);
nand UO_955 (O_955,N_9727,N_9858);
or UO_956 (O_956,N_9844,N_9540);
and UO_957 (O_957,N_9991,N_9756);
or UO_958 (O_958,N_9538,N_9994);
or UO_959 (O_959,N_9545,N_9757);
and UO_960 (O_960,N_9739,N_9923);
nand UO_961 (O_961,N_9546,N_9926);
nand UO_962 (O_962,N_9580,N_9735);
nor UO_963 (O_963,N_9628,N_9936);
nand UO_964 (O_964,N_9857,N_9982);
nor UO_965 (O_965,N_9966,N_9581);
and UO_966 (O_966,N_9916,N_9897);
nor UO_967 (O_967,N_9684,N_9562);
or UO_968 (O_968,N_9676,N_9724);
nor UO_969 (O_969,N_9936,N_9807);
and UO_970 (O_970,N_9846,N_9502);
nor UO_971 (O_971,N_9578,N_9807);
nor UO_972 (O_972,N_9564,N_9774);
nor UO_973 (O_973,N_9557,N_9838);
nand UO_974 (O_974,N_9589,N_9581);
nand UO_975 (O_975,N_9982,N_9629);
nand UO_976 (O_976,N_9735,N_9551);
xor UO_977 (O_977,N_9518,N_9809);
nand UO_978 (O_978,N_9651,N_9706);
nor UO_979 (O_979,N_9947,N_9856);
and UO_980 (O_980,N_9802,N_9633);
nand UO_981 (O_981,N_9895,N_9873);
and UO_982 (O_982,N_9899,N_9704);
nand UO_983 (O_983,N_9807,N_9924);
nor UO_984 (O_984,N_9851,N_9951);
and UO_985 (O_985,N_9604,N_9524);
nor UO_986 (O_986,N_9715,N_9726);
nor UO_987 (O_987,N_9507,N_9794);
and UO_988 (O_988,N_9539,N_9530);
nand UO_989 (O_989,N_9639,N_9928);
and UO_990 (O_990,N_9915,N_9923);
and UO_991 (O_991,N_9599,N_9618);
nor UO_992 (O_992,N_9604,N_9728);
nand UO_993 (O_993,N_9704,N_9664);
xnor UO_994 (O_994,N_9767,N_9864);
nand UO_995 (O_995,N_9913,N_9784);
nor UO_996 (O_996,N_9985,N_9722);
or UO_997 (O_997,N_9606,N_9979);
or UO_998 (O_998,N_9658,N_9870);
and UO_999 (O_999,N_9639,N_9615);
nand UO_1000 (O_1000,N_9660,N_9870);
nand UO_1001 (O_1001,N_9787,N_9576);
nand UO_1002 (O_1002,N_9575,N_9756);
nor UO_1003 (O_1003,N_9636,N_9828);
xor UO_1004 (O_1004,N_9833,N_9700);
nand UO_1005 (O_1005,N_9798,N_9515);
and UO_1006 (O_1006,N_9642,N_9579);
nand UO_1007 (O_1007,N_9840,N_9932);
nor UO_1008 (O_1008,N_9638,N_9606);
or UO_1009 (O_1009,N_9936,N_9713);
or UO_1010 (O_1010,N_9639,N_9590);
or UO_1011 (O_1011,N_9779,N_9781);
and UO_1012 (O_1012,N_9775,N_9934);
and UO_1013 (O_1013,N_9911,N_9989);
nor UO_1014 (O_1014,N_9737,N_9656);
nand UO_1015 (O_1015,N_9765,N_9753);
nor UO_1016 (O_1016,N_9603,N_9743);
nor UO_1017 (O_1017,N_9502,N_9563);
and UO_1018 (O_1018,N_9773,N_9905);
nor UO_1019 (O_1019,N_9781,N_9771);
and UO_1020 (O_1020,N_9891,N_9985);
nand UO_1021 (O_1021,N_9579,N_9944);
nor UO_1022 (O_1022,N_9982,N_9914);
nor UO_1023 (O_1023,N_9692,N_9888);
nor UO_1024 (O_1024,N_9517,N_9832);
or UO_1025 (O_1025,N_9640,N_9953);
nand UO_1026 (O_1026,N_9685,N_9965);
or UO_1027 (O_1027,N_9703,N_9986);
or UO_1028 (O_1028,N_9875,N_9591);
xnor UO_1029 (O_1029,N_9949,N_9796);
and UO_1030 (O_1030,N_9656,N_9513);
or UO_1031 (O_1031,N_9924,N_9547);
nor UO_1032 (O_1032,N_9646,N_9884);
or UO_1033 (O_1033,N_9955,N_9695);
or UO_1034 (O_1034,N_9573,N_9847);
or UO_1035 (O_1035,N_9856,N_9589);
nor UO_1036 (O_1036,N_9764,N_9767);
nor UO_1037 (O_1037,N_9867,N_9592);
and UO_1038 (O_1038,N_9617,N_9855);
or UO_1039 (O_1039,N_9537,N_9774);
and UO_1040 (O_1040,N_9627,N_9847);
nand UO_1041 (O_1041,N_9977,N_9757);
nor UO_1042 (O_1042,N_9844,N_9565);
nor UO_1043 (O_1043,N_9985,N_9948);
nand UO_1044 (O_1044,N_9651,N_9951);
nor UO_1045 (O_1045,N_9525,N_9737);
nor UO_1046 (O_1046,N_9721,N_9784);
and UO_1047 (O_1047,N_9754,N_9721);
and UO_1048 (O_1048,N_9671,N_9538);
nand UO_1049 (O_1049,N_9576,N_9763);
nor UO_1050 (O_1050,N_9594,N_9822);
and UO_1051 (O_1051,N_9630,N_9700);
nand UO_1052 (O_1052,N_9549,N_9731);
nor UO_1053 (O_1053,N_9650,N_9593);
and UO_1054 (O_1054,N_9960,N_9662);
and UO_1055 (O_1055,N_9733,N_9846);
nor UO_1056 (O_1056,N_9533,N_9921);
nor UO_1057 (O_1057,N_9870,N_9737);
and UO_1058 (O_1058,N_9699,N_9852);
or UO_1059 (O_1059,N_9902,N_9515);
and UO_1060 (O_1060,N_9997,N_9958);
nand UO_1061 (O_1061,N_9920,N_9934);
and UO_1062 (O_1062,N_9801,N_9740);
or UO_1063 (O_1063,N_9557,N_9896);
nor UO_1064 (O_1064,N_9983,N_9906);
or UO_1065 (O_1065,N_9785,N_9812);
nand UO_1066 (O_1066,N_9768,N_9978);
or UO_1067 (O_1067,N_9915,N_9639);
and UO_1068 (O_1068,N_9702,N_9519);
nand UO_1069 (O_1069,N_9516,N_9570);
nand UO_1070 (O_1070,N_9963,N_9869);
and UO_1071 (O_1071,N_9709,N_9894);
nor UO_1072 (O_1072,N_9664,N_9991);
nand UO_1073 (O_1073,N_9597,N_9939);
and UO_1074 (O_1074,N_9895,N_9863);
nand UO_1075 (O_1075,N_9762,N_9757);
or UO_1076 (O_1076,N_9693,N_9707);
nor UO_1077 (O_1077,N_9605,N_9950);
or UO_1078 (O_1078,N_9685,N_9618);
nor UO_1079 (O_1079,N_9831,N_9982);
nand UO_1080 (O_1080,N_9685,N_9591);
or UO_1081 (O_1081,N_9768,N_9635);
xnor UO_1082 (O_1082,N_9810,N_9669);
xor UO_1083 (O_1083,N_9956,N_9541);
nand UO_1084 (O_1084,N_9615,N_9848);
and UO_1085 (O_1085,N_9653,N_9612);
xnor UO_1086 (O_1086,N_9645,N_9905);
or UO_1087 (O_1087,N_9511,N_9891);
and UO_1088 (O_1088,N_9948,N_9817);
nand UO_1089 (O_1089,N_9823,N_9772);
or UO_1090 (O_1090,N_9630,N_9646);
nand UO_1091 (O_1091,N_9662,N_9947);
and UO_1092 (O_1092,N_9726,N_9629);
nand UO_1093 (O_1093,N_9601,N_9634);
nor UO_1094 (O_1094,N_9901,N_9802);
nand UO_1095 (O_1095,N_9713,N_9633);
or UO_1096 (O_1096,N_9814,N_9534);
nor UO_1097 (O_1097,N_9910,N_9781);
nand UO_1098 (O_1098,N_9571,N_9531);
or UO_1099 (O_1099,N_9918,N_9880);
nand UO_1100 (O_1100,N_9694,N_9934);
or UO_1101 (O_1101,N_9698,N_9987);
or UO_1102 (O_1102,N_9665,N_9820);
or UO_1103 (O_1103,N_9571,N_9715);
or UO_1104 (O_1104,N_9939,N_9719);
and UO_1105 (O_1105,N_9668,N_9661);
or UO_1106 (O_1106,N_9727,N_9874);
or UO_1107 (O_1107,N_9948,N_9944);
and UO_1108 (O_1108,N_9699,N_9905);
nand UO_1109 (O_1109,N_9527,N_9878);
or UO_1110 (O_1110,N_9570,N_9645);
nor UO_1111 (O_1111,N_9876,N_9705);
nand UO_1112 (O_1112,N_9570,N_9934);
nand UO_1113 (O_1113,N_9752,N_9627);
nor UO_1114 (O_1114,N_9828,N_9548);
nor UO_1115 (O_1115,N_9752,N_9774);
nor UO_1116 (O_1116,N_9729,N_9922);
and UO_1117 (O_1117,N_9790,N_9665);
nand UO_1118 (O_1118,N_9937,N_9751);
nand UO_1119 (O_1119,N_9792,N_9980);
and UO_1120 (O_1120,N_9676,N_9814);
or UO_1121 (O_1121,N_9695,N_9992);
and UO_1122 (O_1122,N_9624,N_9694);
nand UO_1123 (O_1123,N_9563,N_9612);
and UO_1124 (O_1124,N_9682,N_9948);
or UO_1125 (O_1125,N_9512,N_9631);
nand UO_1126 (O_1126,N_9674,N_9830);
or UO_1127 (O_1127,N_9501,N_9592);
and UO_1128 (O_1128,N_9981,N_9966);
xnor UO_1129 (O_1129,N_9639,N_9973);
or UO_1130 (O_1130,N_9798,N_9639);
nand UO_1131 (O_1131,N_9660,N_9580);
nand UO_1132 (O_1132,N_9862,N_9582);
nand UO_1133 (O_1133,N_9656,N_9733);
nor UO_1134 (O_1134,N_9723,N_9606);
nor UO_1135 (O_1135,N_9692,N_9512);
nand UO_1136 (O_1136,N_9846,N_9847);
or UO_1137 (O_1137,N_9825,N_9667);
and UO_1138 (O_1138,N_9940,N_9534);
and UO_1139 (O_1139,N_9882,N_9517);
nand UO_1140 (O_1140,N_9866,N_9526);
and UO_1141 (O_1141,N_9801,N_9525);
nand UO_1142 (O_1142,N_9603,N_9901);
xor UO_1143 (O_1143,N_9710,N_9880);
nand UO_1144 (O_1144,N_9861,N_9619);
nand UO_1145 (O_1145,N_9969,N_9923);
or UO_1146 (O_1146,N_9926,N_9945);
or UO_1147 (O_1147,N_9761,N_9929);
nand UO_1148 (O_1148,N_9805,N_9573);
and UO_1149 (O_1149,N_9533,N_9797);
nand UO_1150 (O_1150,N_9791,N_9608);
nor UO_1151 (O_1151,N_9754,N_9875);
nand UO_1152 (O_1152,N_9905,N_9660);
nand UO_1153 (O_1153,N_9781,N_9727);
or UO_1154 (O_1154,N_9745,N_9951);
nand UO_1155 (O_1155,N_9596,N_9734);
and UO_1156 (O_1156,N_9987,N_9772);
nor UO_1157 (O_1157,N_9958,N_9753);
or UO_1158 (O_1158,N_9799,N_9631);
and UO_1159 (O_1159,N_9963,N_9890);
xor UO_1160 (O_1160,N_9738,N_9856);
or UO_1161 (O_1161,N_9852,N_9809);
and UO_1162 (O_1162,N_9682,N_9626);
and UO_1163 (O_1163,N_9735,N_9887);
and UO_1164 (O_1164,N_9594,N_9681);
and UO_1165 (O_1165,N_9911,N_9934);
and UO_1166 (O_1166,N_9988,N_9849);
nor UO_1167 (O_1167,N_9631,N_9513);
nand UO_1168 (O_1168,N_9978,N_9983);
and UO_1169 (O_1169,N_9581,N_9835);
or UO_1170 (O_1170,N_9706,N_9525);
and UO_1171 (O_1171,N_9898,N_9690);
nor UO_1172 (O_1172,N_9893,N_9679);
nor UO_1173 (O_1173,N_9728,N_9713);
nor UO_1174 (O_1174,N_9537,N_9636);
or UO_1175 (O_1175,N_9671,N_9694);
nand UO_1176 (O_1176,N_9716,N_9728);
nand UO_1177 (O_1177,N_9683,N_9675);
nor UO_1178 (O_1178,N_9587,N_9707);
xor UO_1179 (O_1179,N_9586,N_9955);
and UO_1180 (O_1180,N_9737,N_9604);
or UO_1181 (O_1181,N_9906,N_9849);
and UO_1182 (O_1182,N_9700,N_9858);
nand UO_1183 (O_1183,N_9590,N_9773);
and UO_1184 (O_1184,N_9844,N_9840);
nand UO_1185 (O_1185,N_9891,N_9863);
xnor UO_1186 (O_1186,N_9725,N_9817);
and UO_1187 (O_1187,N_9837,N_9625);
nor UO_1188 (O_1188,N_9993,N_9515);
or UO_1189 (O_1189,N_9746,N_9661);
or UO_1190 (O_1190,N_9833,N_9703);
nor UO_1191 (O_1191,N_9619,N_9792);
nand UO_1192 (O_1192,N_9654,N_9562);
or UO_1193 (O_1193,N_9898,N_9830);
nor UO_1194 (O_1194,N_9631,N_9675);
or UO_1195 (O_1195,N_9552,N_9741);
or UO_1196 (O_1196,N_9594,N_9528);
nand UO_1197 (O_1197,N_9849,N_9699);
nor UO_1198 (O_1198,N_9755,N_9607);
and UO_1199 (O_1199,N_9891,N_9515);
and UO_1200 (O_1200,N_9901,N_9805);
nand UO_1201 (O_1201,N_9675,N_9760);
or UO_1202 (O_1202,N_9624,N_9838);
nor UO_1203 (O_1203,N_9693,N_9935);
nor UO_1204 (O_1204,N_9878,N_9558);
nor UO_1205 (O_1205,N_9849,N_9586);
nor UO_1206 (O_1206,N_9720,N_9538);
nand UO_1207 (O_1207,N_9769,N_9716);
nor UO_1208 (O_1208,N_9586,N_9837);
and UO_1209 (O_1209,N_9664,N_9714);
or UO_1210 (O_1210,N_9884,N_9909);
nand UO_1211 (O_1211,N_9665,N_9919);
or UO_1212 (O_1212,N_9684,N_9974);
nand UO_1213 (O_1213,N_9989,N_9555);
nand UO_1214 (O_1214,N_9887,N_9890);
or UO_1215 (O_1215,N_9921,N_9843);
or UO_1216 (O_1216,N_9607,N_9697);
nor UO_1217 (O_1217,N_9586,N_9892);
nand UO_1218 (O_1218,N_9571,N_9925);
or UO_1219 (O_1219,N_9616,N_9988);
and UO_1220 (O_1220,N_9820,N_9801);
and UO_1221 (O_1221,N_9955,N_9949);
and UO_1222 (O_1222,N_9684,N_9580);
and UO_1223 (O_1223,N_9920,N_9812);
or UO_1224 (O_1224,N_9794,N_9625);
nand UO_1225 (O_1225,N_9631,N_9648);
and UO_1226 (O_1226,N_9915,N_9772);
nor UO_1227 (O_1227,N_9661,N_9644);
or UO_1228 (O_1228,N_9729,N_9980);
nand UO_1229 (O_1229,N_9914,N_9787);
and UO_1230 (O_1230,N_9997,N_9803);
nor UO_1231 (O_1231,N_9975,N_9742);
nor UO_1232 (O_1232,N_9886,N_9825);
and UO_1233 (O_1233,N_9910,N_9775);
and UO_1234 (O_1234,N_9909,N_9517);
and UO_1235 (O_1235,N_9594,N_9878);
or UO_1236 (O_1236,N_9906,N_9635);
or UO_1237 (O_1237,N_9748,N_9933);
or UO_1238 (O_1238,N_9554,N_9655);
or UO_1239 (O_1239,N_9783,N_9661);
or UO_1240 (O_1240,N_9778,N_9871);
and UO_1241 (O_1241,N_9610,N_9554);
nand UO_1242 (O_1242,N_9911,N_9917);
nand UO_1243 (O_1243,N_9904,N_9721);
nor UO_1244 (O_1244,N_9905,N_9849);
nor UO_1245 (O_1245,N_9562,N_9660);
or UO_1246 (O_1246,N_9907,N_9799);
and UO_1247 (O_1247,N_9878,N_9635);
nand UO_1248 (O_1248,N_9708,N_9878);
or UO_1249 (O_1249,N_9832,N_9532);
nor UO_1250 (O_1250,N_9909,N_9928);
or UO_1251 (O_1251,N_9512,N_9880);
or UO_1252 (O_1252,N_9711,N_9818);
nand UO_1253 (O_1253,N_9976,N_9555);
xnor UO_1254 (O_1254,N_9686,N_9658);
nand UO_1255 (O_1255,N_9552,N_9970);
or UO_1256 (O_1256,N_9830,N_9924);
nand UO_1257 (O_1257,N_9607,N_9557);
or UO_1258 (O_1258,N_9567,N_9919);
and UO_1259 (O_1259,N_9782,N_9675);
and UO_1260 (O_1260,N_9557,N_9975);
and UO_1261 (O_1261,N_9867,N_9753);
nand UO_1262 (O_1262,N_9678,N_9708);
nand UO_1263 (O_1263,N_9569,N_9871);
nor UO_1264 (O_1264,N_9616,N_9786);
or UO_1265 (O_1265,N_9812,N_9501);
and UO_1266 (O_1266,N_9599,N_9839);
and UO_1267 (O_1267,N_9911,N_9736);
and UO_1268 (O_1268,N_9686,N_9826);
and UO_1269 (O_1269,N_9849,N_9735);
and UO_1270 (O_1270,N_9557,N_9732);
nor UO_1271 (O_1271,N_9963,N_9990);
nand UO_1272 (O_1272,N_9879,N_9668);
or UO_1273 (O_1273,N_9725,N_9762);
xnor UO_1274 (O_1274,N_9927,N_9980);
nand UO_1275 (O_1275,N_9766,N_9610);
and UO_1276 (O_1276,N_9528,N_9759);
nor UO_1277 (O_1277,N_9711,N_9997);
nor UO_1278 (O_1278,N_9893,N_9656);
and UO_1279 (O_1279,N_9894,N_9863);
xnor UO_1280 (O_1280,N_9500,N_9720);
xnor UO_1281 (O_1281,N_9797,N_9912);
and UO_1282 (O_1282,N_9692,N_9676);
nand UO_1283 (O_1283,N_9550,N_9693);
nor UO_1284 (O_1284,N_9516,N_9901);
or UO_1285 (O_1285,N_9679,N_9808);
nand UO_1286 (O_1286,N_9779,N_9850);
or UO_1287 (O_1287,N_9950,N_9500);
or UO_1288 (O_1288,N_9847,N_9669);
or UO_1289 (O_1289,N_9631,N_9968);
and UO_1290 (O_1290,N_9948,N_9827);
nand UO_1291 (O_1291,N_9999,N_9660);
and UO_1292 (O_1292,N_9836,N_9985);
and UO_1293 (O_1293,N_9663,N_9676);
and UO_1294 (O_1294,N_9567,N_9971);
nand UO_1295 (O_1295,N_9749,N_9980);
or UO_1296 (O_1296,N_9651,N_9809);
and UO_1297 (O_1297,N_9954,N_9724);
nand UO_1298 (O_1298,N_9977,N_9826);
and UO_1299 (O_1299,N_9947,N_9935);
nor UO_1300 (O_1300,N_9840,N_9804);
nand UO_1301 (O_1301,N_9613,N_9983);
nand UO_1302 (O_1302,N_9856,N_9673);
and UO_1303 (O_1303,N_9769,N_9724);
nor UO_1304 (O_1304,N_9661,N_9624);
nand UO_1305 (O_1305,N_9619,N_9991);
nand UO_1306 (O_1306,N_9736,N_9928);
nand UO_1307 (O_1307,N_9624,N_9710);
nor UO_1308 (O_1308,N_9591,N_9552);
or UO_1309 (O_1309,N_9594,N_9586);
nand UO_1310 (O_1310,N_9724,N_9672);
nand UO_1311 (O_1311,N_9886,N_9684);
and UO_1312 (O_1312,N_9507,N_9907);
or UO_1313 (O_1313,N_9991,N_9794);
xor UO_1314 (O_1314,N_9767,N_9830);
nor UO_1315 (O_1315,N_9816,N_9513);
and UO_1316 (O_1316,N_9801,N_9866);
or UO_1317 (O_1317,N_9985,N_9699);
nor UO_1318 (O_1318,N_9522,N_9997);
and UO_1319 (O_1319,N_9530,N_9875);
nor UO_1320 (O_1320,N_9696,N_9963);
nand UO_1321 (O_1321,N_9584,N_9571);
nor UO_1322 (O_1322,N_9921,N_9872);
and UO_1323 (O_1323,N_9865,N_9792);
and UO_1324 (O_1324,N_9518,N_9811);
and UO_1325 (O_1325,N_9901,N_9714);
xor UO_1326 (O_1326,N_9941,N_9699);
or UO_1327 (O_1327,N_9691,N_9981);
and UO_1328 (O_1328,N_9746,N_9893);
or UO_1329 (O_1329,N_9942,N_9952);
or UO_1330 (O_1330,N_9592,N_9728);
or UO_1331 (O_1331,N_9626,N_9529);
nand UO_1332 (O_1332,N_9701,N_9510);
nand UO_1333 (O_1333,N_9550,N_9664);
nor UO_1334 (O_1334,N_9861,N_9533);
or UO_1335 (O_1335,N_9904,N_9760);
or UO_1336 (O_1336,N_9532,N_9542);
or UO_1337 (O_1337,N_9720,N_9946);
or UO_1338 (O_1338,N_9891,N_9944);
or UO_1339 (O_1339,N_9790,N_9818);
nor UO_1340 (O_1340,N_9925,N_9980);
or UO_1341 (O_1341,N_9526,N_9501);
nand UO_1342 (O_1342,N_9639,N_9773);
and UO_1343 (O_1343,N_9591,N_9898);
and UO_1344 (O_1344,N_9552,N_9549);
and UO_1345 (O_1345,N_9952,N_9724);
nand UO_1346 (O_1346,N_9616,N_9955);
nor UO_1347 (O_1347,N_9991,N_9890);
or UO_1348 (O_1348,N_9510,N_9545);
or UO_1349 (O_1349,N_9744,N_9735);
or UO_1350 (O_1350,N_9949,N_9686);
xor UO_1351 (O_1351,N_9701,N_9555);
nand UO_1352 (O_1352,N_9548,N_9802);
nor UO_1353 (O_1353,N_9752,N_9619);
nand UO_1354 (O_1354,N_9575,N_9988);
nand UO_1355 (O_1355,N_9934,N_9649);
or UO_1356 (O_1356,N_9562,N_9969);
nand UO_1357 (O_1357,N_9876,N_9883);
nor UO_1358 (O_1358,N_9698,N_9812);
and UO_1359 (O_1359,N_9922,N_9945);
xnor UO_1360 (O_1360,N_9572,N_9562);
and UO_1361 (O_1361,N_9559,N_9529);
nor UO_1362 (O_1362,N_9556,N_9685);
nand UO_1363 (O_1363,N_9600,N_9882);
and UO_1364 (O_1364,N_9760,N_9523);
or UO_1365 (O_1365,N_9617,N_9976);
nor UO_1366 (O_1366,N_9916,N_9526);
and UO_1367 (O_1367,N_9932,N_9917);
nand UO_1368 (O_1368,N_9527,N_9607);
or UO_1369 (O_1369,N_9822,N_9846);
or UO_1370 (O_1370,N_9875,N_9566);
and UO_1371 (O_1371,N_9591,N_9892);
nor UO_1372 (O_1372,N_9579,N_9617);
nand UO_1373 (O_1373,N_9964,N_9951);
nor UO_1374 (O_1374,N_9641,N_9952);
and UO_1375 (O_1375,N_9645,N_9769);
or UO_1376 (O_1376,N_9705,N_9679);
or UO_1377 (O_1377,N_9780,N_9857);
or UO_1378 (O_1378,N_9692,N_9768);
nor UO_1379 (O_1379,N_9858,N_9766);
or UO_1380 (O_1380,N_9887,N_9617);
or UO_1381 (O_1381,N_9693,N_9593);
and UO_1382 (O_1382,N_9678,N_9723);
or UO_1383 (O_1383,N_9578,N_9862);
and UO_1384 (O_1384,N_9969,N_9551);
or UO_1385 (O_1385,N_9601,N_9890);
and UO_1386 (O_1386,N_9577,N_9552);
nor UO_1387 (O_1387,N_9966,N_9670);
nand UO_1388 (O_1388,N_9671,N_9618);
nor UO_1389 (O_1389,N_9916,N_9975);
nor UO_1390 (O_1390,N_9931,N_9764);
nand UO_1391 (O_1391,N_9858,N_9853);
nor UO_1392 (O_1392,N_9513,N_9599);
and UO_1393 (O_1393,N_9581,N_9752);
or UO_1394 (O_1394,N_9867,N_9998);
nand UO_1395 (O_1395,N_9502,N_9747);
nand UO_1396 (O_1396,N_9737,N_9740);
nor UO_1397 (O_1397,N_9596,N_9992);
or UO_1398 (O_1398,N_9704,N_9914);
and UO_1399 (O_1399,N_9985,N_9963);
and UO_1400 (O_1400,N_9635,N_9643);
and UO_1401 (O_1401,N_9606,N_9631);
or UO_1402 (O_1402,N_9568,N_9714);
or UO_1403 (O_1403,N_9947,N_9553);
or UO_1404 (O_1404,N_9830,N_9811);
or UO_1405 (O_1405,N_9528,N_9652);
nor UO_1406 (O_1406,N_9867,N_9877);
nand UO_1407 (O_1407,N_9630,N_9658);
nand UO_1408 (O_1408,N_9840,N_9871);
and UO_1409 (O_1409,N_9715,N_9872);
nand UO_1410 (O_1410,N_9584,N_9956);
or UO_1411 (O_1411,N_9834,N_9869);
and UO_1412 (O_1412,N_9728,N_9717);
nor UO_1413 (O_1413,N_9545,N_9833);
and UO_1414 (O_1414,N_9830,N_9661);
or UO_1415 (O_1415,N_9574,N_9999);
nand UO_1416 (O_1416,N_9633,N_9566);
and UO_1417 (O_1417,N_9706,N_9657);
or UO_1418 (O_1418,N_9709,N_9900);
nand UO_1419 (O_1419,N_9727,N_9932);
nor UO_1420 (O_1420,N_9608,N_9796);
nand UO_1421 (O_1421,N_9693,N_9583);
or UO_1422 (O_1422,N_9567,N_9852);
nor UO_1423 (O_1423,N_9821,N_9510);
nor UO_1424 (O_1424,N_9965,N_9708);
nand UO_1425 (O_1425,N_9750,N_9862);
or UO_1426 (O_1426,N_9679,N_9875);
nand UO_1427 (O_1427,N_9668,N_9991);
and UO_1428 (O_1428,N_9634,N_9713);
nor UO_1429 (O_1429,N_9526,N_9602);
nor UO_1430 (O_1430,N_9620,N_9788);
nor UO_1431 (O_1431,N_9528,N_9860);
nand UO_1432 (O_1432,N_9749,N_9658);
nand UO_1433 (O_1433,N_9811,N_9582);
xor UO_1434 (O_1434,N_9726,N_9986);
and UO_1435 (O_1435,N_9817,N_9516);
and UO_1436 (O_1436,N_9601,N_9868);
nand UO_1437 (O_1437,N_9682,N_9734);
nor UO_1438 (O_1438,N_9934,N_9724);
or UO_1439 (O_1439,N_9597,N_9899);
nor UO_1440 (O_1440,N_9781,N_9977);
nand UO_1441 (O_1441,N_9771,N_9647);
xor UO_1442 (O_1442,N_9970,N_9529);
nor UO_1443 (O_1443,N_9727,N_9840);
or UO_1444 (O_1444,N_9805,N_9544);
nor UO_1445 (O_1445,N_9550,N_9695);
nor UO_1446 (O_1446,N_9849,N_9896);
and UO_1447 (O_1447,N_9586,N_9721);
or UO_1448 (O_1448,N_9863,N_9782);
nor UO_1449 (O_1449,N_9623,N_9530);
nor UO_1450 (O_1450,N_9775,N_9546);
and UO_1451 (O_1451,N_9609,N_9585);
nand UO_1452 (O_1452,N_9620,N_9918);
and UO_1453 (O_1453,N_9724,N_9691);
or UO_1454 (O_1454,N_9613,N_9996);
nand UO_1455 (O_1455,N_9868,N_9668);
or UO_1456 (O_1456,N_9842,N_9896);
and UO_1457 (O_1457,N_9509,N_9703);
nor UO_1458 (O_1458,N_9673,N_9654);
nand UO_1459 (O_1459,N_9656,N_9505);
nor UO_1460 (O_1460,N_9952,N_9800);
nor UO_1461 (O_1461,N_9597,N_9861);
nand UO_1462 (O_1462,N_9951,N_9796);
nor UO_1463 (O_1463,N_9665,N_9746);
or UO_1464 (O_1464,N_9933,N_9907);
nand UO_1465 (O_1465,N_9839,N_9575);
xnor UO_1466 (O_1466,N_9520,N_9507);
nand UO_1467 (O_1467,N_9787,N_9793);
and UO_1468 (O_1468,N_9902,N_9612);
nand UO_1469 (O_1469,N_9811,N_9719);
and UO_1470 (O_1470,N_9976,N_9983);
and UO_1471 (O_1471,N_9590,N_9696);
nor UO_1472 (O_1472,N_9503,N_9500);
nor UO_1473 (O_1473,N_9780,N_9764);
nand UO_1474 (O_1474,N_9720,N_9629);
nand UO_1475 (O_1475,N_9881,N_9646);
or UO_1476 (O_1476,N_9796,N_9959);
and UO_1477 (O_1477,N_9574,N_9950);
nand UO_1478 (O_1478,N_9866,N_9787);
nor UO_1479 (O_1479,N_9564,N_9770);
nand UO_1480 (O_1480,N_9786,N_9590);
and UO_1481 (O_1481,N_9775,N_9744);
nand UO_1482 (O_1482,N_9647,N_9774);
nor UO_1483 (O_1483,N_9570,N_9550);
nor UO_1484 (O_1484,N_9519,N_9781);
nand UO_1485 (O_1485,N_9719,N_9678);
nand UO_1486 (O_1486,N_9845,N_9842);
and UO_1487 (O_1487,N_9626,N_9799);
nand UO_1488 (O_1488,N_9839,N_9618);
and UO_1489 (O_1489,N_9982,N_9991);
and UO_1490 (O_1490,N_9845,N_9599);
nor UO_1491 (O_1491,N_9942,N_9767);
nor UO_1492 (O_1492,N_9919,N_9892);
nand UO_1493 (O_1493,N_9759,N_9563);
nand UO_1494 (O_1494,N_9691,N_9726);
nor UO_1495 (O_1495,N_9852,N_9715);
xor UO_1496 (O_1496,N_9533,N_9754);
or UO_1497 (O_1497,N_9834,N_9743);
or UO_1498 (O_1498,N_9937,N_9530);
nand UO_1499 (O_1499,N_9610,N_9896);
endmodule