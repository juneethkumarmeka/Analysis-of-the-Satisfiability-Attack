module basic_500_3000_500_6_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_405,In_245);
nand U1 (N_1,In_393,In_208);
and U2 (N_2,In_427,In_314);
or U3 (N_3,In_154,In_97);
nor U4 (N_4,In_306,In_143);
and U5 (N_5,In_167,In_230);
nand U6 (N_6,In_441,In_304);
and U7 (N_7,In_300,In_342);
or U8 (N_8,In_161,In_407);
nor U9 (N_9,In_163,In_11);
nand U10 (N_10,In_267,In_364);
or U11 (N_11,In_9,In_375);
or U12 (N_12,In_225,In_212);
xor U13 (N_13,In_8,In_6);
nand U14 (N_14,In_403,In_482);
and U15 (N_15,In_265,In_30);
or U16 (N_16,In_88,In_247);
and U17 (N_17,In_79,In_384);
nor U18 (N_18,In_246,In_227);
nor U19 (N_19,In_328,In_148);
or U20 (N_20,In_268,In_372);
nor U21 (N_21,In_138,In_293);
and U22 (N_22,In_152,In_63);
nor U23 (N_23,In_471,In_305);
or U24 (N_24,In_32,In_447);
nand U25 (N_25,In_68,In_62);
nor U26 (N_26,In_254,In_318);
nor U27 (N_27,In_186,In_81);
and U28 (N_28,In_307,In_111);
and U29 (N_29,In_324,In_192);
nor U30 (N_30,In_7,In_402);
and U31 (N_31,In_121,In_115);
nand U32 (N_32,In_353,In_223);
nor U33 (N_33,In_90,In_352);
or U34 (N_34,In_224,In_359);
and U35 (N_35,In_43,In_50);
and U36 (N_36,In_363,In_101);
or U37 (N_37,In_226,In_423);
nand U38 (N_38,In_426,In_58);
or U39 (N_39,In_432,In_151);
nor U40 (N_40,In_128,In_309);
nor U41 (N_41,In_477,In_44);
nor U42 (N_42,In_467,In_140);
nor U43 (N_43,In_498,In_462);
or U44 (N_44,In_214,In_181);
nand U45 (N_45,In_253,In_455);
and U46 (N_46,In_266,In_459);
nand U47 (N_47,In_70,In_345);
and U48 (N_48,In_136,In_395);
or U49 (N_49,In_271,In_178);
or U50 (N_50,In_234,In_237);
nor U51 (N_51,In_67,In_458);
or U52 (N_52,In_53,In_107);
nor U53 (N_53,In_415,In_145);
nand U54 (N_54,In_380,In_262);
and U55 (N_55,In_4,In_84);
or U56 (N_56,In_444,In_366);
nor U57 (N_57,In_40,In_59);
nand U58 (N_58,In_113,In_235);
nand U59 (N_59,In_220,In_326);
nor U60 (N_60,In_48,In_311);
and U61 (N_61,In_292,In_313);
and U62 (N_62,In_41,In_85);
nor U63 (N_63,In_75,In_351);
and U64 (N_64,In_382,In_346);
or U65 (N_65,In_485,In_171);
or U66 (N_66,In_1,In_422);
nand U67 (N_67,In_492,In_57);
or U68 (N_68,In_93,In_408);
or U69 (N_69,In_396,In_21);
or U70 (N_70,In_451,In_251);
and U71 (N_71,In_103,In_435);
nand U72 (N_72,In_312,In_199);
or U73 (N_73,In_406,In_46);
nor U74 (N_74,In_184,In_404);
or U75 (N_75,In_26,In_179);
and U76 (N_76,In_278,In_474);
and U77 (N_77,In_157,In_155);
and U78 (N_78,In_187,In_277);
or U79 (N_79,In_218,In_0);
or U80 (N_80,In_259,In_354);
and U81 (N_81,In_95,In_117);
and U82 (N_82,In_490,In_164);
and U83 (N_83,In_159,In_409);
nand U84 (N_84,In_219,In_410);
or U85 (N_85,In_196,In_487);
nor U86 (N_86,In_344,In_373);
nand U87 (N_87,In_130,In_466);
and U88 (N_88,In_499,In_340);
and U89 (N_89,In_480,In_213);
nor U90 (N_90,In_54,In_102);
and U91 (N_91,In_486,In_473);
nand U92 (N_92,In_80,In_98);
nand U93 (N_93,In_356,In_270);
and U94 (N_94,In_478,In_190);
nor U95 (N_95,In_185,In_453);
nand U96 (N_96,In_420,In_132);
and U97 (N_97,In_35,In_24);
nand U98 (N_98,In_83,In_329);
nand U99 (N_99,In_233,In_289);
nand U100 (N_100,In_175,In_39);
nor U101 (N_101,In_169,In_29);
nand U102 (N_102,In_436,In_442);
or U103 (N_103,In_371,In_193);
and U104 (N_104,In_51,In_123);
nor U105 (N_105,In_394,In_446);
nor U106 (N_106,In_82,In_149);
and U107 (N_107,In_495,In_18);
nor U108 (N_108,In_460,In_298);
nor U109 (N_109,In_3,In_338);
nand U110 (N_110,In_28,In_481);
or U111 (N_111,In_355,In_135);
nor U112 (N_112,In_286,In_476);
or U113 (N_113,In_86,In_288);
nand U114 (N_114,In_176,In_64);
and U115 (N_115,In_74,In_147);
nor U116 (N_116,In_20,In_320);
or U117 (N_117,In_78,In_217);
nand U118 (N_118,In_461,In_439);
and U119 (N_119,In_379,In_378);
nor U120 (N_120,In_114,In_390);
or U121 (N_121,In_297,In_470);
or U122 (N_122,In_189,In_2);
or U123 (N_123,In_183,In_391);
and U124 (N_124,In_285,In_291);
or U125 (N_125,In_308,In_197);
xnor U126 (N_126,In_469,In_388);
and U127 (N_127,In_129,In_445);
or U128 (N_128,In_367,In_15);
nor U129 (N_129,In_350,In_489);
nor U130 (N_130,In_456,In_497);
and U131 (N_131,In_399,In_437);
nand U132 (N_132,In_66,In_116);
and U133 (N_133,In_331,In_448);
or U134 (N_134,In_295,In_60);
and U135 (N_135,In_413,In_238);
or U136 (N_136,In_330,In_275);
nand U137 (N_137,In_216,In_258);
xnor U138 (N_138,In_87,In_463);
nand U139 (N_139,In_398,In_494);
and U140 (N_140,In_207,In_210);
or U141 (N_141,In_411,In_142);
nor U142 (N_142,In_333,In_301);
or U143 (N_143,In_170,In_177);
nand U144 (N_144,In_61,In_110);
and U145 (N_145,In_269,In_325);
or U146 (N_146,In_284,In_361);
nand U147 (N_147,In_72,In_17);
nor U148 (N_148,In_194,In_434);
nor U149 (N_149,In_209,In_389);
or U150 (N_150,In_249,In_200);
and U151 (N_151,In_335,In_174);
nor U152 (N_152,In_488,In_464);
and U153 (N_153,In_141,In_12);
and U154 (N_154,In_47,In_430);
or U155 (N_155,In_369,In_457);
nand U156 (N_156,In_228,In_341);
nand U157 (N_157,In_358,In_336);
or U158 (N_158,In_45,In_133);
nand U159 (N_159,In_146,In_180);
and U160 (N_160,In_160,In_118);
or U161 (N_161,In_315,In_374);
nor U162 (N_162,In_401,In_438);
nor U163 (N_163,In_327,In_440);
or U164 (N_164,In_250,In_112);
nor U165 (N_165,In_5,In_319);
nor U166 (N_166,In_376,In_365);
nand U167 (N_167,In_263,In_303);
nor U168 (N_168,In_222,In_198);
nand U169 (N_169,In_243,In_387);
or U170 (N_170,In_424,In_317);
or U171 (N_171,In_27,In_281);
or U172 (N_172,In_362,In_491);
or U173 (N_173,In_96,In_13);
or U174 (N_174,In_231,In_195);
and U175 (N_175,In_450,In_120);
nor U176 (N_176,In_343,In_19);
nand U177 (N_177,In_273,In_418);
or U178 (N_178,In_125,In_144);
or U179 (N_179,In_465,In_412);
nor U180 (N_180,In_261,In_274);
or U181 (N_181,In_472,In_256);
nor U182 (N_182,In_139,In_166);
nand U183 (N_183,In_377,In_240);
and U184 (N_184,In_165,In_153);
nand U185 (N_185,In_36,In_94);
nor U186 (N_186,In_202,In_236);
or U187 (N_187,In_443,In_150);
nor U188 (N_188,In_201,In_119);
nand U189 (N_189,In_334,In_203);
nor U190 (N_190,In_14,In_56);
xnor U191 (N_191,In_299,In_414);
nand U192 (N_192,In_484,In_386);
or U193 (N_193,In_349,In_296);
nand U194 (N_194,In_23,In_272);
nand U195 (N_195,In_204,In_429);
or U196 (N_196,In_321,In_134);
nor U197 (N_197,In_156,In_168);
or U198 (N_198,In_348,In_105);
nor U199 (N_199,In_25,In_126);
and U200 (N_200,In_280,In_357);
nor U201 (N_201,In_10,In_34);
and U202 (N_202,In_158,In_22);
or U203 (N_203,In_323,In_241);
or U204 (N_204,In_496,In_475);
nand U205 (N_205,In_479,In_287);
and U206 (N_206,In_232,In_173);
nor U207 (N_207,In_428,In_392);
nor U208 (N_208,In_124,In_73);
or U209 (N_209,In_127,In_322);
or U210 (N_210,In_221,In_360);
or U211 (N_211,In_255,In_182);
nor U212 (N_212,In_122,In_417);
or U213 (N_213,In_76,In_172);
nand U214 (N_214,In_421,In_37);
and U215 (N_215,In_65,In_91);
and U216 (N_216,In_452,In_493);
nor U217 (N_217,In_397,In_248);
nor U218 (N_218,In_400,In_191);
and U219 (N_219,In_282,In_211);
nand U220 (N_220,In_468,In_483);
nor U221 (N_221,In_381,In_310);
nand U222 (N_222,In_215,In_108);
nand U223 (N_223,In_279,In_283);
and U224 (N_224,In_42,In_416);
or U225 (N_225,In_52,In_260);
or U226 (N_226,In_89,In_38);
or U227 (N_227,In_370,In_229);
and U228 (N_228,In_454,In_162);
nand U229 (N_229,In_239,In_109);
and U230 (N_230,In_431,In_383);
nor U231 (N_231,In_332,In_316);
nand U232 (N_232,In_264,In_419);
and U233 (N_233,In_100,In_276);
nand U234 (N_234,In_92,In_69);
or U235 (N_235,In_425,In_77);
xor U236 (N_236,In_337,In_104);
and U237 (N_237,In_206,In_368);
nand U238 (N_238,In_290,In_137);
nor U239 (N_239,In_55,In_433);
and U240 (N_240,In_385,In_99);
or U241 (N_241,In_339,In_294);
nand U242 (N_242,In_244,In_131);
nor U243 (N_243,In_347,In_302);
nand U244 (N_244,In_257,In_106);
and U245 (N_245,In_188,In_449);
or U246 (N_246,In_252,In_49);
nand U247 (N_247,In_16,In_205);
nor U248 (N_248,In_242,In_71);
and U249 (N_249,In_31,In_33);
nand U250 (N_250,In_68,In_474);
nand U251 (N_251,In_410,In_115);
nand U252 (N_252,In_420,In_156);
and U253 (N_253,In_438,In_330);
nand U254 (N_254,In_311,In_481);
and U255 (N_255,In_48,In_315);
xor U256 (N_256,In_426,In_113);
nand U257 (N_257,In_31,In_60);
xnor U258 (N_258,In_420,In_416);
or U259 (N_259,In_240,In_301);
and U260 (N_260,In_39,In_463);
or U261 (N_261,In_257,In_346);
or U262 (N_262,In_20,In_280);
xor U263 (N_263,In_23,In_29);
nor U264 (N_264,In_314,In_381);
or U265 (N_265,In_248,In_112);
and U266 (N_266,In_482,In_203);
and U267 (N_267,In_418,In_20);
nor U268 (N_268,In_443,In_166);
or U269 (N_269,In_243,In_217);
or U270 (N_270,In_266,In_358);
and U271 (N_271,In_41,In_483);
nor U272 (N_272,In_342,In_61);
or U273 (N_273,In_391,In_474);
nand U274 (N_274,In_427,In_131);
nor U275 (N_275,In_61,In_251);
or U276 (N_276,In_232,In_268);
or U277 (N_277,In_28,In_222);
and U278 (N_278,In_304,In_15);
nand U279 (N_279,In_138,In_291);
nor U280 (N_280,In_291,In_19);
and U281 (N_281,In_105,In_260);
nor U282 (N_282,In_311,In_497);
or U283 (N_283,In_338,In_349);
or U284 (N_284,In_46,In_201);
or U285 (N_285,In_347,In_380);
or U286 (N_286,In_155,In_425);
and U287 (N_287,In_416,In_146);
and U288 (N_288,In_71,In_102);
or U289 (N_289,In_331,In_219);
nand U290 (N_290,In_217,In_153);
nand U291 (N_291,In_13,In_275);
and U292 (N_292,In_181,In_412);
or U293 (N_293,In_321,In_189);
nor U294 (N_294,In_213,In_301);
and U295 (N_295,In_3,In_410);
or U296 (N_296,In_286,In_326);
nor U297 (N_297,In_396,In_205);
or U298 (N_298,In_189,In_157);
or U299 (N_299,In_63,In_335);
or U300 (N_300,In_281,In_33);
nor U301 (N_301,In_460,In_247);
or U302 (N_302,In_424,In_320);
nand U303 (N_303,In_414,In_225);
and U304 (N_304,In_480,In_162);
and U305 (N_305,In_129,In_134);
nor U306 (N_306,In_189,In_108);
or U307 (N_307,In_219,In_90);
nor U308 (N_308,In_449,In_84);
or U309 (N_309,In_72,In_477);
or U310 (N_310,In_157,In_364);
nor U311 (N_311,In_318,In_442);
nor U312 (N_312,In_377,In_332);
nor U313 (N_313,In_248,In_216);
nor U314 (N_314,In_143,In_405);
nand U315 (N_315,In_475,In_142);
or U316 (N_316,In_52,In_252);
nand U317 (N_317,In_287,In_100);
nand U318 (N_318,In_163,In_337);
and U319 (N_319,In_224,In_87);
or U320 (N_320,In_361,In_20);
and U321 (N_321,In_174,In_61);
nor U322 (N_322,In_234,In_269);
nor U323 (N_323,In_118,In_412);
nand U324 (N_324,In_229,In_206);
or U325 (N_325,In_339,In_156);
or U326 (N_326,In_294,In_61);
nand U327 (N_327,In_412,In_219);
and U328 (N_328,In_256,In_193);
and U329 (N_329,In_375,In_373);
nor U330 (N_330,In_308,In_143);
and U331 (N_331,In_332,In_219);
nor U332 (N_332,In_349,In_66);
nand U333 (N_333,In_334,In_441);
and U334 (N_334,In_215,In_259);
nand U335 (N_335,In_194,In_71);
nand U336 (N_336,In_438,In_394);
nand U337 (N_337,In_151,In_443);
nand U338 (N_338,In_486,In_10);
nand U339 (N_339,In_158,In_320);
nand U340 (N_340,In_302,In_134);
nor U341 (N_341,In_49,In_454);
nor U342 (N_342,In_371,In_416);
nand U343 (N_343,In_339,In_425);
nand U344 (N_344,In_207,In_65);
nor U345 (N_345,In_104,In_272);
or U346 (N_346,In_8,In_365);
and U347 (N_347,In_24,In_44);
nand U348 (N_348,In_72,In_32);
or U349 (N_349,In_203,In_138);
or U350 (N_350,In_243,In_306);
and U351 (N_351,In_16,In_431);
and U352 (N_352,In_209,In_283);
nand U353 (N_353,In_216,In_417);
nand U354 (N_354,In_57,In_384);
nand U355 (N_355,In_250,In_145);
or U356 (N_356,In_411,In_132);
and U357 (N_357,In_53,In_189);
or U358 (N_358,In_240,In_408);
or U359 (N_359,In_485,In_285);
nor U360 (N_360,In_108,In_468);
nor U361 (N_361,In_122,In_111);
nand U362 (N_362,In_317,In_4);
and U363 (N_363,In_106,In_113);
and U364 (N_364,In_10,In_406);
or U365 (N_365,In_325,In_199);
nor U366 (N_366,In_174,In_451);
nand U367 (N_367,In_379,In_26);
nand U368 (N_368,In_324,In_120);
nand U369 (N_369,In_339,In_27);
nand U370 (N_370,In_399,In_356);
xnor U371 (N_371,In_384,In_322);
and U372 (N_372,In_356,In_181);
or U373 (N_373,In_100,In_193);
nand U374 (N_374,In_236,In_176);
nor U375 (N_375,In_53,In_80);
nand U376 (N_376,In_377,In_153);
nor U377 (N_377,In_180,In_318);
nand U378 (N_378,In_423,In_339);
or U379 (N_379,In_71,In_150);
nand U380 (N_380,In_146,In_153);
nand U381 (N_381,In_37,In_69);
and U382 (N_382,In_373,In_226);
and U383 (N_383,In_54,In_31);
nor U384 (N_384,In_221,In_403);
nor U385 (N_385,In_215,In_477);
and U386 (N_386,In_98,In_492);
nor U387 (N_387,In_318,In_458);
and U388 (N_388,In_188,In_467);
and U389 (N_389,In_336,In_430);
nand U390 (N_390,In_114,In_90);
or U391 (N_391,In_67,In_401);
or U392 (N_392,In_292,In_68);
nor U393 (N_393,In_326,In_459);
or U394 (N_394,In_481,In_137);
nand U395 (N_395,In_4,In_213);
nor U396 (N_396,In_186,In_79);
nor U397 (N_397,In_303,In_88);
or U398 (N_398,In_427,In_363);
or U399 (N_399,In_219,In_45);
nand U400 (N_400,In_348,In_404);
or U401 (N_401,In_368,In_461);
and U402 (N_402,In_19,In_101);
and U403 (N_403,In_18,In_200);
or U404 (N_404,In_94,In_35);
nor U405 (N_405,In_317,In_292);
or U406 (N_406,In_385,In_281);
or U407 (N_407,In_369,In_463);
and U408 (N_408,In_49,In_358);
nor U409 (N_409,In_165,In_403);
and U410 (N_410,In_222,In_448);
nand U411 (N_411,In_145,In_381);
nand U412 (N_412,In_98,In_489);
and U413 (N_413,In_421,In_310);
and U414 (N_414,In_10,In_489);
nor U415 (N_415,In_56,In_289);
nand U416 (N_416,In_71,In_406);
and U417 (N_417,In_144,In_250);
and U418 (N_418,In_374,In_245);
and U419 (N_419,In_446,In_270);
nand U420 (N_420,In_435,In_98);
or U421 (N_421,In_362,In_385);
nand U422 (N_422,In_316,In_250);
or U423 (N_423,In_418,In_129);
nand U424 (N_424,In_454,In_369);
nand U425 (N_425,In_463,In_440);
or U426 (N_426,In_357,In_194);
nand U427 (N_427,In_315,In_361);
nand U428 (N_428,In_397,In_259);
or U429 (N_429,In_234,In_253);
or U430 (N_430,In_144,In_342);
or U431 (N_431,In_279,In_62);
nor U432 (N_432,In_342,In_485);
or U433 (N_433,In_67,In_222);
nor U434 (N_434,In_437,In_206);
or U435 (N_435,In_482,In_287);
nor U436 (N_436,In_227,In_292);
nor U437 (N_437,In_188,In_377);
and U438 (N_438,In_297,In_137);
and U439 (N_439,In_312,In_70);
nand U440 (N_440,In_296,In_309);
nand U441 (N_441,In_139,In_302);
nor U442 (N_442,In_27,In_404);
and U443 (N_443,In_224,In_4);
or U444 (N_444,In_243,In_8);
xnor U445 (N_445,In_456,In_354);
and U446 (N_446,In_102,In_206);
xor U447 (N_447,In_63,In_175);
and U448 (N_448,In_353,In_452);
nand U449 (N_449,In_77,In_254);
nor U450 (N_450,In_314,In_179);
nor U451 (N_451,In_244,In_128);
or U452 (N_452,In_165,In_362);
nor U453 (N_453,In_53,In_371);
and U454 (N_454,In_253,In_383);
nor U455 (N_455,In_319,In_480);
nor U456 (N_456,In_200,In_47);
or U457 (N_457,In_86,In_358);
or U458 (N_458,In_80,In_443);
or U459 (N_459,In_166,In_309);
and U460 (N_460,In_58,In_320);
nand U461 (N_461,In_178,In_5);
nand U462 (N_462,In_119,In_21);
or U463 (N_463,In_20,In_4);
and U464 (N_464,In_46,In_132);
and U465 (N_465,In_114,In_231);
nor U466 (N_466,In_42,In_196);
or U467 (N_467,In_472,In_67);
nand U468 (N_468,In_443,In_2);
and U469 (N_469,In_338,In_100);
and U470 (N_470,In_21,In_309);
and U471 (N_471,In_94,In_435);
or U472 (N_472,In_467,In_405);
nand U473 (N_473,In_296,In_390);
and U474 (N_474,In_180,In_8);
and U475 (N_475,In_160,In_15);
or U476 (N_476,In_186,In_288);
and U477 (N_477,In_294,In_126);
nand U478 (N_478,In_472,In_411);
nor U479 (N_479,In_491,In_457);
nor U480 (N_480,In_33,In_144);
or U481 (N_481,In_152,In_493);
nor U482 (N_482,In_250,In_476);
nor U483 (N_483,In_284,In_115);
nor U484 (N_484,In_220,In_320);
nor U485 (N_485,In_176,In_377);
and U486 (N_486,In_331,In_451);
and U487 (N_487,In_145,In_176);
nor U488 (N_488,In_206,In_413);
or U489 (N_489,In_376,In_486);
or U490 (N_490,In_324,In_227);
or U491 (N_491,In_106,In_146);
and U492 (N_492,In_85,In_419);
or U493 (N_493,In_109,In_374);
nand U494 (N_494,In_13,In_367);
nor U495 (N_495,In_244,In_414);
nand U496 (N_496,In_332,In_438);
or U497 (N_497,In_139,In_174);
or U498 (N_498,In_262,In_171);
or U499 (N_499,In_310,In_220);
nand U500 (N_500,N_188,N_143);
or U501 (N_501,N_449,N_39);
nand U502 (N_502,N_339,N_44);
and U503 (N_503,N_483,N_231);
or U504 (N_504,N_368,N_267);
or U505 (N_505,N_302,N_111);
nor U506 (N_506,N_216,N_276);
or U507 (N_507,N_142,N_460);
nor U508 (N_508,N_357,N_319);
or U509 (N_509,N_448,N_346);
or U510 (N_510,N_380,N_323);
and U511 (N_511,N_164,N_22);
nor U512 (N_512,N_140,N_467);
and U513 (N_513,N_63,N_94);
nor U514 (N_514,N_208,N_107);
or U515 (N_515,N_345,N_292);
nand U516 (N_516,N_64,N_69);
and U517 (N_517,N_281,N_24);
and U518 (N_518,N_401,N_468);
nor U519 (N_519,N_415,N_322);
nand U520 (N_520,N_2,N_362);
nor U521 (N_521,N_106,N_241);
and U522 (N_522,N_299,N_251);
nor U523 (N_523,N_383,N_439);
nand U524 (N_524,N_489,N_77);
and U525 (N_525,N_366,N_156);
nand U526 (N_526,N_436,N_193);
nand U527 (N_527,N_286,N_414);
nor U528 (N_528,N_284,N_354);
or U529 (N_529,N_256,N_257);
or U530 (N_530,N_58,N_253);
nor U531 (N_531,N_499,N_228);
nand U532 (N_532,N_91,N_169);
and U533 (N_533,N_96,N_147);
and U534 (N_534,N_25,N_19);
or U535 (N_535,N_237,N_29);
or U536 (N_536,N_128,N_76);
nand U537 (N_537,N_78,N_443);
nor U538 (N_538,N_430,N_438);
nor U539 (N_539,N_240,N_360);
nand U540 (N_540,N_220,N_341);
or U541 (N_541,N_172,N_309);
nand U542 (N_542,N_297,N_125);
or U543 (N_543,N_325,N_373);
and U544 (N_544,N_60,N_494);
nand U545 (N_545,N_327,N_226);
nand U546 (N_546,N_404,N_173);
nand U547 (N_547,N_273,N_272);
nand U548 (N_548,N_264,N_202);
and U549 (N_549,N_308,N_334);
or U550 (N_550,N_459,N_473);
nand U551 (N_551,N_223,N_315);
nand U552 (N_552,N_218,N_375);
nand U553 (N_553,N_396,N_185);
or U554 (N_554,N_261,N_168);
or U555 (N_555,N_398,N_191);
and U556 (N_556,N_180,N_379);
and U557 (N_557,N_32,N_472);
or U558 (N_558,N_420,N_456);
nand U559 (N_559,N_303,N_392);
nand U560 (N_560,N_126,N_12);
nand U561 (N_561,N_498,N_482);
or U562 (N_562,N_219,N_310);
or U563 (N_563,N_407,N_381);
nand U564 (N_564,N_0,N_455);
or U565 (N_565,N_301,N_6);
or U566 (N_566,N_49,N_418);
or U567 (N_567,N_153,N_109);
or U568 (N_568,N_50,N_112);
nor U569 (N_569,N_217,N_38);
and U570 (N_570,N_440,N_386);
or U571 (N_571,N_409,N_437);
and U572 (N_572,N_361,N_464);
nand U573 (N_573,N_492,N_115);
nor U574 (N_574,N_119,N_283);
and U575 (N_575,N_422,N_305);
or U576 (N_576,N_210,N_350);
nand U577 (N_577,N_290,N_424);
nand U578 (N_578,N_141,N_371);
and U579 (N_579,N_213,N_389);
nor U580 (N_580,N_235,N_88);
nor U581 (N_581,N_83,N_280);
and U582 (N_582,N_453,N_470);
or U583 (N_583,N_26,N_127);
nand U584 (N_584,N_214,N_471);
nand U585 (N_585,N_197,N_461);
and U586 (N_586,N_356,N_355);
and U587 (N_587,N_16,N_313);
nand U588 (N_588,N_194,N_458);
nand U589 (N_589,N_203,N_370);
nor U590 (N_590,N_33,N_255);
nand U591 (N_591,N_137,N_359);
nand U592 (N_592,N_426,N_68);
nor U593 (N_593,N_87,N_343);
or U594 (N_594,N_433,N_377);
or U595 (N_595,N_4,N_340);
nand U596 (N_596,N_314,N_84);
or U597 (N_597,N_85,N_224);
or U598 (N_598,N_263,N_92);
and U599 (N_599,N_242,N_465);
nor U600 (N_600,N_363,N_417);
or U601 (N_601,N_294,N_42);
and U602 (N_602,N_174,N_189);
or U603 (N_603,N_55,N_3);
nor U604 (N_604,N_485,N_130);
or U605 (N_605,N_13,N_198);
nand U606 (N_606,N_333,N_391);
or U607 (N_607,N_387,N_411);
nand U608 (N_608,N_209,N_211);
nor U609 (N_609,N_56,N_104);
nor U610 (N_610,N_278,N_452);
nand U611 (N_611,N_488,N_479);
nor U612 (N_612,N_48,N_131);
nor U613 (N_613,N_221,N_434);
or U614 (N_614,N_116,N_187);
nand U615 (N_615,N_43,N_410);
and U616 (N_616,N_451,N_71);
nand U617 (N_617,N_167,N_195);
nor U618 (N_618,N_412,N_166);
nor U619 (N_619,N_178,N_245);
nor U620 (N_620,N_466,N_121);
and U621 (N_621,N_432,N_328);
nor U622 (N_622,N_306,N_154);
nor U623 (N_623,N_150,N_227);
nor U624 (N_624,N_399,N_484);
nor U625 (N_625,N_329,N_384);
nor U626 (N_626,N_457,N_159);
or U627 (N_627,N_160,N_10);
nor U628 (N_628,N_337,N_122);
nand U629 (N_629,N_165,N_408);
or U630 (N_630,N_332,N_120);
or U631 (N_631,N_136,N_249);
or U632 (N_632,N_289,N_490);
xor U633 (N_633,N_338,N_291);
nor U634 (N_634,N_177,N_207);
or U635 (N_635,N_474,N_271);
nand U636 (N_636,N_47,N_385);
and U637 (N_637,N_72,N_405);
and U638 (N_638,N_427,N_421);
or U639 (N_639,N_66,N_46);
and U640 (N_640,N_394,N_419);
nand U641 (N_641,N_236,N_206);
and U642 (N_642,N_36,N_365);
and U643 (N_643,N_446,N_390);
nand U644 (N_644,N_258,N_201);
nor U645 (N_645,N_425,N_145);
nor U646 (N_646,N_93,N_266);
nand U647 (N_647,N_311,N_254);
nor U648 (N_648,N_316,N_37);
or U649 (N_649,N_476,N_320);
nor U650 (N_650,N_15,N_183);
nor U651 (N_651,N_296,N_65);
or U652 (N_652,N_212,N_374);
nor U653 (N_653,N_288,N_435);
and U654 (N_654,N_133,N_59);
nor U655 (N_655,N_246,N_369);
xnor U656 (N_656,N_148,N_200);
and U657 (N_657,N_238,N_335);
nor U658 (N_658,N_11,N_428);
nand U659 (N_659,N_352,N_324);
nor U660 (N_660,N_139,N_239);
or U661 (N_661,N_9,N_395);
nor U662 (N_662,N_270,N_268);
nand U663 (N_663,N_454,N_393);
nor U664 (N_664,N_181,N_234);
nor U665 (N_665,N_232,N_481);
or U666 (N_666,N_30,N_113);
nand U667 (N_667,N_108,N_82);
or U668 (N_668,N_233,N_244);
nand U669 (N_669,N_250,N_486);
nor U670 (N_670,N_243,N_158);
nor U671 (N_671,N_31,N_259);
or U672 (N_672,N_28,N_469);
or U673 (N_673,N_20,N_182);
or U674 (N_674,N_372,N_34);
nor U675 (N_675,N_269,N_496);
nor U676 (N_676,N_493,N_51);
or U677 (N_677,N_17,N_406);
nor U678 (N_678,N_151,N_123);
nand U679 (N_679,N_230,N_57);
nand U680 (N_680,N_79,N_199);
nor U681 (N_681,N_388,N_40);
and U682 (N_682,N_215,N_429);
nand U683 (N_683,N_103,N_318);
nand U684 (N_684,N_248,N_70);
nand U685 (N_685,N_162,N_367);
and U686 (N_686,N_497,N_18);
or U687 (N_687,N_129,N_295);
nand U688 (N_688,N_447,N_14);
or U689 (N_689,N_382,N_229);
nand U690 (N_690,N_23,N_155);
and U691 (N_691,N_186,N_101);
nor U692 (N_692,N_348,N_347);
nand U693 (N_693,N_95,N_205);
or U694 (N_694,N_86,N_184);
nand U695 (N_695,N_45,N_7);
or U696 (N_696,N_431,N_416);
and U697 (N_697,N_252,N_358);
or U698 (N_698,N_98,N_402);
and U699 (N_699,N_376,N_105);
or U700 (N_700,N_204,N_152);
nor U701 (N_701,N_364,N_342);
or U702 (N_702,N_331,N_279);
or U703 (N_703,N_175,N_62);
nand U704 (N_704,N_442,N_190);
nand U705 (N_705,N_114,N_312);
or U706 (N_706,N_1,N_144);
nor U707 (N_707,N_277,N_491);
or U708 (N_708,N_61,N_225);
nand U709 (N_709,N_117,N_161);
and U710 (N_710,N_196,N_260);
and U711 (N_711,N_285,N_192);
and U712 (N_712,N_171,N_110);
nor U713 (N_713,N_179,N_27);
nand U714 (N_714,N_146,N_99);
nor U715 (N_715,N_463,N_330);
and U716 (N_716,N_41,N_282);
nand U717 (N_717,N_287,N_35);
nor U718 (N_718,N_326,N_450);
nand U719 (N_719,N_293,N_487);
nor U720 (N_720,N_124,N_134);
nor U721 (N_721,N_403,N_441);
and U722 (N_722,N_351,N_90);
nor U723 (N_723,N_321,N_75);
nand U724 (N_724,N_300,N_304);
and U725 (N_725,N_118,N_176);
nand U726 (N_726,N_5,N_344);
or U727 (N_727,N_307,N_477);
and U728 (N_728,N_53,N_475);
nor U729 (N_729,N_138,N_298);
nand U730 (N_730,N_413,N_400);
or U731 (N_731,N_52,N_317);
and U732 (N_732,N_265,N_170);
or U733 (N_733,N_445,N_336);
nor U734 (N_734,N_132,N_102);
nor U735 (N_735,N_97,N_353);
and U736 (N_736,N_495,N_89);
nand U737 (N_737,N_349,N_423);
or U738 (N_738,N_81,N_100);
nor U739 (N_739,N_247,N_54);
nand U740 (N_740,N_274,N_80);
nor U741 (N_741,N_8,N_163);
or U742 (N_742,N_444,N_149);
or U743 (N_743,N_397,N_135);
nand U744 (N_744,N_157,N_67);
and U745 (N_745,N_478,N_222);
or U746 (N_746,N_21,N_480);
nand U747 (N_747,N_462,N_275);
nand U748 (N_748,N_73,N_378);
xor U749 (N_749,N_74,N_262);
or U750 (N_750,N_279,N_271);
nor U751 (N_751,N_359,N_19);
and U752 (N_752,N_184,N_110);
nor U753 (N_753,N_91,N_353);
or U754 (N_754,N_112,N_206);
nor U755 (N_755,N_249,N_485);
nand U756 (N_756,N_11,N_448);
nor U757 (N_757,N_238,N_489);
or U758 (N_758,N_116,N_324);
nor U759 (N_759,N_10,N_244);
nor U760 (N_760,N_398,N_175);
nand U761 (N_761,N_307,N_12);
and U762 (N_762,N_407,N_116);
or U763 (N_763,N_333,N_49);
and U764 (N_764,N_203,N_183);
nand U765 (N_765,N_139,N_332);
and U766 (N_766,N_108,N_170);
or U767 (N_767,N_245,N_182);
nor U768 (N_768,N_87,N_395);
or U769 (N_769,N_432,N_126);
nor U770 (N_770,N_350,N_424);
and U771 (N_771,N_173,N_146);
nand U772 (N_772,N_25,N_365);
and U773 (N_773,N_470,N_94);
nand U774 (N_774,N_316,N_34);
and U775 (N_775,N_280,N_451);
nor U776 (N_776,N_248,N_383);
or U777 (N_777,N_339,N_252);
and U778 (N_778,N_332,N_465);
or U779 (N_779,N_412,N_258);
or U780 (N_780,N_480,N_401);
and U781 (N_781,N_383,N_8);
or U782 (N_782,N_446,N_228);
or U783 (N_783,N_142,N_194);
nand U784 (N_784,N_320,N_493);
and U785 (N_785,N_226,N_465);
nand U786 (N_786,N_486,N_39);
nor U787 (N_787,N_315,N_167);
or U788 (N_788,N_319,N_56);
and U789 (N_789,N_353,N_402);
nor U790 (N_790,N_0,N_279);
nand U791 (N_791,N_91,N_223);
and U792 (N_792,N_157,N_279);
or U793 (N_793,N_332,N_277);
nor U794 (N_794,N_47,N_434);
or U795 (N_795,N_445,N_120);
nor U796 (N_796,N_207,N_80);
or U797 (N_797,N_117,N_445);
and U798 (N_798,N_21,N_219);
nand U799 (N_799,N_301,N_103);
nand U800 (N_800,N_198,N_243);
or U801 (N_801,N_178,N_213);
and U802 (N_802,N_452,N_415);
nand U803 (N_803,N_382,N_8);
or U804 (N_804,N_373,N_272);
xor U805 (N_805,N_59,N_207);
and U806 (N_806,N_133,N_372);
and U807 (N_807,N_47,N_441);
or U808 (N_808,N_108,N_297);
nand U809 (N_809,N_435,N_32);
nand U810 (N_810,N_387,N_58);
nand U811 (N_811,N_299,N_51);
and U812 (N_812,N_104,N_427);
nand U813 (N_813,N_46,N_20);
nor U814 (N_814,N_15,N_132);
and U815 (N_815,N_254,N_252);
nor U816 (N_816,N_437,N_30);
nor U817 (N_817,N_92,N_368);
nor U818 (N_818,N_72,N_123);
nand U819 (N_819,N_228,N_251);
or U820 (N_820,N_434,N_416);
or U821 (N_821,N_282,N_441);
nor U822 (N_822,N_62,N_382);
nand U823 (N_823,N_148,N_163);
nand U824 (N_824,N_203,N_473);
and U825 (N_825,N_124,N_91);
nor U826 (N_826,N_43,N_165);
and U827 (N_827,N_244,N_101);
nand U828 (N_828,N_142,N_104);
nor U829 (N_829,N_294,N_273);
and U830 (N_830,N_72,N_151);
and U831 (N_831,N_7,N_433);
nor U832 (N_832,N_106,N_352);
nand U833 (N_833,N_124,N_43);
nor U834 (N_834,N_28,N_110);
nor U835 (N_835,N_495,N_236);
nor U836 (N_836,N_494,N_335);
and U837 (N_837,N_406,N_309);
nand U838 (N_838,N_279,N_128);
or U839 (N_839,N_152,N_391);
and U840 (N_840,N_99,N_241);
and U841 (N_841,N_428,N_201);
nor U842 (N_842,N_453,N_447);
nand U843 (N_843,N_336,N_77);
nand U844 (N_844,N_18,N_221);
nor U845 (N_845,N_250,N_227);
nand U846 (N_846,N_72,N_188);
or U847 (N_847,N_286,N_221);
and U848 (N_848,N_328,N_389);
nand U849 (N_849,N_124,N_53);
nand U850 (N_850,N_358,N_39);
nor U851 (N_851,N_56,N_219);
and U852 (N_852,N_306,N_46);
nor U853 (N_853,N_91,N_113);
and U854 (N_854,N_293,N_67);
nor U855 (N_855,N_207,N_471);
nor U856 (N_856,N_191,N_454);
and U857 (N_857,N_413,N_387);
nand U858 (N_858,N_87,N_101);
or U859 (N_859,N_109,N_425);
or U860 (N_860,N_176,N_394);
nand U861 (N_861,N_167,N_389);
or U862 (N_862,N_314,N_145);
and U863 (N_863,N_426,N_335);
and U864 (N_864,N_90,N_252);
and U865 (N_865,N_63,N_313);
and U866 (N_866,N_365,N_389);
nand U867 (N_867,N_222,N_448);
or U868 (N_868,N_64,N_42);
nor U869 (N_869,N_253,N_303);
nand U870 (N_870,N_96,N_304);
nand U871 (N_871,N_431,N_51);
nor U872 (N_872,N_272,N_243);
or U873 (N_873,N_173,N_289);
nand U874 (N_874,N_182,N_263);
nor U875 (N_875,N_263,N_38);
or U876 (N_876,N_492,N_122);
nor U877 (N_877,N_451,N_298);
nor U878 (N_878,N_315,N_109);
or U879 (N_879,N_485,N_409);
and U880 (N_880,N_278,N_318);
or U881 (N_881,N_9,N_444);
nand U882 (N_882,N_321,N_103);
and U883 (N_883,N_321,N_124);
or U884 (N_884,N_256,N_217);
or U885 (N_885,N_3,N_212);
nor U886 (N_886,N_430,N_122);
or U887 (N_887,N_55,N_247);
nand U888 (N_888,N_231,N_60);
and U889 (N_889,N_123,N_132);
nand U890 (N_890,N_375,N_293);
and U891 (N_891,N_368,N_142);
nand U892 (N_892,N_181,N_74);
nand U893 (N_893,N_169,N_134);
nor U894 (N_894,N_346,N_219);
or U895 (N_895,N_440,N_366);
or U896 (N_896,N_100,N_405);
nand U897 (N_897,N_42,N_126);
and U898 (N_898,N_32,N_270);
nor U899 (N_899,N_163,N_236);
nor U900 (N_900,N_179,N_287);
and U901 (N_901,N_262,N_169);
or U902 (N_902,N_468,N_16);
and U903 (N_903,N_26,N_72);
nand U904 (N_904,N_131,N_180);
and U905 (N_905,N_69,N_389);
and U906 (N_906,N_228,N_42);
nand U907 (N_907,N_173,N_123);
nand U908 (N_908,N_157,N_36);
and U909 (N_909,N_218,N_423);
nand U910 (N_910,N_404,N_312);
nor U911 (N_911,N_297,N_486);
and U912 (N_912,N_152,N_53);
nand U913 (N_913,N_154,N_70);
or U914 (N_914,N_478,N_302);
or U915 (N_915,N_345,N_130);
and U916 (N_916,N_146,N_358);
or U917 (N_917,N_178,N_252);
and U918 (N_918,N_50,N_115);
nand U919 (N_919,N_220,N_461);
nand U920 (N_920,N_491,N_208);
and U921 (N_921,N_53,N_454);
or U922 (N_922,N_485,N_1);
nand U923 (N_923,N_51,N_232);
and U924 (N_924,N_52,N_281);
nor U925 (N_925,N_81,N_280);
nor U926 (N_926,N_355,N_457);
nand U927 (N_927,N_64,N_477);
nor U928 (N_928,N_13,N_98);
nor U929 (N_929,N_452,N_181);
nor U930 (N_930,N_322,N_346);
nand U931 (N_931,N_350,N_216);
or U932 (N_932,N_455,N_271);
nor U933 (N_933,N_499,N_415);
nand U934 (N_934,N_349,N_146);
nor U935 (N_935,N_194,N_5);
or U936 (N_936,N_343,N_440);
nor U937 (N_937,N_249,N_43);
or U938 (N_938,N_288,N_451);
and U939 (N_939,N_354,N_49);
or U940 (N_940,N_294,N_203);
or U941 (N_941,N_312,N_309);
nand U942 (N_942,N_211,N_274);
or U943 (N_943,N_392,N_198);
nand U944 (N_944,N_493,N_52);
nand U945 (N_945,N_17,N_331);
nand U946 (N_946,N_108,N_178);
nor U947 (N_947,N_448,N_361);
or U948 (N_948,N_369,N_125);
or U949 (N_949,N_460,N_371);
and U950 (N_950,N_254,N_173);
and U951 (N_951,N_297,N_63);
nor U952 (N_952,N_168,N_367);
nand U953 (N_953,N_373,N_192);
nor U954 (N_954,N_472,N_282);
nand U955 (N_955,N_173,N_447);
nor U956 (N_956,N_195,N_404);
and U957 (N_957,N_97,N_23);
nor U958 (N_958,N_267,N_111);
nor U959 (N_959,N_205,N_2);
nor U960 (N_960,N_408,N_460);
nand U961 (N_961,N_395,N_115);
or U962 (N_962,N_192,N_222);
and U963 (N_963,N_461,N_84);
nand U964 (N_964,N_359,N_370);
and U965 (N_965,N_73,N_263);
and U966 (N_966,N_263,N_240);
or U967 (N_967,N_190,N_377);
or U968 (N_968,N_175,N_121);
nor U969 (N_969,N_466,N_116);
or U970 (N_970,N_404,N_224);
and U971 (N_971,N_259,N_414);
and U972 (N_972,N_334,N_191);
nor U973 (N_973,N_195,N_435);
nor U974 (N_974,N_447,N_495);
nor U975 (N_975,N_347,N_338);
nand U976 (N_976,N_50,N_139);
nand U977 (N_977,N_443,N_225);
and U978 (N_978,N_43,N_320);
and U979 (N_979,N_150,N_84);
nor U980 (N_980,N_39,N_108);
and U981 (N_981,N_467,N_488);
nor U982 (N_982,N_130,N_231);
nor U983 (N_983,N_167,N_148);
nor U984 (N_984,N_245,N_335);
nand U985 (N_985,N_126,N_18);
xnor U986 (N_986,N_398,N_166);
nor U987 (N_987,N_402,N_317);
nor U988 (N_988,N_399,N_19);
or U989 (N_989,N_2,N_28);
nand U990 (N_990,N_297,N_260);
nand U991 (N_991,N_75,N_120);
nor U992 (N_992,N_427,N_174);
or U993 (N_993,N_383,N_41);
nor U994 (N_994,N_382,N_266);
and U995 (N_995,N_228,N_448);
nor U996 (N_996,N_190,N_332);
or U997 (N_997,N_274,N_43);
and U998 (N_998,N_472,N_110);
nor U999 (N_999,N_20,N_149);
nand U1000 (N_1000,N_945,N_913);
or U1001 (N_1001,N_952,N_600);
or U1002 (N_1002,N_958,N_699);
or U1003 (N_1003,N_921,N_638);
xnor U1004 (N_1004,N_550,N_658);
and U1005 (N_1005,N_647,N_525);
nand U1006 (N_1006,N_665,N_948);
nor U1007 (N_1007,N_846,N_552);
and U1008 (N_1008,N_624,N_907);
nor U1009 (N_1009,N_816,N_875);
nor U1010 (N_1010,N_575,N_643);
and U1011 (N_1011,N_630,N_605);
or U1012 (N_1012,N_912,N_750);
and U1013 (N_1013,N_946,N_668);
nor U1014 (N_1014,N_740,N_811);
nor U1015 (N_1015,N_863,N_723);
nor U1016 (N_1016,N_993,N_865);
and U1017 (N_1017,N_814,N_854);
and U1018 (N_1018,N_579,N_646);
or U1019 (N_1019,N_978,N_687);
nor U1020 (N_1020,N_695,N_726);
or U1021 (N_1021,N_756,N_562);
or U1022 (N_1022,N_663,N_753);
nand U1023 (N_1023,N_804,N_793);
nand U1024 (N_1024,N_620,N_901);
nor U1025 (N_1025,N_654,N_971);
nand U1026 (N_1026,N_869,N_806);
or U1027 (N_1027,N_965,N_634);
and U1028 (N_1028,N_724,N_833);
and U1029 (N_1029,N_932,N_760);
and U1030 (N_1030,N_610,N_531);
or U1031 (N_1031,N_914,N_559);
or U1032 (N_1032,N_789,N_836);
nor U1033 (N_1033,N_761,N_714);
or U1034 (N_1034,N_955,N_547);
nand U1035 (N_1035,N_848,N_573);
nand U1036 (N_1036,N_902,N_667);
or U1037 (N_1037,N_651,N_784);
nor U1038 (N_1038,N_669,N_815);
nand U1039 (N_1039,N_592,N_617);
or U1040 (N_1040,N_953,N_572);
nor U1041 (N_1041,N_877,N_904);
nor U1042 (N_1042,N_515,N_922);
and U1043 (N_1043,N_960,N_765);
and U1044 (N_1044,N_707,N_650);
nor U1045 (N_1045,N_888,N_763);
nand U1046 (N_1046,N_596,N_995);
nand U1047 (N_1047,N_749,N_856);
and U1048 (N_1048,N_659,N_839);
and U1049 (N_1049,N_817,N_867);
and U1050 (N_1050,N_641,N_849);
or U1051 (N_1051,N_537,N_717);
and U1052 (N_1052,N_631,N_551);
or U1053 (N_1053,N_535,N_589);
nand U1054 (N_1054,N_544,N_940);
nand U1055 (N_1055,N_770,N_671);
nand U1056 (N_1056,N_871,N_801);
or U1057 (N_1057,N_564,N_734);
nor U1058 (N_1058,N_730,N_838);
or U1059 (N_1059,N_616,N_673);
nand U1060 (N_1060,N_924,N_644);
nor U1061 (N_1061,N_529,N_937);
nor U1062 (N_1062,N_794,N_949);
nand U1063 (N_1063,N_828,N_969);
or U1064 (N_1064,N_516,N_633);
or U1065 (N_1065,N_582,N_601);
nor U1066 (N_1066,N_766,N_825);
nand U1067 (N_1067,N_686,N_855);
or U1068 (N_1068,N_892,N_521);
or U1069 (N_1069,N_927,N_786);
or U1070 (N_1070,N_731,N_994);
or U1071 (N_1071,N_859,N_939);
or U1072 (N_1072,N_858,N_983);
nand U1073 (N_1073,N_632,N_762);
nand U1074 (N_1074,N_788,N_956);
nand U1075 (N_1075,N_915,N_626);
nand U1076 (N_1076,N_870,N_660);
and U1077 (N_1077,N_712,N_885);
nor U1078 (N_1078,N_951,N_853);
nor U1079 (N_1079,N_557,N_581);
or U1080 (N_1080,N_539,N_519);
nand U1081 (N_1081,N_841,N_934);
nand U1082 (N_1082,N_642,N_501);
nor U1083 (N_1083,N_942,N_840);
nand U1084 (N_1084,N_505,N_586);
nor U1085 (N_1085,N_925,N_664);
and U1086 (N_1086,N_874,N_889);
nand U1087 (N_1087,N_908,N_797);
or U1088 (N_1088,N_536,N_943);
nor U1089 (N_1089,N_688,N_742);
nand U1090 (N_1090,N_694,N_812);
or U1091 (N_1091,N_928,N_670);
nand U1092 (N_1092,N_509,N_523);
or U1093 (N_1093,N_627,N_987);
and U1094 (N_1094,N_538,N_984);
and U1095 (N_1095,N_612,N_944);
or U1096 (N_1096,N_549,N_713);
xnor U1097 (N_1097,N_795,N_689);
nand U1098 (N_1098,N_615,N_530);
and U1099 (N_1099,N_502,N_704);
or U1100 (N_1100,N_703,N_852);
and U1101 (N_1101,N_567,N_798);
or U1102 (N_1102,N_974,N_999);
nor U1103 (N_1103,N_648,N_986);
or U1104 (N_1104,N_662,N_998);
and U1105 (N_1105,N_716,N_819);
nor U1106 (N_1106,N_866,N_963);
or U1107 (N_1107,N_930,N_850);
nor U1108 (N_1108,N_781,N_935);
nand U1109 (N_1109,N_653,N_533);
nand U1110 (N_1110,N_715,N_560);
or U1111 (N_1111,N_861,N_792);
or U1112 (N_1112,N_545,N_520);
or U1113 (N_1113,N_656,N_543);
or U1114 (N_1114,N_918,N_843);
nor U1115 (N_1115,N_587,N_973);
nor U1116 (N_1116,N_732,N_903);
nand U1117 (N_1117,N_504,N_628);
nand U1118 (N_1118,N_968,N_639);
nand U1119 (N_1119,N_692,N_678);
and U1120 (N_1120,N_837,N_893);
nor U1121 (N_1121,N_542,N_540);
xnor U1122 (N_1122,N_618,N_873);
and U1123 (N_1123,N_500,N_748);
nand U1124 (N_1124,N_896,N_611);
nand U1125 (N_1125,N_566,N_820);
and U1126 (N_1126,N_778,N_807);
nand U1127 (N_1127,N_823,N_972);
and U1128 (N_1128,N_959,N_844);
and U1129 (N_1129,N_541,N_556);
and U1130 (N_1130,N_595,N_782);
or U1131 (N_1131,N_558,N_751);
and U1132 (N_1132,N_708,N_554);
nand U1133 (N_1133,N_752,N_758);
and U1134 (N_1134,N_696,N_623);
nor U1135 (N_1135,N_739,N_805);
nand U1136 (N_1136,N_926,N_906);
or U1137 (N_1137,N_936,N_982);
and U1138 (N_1138,N_777,N_599);
or U1139 (N_1139,N_706,N_591);
or U1140 (N_1140,N_517,N_961);
nor U1141 (N_1141,N_813,N_603);
or U1142 (N_1142,N_933,N_964);
nand U1143 (N_1143,N_950,N_503);
or U1144 (N_1144,N_609,N_773);
nand U1145 (N_1145,N_733,N_677);
nor U1146 (N_1146,N_923,N_897);
nand U1147 (N_1147,N_736,N_929);
and U1148 (N_1148,N_649,N_868);
nor U1149 (N_1149,N_808,N_512);
nor U1150 (N_1150,N_818,N_569);
and U1151 (N_1151,N_976,N_744);
nand U1152 (N_1152,N_685,N_755);
and U1153 (N_1153,N_661,N_507);
nor U1154 (N_1154,N_842,N_637);
or U1155 (N_1155,N_879,N_718);
nand U1156 (N_1156,N_719,N_947);
nand U1157 (N_1157,N_791,N_872);
and U1158 (N_1158,N_655,N_992);
nor U1159 (N_1159,N_776,N_996);
nor U1160 (N_1160,N_796,N_511);
or U1161 (N_1161,N_743,N_576);
nand U1162 (N_1162,N_675,N_821);
nor U1163 (N_1163,N_565,N_553);
or U1164 (N_1164,N_790,N_787);
and U1165 (N_1165,N_767,N_698);
and U1166 (N_1166,N_916,N_622);
nor U1167 (N_1167,N_580,N_709);
nor U1168 (N_1168,N_590,N_693);
nand U1169 (N_1169,N_571,N_720);
nand U1170 (N_1170,N_705,N_985);
or U1171 (N_1171,N_988,N_727);
or U1172 (N_1172,N_822,N_514);
nor U1173 (N_1173,N_508,N_584);
nand U1174 (N_1174,N_997,N_779);
and U1175 (N_1175,N_657,N_561);
or U1176 (N_1176,N_722,N_886);
or U1177 (N_1177,N_803,N_895);
or U1178 (N_1178,N_606,N_759);
and U1179 (N_1179,N_522,N_883);
and U1180 (N_1180,N_954,N_768);
nor U1181 (N_1181,N_546,N_754);
nor U1182 (N_1182,N_917,N_593);
nor U1183 (N_1183,N_635,N_683);
and U1184 (N_1184,N_728,N_887);
nor U1185 (N_1185,N_532,N_607);
and U1186 (N_1186,N_800,N_991);
nor U1187 (N_1187,N_824,N_518);
or U1188 (N_1188,N_802,N_774);
nand U1189 (N_1189,N_555,N_826);
nand U1190 (N_1190,N_764,N_741);
or U1191 (N_1191,N_891,N_911);
and U1192 (N_1192,N_977,N_894);
and U1193 (N_1193,N_882,N_691);
and U1194 (N_1194,N_831,N_769);
or U1195 (N_1195,N_585,N_676);
nor U1196 (N_1196,N_941,N_864);
nand U1197 (N_1197,N_931,N_681);
and U1198 (N_1198,N_979,N_568);
or U1199 (N_1199,N_785,N_588);
nor U1200 (N_1200,N_563,N_711);
nor U1201 (N_1201,N_710,N_721);
and U1202 (N_1202,N_598,N_899);
and U1203 (N_1203,N_890,N_702);
or U1204 (N_1204,N_847,N_857);
or U1205 (N_1205,N_613,N_898);
or U1206 (N_1206,N_666,N_725);
nand U1207 (N_1207,N_970,N_957);
and U1208 (N_1208,N_701,N_737);
nand U1209 (N_1209,N_597,N_827);
nand U1210 (N_1210,N_738,N_860);
or U1211 (N_1211,N_594,N_684);
nand U1212 (N_1212,N_909,N_636);
nand U1213 (N_1213,N_829,N_845);
nand U1214 (N_1214,N_548,N_851);
and U1215 (N_1215,N_966,N_905);
and U1216 (N_1216,N_640,N_672);
or U1217 (N_1217,N_527,N_772);
or U1218 (N_1218,N_799,N_783);
nand U1219 (N_1219,N_881,N_506);
or U1220 (N_1220,N_745,N_578);
nor U1221 (N_1221,N_679,N_810);
and U1222 (N_1222,N_528,N_775);
or U1223 (N_1223,N_876,N_700);
or U1224 (N_1224,N_629,N_771);
nor U1225 (N_1225,N_834,N_938);
and U1226 (N_1226,N_757,N_980);
nand U1227 (N_1227,N_625,N_920);
nand U1228 (N_1228,N_900,N_674);
nand U1229 (N_1229,N_835,N_510);
or U1230 (N_1230,N_990,N_602);
nor U1231 (N_1231,N_526,N_608);
or U1232 (N_1232,N_534,N_619);
nor U1233 (N_1233,N_697,N_878);
xnor U1234 (N_1234,N_690,N_729);
or U1235 (N_1235,N_884,N_513);
and U1236 (N_1236,N_604,N_967);
or U1237 (N_1237,N_682,N_583);
nor U1238 (N_1238,N_862,N_652);
and U1239 (N_1239,N_645,N_574);
nor U1240 (N_1240,N_910,N_577);
or U1241 (N_1241,N_614,N_962);
and U1242 (N_1242,N_746,N_830);
and U1243 (N_1243,N_570,N_919);
and U1244 (N_1244,N_975,N_747);
nand U1245 (N_1245,N_621,N_524);
or U1246 (N_1246,N_780,N_809);
nor U1247 (N_1247,N_880,N_832);
nor U1248 (N_1248,N_735,N_680);
nor U1249 (N_1249,N_989,N_981);
nor U1250 (N_1250,N_691,N_587);
or U1251 (N_1251,N_666,N_546);
and U1252 (N_1252,N_999,N_693);
nand U1253 (N_1253,N_937,N_604);
nand U1254 (N_1254,N_951,N_874);
nor U1255 (N_1255,N_546,N_564);
and U1256 (N_1256,N_884,N_719);
and U1257 (N_1257,N_632,N_989);
nor U1258 (N_1258,N_638,N_914);
or U1259 (N_1259,N_711,N_512);
xor U1260 (N_1260,N_756,N_672);
or U1261 (N_1261,N_806,N_902);
and U1262 (N_1262,N_884,N_839);
and U1263 (N_1263,N_828,N_641);
nor U1264 (N_1264,N_735,N_536);
and U1265 (N_1265,N_892,N_786);
or U1266 (N_1266,N_818,N_808);
nor U1267 (N_1267,N_741,N_811);
or U1268 (N_1268,N_994,N_861);
and U1269 (N_1269,N_757,N_534);
nor U1270 (N_1270,N_734,N_651);
or U1271 (N_1271,N_739,N_773);
or U1272 (N_1272,N_951,N_532);
nand U1273 (N_1273,N_938,N_836);
nor U1274 (N_1274,N_594,N_955);
and U1275 (N_1275,N_853,N_528);
nor U1276 (N_1276,N_603,N_605);
nand U1277 (N_1277,N_779,N_736);
nand U1278 (N_1278,N_845,N_823);
nor U1279 (N_1279,N_945,N_989);
nor U1280 (N_1280,N_745,N_571);
nand U1281 (N_1281,N_901,N_715);
nor U1282 (N_1282,N_847,N_650);
or U1283 (N_1283,N_922,N_594);
nor U1284 (N_1284,N_607,N_979);
nand U1285 (N_1285,N_636,N_873);
nand U1286 (N_1286,N_864,N_844);
and U1287 (N_1287,N_992,N_882);
nand U1288 (N_1288,N_939,N_668);
and U1289 (N_1289,N_891,N_895);
nor U1290 (N_1290,N_943,N_801);
nor U1291 (N_1291,N_765,N_800);
or U1292 (N_1292,N_981,N_999);
nor U1293 (N_1293,N_595,N_662);
nor U1294 (N_1294,N_895,N_722);
or U1295 (N_1295,N_681,N_790);
and U1296 (N_1296,N_926,N_518);
nand U1297 (N_1297,N_989,N_851);
and U1298 (N_1298,N_714,N_762);
nand U1299 (N_1299,N_815,N_553);
nor U1300 (N_1300,N_544,N_835);
nand U1301 (N_1301,N_676,N_787);
or U1302 (N_1302,N_556,N_641);
nor U1303 (N_1303,N_619,N_825);
and U1304 (N_1304,N_893,N_999);
nor U1305 (N_1305,N_816,N_615);
or U1306 (N_1306,N_904,N_846);
and U1307 (N_1307,N_991,N_702);
or U1308 (N_1308,N_528,N_659);
nand U1309 (N_1309,N_847,N_889);
nand U1310 (N_1310,N_986,N_851);
or U1311 (N_1311,N_527,N_969);
or U1312 (N_1312,N_734,N_549);
or U1313 (N_1313,N_908,N_668);
and U1314 (N_1314,N_681,N_531);
and U1315 (N_1315,N_879,N_731);
or U1316 (N_1316,N_883,N_659);
or U1317 (N_1317,N_980,N_951);
nand U1318 (N_1318,N_554,N_682);
nand U1319 (N_1319,N_500,N_567);
nand U1320 (N_1320,N_743,N_726);
nand U1321 (N_1321,N_651,N_904);
nor U1322 (N_1322,N_588,N_817);
or U1323 (N_1323,N_720,N_916);
nor U1324 (N_1324,N_738,N_701);
nor U1325 (N_1325,N_535,N_857);
nor U1326 (N_1326,N_736,N_764);
nand U1327 (N_1327,N_768,N_537);
or U1328 (N_1328,N_704,N_841);
nor U1329 (N_1329,N_771,N_878);
or U1330 (N_1330,N_979,N_906);
and U1331 (N_1331,N_699,N_663);
or U1332 (N_1332,N_560,N_622);
nor U1333 (N_1333,N_739,N_885);
and U1334 (N_1334,N_508,N_738);
nor U1335 (N_1335,N_699,N_743);
or U1336 (N_1336,N_938,N_868);
nor U1337 (N_1337,N_731,N_918);
xor U1338 (N_1338,N_717,N_979);
nor U1339 (N_1339,N_577,N_869);
nor U1340 (N_1340,N_618,N_796);
or U1341 (N_1341,N_880,N_752);
and U1342 (N_1342,N_808,N_903);
and U1343 (N_1343,N_680,N_616);
and U1344 (N_1344,N_861,N_869);
or U1345 (N_1345,N_719,N_999);
or U1346 (N_1346,N_734,N_566);
nand U1347 (N_1347,N_988,N_782);
nor U1348 (N_1348,N_616,N_911);
nor U1349 (N_1349,N_946,N_980);
nor U1350 (N_1350,N_978,N_683);
or U1351 (N_1351,N_578,N_887);
nand U1352 (N_1352,N_546,N_662);
nand U1353 (N_1353,N_932,N_992);
and U1354 (N_1354,N_638,N_560);
or U1355 (N_1355,N_912,N_527);
nand U1356 (N_1356,N_709,N_918);
nor U1357 (N_1357,N_549,N_502);
or U1358 (N_1358,N_656,N_761);
or U1359 (N_1359,N_993,N_697);
nor U1360 (N_1360,N_733,N_846);
or U1361 (N_1361,N_881,N_599);
nand U1362 (N_1362,N_653,N_786);
nor U1363 (N_1363,N_545,N_897);
or U1364 (N_1364,N_745,N_562);
and U1365 (N_1365,N_786,N_640);
and U1366 (N_1366,N_867,N_895);
nor U1367 (N_1367,N_850,N_721);
nor U1368 (N_1368,N_509,N_646);
nor U1369 (N_1369,N_923,N_857);
nor U1370 (N_1370,N_871,N_872);
nand U1371 (N_1371,N_536,N_909);
or U1372 (N_1372,N_709,N_800);
nand U1373 (N_1373,N_706,N_821);
or U1374 (N_1374,N_795,N_807);
or U1375 (N_1375,N_537,N_715);
and U1376 (N_1376,N_651,N_500);
or U1377 (N_1377,N_993,N_507);
and U1378 (N_1378,N_946,N_632);
nand U1379 (N_1379,N_773,N_987);
nand U1380 (N_1380,N_817,N_740);
and U1381 (N_1381,N_851,N_642);
nor U1382 (N_1382,N_792,N_991);
nand U1383 (N_1383,N_702,N_942);
or U1384 (N_1384,N_909,N_731);
nand U1385 (N_1385,N_843,N_536);
nand U1386 (N_1386,N_532,N_790);
nor U1387 (N_1387,N_770,N_951);
and U1388 (N_1388,N_976,N_861);
or U1389 (N_1389,N_767,N_869);
and U1390 (N_1390,N_501,N_626);
and U1391 (N_1391,N_521,N_691);
nor U1392 (N_1392,N_851,N_691);
or U1393 (N_1393,N_619,N_704);
nand U1394 (N_1394,N_824,N_744);
nand U1395 (N_1395,N_892,N_574);
or U1396 (N_1396,N_891,N_552);
and U1397 (N_1397,N_717,N_930);
nor U1398 (N_1398,N_818,N_706);
and U1399 (N_1399,N_572,N_903);
nor U1400 (N_1400,N_981,N_632);
or U1401 (N_1401,N_536,N_687);
nand U1402 (N_1402,N_697,N_739);
or U1403 (N_1403,N_969,N_954);
nor U1404 (N_1404,N_650,N_761);
nand U1405 (N_1405,N_532,N_784);
and U1406 (N_1406,N_850,N_993);
and U1407 (N_1407,N_913,N_829);
and U1408 (N_1408,N_963,N_510);
nor U1409 (N_1409,N_587,N_947);
nand U1410 (N_1410,N_658,N_769);
and U1411 (N_1411,N_596,N_512);
nand U1412 (N_1412,N_688,N_547);
nor U1413 (N_1413,N_786,N_789);
or U1414 (N_1414,N_785,N_866);
or U1415 (N_1415,N_846,N_985);
and U1416 (N_1416,N_525,N_690);
nor U1417 (N_1417,N_860,N_693);
nand U1418 (N_1418,N_905,N_931);
and U1419 (N_1419,N_606,N_608);
or U1420 (N_1420,N_731,N_632);
or U1421 (N_1421,N_981,N_539);
nor U1422 (N_1422,N_768,N_680);
and U1423 (N_1423,N_723,N_807);
nand U1424 (N_1424,N_647,N_786);
and U1425 (N_1425,N_642,N_827);
nor U1426 (N_1426,N_759,N_669);
or U1427 (N_1427,N_795,N_820);
nor U1428 (N_1428,N_893,N_730);
nand U1429 (N_1429,N_689,N_504);
or U1430 (N_1430,N_658,N_768);
and U1431 (N_1431,N_575,N_683);
nor U1432 (N_1432,N_639,N_862);
nor U1433 (N_1433,N_596,N_953);
nor U1434 (N_1434,N_551,N_954);
or U1435 (N_1435,N_629,N_829);
or U1436 (N_1436,N_612,N_611);
or U1437 (N_1437,N_649,N_874);
or U1438 (N_1438,N_989,N_842);
nand U1439 (N_1439,N_546,N_944);
and U1440 (N_1440,N_739,N_681);
or U1441 (N_1441,N_907,N_634);
nand U1442 (N_1442,N_974,N_618);
nand U1443 (N_1443,N_811,N_746);
nor U1444 (N_1444,N_744,N_860);
or U1445 (N_1445,N_677,N_929);
or U1446 (N_1446,N_800,N_823);
nor U1447 (N_1447,N_936,N_675);
or U1448 (N_1448,N_586,N_869);
nor U1449 (N_1449,N_700,N_832);
nand U1450 (N_1450,N_532,N_689);
or U1451 (N_1451,N_648,N_963);
and U1452 (N_1452,N_909,N_793);
or U1453 (N_1453,N_670,N_824);
and U1454 (N_1454,N_960,N_885);
and U1455 (N_1455,N_765,N_733);
nand U1456 (N_1456,N_668,N_938);
and U1457 (N_1457,N_830,N_692);
or U1458 (N_1458,N_896,N_683);
nor U1459 (N_1459,N_607,N_847);
nor U1460 (N_1460,N_938,N_654);
nor U1461 (N_1461,N_720,N_817);
and U1462 (N_1462,N_894,N_792);
nand U1463 (N_1463,N_833,N_945);
nand U1464 (N_1464,N_550,N_924);
nand U1465 (N_1465,N_637,N_764);
nand U1466 (N_1466,N_628,N_649);
nor U1467 (N_1467,N_611,N_763);
nand U1468 (N_1468,N_968,N_755);
nor U1469 (N_1469,N_654,N_681);
or U1470 (N_1470,N_830,N_924);
nand U1471 (N_1471,N_726,N_530);
nor U1472 (N_1472,N_695,N_648);
or U1473 (N_1473,N_906,N_809);
or U1474 (N_1474,N_613,N_806);
and U1475 (N_1475,N_547,N_917);
nor U1476 (N_1476,N_903,N_692);
and U1477 (N_1477,N_875,N_898);
nor U1478 (N_1478,N_735,N_514);
xnor U1479 (N_1479,N_915,N_630);
nand U1480 (N_1480,N_939,N_653);
and U1481 (N_1481,N_819,N_540);
and U1482 (N_1482,N_520,N_746);
nand U1483 (N_1483,N_842,N_531);
and U1484 (N_1484,N_683,N_745);
nand U1485 (N_1485,N_953,N_839);
and U1486 (N_1486,N_658,N_915);
nand U1487 (N_1487,N_775,N_568);
nand U1488 (N_1488,N_708,N_503);
nand U1489 (N_1489,N_672,N_566);
nand U1490 (N_1490,N_854,N_846);
nor U1491 (N_1491,N_725,N_964);
and U1492 (N_1492,N_629,N_692);
and U1493 (N_1493,N_843,N_668);
or U1494 (N_1494,N_582,N_906);
nor U1495 (N_1495,N_847,N_843);
and U1496 (N_1496,N_688,N_573);
xor U1497 (N_1497,N_680,N_634);
and U1498 (N_1498,N_677,N_856);
or U1499 (N_1499,N_624,N_933);
nor U1500 (N_1500,N_1375,N_1044);
or U1501 (N_1501,N_1015,N_1325);
or U1502 (N_1502,N_1076,N_1132);
and U1503 (N_1503,N_1465,N_1408);
nor U1504 (N_1504,N_1226,N_1394);
or U1505 (N_1505,N_1298,N_1324);
nor U1506 (N_1506,N_1316,N_1145);
nor U1507 (N_1507,N_1405,N_1430);
or U1508 (N_1508,N_1191,N_1498);
nand U1509 (N_1509,N_1342,N_1002);
nor U1510 (N_1510,N_1222,N_1173);
nor U1511 (N_1511,N_1120,N_1403);
or U1512 (N_1512,N_1140,N_1420);
nand U1513 (N_1513,N_1041,N_1082);
nor U1514 (N_1514,N_1409,N_1292);
nor U1515 (N_1515,N_1458,N_1205);
and U1516 (N_1516,N_1242,N_1429);
nor U1517 (N_1517,N_1037,N_1443);
nor U1518 (N_1518,N_1457,N_1167);
and U1519 (N_1519,N_1014,N_1255);
nor U1520 (N_1520,N_1163,N_1105);
nor U1521 (N_1521,N_1006,N_1404);
nand U1522 (N_1522,N_1371,N_1490);
and U1523 (N_1523,N_1344,N_1437);
or U1524 (N_1524,N_1389,N_1146);
nand U1525 (N_1525,N_1338,N_1266);
nor U1526 (N_1526,N_1286,N_1483);
or U1527 (N_1527,N_1354,N_1312);
and U1528 (N_1528,N_1350,N_1060);
or U1529 (N_1529,N_1313,N_1072);
or U1530 (N_1530,N_1155,N_1412);
nand U1531 (N_1531,N_1017,N_1165);
or U1532 (N_1532,N_1449,N_1094);
nand U1533 (N_1533,N_1080,N_1178);
and U1534 (N_1534,N_1129,N_1306);
nor U1535 (N_1535,N_1198,N_1398);
or U1536 (N_1536,N_1453,N_1307);
nor U1537 (N_1537,N_1265,N_1168);
nand U1538 (N_1538,N_1439,N_1180);
nor U1539 (N_1539,N_1194,N_1023);
nand U1540 (N_1540,N_1235,N_1141);
nor U1541 (N_1541,N_1393,N_1410);
nand U1542 (N_1542,N_1374,N_1133);
or U1543 (N_1543,N_1149,N_1181);
or U1544 (N_1544,N_1471,N_1013);
nor U1545 (N_1545,N_1033,N_1386);
and U1546 (N_1546,N_1110,N_1278);
nand U1547 (N_1547,N_1323,N_1030);
nand U1548 (N_1548,N_1209,N_1282);
nor U1549 (N_1549,N_1433,N_1000);
and U1550 (N_1550,N_1438,N_1124);
nor U1551 (N_1551,N_1474,N_1150);
and U1552 (N_1552,N_1010,N_1097);
nor U1553 (N_1553,N_1111,N_1213);
or U1554 (N_1554,N_1179,N_1311);
or U1555 (N_1555,N_1204,N_1134);
nor U1556 (N_1556,N_1159,N_1304);
nand U1557 (N_1557,N_1492,N_1053);
nor U1558 (N_1558,N_1416,N_1388);
and U1559 (N_1559,N_1096,N_1031);
nand U1560 (N_1560,N_1079,N_1480);
or U1561 (N_1561,N_1363,N_1005);
nand U1562 (N_1562,N_1297,N_1123);
or U1563 (N_1563,N_1333,N_1143);
or U1564 (N_1564,N_1425,N_1249);
nand U1565 (N_1565,N_1225,N_1463);
nor U1566 (N_1566,N_1075,N_1296);
or U1567 (N_1567,N_1455,N_1218);
nand U1568 (N_1568,N_1026,N_1478);
nand U1569 (N_1569,N_1305,N_1277);
nor U1570 (N_1570,N_1216,N_1007);
or U1571 (N_1571,N_1495,N_1435);
nor U1572 (N_1572,N_1067,N_1185);
xor U1573 (N_1573,N_1318,N_1239);
and U1574 (N_1574,N_1035,N_1351);
nand U1575 (N_1575,N_1361,N_1252);
or U1576 (N_1576,N_1320,N_1059);
nand U1577 (N_1577,N_1004,N_1308);
nor U1578 (N_1578,N_1202,N_1248);
nand U1579 (N_1579,N_1104,N_1217);
or U1580 (N_1580,N_1291,N_1415);
and U1581 (N_1581,N_1088,N_1024);
nor U1582 (N_1582,N_1263,N_1419);
nand U1583 (N_1583,N_1112,N_1244);
or U1584 (N_1584,N_1171,N_1040);
and U1585 (N_1585,N_1328,N_1074);
and U1586 (N_1586,N_1379,N_1175);
or U1587 (N_1587,N_1290,N_1161);
nand U1588 (N_1588,N_1245,N_1347);
nand U1589 (N_1589,N_1227,N_1211);
or U1590 (N_1590,N_1025,N_1481);
or U1591 (N_1591,N_1220,N_1269);
or U1592 (N_1592,N_1052,N_1329);
or U1593 (N_1593,N_1012,N_1496);
nor U1594 (N_1594,N_1116,N_1195);
nor U1595 (N_1595,N_1479,N_1261);
nor U1596 (N_1596,N_1034,N_1341);
nand U1597 (N_1597,N_1396,N_1190);
or U1598 (N_1598,N_1369,N_1048);
nor U1599 (N_1599,N_1151,N_1270);
nor U1600 (N_1600,N_1203,N_1135);
and U1601 (N_1601,N_1285,N_1106);
nor U1602 (N_1602,N_1071,N_1456);
and U1603 (N_1603,N_1497,N_1421);
nand U1604 (N_1604,N_1336,N_1130);
nor U1605 (N_1605,N_1322,N_1138);
or U1606 (N_1606,N_1339,N_1381);
or U1607 (N_1607,N_1314,N_1493);
nand U1608 (N_1608,N_1170,N_1128);
and U1609 (N_1609,N_1289,N_1118);
and U1610 (N_1610,N_1207,N_1064);
or U1611 (N_1611,N_1377,N_1272);
or U1612 (N_1612,N_1090,N_1224);
or U1613 (N_1613,N_1029,N_1114);
or U1614 (N_1614,N_1450,N_1357);
nand U1615 (N_1615,N_1022,N_1231);
nor U1616 (N_1616,N_1233,N_1462);
or U1617 (N_1617,N_1020,N_1230);
nand U1618 (N_1618,N_1319,N_1414);
or U1619 (N_1619,N_1295,N_1160);
nand U1620 (N_1620,N_1491,N_1056);
and U1621 (N_1621,N_1137,N_1147);
nand U1622 (N_1622,N_1008,N_1027);
nor U1623 (N_1623,N_1383,N_1085);
xor U1624 (N_1624,N_1432,N_1426);
nand U1625 (N_1625,N_1434,N_1201);
nand U1626 (N_1626,N_1069,N_1424);
and U1627 (N_1627,N_1452,N_1436);
and U1628 (N_1628,N_1055,N_1358);
or U1629 (N_1629,N_1395,N_1062);
or U1630 (N_1630,N_1018,N_1407);
and U1631 (N_1631,N_1045,N_1247);
nand U1632 (N_1632,N_1142,N_1061);
nand U1633 (N_1633,N_1353,N_1442);
nor U1634 (N_1634,N_1193,N_1302);
nand U1635 (N_1635,N_1460,N_1042);
nand U1636 (N_1636,N_1065,N_1127);
nor U1637 (N_1637,N_1073,N_1273);
or U1638 (N_1638,N_1340,N_1221);
and U1639 (N_1639,N_1356,N_1232);
and U1640 (N_1640,N_1084,N_1258);
nand U1641 (N_1641,N_1210,N_1335);
or U1642 (N_1642,N_1139,N_1310);
xnor U1643 (N_1643,N_1337,N_1229);
or U1644 (N_1644,N_1259,N_1468);
nand U1645 (N_1645,N_1077,N_1189);
nand U1646 (N_1646,N_1066,N_1387);
nand U1647 (N_1647,N_1472,N_1078);
nor U1648 (N_1648,N_1153,N_1199);
or U1649 (N_1649,N_1240,N_1267);
and U1650 (N_1650,N_1122,N_1422);
nand U1651 (N_1651,N_1003,N_1376);
nand U1652 (N_1652,N_1051,N_1241);
and U1653 (N_1653,N_1016,N_1043);
or U1654 (N_1654,N_1345,N_1098);
and U1655 (N_1655,N_1367,N_1299);
and U1656 (N_1656,N_1115,N_1152);
and U1657 (N_1657,N_1162,N_1406);
nand U1658 (N_1658,N_1476,N_1390);
and U1659 (N_1659,N_1107,N_1081);
nand U1660 (N_1660,N_1215,N_1136);
or U1661 (N_1661,N_1011,N_1373);
and U1662 (N_1662,N_1251,N_1184);
nand U1663 (N_1663,N_1359,N_1268);
or U1664 (N_1664,N_1121,N_1169);
or U1665 (N_1665,N_1378,N_1236);
nor U1666 (N_1666,N_1392,N_1117);
and U1667 (N_1667,N_1413,N_1482);
nand U1668 (N_1668,N_1362,N_1206);
and U1669 (N_1669,N_1448,N_1102);
nand U1670 (N_1670,N_1253,N_1469);
and U1671 (N_1671,N_1046,N_1164);
nand U1672 (N_1672,N_1315,N_1070);
and U1673 (N_1673,N_1257,N_1228);
nor U1674 (N_1674,N_1208,N_1036);
nor U1675 (N_1675,N_1327,N_1086);
nand U1676 (N_1676,N_1275,N_1279);
nand U1677 (N_1677,N_1431,N_1461);
or U1678 (N_1678,N_1038,N_1473);
and U1679 (N_1679,N_1246,N_1451);
nor U1680 (N_1680,N_1192,N_1303);
and U1681 (N_1681,N_1126,N_1467);
nor U1682 (N_1682,N_1197,N_1428);
or U1683 (N_1683,N_1317,N_1447);
nor U1684 (N_1684,N_1214,N_1166);
and U1685 (N_1685,N_1243,N_1050);
or U1686 (N_1686,N_1196,N_1028);
or U1687 (N_1687,N_1083,N_1177);
or U1688 (N_1688,N_1459,N_1119);
nand U1689 (N_1689,N_1058,N_1254);
and U1690 (N_1690,N_1274,N_1186);
nor U1691 (N_1691,N_1212,N_1262);
nand U1692 (N_1692,N_1009,N_1125);
and U1693 (N_1693,N_1049,N_1444);
nand U1694 (N_1694,N_1219,N_1454);
or U1695 (N_1695,N_1399,N_1301);
nand U1696 (N_1696,N_1370,N_1099);
and U1697 (N_1697,N_1402,N_1188);
or U1698 (N_1698,N_1223,N_1200);
nand U1699 (N_1699,N_1032,N_1384);
nand U1700 (N_1700,N_1087,N_1054);
or U1701 (N_1701,N_1488,N_1427);
nor U1702 (N_1702,N_1047,N_1464);
nor U1703 (N_1703,N_1348,N_1256);
or U1704 (N_1704,N_1237,N_1187);
nor U1705 (N_1705,N_1440,N_1144);
nand U1706 (N_1706,N_1182,N_1401);
nor U1707 (N_1707,N_1331,N_1176);
and U1708 (N_1708,N_1093,N_1103);
nor U1709 (N_1709,N_1109,N_1466);
nand U1710 (N_1710,N_1294,N_1486);
and U1711 (N_1711,N_1131,N_1108);
and U1712 (N_1712,N_1039,N_1234);
nand U1713 (N_1713,N_1485,N_1293);
nand U1714 (N_1714,N_1100,N_1156);
and U1715 (N_1715,N_1321,N_1068);
or U1716 (N_1716,N_1417,N_1489);
nor U1717 (N_1717,N_1397,N_1021);
or U1718 (N_1718,N_1280,N_1380);
and U1719 (N_1719,N_1355,N_1264);
nor U1720 (N_1720,N_1499,N_1346);
and U1721 (N_1721,N_1271,N_1154);
nor U1722 (N_1722,N_1283,N_1368);
nor U1723 (N_1723,N_1364,N_1366);
or U1724 (N_1724,N_1091,N_1360);
or U1725 (N_1725,N_1284,N_1475);
nand U1726 (N_1726,N_1157,N_1330);
nand U1727 (N_1727,N_1238,N_1372);
nor U1728 (N_1728,N_1365,N_1477);
nand U1729 (N_1729,N_1309,N_1276);
or U1730 (N_1730,N_1352,N_1300);
nand U1731 (N_1731,N_1418,N_1349);
nand U1732 (N_1732,N_1287,N_1445);
and U1733 (N_1733,N_1423,N_1001);
or U1734 (N_1734,N_1148,N_1281);
and U1735 (N_1735,N_1174,N_1441);
or U1736 (N_1736,N_1089,N_1332);
and U1737 (N_1737,N_1382,N_1385);
nand U1738 (N_1738,N_1334,N_1057);
or U1739 (N_1739,N_1092,N_1470);
nand U1740 (N_1740,N_1158,N_1343);
or U1741 (N_1741,N_1400,N_1095);
nor U1742 (N_1742,N_1411,N_1391);
nand U1743 (N_1743,N_1113,N_1183);
nor U1744 (N_1744,N_1101,N_1494);
nor U1745 (N_1745,N_1484,N_1326);
and U1746 (N_1746,N_1250,N_1288);
nand U1747 (N_1747,N_1172,N_1019);
nand U1748 (N_1748,N_1260,N_1487);
nand U1749 (N_1749,N_1063,N_1446);
or U1750 (N_1750,N_1077,N_1224);
or U1751 (N_1751,N_1377,N_1040);
and U1752 (N_1752,N_1166,N_1152);
and U1753 (N_1753,N_1098,N_1323);
nor U1754 (N_1754,N_1179,N_1106);
nand U1755 (N_1755,N_1061,N_1028);
nor U1756 (N_1756,N_1493,N_1110);
nand U1757 (N_1757,N_1051,N_1182);
and U1758 (N_1758,N_1439,N_1373);
nand U1759 (N_1759,N_1253,N_1036);
and U1760 (N_1760,N_1249,N_1494);
and U1761 (N_1761,N_1439,N_1476);
nand U1762 (N_1762,N_1031,N_1063);
or U1763 (N_1763,N_1425,N_1374);
nand U1764 (N_1764,N_1195,N_1229);
nand U1765 (N_1765,N_1181,N_1333);
or U1766 (N_1766,N_1040,N_1251);
nand U1767 (N_1767,N_1443,N_1432);
or U1768 (N_1768,N_1153,N_1077);
and U1769 (N_1769,N_1391,N_1479);
and U1770 (N_1770,N_1025,N_1491);
or U1771 (N_1771,N_1289,N_1310);
and U1772 (N_1772,N_1499,N_1063);
nor U1773 (N_1773,N_1368,N_1294);
nand U1774 (N_1774,N_1107,N_1346);
nand U1775 (N_1775,N_1217,N_1376);
nor U1776 (N_1776,N_1040,N_1243);
or U1777 (N_1777,N_1126,N_1408);
or U1778 (N_1778,N_1195,N_1101);
or U1779 (N_1779,N_1109,N_1486);
nor U1780 (N_1780,N_1345,N_1216);
or U1781 (N_1781,N_1447,N_1389);
or U1782 (N_1782,N_1244,N_1249);
and U1783 (N_1783,N_1096,N_1019);
and U1784 (N_1784,N_1283,N_1073);
or U1785 (N_1785,N_1189,N_1062);
or U1786 (N_1786,N_1166,N_1315);
and U1787 (N_1787,N_1131,N_1301);
nand U1788 (N_1788,N_1378,N_1114);
or U1789 (N_1789,N_1477,N_1467);
nand U1790 (N_1790,N_1493,N_1006);
and U1791 (N_1791,N_1490,N_1296);
and U1792 (N_1792,N_1026,N_1072);
and U1793 (N_1793,N_1222,N_1398);
and U1794 (N_1794,N_1361,N_1155);
nor U1795 (N_1795,N_1258,N_1331);
and U1796 (N_1796,N_1301,N_1431);
nor U1797 (N_1797,N_1213,N_1083);
and U1798 (N_1798,N_1162,N_1344);
xnor U1799 (N_1799,N_1311,N_1093);
or U1800 (N_1800,N_1338,N_1231);
and U1801 (N_1801,N_1208,N_1087);
and U1802 (N_1802,N_1202,N_1134);
nor U1803 (N_1803,N_1172,N_1016);
and U1804 (N_1804,N_1396,N_1048);
or U1805 (N_1805,N_1363,N_1134);
nand U1806 (N_1806,N_1254,N_1250);
and U1807 (N_1807,N_1298,N_1102);
nand U1808 (N_1808,N_1322,N_1010);
or U1809 (N_1809,N_1254,N_1233);
and U1810 (N_1810,N_1299,N_1429);
or U1811 (N_1811,N_1305,N_1190);
and U1812 (N_1812,N_1131,N_1064);
or U1813 (N_1813,N_1139,N_1331);
nor U1814 (N_1814,N_1063,N_1247);
or U1815 (N_1815,N_1312,N_1255);
nand U1816 (N_1816,N_1018,N_1438);
nand U1817 (N_1817,N_1169,N_1136);
nor U1818 (N_1818,N_1258,N_1016);
nor U1819 (N_1819,N_1311,N_1374);
and U1820 (N_1820,N_1095,N_1029);
nor U1821 (N_1821,N_1404,N_1414);
or U1822 (N_1822,N_1321,N_1251);
nand U1823 (N_1823,N_1494,N_1187);
or U1824 (N_1824,N_1427,N_1013);
nand U1825 (N_1825,N_1182,N_1018);
nor U1826 (N_1826,N_1456,N_1412);
or U1827 (N_1827,N_1436,N_1349);
nor U1828 (N_1828,N_1379,N_1085);
nand U1829 (N_1829,N_1149,N_1462);
and U1830 (N_1830,N_1034,N_1143);
nor U1831 (N_1831,N_1243,N_1483);
nor U1832 (N_1832,N_1240,N_1401);
or U1833 (N_1833,N_1066,N_1368);
nand U1834 (N_1834,N_1203,N_1037);
nor U1835 (N_1835,N_1194,N_1054);
nor U1836 (N_1836,N_1245,N_1498);
and U1837 (N_1837,N_1305,N_1129);
nand U1838 (N_1838,N_1424,N_1362);
nand U1839 (N_1839,N_1286,N_1447);
and U1840 (N_1840,N_1049,N_1056);
nor U1841 (N_1841,N_1302,N_1407);
or U1842 (N_1842,N_1414,N_1182);
or U1843 (N_1843,N_1358,N_1234);
nand U1844 (N_1844,N_1173,N_1303);
nor U1845 (N_1845,N_1100,N_1231);
nand U1846 (N_1846,N_1390,N_1203);
and U1847 (N_1847,N_1333,N_1350);
or U1848 (N_1848,N_1311,N_1292);
nand U1849 (N_1849,N_1103,N_1011);
or U1850 (N_1850,N_1380,N_1067);
or U1851 (N_1851,N_1385,N_1483);
or U1852 (N_1852,N_1049,N_1189);
and U1853 (N_1853,N_1074,N_1198);
nand U1854 (N_1854,N_1085,N_1481);
nor U1855 (N_1855,N_1403,N_1327);
nand U1856 (N_1856,N_1107,N_1343);
nor U1857 (N_1857,N_1257,N_1081);
nor U1858 (N_1858,N_1469,N_1227);
nor U1859 (N_1859,N_1415,N_1227);
nand U1860 (N_1860,N_1079,N_1418);
or U1861 (N_1861,N_1055,N_1336);
and U1862 (N_1862,N_1321,N_1179);
nand U1863 (N_1863,N_1262,N_1371);
and U1864 (N_1864,N_1236,N_1183);
or U1865 (N_1865,N_1329,N_1150);
or U1866 (N_1866,N_1464,N_1015);
and U1867 (N_1867,N_1378,N_1210);
nand U1868 (N_1868,N_1461,N_1213);
nor U1869 (N_1869,N_1393,N_1416);
or U1870 (N_1870,N_1051,N_1101);
nor U1871 (N_1871,N_1084,N_1110);
and U1872 (N_1872,N_1219,N_1128);
nand U1873 (N_1873,N_1081,N_1464);
or U1874 (N_1874,N_1279,N_1325);
nand U1875 (N_1875,N_1358,N_1081);
or U1876 (N_1876,N_1405,N_1129);
nor U1877 (N_1877,N_1051,N_1171);
and U1878 (N_1878,N_1387,N_1411);
nor U1879 (N_1879,N_1366,N_1457);
nor U1880 (N_1880,N_1454,N_1266);
or U1881 (N_1881,N_1061,N_1427);
nand U1882 (N_1882,N_1144,N_1316);
and U1883 (N_1883,N_1435,N_1380);
nand U1884 (N_1884,N_1220,N_1249);
xor U1885 (N_1885,N_1191,N_1448);
xor U1886 (N_1886,N_1179,N_1433);
and U1887 (N_1887,N_1401,N_1076);
nand U1888 (N_1888,N_1160,N_1492);
and U1889 (N_1889,N_1426,N_1171);
nand U1890 (N_1890,N_1006,N_1499);
nand U1891 (N_1891,N_1432,N_1182);
or U1892 (N_1892,N_1352,N_1225);
nor U1893 (N_1893,N_1443,N_1324);
or U1894 (N_1894,N_1028,N_1472);
nor U1895 (N_1895,N_1118,N_1294);
or U1896 (N_1896,N_1441,N_1490);
or U1897 (N_1897,N_1179,N_1450);
and U1898 (N_1898,N_1118,N_1447);
or U1899 (N_1899,N_1320,N_1469);
nor U1900 (N_1900,N_1194,N_1001);
or U1901 (N_1901,N_1280,N_1447);
nand U1902 (N_1902,N_1302,N_1366);
nor U1903 (N_1903,N_1222,N_1203);
and U1904 (N_1904,N_1349,N_1355);
and U1905 (N_1905,N_1341,N_1253);
nor U1906 (N_1906,N_1415,N_1230);
nor U1907 (N_1907,N_1396,N_1215);
or U1908 (N_1908,N_1033,N_1486);
or U1909 (N_1909,N_1041,N_1473);
nor U1910 (N_1910,N_1476,N_1255);
nor U1911 (N_1911,N_1273,N_1350);
and U1912 (N_1912,N_1273,N_1266);
nor U1913 (N_1913,N_1159,N_1107);
or U1914 (N_1914,N_1287,N_1043);
nand U1915 (N_1915,N_1049,N_1485);
nand U1916 (N_1916,N_1335,N_1404);
nor U1917 (N_1917,N_1491,N_1173);
nand U1918 (N_1918,N_1264,N_1434);
nand U1919 (N_1919,N_1363,N_1131);
or U1920 (N_1920,N_1387,N_1226);
and U1921 (N_1921,N_1066,N_1139);
nor U1922 (N_1922,N_1267,N_1010);
nor U1923 (N_1923,N_1218,N_1284);
nor U1924 (N_1924,N_1214,N_1346);
nand U1925 (N_1925,N_1308,N_1241);
and U1926 (N_1926,N_1241,N_1401);
nand U1927 (N_1927,N_1369,N_1145);
nand U1928 (N_1928,N_1466,N_1431);
or U1929 (N_1929,N_1012,N_1104);
and U1930 (N_1930,N_1313,N_1076);
and U1931 (N_1931,N_1286,N_1147);
nor U1932 (N_1932,N_1333,N_1349);
and U1933 (N_1933,N_1274,N_1317);
or U1934 (N_1934,N_1123,N_1204);
nand U1935 (N_1935,N_1169,N_1328);
and U1936 (N_1936,N_1013,N_1022);
nor U1937 (N_1937,N_1205,N_1324);
and U1938 (N_1938,N_1116,N_1286);
and U1939 (N_1939,N_1323,N_1010);
or U1940 (N_1940,N_1495,N_1479);
and U1941 (N_1941,N_1483,N_1407);
and U1942 (N_1942,N_1225,N_1279);
and U1943 (N_1943,N_1399,N_1297);
nand U1944 (N_1944,N_1191,N_1307);
nor U1945 (N_1945,N_1064,N_1217);
nand U1946 (N_1946,N_1328,N_1253);
and U1947 (N_1947,N_1144,N_1220);
nand U1948 (N_1948,N_1007,N_1473);
nor U1949 (N_1949,N_1493,N_1234);
and U1950 (N_1950,N_1128,N_1022);
and U1951 (N_1951,N_1333,N_1452);
or U1952 (N_1952,N_1355,N_1302);
nor U1953 (N_1953,N_1457,N_1395);
and U1954 (N_1954,N_1032,N_1335);
and U1955 (N_1955,N_1386,N_1263);
or U1956 (N_1956,N_1191,N_1163);
or U1957 (N_1957,N_1164,N_1307);
and U1958 (N_1958,N_1042,N_1131);
or U1959 (N_1959,N_1044,N_1444);
and U1960 (N_1960,N_1210,N_1282);
and U1961 (N_1961,N_1410,N_1456);
nand U1962 (N_1962,N_1087,N_1466);
and U1963 (N_1963,N_1048,N_1374);
nor U1964 (N_1964,N_1314,N_1272);
and U1965 (N_1965,N_1067,N_1165);
and U1966 (N_1966,N_1437,N_1203);
nand U1967 (N_1967,N_1166,N_1177);
xor U1968 (N_1968,N_1310,N_1399);
nand U1969 (N_1969,N_1483,N_1484);
nand U1970 (N_1970,N_1212,N_1476);
or U1971 (N_1971,N_1039,N_1175);
or U1972 (N_1972,N_1380,N_1135);
and U1973 (N_1973,N_1346,N_1449);
nand U1974 (N_1974,N_1336,N_1086);
or U1975 (N_1975,N_1268,N_1311);
nor U1976 (N_1976,N_1334,N_1046);
or U1977 (N_1977,N_1208,N_1028);
nand U1978 (N_1978,N_1422,N_1044);
nor U1979 (N_1979,N_1122,N_1096);
or U1980 (N_1980,N_1467,N_1468);
nor U1981 (N_1981,N_1282,N_1305);
or U1982 (N_1982,N_1370,N_1278);
nor U1983 (N_1983,N_1237,N_1254);
nor U1984 (N_1984,N_1481,N_1447);
and U1985 (N_1985,N_1006,N_1254);
or U1986 (N_1986,N_1315,N_1418);
and U1987 (N_1987,N_1103,N_1361);
nand U1988 (N_1988,N_1296,N_1426);
or U1989 (N_1989,N_1308,N_1136);
or U1990 (N_1990,N_1324,N_1178);
or U1991 (N_1991,N_1106,N_1191);
nor U1992 (N_1992,N_1265,N_1157);
nor U1993 (N_1993,N_1199,N_1321);
and U1994 (N_1994,N_1104,N_1470);
nor U1995 (N_1995,N_1286,N_1471);
or U1996 (N_1996,N_1490,N_1410);
nand U1997 (N_1997,N_1051,N_1160);
or U1998 (N_1998,N_1349,N_1062);
and U1999 (N_1999,N_1449,N_1092);
nor U2000 (N_2000,N_1650,N_1710);
and U2001 (N_2001,N_1885,N_1584);
nand U2002 (N_2002,N_1819,N_1679);
nand U2003 (N_2003,N_1605,N_1896);
nor U2004 (N_2004,N_1730,N_1872);
or U2005 (N_2005,N_1835,N_1691);
and U2006 (N_2006,N_1845,N_1652);
nor U2007 (N_2007,N_1798,N_1911);
nand U2008 (N_2008,N_1856,N_1703);
nand U2009 (N_2009,N_1894,N_1723);
nand U2010 (N_2010,N_1604,N_1561);
nor U2011 (N_2011,N_1810,N_1744);
or U2012 (N_2012,N_1895,N_1899);
and U2013 (N_2013,N_1646,N_1775);
and U2014 (N_2014,N_1581,N_1992);
nor U2015 (N_2015,N_1824,N_1714);
nand U2016 (N_2016,N_1715,N_1544);
and U2017 (N_2017,N_1915,N_1566);
nand U2018 (N_2018,N_1955,N_1512);
and U2019 (N_2019,N_1971,N_1893);
nor U2020 (N_2020,N_1532,N_1913);
nand U2021 (N_2021,N_1695,N_1941);
nor U2022 (N_2022,N_1559,N_1700);
or U2023 (N_2023,N_1681,N_1929);
nand U2024 (N_2024,N_1656,N_1667);
nand U2025 (N_2025,N_1944,N_1828);
or U2026 (N_2026,N_1540,N_1623);
nand U2027 (N_2027,N_1582,N_1545);
nand U2028 (N_2028,N_1866,N_1757);
nand U2029 (N_2029,N_1843,N_1501);
and U2030 (N_2030,N_1928,N_1610);
nand U2031 (N_2031,N_1634,N_1751);
or U2032 (N_2032,N_1717,N_1585);
nor U2033 (N_2033,N_1517,N_1621);
nand U2034 (N_2034,N_1510,N_1597);
nand U2035 (N_2035,N_1921,N_1905);
and U2036 (N_2036,N_1882,N_1603);
nand U2037 (N_2037,N_1937,N_1945);
and U2038 (N_2038,N_1556,N_1965);
and U2039 (N_2039,N_1592,N_1541);
nand U2040 (N_2040,N_1740,N_1830);
nor U2041 (N_2041,N_1979,N_1909);
or U2042 (N_2042,N_1522,N_1551);
nor U2043 (N_2043,N_1811,N_1966);
nor U2044 (N_2044,N_1755,N_1675);
and U2045 (N_2045,N_1553,N_1914);
nand U2046 (N_2046,N_1814,N_1586);
nand U2047 (N_2047,N_1794,N_1699);
nand U2048 (N_2048,N_1785,N_1972);
and U2049 (N_2049,N_1837,N_1764);
nor U2050 (N_2050,N_1642,N_1773);
and U2051 (N_2051,N_1879,N_1840);
and U2052 (N_2052,N_1538,N_1687);
nor U2053 (N_2053,N_1977,N_1509);
or U2054 (N_2054,N_1622,N_1564);
nor U2055 (N_2055,N_1734,N_1784);
or U2056 (N_2056,N_1518,N_1549);
nand U2057 (N_2057,N_1953,N_1865);
or U2058 (N_2058,N_1827,N_1708);
nand U2059 (N_2059,N_1555,N_1528);
nor U2060 (N_2060,N_1758,N_1658);
or U2061 (N_2061,N_1959,N_1782);
nand U2062 (N_2062,N_1500,N_1735);
or U2063 (N_2063,N_1690,N_1875);
nor U2064 (N_2064,N_1906,N_1632);
nor U2065 (N_2065,N_1546,N_1779);
nand U2066 (N_2066,N_1996,N_1833);
or U2067 (N_2067,N_1521,N_1860);
nand U2068 (N_2068,N_1575,N_1548);
nand U2069 (N_2069,N_1737,N_1961);
nand U2070 (N_2070,N_1578,N_1838);
or U2071 (N_2071,N_1560,N_1907);
or U2072 (N_2072,N_1728,N_1672);
nor U2073 (N_2073,N_1981,N_1797);
and U2074 (N_2074,N_1869,N_1676);
or U2075 (N_2075,N_1647,N_1883);
nand U2076 (N_2076,N_1759,N_1884);
or U2077 (N_2077,N_1630,N_1858);
or U2078 (N_2078,N_1697,N_1673);
nand U2079 (N_2079,N_1611,N_1917);
or U2080 (N_2080,N_1653,N_1813);
or U2081 (N_2081,N_1631,N_1507);
or U2082 (N_2082,N_1624,N_1962);
nor U2083 (N_2083,N_1638,N_1857);
nor U2084 (N_2084,N_1557,N_1800);
or U2085 (N_2085,N_1666,N_1982);
or U2086 (N_2086,N_1602,N_1671);
nand U2087 (N_2087,N_1776,N_1766);
and U2088 (N_2088,N_1573,N_1524);
and U2089 (N_2089,N_1851,N_1807);
nor U2090 (N_2090,N_1748,N_1788);
nor U2091 (N_2091,N_1503,N_1892);
nor U2092 (N_2092,N_1946,N_1725);
or U2093 (N_2093,N_1781,N_1635);
and U2094 (N_2094,N_1645,N_1821);
and U2095 (N_2095,N_1829,N_1786);
nand U2096 (N_2096,N_1628,N_1854);
nand U2097 (N_2097,N_1760,N_1763);
and U2098 (N_2098,N_1599,N_1562);
nand U2099 (N_2099,N_1808,N_1940);
or U2100 (N_2100,N_1983,N_1743);
nor U2101 (N_2101,N_1570,N_1682);
and U2102 (N_2102,N_1591,N_1741);
nand U2103 (N_2103,N_1926,N_1769);
or U2104 (N_2104,N_1537,N_1505);
nand U2105 (N_2105,N_1629,N_1799);
and U2106 (N_2106,N_1665,N_1890);
or U2107 (N_2107,N_1519,N_1689);
nor U2108 (N_2108,N_1900,N_1729);
nor U2109 (N_2109,N_1816,N_1956);
and U2110 (N_2110,N_1749,N_1620);
or U2111 (N_2111,N_1772,N_1831);
and U2112 (N_2112,N_1904,N_1711);
nand U2113 (N_2113,N_1873,N_1637);
nand U2114 (N_2114,N_1738,N_1600);
nand U2115 (N_2115,N_1754,N_1565);
nor U2116 (N_2116,N_1934,N_1792);
nand U2117 (N_2117,N_1952,N_1598);
nor U2118 (N_2118,N_1790,N_1720);
nor U2119 (N_2119,N_1722,N_1947);
nor U2120 (N_2120,N_1614,N_1696);
and U2121 (N_2121,N_1579,N_1832);
nor U2122 (N_2122,N_1973,N_1948);
nor U2123 (N_2123,N_1815,N_1664);
nor U2124 (N_2124,N_1862,N_1593);
nand U2125 (N_2125,N_1716,N_1849);
nor U2126 (N_2126,N_1712,N_1770);
and U2127 (N_2127,N_1806,N_1826);
or U2128 (N_2128,N_1818,N_1932);
or U2129 (N_2129,N_1943,N_1942);
and U2130 (N_2130,N_1567,N_1726);
and U2131 (N_2131,N_1791,N_1783);
and U2132 (N_2132,N_1662,N_1569);
nand U2133 (N_2133,N_1721,N_1853);
or U2134 (N_2134,N_1850,N_1935);
nand U2135 (N_2135,N_1516,N_1999);
or U2136 (N_2136,N_1502,N_1706);
or U2137 (N_2137,N_1713,N_1677);
or U2138 (N_2138,N_1767,N_1587);
nand U2139 (N_2139,N_1694,N_1756);
and U2140 (N_2140,N_1871,N_1823);
nor U2141 (N_2141,N_1848,N_1918);
and U2142 (N_2142,N_1732,N_1644);
nand U2143 (N_2143,N_1612,N_1702);
nand U2144 (N_2144,N_1964,N_1731);
nor U2145 (N_2145,N_1825,N_1513);
nand U2146 (N_2146,N_1891,N_1912);
nor U2147 (N_2147,N_1771,N_1719);
nand U2148 (N_2148,N_1985,N_1616);
and U2149 (N_2149,N_1844,N_1601);
or U2150 (N_2150,N_1588,N_1901);
or U2151 (N_2151,N_1609,N_1508);
or U2152 (N_2152,N_1654,N_1868);
or U2153 (N_2153,N_1615,N_1889);
or U2154 (N_2154,N_1657,N_1685);
nor U2155 (N_2155,N_1527,N_1916);
nand U2156 (N_2156,N_1554,N_1698);
and U2157 (N_2157,N_1649,N_1514);
or U2158 (N_2158,N_1558,N_1704);
or U2159 (N_2159,N_1789,N_1577);
and U2160 (N_2160,N_1761,N_1778);
and U2161 (N_2161,N_1836,N_1668);
nand U2162 (N_2162,N_1796,N_1878);
nor U2163 (N_2163,N_1547,N_1692);
or U2164 (N_2164,N_1701,N_1903);
nand U2165 (N_2165,N_1951,N_1563);
or U2166 (N_2166,N_1957,N_1861);
and U2167 (N_2167,N_1908,N_1997);
or U2168 (N_2168,N_1968,N_1793);
or U2169 (N_2169,N_1536,N_1841);
and U2170 (N_2170,N_1580,N_1762);
or U2171 (N_2171,N_1627,N_1750);
or U2172 (N_2172,N_1842,N_1963);
or U2173 (N_2173,N_1626,N_1958);
or U2174 (N_2174,N_1874,N_1534);
nor U2175 (N_2175,N_1847,N_1902);
or U2176 (N_2176,N_1688,N_1930);
and U2177 (N_2177,N_1897,N_1984);
nand U2178 (N_2178,N_1804,N_1552);
xnor U2179 (N_2179,N_1880,N_1660);
or U2180 (N_2180,N_1927,N_1970);
nand U2181 (N_2181,N_1625,N_1768);
nand U2182 (N_2182,N_1727,N_1925);
and U2183 (N_2183,N_1938,N_1684);
or U2184 (N_2184,N_1742,N_1994);
nand U2185 (N_2185,N_1787,N_1693);
or U2186 (N_2186,N_1765,N_1998);
xnor U2187 (N_2187,N_1949,N_1867);
and U2188 (N_2188,N_1618,N_1533);
nand U2189 (N_2189,N_1801,N_1595);
nor U2190 (N_2190,N_1933,N_1659);
or U2191 (N_2191,N_1886,N_1739);
or U2192 (N_2192,N_1529,N_1669);
or U2193 (N_2193,N_1535,N_1543);
nor U2194 (N_2194,N_1745,N_1777);
or U2195 (N_2195,N_1922,N_1594);
and U2196 (N_2196,N_1617,N_1753);
nand U2197 (N_2197,N_1923,N_1931);
nand U2198 (N_2198,N_1639,N_1606);
and U2199 (N_2199,N_1812,N_1920);
nor U2200 (N_2200,N_1863,N_1993);
nor U2201 (N_2201,N_1520,N_1795);
and U2202 (N_2202,N_1990,N_1995);
and U2203 (N_2203,N_1980,N_1709);
or U2204 (N_2204,N_1802,N_1680);
nor U2205 (N_2205,N_1705,N_1989);
and U2206 (N_2206,N_1974,N_1619);
and U2207 (N_2207,N_1939,N_1636);
nand U2208 (N_2208,N_1674,N_1511);
or U2209 (N_2209,N_1542,N_1733);
and U2210 (N_2210,N_1607,N_1747);
nor U2211 (N_2211,N_1820,N_1987);
or U2212 (N_2212,N_1651,N_1608);
and U2213 (N_2213,N_1887,N_1640);
or U2214 (N_2214,N_1736,N_1724);
nor U2215 (N_2215,N_1523,N_1950);
nand U2216 (N_2216,N_1881,N_1752);
or U2217 (N_2217,N_1678,N_1531);
and U2218 (N_2218,N_1530,N_1954);
nand U2219 (N_2219,N_1975,N_1924);
nand U2220 (N_2220,N_1504,N_1613);
and U2221 (N_2221,N_1550,N_1643);
and U2222 (N_2222,N_1670,N_1803);
and U2223 (N_2223,N_1834,N_1969);
xnor U2224 (N_2224,N_1576,N_1967);
nand U2225 (N_2225,N_1910,N_1661);
or U2226 (N_2226,N_1870,N_1978);
nand U2227 (N_2227,N_1683,N_1525);
and U2228 (N_2228,N_1574,N_1936);
and U2229 (N_2229,N_1859,N_1774);
or U2230 (N_2230,N_1877,N_1663);
nor U2231 (N_2231,N_1572,N_1746);
or U2232 (N_2232,N_1855,N_1596);
nand U2233 (N_2233,N_1839,N_1809);
nor U2234 (N_2234,N_1539,N_1822);
or U2235 (N_2235,N_1641,N_1655);
nand U2236 (N_2236,N_1805,N_1568);
nor U2237 (N_2237,N_1876,N_1589);
and U2238 (N_2238,N_1515,N_1571);
nand U2239 (N_2239,N_1707,N_1780);
or U2240 (N_2240,N_1988,N_1888);
or U2241 (N_2241,N_1986,N_1590);
or U2242 (N_2242,N_1686,N_1506);
nand U2243 (N_2243,N_1817,N_1633);
or U2244 (N_2244,N_1898,N_1864);
or U2245 (N_2245,N_1718,N_1960);
and U2246 (N_2246,N_1852,N_1991);
xnor U2247 (N_2247,N_1846,N_1583);
or U2248 (N_2248,N_1919,N_1526);
and U2249 (N_2249,N_1648,N_1976);
and U2250 (N_2250,N_1871,N_1877);
nand U2251 (N_2251,N_1814,N_1747);
or U2252 (N_2252,N_1990,N_1695);
and U2253 (N_2253,N_1848,N_1826);
and U2254 (N_2254,N_1851,N_1512);
and U2255 (N_2255,N_1998,N_1592);
nand U2256 (N_2256,N_1672,N_1963);
xor U2257 (N_2257,N_1772,N_1931);
and U2258 (N_2258,N_1981,N_1573);
nor U2259 (N_2259,N_1947,N_1948);
or U2260 (N_2260,N_1988,N_1699);
nor U2261 (N_2261,N_1708,N_1804);
nand U2262 (N_2262,N_1797,N_1697);
or U2263 (N_2263,N_1738,N_1858);
or U2264 (N_2264,N_1779,N_1643);
nor U2265 (N_2265,N_1741,N_1998);
and U2266 (N_2266,N_1679,N_1969);
nand U2267 (N_2267,N_1883,N_1643);
and U2268 (N_2268,N_1803,N_1687);
nor U2269 (N_2269,N_1902,N_1537);
and U2270 (N_2270,N_1759,N_1708);
and U2271 (N_2271,N_1758,N_1683);
nor U2272 (N_2272,N_1559,N_1772);
and U2273 (N_2273,N_1941,N_1823);
or U2274 (N_2274,N_1608,N_1784);
nor U2275 (N_2275,N_1526,N_1547);
nand U2276 (N_2276,N_1705,N_1778);
and U2277 (N_2277,N_1942,N_1830);
nand U2278 (N_2278,N_1701,N_1838);
or U2279 (N_2279,N_1928,N_1911);
and U2280 (N_2280,N_1629,N_1847);
or U2281 (N_2281,N_1565,N_1868);
nand U2282 (N_2282,N_1542,N_1774);
nor U2283 (N_2283,N_1965,N_1659);
or U2284 (N_2284,N_1824,N_1634);
nor U2285 (N_2285,N_1965,N_1718);
or U2286 (N_2286,N_1598,N_1590);
and U2287 (N_2287,N_1880,N_1697);
nor U2288 (N_2288,N_1620,N_1796);
or U2289 (N_2289,N_1676,N_1811);
and U2290 (N_2290,N_1795,N_1840);
nand U2291 (N_2291,N_1724,N_1671);
and U2292 (N_2292,N_1908,N_1550);
or U2293 (N_2293,N_1798,N_1581);
nand U2294 (N_2294,N_1654,N_1516);
and U2295 (N_2295,N_1993,N_1841);
nor U2296 (N_2296,N_1623,N_1770);
and U2297 (N_2297,N_1819,N_1996);
nand U2298 (N_2298,N_1871,N_1896);
nand U2299 (N_2299,N_1807,N_1532);
nor U2300 (N_2300,N_1557,N_1628);
and U2301 (N_2301,N_1895,N_1958);
nand U2302 (N_2302,N_1668,N_1989);
and U2303 (N_2303,N_1672,N_1629);
or U2304 (N_2304,N_1650,N_1691);
or U2305 (N_2305,N_1703,N_1666);
and U2306 (N_2306,N_1514,N_1648);
nand U2307 (N_2307,N_1968,N_1842);
nand U2308 (N_2308,N_1685,N_1936);
nor U2309 (N_2309,N_1581,N_1624);
nor U2310 (N_2310,N_1677,N_1862);
and U2311 (N_2311,N_1831,N_1929);
or U2312 (N_2312,N_1778,N_1516);
nor U2313 (N_2313,N_1906,N_1865);
and U2314 (N_2314,N_1869,N_1518);
nor U2315 (N_2315,N_1823,N_1672);
nor U2316 (N_2316,N_1947,N_1746);
nand U2317 (N_2317,N_1682,N_1534);
nand U2318 (N_2318,N_1929,N_1795);
and U2319 (N_2319,N_1613,N_1783);
nor U2320 (N_2320,N_1751,N_1801);
nand U2321 (N_2321,N_1766,N_1562);
and U2322 (N_2322,N_1706,N_1832);
and U2323 (N_2323,N_1761,N_1608);
xnor U2324 (N_2324,N_1806,N_1530);
nand U2325 (N_2325,N_1988,N_1509);
or U2326 (N_2326,N_1721,N_1732);
nor U2327 (N_2327,N_1937,N_1769);
and U2328 (N_2328,N_1764,N_1819);
xnor U2329 (N_2329,N_1675,N_1895);
or U2330 (N_2330,N_1568,N_1672);
nand U2331 (N_2331,N_1563,N_1872);
nand U2332 (N_2332,N_1746,N_1545);
nand U2333 (N_2333,N_1843,N_1626);
nand U2334 (N_2334,N_1989,N_1947);
or U2335 (N_2335,N_1786,N_1591);
nand U2336 (N_2336,N_1657,N_1879);
and U2337 (N_2337,N_1877,N_1872);
nand U2338 (N_2338,N_1599,N_1732);
nand U2339 (N_2339,N_1712,N_1829);
nor U2340 (N_2340,N_1872,N_1685);
nor U2341 (N_2341,N_1567,N_1532);
or U2342 (N_2342,N_1794,N_1911);
nor U2343 (N_2343,N_1743,N_1529);
or U2344 (N_2344,N_1717,N_1864);
nor U2345 (N_2345,N_1881,N_1884);
nor U2346 (N_2346,N_1990,N_1504);
nor U2347 (N_2347,N_1978,N_1703);
and U2348 (N_2348,N_1827,N_1527);
nand U2349 (N_2349,N_1886,N_1701);
nand U2350 (N_2350,N_1614,N_1588);
nor U2351 (N_2351,N_1585,N_1589);
nor U2352 (N_2352,N_1964,N_1599);
or U2353 (N_2353,N_1886,N_1699);
nand U2354 (N_2354,N_1651,N_1553);
nand U2355 (N_2355,N_1682,N_1689);
or U2356 (N_2356,N_1945,N_1748);
and U2357 (N_2357,N_1868,N_1780);
nand U2358 (N_2358,N_1668,N_1747);
and U2359 (N_2359,N_1955,N_1768);
nor U2360 (N_2360,N_1516,N_1805);
or U2361 (N_2361,N_1609,N_1557);
and U2362 (N_2362,N_1545,N_1717);
nor U2363 (N_2363,N_1805,N_1667);
nand U2364 (N_2364,N_1768,N_1852);
nor U2365 (N_2365,N_1555,N_1567);
nand U2366 (N_2366,N_1902,N_1987);
and U2367 (N_2367,N_1939,N_1666);
or U2368 (N_2368,N_1906,N_1817);
nand U2369 (N_2369,N_1630,N_1658);
nand U2370 (N_2370,N_1610,N_1702);
nor U2371 (N_2371,N_1525,N_1709);
nand U2372 (N_2372,N_1777,N_1514);
and U2373 (N_2373,N_1807,N_1742);
nor U2374 (N_2374,N_1791,N_1935);
or U2375 (N_2375,N_1821,N_1796);
or U2376 (N_2376,N_1592,N_1754);
nand U2377 (N_2377,N_1648,N_1686);
or U2378 (N_2378,N_1845,N_1627);
nor U2379 (N_2379,N_1558,N_1700);
and U2380 (N_2380,N_1960,N_1918);
nand U2381 (N_2381,N_1733,N_1694);
and U2382 (N_2382,N_1893,N_1834);
nand U2383 (N_2383,N_1677,N_1661);
and U2384 (N_2384,N_1786,N_1842);
or U2385 (N_2385,N_1814,N_1702);
nand U2386 (N_2386,N_1828,N_1696);
or U2387 (N_2387,N_1578,N_1757);
nor U2388 (N_2388,N_1787,N_1943);
nand U2389 (N_2389,N_1650,N_1613);
nor U2390 (N_2390,N_1998,N_1639);
and U2391 (N_2391,N_1720,N_1962);
or U2392 (N_2392,N_1931,N_1990);
nand U2393 (N_2393,N_1933,N_1793);
and U2394 (N_2394,N_1741,N_1569);
and U2395 (N_2395,N_1608,N_1952);
nand U2396 (N_2396,N_1562,N_1882);
nand U2397 (N_2397,N_1818,N_1550);
and U2398 (N_2398,N_1909,N_1843);
and U2399 (N_2399,N_1724,N_1532);
nand U2400 (N_2400,N_1760,N_1983);
nor U2401 (N_2401,N_1918,N_1666);
or U2402 (N_2402,N_1912,N_1818);
and U2403 (N_2403,N_1590,N_1903);
and U2404 (N_2404,N_1736,N_1773);
or U2405 (N_2405,N_1761,N_1819);
or U2406 (N_2406,N_1535,N_1605);
or U2407 (N_2407,N_1864,N_1570);
nor U2408 (N_2408,N_1583,N_1731);
nor U2409 (N_2409,N_1905,N_1662);
or U2410 (N_2410,N_1726,N_1778);
and U2411 (N_2411,N_1520,N_1732);
nor U2412 (N_2412,N_1923,N_1594);
or U2413 (N_2413,N_1503,N_1627);
nor U2414 (N_2414,N_1700,N_1721);
and U2415 (N_2415,N_1890,N_1580);
nor U2416 (N_2416,N_1606,N_1659);
and U2417 (N_2417,N_1598,N_1825);
and U2418 (N_2418,N_1977,N_1848);
nor U2419 (N_2419,N_1939,N_1540);
nor U2420 (N_2420,N_1801,N_1835);
or U2421 (N_2421,N_1622,N_1635);
nor U2422 (N_2422,N_1961,N_1946);
or U2423 (N_2423,N_1745,N_1905);
xor U2424 (N_2424,N_1563,N_1755);
nor U2425 (N_2425,N_1845,N_1790);
nand U2426 (N_2426,N_1940,N_1863);
nor U2427 (N_2427,N_1791,N_1853);
or U2428 (N_2428,N_1803,N_1715);
or U2429 (N_2429,N_1991,N_1942);
or U2430 (N_2430,N_1914,N_1788);
nand U2431 (N_2431,N_1580,N_1968);
nand U2432 (N_2432,N_1604,N_1713);
nand U2433 (N_2433,N_1753,N_1510);
and U2434 (N_2434,N_1969,N_1682);
nand U2435 (N_2435,N_1657,N_1721);
nand U2436 (N_2436,N_1545,N_1975);
nor U2437 (N_2437,N_1669,N_1710);
or U2438 (N_2438,N_1612,N_1773);
or U2439 (N_2439,N_1785,N_1644);
and U2440 (N_2440,N_1923,N_1800);
nor U2441 (N_2441,N_1646,N_1700);
or U2442 (N_2442,N_1570,N_1801);
and U2443 (N_2443,N_1926,N_1826);
nand U2444 (N_2444,N_1835,N_1993);
or U2445 (N_2445,N_1919,N_1992);
xor U2446 (N_2446,N_1674,N_1978);
nor U2447 (N_2447,N_1896,N_1944);
or U2448 (N_2448,N_1622,N_1785);
nor U2449 (N_2449,N_1944,N_1696);
nor U2450 (N_2450,N_1974,N_1554);
nor U2451 (N_2451,N_1700,N_1879);
or U2452 (N_2452,N_1611,N_1816);
or U2453 (N_2453,N_1980,N_1714);
nor U2454 (N_2454,N_1528,N_1664);
nand U2455 (N_2455,N_1780,N_1909);
and U2456 (N_2456,N_1752,N_1699);
or U2457 (N_2457,N_1816,N_1725);
nand U2458 (N_2458,N_1867,N_1698);
nor U2459 (N_2459,N_1748,N_1642);
and U2460 (N_2460,N_1525,N_1857);
nor U2461 (N_2461,N_1964,N_1637);
and U2462 (N_2462,N_1600,N_1604);
nor U2463 (N_2463,N_1908,N_1573);
or U2464 (N_2464,N_1588,N_1970);
nand U2465 (N_2465,N_1536,N_1676);
or U2466 (N_2466,N_1531,N_1675);
or U2467 (N_2467,N_1930,N_1585);
and U2468 (N_2468,N_1870,N_1614);
nand U2469 (N_2469,N_1592,N_1556);
and U2470 (N_2470,N_1958,N_1728);
nor U2471 (N_2471,N_1619,N_1572);
or U2472 (N_2472,N_1736,N_1512);
and U2473 (N_2473,N_1876,N_1791);
and U2474 (N_2474,N_1786,N_1699);
nand U2475 (N_2475,N_1965,N_1645);
and U2476 (N_2476,N_1756,N_1994);
or U2477 (N_2477,N_1761,N_1683);
nor U2478 (N_2478,N_1591,N_1929);
nor U2479 (N_2479,N_1973,N_1783);
nand U2480 (N_2480,N_1931,N_1968);
and U2481 (N_2481,N_1510,N_1647);
nand U2482 (N_2482,N_1644,N_1813);
or U2483 (N_2483,N_1952,N_1923);
and U2484 (N_2484,N_1622,N_1694);
and U2485 (N_2485,N_1944,N_1848);
and U2486 (N_2486,N_1612,N_1689);
nor U2487 (N_2487,N_1621,N_1504);
or U2488 (N_2488,N_1991,N_1559);
nand U2489 (N_2489,N_1771,N_1765);
or U2490 (N_2490,N_1970,N_1632);
nand U2491 (N_2491,N_1829,N_1572);
nor U2492 (N_2492,N_1672,N_1593);
nand U2493 (N_2493,N_1708,N_1828);
and U2494 (N_2494,N_1865,N_1987);
and U2495 (N_2495,N_1796,N_1552);
or U2496 (N_2496,N_1783,N_1935);
nor U2497 (N_2497,N_1578,N_1508);
nor U2498 (N_2498,N_1977,N_1624);
and U2499 (N_2499,N_1910,N_1680);
or U2500 (N_2500,N_2163,N_2216);
nor U2501 (N_2501,N_2347,N_2098);
nor U2502 (N_2502,N_2240,N_2052);
or U2503 (N_2503,N_2110,N_2397);
nor U2504 (N_2504,N_2144,N_2094);
nor U2505 (N_2505,N_2318,N_2349);
and U2506 (N_2506,N_2197,N_2461);
nand U2507 (N_2507,N_2372,N_2267);
or U2508 (N_2508,N_2403,N_2259);
and U2509 (N_2509,N_2025,N_2458);
and U2510 (N_2510,N_2235,N_2096);
or U2511 (N_2511,N_2380,N_2361);
nor U2512 (N_2512,N_2463,N_2258);
nor U2513 (N_2513,N_2445,N_2362);
or U2514 (N_2514,N_2152,N_2474);
or U2515 (N_2515,N_2135,N_2138);
nand U2516 (N_2516,N_2172,N_2218);
nand U2517 (N_2517,N_2151,N_2333);
nor U2518 (N_2518,N_2285,N_2367);
nand U2519 (N_2519,N_2228,N_2226);
nor U2520 (N_2520,N_2194,N_2428);
nor U2521 (N_2521,N_2350,N_2462);
and U2522 (N_2522,N_2024,N_2336);
nand U2523 (N_2523,N_2198,N_2112);
and U2524 (N_2524,N_2328,N_2100);
or U2525 (N_2525,N_2124,N_2008);
nand U2526 (N_2526,N_2447,N_2479);
nand U2527 (N_2527,N_2232,N_2210);
or U2528 (N_2528,N_2014,N_2066);
nor U2529 (N_2529,N_2296,N_2407);
or U2530 (N_2530,N_2340,N_2208);
and U2531 (N_2531,N_2242,N_2034);
or U2532 (N_2532,N_2396,N_2060);
or U2533 (N_2533,N_2040,N_2436);
or U2534 (N_2534,N_2455,N_2320);
nor U2535 (N_2535,N_2425,N_2414);
nand U2536 (N_2536,N_2215,N_2246);
and U2537 (N_2537,N_2290,N_2472);
nand U2538 (N_2538,N_2103,N_2076);
or U2539 (N_2539,N_2402,N_2257);
nand U2540 (N_2540,N_2494,N_2492);
nand U2541 (N_2541,N_2074,N_2470);
and U2542 (N_2542,N_2199,N_2297);
or U2543 (N_2543,N_2227,N_2239);
nor U2544 (N_2544,N_2013,N_2128);
nor U2545 (N_2545,N_2377,N_2272);
nor U2546 (N_2546,N_2373,N_2130);
or U2547 (N_2547,N_2062,N_2486);
and U2548 (N_2548,N_2450,N_2145);
nand U2549 (N_2549,N_2324,N_2108);
nand U2550 (N_2550,N_2159,N_2121);
nand U2551 (N_2551,N_2248,N_2260);
nor U2552 (N_2552,N_2263,N_2497);
or U2553 (N_2553,N_2287,N_2408);
nor U2554 (N_2554,N_2048,N_2203);
nor U2555 (N_2555,N_2384,N_2453);
and U2556 (N_2556,N_2075,N_2432);
nor U2557 (N_2557,N_2224,N_2344);
or U2558 (N_2558,N_2002,N_2032);
nand U2559 (N_2559,N_2165,N_2393);
nor U2560 (N_2560,N_2019,N_2104);
or U2561 (N_2561,N_2120,N_2327);
or U2562 (N_2562,N_2271,N_2364);
nor U2563 (N_2563,N_2038,N_2469);
and U2564 (N_2564,N_2390,N_2378);
nand U2565 (N_2565,N_2427,N_2478);
nand U2566 (N_2566,N_2091,N_2289);
nand U2567 (N_2567,N_2437,N_2017);
nor U2568 (N_2568,N_2173,N_2241);
nor U2569 (N_2569,N_2326,N_2411);
and U2570 (N_2570,N_2149,N_2186);
or U2571 (N_2571,N_2277,N_2119);
nand U2572 (N_2572,N_2348,N_2311);
nor U2573 (N_2573,N_2345,N_2387);
or U2574 (N_2574,N_2442,N_2045);
nor U2575 (N_2575,N_2078,N_2404);
and U2576 (N_2576,N_2280,N_2175);
nor U2577 (N_2577,N_2351,N_2398);
and U2578 (N_2578,N_2243,N_2471);
and U2579 (N_2579,N_2319,N_2370);
nor U2580 (N_2580,N_2132,N_2150);
nand U2581 (N_2581,N_2230,N_2485);
nor U2582 (N_2582,N_2219,N_2309);
nor U2583 (N_2583,N_2214,N_2026);
and U2584 (N_2584,N_2446,N_2368);
nor U2585 (N_2585,N_2421,N_2092);
and U2586 (N_2586,N_2109,N_2449);
nor U2587 (N_2587,N_2457,N_2483);
and U2588 (N_2588,N_2430,N_2031);
or U2589 (N_2589,N_2381,N_2001);
and U2590 (N_2590,N_2256,N_2346);
nor U2591 (N_2591,N_2033,N_2426);
and U2592 (N_2592,N_2184,N_2054);
nand U2593 (N_2593,N_2047,N_2383);
or U2594 (N_2594,N_2342,N_2077);
nand U2595 (N_2595,N_2269,N_2134);
nand U2596 (N_2596,N_2468,N_2356);
or U2597 (N_2597,N_2312,N_2190);
nor U2598 (N_2598,N_2015,N_2394);
nand U2599 (N_2599,N_2391,N_2238);
and U2600 (N_2600,N_2354,N_2058);
or U2601 (N_2601,N_2366,N_2053);
nand U2602 (N_2602,N_2212,N_2051);
and U2603 (N_2603,N_2231,N_2386);
and U2604 (N_2604,N_2050,N_2160);
nor U2605 (N_2605,N_2106,N_2116);
nor U2606 (N_2606,N_2322,N_2295);
nand U2607 (N_2607,N_2292,N_2089);
and U2608 (N_2608,N_2400,N_2158);
and U2609 (N_2609,N_2187,N_2438);
and U2610 (N_2610,N_2064,N_2482);
nand U2611 (N_2611,N_2082,N_2448);
nand U2612 (N_2612,N_2299,N_2087);
nand U2613 (N_2613,N_2360,N_2358);
nand U2614 (N_2614,N_2480,N_2395);
and U2615 (N_2615,N_2245,N_2170);
and U2616 (N_2616,N_2489,N_2374);
and U2617 (N_2617,N_2185,N_2022);
or U2618 (N_2618,N_2417,N_2274);
or U2619 (N_2619,N_2084,N_2466);
nor U2620 (N_2620,N_2423,N_2443);
nor U2621 (N_2621,N_2371,N_2205);
nor U2622 (N_2622,N_2140,N_2307);
nor U2623 (N_2623,N_2379,N_2255);
and U2624 (N_2624,N_2069,N_2491);
and U2625 (N_2625,N_2357,N_2016);
or U2626 (N_2626,N_2153,N_2169);
nand U2627 (N_2627,N_2117,N_2420);
nor U2628 (N_2628,N_2389,N_2063);
nor U2629 (N_2629,N_2317,N_2057);
or U2630 (N_2630,N_2085,N_2353);
and U2631 (N_2631,N_2018,N_2209);
nor U2632 (N_2632,N_2288,N_2382);
nand U2633 (N_2633,N_2441,N_2065);
nand U2634 (N_2634,N_2028,N_2416);
and U2635 (N_2635,N_2237,N_2476);
and U2636 (N_2636,N_2473,N_2095);
and U2637 (N_2637,N_2192,N_2496);
nand U2638 (N_2638,N_2131,N_2464);
nor U2639 (N_2639,N_2102,N_2337);
nor U2640 (N_2640,N_2306,N_2467);
nor U2641 (N_2641,N_2335,N_2139);
nor U2642 (N_2642,N_2189,N_2298);
and U2643 (N_2643,N_2315,N_2101);
nor U2644 (N_2644,N_2451,N_2422);
and U2645 (N_2645,N_2141,N_2343);
nor U2646 (N_2646,N_2253,N_2266);
nand U2647 (N_2647,N_2431,N_2167);
or U2648 (N_2648,N_2251,N_2093);
or U2649 (N_2649,N_2409,N_2369);
nor U2650 (N_2650,N_2113,N_2376);
or U2651 (N_2651,N_2174,N_2146);
nand U2652 (N_2652,N_2495,N_2148);
or U2653 (N_2653,N_2155,N_2250);
nor U2654 (N_2654,N_2433,N_2142);
or U2655 (N_2655,N_2196,N_2268);
or U2656 (N_2656,N_2080,N_2122);
nor U2657 (N_2657,N_2254,N_2365);
nand U2658 (N_2658,N_2329,N_2073);
or U2659 (N_2659,N_2083,N_2180);
nor U2660 (N_2660,N_2162,N_2294);
nand U2661 (N_2661,N_2452,N_2071);
nor U2662 (N_2662,N_2207,N_2410);
nand U2663 (N_2663,N_2265,N_2157);
and U2664 (N_2664,N_2308,N_2392);
nand U2665 (N_2665,N_2220,N_2359);
or U2666 (N_2666,N_2156,N_2178);
or U2667 (N_2667,N_2118,N_2213);
or U2668 (N_2668,N_2275,N_2042);
or U2669 (N_2669,N_2081,N_2202);
or U2670 (N_2670,N_2041,N_2123);
and U2671 (N_2671,N_2114,N_2481);
and U2672 (N_2672,N_2206,N_2284);
or U2673 (N_2673,N_2126,N_2097);
and U2674 (N_2674,N_2136,N_2044);
nand U2675 (N_2675,N_2221,N_2176);
nand U2676 (N_2676,N_2477,N_2279);
nor U2677 (N_2677,N_2424,N_2046);
or U2678 (N_2678,N_2105,N_2043);
nand U2679 (N_2679,N_2171,N_2456);
or U2680 (N_2680,N_2493,N_2107);
or U2681 (N_2681,N_2070,N_2401);
and U2682 (N_2682,N_2222,N_2177);
and U2683 (N_2683,N_2023,N_2183);
nand U2684 (N_2684,N_2475,N_2303);
or U2685 (N_2685,N_2440,N_2300);
nand U2686 (N_2686,N_2059,N_2498);
or U2687 (N_2687,N_2049,N_2405);
nor U2688 (N_2688,N_2161,N_2278);
nor U2689 (N_2689,N_2164,N_2444);
nand U2690 (N_2690,N_2154,N_2276);
nor U2691 (N_2691,N_2166,N_2439);
nor U2692 (N_2692,N_2434,N_2419);
and U2693 (N_2693,N_2191,N_2286);
nor U2694 (N_2694,N_2454,N_2027);
nor U2695 (N_2695,N_2168,N_2030);
nor U2696 (N_2696,N_2037,N_2282);
or U2697 (N_2697,N_2301,N_2325);
or U2698 (N_2698,N_2460,N_2007);
nand U2699 (N_2699,N_2039,N_2035);
or U2700 (N_2700,N_2127,N_2310);
nor U2701 (N_2701,N_2399,N_2252);
or U2702 (N_2702,N_2143,N_2179);
nand U2703 (N_2703,N_2003,N_2200);
and U2704 (N_2704,N_2264,N_2204);
and U2705 (N_2705,N_2293,N_2339);
nor U2706 (N_2706,N_2036,N_2261);
nand U2707 (N_2707,N_2262,N_2385);
nor U2708 (N_2708,N_2217,N_2316);
or U2709 (N_2709,N_2321,N_2195);
or U2710 (N_2710,N_2229,N_2029);
nand U2711 (N_2711,N_2193,N_2247);
nand U2712 (N_2712,N_2465,N_2188);
and U2713 (N_2713,N_2270,N_2413);
nand U2714 (N_2714,N_2225,N_2484);
nor U2715 (N_2715,N_2459,N_2090);
and U2716 (N_2716,N_2061,N_2223);
and U2717 (N_2717,N_2236,N_2291);
or U2718 (N_2718,N_2012,N_2115);
or U2719 (N_2719,N_2020,N_2305);
nand U2720 (N_2720,N_2375,N_2137);
xnor U2721 (N_2721,N_2182,N_2006);
and U2722 (N_2722,N_2429,N_2129);
nand U2723 (N_2723,N_2133,N_2181);
and U2724 (N_2724,N_2211,N_2338);
nand U2725 (N_2725,N_2283,N_2233);
and U2726 (N_2726,N_2304,N_2011);
nor U2727 (N_2727,N_2435,N_2088);
and U2728 (N_2728,N_2147,N_2249);
and U2729 (N_2729,N_2334,N_2099);
nor U2730 (N_2730,N_2125,N_2488);
or U2731 (N_2731,N_2352,N_2000);
nor U2732 (N_2732,N_2234,N_2314);
nand U2733 (N_2733,N_2281,N_2004);
nand U2734 (N_2734,N_2067,N_2010);
and U2735 (N_2735,N_2302,N_2363);
or U2736 (N_2736,N_2021,N_2406);
and U2737 (N_2737,N_2273,N_2313);
and U2738 (N_2738,N_2086,N_2388);
and U2739 (N_2739,N_2355,N_2499);
nand U2740 (N_2740,N_2418,N_2009);
nor U2741 (N_2741,N_2244,N_2490);
nand U2742 (N_2742,N_2056,N_2068);
or U2743 (N_2743,N_2332,N_2415);
or U2744 (N_2744,N_2412,N_2055);
nand U2745 (N_2745,N_2341,N_2072);
nor U2746 (N_2746,N_2005,N_2487);
nand U2747 (N_2747,N_2111,N_2201);
nor U2748 (N_2748,N_2079,N_2330);
nor U2749 (N_2749,N_2323,N_2331);
nand U2750 (N_2750,N_2036,N_2417);
and U2751 (N_2751,N_2083,N_2168);
nand U2752 (N_2752,N_2485,N_2447);
nand U2753 (N_2753,N_2300,N_2066);
nor U2754 (N_2754,N_2035,N_2442);
nor U2755 (N_2755,N_2212,N_2118);
nor U2756 (N_2756,N_2277,N_2483);
nand U2757 (N_2757,N_2395,N_2498);
nand U2758 (N_2758,N_2060,N_2161);
nand U2759 (N_2759,N_2297,N_2362);
nand U2760 (N_2760,N_2439,N_2323);
or U2761 (N_2761,N_2190,N_2067);
nand U2762 (N_2762,N_2217,N_2141);
or U2763 (N_2763,N_2469,N_2113);
and U2764 (N_2764,N_2114,N_2267);
nand U2765 (N_2765,N_2056,N_2185);
and U2766 (N_2766,N_2185,N_2119);
nor U2767 (N_2767,N_2034,N_2234);
and U2768 (N_2768,N_2004,N_2230);
nor U2769 (N_2769,N_2476,N_2034);
or U2770 (N_2770,N_2291,N_2133);
or U2771 (N_2771,N_2074,N_2027);
and U2772 (N_2772,N_2382,N_2191);
or U2773 (N_2773,N_2174,N_2243);
nor U2774 (N_2774,N_2447,N_2250);
and U2775 (N_2775,N_2348,N_2467);
and U2776 (N_2776,N_2198,N_2208);
nor U2777 (N_2777,N_2376,N_2145);
nor U2778 (N_2778,N_2240,N_2394);
nand U2779 (N_2779,N_2282,N_2286);
and U2780 (N_2780,N_2270,N_2324);
or U2781 (N_2781,N_2235,N_2210);
nor U2782 (N_2782,N_2272,N_2450);
and U2783 (N_2783,N_2144,N_2148);
nand U2784 (N_2784,N_2335,N_2086);
and U2785 (N_2785,N_2234,N_2125);
nand U2786 (N_2786,N_2389,N_2381);
nor U2787 (N_2787,N_2084,N_2139);
nand U2788 (N_2788,N_2174,N_2396);
nor U2789 (N_2789,N_2004,N_2162);
nor U2790 (N_2790,N_2384,N_2128);
and U2791 (N_2791,N_2401,N_2288);
or U2792 (N_2792,N_2372,N_2074);
nor U2793 (N_2793,N_2051,N_2338);
or U2794 (N_2794,N_2061,N_2199);
or U2795 (N_2795,N_2346,N_2146);
nand U2796 (N_2796,N_2220,N_2165);
or U2797 (N_2797,N_2324,N_2074);
nor U2798 (N_2798,N_2465,N_2135);
nand U2799 (N_2799,N_2238,N_2118);
nor U2800 (N_2800,N_2128,N_2322);
nor U2801 (N_2801,N_2152,N_2148);
or U2802 (N_2802,N_2198,N_2325);
nor U2803 (N_2803,N_2220,N_2248);
nor U2804 (N_2804,N_2098,N_2247);
or U2805 (N_2805,N_2137,N_2202);
nor U2806 (N_2806,N_2140,N_2091);
xor U2807 (N_2807,N_2014,N_2097);
and U2808 (N_2808,N_2229,N_2240);
and U2809 (N_2809,N_2441,N_2452);
or U2810 (N_2810,N_2369,N_2258);
nand U2811 (N_2811,N_2396,N_2251);
nor U2812 (N_2812,N_2105,N_2427);
nand U2813 (N_2813,N_2422,N_2364);
nor U2814 (N_2814,N_2078,N_2422);
or U2815 (N_2815,N_2079,N_2178);
and U2816 (N_2816,N_2493,N_2294);
or U2817 (N_2817,N_2458,N_2206);
nand U2818 (N_2818,N_2275,N_2192);
and U2819 (N_2819,N_2091,N_2259);
and U2820 (N_2820,N_2138,N_2471);
and U2821 (N_2821,N_2155,N_2192);
or U2822 (N_2822,N_2325,N_2433);
or U2823 (N_2823,N_2068,N_2211);
or U2824 (N_2824,N_2109,N_2485);
or U2825 (N_2825,N_2456,N_2432);
nand U2826 (N_2826,N_2499,N_2371);
and U2827 (N_2827,N_2150,N_2127);
or U2828 (N_2828,N_2215,N_2355);
or U2829 (N_2829,N_2166,N_2126);
nor U2830 (N_2830,N_2389,N_2335);
nand U2831 (N_2831,N_2111,N_2048);
and U2832 (N_2832,N_2352,N_2260);
nor U2833 (N_2833,N_2276,N_2484);
or U2834 (N_2834,N_2382,N_2343);
nand U2835 (N_2835,N_2191,N_2264);
nand U2836 (N_2836,N_2435,N_2362);
nor U2837 (N_2837,N_2203,N_2120);
nor U2838 (N_2838,N_2335,N_2218);
nand U2839 (N_2839,N_2110,N_2145);
or U2840 (N_2840,N_2298,N_2494);
and U2841 (N_2841,N_2134,N_2484);
and U2842 (N_2842,N_2332,N_2491);
and U2843 (N_2843,N_2216,N_2071);
nand U2844 (N_2844,N_2314,N_2355);
or U2845 (N_2845,N_2468,N_2038);
or U2846 (N_2846,N_2439,N_2006);
nand U2847 (N_2847,N_2442,N_2360);
or U2848 (N_2848,N_2446,N_2111);
or U2849 (N_2849,N_2490,N_2383);
nand U2850 (N_2850,N_2449,N_2086);
or U2851 (N_2851,N_2128,N_2490);
and U2852 (N_2852,N_2473,N_2027);
nor U2853 (N_2853,N_2255,N_2082);
nand U2854 (N_2854,N_2092,N_2482);
nand U2855 (N_2855,N_2155,N_2336);
nor U2856 (N_2856,N_2108,N_2275);
nand U2857 (N_2857,N_2443,N_2394);
nand U2858 (N_2858,N_2309,N_2408);
nand U2859 (N_2859,N_2240,N_2177);
nor U2860 (N_2860,N_2417,N_2065);
and U2861 (N_2861,N_2398,N_2103);
and U2862 (N_2862,N_2452,N_2498);
or U2863 (N_2863,N_2480,N_2188);
nand U2864 (N_2864,N_2425,N_2355);
nor U2865 (N_2865,N_2104,N_2064);
and U2866 (N_2866,N_2135,N_2014);
nand U2867 (N_2867,N_2156,N_2431);
and U2868 (N_2868,N_2401,N_2440);
or U2869 (N_2869,N_2489,N_2499);
nand U2870 (N_2870,N_2004,N_2033);
nand U2871 (N_2871,N_2371,N_2461);
and U2872 (N_2872,N_2031,N_2474);
xnor U2873 (N_2873,N_2345,N_2477);
nor U2874 (N_2874,N_2425,N_2204);
and U2875 (N_2875,N_2002,N_2222);
nand U2876 (N_2876,N_2124,N_2025);
nand U2877 (N_2877,N_2014,N_2039);
and U2878 (N_2878,N_2087,N_2437);
nand U2879 (N_2879,N_2091,N_2125);
nor U2880 (N_2880,N_2330,N_2105);
nand U2881 (N_2881,N_2338,N_2322);
nand U2882 (N_2882,N_2164,N_2003);
or U2883 (N_2883,N_2302,N_2378);
or U2884 (N_2884,N_2309,N_2250);
or U2885 (N_2885,N_2369,N_2039);
nand U2886 (N_2886,N_2090,N_2184);
nor U2887 (N_2887,N_2077,N_2000);
nor U2888 (N_2888,N_2472,N_2441);
xor U2889 (N_2889,N_2471,N_2049);
and U2890 (N_2890,N_2322,N_2455);
nor U2891 (N_2891,N_2262,N_2165);
and U2892 (N_2892,N_2319,N_2084);
and U2893 (N_2893,N_2310,N_2285);
nor U2894 (N_2894,N_2192,N_2106);
nor U2895 (N_2895,N_2381,N_2154);
nor U2896 (N_2896,N_2165,N_2058);
nor U2897 (N_2897,N_2408,N_2143);
nand U2898 (N_2898,N_2013,N_2061);
nor U2899 (N_2899,N_2454,N_2268);
nand U2900 (N_2900,N_2038,N_2422);
nor U2901 (N_2901,N_2177,N_2255);
nor U2902 (N_2902,N_2127,N_2132);
and U2903 (N_2903,N_2133,N_2245);
nor U2904 (N_2904,N_2275,N_2480);
nand U2905 (N_2905,N_2302,N_2384);
or U2906 (N_2906,N_2372,N_2342);
nor U2907 (N_2907,N_2131,N_2251);
and U2908 (N_2908,N_2105,N_2279);
and U2909 (N_2909,N_2453,N_2239);
nand U2910 (N_2910,N_2259,N_2452);
or U2911 (N_2911,N_2159,N_2436);
or U2912 (N_2912,N_2460,N_2240);
nand U2913 (N_2913,N_2118,N_2229);
nand U2914 (N_2914,N_2448,N_2081);
nand U2915 (N_2915,N_2205,N_2054);
nor U2916 (N_2916,N_2034,N_2455);
nand U2917 (N_2917,N_2027,N_2462);
nand U2918 (N_2918,N_2234,N_2069);
or U2919 (N_2919,N_2332,N_2371);
or U2920 (N_2920,N_2044,N_2010);
and U2921 (N_2921,N_2449,N_2074);
or U2922 (N_2922,N_2195,N_2329);
and U2923 (N_2923,N_2220,N_2333);
or U2924 (N_2924,N_2495,N_2486);
and U2925 (N_2925,N_2163,N_2224);
and U2926 (N_2926,N_2035,N_2106);
or U2927 (N_2927,N_2369,N_2200);
and U2928 (N_2928,N_2008,N_2322);
or U2929 (N_2929,N_2100,N_2041);
nor U2930 (N_2930,N_2268,N_2328);
nor U2931 (N_2931,N_2179,N_2475);
or U2932 (N_2932,N_2061,N_2363);
nor U2933 (N_2933,N_2077,N_2004);
and U2934 (N_2934,N_2281,N_2331);
nand U2935 (N_2935,N_2069,N_2077);
and U2936 (N_2936,N_2096,N_2457);
nor U2937 (N_2937,N_2145,N_2486);
nand U2938 (N_2938,N_2160,N_2381);
nand U2939 (N_2939,N_2002,N_2463);
nand U2940 (N_2940,N_2431,N_2418);
or U2941 (N_2941,N_2235,N_2315);
nor U2942 (N_2942,N_2164,N_2110);
nand U2943 (N_2943,N_2313,N_2202);
or U2944 (N_2944,N_2286,N_2434);
or U2945 (N_2945,N_2169,N_2480);
and U2946 (N_2946,N_2171,N_2434);
nand U2947 (N_2947,N_2047,N_2479);
and U2948 (N_2948,N_2438,N_2302);
nor U2949 (N_2949,N_2102,N_2394);
and U2950 (N_2950,N_2375,N_2463);
and U2951 (N_2951,N_2446,N_2195);
nand U2952 (N_2952,N_2320,N_2069);
or U2953 (N_2953,N_2192,N_2238);
and U2954 (N_2954,N_2406,N_2127);
nor U2955 (N_2955,N_2376,N_2193);
nand U2956 (N_2956,N_2436,N_2134);
and U2957 (N_2957,N_2171,N_2125);
nand U2958 (N_2958,N_2000,N_2439);
nor U2959 (N_2959,N_2084,N_2409);
nor U2960 (N_2960,N_2183,N_2406);
nand U2961 (N_2961,N_2086,N_2305);
and U2962 (N_2962,N_2227,N_2065);
nor U2963 (N_2963,N_2108,N_2086);
nand U2964 (N_2964,N_2155,N_2387);
nand U2965 (N_2965,N_2268,N_2462);
or U2966 (N_2966,N_2196,N_2054);
nor U2967 (N_2967,N_2150,N_2233);
nor U2968 (N_2968,N_2437,N_2285);
or U2969 (N_2969,N_2189,N_2423);
and U2970 (N_2970,N_2375,N_2073);
nor U2971 (N_2971,N_2464,N_2490);
and U2972 (N_2972,N_2499,N_2303);
nor U2973 (N_2973,N_2220,N_2197);
or U2974 (N_2974,N_2292,N_2180);
nor U2975 (N_2975,N_2175,N_2122);
nand U2976 (N_2976,N_2257,N_2325);
or U2977 (N_2977,N_2495,N_2068);
and U2978 (N_2978,N_2020,N_2152);
and U2979 (N_2979,N_2303,N_2462);
nand U2980 (N_2980,N_2321,N_2137);
nor U2981 (N_2981,N_2489,N_2185);
nor U2982 (N_2982,N_2381,N_2316);
or U2983 (N_2983,N_2369,N_2017);
nor U2984 (N_2984,N_2337,N_2302);
nor U2985 (N_2985,N_2201,N_2498);
nand U2986 (N_2986,N_2007,N_2293);
nor U2987 (N_2987,N_2120,N_2053);
nor U2988 (N_2988,N_2277,N_2034);
nor U2989 (N_2989,N_2164,N_2448);
or U2990 (N_2990,N_2021,N_2422);
nor U2991 (N_2991,N_2038,N_2124);
or U2992 (N_2992,N_2416,N_2459);
or U2993 (N_2993,N_2444,N_2286);
and U2994 (N_2994,N_2390,N_2071);
and U2995 (N_2995,N_2139,N_2451);
or U2996 (N_2996,N_2216,N_2276);
or U2997 (N_2997,N_2295,N_2431);
nand U2998 (N_2998,N_2390,N_2423);
or U2999 (N_2999,N_2075,N_2273);
nor UO_0 (O_0,N_2789,N_2618);
and UO_1 (O_1,N_2508,N_2562);
and UO_2 (O_2,N_2863,N_2503);
nor UO_3 (O_3,N_2895,N_2864);
and UO_4 (O_4,N_2719,N_2885);
nand UO_5 (O_5,N_2581,N_2910);
nor UO_6 (O_6,N_2643,N_2966);
or UO_7 (O_7,N_2671,N_2753);
or UO_8 (O_8,N_2665,N_2927);
and UO_9 (O_9,N_2876,N_2920);
or UO_10 (O_10,N_2994,N_2820);
nand UO_11 (O_11,N_2795,N_2999);
nor UO_12 (O_12,N_2914,N_2855);
and UO_13 (O_13,N_2575,N_2580);
nor UO_14 (O_14,N_2611,N_2880);
and UO_15 (O_15,N_2942,N_2934);
nand UO_16 (O_16,N_2757,N_2916);
or UO_17 (O_17,N_2553,N_2869);
or UO_18 (O_18,N_2722,N_2590);
or UO_19 (O_19,N_2653,N_2632);
or UO_20 (O_20,N_2662,N_2735);
and UO_21 (O_21,N_2793,N_2734);
nor UO_22 (O_22,N_2723,N_2774);
nor UO_23 (O_23,N_2906,N_2560);
and UO_24 (O_24,N_2597,N_2955);
and UO_25 (O_25,N_2993,N_2752);
nand UO_26 (O_26,N_2658,N_2822);
nand UO_27 (O_27,N_2799,N_2677);
nand UO_28 (O_28,N_2907,N_2610);
nor UO_29 (O_29,N_2992,N_2633);
and UO_30 (O_30,N_2782,N_2511);
or UO_31 (O_31,N_2804,N_2787);
nor UO_32 (O_32,N_2932,N_2681);
nor UO_33 (O_33,N_2922,N_2856);
nand UO_34 (O_34,N_2529,N_2981);
and UO_35 (O_35,N_2741,N_2814);
nor UO_36 (O_36,N_2953,N_2800);
nor UO_37 (O_37,N_2680,N_2874);
nand UO_38 (O_38,N_2840,N_2860);
nand UO_39 (O_39,N_2875,N_2641);
nand UO_40 (O_40,N_2850,N_2768);
or UO_41 (O_41,N_2656,N_2939);
nor UO_42 (O_42,N_2829,N_2563);
or UO_43 (O_43,N_2520,N_2676);
nand UO_44 (O_44,N_2565,N_2531);
nand UO_45 (O_45,N_2970,N_2644);
nor UO_46 (O_46,N_2646,N_2550);
or UO_47 (O_47,N_2897,N_2724);
and UO_48 (O_48,N_2542,N_2851);
and UO_49 (O_49,N_2688,N_2728);
nand UO_50 (O_50,N_2823,N_2758);
or UO_51 (O_51,N_2903,N_2819);
and UO_52 (O_52,N_2890,N_2905);
nand UO_53 (O_53,N_2978,N_2504);
nand UO_54 (O_54,N_2926,N_2586);
or UO_55 (O_55,N_2567,N_2852);
and UO_56 (O_56,N_2969,N_2501);
nand UO_57 (O_57,N_2938,N_2522);
or UO_58 (O_58,N_2766,N_2785);
nor UO_59 (O_59,N_2614,N_2996);
or UO_60 (O_60,N_2568,N_2647);
nand UO_61 (O_61,N_2594,N_2783);
nor UO_62 (O_62,N_2827,N_2990);
or UO_63 (O_63,N_2691,N_2579);
nand UO_64 (O_64,N_2767,N_2866);
nand UO_65 (O_65,N_2651,N_2726);
nor UO_66 (O_66,N_2527,N_2925);
nand UO_67 (O_67,N_2707,N_2849);
and UO_68 (O_68,N_2941,N_2976);
and UO_69 (O_69,N_2837,N_2745);
nand UO_70 (O_70,N_2909,N_2507);
nand UO_71 (O_71,N_2652,N_2937);
nor UO_72 (O_72,N_2929,N_2685);
or UO_73 (O_73,N_2603,N_2706);
nand UO_74 (O_74,N_2986,N_2912);
nor UO_75 (O_75,N_2718,N_2818);
and UO_76 (O_76,N_2877,N_2900);
nand UO_77 (O_77,N_2985,N_2500);
and UO_78 (O_78,N_2606,N_2975);
nand UO_79 (O_79,N_2773,N_2808);
and UO_80 (O_80,N_2601,N_2868);
nand UO_81 (O_81,N_2881,N_2809);
nand UO_82 (O_82,N_2836,N_2779);
or UO_83 (O_83,N_2589,N_2843);
and UO_84 (O_84,N_2729,N_2502);
and UO_85 (O_85,N_2667,N_2867);
nor UO_86 (O_86,N_2695,N_2626);
xnor UO_87 (O_87,N_2845,N_2694);
and UO_88 (O_88,N_2717,N_2893);
or UO_89 (O_89,N_2748,N_2648);
nor UO_90 (O_90,N_2564,N_2620);
nor UO_91 (O_91,N_2515,N_2848);
xnor UO_92 (O_92,N_2525,N_2742);
nor UO_93 (O_93,N_2721,N_2596);
nand UO_94 (O_94,N_2842,N_2991);
nand UO_95 (O_95,N_2540,N_2640);
nand UO_96 (O_96,N_2805,N_2740);
nand UO_97 (O_97,N_2686,N_2655);
nand UO_98 (O_98,N_2796,N_2664);
and UO_99 (O_99,N_2810,N_2638);
nand UO_100 (O_100,N_2858,N_2760);
nand UO_101 (O_101,N_2791,N_2730);
nand UO_102 (O_102,N_2621,N_2672);
or UO_103 (O_103,N_2624,N_2687);
nand UO_104 (O_104,N_2835,N_2576);
nor UO_105 (O_105,N_2534,N_2595);
or UO_106 (O_106,N_2551,N_2790);
nor UO_107 (O_107,N_2711,N_2702);
and UO_108 (O_108,N_2798,N_2678);
xnor UO_109 (O_109,N_2746,N_2547);
or UO_110 (O_110,N_2598,N_2593);
nor UO_111 (O_111,N_2983,N_2612);
nor UO_112 (O_112,N_2519,N_2518);
or UO_113 (O_113,N_2965,N_2698);
or UO_114 (O_114,N_2727,N_2764);
or UO_115 (O_115,N_2731,N_2821);
and UO_116 (O_116,N_2961,N_2585);
and UO_117 (O_117,N_2803,N_2539);
or UO_118 (O_118,N_2923,N_2548);
nor UO_119 (O_119,N_2936,N_2989);
and UO_120 (O_120,N_2960,N_2627);
nand UO_121 (O_121,N_2919,N_2962);
nand UO_122 (O_122,N_2716,N_2878);
nand UO_123 (O_123,N_2904,N_2571);
and UO_124 (O_124,N_2690,N_2834);
and UO_125 (O_125,N_2888,N_2535);
nand UO_126 (O_126,N_2988,N_2951);
nor UO_127 (O_127,N_2908,N_2675);
nand UO_128 (O_128,N_2754,N_2898);
nor UO_129 (O_129,N_2591,N_2533);
nor UO_130 (O_130,N_2668,N_2846);
and UO_131 (O_131,N_2733,N_2825);
nand UO_132 (O_132,N_2870,N_2736);
nand UO_133 (O_133,N_2543,N_2854);
and UO_134 (O_134,N_2549,N_2828);
nor UO_135 (O_135,N_2604,N_2639);
or UO_136 (O_136,N_2645,N_2913);
nor UO_137 (O_137,N_2725,N_2708);
or UO_138 (O_138,N_2657,N_2714);
or UO_139 (O_139,N_2583,N_2882);
and UO_140 (O_140,N_2894,N_2781);
nand UO_141 (O_141,N_2710,N_2896);
nand UO_142 (O_142,N_2873,N_2984);
nand UO_143 (O_143,N_2801,N_2756);
nor UO_144 (O_144,N_2578,N_2751);
nand UO_145 (O_145,N_2931,N_2509);
nor UO_146 (O_146,N_2683,N_2972);
or UO_147 (O_147,N_2924,N_2552);
nand UO_148 (O_148,N_2577,N_2505);
and UO_149 (O_149,N_2968,N_2744);
or UO_150 (O_150,N_2623,N_2602);
or UO_151 (O_151,N_2634,N_2699);
or UO_152 (O_152,N_2964,N_2977);
and UO_153 (O_153,N_2949,N_2556);
or UO_154 (O_154,N_2609,N_2558);
or UO_155 (O_155,N_2701,N_2523);
or UO_156 (O_156,N_2940,N_2625);
nor UO_157 (O_157,N_2689,N_2802);
nand UO_158 (O_158,N_2629,N_2713);
nand UO_159 (O_159,N_2792,N_2546);
nand UO_160 (O_160,N_2738,N_2622);
and UO_161 (O_161,N_2899,N_2739);
or UO_162 (O_162,N_2831,N_2732);
nand UO_163 (O_163,N_2998,N_2636);
nor UO_164 (O_164,N_2862,N_2559);
nor UO_165 (O_165,N_2737,N_2514);
nand UO_166 (O_166,N_2945,N_2704);
nand UO_167 (O_167,N_2824,N_2761);
nand UO_168 (O_168,N_2588,N_2765);
or UO_169 (O_169,N_2812,N_2649);
nand UO_170 (O_170,N_2911,N_2884);
nand UO_171 (O_171,N_2816,N_2660);
nand UO_172 (O_172,N_2817,N_2510);
nor UO_173 (O_173,N_2599,N_2674);
and UO_174 (O_174,N_2679,N_2715);
nor UO_175 (O_175,N_2947,N_2918);
or UO_176 (O_176,N_2669,N_2616);
or UO_177 (O_177,N_2631,N_2815);
nor UO_178 (O_178,N_2743,N_2794);
nor UO_179 (O_179,N_2592,N_2557);
or UO_180 (O_180,N_2720,N_2666);
and UO_181 (O_181,N_2569,N_2974);
or UO_182 (O_182,N_2784,N_2630);
and UO_183 (O_183,N_2865,N_2959);
nand UO_184 (O_184,N_2997,N_2703);
and UO_185 (O_185,N_2524,N_2747);
nand UO_186 (O_186,N_2635,N_2692);
nor UO_187 (O_187,N_2709,N_2830);
and UO_188 (O_188,N_2617,N_2980);
nand UO_189 (O_189,N_2750,N_2570);
nand UO_190 (O_190,N_2544,N_2841);
and UO_191 (O_191,N_2826,N_2807);
xnor UO_192 (O_192,N_2554,N_2513);
nand UO_193 (O_193,N_2697,N_2987);
nor UO_194 (O_194,N_2853,N_2693);
nor UO_195 (O_195,N_2573,N_2839);
nor UO_196 (O_196,N_2545,N_2654);
or UO_197 (O_197,N_2861,N_2526);
xor UO_198 (O_198,N_2628,N_2917);
nand UO_199 (O_199,N_2541,N_2771);
nand UO_200 (O_200,N_2650,N_2901);
or UO_201 (O_201,N_2883,N_2673);
nand UO_202 (O_202,N_2517,N_2608);
nand UO_203 (O_203,N_2770,N_2956);
nor UO_204 (O_204,N_2670,N_2530);
and UO_205 (O_205,N_2950,N_2682);
nor UO_206 (O_206,N_2538,N_2892);
nand UO_207 (O_207,N_2948,N_2619);
nor UO_208 (O_208,N_2933,N_2555);
and UO_209 (O_209,N_2712,N_2561);
or UO_210 (O_210,N_2776,N_2661);
or UO_211 (O_211,N_2944,N_2973);
nor UO_212 (O_212,N_2642,N_2512);
nor UO_213 (O_213,N_2763,N_2982);
and UO_214 (O_214,N_2921,N_2684);
nor UO_215 (O_215,N_2777,N_2943);
or UO_216 (O_216,N_2755,N_2915);
nand UO_217 (O_217,N_2607,N_2946);
xnor UO_218 (O_218,N_2957,N_2537);
or UO_219 (O_219,N_2600,N_2952);
nand UO_220 (O_220,N_2582,N_2887);
nand UO_221 (O_221,N_2963,N_2954);
and UO_222 (O_222,N_2700,N_2902);
and UO_223 (O_223,N_2615,N_2847);
xor UO_224 (O_224,N_2572,N_2786);
and UO_225 (O_225,N_2775,N_2780);
nor UO_226 (O_226,N_2659,N_2979);
nor UO_227 (O_227,N_2971,N_2872);
nand UO_228 (O_228,N_2528,N_2566);
nor UO_229 (O_229,N_2705,N_2613);
or UO_230 (O_230,N_2769,N_2813);
and UO_231 (O_231,N_2532,N_2759);
nor UO_232 (O_232,N_2833,N_2844);
and UO_233 (O_233,N_2521,N_2762);
or UO_234 (O_234,N_2832,N_2838);
and UO_235 (O_235,N_2749,N_2584);
nor UO_236 (O_236,N_2891,N_2928);
or UO_237 (O_237,N_2637,N_2772);
and UO_238 (O_238,N_2886,N_2506);
or UO_239 (O_239,N_2859,N_2516);
or UO_240 (O_240,N_2536,N_2574);
nand UO_241 (O_241,N_2696,N_2587);
nand UO_242 (O_242,N_2958,N_2879);
or UO_243 (O_243,N_2995,N_2806);
or UO_244 (O_244,N_2871,N_2663);
and UO_245 (O_245,N_2811,N_2778);
nand UO_246 (O_246,N_2857,N_2967);
nand UO_247 (O_247,N_2889,N_2797);
nand UO_248 (O_248,N_2788,N_2605);
nand UO_249 (O_249,N_2935,N_2930);
or UO_250 (O_250,N_2642,N_2909);
xor UO_251 (O_251,N_2906,N_2864);
and UO_252 (O_252,N_2994,N_2506);
and UO_253 (O_253,N_2938,N_2680);
and UO_254 (O_254,N_2941,N_2903);
nor UO_255 (O_255,N_2885,N_2854);
nor UO_256 (O_256,N_2632,N_2559);
and UO_257 (O_257,N_2567,N_2787);
and UO_258 (O_258,N_2770,N_2633);
nand UO_259 (O_259,N_2869,N_2899);
nor UO_260 (O_260,N_2812,N_2752);
nand UO_261 (O_261,N_2720,N_2999);
or UO_262 (O_262,N_2976,N_2500);
nand UO_263 (O_263,N_2551,N_2748);
or UO_264 (O_264,N_2937,N_2785);
nor UO_265 (O_265,N_2668,N_2906);
nand UO_266 (O_266,N_2512,N_2552);
nor UO_267 (O_267,N_2825,N_2799);
nor UO_268 (O_268,N_2545,N_2845);
or UO_269 (O_269,N_2636,N_2818);
and UO_270 (O_270,N_2698,N_2582);
and UO_271 (O_271,N_2615,N_2568);
nand UO_272 (O_272,N_2681,N_2741);
or UO_273 (O_273,N_2576,N_2949);
nand UO_274 (O_274,N_2884,N_2813);
and UO_275 (O_275,N_2966,N_2752);
and UO_276 (O_276,N_2843,N_2941);
nor UO_277 (O_277,N_2827,N_2648);
and UO_278 (O_278,N_2585,N_2731);
and UO_279 (O_279,N_2585,N_2584);
or UO_280 (O_280,N_2713,N_2721);
and UO_281 (O_281,N_2829,N_2853);
and UO_282 (O_282,N_2912,N_2562);
nand UO_283 (O_283,N_2651,N_2607);
nand UO_284 (O_284,N_2586,N_2895);
and UO_285 (O_285,N_2720,N_2751);
or UO_286 (O_286,N_2951,N_2616);
xor UO_287 (O_287,N_2948,N_2729);
nand UO_288 (O_288,N_2737,N_2850);
nand UO_289 (O_289,N_2664,N_2744);
or UO_290 (O_290,N_2735,N_2645);
nand UO_291 (O_291,N_2804,N_2983);
and UO_292 (O_292,N_2515,N_2569);
or UO_293 (O_293,N_2683,N_2597);
or UO_294 (O_294,N_2541,N_2942);
nand UO_295 (O_295,N_2543,N_2768);
and UO_296 (O_296,N_2684,N_2841);
or UO_297 (O_297,N_2638,N_2855);
nor UO_298 (O_298,N_2676,N_2883);
or UO_299 (O_299,N_2933,N_2558);
xnor UO_300 (O_300,N_2908,N_2692);
nor UO_301 (O_301,N_2617,N_2572);
nand UO_302 (O_302,N_2934,N_2622);
nand UO_303 (O_303,N_2868,N_2830);
and UO_304 (O_304,N_2606,N_2609);
nand UO_305 (O_305,N_2718,N_2909);
nor UO_306 (O_306,N_2692,N_2859);
or UO_307 (O_307,N_2838,N_2741);
or UO_308 (O_308,N_2633,N_2639);
or UO_309 (O_309,N_2729,N_2895);
or UO_310 (O_310,N_2596,N_2775);
nand UO_311 (O_311,N_2637,N_2620);
nor UO_312 (O_312,N_2978,N_2790);
nor UO_313 (O_313,N_2999,N_2506);
nand UO_314 (O_314,N_2834,N_2810);
nor UO_315 (O_315,N_2638,N_2928);
nor UO_316 (O_316,N_2606,N_2947);
nand UO_317 (O_317,N_2757,N_2967);
and UO_318 (O_318,N_2540,N_2670);
or UO_319 (O_319,N_2839,N_2867);
and UO_320 (O_320,N_2995,N_2793);
nor UO_321 (O_321,N_2712,N_2519);
nand UO_322 (O_322,N_2930,N_2568);
xor UO_323 (O_323,N_2953,N_2944);
nand UO_324 (O_324,N_2698,N_2710);
or UO_325 (O_325,N_2675,N_2724);
nor UO_326 (O_326,N_2755,N_2981);
nand UO_327 (O_327,N_2565,N_2888);
nor UO_328 (O_328,N_2993,N_2666);
or UO_329 (O_329,N_2967,N_2703);
and UO_330 (O_330,N_2838,N_2694);
nand UO_331 (O_331,N_2587,N_2868);
nand UO_332 (O_332,N_2687,N_2700);
and UO_333 (O_333,N_2859,N_2915);
nor UO_334 (O_334,N_2916,N_2654);
xor UO_335 (O_335,N_2551,N_2871);
and UO_336 (O_336,N_2755,N_2773);
or UO_337 (O_337,N_2765,N_2981);
nand UO_338 (O_338,N_2756,N_2908);
and UO_339 (O_339,N_2715,N_2910);
nor UO_340 (O_340,N_2631,N_2937);
and UO_341 (O_341,N_2505,N_2795);
and UO_342 (O_342,N_2738,N_2906);
nor UO_343 (O_343,N_2631,N_2944);
and UO_344 (O_344,N_2743,N_2913);
nand UO_345 (O_345,N_2626,N_2551);
or UO_346 (O_346,N_2823,N_2581);
and UO_347 (O_347,N_2555,N_2636);
and UO_348 (O_348,N_2835,N_2894);
or UO_349 (O_349,N_2989,N_2826);
and UO_350 (O_350,N_2749,N_2967);
nor UO_351 (O_351,N_2620,N_2884);
nand UO_352 (O_352,N_2688,N_2694);
nor UO_353 (O_353,N_2965,N_2692);
and UO_354 (O_354,N_2839,N_2686);
nor UO_355 (O_355,N_2924,N_2706);
and UO_356 (O_356,N_2593,N_2941);
and UO_357 (O_357,N_2804,N_2584);
or UO_358 (O_358,N_2780,N_2945);
nor UO_359 (O_359,N_2757,N_2529);
nor UO_360 (O_360,N_2879,N_2637);
or UO_361 (O_361,N_2842,N_2796);
and UO_362 (O_362,N_2936,N_2894);
or UO_363 (O_363,N_2721,N_2710);
nor UO_364 (O_364,N_2518,N_2835);
nand UO_365 (O_365,N_2517,N_2999);
nand UO_366 (O_366,N_2923,N_2657);
and UO_367 (O_367,N_2694,N_2650);
nor UO_368 (O_368,N_2698,N_2614);
and UO_369 (O_369,N_2720,N_2500);
nand UO_370 (O_370,N_2646,N_2712);
or UO_371 (O_371,N_2545,N_2655);
nor UO_372 (O_372,N_2651,N_2664);
nor UO_373 (O_373,N_2652,N_2799);
and UO_374 (O_374,N_2682,N_2528);
and UO_375 (O_375,N_2830,N_2535);
and UO_376 (O_376,N_2897,N_2618);
nand UO_377 (O_377,N_2578,N_2569);
nor UO_378 (O_378,N_2863,N_2698);
and UO_379 (O_379,N_2832,N_2572);
or UO_380 (O_380,N_2690,N_2898);
and UO_381 (O_381,N_2726,N_2641);
or UO_382 (O_382,N_2856,N_2538);
nand UO_383 (O_383,N_2697,N_2897);
nand UO_384 (O_384,N_2971,N_2874);
and UO_385 (O_385,N_2973,N_2512);
or UO_386 (O_386,N_2939,N_2797);
and UO_387 (O_387,N_2951,N_2884);
nor UO_388 (O_388,N_2660,N_2997);
nor UO_389 (O_389,N_2722,N_2789);
nand UO_390 (O_390,N_2719,N_2607);
xnor UO_391 (O_391,N_2820,N_2570);
nand UO_392 (O_392,N_2540,N_2591);
nor UO_393 (O_393,N_2905,N_2968);
nand UO_394 (O_394,N_2831,N_2942);
or UO_395 (O_395,N_2863,N_2965);
or UO_396 (O_396,N_2822,N_2943);
nand UO_397 (O_397,N_2955,N_2604);
and UO_398 (O_398,N_2811,N_2762);
nand UO_399 (O_399,N_2879,N_2722);
or UO_400 (O_400,N_2702,N_2723);
nand UO_401 (O_401,N_2696,N_2519);
nand UO_402 (O_402,N_2887,N_2550);
nor UO_403 (O_403,N_2623,N_2783);
and UO_404 (O_404,N_2745,N_2776);
nor UO_405 (O_405,N_2625,N_2710);
and UO_406 (O_406,N_2507,N_2778);
nand UO_407 (O_407,N_2946,N_2701);
and UO_408 (O_408,N_2613,N_2614);
or UO_409 (O_409,N_2790,N_2519);
or UO_410 (O_410,N_2726,N_2563);
and UO_411 (O_411,N_2993,N_2958);
nand UO_412 (O_412,N_2971,N_2735);
nand UO_413 (O_413,N_2778,N_2815);
or UO_414 (O_414,N_2825,N_2614);
or UO_415 (O_415,N_2832,N_2670);
nor UO_416 (O_416,N_2965,N_2997);
nand UO_417 (O_417,N_2854,N_2876);
or UO_418 (O_418,N_2678,N_2683);
and UO_419 (O_419,N_2521,N_2799);
and UO_420 (O_420,N_2852,N_2866);
or UO_421 (O_421,N_2978,N_2957);
nand UO_422 (O_422,N_2960,N_2616);
and UO_423 (O_423,N_2609,N_2820);
nand UO_424 (O_424,N_2615,N_2746);
nor UO_425 (O_425,N_2944,N_2814);
nand UO_426 (O_426,N_2911,N_2666);
nand UO_427 (O_427,N_2963,N_2872);
and UO_428 (O_428,N_2930,N_2776);
or UO_429 (O_429,N_2860,N_2662);
and UO_430 (O_430,N_2669,N_2583);
and UO_431 (O_431,N_2999,N_2992);
and UO_432 (O_432,N_2940,N_2617);
and UO_433 (O_433,N_2533,N_2950);
xnor UO_434 (O_434,N_2653,N_2719);
or UO_435 (O_435,N_2618,N_2567);
or UO_436 (O_436,N_2711,N_2584);
and UO_437 (O_437,N_2823,N_2833);
xor UO_438 (O_438,N_2622,N_2505);
nand UO_439 (O_439,N_2851,N_2780);
nor UO_440 (O_440,N_2556,N_2532);
nor UO_441 (O_441,N_2667,N_2770);
nor UO_442 (O_442,N_2768,N_2798);
nor UO_443 (O_443,N_2610,N_2771);
nor UO_444 (O_444,N_2773,N_2541);
or UO_445 (O_445,N_2555,N_2984);
nor UO_446 (O_446,N_2755,N_2931);
nor UO_447 (O_447,N_2739,N_2947);
and UO_448 (O_448,N_2510,N_2600);
xnor UO_449 (O_449,N_2740,N_2598);
or UO_450 (O_450,N_2606,N_2894);
nor UO_451 (O_451,N_2851,N_2921);
or UO_452 (O_452,N_2857,N_2947);
or UO_453 (O_453,N_2603,N_2536);
nand UO_454 (O_454,N_2740,N_2943);
nor UO_455 (O_455,N_2997,N_2783);
nand UO_456 (O_456,N_2505,N_2916);
nor UO_457 (O_457,N_2931,N_2693);
and UO_458 (O_458,N_2706,N_2913);
nand UO_459 (O_459,N_2823,N_2641);
nor UO_460 (O_460,N_2844,N_2669);
and UO_461 (O_461,N_2561,N_2750);
nor UO_462 (O_462,N_2765,N_2884);
nand UO_463 (O_463,N_2541,N_2743);
and UO_464 (O_464,N_2570,N_2832);
or UO_465 (O_465,N_2511,N_2534);
nor UO_466 (O_466,N_2533,N_2859);
and UO_467 (O_467,N_2527,N_2799);
nor UO_468 (O_468,N_2850,N_2754);
and UO_469 (O_469,N_2698,N_2656);
and UO_470 (O_470,N_2600,N_2541);
or UO_471 (O_471,N_2702,N_2785);
or UO_472 (O_472,N_2543,N_2969);
nand UO_473 (O_473,N_2967,N_2644);
and UO_474 (O_474,N_2776,N_2759);
or UO_475 (O_475,N_2824,N_2921);
or UO_476 (O_476,N_2594,N_2619);
nor UO_477 (O_477,N_2675,N_2596);
nor UO_478 (O_478,N_2764,N_2969);
nand UO_479 (O_479,N_2811,N_2579);
nand UO_480 (O_480,N_2954,N_2588);
nand UO_481 (O_481,N_2507,N_2855);
and UO_482 (O_482,N_2675,N_2587);
nor UO_483 (O_483,N_2588,N_2768);
or UO_484 (O_484,N_2833,N_2709);
or UO_485 (O_485,N_2525,N_2738);
or UO_486 (O_486,N_2510,N_2782);
or UO_487 (O_487,N_2668,N_2985);
nand UO_488 (O_488,N_2975,N_2683);
nor UO_489 (O_489,N_2653,N_2866);
nor UO_490 (O_490,N_2914,N_2650);
or UO_491 (O_491,N_2880,N_2640);
or UO_492 (O_492,N_2732,N_2530);
or UO_493 (O_493,N_2786,N_2651);
or UO_494 (O_494,N_2632,N_2940);
and UO_495 (O_495,N_2982,N_2932);
and UO_496 (O_496,N_2586,N_2971);
and UO_497 (O_497,N_2984,N_2910);
nor UO_498 (O_498,N_2623,N_2611);
nor UO_499 (O_499,N_2595,N_2501);
endmodule