module basic_1500_15000_2000_75_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_285,In_1390);
nor U1 (N_1,In_8,In_1410);
and U2 (N_2,In_1159,In_1278);
nor U3 (N_3,In_62,In_1258);
xor U4 (N_4,In_122,In_637);
nor U5 (N_5,In_348,In_469);
nor U6 (N_6,In_118,In_899);
and U7 (N_7,In_1094,In_464);
or U8 (N_8,In_1270,In_289);
nor U9 (N_9,In_935,In_384);
xnor U10 (N_10,In_956,In_1380);
or U11 (N_11,In_1028,In_1020);
and U12 (N_12,In_23,In_372);
nand U13 (N_13,In_914,In_810);
nand U14 (N_14,In_25,In_1375);
nor U15 (N_15,In_1205,In_1301);
and U16 (N_16,In_107,In_37);
or U17 (N_17,In_1180,In_1470);
and U18 (N_18,In_1243,In_1035);
or U19 (N_19,In_1150,In_772);
nand U20 (N_20,In_214,In_254);
xnor U21 (N_21,In_120,In_79);
or U22 (N_22,In_425,In_243);
xnor U23 (N_23,In_19,In_476);
xnor U24 (N_24,In_445,In_465);
nor U25 (N_25,In_1490,In_1385);
xor U26 (N_26,In_178,In_724);
nand U27 (N_27,In_101,In_752);
and U28 (N_28,In_433,In_435);
and U29 (N_29,In_807,In_1255);
and U30 (N_30,In_437,In_987);
xor U31 (N_31,In_738,In_1177);
nand U32 (N_32,In_1108,In_357);
or U33 (N_33,In_121,In_351);
nor U34 (N_34,In_96,In_216);
and U35 (N_35,In_74,In_554);
or U36 (N_36,In_809,In_683);
xnor U37 (N_37,In_1325,In_570);
xor U38 (N_38,In_561,In_538);
xnor U39 (N_39,In_1396,In_184);
or U40 (N_40,In_1169,In_1224);
and U41 (N_41,In_1005,In_166);
nand U42 (N_42,In_658,In_1452);
nor U43 (N_43,In_1382,In_1154);
xnor U44 (N_44,In_207,In_1140);
or U45 (N_45,In_479,In_547);
and U46 (N_46,In_495,In_1231);
nand U47 (N_47,In_1336,In_453);
xnor U48 (N_48,In_1013,In_599);
xor U49 (N_49,In_280,In_135);
nand U50 (N_50,In_1326,In_584);
and U51 (N_51,In_848,In_632);
nand U52 (N_52,In_317,In_603);
and U53 (N_53,In_201,In_405);
nand U54 (N_54,In_410,In_1081);
xnor U55 (N_55,In_1304,In_1040);
nor U56 (N_56,In_869,In_151);
nand U57 (N_57,In_705,In_106);
and U58 (N_58,In_635,In_1473);
nor U59 (N_59,In_237,In_936);
nand U60 (N_60,In_607,In_394);
and U61 (N_61,In_1386,In_981);
nor U62 (N_62,In_1161,In_877);
xor U63 (N_63,In_979,In_845);
xnor U64 (N_64,In_745,In_1234);
or U65 (N_65,In_10,In_268);
xor U66 (N_66,In_1026,In_910);
and U67 (N_67,In_198,In_99);
nand U68 (N_68,In_229,In_879);
nand U69 (N_69,In_939,In_1277);
xor U70 (N_70,In_729,In_620);
or U71 (N_71,In_4,In_1210);
nor U72 (N_72,In_466,In_1455);
xor U73 (N_73,In_129,In_903);
nand U74 (N_74,In_245,In_741);
and U75 (N_75,In_639,In_1105);
and U76 (N_76,In_130,In_842);
nand U77 (N_77,In_292,In_1459);
and U78 (N_78,In_827,In_1126);
xnor U79 (N_79,In_1055,In_385);
and U80 (N_80,In_1286,In_168);
nand U81 (N_81,In_81,In_139);
nor U82 (N_82,In_1297,In_1249);
xor U83 (N_83,In_1497,In_1416);
nor U84 (N_84,In_962,In_596);
nand U85 (N_85,In_984,In_391);
xnor U86 (N_86,In_1137,In_463);
xor U87 (N_87,In_559,In_1010);
nor U88 (N_88,In_978,In_1285);
and U89 (N_89,In_224,In_1139);
xor U90 (N_90,In_21,In_1246);
xor U91 (N_91,In_1371,In_155);
nand U92 (N_92,In_258,In_1064);
nor U93 (N_93,In_206,In_36);
nand U94 (N_94,In_997,In_446);
and U95 (N_95,In_393,In_713);
xnor U96 (N_96,In_998,In_1495);
or U97 (N_97,In_1148,In_17);
and U98 (N_98,In_1025,In_419);
nor U99 (N_99,In_860,In_544);
and U100 (N_100,In_18,In_1237);
and U101 (N_101,In_146,In_1412);
xnor U102 (N_102,In_261,In_449);
nand U103 (N_103,In_91,In_1118);
nor U104 (N_104,In_450,In_595);
and U105 (N_105,In_109,In_167);
xor U106 (N_106,In_92,In_600);
nand U107 (N_107,In_43,In_376);
xnor U108 (N_108,In_1049,In_1492);
nor U109 (N_109,In_926,In_1404);
nand U110 (N_110,In_1256,In_363);
xnor U111 (N_111,In_916,In_1075);
nand U112 (N_112,In_325,In_725);
and U113 (N_113,In_698,In_440);
and U114 (N_114,In_474,In_455);
nor U115 (N_115,In_761,In_1117);
and U116 (N_116,In_1349,In_1310);
nor U117 (N_117,In_1352,In_1467);
nand U118 (N_118,In_271,In_780);
nor U119 (N_119,In_182,In_753);
and U120 (N_120,In_1288,In_555);
and U121 (N_121,In_988,In_861);
nand U122 (N_122,In_347,In_950);
and U123 (N_123,In_170,In_1024);
xor U124 (N_124,In_190,In_886);
or U125 (N_125,In_248,In_526);
or U126 (N_126,In_884,In_30);
or U127 (N_127,In_160,In_1446);
or U128 (N_128,In_1052,In_5);
nand U129 (N_129,In_806,In_335);
or U130 (N_130,In_576,In_1319);
or U131 (N_131,In_204,In_1238);
and U132 (N_132,In_684,In_647);
xor U133 (N_133,In_1261,In_579);
or U134 (N_134,In_605,In_768);
nor U135 (N_135,In_965,In_550);
or U136 (N_136,In_623,In_1187);
or U137 (N_137,In_378,In_720);
or U138 (N_138,In_704,In_868);
xor U139 (N_139,In_390,In_1147);
nor U140 (N_140,In_1477,In_734);
or U141 (N_141,In_718,In_609);
nor U142 (N_142,In_706,In_218);
nand U143 (N_143,In_699,In_1109);
and U144 (N_144,In_294,In_203);
and U145 (N_145,In_850,In_119);
nand U146 (N_146,In_627,In_1122);
or U147 (N_147,In_814,In_368);
nor U148 (N_148,In_478,In_908);
and U149 (N_149,In_1134,In_661);
xor U150 (N_150,In_374,In_485);
xor U151 (N_151,In_164,In_568);
or U152 (N_152,In_1207,In_117);
or U153 (N_153,In_1044,In_1219);
or U154 (N_154,In_755,In_1327);
nor U155 (N_155,In_171,In_1119);
xor U156 (N_156,In_140,In_24);
nor U157 (N_157,In_1209,In_1287);
xnor U158 (N_158,In_1215,In_187);
or U159 (N_159,In_836,In_161);
and U160 (N_160,In_1340,In_928);
or U161 (N_161,In_11,In_77);
and U162 (N_162,In_1398,In_516);
and U163 (N_163,In_165,In_1115);
xnor U164 (N_164,In_442,In_159);
or U165 (N_165,In_883,In_176);
nand U166 (N_166,In_833,In_341);
nor U167 (N_167,In_1206,In_675);
nand U168 (N_168,In_138,In_227);
or U169 (N_169,In_219,In_687);
nor U170 (N_170,In_361,In_483);
and U171 (N_171,In_1351,In_1014);
and U172 (N_172,In_33,In_1050);
and U173 (N_173,In_1103,In_940);
nor U174 (N_174,In_1464,In_714);
nand U175 (N_175,In_918,In_583);
xor U176 (N_176,In_668,In_1242);
and U177 (N_177,In_486,In_1063);
and U178 (N_178,In_86,In_1156);
nor U179 (N_179,In_749,In_403);
and U180 (N_180,In_512,In_530);
nand U181 (N_181,In_1008,In_1107);
or U182 (N_182,In_856,In_970);
nor U183 (N_183,In_580,In_352);
xnor U184 (N_184,In_1053,In_1083);
nor U185 (N_185,In_626,In_934);
nand U186 (N_186,In_269,In_489);
and U187 (N_187,In_959,In_641);
xor U188 (N_188,In_221,In_1273);
nand U189 (N_189,In_298,In_1415);
xnor U190 (N_190,In_1370,In_1060);
nor U191 (N_191,In_175,In_947);
nor U192 (N_192,In_1068,In_710);
or U193 (N_193,In_148,In_452);
nand U194 (N_194,In_222,In_1182);
nor U195 (N_195,In_1337,In_894);
nor U196 (N_196,In_983,In_125);
xnor U197 (N_197,In_1476,In_1401);
and U198 (N_198,In_1399,In_1172);
or U199 (N_199,In_1474,In_931);
nand U200 (N_200,N_37,In_905);
xor U201 (N_201,In_284,In_158);
nor U202 (N_202,In_1289,In_27);
nand U203 (N_203,In_327,In_1096);
xor U204 (N_204,N_183,N_58);
nor U205 (N_205,In_231,In_765);
or U206 (N_206,In_515,N_23);
nand U207 (N_207,In_996,N_89);
nand U208 (N_208,In_1491,In_177);
nor U209 (N_209,In_270,In_228);
or U210 (N_210,In_97,In_304);
nand U211 (N_211,N_48,In_186);
xor U212 (N_212,In_737,In_678);
nor U213 (N_213,In_286,In_262);
and U214 (N_214,In_472,In_392);
xor U215 (N_215,In_264,In_1221);
and U216 (N_216,In_290,In_703);
and U217 (N_217,In_157,In_993);
or U218 (N_218,In_239,In_565);
and U219 (N_219,In_813,In_1127);
and U220 (N_220,In_542,In_758);
and U221 (N_221,In_840,In_1051);
nor U222 (N_222,In_723,In_46);
nand U223 (N_223,In_712,In_42);
or U224 (N_224,In_497,In_1485);
xnor U225 (N_225,In_975,In_1208);
nand U226 (N_226,In_1007,In_147);
nand U227 (N_227,N_148,In_1358);
nor U228 (N_228,In_977,In_1295);
nor U229 (N_229,In_1070,In_417);
or U230 (N_230,In_1489,In_1157);
xor U231 (N_231,In_309,In_67);
nand U232 (N_232,In_451,In_898);
or U233 (N_233,N_50,In_334);
or U234 (N_234,N_79,In_1417);
and U235 (N_235,In_514,In_112);
xor U236 (N_236,In_503,In_383);
nand U237 (N_237,In_921,In_951);
nand U238 (N_238,N_62,In_481);
nand U239 (N_239,In_509,N_177);
or U240 (N_240,In_132,In_1091);
nor U241 (N_241,In_851,In_517);
nand U242 (N_242,In_45,In_1003);
nor U243 (N_243,In_913,In_1447);
and U244 (N_244,In_828,In_342);
nand U245 (N_245,In_823,In_35);
nor U246 (N_246,In_400,In_1283);
xor U247 (N_247,In_566,In_982);
and U248 (N_248,In_1197,In_257);
or U249 (N_249,In_930,In_1403);
nor U250 (N_250,In_448,In_240);
or U251 (N_251,In_1136,In_625);
xnor U252 (N_252,In_211,In_1056);
xor U253 (N_253,In_777,N_139);
and U254 (N_254,N_130,In_591);
and U255 (N_255,N_74,In_799);
or U256 (N_256,In_890,In_735);
or U257 (N_257,In_1184,In_1343);
xnor U258 (N_258,In_1213,In_1259);
nand U259 (N_259,In_1484,In_266);
or U260 (N_260,In_246,N_51);
nor U261 (N_261,In_1240,In_1226);
nor U262 (N_262,In_610,N_196);
nand U263 (N_263,In_907,In_1335);
or U264 (N_264,In_598,N_149);
xnor U265 (N_265,In_379,N_103);
and U266 (N_266,In_1482,N_119);
and U267 (N_267,In_980,In_1178);
xnor U268 (N_268,In_436,In_84);
xnor U269 (N_269,In_142,In_1338);
and U270 (N_270,N_6,In_1479);
nand U271 (N_271,In_128,In_69);
nor U272 (N_272,In_1293,In_1284);
or U273 (N_273,In_312,N_91);
and U274 (N_274,In_1407,In_316);
or U275 (N_275,In_532,In_1279);
and U276 (N_276,In_336,In_657);
nand U277 (N_277,In_708,In_671);
xnor U278 (N_278,In_917,In_212);
xnor U279 (N_279,In_1229,In_1394);
and U280 (N_280,In_1100,N_88);
nor U281 (N_281,In_60,In_195);
xor U282 (N_282,In_1457,In_937);
nor U283 (N_283,In_1430,In_1406);
or U284 (N_284,In_1162,In_876);
xnor U285 (N_285,In_617,In_1130);
nor U286 (N_286,In_1376,In_776);
and U287 (N_287,In_225,In_13);
nand U288 (N_288,In_1269,In_344);
or U289 (N_289,N_185,In_295);
and U290 (N_290,In_781,In_785);
nor U291 (N_291,In_518,In_945);
xor U292 (N_292,In_1186,In_1202);
nor U293 (N_293,In_1441,In_1395);
xnor U294 (N_294,In_1369,In_622);
and U295 (N_295,In_665,In_1129);
or U296 (N_296,In_1361,In_1264);
and U297 (N_297,N_152,In_1423);
and U298 (N_298,In_577,In_679);
xnor U299 (N_299,In_674,N_169);
xor U300 (N_300,In_646,In_540);
nand U301 (N_301,N_57,In_456);
and U302 (N_302,In_731,In_636);
and U303 (N_303,In_1333,In_1036);
nor U304 (N_304,In_797,In_867);
or U305 (N_305,In_1414,In_193);
nand U306 (N_306,In_923,In_739);
nand U307 (N_307,In_792,N_186);
or U308 (N_308,In_1329,In_1006);
or U309 (N_309,In_1313,In_841);
and U310 (N_310,N_41,In_1176);
nand U311 (N_311,N_197,In_302);
nand U312 (N_312,N_161,In_1276);
or U313 (N_313,In_644,In_502);
xor U314 (N_314,In_901,In_162);
nor U315 (N_315,In_621,In_1453);
nor U316 (N_316,In_126,In_188);
nand U317 (N_317,In_424,In_685);
or U318 (N_318,In_1165,N_135);
xor U319 (N_319,In_1280,N_122);
nand U320 (N_320,In_1469,In_1015);
nand U321 (N_321,In_832,In_1179);
or U322 (N_322,N_132,N_78);
or U323 (N_323,In_733,In_1450);
nand U324 (N_324,In_629,In_1373);
nor U325 (N_325,In_366,In_1486);
nor U326 (N_326,N_190,In_427);
nand U327 (N_327,In_1065,In_594);
nor U328 (N_328,In_938,In_447);
or U329 (N_329,N_26,N_158);
nor U330 (N_330,In_1451,In_137);
nor U331 (N_331,In_273,In_766);
xnor U332 (N_332,In_1468,In_1223);
nor U333 (N_333,In_47,In_1043);
xor U334 (N_334,In_1124,N_101);
xor U335 (N_335,In_1042,In_1123);
xor U336 (N_336,N_80,N_81);
and U337 (N_337,In_1445,In_202);
nand U338 (N_338,In_149,In_858);
nand U339 (N_339,In_1381,In_324);
or U340 (N_340,N_109,In_356);
or U341 (N_341,In_1321,In_1438);
or U342 (N_342,In_242,In_215);
and U343 (N_343,N_189,In_533);
and U344 (N_344,N_44,In_722);
or U345 (N_345,In_1436,In_200);
and U346 (N_346,In_457,In_1334);
and U347 (N_347,In_721,N_164);
nand U348 (N_348,In_499,In_396);
or U349 (N_349,In_1443,In_656);
xnor U350 (N_350,In_287,In_608);
nor U351 (N_351,In_727,In_783);
nor U352 (N_352,N_166,N_159);
xor U353 (N_353,N_70,In_55);
xnor U354 (N_354,In_369,In_1188);
nand U355 (N_355,In_1151,In_83);
nand U356 (N_356,In_172,In_545);
nor U357 (N_357,N_170,In_300);
xor U358 (N_358,In_1323,In_1183);
or U359 (N_359,In_1377,In_1413);
nor U360 (N_360,In_1252,In_551);
or U361 (N_361,In_253,N_75);
xnor U362 (N_362,In_364,N_104);
nor U363 (N_363,In_278,In_1324);
nor U364 (N_364,In_1408,In_866);
nor U365 (N_365,In_587,In_895);
nand U366 (N_366,In_527,N_155);
nand U367 (N_367,In_920,In_655);
xnor U368 (N_368,In_795,In_885);
and U369 (N_369,In_1047,N_76);
nor U370 (N_370,In_428,In_412);
xor U371 (N_371,In_585,In_838);
and U372 (N_372,In_811,In_1409);
nor U373 (N_373,In_902,In_1348);
xor U374 (N_374,In_1120,In_602);
and U375 (N_375,N_11,In_249);
and U376 (N_376,N_138,In_1031);
xor U377 (N_377,N_118,N_4);
nor U378 (N_378,In_1095,In_941);
nand U379 (N_379,In_943,In_520);
xor U380 (N_380,In_770,In_794);
or U381 (N_381,In_1090,N_144);
and U382 (N_382,In_1461,In_460);
xnor U383 (N_383,In_51,In_401);
nand U384 (N_384,In_32,In_893);
nand U385 (N_385,In_1316,In_693);
nor U386 (N_386,In_1191,N_100);
and U387 (N_387,In_1203,In_728);
or U388 (N_388,In_471,N_60);
xor U389 (N_389,In_65,In_990);
and U390 (N_390,In_1367,In_480);
xnor U391 (N_391,In_1102,In_677);
and U392 (N_392,In_429,In_1425);
nand U393 (N_393,In_1037,In_462);
and U394 (N_394,In_1201,In_467);
xnor U395 (N_395,In_697,In_649);
and U396 (N_396,In_34,N_66);
or U397 (N_397,In_616,In_28);
nand U398 (N_398,In_853,In_992);
xnor U399 (N_399,In_434,In_1434);
nor U400 (N_400,In_1366,N_117);
nor U401 (N_401,N_35,N_303);
xor U402 (N_402,N_5,In_812);
or U403 (N_403,In_1086,In_277);
nor U404 (N_404,In_1355,In_1142);
or U405 (N_405,In_1168,In_1078);
or U406 (N_406,In_1158,N_294);
nand U407 (N_407,In_265,In_1294);
and U408 (N_408,N_178,In_89);
or U409 (N_409,In_57,In_6);
or U410 (N_410,N_291,In_1239);
xnor U411 (N_411,In_606,In_952);
or U412 (N_412,In_1125,N_53);
nor U413 (N_413,In_473,N_350);
nor U414 (N_414,N_8,N_237);
nor U415 (N_415,In_863,N_38);
xor U416 (N_416,In_38,N_46);
xor U417 (N_417,N_56,In_750);
nand U418 (N_418,In_673,N_389);
or U419 (N_419,In_1302,In_872);
nor U420 (N_420,N_345,In_64);
nor U421 (N_421,In_331,In_522);
nand U422 (N_422,N_10,In_404);
xnor U423 (N_423,N_388,In_328);
xnor U424 (N_424,In_645,In_946);
or U425 (N_425,In_310,In_326);
or U426 (N_426,In_333,N_259);
or U427 (N_427,In_778,In_1462);
or U428 (N_428,In_844,In_1439);
nand U429 (N_429,In_826,N_110);
nor U430 (N_430,In_1093,In_1077);
and U431 (N_431,In_686,N_250);
xor U432 (N_432,In_651,In_1496);
xnor U433 (N_433,N_142,N_200);
xor U434 (N_434,N_374,In_299);
or U435 (N_435,In_662,N_198);
and U436 (N_436,In_791,N_64);
and U437 (N_437,N_173,N_199);
xor U438 (N_438,In_653,In_556);
nand U439 (N_439,N_372,In_912);
or U440 (N_440,N_378,In_694);
or U441 (N_441,N_77,In_422);
xor U442 (N_442,N_364,N_204);
nand U443 (N_443,In_100,In_767);
xnor U444 (N_444,In_53,In_443);
or U445 (N_445,In_1076,N_324);
xnor U446 (N_446,In_1073,N_396);
xor U447 (N_447,In_371,In_470);
nor U448 (N_448,In_1164,N_307);
and U449 (N_449,N_279,N_330);
nor U450 (N_450,In_628,N_329);
nand U451 (N_451,N_249,In_573);
nand U452 (N_452,In_1017,In_438);
nor U453 (N_453,In_272,In_500);
and U454 (N_454,N_341,In_973);
nand U455 (N_455,N_293,In_747);
xnor U456 (N_456,N_224,In_49);
nor U457 (N_457,In_1475,In_717);
xor U458 (N_458,In_995,In_388);
nand U459 (N_459,In_1347,N_131);
xnor U460 (N_460,N_182,N_243);
nand U461 (N_461,In_815,N_42);
xnor U462 (N_462,In_1163,In_1089);
nand U463 (N_463,In_971,N_3);
nor U464 (N_464,N_271,In_571);
nand U465 (N_465,N_15,In_244);
or U466 (N_466,In_589,N_277);
and U467 (N_467,In_798,N_40);
nand U468 (N_468,In_967,N_59);
nand U469 (N_469,In_1384,N_32);
and U470 (N_470,In_553,In_543);
nor U471 (N_471,In_624,N_205);
xnor U472 (N_472,In_1392,In_835);
nor U473 (N_473,In_274,In_241);
and U474 (N_474,In_362,N_241);
nand U475 (N_475,N_227,N_240);
nor U476 (N_476,In_927,In_839);
or U477 (N_477,In_256,In_1391);
nor U478 (N_478,N_298,In_702);
xor U479 (N_479,In_7,In_381);
nand U480 (N_480,In_169,In_1146);
nand U481 (N_481,N_112,In_426);
and U482 (N_482,In_790,In_1303);
or U483 (N_483,In_779,In_76);
nand U484 (N_484,In_1248,In_972);
or U485 (N_485,In_1250,In_746);
or U486 (N_486,In_654,In_1192);
nand U487 (N_487,In_1431,In_1067);
nor U488 (N_488,In_830,N_383);
nand U489 (N_489,N_73,In_402);
nand U490 (N_490,In_942,N_107);
nand U491 (N_491,N_172,N_54);
nand U492 (N_492,In_865,N_358);
nor U493 (N_493,In_1212,In_209);
or U494 (N_494,In_1041,N_349);
nand U495 (N_495,N_102,In_822);
or U496 (N_496,In_1200,N_0);
xor U497 (N_497,In_275,In_323);
nor U498 (N_498,In_680,N_165);
nand U499 (N_499,In_1141,In_1198);
or U500 (N_500,N_269,In_1171);
xnor U501 (N_501,N_284,In_888);
nor U502 (N_502,In_578,In_513);
xor U503 (N_503,N_30,N_275);
and U504 (N_504,N_242,In_986);
and U505 (N_505,N_226,In_689);
or U506 (N_506,N_43,In_769);
xnor U507 (N_507,In_744,N_251);
and U508 (N_508,N_267,In_370);
and U509 (N_509,In_1345,In_1220);
and U510 (N_510,In_534,N_233);
nor U511 (N_511,N_136,In_131);
xor U512 (N_512,In_196,In_181);
nor U513 (N_513,N_116,In_1356);
nand U514 (N_514,In_1266,In_191);
or U515 (N_515,In_1499,In_618);
nand U516 (N_516,In_1079,In_1307);
xor U517 (N_517,In_1272,In_1131);
nand U518 (N_518,In_1435,In_1332);
or U519 (N_519,N_206,In_441);
or U520 (N_520,N_362,In_1383);
or U521 (N_521,N_235,In_1465);
nand U522 (N_522,N_367,In_805);
or U523 (N_523,In_817,In_260);
xnor U524 (N_524,In_726,In_818);
nor U525 (N_525,In_613,In_743);
nor U526 (N_526,In_296,N_72);
xnor U527 (N_527,In_1016,In_802);
nand U528 (N_528,N_1,In_1216);
xnor U529 (N_529,In_896,N_108);
and U530 (N_530,N_137,In_1048);
xnor U531 (N_531,In_144,In_961);
nand U532 (N_532,In_1251,In_418);
xnor U533 (N_533,In_1331,N_22);
xnor U534 (N_534,In_41,In_199);
or U535 (N_535,In_682,In_345);
xnor U536 (N_536,In_994,In_1344);
nor U537 (N_537,In_281,In_90);
nor U538 (N_538,In_1298,In_1493);
xnor U539 (N_539,N_92,N_268);
nor U540 (N_540,In_1471,In_669);
nor U541 (N_541,In_1339,In_1113);
nand U542 (N_542,N_71,In_338);
xor U543 (N_543,In_1145,In_407);
xnor U544 (N_544,N_248,In_85);
or U545 (N_545,In_1472,In_964);
xnor U546 (N_546,N_333,In_39);
or U547 (N_547,In_377,In_44);
xor U548 (N_548,In_133,N_339);
nor U549 (N_549,N_391,N_212);
xnor U550 (N_550,In_355,In_380);
nand U551 (N_551,In_1022,N_29);
xnor U552 (N_552,In_1084,In_1357);
nand U553 (N_553,In_1442,In_1128);
and U554 (N_554,In_1133,N_318);
xor U555 (N_555,In_948,In_1085);
xor U556 (N_556,In_871,N_145);
nand U557 (N_557,In_420,N_246);
and U558 (N_558,In_1166,N_278);
nor U559 (N_559,In_1038,N_338);
and U560 (N_560,In_163,In_1444);
nand U561 (N_561,N_25,In_1483);
xor U562 (N_562,N_386,N_288);
nand U563 (N_563,In_688,N_39);
xor U564 (N_564,In_1420,In_506);
nor U565 (N_565,In_1218,In_963);
nor U566 (N_566,In_72,N_353);
nor U567 (N_567,N_263,In_524);
xnor U568 (N_568,In_763,In_1481);
nand U569 (N_569,In_397,In_870);
nand U570 (N_570,In_444,In_659);
nor U571 (N_571,N_24,In_1000);
nand U572 (N_572,N_18,In_824);
nand U573 (N_573,N_295,In_382);
and U574 (N_574,In_1466,N_192);
or U575 (N_575,In_696,In_1267);
nor U576 (N_576,In_619,N_346);
nand U577 (N_577,In_634,N_302);
or U578 (N_578,N_310,N_114);
and U579 (N_579,N_225,In_786);
or U580 (N_580,In_1426,In_652);
or U581 (N_581,N_157,N_133);
nor U582 (N_582,In_291,In_1312);
and U583 (N_583,In_762,In_1299);
nand U584 (N_584,In_1149,N_384);
and U585 (N_585,In_663,In_528);
and U586 (N_586,N_219,In_643);
xnor U587 (N_587,In_124,In_1135);
xor U588 (N_588,N_211,In_771);
or U589 (N_589,In_314,In_759);
or U590 (N_590,In_1082,N_201);
xor U591 (N_591,In_796,In_1241);
nor U592 (N_592,In_1454,N_292);
or U593 (N_593,In_1106,In_173);
nor U594 (N_594,In_421,In_1235);
nand U595 (N_595,In_592,In_329);
nor U596 (N_596,In_1092,In_375);
nor U597 (N_597,N_322,In_1045);
or U598 (N_598,In_922,N_93);
and U599 (N_599,N_65,In_874);
nand U600 (N_600,In_1363,In_523);
nand U601 (N_601,N_584,In_1232);
nand U602 (N_602,N_504,In_507);
xor U603 (N_603,N_598,In_78);
nand U604 (N_604,N_257,In_113);
or U605 (N_605,In_306,N_426);
and U606 (N_606,N_516,N_528);
xor U607 (N_607,In_567,N_52);
nand U608 (N_608,In_102,In_1488);
nand U609 (N_609,N_85,In_1368);
xnor U610 (N_610,In_1315,In_881);
nor U611 (N_611,In_1111,N_427);
nor U612 (N_612,In_431,N_168);
nor U613 (N_613,N_281,In_552);
and U614 (N_614,N_481,In_1228);
nand U615 (N_615,In_1194,In_75);
xnor U616 (N_616,In_1405,N_409);
nor U617 (N_617,In_736,In_582);
xor U618 (N_618,In_332,In_1300);
or U619 (N_619,N_524,In_966);
and U620 (N_620,In_414,In_1257);
xor U621 (N_621,N_449,N_83);
nand U622 (N_622,In_681,N_381);
and U623 (N_623,In_482,In_1456);
nor U624 (N_624,In_408,In_297);
and U625 (N_625,In_707,In_61);
xor U626 (N_626,N_213,In_29);
nor U627 (N_627,N_45,In_255);
and U628 (N_628,N_540,In_288);
nand U629 (N_629,In_230,N_289);
nand U630 (N_630,N_304,N_124);
or U631 (N_631,N_332,N_405);
and U632 (N_632,In_197,In_932);
or U633 (N_633,N_547,In_700);
nor U634 (N_634,N_262,In_423);
or U635 (N_635,N_340,N_412);
xnor U636 (N_636,In_588,N_285);
or U637 (N_637,N_121,N_489);
and U638 (N_638,N_484,In_929);
xor U639 (N_639,N_425,In_127);
or U640 (N_640,N_238,In_1071);
and U641 (N_641,In_944,N_223);
nand U642 (N_642,In_843,In_968);
nand U643 (N_643,In_194,N_184);
nor U644 (N_644,N_556,In_816);
nand U645 (N_645,In_1227,In_360);
or U646 (N_646,In_233,In_103);
xor U647 (N_647,N_361,N_296);
or U648 (N_648,In_1027,N_244);
and U649 (N_649,N_585,In_398);
xnor U650 (N_650,In_1110,N_413);
nor U651 (N_651,In_1254,N_573);
xor U652 (N_652,N_67,N_548);
and U653 (N_653,In_1360,In_354);
xor U654 (N_654,In_574,In_716);
nor U655 (N_655,In_143,N_297);
xnor U656 (N_656,N_216,N_210);
xor U657 (N_657,In_690,In_1104);
xnor U658 (N_658,N_258,N_97);
nor U659 (N_659,N_230,N_402);
nand U660 (N_660,In_251,In_640);
and U661 (N_661,N_188,In_223);
or U662 (N_662,In_40,In_95);
xnor U663 (N_663,In_638,In_58);
xor U664 (N_664,In_1291,In_1247);
xor U665 (N_665,In_68,N_400);
nand U666 (N_666,In_1217,N_582);
xor U667 (N_667,In_1018,N_126);
nor U668 (N_668,In_1012,In_145);
nor U669 (N_669,In_1342,N_436);
nor U670 (N_670,N_520,N_510);
nand U671 (N_671,In_232,In_581);
xnor U672 (N_672,N_570,N_473);
nand U673 (N_673,In_315,In_56);
and U674 (N_674,N_589,In_1155);
and U675 (N_675,In_667,N_379);
xnor U676 (N_676,In_154,N_496);
and U677 (N_677,N_160,In_508);
or U678 (N_678,N_220,In_1112);
nand U679 (N_679,In_715,In_1328);
xor U680 (N_680,N_502,In_732);
or U681 (N_681,N_492,N_467);
nand U682 (N_682,In_1072,N_90);
nor U683 (N_683,N_475,In_493);
and U684 (N_684,N_369,N_515);
and U685 (N_685,In_925,In_1244);
nor U686 (N_686,In_189,N_401);
xor U687 (N_687,In_672,N_562);
nor U688 (N_688,In_1374,In_153);
nor U689 (N_689,N_208,N_416);
xor U690 (N_690,N_355,In_701);
or U691 (N_691,In_247,In_12);
xor U692 (N_692,N_513,In_1153);
xor U693 (N_693,In_1069,N_529);
xnor U694 (N_694,N_522,In_283);
xnor U695 (N_695,N_193,N_343);
or U696 (N_696,In_477,N_382);
nand U697 (N_697,N_406,N_443);
nor U698 (N_698,N_534,In_1309);
xor U699 (N_699,In_510,In_1253);
nor U700 (N_700,In_1290,In_1074);
and U701 (N_701,N_577,N_99);
nor U702 (N_702,In_650,N_61);
and U703 (N_703,N_435,N_229);
nand U704 (N_704,In_1167,In_1292);
or U705 (N_705,N_156,In_305);
nor U706 (N_706,In_1054,In_748);
or U707 (N_707,N_334,N_519);
and U708 (N_708,In_1,In_590);
nor U709 (N_709,In_491,N_571);
and U710 (N_710,In_614,In_1029);
nand U711 (N_711,In_192,In_906);
or U712 (N_712,In_1062,In_855);
nand U713 (N_713,In_820,In_531);
or U714 (N_714,N_477,In_340);
or U715 (N_715,In_924,In_676);
nand U716 (N_716,In_666,N_373);
or U717 (N_717,N_253,In_1478);
xor U718 (N_718,N_228,In_293);
or U719 (N_719,In_949,In_803);
xor U720 (N_720,In_969,In_1144);
nor U721 (N_721,In_1306,In_1023);
nand U722 (N_722,In_1138,In_359);
or U723 (N_723,In_71,In_226);
xor U724 (N_724,N_495,N_256);
nor U725 (N_725,In_54,In_111);
and U726 (N_726,In_557,N_55);
xnor U727 (N_727,In_711,N_320);
or U728 (N_728,N_583,In_900);
xor U729 (N_729,N_479,In_307);
or U730 (N_730,In_1114,In_330);
or U731 (N_731,N_575,N_12);
nand U732 (N_732,In_648,N_453);
xnor U733 (N_733,In_16,In_461);
nand U734 (N_734,In_496,N_415);
xor U735 (N_735,N_526,N_459);
and U736 (N_736,In_536,N_94);
or U737 (N_737,N_47,In_873);
or U738 (N_738,In_1143,N_264);
nor U739 (N_739,In_1397,N_335);
xor U740 (N_740,N_163,N_596);
and U741 (N_741,N_375,In_115);
nand U742 (N_742,N_221,N_505);
xnor U743 (N_743,N_586,In_9);
nand U744 (N_744,N_20,In_415);
nor U745 (N_745,N_460,N_446);
xnor U746 (N_746,In_358,N_214);
or U747 (N_747,In_597,In_2);
xnor U748 (N_748,In_958,N_218);
xor U749 (N_749,In_1199,N_16);
xor U750 (N_750,N_404,In_1039);
xor U751 (N_751,In_1317,In_234);
nor U752 (N_752,N_448,In_1314);
nor U753 (N_753,In_311,N_499);
or U754 (N_754,In_572,N_521);
nand U755 (N_755,N_115,In_1236);
or U756 (N_756,N_87,N_565);
nand U757 (N_757,In_1372,N_555);
xor U758 (N_758,In_1245,N_327);
nand U759 (N_759,N_500,N_317);
nand U760 (N_760,In_954,In_821);
and U761 (N_761,In_308,In_740);
nor U762 (N_762,N_518,In_549);
nor U763 (N_763,N_506,In_1274);
nand U764 (N_764,In_59,In_782);
or U765 (N_765,In_252,In_156);
or U766 (N_766,In_695,N_597);
xnor U767 (N_767,In_1440,In_1009);
and U768 (N_768,In_541,In_208);
or U769 (N_769,N_377,In_563);
nand U770 (N_770,N_28,In_1196);
xnor U771 (N_771,In_1189,In_955);
xnor U772 (N_772,N_273,N_403);
or U773 (N_773,In_494,In_801);
nor U774 (N_774,In_1058,In_800);
and U775 (N_775,In_365,In_238);
xnor U776 (N_776,In_459,In_846);
or U777 (N_777,N_363,In_1387);
nand U778 (N_778,In_1389,N_113);
or U779 (N_779,N_527,In_1379);
nor U780 (N_780,In_664,In_389);
xnor U781 (N_781,In_691,N_414);
nor U782 (N_782,N_95,N_398);
or U783 (N_783,N_517,N_395);
xor U784 (N_784,In_593,N_328);
and U785 (N_785,In_775,In_1318);
nor U786 (N_786,N_9,In_1088);
xor U787 (N_787,In_789,In_1320);
and U788 (N_788,In_1214,N_123);
nor U789 (N_789,N_111,In_784);
nand U790 (N_790,N_411,In_892);
or U791 (N_791,In_313,In_82);
nor U792 (N_792,N_252,N_490);
and U793 (N_793,N_471,In_991);
nor U794 (N_794,N_559,N_394);
xor U795 (N_795,In_586,N_433);
and U796 (N_796,In_1004,In_1099);
nor U797 (N_797,N_444,In_754);
nor U798 (N_798,In_1341,N_106);
and U799 (N_799,In_1204,In_709);
and U800 (N_800,In_1116,N_668);
nor U801 (N_801,N_301,In_498);
or U802 (N_802,N_483,N_311);
and U803 (N_803,N_129,In_757);
xnor U804 (N_804,N_342,N_657);
xnor U805 (N_805,In_50,N_550);
xor U806 (N_806,N_758,In_1034);
or U807 (N_807,In_321,In_373);
nand U808 (N_808,N_215,In_1458);
xnor U809 (N_809,N_171,In_1193);
or U810 (N_810,N_660,N_503);
or U811 (N_811,In_353,N_175);
nand U812 (N_812,N_428,In_1463);
nand U813 (N_813,N_731,In_875);
or U814 (N_814,In_31,N_541);
xnor U815 (N_815,N_590,N_760);
nor U816 (N_816,N_154,In_1275);
and U817 (N_817,In_529,In_346);
and U818 (N_818,N_704,N_439);
nand U819 (N_819,N_419,N_725);
xnor U820 (N_820,In_63,N_788);
nand U821 (N_821,N_711,N_509);
nor U822 (N_822,N_719,N_620);
or U823 (N_823,In_787,N_689);
xor U824 (N_824,In_454,N_635);
and U825 (N_825,N_702,In_1362);
nand U826 (N_826,In_1059,N_629);
nor U827 (N_827,N_781,In_504);
and U828 (N_828,N_676,In_259);
xor U829 (N_829,N_410,N_234);
or U830 (N_830,In_322,N_755);
or U831 (N_831,In_1346,In_488);
and U832 (N_832,In_825,In_73);
nor U833 (N_833,In_560,In_756);
and U834 (N_834,N_537,N_773);
and U835 (N_835,In_882,N_336);
nor U836 (N_836,In_854,N_356);
nand U837 (N_837,N_308,N_688);
nor U838 (N_838,N_33,N_316);
and U839 (N_839,N_790,N_640);
xnor U840 (N_840,In_878,N_331);
xnor U841 (N_841,N_543,N_651);
nand U842 (N_842,N_314,N_618);
or U843 (N_843,N_207,In_539);
nor U844 (N_844,In_601,N_430);
xnor U845 (N_845,In_1308,N_796);
and U846 (N_846,N_558,N_417);
and U847 (N_847,In_887,In_87);
nand U848 (N_848,N_424,N_162);
nand U849 (N_849,N_247,N_147);
and U850 (N_850,In_730,In_105);
xor U851 (N_851,In_339,N_709);
and U852 (N_852,In_834,N_21);
nor U853 (N_853,In_742,In_1152);
or U854 (N_854,In_1268,N_365);
or U855 (N_855,In_985,In_1057);
or U856 (N_856,N_601,N_680);
and U857 (N_857,N_366,In_1001);
xor U858 (N_858,N_437,In_1121);
nand U859 (N_859,N_319,N_525);
or U860 (N_860,In_1262,N_472);
or U861 (N_861,N_452,N_354);
or U862 (N_862,N_167,N_606);
nand U863 (N_863,N_68,N_744);
and U864 (N_864,N_494,N_429);
and U865 (N_865,N_636,N_96);
nor U866 (N_866,N_560,N_686);
xnor U867 (N_867,N_348,N_581);
xnor U868 (N_868,N_721,In_1190);
xnor U869 (N_869,N_756,In_1359);
nand U870 (N_870,N_765,N_748);
nor U871 (N_871,N_536,N_127);
and U872 (N_872,N_623,In_764);
or U873 (N_873,N_768,N_455);
xnor U874 (N_874,N_287,N_458);
nor U875 (N_875,In_1353,N_265);
nand U876 (N_876,N_682,In_1211);
or U877 (N_877,In_1098,N_650);
xnor U878 (N_878,In_546,In_386);
and U879 (N_879,In_1175,In_263);
or U880 (N_880,N_673,N_666);
and U881 (N_881,N_587,N_663);
nand U882 (N_882,N_86,N_397);
xnor U883 (N_883,N_659,N_566);
or U884 (N_884,In_413,N_656);
xnor U885 (N_885,In_15,In_123);
and U886 (N_886,N_120,In_1174);
or U887 (N_887,In_989,N_464);
or U888 (N_888,N_786,In_1311);
or U889 (N_889,N_690,In_1419);
nand U890 (N_890,In_719,N_639);
nor U891 (N_891,N_578,N_462);
xor U892 (N_892,In_236,N_767);
xnor U893 (N_893,In_1160,N_714);
nor U894 (N_894,N_456,N_605);
and U895 (N_895,N_306,N_270);
and U896 (N_896,N_440,N_181);
and U897 (N_897,In_409,N_647);
or U898 (N_898,In_70,N_729);
and U899 (N_899,In_416,In_26);
and U900 (N_900,N_572,N_608);
and U901 (N_901,N_7,In_349);
nor U902 (N_902,N_14,In_501);
xor U903 (N_903,In_976,In_1225);
and U904 (N_904,In_180,N_187);
or U905 (N_905,N_634,N_533);
xnor U906 (N_906,In_1222,N_661);
xor U907 (N_907,N_580,N_447);
and U908 (N_908,In_1019,In_521);
nor U909 (N_909,N_508,In_829);
nor U910 (N_910,In_558,N_681);
xor U911 (N_911,N_399,In_1364);
xor U912 (N_912,N_576,In_387);
xor U913 (N_913,In_519,N_715);
or U914 (N_914,N_357,In_660);
or U915 (N_915,N_98,N_376);
and U916 (N_916,N_664,N_476);
xor U917 (N_917,In_439,N_290);
nand U918 (N_918,N_724,N_261);
xor U919 (N_919,N_648,In_492);
xor U920 (N_920,In_891,N_769);
nand U921 (N_921,In_1449,N_665);
nand U922 (N_922,In_205,N_784);
or U923 (N_923,In_692,N_13);
nor U924 (N_924,N_231,N_344);
nor U925 (N_925,In_611,N_780);
or U926 (N_926,In_1433,In_909);
or U927 (N_927,N_27,N_554);
or U928 (N_928,In_974,N_698);
nand U929 (N_929,N_604,N_478);
xor U930 (N_930,N_746,In_1181);
nand U931 (N_931,N_360,In_615);
xor U932 (N_932,N_610,In_1185);
nor U933 (N_933,In_1011,N_84);
nor U934 (N_934,In_14,N_699);
xnor U935 (N_935,N_557,N_779);
or U936 (N_936,N_785,N_423);
and U937 (N_937,In_411,N_691);
and U938 (N_938,In_484,N_19);
and U939 (N_939,N_612,N_563);
and U940 (N_940,N_726,In_1448);
nand U941 (N_941,N_684,N_283);
or U942 (N_942,N_323,In_1233);
and U943 (N_943,In_1354,In_960);
nor U944 (N_944,N_789,In_468);
or U945 (N_945,N_498,N_754);
nor U946 (N_946,N_514,In_1296);
nor U947 (N_947,N_593,In_110);
xnor U948 (N_948,In_1097,N_36);
nand U949 (N_949,In_0,N_783);
nor U950 (N_950,N_734,N_511);
or U951 (N_951,N_772,N_619);
or U952 (N_952,N_701,N_643);
nand U953 (N_953,N_759,In_1427);
nand U954 (N_954,In_367,In_1260);
nand U955 (N_955,N_607,N_274);
or U956 (N_956,In_475,N_737);
xnor U957 (N_957,In_1487,N_134);
nand U958 (N_958,In_1033,N_282);
and U959 (N_959,N_549,In_1365);
or U960 (N_960,In_911,N_614);
or U961 (N_961,N_670,N_649);
nor U962 (N_962,In_52,N_245);
xnor U963 (N_963,N_551,N_497);
nand U964 (N_964,N_217,In_1322);
nand U965 (N_965,In_1421,In_1411);
and U966 (N_966,N_254,N_778);
xor U967 (N_967,N_491,N_777);
nor U968 (N_968,N_180,N_561);
xnor U969 (N_969,In_179,In_136);
xor U970 (N_970,N_717,In_337);
or U971 (N_971,N_564,In_66);
and U972 (N_972,In_505,N_286);
or U973 (N_973,N_392,N_574);
nand U974 (N_974,N_195,N_644);
or U975 (N_975,In_859,N_532);
or U976 (N_976,In_857,N_708);
and U977 (N_977,N_736,In_1330);
or U978 (N_978,N_312,N_387);
and U979 (N_979,N_530,N_615);
or U980 (N_980,In_904,In_852);
xor U981 (N_981,N_487,N_642);
nand U982 (N_982,N_653,In_318);
nand U983 (N_983,N_280,In_788);
nor U984 (N_984,N_627,In_862);
nand U985 (N_985,N_140,In_915);
nand U986 (N_986,N_685,N_501);
nor U987 (N_987,N_385,N_747);
xnor U988 (N_988,N_337,In_631);
nand U989 (N_989,In_1271,In_1432);
or U990 (N_990,N_315,In_1350);
xnor U991 (N_991,N_621,N_545);
nand U992 (N_992,N_146,N_209);
and U993 (N_993,N_774,In_889);
and U994 (N_994,N_603,N_672);
xnor U995 (N_995,In_217,N_678);
or U996 (N_996,In_279,In_319);
xnor U997 (N_997,In_183,N_370);
and U998 (N_998,In_793,N_579);
nand U999 (N_999,In_490,N_703);
xor U1000 (N_1000,N_878,In_3);
or U1001 (N_1001,N_985,N_671);
and U1002 (N_1002,N_569,N_936);
or U1003 (N_1003,N_823,In_831);
nand U1004 (N_1004,N_885,N_914);
or U1005 (N_1005,N_710,N_827);
and U1006 (N_1006,N_626,N_907);
xnor U1007 (N_1007,N_602,N_761);
and U1008 (N_1008,N_920,N_368);
and U1009 (N_1009,N_952,N_908);
nand U1010 (N_1010,In_1402,N_857);
nand U1011 (N_1011,N_804,N_309);
xor U1012 (N_1012,N_69,N_960);
and U1013 (N_1013,N_882,N_272);
xnor U1014 (N_1014,N_260,In_116);
and U1015 (N_1015,N_963,In_406);
or U1016 (N_1016,N_749,N_951);
nor U1017 (N_1017,N_870,N_2);
or U1018 (N_1018,N_893,N_628);
nor U1019 (N_1019,In_897,N_631);
nor U1020 (N_1020,N_888,In_774);
xor U1021 (N_1021,N_900,In_633);
nand U1022 (N_1022,N_828,N_432);
nor U1023 (N_1023,In_1424,N_485);
or U1024 (N_1024,In_343,N_512);
nand U1025 (N_1025,N_125,N_630);
and U1026 (N_1026,N_901,N_921);
or U1027 (N_1027,In_88,N_990);
xor U1028 (N_1028,In_1494,In_430);
xnor U1029 (N_1029,N_854,In_1230);
xnor U1030 (N_1030,N_552,N_807);
or U1031 (N_1031,N_838,N_876);
and U1032 (N_1032,N_683,N_845);
nand U1033 (N_1033,In_1418,N_646);
or U1034 (N_1034,N_757,In_1101);
nand U1035 (N_1035,N_461,In_575);
or U1036 (N_1036,N_962,In_152);
and U1037 (N_1037,N_968,N_733);
or U1038 (N_1038,N_808,N_816);
or U1039 (N_1039,N_202,N_800);
nor U1040 (N_1040,In_185,In_760);
xnor U1041 (N_1041,N_841,N_794);
xnor U1042 (N_1042,In_1429,In_1393);
or U1043 (N_1043,N_222,N_740);
nand U1044 (N_1044,N_873,N_822);
nand U1045 (N_1045,In_630,N_609);
or U1046 (N_1046,N_813,N_441);
nor U1047 (N_1047,N_695,N_847);
or U1048 (N_1048,N_846,N_299);
or U1049 (N_1049,N_17,In_1263);
nand U1050 (N_1050,In_1080,N_625);
and U1051 (N_1051,N_879,N_811);
nand U1052 (N_1052,N_815,N_730);
or U1053 (N_1053,N_909,N_961);
xnor U1054 (N_1054,In_847,N_843);
nand U1055 (N_1055,N_63,N_812);
xnor U1056 (N_1056,N_421,N_450);
nand U1057 (N_1057,N_851,N_654);
nand U1058 (N_1058,In_564,N_588);
xor U1059 (N_1059,N_874,N_697);
and U1060 (N_1060,N_809,N_735);
and U1061 (N_1061,N_896,N_938);
nand U1062 (N_1062,N_996,In_98);
nand U1063 (N_1063,N_713,N_924);
nand U1064 (N_1064,N_867,N_949);
and U1065 (N_1065,N_465,N_934);
nand U1066 (N_1066,N_953,In_93);
xor U1067 (N_1067,N_707,N_821);
nor U1068 (N_1068,In_919,In_670);
xor U1069 (N_1069,N_633,N_49);
xor U1070 (N_1070,N_128,N_799);
nor U1071 (N_1071,N_913,N_944);
or U1072 (N_1072,In_1032,N_352);
nand U1073 (N_1073,N_844,N_972);
xnor U1074 (N_1074,N_438,In_1066);
or U1075 (N_1075,N_967,N_743);
and U1076 (N_1076,N_143,N_687);
nand U1077 (N_1077,N_632,N_928);
and U1078 (N_1078,In_350,N_852);
or U1079 (N_1079,N_959,N_712);
nand U1080 (N_1080,N_916,N_925);
and U1081 (N_1081,In_1002,N_313);
or U1082 (N_1082,N_892,In_235);
nor U1083 (N_1083,N_466,N_999);
or U1084 (N_1084,N_919,In_569);
and U1085 (N_1085,N_834,N_766);
and U1086 (N_1086,In_1480,In_1422);
xnor U1087 (N_1087,N_947,N_958);
or U1088 (N_1088,N_964,N_880);
or U1089 (N_1089,N_992,N_956);
nand U1090 (N_1090,N_818,N_869);
and U1091 (N_1091,N_82,N_638);
and U1092 (N_1092,N_745,N_825);
xnor U1093 (N_1093,N_191,N_591);
nand U1094 (N_1094,In_1281,N_830);
and U1095 (N_1095,In_1498,In_220);
and U1096 (N_1096,N_863,N_832);
nand U1097 (N_1097,In_1460,N_624);
xor U1098 (N_1098,In_864,N_700);
nand U1099 (N_1099,N_877,In_511);
and U1100 (N_1100,N_770,In_303);
or U1101 (N_1101,N_911,N_973);
and U1102 (N_1102,N_718,In_1087);
xnor U1103 (N_1103,N_720,N_347);
or U1104 (N_1104,N_997,N_970);
and U1105 (N_1105,N_480,In_114);
nor U1106 (N_1106,N_408,N_829);
nand U1107 (N_1107,N_883,N_984);
nand U1108 (N_1108,In_1021,N_775);
and U1109 (N_1109,N_810,N_325);
and U1110 (N_1110,N_897,N_390);
and U1111 (N_1111,N_538,N_903);
and U1112 (N_1112,N_969,N_932);
and U1113 (N_1113,In_141,N_998);
and U1114 (N_1114,N_407,N_929);
and U1115 (N_1115,N_652,N_871);
and U1116 (N_1116,N_803,N_941);
or U1117 (N_1117,N_669,N_872);
and U1118 (N_1118,In_94,N_986);
and U1119 (N_1119,N_837,N_965);
or U1120 (N_1120,In_301,N_886);
and U1121 (N_1121,N_795,N_995);
nand U1122 (N_1122,N_266,N_884);
or U1123 (N_1123,In_1437,N_943);
and U1124 (N_1124,In_432,In_1030);
and U1125 (N_1125,In_1061,N_875);
nand U1126 (N_1126,N_946,In_134);
nand U1127 (N_1127,N_753,N_727);
xor U1128 (N_1128,N_860,N_927);
or U1129 (N_1129,N_599,N_842);
nor U1130 (N_1130,N_817,N_894);
xor U1131 (N_1131,In_837,N_470);
xnor U1132 (N_1132,N_716,In_48);
xnor U1133 (N_1133,N_741,In_1132);
or U1134 (N_1134,In_525,N_637);
xor U1135 (N_1135,N_915,N_887);
nor U1136 (N_1136,N_723,In_213);
or U1137 (N_1137,N_820,N_420);
and U1138 (N_1138,N_300,N_782);
nor U1139 (N_1139,N_819,N_542);
xor U1140 (N_1140,N_912,N_994);
xor U1141 (N_1141,N_594,In_1400);
nand U1142 (N_1142,In_642,N_474);
or U1143 (N_1143,N_531,N_655);
or U1144 (N_1144,N_930,N_677);
or U1145 (N_1145,N_434,N_592);
or U1146 (N_1146,N_722,In_174);
or U1147 (N_1147,In_1265,N_174);
and U1148 (N_1148,N_750,In_250);
nor U1149 (N_1149,N_974,N_732);
nand U1150 (N_1150,In_562,N_983);
and U1151 (N_1151,N_917,N_371);
nand U1152 (N_1152,N_645,N_482);
nand U1153 (N_1153,N_801,N_738);
and U1154 (N_1154,In_933,N_826);
xor U1155 (N_1155,In_395,N_728);
nor U1156 (N_1156,In_1046,N_151);
and U1157 (N_1157,N_792,N_674);
xor U1158 (N_1158,N_568,N_948);
nand U1159 (N_1159,N_179,N_805);
xor U1160 (N_1160,N_931,N_989);
and U1161 (N_1161,N_763,N_600);
or U1162 (N_1162,N_942,N_445);
nor U1163 (N_1163,In_1305,N_868);
xnor U1164 (N_1164,In_773,N_622);
nor U1165 (N_1165,N_616,N_431);
xnor U1166 (N_1166,N_667,N_764);
and U1167 (N_1167,N_422,N_31);
nor U1168 (N_1168,N_881,N_945);
nand U1169 (N_1169,N_987,N_864);
and U1170 (N_1170,N_891,N_939);
xnor U1171 (N_1171,N_979,N_507);
or U1172 (N_1172,N_762,In_104);
nor U1173 (N_1173,N_988,In_535);
and U1174 (N_1174,N_305,N_977);
or U1175 (N_1175,N_980,N_814);
nand U1176 (N_1176,N_141,In_1388);
nand U1177 (N_1177,In_1195,In_548);
nor U1178 (N_1178,N_662,In_1170);
xnor U1179 (N_1179,N_890,N_978);
or U1180 (N_1180,N_861,N_856);
nand U1181 (N_1181,N_176,N_546);
xnor U1182 (N_1182,N_853,In_604);
xnor U1183 (N_1183,In_751,N_955);
nand U1184 (N_1184,N_442,N_923);
xor U1185 (N_1185,In_612,N_694);
nor U1186 (N_1186,N_898,In_880);
or U1187 (N_1187,N_567,N_321);
xor U1188 (N_1188,N_976,N_239);
nor U1189 (N_1189,N_865,N_918);
nand U1190 (N_1190,N_910,In_80);
nand U1191 (N_1191,In_108,N_922);
or U1192 (N_1192,In_22,N_679);
nor U1193 (N_1193,N_971,N_380);
and U1194 (N_1194,N_848,N_326);
or U1195 (N_1195,N_840,N_906);
nor U1196 (N_1196,N_833,N_902);
nor U1197 (N_1197,In_999,N_351);
or U1198 (N_1198,N_802,N_798);
nand U1199 (N_1199,N_194,N_991);
nand U1200 (N_1200,N_1065,N_1017);
and U1201 (N_1201,N_153,N_1133);
nor U1202 (N_1202,N_1118,N_1126);
nor U1203 (N_1203,N_862,N_454);
nor U1204 (N_1204,N_1185,N_1087);
xor U1205 (N_1205,N_1004,N_1063);
nor U1206 (N_1206,N_1135,N_1192);
or U1207 (N_1207,N_1136,N_1188);
nor U1208 (N_1208,N_1112,N_835);
and U1209 (N_1209,N_1037,N_1138);
and U1210 (N_1210,N_1158,In_953);
and U1211 (N_1211,N_895,N_1179);
xor U1212 (N_1212,N_797,N_1038);
or U1213 (N_1213,N_993,N_1080);
or U1214 (N_1214,N_1100,N_866);
xor U1215 (N_1215,N_150,N_1102);
and U1216 (N_1216,N_693,N_1069);
or U1217 (N_1217,N_1098,N_486);
or U1218 (N_1218,N_831,N_1071);
and U1219 (N_1219,N_1083,In_537);
or U1220 (N_1220,N_1095,N_1161);
and U1221 (N_1221,N_1084,N_791);
nor U1222 (N_1222,N_1131,N_1175);
xor U1223 (N_1223,N_613,N_1043);
xor U1224 (N_1224,N_1048,N_463);
nand U1225 (N_1225,N_1127,In_487);
nand U1226 (N_1226,N_1040,N_1107);
nand U1227 (N_1227,N_859,N_1111);
or U1228 (N_1228,N_1020,N_1047);
or U1229 (N_1229,N_1093,N_1097);
nor U1230 (N_1230,N_1142,N_1176);
nor U1231 (N_1231,N_1180,N_1064);
or U1232 (N_1232,N_1125,In_20);
and U1233 (N_1233,N_1195,In_1282);
and U1234 (N_1234,N_1077,N_1061);
or U1235 (N_1235,N_824,N_595);
or U1236 (N_1236,N_904,N_1166);
nand U1237 (N_1237,N_1010,N_1003);
nand U1238 (N_1238,N_1181,N_1058);
and U1239 (N_1239,N_742,In_276);
xor U1240 (N_1240,N_1025,In_320);
nand U1241 (N_1241,N_692,N_418);
and U1242 (N_1242,In_957,N_1150);
xor U1243 (N_1243,N_1117,N_34);
and U1244 (N_1244,N_488,N_1105);
and U1245 (N_1245,N_771,N_1006);
nand U1246 (N_1246,N_1089,N_493);
or U1247 (N_1247,N_1066,N_1120);
nand U1248 (N_1248,N_1073,N_1169);
or U1249 (N_1249,N_1113,N_1018);
xor U1250 (N_1250,In_1428,N_1092);
or U1251 (N_1251,N_1021,N_1094);
or U1252 (N_1252,N_1193,N_1050);
xor U1253 (N_1253,N_696,N_899);
and U1254 (N_1254,N_1143,N_1075);
or U1255 (N_1255,N_1148,N_1076);
xor U1256 (N_1256,N_1088,N_1140);
and U1257 (N_1257,N_1044,In_808);
xnor U1258 (N_1258,In_399,N_1191);
nor U1259 (N_1259,N_1168,N_617);
xnor U1260 (N_1260,N_611,N_1055);
or U1261 (N_1261,N_1051,N_359);
or U1262 (N_1262,N_926,N_905);
or U1263 (N_1263,N_1114,N_1005);
nand U1264 (N_1264,N_705,N_1034);
or U1265 (N_1265,N_539,N_675);
xnor U1266 (N_1266,In_1173,N_1163);
and U1267 (N_1267,N_855,N_1057);
or U1268 (N_1268,N_1041,N_954);
or U1269 (N_1269,In_282,N_1015);
nor U1270 (N_1270,N_1178,N_451);
nand U1271 (N_1271,N_1035,N_1000);
and U1272 (N_1272,N_1108,N_1183);
or U1273 (N_1273,N_1170,N_1164);
nor U1274 (N_1274,N_1198,In_267);
xor U1275 (N_1275,N_1130,N_975);
nand U1276 (N_1276,In_150,N_1062);
nand U1277 (N_1277,N_276,N_1123);
xor U1278 (N_1278,N_1144,N_950);
or U1279 (N_1279,In_210,N_1106);
and U1280 (N_1280,N_940,In_458);
or U1281 (N_1281,N_1039,N_933);
xnor U1282 (N_1282,N_1026,N_1174);
nand U1283 (N_1283,N_836,N_1159);
nand U1284 (N_1284,N_739,N_1008);
nor U1285 (N_1285,N_1036,N_981);
xnor U1286 (N_1286,N_937,N_1019);
or U1287 (N_1287,N_1001,N_1110);
nor U1288 (N_1288,N_1134,N_1099);
xor U1289 (N_1289,N_468,N_1129);
and U1290 (N_1290,N_1009,N_1104);
or U1291 (N_1291,N_1033,N_1060);
nor U1292 (N_1292,N_1156,N_1141);
nand U1293 (N_1293,N_1160,N_1184);
xnor U1294 (N_1294,N_1028,N_1096);
or U1295 (N_1295,N_1189,N_1042);
nor U1296 (N_1296,N_1059,N_1086);
nor U1297 (N_1297,N_1085,N_457);
xor U1298 (N_1298,N_535,N_1024);
and U1299 (N_1299,N_1146,N_105);
xnor U1300 (N_1300,N_776,In_1378);
nor U1301 (N_1301,N_787,N_1022);
nor U1302 (N_1302,N_1171,N_1072);
and U1303 (N_1303,N_1103,N_1013);
xor U1304 (N_1304,N_1002,N_469);
xnor U1305 (N_1305,N_1145,N_1091);
or U1306 (N_1306,N_982,N_1116);
and U1307 (N_1307,N_850,N_1011);
and U1308 (N_1308,N_889,N_1070);
xor U1309 (N_1309,N_839,N_806);
nand U1310 (N_1310,N_1032,N_1172);
nor U1311 (N_1311,N_849,N_553);
and U1312 (N_1312,N_1082,N_1078);
or U1313 (N_1313,N_1197,N_1154);
nor U1314 (N_1314,N_1153,N_1122);
nor U1315 (N_1315,In_849,N_393);
nand U1316 (N_1316,N_1173,N_1139);
and U1317 (N_1317,N_1101,In_804);
nand U1318 (N_1318,N_641,N_1016);
and U1319 (N_1319,N_658,N_1079);
nand U1320 (N_1320,N_1031,N_1029);
and U1321 (N_1321,N_1132,N_1196);
or U1322 (N_1322,N_1049,N_1187);
xor U1323 (N_1323,N_1151,N_232);
or U1324 (N_1324,N_1124,N_1053);
or U1325 (N_1325,N_203,N_1137);
xnor U1326 (N_1326,N_1147,N_255);
nor U1327 (N_1327,N_236,In_819);
nor U1328 (N_1328,N_1012,N_966);
and U1329 (N_1329,N_1119,N_1074);
nand U1330 (N_1330,N_751,N_1162);
xnor U1331 (N_1331,N_1014,N_1199);
nor U1332 (N_1332,N_858,N_1056);
xnor U1333 (N_1333,N_1177,N_1023);
or U1334 (N_1334,N_1052,N_1030);
or U1335 (N_1335,N_1068,N_1194);
xnor U1336 (N_1336,N_1155,N_1046);
nand U1337 (N_1337,N_1045,N_1167);
nand U1338 (N_1338,N_935,N_544);
nor U1339 (N_1339,N_957,N_1081);
xnor U1340 (N_1340,N_1067,N_1109);
xor U1341 (N_1341,N_1182,N_1115);
xnor U1342 (N_1342,N_1190,N_1121);
or U1343 (N_1343,N_1152,N_1157);
nor U1344 (N_1344,N_752,N_1054);
and U1345 (N_1345,N_1149,N_793);
or U1346 (N_1346,N_1165,N_1128);
and U1347 (N_1347,N_1007,N_523);
or U1348 (N_1348,N_706,N_1186);
nand U1349 (N_1349,N_1090,N_1027);
and U1350 (N_1350,N_1113,N_1179);
nand U1351 (N_1351,In_282,N_1075);
xnor U1352 (N_1352,N_1124,N_824);
xor U1353 (N_1353,N_1135,N_1098);
xor U1354 (N_1354,N_1007,N_1180);
xnor U1355 (N_1355,N_1030,N_1000);
nand U1356 (N_1356,N_1094,N_693);
xnor U1357 (N_1357,N_1191,N_1001);
and U1358 (N_1358,N_866,In_1378);
xor U1359 (N_1359,N_1127,N_1019);
nand U1360 (N_1360,In_282,N_797);
and U1361 (N_1361,N_859,N_1002);
nor U1362 (N_1362,N_1022,In_1378);
and U1363 (N_1363,N_1078,N_1107);
and U1364 (N_1364,N_1030,N_739);
and U1365 (N_1365,N_1037,N_1133);
xnor U1366 (N_1366,N_1088,N_937);
xor U1367 (N_1367,N_675,N_1063);
xnor U1368 (N_1368,N_1097,N_1000);
nor U1369 (N_1369,N_1076,N_935);
nor U1370 (N_1370,N_1135,N_1125);
nand U1371 (N_1371,N_752,In_1378);
xor U1372 (N_1372,N_1152,N_150);
and U1373 (N_1373,N_1192,N_153);
and U1374 (N_1374,N_771,N_1070);
nor U1375 (N_1375,N_1091,N_1122);
nand U1376 (N_1376,N_1003,N_1033);
or U1377 (N_1377,N_1054,N_1106);
nor U1378 (N_1378,N_1133,N_1095);
and U1379 (N_1379,N_1048,N_862);
nand U1380 (N_1380,N_1166,N_1151);
or U1381 (N_1381,N_1177,N_1076);
nor U1382 (N_1382,N_1056,N_1067);
nor U1383 (N_1383,N_1065,N_595);
or U1384 (N_1384,N_1089,N_1024);
xnor U1385 (N_1385,N_1183,N_1008);
xor U1386 (N_1386,N_1088,N_1127);
and U1387 (N_1387,N_1199,N_1137);
nand U1388 (N_1388,N_1143,N_1172);
nand U1389 (N_1389,N_658,N_1154);
and U1390 (N_1390,N_706,N_1126);
and U1391 (N_1391,N_523,N_981);
nor U1392 (N_1392,N_469,N_544);
nor U1393 (N_1393,N_493,N_1176);
or U1394 (N_1394,N_950,N_1119);
and U1395 (N_1395,N_1022,N_1088);
xor U1396 (N_1396,N_1049,N_1164);
nor U1397 (N_1397,N_1049,N_544);
and U1398 (N_1398,N_1069,N_1029);
and U1399 (N_1399,N_975,N_899);
and U1400 (N_1400,N_1351,N_1303);
and U1401 (N_1401,N_1239,N_1343);
nor U1402 (N_1402,N_1367,N_1387);
and U1403 (N_1403,N_1368,N_1372);
xnor U1404 (N_1404,N_1383,N_1398);
and U1405 (N_1405,N_1201,N_1318);
xnor U1406 (N_1406,N_1245,N_1207);
and U1407 (N_1407,N_1344,N_1250);
and U1408 (N_1408,N_1355,N_1249);
xor U1409 (N_1409,N_1257,N_1311);
nand U1410 (N_1410,N_1271,N_1347);
nor U1411 (N_1411,N_1206,N_1366);
xnor U1412 (N_1412,N_1334,N_1302);
nor U1413 (N_1413,N_1342,N_1229);
or U1414 (N_1414,N_1220,N_1396);
nand U1415 (N_1415,N_1376,N_1270);
xnor U1416 (N_1416,N_1277,N_1203);
xnor U1417 (N_1417,N_1269,N_1228);
nand U1418 (N_1418,N_1314,N_1328);
nand U1419 (N_1419,N_1247,N_1246);
and U1420 (N_1420,N_1236,N_1352);
xor U1421 (N_1421,N_1231,N_1253);
and U1422 (N_1422,N_1258,N_1243);
nand U1423 (N_1423,N_1373,N_1320);
xnor U1424 (N_1424,N_1293,N_1386);
nand U1425 (N_1425,N_1210,N_1323);
and U1426 (N_1426,N_1362,N_1345);
xor U1427 (N_1427,N_1268,N_1370);
nor U1428 (N_1428,N_1297,N_1260);
nor U1429 (N_1429,N_1313,N_1224);
nand U1430 (N_1430,N_1321,N_1391);
xnor U1431 (N_1431,N_1256,N_1209);
and U1432 (N_1432,N_1353,N_1255);
xor U1433 (N_1433,N_1213,N_1218);
nand U1434 (N_1434,N_1287,N_1369);
nand U1435 (N_1435,N_1278,N_1230);
and U1436 (N_1436,N_1300,N_1291);
nor U1437 (N_1437,N_1374,N_1350);
nand U1438 (N_1438,N_1216,N_1379);
nand U1439 (N_1439,N_1381,N_1215);
nand U1440 (N_1440,N_1290,N_1358);
nand U1441 (N_1441,N_1332,N_1251);
xor U1442 (N_1442,N_1208,N_1326);
nand U1443 (N_1443,N_1262,N_1275);
or U1444 (N_1444,N_1272,N_1346);
or U1445 (N_1445,N_1283,N_1382);
nand U1446 (N_1446,N_1338,N_1325);
xnor U1447 (N_1447,N_1299,N_1312);
nand U1448 (N_1448,N_1307,N_1248);
nor U1449 (N_1449,N_1306,N_1254);
xor U1450 (N_1450,N_1324,N_1341);
and U1451 (N_1451,N_1298,N_1214);
or U1452 (N_1452,N_1288,N_1319);
nor U1453 (N_1453,N_1392,N_1223);
xnor U1454 (N_1454,N_1237,N_1294);
xor U1455 (N_1455,N_1265,N_1394);
and U1456 (N_1456,N_1317,N_1333);
nor U1457 (N_1457,N_1361,N_1322);
nand U1458 (N_1458,N_1327,N_1227);
or U1459 (N_1459,N_1356,N_1371);
and U1460 (N_1460,N_1360,N_1395);
and U1461 (N_1461,N_1388,N_1292);
xor U1462 (N_1462,N_1259,N_1305);
nand U1463 (N_1463,N_1393,N_1232);
nand U1464 (N_1464,N_1284,N_1289);
nand U1465 (N_1465,N_1357,N_1222);
and U1466 (N_1466,N_1263,N_1349);
nor U1467 (N_1467,N_1205,N_1380);
nand U1468 (N_1468,N_1244,N_1264);
and U1469 (N_1469,N_1281,N_1336);
and U1470 (N_1470,N_1384,N_1363);
nand U1471 (N_1471,N_1339,N_1241);
xnor U1472 (N_1472,N_1340,N_1375);
or U1473 (N_1473,N_1279,N_1252);
nand U1474 (N_1474,N_1308,N_1359);
and U1475 (N_1475,N_1309,N_1389);
or U1476 (N_1476,N_1286,N_1304);
and U1477 (N_1477,N_1365,N_1219);
nand U1478 (N_1478,N_1282,N_1240);
nand U1479 (N_1479,N_1285,N_1266);
or U1480 (N_1480,N_1238,N_1295);
nand U1481 (N_1481,N_1390,N_1364);
and U1482 (N_1482,N_1225,N_1377);
nand U1483 (N_1483,N_1221,N_1397);
nor U1484 (N_1484,N_1399,N_1315);
or U1485 (N_1485,N_1211,N_1316);
nor U1486 (N_1486,N_1378,N_1310);
nor U1487 (N_1487,N_1330,N_1280);
nand U1488 (N_1488,N_1274,N_1202);
nor U1489 (N_1489,N_1261,N_1212);
and U1490 (N_1490,N_1296,N_1331);
nor U1491 (N_1491,N_1348,N_1200);
and U1492 (N_1492,N_1385,N_1354);
xor U1493 (N_1493,N_1337,N_1329);
nor U1494 (N_1494,N_1226,N_1267);
nand U1495 (N_1495,N_1235,N_1276);
and U1496 (N_1496,N_1335,N_1301);
and U1497 (N_1497,N_1234,N_1242);
and U1498 (N_1498,N_1204,N_1217);
nand U1499 (N_1499,N_1233,N_1273);
or U1500 (N_1500,N_1239,N_1205);
nor U1501 (N_1501,N_1311,N_1203);
and U1502 (N_1502,N_1378,N_1226);
and U1503 (N_1503,N_1251,N_1290);
xnor U1504 (N_1504,N_1349,N_1294);
nand U1505 (N_1505,N_1214,N_1387);
and U1506 (N_1506,N_1201,N_1243);
xor U1507 (N_1507,N_1294,N_1265);
xnor U1508 (N_1508,N_1369,N_1321);
or U1509 (N_1509,N_1258,N_1398);
nand U1510 (N_1510,N_1311,N_1224);
xnor U1511 (N_1511,N_1342,N_1301);
and U1512 (N_1512,N_1366,N_1302);
nand U1513 (N_1513,N_1359,N_1224);
nor U1514 (N_1514,N_1222,N_1233);
xnor U1515 (N_1515,N_1359,N_1273);
nor U1516 (N_1516,N_1216,N_1334);
nor U1517 (N_1517,N_1205,N_1393);
xnor U1518 (N_1518,N_1218,N_1269);
nor U1519 (N_1519,N_1338,N_1323);
and U1520 (N_1520,N_1343,N_1270);
and U1521 (N_1521,N_1319,N_1308);
xor U1522 (N_1522,N_1255,N_1335);
and U1523 (N_1523,N_1391,N_1282);
nor U1524 (N_1524,N_1241,N_1283);
nand U1525 (N_1525,N_1358,N_1355);
xnor U1526 (N_1526,N_1215,N_1324);
and U1527 (N_1527,N_1202,N_1209);
and U1528 (N_1528,N_1212,N_1323);
nand U1529 (N_1529,N_1319,N_1350);
or U1530 (N_1530,N_1201,N_1251);
nand U1531 (N_1531,N_1323,N_1301);
and U1532 (N_1532,N_1395,N_1216);
nand U1533 (N_1533,N_1347,N_1261);
and U1534 (N_1534,N_1271,N_1329);
nand U1535 (N_1535,N_1342,N_1387);
xnor U1536 (N_1536,N_1330,N_1344);
nor U1537 (N_1537,N_1293,N_1207);
nor U1538 (N_1538,N_1280,N_1301);
xor U1539 (N_1539,N_1248,N_1344);
or U1540 (N_1540,N_1308,N_1399);
and U1541 (N_1541,N_1387,N_1329);
xnor U1542 (N_1542,N_1355,N_1335);
nand U1543 (N_1543,N_1333,N_1237);
and U1544 (N_1544,N_1306,N_1310);
and U1545 (N_1545,N_1326,N_1376);
xnor U1546 (N_1546,N_1357,N_1275);
or U1547 (N_1547,N_1302,N_1382);
nand U1548 (N_1548,N_1220,N_1354);
and U1549 (N_1549,N_1221,N_1218);
nor U1550 (N_1550,N_1266,N_1240);
nor U1551 (N_1551,N_1372,N_1233);
nand U1552 (N_1552,N_1224,N_1290);
nor U1553 (N_1553,N_1375,N_1266);
nor U1554 (N_1554,N_1287,N_1368);
xnor U1555 (N_1555,N_1344,N_1332);
nand U1556 (N_1556,N_1324,N_1374);
nor U1557 (N_1557,N_1210,N_1373);
xor U1558 (N_1558,N_1286,N_1250);
xor U1559 (N_1559,N_1313,N_1356);
nand U1560 (N_1560,N_1350,N_1217);
or U1561 (N_1561,N_1220,N_1269);
nor U1562 (N_1562,N_1331,N_1294);
or U1563 (N_1563,N_1247,N_1308);
nand U1564 (N_1564,N_1244,N_1361);
xor U1565 (N_1565,N_1206,N_1242);
nand U1566 (N_1566,N_1241,N_1226);
nand U1567 (N_1567,N_1207,N_1371);
xnor U1568 (N_1568,N_1257,N_1378);
and U1569 (N_1569,N_1215,N_1335);
nor U1570 (N_1570,N_1261,N_1283);
or U1571 (N_1571,N_1310,N_1329);
nor U1572 (N_1572,N_1334,N_1368);
or U1573 (N_1573,N_1266,N_1380);
xor U1574 (N_1574,N_1262,N_1240);
nand U1575 (N_1575,N_1288,N_1360);
nand U1576 (N_1576,N_1390,N_1237);
nand U1577 (N_1577,N_1240,N_1292);
and U1578 (N_1578,N_1235,N_1308);
nand U1579 (N_1579,N_1254,N_1277);
nand U1580 (N_1580,N_1240,N_1255);
or U1581 (N_1581,N_1233,N_1235);
xnor U1582 (N_1582,N_1278,N_1295);
and U1583 (N_1583,N_1371,N_1257);
nand U1584 (N_1584,N_1235,N_1346);
xnor U1585 (N_1585,N_1391,N_1296);
and U1586 (N_1586,N_1211,N_1317);
or U1587 (N_1587,N_1346,N_1260);
nand U1588 (N_1588,N_1354,N_1377);
nor U1589 (N_1589,N_1395,N_1290);
xnor U1590 (N_1590,N_1364,N_1249);
xnor U1591 (N_1591,N_1371,N_1296);
xnor U1592 (N_1592,N_1358,N_1292);
xnor U1593 (N_1593,N_1200,N_1282);
or U1594 (N_1594,N_1368,N_1211);
and U1595 (N_1595,N_1242,N_1336);
and U1596 (N_1596,N_1337,N_1292);
or U1597 (N_1597,N_1394,N_1275);
and U1598 (N_1598,N_1253,N_1218);
and U1599 (N_1599,N_1313,N_1331);
or U1600 (N_1600,N_1413,N_1596);
or U1601 (N_1601,N_1573,N_1575);
and U1602 (N_1602,N_1507,N_1496);
and U1603 (N_1603,N_1581,N_1543);
nor U1604 (N_1604,N_1571,N_1560);
nand U1605 (N_1605,N_1487,N_1480);
or U1606 (N_1606,N_1474,N_1556);
or U1607 (N_1607,N_1422,N_1586);
nand U1608 (N_1608,N_1448,N_1438);
or U1609 (N_1609,N_1419,N_1404);
and U1610 (N_1610,N_1436,N_1595);
or U1611 (N_1611,N_1473,N_1454);
and U1612 (N_1612,N_1402,N_1488);
or U1613 (N_1613,N_1457,N_1555);
nor U1614 (N_1614,N_1443,N_1501);
nor U1615 (N_1615,N_1461,N_1572);
nor U1616 (N_1616,N_1414,N_1500);
or U1617 (N_1617,N_1551,N_1462);
nor U1618 (N_1618,N_1511,N_1469);
nor U1619 (N_1619,N_1431,N_1442);
and U1620 (N_1620,N_1456,N_1441);
and U1621 (N_1621,N_1528,N_1499);
nor U1622 (N_1622,N_1524,N_1517);
xnor U1623 (N_1623,N_1439,N_1411);
nand U1624 (N_1624,N_1460,N_1588);
and U1625 (N_1625,N_1493,N_1545);
nor U1626 (N_1626,N_1550,N_1599);
nor U1627 (N_1627,N_1526,N_1435);
nand U1628 (N_1628,N_1428,N_1475);
xor U1629 (N_1629,N_1522,N_1564);
xnor U1630 (N_1630,N_1514,N_1536);
nor U1631 (N_1631,N_1486,N_1531);
or U1632 (N_1632,N_1539,N_1446);
and U1633 (N_1633,N_1598,N_1447);
nand U1634 (N_1634,N_1585,N_1544);
nand U1635 (N_1635,N_1540,N_1410);
and U1636 (N_1636,N_1466,N_1542);
nand U1637 (N_1637,N_1532,N_1527);
and U1638 (N_1638,N_1465,N_1403);
or U1639 (N_1639,N_1587,N_1491);
nand U1640 (N_1640,N_1459,N_1429);
and U1641 (N_1641,N_1518,N_1502);
or U1642 (N_1642,N_1440,N_1521);
xor U1643 (N_1643,N_1558,N_1415);
and U1644 (N_1644,N_1552,N_1437);
and U1645 (N_1645,N_1497,N_1568);
xor U1646 (N_1646,N_1567,N_1516);
nor U1647 (N_1647,N_1453,N_1452);
nor U1648 (N_1648,N_1510,N_1530);
xnor U1649 (N_1649,N_1503,N_1546);
nor U1650 (N_1650,N_1405,N_1471);
nand U1651 (N_1651,N_1504,N_1467);
and U1652 (N_1652,N_1538,N_1498);
or U1653 (N_1653,N_1529,N_1570);
nor U1654 (N_1654,N_1478,N_1458);
xor U1655 (N_1655,N_1432,N_1424);
or U1656 (N_1656,N_1508,N_1485);
nand U1657 (N_1657,N_1434,N_1463);
xor U1658 (N_1658,N_1548,N_1512);
or U1659 (N_1659,N_1583,N_1579);
xnor U1660 (N_1660,N_1576,N_1561);
xnor U1661 (N_1661,N_1477,N_1569);
xnor U1662 (N_1662,N_1574,N_1563);
nor U1663 (N_1663,N_1554,N_1597);
and U1664 (N_1664,N_1408,N_1580);
and U1665 (N_1665,N_1594,N_1451);
nand U1666 (N_1666,N_1534,N_1505);
or U1667 (N_1667,N_1406,N_1407);
xnor U1668 (N_1668,N_1523,N_1557);
nand U1669 (N_1669,N_1430,N_1520);
and U1670 (N_1670,N_1578,N_1455);
or U1671 (N_1671,N_1515,N_1450);
or U1672 (N_1672,N_1417,N_1418);
and U1673 (N_1673,N_1470,N_1547);
or U1674 (N_1674,N_1412,N_1553);
or U1675 (N_1675,N_1590,N_1489);
nor U1676 (N_1676,N_1400,N_1562);
nand U1677 (N_1677,N_1484,N_1535);
nand U1678 (N_1678,N_1409,N_1577);
xor U1679 (N_1679,N_1589,N_1537);
and U1680 (N_1680,N_1565,N_1479);
nor U1681 (N_1681,N_1416,N_1427);
and U1682 (N_1682,N_1519,N_1433);
nand U1683 (N_1683,N_1513,N_1566);
and U1684 (N_1684,N_1506,N_1449);
xnor U1685 (N_1685,N_1445,N_1509);
xor U1686 (N_1686,N_1533,N_1494);
nand U1687 (N_1687,N_1423,N_1426);
nor U1688 (N_1688,N_1401,N_1541);
nand U1689 (N_1689,N_1592,N_1425);
nor U1690 (N_1690,N_1584,N_1420);
nand U1691 (N_1691,N_1468,N_1490);
or U1692 (N_1692,N_1472,N_1549);
nand U1693 (N_1693,N_1476,N_1482);
xnor U1694 (N_1694,N_1495,N_1481);
nand U1695 (N_1695,N_1492,N_1593);
xor U1696 (N_1696,N_1591,N_1582);
xor U1697 (N_1697,N_1464,N_1559);
and U1698 (N_1698,N_1444,N_1525);
nand U1699 (N_1699,N_1421,N_1483);
nand U1700 (N_1700,N_1565,N_1499);
or U1701 (N_1701,N_1407,N_1466);
nor U1702 (N_1702,N_1590,N_1503);
nand U1703 (N_1703,N_1527,N_1564);
nand U1704 (N_1704,N_1514,N_1479);
or U1705 (N_1705,N_1404,N_1407);
nand U1706 (N_1706,N_1542,N_1490);
xnor U1707 (N_1707,N_1500,N_1456);
nand U1708 (N_1708,N_1565,N_1502);
xor U1709 (N_1709,N_1522,N_1484);
or U1710 (N_1710,N_1578,N_1540);
and U1711 (N_1711,N_1544,N_1524);
nor U1712 (N_1712,N_1550,N_1426);
and U1713 (N_1713,N_1574,N_1454);
nor U1714 (N_1714,N_1588,N_1430);
and U1715 (N_1715,N_1526,N_1510);
nand U1716 (N_1716,N_1543,N_1517);
nor U1717 (N_1717,N_1467,N_1450);
xor U1718 (N_1718,N_1431,N_1465);
or U1719 (N_1719,N_1569,N_1419);
nand U1720 (N_1720,N_1452,N_1467);
and U1721 (N_1721,N_1483,N_1448);
and U1722 (N_1722,N_1403,N_1551);
and U1723 (N_1723,N_1410,N_1455);
nor U1724 (N_1724,N_1486,N_1481);
and U1725 (N_1725,N_1576,N_1411);
or U1726 (N_1726,N_1457,N_1541);
or U1727 (N_1727,N_1524,N_1473);
or U1728 (N_1728,N_1458,N_1511);
nand U1729 (N_1729,N_1464,N_1447);
and U1730 (N_1730,N_1460,N_1410);
nor U1731 (N_1731,N_1462,N_1413);
nor U1732 (N_1732,N_1421,N_1498);
or U1733 (N_1733,N_1464,N_1451);
or U1734 (N_1734,N_1472,N_1440);
nand U1735 (N_1735,N_1420,N_1538);
and U1736 (N_1736,N_1578,N_1457);
or U1737 (N_1737,N_1511,N_1420);
or U1738 (N_1738,N_1558,N_1465);
nor U1739 (N_1739,N_1495,N_1470);
xor U1740 (N_1740,N_1510,N_1567);
and U1741 (N_1741,N_1586,N_1430);
or U1742 (N_1742,N_1550,N_1490);
nand U1743 (N_1743,N_1410,N_1432);
and U1744 (N_1744,N_1407,N_1551);
nand U1745 (N_1745,N_1466,N_1565);
nor U1746 (N_1746,N_1494,N_1588);
xor U1747 (N_1747,N_1453,N_1507);
nor U1748 (N_1748,N_1442,N_1592);
and U1749 (N_1749,N_1550,N_1475);
and U1750 (N_1750,N_1551,N_1527);
or U1751 (N_1751,N_1598,N_1509);
nor U1752 (N_1752,N_1439,N_1476);
and U1753 (N_1753,N_1518,N_1415);
or U1754 (N_1754,N_1561,N_1495);
xnor U1755 (N_1755,N_1460,N_1498);
and U1756 (N_1756,N_1483,N_1460);
nand U1757 (N_1757,N_1404,N_1532);
or U1758 (N_1758,N_1426,N_1458);
xor U1759 (N_1759,N_1509,N_1494);
xor U1760 (N_1760,N_1555,N_1554);
xor U1761 (N_1761,N_1478,N_1468);
xor U1762 (N_1762,N_1403,N_1458);
nand U1763 (N_1763,N_1531,N_1548);
nand U1764 (N_1764,N_1439,N_1457);
xnor U1765 (N_1765,N_1424,N_1501);
xor U1766 (N_1766,N_1570,N_1508);
nor U1767 (N_1767,N_1562,N_1432);
nor U1768 (N_1768,N_1483,N_1522);
and U1769 (N_1769,N_1574,N_1517);
nand U1770 (N_1770,N_1553,N_1454);
nor U1771 (N_1771,N_1415,N_1492);
and U1772 (N_1772,N_1423,N_1528);
nor U1773 (N_1773,N_1468,N_1543);
nand U1774 (N_1774,N_1463,N_1568);
and U1775 (N_1775,N_1528,N_1565);
nand U1776 (N_1776,N_1494,N_1593);
xor U1777 (N_1777,N_1413,N_1580);
or U1778 (N_1778,N_1472,N_1540);
nor U1779 (N_1779,N_1424,N_1580);
xnor U1780 (N_1780,N_1508,N_1425);
xor U1781 (N_1781,N_1507,N_1511);
or U1782 (N_1782,N_1537,N_1461);
or U1783 (N_1783,N_1433,N_1507);
xnor U1784 (N_1784,N_1533,N_1566);
nor U1785 (N_1785,N_1424,N_1596);
and U1786 (N_1786,N_1520,N_1546);
xnor U1787 (N_1787,N_1510,N_1493);
nand U1788 (N_1788,N_1468,N_1527);
or U1789 (N_1789,N_1519,N_1500);
or U1790 (N_1790,N_1551,N_1482);
or U1791 (N_1791,N_1430,N_1423);
xnor U1792 (N_1792,N_1548,N_1564);
xor U1793 (N_1793,N_1569,N_1585);
nand U1794 (N_1794,N_1553,N_1445);
xnor U1795 (N_1795,N_1437,N_1525);
xnor U1796 (N_1796,N_1410,N_1418);
or U1797 (N_1797,N_1444,N_1598);
or U1798 (N_1798,N_1599,N_1428);
nor U1799 (N_1799,N_1506,N_1505);
nor U1800 (N_1800,N_1763,N_1650);
or U1801 (N_1801,N_1607,N_1781);
xor U1802 (N_1802,N_1647,N_1728);
and U1803 (N_1803,N_1768,N_1686);
nor U1804 (N_1804,N_1762,N_1672);
or U1805 (N_1805,N_1644,N_1670);
xnor U1806 (N_1806,N_1733,N_1614);
nand U1807 (N_1807,N_1677,N_1664);
nor U1808 (N_1808,N_1718,N_1641);
or U1809 (N_1809,N_1639,N_1631);
or U1810 (N_1810,N_1694,N_1642);
xnor U1811 (N_1811,N_1712,N_1615);
nand U1812 (N_1812,N_1788,N_1674);
xnor U1813 (N_1813,N_1665,N_1721);
xnor U1814 (N_1814,N_1635,N_1740);
nor U1815 (N_1815,N_1692,N_1743);
or U1816 (N_1816,N_1629,N_1682);
or U1817 (N_1817,N_1722,N_1778);
and U1818 (N_1818,N_1796,N_1646);
nand U1819 (N_1819,N_1734,N_1689);
nand U1820 (N_1820,N_1774,N_1754);
nor U1821 (N_1821,N_1795,N_1640);
nand U1822 (N_1822,N_1663,N_1704);
and U1823 (N_1823,N_1643,N_1793);
and U1824 (N_1824,N_1693,N_1736);
nand U1825 (N_1825,N_1758,N_1726);
xnor U1826 (N_1826,N_1713,N_1764);
xnor U1827 (N_1827,N_1730,N_1619);
or U1828 (N_1828,N_1747,N_1741);
nand U1829 (N_1829,N_1746,N_1757);
nand U1830 (N_1830,N_1691,N_1675);
and U1831 (N_1831,N_1613,N_1794);
or U1832 (N_1832,N_1773,N_1652);
and U1833 (N_1833,N_1779,N_1661);
nor U1834 (N_1834,N_1751,N_1777);
and U1835 (N_1835,N_1660,N_1784);
xor U1836 (N_1836,N_1605,N_1749);
nor U1837 (N_1837,N_1767,N_1761);
xor U1838 (N_1838,N_1739,N_1744);
or U1839 (N_1839,N_1703,N_1604);
and U1840 (N_1840,N_1628,N_1745);
nor U1841 (N_1841,N_1676,N_1798);
and U1842 (N_1842,N_1651,N_1624);
nand U1843 (N_1843,N_1667,N_1603);
xnor U1844 (N_1844,N_1632,N_1708);
xnor U1845 (N_1845,N_1699,N_1627);
nand U1846 (N_1846,N_1724,N_1750);
or U1847 (N_1847,N_1732,N_1654);
nor U1848 (N_1848,N_1620,N_1738);
nand U1849 (N_1849,N_1707,N_1702);
xnor U1850 (N_1850,N_1717,N_1797);
or U1851 (N_1851,N_1709,N_1601);
nand U1852 (N_1852,N_1617,N_1727);
xor U1853 (N_1853,N_1659,N_1714);
nand U1854 (N_1854,N_1690,N_1783);
or U1855 (N_1855,N_1716,N_1671);
and U1856 (N_1856,N_1785,N_1735);
nor U1857 (N_1857,N_1656,N_1658);
nand U1858 (N_1858,N_1678,N_1600);
nor U1859 (N_1859,N_1633,N_1759);
nor U1860 (N_1860,N_1683,N_1696);
nor U1861 (N_1861,N_1653,N_1711);
nand U1862 (N_1862,N_1637,N_1799);
nand U1863 (N_1863,N_1725,N_1706);
or U1864 (N_1864,N_1657,N_1772);
and U1865 (N_1865,N_1681,N_1748);
xor U1866 (N_1866,N_1623,N_1626);
xnor U1867 (N_1867,N_1634,N_1723);
nor U1868 (N_1868,N_1737,N_1775);
or U1869 (N_1869,N_1679,N_1780);
nor U1870 (N_1870,N_1666,N_1755);
xor U1871 (N_1871,N_1770,N_1673);
xor U1872 (N_1872,N_1752,N_1649);
and U1873 (N_1873,N_1610,N_1792);
nand U1874 (N_1874,N_1606,N_1729);
nor U1875 (N_1875,N_1645,N_1700);
xnor U1876 (N_1876,N_1612,N_1611);
nor U1877 (N_1877,N_1636,N_1687);
nor U1878 (N_1878,N_1662,N_1705);
or U1879 (N_1879,N_1715,N_1622);
nor U1880 (N_1880,N_1688,N_1731);
or U1881 (N_1881,N_1720,N_1680);
or U1882 (N_1882,N_1791,N_1602);
nor U1883 (N_1883,N_1685,N_1765);
xor U1884 (N_1884,N_1608,N_1766);
nor U1885 (N_1885,N_1790,N_1756);
xor U1886 (N_1886,N_1753,N_1668);
nand U1887 (N_1887,N_1776,N_1698);
or U1888 (N_1888,N_1625,N_1648);
and U1889 (N_1889,N_1655,N_1669);
or U1890 (N_1890,N_1782,N_1769);
xnor U1891 (N_1891,N_1760,N_1786);
or U1892 (N_1892,N_1701,N_1719);
xnor U1893 (N_1893,N_1695,N_1609);
and U1894 (N_1894,N_1771,N_1621);
nand U1895 (N_1895,N_1742,N_1630);
or U1896 (N_1896,N_1710,N_1638);
xor U1897 (N_1897,N_1789,N_1618);
nand U1898 (N_1898,N_1787,N_1616);
or U1899 (N_1899,N_1684,N_1697);
nor U1900 (N_1900,N_1731,N_1601);
or U1901 (N_1901,N_1745,N_1728);
nand U1902 (N_1902,N_1679,N_1645);
xnor U1903 (N_1903,N_1783,N_1705);
xnor U1904 (N_1904,N_1763,N_1743);
xnor U1905 (N_1905,N_1672,N_1736);
xor U1906 (N_1906,N_1760,N_1700);
nor U1907 (N_1907,N_1766,N_1698);
nand U1908 (N_1908,N_1666,N_1727);
or U1909 (N_1909,N_1619,N_1773);
nor U1910 (N_1910,N_1612,N_1693);
or U1911 (N_1911,N_1700,N_1661);
xnor U1912 (N_1912,N_1629,N_1698);
nor U1913 (N_1913,N_1626,N_1647);
nand U1914 (N_1914,N_1656,N_1769);
or U1915 (N_1915,N_1717,N_1669);
xor U1916 (N_1916,N_1615,N_1794);
and U1917 (N_1917,N_1775,N_1781);
and U1918 (N_1918,N_1794,N_1682);
xor U1919 (N_1919,N_1638,N_1628);
nor U1920 (N_1920,N_1646,N_1604);
or U1921 (N_1921,N_1600,N_1617);
nor U1922 (N_1922,N_1625,N_1668);
or U1923 (N_1923,N_1722,N_1718);
xor U1924 (N_1924,N_1689,N_1703);
or U1925 (N_1925,N_1698,N_1792);
and U1926 (N_1926,N_1679,N_1717);
nor U1927 (N_1927,N_1787,N_1673);
nand U1928 (N_1928,N_1724,N_1785);
or U1929 (N_1929,N_1630,N_1741);
nor U1930 (N_1930,N_1773,N_1662);
or U1931 (N_1931,N_1785,N_1687);
or U1932 (N_1932,N_1750,N_1628);
nand U1933 (N_1933,N_1728,N_1765);
or U1934 (N_1934,N_1797,N_1781);
nor U1935 (N_1935,N_1676,N_1664);
xor U1936 (N_1936,N_1609,N_1765);
nand U1937 (N_1937,N_1666,N_1723);
or U1938 (N_1938,N_1768,N_1718);
or U1939 (N_1939,N_1684,N_1688);
xnor U1940 (N_1940,N_1747,N_1613);
xnor U1941 (N_1941,N_1722,N_1782);
xor U1942 (N_1942,N_1615,N_1620);
xnor U1943 (N_1943,N_1774,N_1705);
nand U1944 (N_1944,N_1740,N_1788);
and U1945 (N_1945,N_1666,N_1753);
nor U1946 (N_1946,N_1766,N_1691);
xnor U1947 (N_1947,N_1673,N_1680);
nand U1948 (N_1948,N_1761,N_1783);
and U1949 (N_1949,N_1707,N_1681);
xor U1950 (N_1950,N_1651,N_1640);
nand U1951 (N_1951,N_1671,N_1774);
or U1952 (N_1952,N_1618,N_1794);
or U1953 (N_1953,N_1713,N_1681);
xor U1954 (N_1954,N_1694,N_1725);
nor U1955 (N_1955,N_1748,N_1728);
xnor U1956 (N_1956,N_1666,N_1678);
xnor U1957 (N_1957,N_1792,N_1681);
and U1958 (N_1958,N_1783,N_1620);
and U1959 (N_1959,N_1749,N_1643);
or U1960 (N_1960,N_1797,N_1778);
and U1961 (N_1961,N_1672,N_1758);
nor U1962 (N_1962,N_1781,N_1637);
nor U1963 (N_1963,N_1676,N_1797);
or U1964 (N_1964,N_1601,N_1621);
xor U1965 (N_1965,N_1776,N_1673);
xor U1966 (N_1966,N_1790,N_1775);
and U1967 (N_1967,N_1756,N_1635);
xnor U1968 (N_1968,N_1757,N_1641);
nand U1969 (N_1969,N_1718,N_1640);
and U1970 (N_1970,N_1637,N_1674);
or U1971 (N_1971,N_1692,N_1760);
or U1972 (N_1972,N_1727,N_1642);
or U1973 (N_1973,N_1759,N_1674);
or U1974 (N_1974,N_1691,N_1795);
xnor U1975 (N_1975,N_1630,N_1603);
and U1976 (N_1976,N_1622,N_1745);
xnor U1977 (N_1977,N_1730,N_1742);
xor U1978 (N_1978,N_1626,N_1778);
nand U1979 (N_1979,N_1715,N_1781);
and U1980 (N_1980,N_1617,N_1768);
or U1981 (N_1981,N_1621,N_1712);
nor U1982 (N_1982,N_1768,N_1794);
or U1983 (N_1983,N_1605,N_1607);
nor U1984 (N_1984,N_1652,N_1690);
and U1985 (N_1985,N_1777,N_1654);
nor U1986 (N_1986,N_1742,N_1645);
xnor U1987 (N_1987,N_1742,N_1702);
nand U1988 (N_1988,N_1737,N_1647);
nor U1989 (N_1989,N_1761,N_1670);
and U1990 (N_1990,N_1759,N_1762);
and U1991 (N_1991,N_1603,N_1777);
nor U1992 (N_1992,N_1630,N_1665);
or U1993 (N_1993,N_1652,N_1745);
or U1994 (N_1994,N_1743,N_1752);
nand U1995 (N_1995,N_1624,N_1763);
nand U1996 (N_1996,N_1779,N_1636);
or U1997 (N_1997,N_1699,N_1758);
nand U1998 (N_1998,N_1789,N_1651);
nor U1999 (N_1999,N_1647,N_1684);
or U2000 (N_2000,N_1846,N_1928);
or U2001 (N_2001,N_1946,N_1857);
nor U2002 (N_2002,N_1934,N_1949);
nand U2003 (N_2003,N_1966,N_1840);
and U2004 (N_2004,N_1850,N_1969);
nand U2005 (N_2005,N_1999,N_1916);
nand U2006 (N_2006,N_1906,N_1953);
and U2007 (N_2007,N_1835,N_1820);
and U2008 (N_2008,N_1829,N_1825);
or U2009 (N_2009,N_1819,N_1903);
xnor U2010 (N_2010,N_1871,N_1849);
xor U2011 (N_2011,N_1884,N_1833);
nand U2012 (N_2012,N_1892,N_1875);
nor U2013 (N_2013,N_1831,N_1885);
and U2014 (N_2014,N_1910,N_1826);
or U2015 (N_2015,N_1914,N_1842);
nor U2016 (N_2016,N_1948,N_1951);
and U2017 (N_2017,N_1919,N_1991);
and U2018 (N_2018,N_1856,N_1872);
nand U2019 (N_2019,N_1974,N_1907);
nor U2020 (N_2020,N_1924,N_1945);
and U2021 (N_2021,N_1947,N_1971);
or U2022 (N_2022,N_1967,N_1808);
and U2023 (N_2023,N_1834,N_1845);
nand U2024 (N_2024,N_1898,N_1930);
nand U2025 (N_2025,N_1902,N_1983);
nor U2026 (N_2026,N_1932,N_1937);
and U2027 (N_2027,N_1848,N_1805);
nor U2028 (N_2028,N_1874,N_1979);
and U2029 (N_2029,N_1844,N_1908);
and U2030 (N_2030,N_1873,N_1896);
and U2031 (N_2031,N_1918,N_1905);
nor U2032 (N_2032,N_1968,N_1801);
xnor U2033 (N_2033,N_1977,N_1922);
or U2034 (N_2034,N_1950,N_1828);
nor U2035 (N_2035,N_1882,N_1994);
nor U2036 (N_2036,N_1867,N_1992);
nand U2037 (N_2037,N_1926,N_1901);
or U2038 (N_2038,N_1890,N_1889);
nor U2039 (N_2039,N_1824,N_1866);
or U2040 (N_2040,N_1847,N_1812);
nor U2041 (N_2041,N_1818,N_1897);
or U2042 (N_2042,N_1855,N_1931);
and U2043 (N_2043,N_1912,N_1927);
and U2044 (N_2044,N_1813,N_1956);
nand U2045 (N_2045,N_1917,N_1870);
and U2046 (N_2046,N_1900,N_1809);
and U2047 (N_2047,N_1864,N_1839);
xnor U2048 (N_2048,N_1877,N_1802);
xnor U2049 (N_2049,N_1958,N_1935);
nor U2050 (N_2050,N_1814,N_1811);
nor U2051 (N_2051,N_1880,N_1806);
nor U2052 (N_2052,N_1942,N_1904);
nor U2053 (N_2053,N_1973,N_1995);
or U2054 (N_2054,N_1876,N_1925);
nand U2055 (N_2055,N_1881,N_1861);
and U2056 (N_2056,N_1920,N_1807);
nand U2057 (N_2057,N_1938,N_1982);
or U2058 (N_2058,N_1888,N_1921);
and U2059 (N_2059,N_1993,N_1827);
nand U2060 (N_2060,N_1954,N_1821);
nor U2061 (N_2061,N_1936,N_1963);
and U2062 (N_2062,N_1998,N_1929);
and U2063 (N_2063,N_1817,N_1863);
and U2064 (N_2064,N_1943,N_1883);
nor U2065 (N_2065,N_1975,N_1838);
or U2066 (N_2066,N_1972,N_1816);
nor U2067 (N_2067,N_1852,N_1862);
xor U2068 (N_2068,N_1894,N_1887);
nor U2069 (N_2069,N_1976,N_1980);
or U2070 (N_2070,N_1803,N_1886);
and U2071 (N_2071,N_1843,N_1981);
xnor U2072 (N_2072,N_1962,N_1990);
xor U2073 (N_2073,N_1899,N_1869);
nor U2074 (N_2074,N_1959,N_1858);
nor U2075 (N_2075,N_1851,N_1957);
nand U2076 (N_2076,N_1815,N_1822);
xnor U2077 (N_2077,N_1961,N_1960);
or U2078 (N_2078,N_1952,N_1800);
nand U2079 (N_2079,N_1923,N_1964);
and U2080 (N_2080,N_1911,N_1988);
nor U2081 (N_2081,N_1804,N_1810);
xor U2082 (N_2082,N_1879,N_1895);
nor U2083 (N_2083,N_1955,N_1891);
nor U2084 (N_2084,N_1933,N_1941);
nor U2085 (N_2085,N_1913,N_1984);
nor U2086 (N_2086,N_1978,N_1985);
nand U2087 (N_2087,N_1996,N_1860);
and U2088 (N_2088,N_1986,N_1832);
nor U2089 (N_2089,N_1893,N_1909);
and U2090 (N_2090,N_1830,N_1965);
nand U2091 (N_2091,N_1865,N_1854);
nor U2092 (N_2092,N_1859,N_1970);
or U2093 (N_2093,N_1853,N_1836);
nand U2094 (N_2094,N_1868,N_1939);
or U2095 (N_2095,N_1841,N_1878);
or U2096 (N_2096,N_1823,N_1987);
xor U2097 (N_2097,N_1997,N_1940);
and U2098 (N_2098,N_1944,N_1915);
nand U2099 (N_2099,N_1837,N_1989);
nor U2100 (N_2100,N_1975,N_1969);
or U2101 (N_2101,N_1884,N_1971);
nand U2102 (N_2102,N_1852,N_1850);
and U2103 (N_2103,N_1987,N_1968);
nand U2104 (N_2104,N_1812,N_1883);
nor U2105 (N_2105,N_1973,N_1849);
and U2106 (N_2106,N_1875,N_1957);
nand U2107 (N_2107,N_1896,N_1812);
or U2108 (N_2108,N_1864,N_1925);
nor U2109 (N_2109,N_1870,N_1876);
or U2110 (N_2110,N_1938,N_1941);
and U2111 (N_2111,N_1973,N_1981);
or U2112 (N_2112,N_1963,N_1907);
or U2113 (N_2113,N_1895,N_1848);
and U2114 (N_2114,N_1814,N_1846);
nand U2115 (N_2115,N_1994,N_1885);
nor U2116 (N_2116,N_1864,N_1947);
or U2117 (N_2117,N_1951,N_1846);
nor U2118 (N_2118,N_1964,N_1957);
nand U2119 (N_2119,N_1993,N_1835);
and U2120 (N_2120,N_1914,N_1812);
nor U2121 (N_2121,N_1825,N_1933);
and U2122 (N_2122,N_1900,N_1800);
nand U2123 (N_2123,N_1861,N_1835);
and U2124 (N_2124,N_1951,N_1910);
nor U2125 (N_2125,N_1980,N_1951);
and U2126 (N_2126,N_1918,N_1965);
xor U2127 (N_2127,N_1956,N_1892);
nand U2128 (N_2128,N_1984,N_1903);
nor U2129 (N_2129,N_1853,N_1834);
nand U2130 (N_2130,N_1925,N_1866);
xnor U2131 (N_2131,N_1874,N_1917);
nand U2132 (N_2132,N_1891,N_1929);
xor U2133 (N_2133,N_1806,N_1879);
or U2134 (N_2134,N_1963,N_1932);
xnor U2135 (N_2135,N_1814,N_1872);
xor U2136 (N_2136,N_1895,N_1974);
or U2137 (N_2137,N_1994,N_1806);
nor U2138 (N_2138,N_1909,N_1913);
and U2139 (N_2139,N_1815,N_1904);
nand U2140 (N_2140,N_1991,N_1974);
nor U2141 (N_2141,N_1918,N_1933);
nand U2142 (N_2142,N_1811,N_1982);
nand U2143 (N_2143,N_1814,N_1915);
or U2144 (N_2144,N_1996,N_1884);
or U2145 (N_2145,N_1932,N_1964);
and U2146 (N_2146,N_1992,N_1887);
xor U2147 (N_2147,N_1986,N_1888);
or U2148 (N_2148,N_1823,N_1990);
xor U2149 (N_2149,N_1935,N_1936);
nand U2150 (N_2150,N_1853,N_1905);
nand U2151 (N_2151,N_1937,N_1997);
and U2152 (N_2152,N_1863,N_1896);
nor U2153 (N_2153,N_1801,N_1958);
or U2154 (N_2154,N_1995,N_1985);
or U2155 (N_2155,N_1931,N_1969);
nor U2156 (N_2156,N_1816,N_1836);
nand U2157 (N_2157,N_1901,N_1933);
or U2158 (N_2158,N_1812,N_1901);
nand U2159 (N_2159,N_1871,N_1938);
nor U2160 (N_2160,N_1949,N_1844);
or U2161 (N_2161,N_1883,N_1907);
nand U2162 (N_2162,N_1829,N_1891);
and U2163 (N_2163,N_1814,N_1951);
and U2164 (N_2164,N_1940,N_1983);
nor U2165 (N_2165,N_1877,N_1892);
xnor U2166 (N_2166,N_1934,N_1886);
nor U2167 (N_2167,N_1962,N_1866);
nand U2168 (N_2168,N_1844,N_1901);
xnor U2169 (N_2169,N_1989,N_1822);
and U2170 (N_2170,N_1940,N_1911);
nor U2171 (N_2171,N_1848,N_1820);
xor U2172 (N_2172,N_1989,N_1883);
nor U2173 (N_2173,N_1938,N_1875);
nor U2174 (N_2174,N_1959,N_1995);
xnor U2175 (N_2175,N_1838,N_1974);
nand U2176 (N_2176,N_1805,N_1995);
nor U2177 (N_2177,N_1942,N_1957);
nand U2178 (N_2178,N_1896,N_1977);
xor U2179 (N_2179,N_1843,N_1855);
xor U2180 (N_2180,N_1926,N_1887);
or U2181 (N_2181,N_1864,N_1934);
nand U2182 (N_2182,N_1814,N_1829);
nand U2183 (N_2183,N_1963,N_1844);
nand U2184 (N_2184,N_1991,N_1806);
nor U2185 (N_2185,N_1881,N_1967);
nor U2186 (N_2186,N_1836,N_1870);
xnor U2187 (N_2187,N_1956,N_1984);
and U2188 (N_2188,N_1934,N_1861);
xor U2189 (N_2189,N_1852,N_1954);
or U2190 (N_2190,N_1975,N_1963);
nor U2191 (N_2191,N_1938,N_1940);
and U2192 (N_2192,N_1855,N_1892);
nor U2193 (N_2193,N_1921,N_1974);
nor U2194 (N_2194,N_1897,N_1827);
nor U2195 (N_2195,N_1862,N_1951);
nand U2196 (N_2196,N_1844,N_1862);
xnor U2197 (N_2197,N_1983,N_1924);
nor U2198 (N_2198,N_1895,N_1983);
or U2199 (N_2199,N_1965,N_1888);
nor U2200 (N_2200,N_2117,N_2155);
xor U2201 (N_2201,N_2104,N_2189);
nand U2202 (N_2202,N_2095,N_2183);
nor U2203 (N_2203,N_2164,N_2100);
or U2204 (N_2204,N_2083,N_2181);
xnor U2205 (N_2205,N_2122,N_2107);
or U2206 (N_2206,N_2076,N_2078);
nor U2207 (N_2207,N_2132,N_2154);
xor U2208 (N_2208,N_2199,N_2144);
xor U2209 (N_2209,N_2035,N_2176);
xnor U2210 (N_2210,N_2065,N_2007);
and U2211 (N_2211,N_2170,N_2111);
nor U2212 (N_2212,N_2055,N_2182);
xnor U2213 (N_2213,N_2038,N_2051);
or U2214 (N_2214,N_2008,N_2019);
nor U2215 (N_2215,N_2151,N_2184);
nand U2216 (N_2216,N_2172,N_2163);
or U2217 (N_2217,N_2090,N_2006);
or U2218 (N_2218,N_2190,N_2198);
nand U2219 (N_2219,N_2021,N_2020);
or U2220 (N_2220,N_2071,N_2092);
or U2221 (N_2221,N_2012,N_2110);
nor U2222 (N_2222,N_2194,N_2015);
nand U2223 (N_2223,N_2033,N_2040);
nor U2224 (N_2224,N_2057,N_2157);
and U2225 (N_2225,N_2150,N_2197);
xnor U2226 (N_2226,N_2102,N_2048);
xnor U2227 (N_2227,N_2084,N_2081);
and U2228 (N_2228,N_2034,N_2074);
nand U2229 (N_2229,N_2106,N_2130);
nor U2230 (N_2230,N_2050,N_2060);
or U2231 (N_2231,N_2041,N_2147);
or U2232 (N_2232,N_2022,N_2175);
nand U2233 (N_2233,N_2113,N_2024);
xnor U2234 (N_2234,N_2016,N_2145);
nand U2235 (N_2235,N_2143,N_2185);
xnor U2236 (N_2236,N_2029,N_2064);
xor U2237 (N_2237,N_2067,N_2077);
or U2238 (N_2238,N_2001,N_2075);
nor U2239 (N_2239,N_2186,N_2085);
and U2240 (N_2240,N_2166,N_2042);
xnor U2241 (N_2241,N_2153,N_2097);
or U2242 (N_2242,N_2121,N_2148);
xnor U2243 (N_2243,N_2003,N_2062);
and U2244 (N_2244,N_2039,N_2037);
or U2245 (N_2245,N_2160,N_2188);
nand U2246 (N_2246,N_2080,N_2125);
and U2247 (N_2247,N_2032,N_2096);
nand U2248 (N_2248,N_2017,N_2168);
xnor U2249 (N_2249,N_2028,N_2049);
nor U2250 (N_2250,N_2103,N_2177);
nor U2251 (N_2251,N_2058,N_2046);
nor U2252 (N_2252,N_2123,N_2192);
or U2253 (N_2253,N_2178,N_2161);
or U2254 (N_2254,N_2089,N_2127);
and U2255 (N_2255,N_2133,N_2066);
nor U2256 (N_2256,N_2099,N_2101);
and U2257 (N_2257,N_2068,N_2180);
xnor U2258 (N_2258,N_2105,N_2138);
nand U2259 (N_2259,N_2027,N_2165);
and U2260 (N_2260,N_2052,N_2069);
nand U2261 (N_2261,N_2093,N_2056);
nor U2262 (N_2262,N_2043,N_2174);
nor U2263 (N_2263,N_2087,N_2082);
nand U2264 (N_2264,N_2005,N_2091);
xor U2265 (N_2265,N_2023,N_2152);
and U2266 (N_2266,N_2094,N_2187);
or U2267 (N_2267,N_2061,N_2010);
nor U2268 (N_2268,N_2169,N_2195);
and U2269 (N_2269,N_2119,N_2004);
and U2270 (N_2270,N_2002,N_2156);
nand U2271 (N_2271,N_2079,N_2129);
nor U2272 (N_2272,N_2149,N_2126);
and U2273 (N_2273,N_2118,N_2128);
or U2274 (N_2274,N_2014,N_2116);
nand U2275 (N_2275,N_2135,N_2109);
nor U2276 (N_2276,N_2011,N_2136);
nand U2277 (N_2277,N_2179,N_2072);
nor U2278 (N_2278,N_2114,N_2086);
xor U2279 (N_2279,N_2025,N_2088);
nor U2280 (N_2280,N_2115,N_2018);
and U2281 (N_2281,N_2070,N_2054);
nor U2282 (N_2282,N_2059,N_2073);
nand U2283 (N_2283,N_2162,N_2026);
xor U2284 (N_2284,N_2013,N_2063);
or U2285 (N_2285,N_2098,N_2139);
nor U2286 (N_2286,N_2036,N_2158);
nand U2287 (N_2287,N_2131,N_2031);
and U2288 (N_2288,N_2124,N_2159);
and U2289 (N_2289,N_2108,N_2009);
nand U2290 (N_2290,N_2140,N_2171);
xnor U2291 (N_2291,N_2030,N_2193);
and U2292 (N_2292,N_2044,N_2000);
nor U2293 (N_2293,N_2141,N_2191);
and U2294 (N_2294,N_2053,N_2112);
nor U2295 (N_2295,N_2134,N_2196);
or U2296 (N_2296,N_2045,N_2047);
nor U2297 (N_2297,N_2142,N_2146);
or U2298 (N_2298,N_2137,N_2173);
or U2299 (N_2299,N_2120,N_2167);
and U2300 (N_2300,N_2173,N_2131);
nand U2301 (N_2301,N_2135,N_2160);
and U2302 (N_2302,N_2190,N_2073);
and U2303 (N_2303,N_2057,N_2092);
nand U2304 (N_2304,N_2129,N_2001);
and U2305 (N_2305,N_2170,N_2086);
nor U2306 (N_2306,N_2158,N_2174);
or U2307 (N_2307,N_2162,N_2172);
nor U2308 (N_2308,N_2030,N_2176);
or U2309 (N_2309,N_2074,N_2190);
nand U2310 (N_2310,N_2031,N_2136);
or U2311 (N_2311,N_2190,N_2100);
or U2312 (N_2312,N_2042,N_2126);
nand U2313 (N_2313,N_2150,N_2194);
and U2314 (N_2314,N_2079,N_2107);
nand U2315 (N_2315,N_2164,N_2009);
and U2316 (N_2316,N_2078,N_2100);
nand U2317 (N_2317,N_2159,N_2180);
nor U2318 (N_2318,N_2108,N_2129);
nand U2319 (N_2319,N_2054,N_2163);
nor U2320 (N_2320,N_2171,N_2153);
xnor U2321 (N_2321,N_2136,N_2034);
xor U2322 (N_2322,N_2045,N_2126);
and U2323 (N_2323,N_2067,N_2193);
and U2324 (N_2324,N_2192,N_2029);
nor U2325 (N_2325,N_2171,N_2024);
nor U2326 (N_2326,N_2038,N_2080);
nor U2327 (N_2327,N_2003,N_2087);
and U2328 (N_2328,N_2085,N_2005);
nor U2329 (N_2329,N_2164,N_2128);
and U2330 (N_2330,N_2123,N_2155);
xor U2331 (N_2331,N_2017,N_2111);
and U2332 (N_2332,N_2185,N_2006);
and U2333 (N_2333,N_2184,N_2043);
or U2334 (N_2334,N_2178,N_2056);
or U2335 (N_2335,N_2085,N_2025);
xnor U2336 (N_2336,N_2092,N_2111);
and U2337 (N_2337,N_2132,N_2139);
nand U2338 (N_2338,N_2029,N_2118);
nand U2339 (N_2339,N_2111,N_2108);
xor U2340 (N_2340,N_2041,N_2189);
and U2341 (N_2341,N_2122,N_2110);
or U2342 (N_2342,N_2000,N_2002);
and U2343 (N_2343,N_2157,N_2100);
nand U2344 (N_2344,N_2002,N_2078);
or U2345 (N_2345,N_2088,N_2143);
xnor U2346 (N_2346,N_2180,N_2121);
nor U2347 (N_2347,N_2136,N_2177);
nand U2348 (N_2348,N_2110,N_2107);
nand U2349 (N_2349,N_2114,N_2012);
and U2350 (N_2350,N_2091,N_2162);
nor U2351 (N_2351,N_2060,N_2072);
nand U2352 (N_2352,N_2077,N_2124);
xor U2353 (N_2353,N_2052,N_2007);
xor U2354 (N_2354,N_2094,N_2106);
nand U2355 (N_2355,N_2066,N_2054);
nand U2356 (N_2356,N_2126,N_2179);
and U2357 (N_2357,N_2178,N_2094);
and U2358 (N_2358,N_2027,N_2082);
nand U2359 (N_2359,N_2039,N_2040);
or U2360 (N_2360,N_2130,N_2177);
nand U2361 (N_2361,N_2004,N_2172);
nand U2362 (N_2362,N_2042,N_2151);
and U2363 (N_2363,N_2001,N_2133);
xnor U2364 (N_2364,N_2125,N_2016);
nor U2365 (N_2365,N_2047,N_2190);
or U2366 (N_2366,N_2020,N_2178);
nand U2367 (N_2367,N_2107,N_2125);
and U2368 (N_2368,N_2031,N_2199);
nand U2369 (N_2369,N_2022,N_2126);
and U2370 (N_2370,N_2197,N_2114);
or U2371 (N_2371,N_2049,N_2146);
xnor U2372 (N_2372,N_2105,N_2119);
nor U2373 (N_2373,N_2072,N_2027);
xnor U2374 (N_2374,N_2107,N_2084);
or U2375 (N_2375,N_2048,N_2095);
nand U2376 (N_2376,N_2183,N_2093);
or U2377 (N_2377,N_2080,N_2133);
xnor U2378 (N_2378,N_2146,N_2038);
nor U2379 (N_2379,N_2054,N_2062);
nor U2380 (N_2380,N_2160,N_2066);
or U2381 (N_2381,N_2089,N_2071);
nor U2382 (N_2382,N_2178,N_2177);
or U2383 (N_2383,N_2067,N_2013);
xnor U2384 (N_2384,N_2061,N_2128);
nand U2385 (N_2385,N_2162,N_2130);
nand U2386 (N_2386,N_2156,N_2131);
nor U2387 (N_2387,N_2100,N_2085);
and U2388 (N_2388,N_2007,N_2016);
xor U2389 (N_2389,N_2117,N_2186);
or U2390 (N_2390,N_2116,N_2155);
and U2391 (N_2391,N_2000,N_2152);
nor U2392 (N_2392,N_2039,N_2098);
or U2393 (N_2393,N_2195,N_2118);
or U2394 (N_2394,N_2031,N_2160);
and U2395 (N_2395,N_2154,N_2104);
nand U2396 (N_2396,N_2159,N_2106);
xor U2397 (N_2397,N_2107,N_2058);
xor U2398 (N_2398,N_2069,N_2041);
nand U2399 (N_2399,N_2142,N_2106);
and U2400 (N_2400,N_2314,N_2323);
or U2401 (N_2401,N_2292,N_2376);
nand U2402 (N_2402,N_2334,N_2367);
nor U2403 (N_2403,N_2229,N_2250);
and U2404 (N_2404,N_2245,N_2386);
nand U2405 (N_2405,N_2224,N_2311);
and U2406 (N_2406,N_2329,N_2393);
nand U2407 (N_2407,N_2330,N_2354);
and U2408 (N_2408,N_2361,N_2228);
and U2409 (N_2409,N_2225,N_2340);
or U2410 (N_2410,N_2304,N_2249);
or U2411 (N_2411,N_2238,N_2379);
xor U2412 (N_2412,N_2370,N_2306);
nor U2413 (N_2413,N_2263,N_2350);
xnor U2414 (N_2414,N_2295,N_2257);
or U2415 (N_2415,N_2273,N_2274);
and U2416 (N_2416,N_2264,N_2384);
xnor U2417 (N_2417,N_2294,N_2365);
xor U2418 (N_2418,N_2328,N_2252);
and U2419 (N_2419,N_2233,N_2355);
or U2420 (N_2420,N_2326,N_2241);
nand U2421 (N_2421,N_2277,N_2254);
nand U2422 (N_2422,N_2286,N_2313);
and U2423 (N_2423,N_2343,N_2259);
nand U2424 (N_2424,N_2247,N_2380);
nor U2425 (N_2425,N_2244,N_2357);
and U2426 (N_2426,N_2303,N_2204);
nor U2427 (N_2427,N_2208,N_2239);
nor U2428 (N_2428,N_2396,N_2375);
nand U2429 (N_2429,N_2287,N_2310);
and U2430 (N_2430,N_2275,N_2280);
and U2431 (N_2431,N_2352,N_2248);
xnor U2432 (N_2432,N_2332,N_2251);
nor U2433 (N_2433,N_2338,N_2305);
and U2434 (N_2434,N_2265,N_2347);
xor U2435 (N_2435,N_2271,N_2337);
xor U2436 (N_2436,N_2267,N_2289);
nor U2437 (N_2437,N_2369,N_2377);
nand U2438 (N_2438,N_2290,N_2363);
nand U2439 (N_2439,N_2336,N_2394);
and U2440 (N_2440,N_2399,N_2344);
xnor U2441 (N_2441,N_2362,N_2381);
or U2442 (N_2442,N_2231,N_2315);
and U2443 (N_2443,N_2378,N_2213);
or U2444 (N_2444,N_2397,N_2335);
xnor U2445 (N_2445,N_2327,N_2206);
or U2446 (N_2446,N_2235,N_2232);
xnor U2447 (N_2447,N_2322,N_2339);
xnor U2448 (N_2448,N_2351,N_2202);
or U2449 (N_2449,N_2388,N_2226);
nand U2450 (N_2450,N_2276,N_2212);
nor U2451 (N_2451,N_2318,N_2308);
and U2452 (N_2452,N_2219,N_2341);
or U2453 (N_2453,N_2392,N_2299);
or U2454 (N_2454,N_2390,N_2227);
or U2455 (N_2455,N_2209,N_2366);
nand U2456 (N_2456,N_2395,N_2266);
xor U2457 (N_2457,N_2312,N_2205);
or U2458 (N_2458,N_2240,N_2359);
xnor U2459 (N_2459,N_2291,N_2372);
nor U2460 (N_2460,N_2391,N_2234);
xnor U2461 (N_2461,N_2387,N_2281);
nand U2462 (N_2462,N_2293,N_2284);
nand U2463 (N_2463,N_2288,N_2298);
nor U2464 (N_2464,N_2279,N_2324);
nand U2465 (N_2465,N_2307,N_2216);
and U2466 (N_2466,N_2223,N_2349);
nand U2467 (N_2467,N_2319,N_2297);
nor U2468 (N_2468,N_2269,N_2382);
or U2469 (N_2469,N_2222,N_2317);
nand U2470 (N_2470,N_2218,N_2353);
xor U2471 (N_2471,N_2220,N_2215);
nor U2472 (N_2472,N_2261,N_2333);
nor U2473 (N_2473,N_2242,N_2368);
or U2474 (N_2474,N_2364,N_2373);
and U2475 (N_2475,N_2296,N_2255);
or U2476 (N_2476,N_2258,N_2383);
nand U2477 (N_2477,N_2316,N_2345);
xnor U2478 (N_2478,N_2360,N_2272);
and U2479 (N_2479,N_2262,N_2270);
xnor U2480 (N_2480,N_2253,N_2260);
and U2481 (N_2481,N_2331,N_2342);
xnor U2482 (N_2482,N_2246,N_2214);
xor U2483 (N_2483,N_2371,N_2309);
or U2484 (N_2484,N_2283,N_2285);
xnor U2485 (N_2485,N_2203,N_2301);
nand U2486 (N_2486,N_2230,N_2217);
and U2487 (N_2487,N_2325,N_2358);
nor U2488 (N_2488,N_2321,N_2243);
nor U2489 (N_2489,N_2320,N_2236);
nor U2490 (N_2490,N_2346,N_2268);
xor U2491 (N_2491,N_2302,N_2282);
or U2492 (N_2492,N_2348,N_2210);
xor U2493 (N_2493,N_2221,N_2200);
and U2494 (N_2494,N_2300,N_2211);
nand U2495 (N_2495,N_2237,N_2389);
nand U2496 (N_2496,N_2256,N_2201);
nand U2497 (N_2497,N_2207,N_2278);
nor U2498 (N_2498,N_2385,N_2398);
or U2499 (N_2499,N_2356,N_2374);
or U2500 (N_2500,N_2232,N_2332);
or U2501 (N_2501,N_2318,N_2270);
nor U2502 (N_2502,N_2363,N_2280);
nor U2503 (N_2503,N_2375,N_2217);
or U2504 (N_2504,N_2237,N_2311);
nand U2505 (N_2505,N_2371,N_2345);
xor U2506 (N_2506,N_2230,N_2283);
nor U2507 (N_2507,N_2293,N_2286);
or U2508 (N_2508,N_2396,N_2394);
nor U2509 (N_2509,N_2352,N_2393);
or U2510 (N_2510,N_2208,N_2323);
nor U2511 (N_2511,N_2341,N_2229);
nor U2512 (N_2512,N_2250,N_2355);
nor U2513 (N_2513,N_2387,N_2279);
and U2514 (N_2514,N_2314,N_2227);
and U2515 (N_2515,N_2304,N_2201);
xor U2516 (N_2516,N_2250,N_2379);
and U2517 (N_2517,N_2212,N_2244);
or U2518 (N_2518,N_2208,N_2214);
nor U2519 (N_2519,N_2227,N_2364);
nand U2520 (N_2520,N_2332,N_2202);
and U2521 (N_2521,N_2368,N_2396);
nor U2522 (N_2522,N_2248,N_2381);
nor U2523 (N_2523,N_2366,N_2230);
nand U2524 (N_2524,N_2205,N_2273);
or U2525 (N_2525,N_2339,N_2203);
or U2526 (N_2526,N_2224,N_2253);
and U2527 (N_2527,N_2324,N_2329);
or U2528 (N_2528,N_2240,N_2323);
nor U2529 (N_2529,N_2268,N_2310);
xor U2530 (N_2530,N_2302,N_2337);
xor U2531 (N_2531,N_2297,N_2280);
xor U2532 (N_2532,N_2208,N_2391);
xnor U2533 (N_2533,N_2339,N_2389);
nand U2534 (N_2534,N_2372,N_2227);
and U2535 (N_2535,N_2335,N_2312);
or U2536 (N_2536,N_2229,N_2331);
or U2537 (N_2537,N_2396,N_2278);
and U2538 (N_2538,N_2376,N_2288);
xnor U2539 (N_2539,N_2368,N_2277);
xnor U2540 (N_2540,N_2328,N_2322);
xor U2541 (N_2541,N_2336,N_2381);
and U2542 (N_2542,N_2286,N_2234);
and U2543 (N_2543,N_2275,N_2346);
nor U2544 (N_2544,N_2229,N_2311);
nand U2545 (N_2545,N_2257,N_2251);
or U2546 (N_2546,N_2271,N_2243);
and U2547 (N_2547,N_2281,N_2265);
and U2548 (N_2548,N_2338,N_2241);
and U2549 (N_2549,N_2212,N_2396);
and U2550 (N_2550,N_2322,N_2211);
nand U2551 (N_2551,N_2250,N_2336);
and U2552 (N_2552,N_2336,N_2327);
nand U2553 (N_2553,N_2395,N_2289);
or U2554 (N_2554,N_2257,N_2256);
xor U2555 (N_2555,N_2364,N_2214);
nor U2556 (N_2556,N_2273,N_2344);
nand U2557 (N_2557,N_2244,N_2373);
or U2558 (N_2558,N_2238,N_2223);
nand U2559 (N_2559,N_2298,N_2259);
nor U2560 (N_2560,N_2362,N_2368);
nor U2561 (N_2561,N_2213,N_2308);
or U2562 (N_2562,N_2344,N_2282);
nand U2563 (N_2563,N_2338,N_2228);
and U2564 (N_2564,N_2270,N_2236);
xnor U2565 (N_2565,N_2216,N_2269);
xnor U2566 (N_2566,N_2381,N_2287);
and U2567 (N_2567,N_2280,N_2397);
nor U2568 (N_2568,N_2230,N_2386);
xor U2569 (N_2569,N_2213,N_2397);
nand U2570 (N_2570,N_2351,N_2233);
nand U2571 (N_2571,N_2206,N_2344);
nand U2572 (N_2572,N_2258,N_2356);
or U2573 (N_2573,N_2248,N_2271);
and U2574 (N_2574,N_2268,N_2236);
nand U2575 (N_2575,N_2337,N_2303);
xnor U2576 (N_2576,N_2294,N_2259);
nand U2577 (N_2577,N_2293,N_2396);
and U2578 (N_2578,N_2353,N_2211);
nor U2579 (N_2579,N_2215,N_2314);
nand U2580 (N_2580,N_2221,N_2344);
and U2581 (N_2581,N_2358,N_2351);
nor U2582 (N_2582,N_2269,N_2220);
or U2583 (N_2583,N_2222,N_2272);
and U2584 (N_2584,N_2309,N_2290);
nor U2585 (N_2585,N_2355,N_2293);
nand U2586 (N_2586,N_2360,N_2280);
and U2587 (N_2587,N_2386,N_2225);
nand U2588 (N_2588,N_2391,N_2255);
xnor U2589 (N_2589,N_2320,N_2327);
and U2590 (N_2590,N_2262,N_2276);
nor U2591 (N_2591,N_2336,N_2259);
nand U2592 (N_2592,N_2349,N_2370);
or U2593 (N_2593,N_2298,N_2339);
and U2594 (N_2594,N_2370,N_2327);
nand U2595 (N_2595,N_2304,N_2275);
nor U2596 (N_2596,N_2228,N_2289);
or U2597 (N_2597,N_2339,N_2321);
nand U2598 (N_2598,N_2259,N_2233);
and U2599 (N_2599,N_2257,N_2264);
or U2600 (N_2600,N_2418,N_2443);
nand U2601 (N_2601,N_2441,N_2448);
nor U2602 (N_2602,N_2425,N_2427);
xnor U2603 (N_2603,N_2562,N_2555);
nor U2604 (N_2604,N_2517,N_2497);
nand U2605 (N_2605,N_2435,N_2505);
or U2606 (N_2606,N_2534,N_2409);
xnor U2607 (N_2607,N_2485,N_2430);
or U2608 (N_2608,N_2402,N_2447);
or U2609 (N_2609,N_2492,N_2501);
or U2610 (N_2610,N_2476,N_2598);
and U2611 (N_2611,N_2493,N_2401);
nand U2612 (N_2612,N_2514,N_2421);
and U2613 (N_2613,N_2454,N_2521);
nand U2614 (N_2614,N_2482,N_2594);
nand U2615 (N_2615,N_2572,N_2439);
nor U2616 (N_2616,N_2446,N_2567);
nor U2617 (N_2617,N_2538,N_2568);
nor U2618 (N_2618,N_2442,N_2532);
xnor U2619 (N_2619,N_2455,N_2563);
or U2620 (N_2620,N_2547,N_2523);
nor U2621 (N_2621,N_2491,N_2431);
nor U2622 (N_2622,N_2434,N_2456);
or U2623 (N_2623,N_2597,N_2500);
nor U2624 (N_2624,N_2524,N_2419);
and U2625 (N_2625,N_2470,N_2490);
xnor U2626 (N_2626,N_2432,N_2483);
nand U2627 (N_2627,N_2513,N_2444);
or U2628 (N_2628,N_2449,N_2460);
xor U2629 (N_2629,N_2400,N_2543);
or U2630 (N_2630,N_2588,N_2411);
nand U2631 (N_2631,N_2551,N_2436);
xor U2632 (N_2632,N_2556,N_2503);
xor U2633 (N_2633,N_2573,N_2403);
nor U2634 (N_2634,N_2465,N_2488);
xnor U2635 (N_2635,N_2528,N_2405);
xor U2636 (N_2636,N_2595,N_2542);
or U2637 (N_2637,N_2437,N_2407);
nand U2638 (N_2638,N_2433,N_2510);
or U2639 (N_2639,N_2489,N_2536);
nand U2640 (N_2640,N_2499,N_2552);
nand U2641 (N_2641,N_2416,N_2496);
xnor U2642 (N_2642,N_2472,N_2565);
or U2643 (N_2643,N_2414,N_2569);
xnor U2644 (N_2644,N_2515,N_2424);
nor U2645 (N_2645,N_2566,N_2423);
nor U2646 (N_2646,N_2559,N_2540);
nor U2647 (N_2647,N_2516,N_2526);
nand U2648 (N_2648,N_2417,N_2557);
nand U2649 (N_2649,N_2531,N_2406);
and U2650 (N_2650,N_2461,N_2554);
xnor U2651 (N_2651,N_2453,N_2466);
and U2652 (N_2652,N_2457,N_2519);
nand U2653 (N_2653,N_2589,N_2428);
or U2654 (N_2654,N_2580,N_2507);
nor U2655 (N_2655,N_2512,N_2404);
and U2656 (N_2656,N_2587,N_2474);
and U2657 (N_2657,N_2475,N_2438);
nand U2658 (N_2658,N_2422,N_2593);
or U2659 (N_2659,N_2509,N_2584);
or U2660 (N_2660,N_2582,N_2506);
or U2661 (N_2661,N_2574,N_2450);
or U2662 (N_2662,N_2412,N_2462);
xnor U2663 (N_2663,N_2458,N_2463);
nand U2664 (N_2664,N_2429,N_2467);
nor U2665 (N_2665,N_2440,N_2494);
nand U2666 (N_2666,N_2544,N_2578);
nand U2667 (N_2667,N_2504,N_2591);
or U2668 (N_2668,N_2498,N_2415);
and U2669 (N_2669,N_2583,N_2520);
and U2670 (N_2670,N_2546,N_2525);
and U2671 (N_2671,N_2571,N_2570);
nor U2672 (N_2672,N_2484,N_2487);
xor U2673 (N_2673,N_2550,N_2558);
or U2674 (N_2674,N_2486,N_2561);
xnor U2675 (N_2675,N_2548,N_2537);
xor U2676 (N_2676,N_2410,N_2579);
or U2677 (N_2677,N_2541,N_2545);
xor U2678 (N_2678,N_2508,N_2479);
xor U2679 (N_2679,N_2511,N_2581);
or U2680 (N_2680,N_2480,N_2452);
and U2681 (N_2681,N_2495,N_2533);
or U2682 (N_2682,N_2473,N_2549);
or U2683 (N_2683,N_2527,N_2530);
xor U2684 (N_2684,N_2408,N_2469);
and U2685 (N_2685,N_2576,N_2535);
nor U2686 (N_2686,N_2420,N_2464);
and U2687 (N_2687,N_2471,N_2459);
xnor U2688 (N_2688,N_2575,N_2468);
or U2689 (N_2689,N_2577,N_2586);
and U2690 (N_2690,N_2585,N_2592);
or U2691 (N_2691,N_2502,N_2445);
nor U2692 (N_2692,N_2518,N_2529);
and U2693 (N_2693,N_2478,N_2539);
and U2694 (N_2694,N_2481,N_2413);
and U2695 (N_2695,N_2477,N_2553);
xnor U2696 (N_2696,N_2564,N_2599);
nand U2697 (N_2697,N_2451,N_2590);
xnor U2698 (N_2698,N_2596,N_2560);
and U2699 (N_2699,N_2522,N_2426);
and U2700 (N_2700,N_2411,N_2575);
or U2701 (N_2701,N_2524,N_2581);
and U2702 (N_2702,N_2400,N_2585);
nand U2703 (N_2703,N_2426,N_2560);
nand U2704 (N_2704,N_2505,N_2594);
nor U2705 (N_2705,N_2579,N_2552);
nor U2706 (N_2706,N_2502,N_2441);
and U2707 (N_2707,N_2515,N_2575);
or U2708 (N_2708,N_2454,N_2408);
xor U2709 (N_2709,N_2587,N_2450);
nand U2710 (N_2710,N_2520,N_2426);
nor U2711 (N_2711,N_2553,N_2578);
and U2712 (N_2712,N_2560,N_2403);
and U2713 (N_2713,N_2510,N_2455);
xnor U2714 (N_2714,N_2539,N_2409);
nor U2715 (N_2715,N_2402,N_2570);
and U2716 (N_2716,N_2412,N_2509);
and U2717 (N_2717,N_2440,N_2414);
nor U2718 (N_2718,N_2517,N_2578);
nor U2719 (N_2719,N_2400,N_2406);
xor U2720 (N_2720,N_2402,N_2424);
nand U2721 (N_2721,N_2488,N_2416);
and U2722 (N_2722,N_2502,N_2411);
nor U2723 (N_2723,N_2534,N_2457);
or U2724 (N_2724,N_2425,N_2492);
nand U2725 (N_2725,N_2532,N_2403);
nand U2726 (N_2726,N_2488,N_2527);
nor U2727 (N_2727,N_2588,N_2447);
or U2728 (N_2728,N_2412,N_2504);
xnor U2729 (N_2729,N_2575,N_2432);
nand U2730 (N_2730,N_2555,N_2553);
or U2731 (N_2731,N_2472,N_2586);
nor U2732 (N_2732,N_2520,N_2478);
and U2733 (N_2733,N_2543,N_2518);
and U2734 (N_2734,N_2481,N_2542);
xor U2735 (N_2735,N_2570,N_2525);
xnor U2736 (N_2736,N_2540,N_2596);
nand U2737 (N_2737,N_2405,N_2450);
nor U2738 (N_2738,N_2598,N_2490);
nor U2739 (N_2739,N_2416,N_2440);
nor U2740 (N_2740,N_2404,N_2449);
and U2741 (N_2741,N_2545,N_2565);
and U2742 (N_2742,N_2477,N_2406);
nor U2743 (N_2743,N_2419,N_2550);
and U2744 (N_2744,N_2494,N_2508);
xnor U2745 (N_2745,N_2472,N_2548);
or U2746 (N_2746,N_2517,N_2507);
and U2747 (N_2747,N_2412,N_2551);
nand U2748 (N_2748,N_2599,N_2511);
or U2749 (N_2749,N_2498,N_2544);
or U2750 (N_2750,N_2578,N_2415);
xor U2751 (N_2751,N_2571,N_2427);
nor U2752 (N_2752,N_2565,N_2597);
nand U2753 (N_2753,N_2547,N_2449);
and U2754 (N_2754,N_2578,N_2424);
or U2755 (N_2755,N_2489,N_2513);
or U2756 (N_2756,N_2554,N_2444);
xnor U2757 (N_2757,N_2463,N_2414);
and U2758 (N_2758,N_2552,N_2465);
and U2759 (N_2759,N_2459,N_2563);
nor U2760 (N_2760,N_2486,N_2436);
nor U2761 (N_2761,N_2433,N_2504);
nand U2762 (N_2762,N_2550,N_2505);
nor U2763 (N_2763,N_2421,N_2593);
and U2764 (N_2764,N_2516,N_2514);
and U2765 (N_2765,N_2528,N_2504);
nand U2766 (N_2766,N_2485,N_2483);
xnor U2767 (N_2767,N_2568,N_2532);
nor U2768 (N_2768,N_2427,N_2573);
nand U2769 (N_2769,N_2409,N_2477);
and U2770 (N_2770,N_2402,N_2583);
and U2771 (N_2771,N_2457,N_2426);
nand U2772 (N_2772,N_2417,N_2486);
and U2773 (N_2773,N_2530,N_2566);
and U2774 (N_2774,N_2571,N_2562);
nor U2775 (N_2775,N_2405,N_2488);
xor U2776 (N_2776,N_2522,N_2542);
nor U2777 (N_2777,N_2550,N_2475);
nor U2778 (N_2778,N_2495,N_2539);
nand U2779 (N_2779,N_2450,N_2539);
nor U2780 (N_2780,N_2519,N_2507);
or U2781 (N_2781,N_2415,N_2481);
xnor U2782 (N_2782,N_2503,N_2409);
nor U2783 (N_2783,N_2569,N_2407);
xnor U2784 (N_2784,N_2506,N_2507);
nor U2785 (N_2785,N_2502,N_2521);
or U2786 (N_2786,N_2504,N_2440);
and U2787 (N_2787,N_2570,N_2462);
or U2788 (N_2788,N_2573,N_2439);
xor U2789 (N_2789,N_2471,N_2440);
and U2790 (N_2790,N_2586,N_2466);
or U2791 (N_2791,N_2571,N_2555);
nand U2792 (N_2792,N_2520,N_2516);
and U2793 (N_2793,N_2457,N_2571);
nand U2794 (N_2794,N_2421,N_2573);
nand U2795 (N_2795,N_2453,N_2406);
and U2796 (N_2796,N_2518,N_2546);
nand U2797 (N_2797,N_2425,N_2592);
and U2798 (N_2798,N_2506,N_2537);
xor U2799 (N_2799,N_2440,N_2463);
nand U2800 (N_2800,N_2712,N_2755);
nor U2801 (N_2801,N_2658,N_2698);
nand U2802 (N_2802,N_2655,N_2685);
and U2803 (N_2803,N_2687,N_2693);
nor U2804 (N_2804,N_2760,N_2785);
or U2805 (N_2805,N_2667,N_2763);
nor U2806 (N_2806,N_2630,N_2627);
or U2807 (N_2807,N_2734,N_2635);
nand U2808 (N_2808,N_2604,N_2794);
nand U2809 (N_2809,N_2740,N_2681);
nand U2810 (N_2810,N_2775,N_2765);
nor U2811 (N_2811,N_2759,N_2735);
nor U2812 (N_2812,N_2676,N_2683);
nor U2813 (N_2813,N_2771,N_2672);
xor U2814 (N_2814,N_2704,N_2787);
and U2815 (N_2815,N_2773,N_2786);
or U2816 (N_2816,N_2719,N_2694);
and U2817 (N_2817,N_2620,N_2644);
xnor U2818 (N_2818,N_2701,N_2690);
nand U2819 (N_2819,N_2741,N_2651);
xor U2820 (N_2820,N_2730,N_2654);
nor U2821 (N_2821,N_2652,N_2772);
nand U2822 (N_2822,N_2709,N_2754);
xnor U2823 (N_2823,N_2789,N_2697);
xor U2824 (N_2824,N_2731,N_2795);
or U2825 (N_2825,N_2799,N_2650);
nand U2826 (N_2826,N_2657,N_2616);
nor U2827 (N_2827,N_2732,N_2792);
xor U2828 (N_2828,N_2796,N_2602);
or U2829 (N_2829,N_2609,N_2737);
or U2830 (N_2830,N_2674,N_2723);
xor U2831 (N_2831,N_2628,N_2728);
nand U2832 (N_2832,N_2626,N_2682);
nor U2833 (N_2833,N_2780,N_2766);
or U2834 (N_2834,N_2727,N_2779);
and U2835 (N_2835,N_2748,N_2758);
and U2836 (N_2836,N_2646,N_2747);
nor U2837 (N_2837,N_2603,N_2661);
and U2838 (N_2838,N_2722,N_2782);
nor U2839 (N_2839,N_2761,N_2633);
nand U2840 (N_2840,N_2739,N_2680);
xnor U2841 (N_2841,N_2714,N_2726);
nor U2842 (N_2842,N_2783,N_2749);
nand U2843 (N_2843,N_2729,N_2798);
nand U2844 (N_2844,N_2797,N_2793);
or U2845 (N_2845,N_2718,N_2753);
nand U2846 (N_2846,N_2611,N_2668);
and U2847 (N_2847,N_2639,N_2671);
xnor U2848 (N_2848,N_2691,N_2623);
xnor U2849 (N_2849,N_2692,N_2664);
or U2850 (N_2850,N_2784,N_2641);
nor U2851 (N_2851,N_2669,N_2660);
or U2852 (N_2852,N_2662,N_2600);
or U2853 (N_2853,N_2770,N_2636);
nand U2854 (N_2854,N_2751,N_2665);
and U2855 (N_2855,N_2643,N_2788);
nor U2856 (N_2856,N_2707,N_2791);
xnor U2857 (N_2857,N_2642,N_2675);
or U2858 (N_2858,N_2713,N_2768);
xor U2859 (N_2859,N_2721,N_2774);
nand U2860 (N_2860,N_2738,N_2743);
and U2861 (N_2861,N_2601,N_2612);
and U2862 (N_2862,N_2618,N_2622);
xnor U2863 (N_2863,N_2645,N_2757);
or U2864 (N_2864,N_2679,N_2608);
and U2865 (N_2865,N_2613,N_2710);
and U2866 (N_2866,N_2678,N_2656);
nand U2867 (N_2867,N_2778,N_2689);
xor U2868 (N_2868,N_2638,N_2720);
xor U2869 (N_2869,N_2663,N_2686);
or U2870 (N_2870,N_2649,N_2724);
xnor U2871 (N_2871,N_2632,N_2708);
xnor U2872 (N_2872,N_2606,N_2653);
and U2873 (N_2873,N_2767,N_2702);
nor U2874 (N_2874,N_2684,N_2631);
and U2875 (N_2875,N_2673,N_2744);
or U2876 (N_2876,N_2688,N_2621);
nor U2877 (N_2877,N_2699,N_2637);
nor U2878 (N_2878,N_2715,N_2717);
and U2879 (N_2879,N_2695,N_2706);
xor U2880 (N_2880,N_2716,N_2610);
nor U2881 (N_2881,N_2607,N_2670);
nand U2882 (N_2882,N_2615,N_2776);
xor U2883 (N_2883,N_2742,N_2733);
or U2884 (N_2884,N_2762,N_2756);
nand U2885 (N_2885,N_2700,N_2705);
nor U2886 (N_2886,N_2617,N_2725);
nor U2887 (N_2887,N_2750,N_2614);
and U2888 (N_2888,N_2711,N_2625);
xnor U2889 (N_2889,N_2769,N_2605);
or U2890 (N_2890,N_2736,N_2696);
or U2891 (N_2891,N_2745,N_2777);
nand U2892 (N_2892,N_2666,N_2677);
or U2893 (N_2893,N_2703,N_2781);
nand U2894 (N_2894,N_2629,N_2752);
xnor U2895 (N_2895,N_2640,N_2647);
nor U2896 (N_2896,N_2648,N_2790);
nor U2897 (N_2897,N_2624,N_2746);
nand U2898 (N_2898,N_2764,N_2619);
nor U2899 (N_2899,N_2659,N_2634);
or U2900 (N_2900,N_2730,N_2616);
nor U2901 (N_2901,N_2726,N_2639);
or U2902 (N_2902,N_2608,N_2661);
or U2903 (N_2903,N_2734,N_2724);
and U2904 (N_2904,N_2757,N_2756);
nand U2905 (N_2905,N_2642,N_2695);
xor U2906 (N_2906,N_2664,N_2616);
nor U2907 (N_2907,N_2620,N_2611);
xor U2908 (N_2908,N_2773,N_2714);
nor U2909 (N_2909,N_2733,N_2600);
nand U2910 (N_2910,N_2601,N_2768);
xor U2911 (N_2911,N_2603,N_2613);
nand U2912 (N_2912,N_2619,N_2771);
and U2913 (N_2913,N_2728,N_2710);
xnor U2914 (N_2914,N_2765,N_2602);
nor U2915 (N_2915,N_2796,N_2679);
and U2916 (N_2916,N_2784,N_2744);
xor U2917 (N_2917,N_2673,N_2697);
or U2918 (N_2918,N_2610,N_2774);
nor U2919 (N_2919,N_2711,N_2607);
nand U2920 (N_2920,N_2738,N_2611);
nor U2921 (N_2921,N_2604,N_2612);
nand U2922 (N_2922,N_2754,N_2674);
and U2923 (N_2923,N_2684,N_2714);
xor U2924 (N_2924,N_2688,N_2722);
or U2925 (N_2925,N_2771,N_2708);
and U2926 (N_2926,N_2723,N_2665);
xor U2927 (N_2927,N_2674,N_2772);
nor U2928 (N_2928,N_2695,N_2626);
xnor U2929 (N_2929,N_2618,N_2703);
or U2930 (N_2930,N_2681,N_2684);
nand U2931 (N_2931,N_2659,N_2708);
nand U2932 (N_2932,N_2668,N_2612);
and U2933 (N_2933,N_2628,N_2770);
and U2934 (N_2934,N_2671,N_2683);
nand U2935 (N_2935,N_2679,N_2699);
or U2936 (N_2936,N_2603,N_2638);
and U2937 (N_2937,N_2619,N_2625);
nor U2938 (N_2938,N_2608,N_2774);
xor U2939 (N_2939,N_2689,N_2694);
nand U2940 (N_2940,N_2727,N_2671);
xnor U2941 (N_2941,N_2676,N_2637);
nand U2942 (N_2942,N_2726,N_2658);
xor U2943 (N_2943,N_2781,N_2754);
xor U2944 (N_2944,N_2668,N_2791);
xnor U2945 (N_2945,N_2696,N_2649);
and U2946 (N_2946,N_2641,N_2706);
xor U2947 (N_2947,N_2633,N_2698);
nor U2948 (N_2948,N_2640,N_2722);
xor U2949 (N_2949,N_2648,N_2764);
nor U2950 (N_2950,N_2693,N_2781);
nand U2951 (N_2951,N_2675,N_2662);
xor U2952 (N_2952,N_2628,N_2659);
or U2953 (N_2953,N_2635,N_2747);
or U2954 (N_2954,N_2723,N_2628);
or U2955 (N_2955,N_2718,N_2729);
xnor U2956 (N_2956,N_2659,N_2700);
nor U2957 (N_2957,N_2712,N_2703);
and U2958 (N_2958,N_2792,N_2755);
and U2959 (N_2959,N_2640,N_2753);
nor U2960 (N_2960,N_2676,N_2793);
nand U2961 (N_2961,N_2799,N_2627);
nor U2962 (N_2962,N_2662,N_2652);
nand U2963 (N_2963,N_2751,N_2780);
or U2964 (N_2964,N_2683,N_2775);
nand U2965 (N_2965,N_2727,N_2651);
or U2966 (N_2966,N_2773,N_2788);
nor U2967 (N_2967,N_2780,N_2659);
nand U2968 (N_2968,N_2720,N_2758);
nand U2969 (N_2969,N_2731,N_2671);
or U2970 (N_2970,N_2635,N_2653);
xor U2971 (N_2971,N_2651,N_2795);
or U2972 (N_2972,N_2680,N_2763);
nand U2973 (N_2973,N_2672,N_2725);
nand U2974 (N_2974,N_2722,N_2603);
xor U2975 (N_2975,N_2623,N_2726);
nand U2976 (N_2976,N_2688,N_2730);
xnor U2977 (N_2977,N_2690,N_2680);
nand U2978 (N_2978,N_2795,N_2688);
nor U2979 (N_2979,N_2691,N_2643);
xnor U2980 (N_2980,N_2648,N_2798);
nor U2981 (N_2981,N_2787,N_2746);
xor U2982 (N_2982,N_2664,N_2603);
nand U2983 (N_2983,N_2692,N_2684);
nand U2984 (N_2984,N_2749,N_2764);
and U2985 (N_2985,N_2644,N_2709);
nor U2986 (N_2986,N_2758,N_2697);
nand U2987 (N_2987,N_2613,N_2784);
nor U2988 (N_2988,N_2646,N_2727);
and U2989 (N_2989,N_2690,N_2788);
nor U2990 (N_2990,N_2781,N_2678);
xnor U2991 (N_2991,N_2629,N_2739);
or U2992 (N_2992,N_2622,N_2781);
nand U2993 (N_2993,N_2638,N_2677);
and U2994 (N_2994,N_2621,N_2632);
and U2995 (N_2995,N_2680,N_2776);
xnor U2996 (N_2996,N_2726,N_2693);
or U2997 (N_2997,N_2669,N_2644);
nand U2998 (N_2998,N_2686,N_2771);
nand U2999 (N_2999,N_2604,N_2610);
xor U3000 (N_3000,N_2863,N_2943);
nor U3001 (N_3001,N_2983,N_2920);
nand U3002 (N_3002,N_2824,N_2929);
xnor U3003 (N_3003,N_2972,N_2960);
xor U3004 (N_3004,N_2978,N_2860);
xnor U3005 (N_3005,N_2956,N_2861);
nor U3006 (N_3006,N_2926,N_2834);
xor U3007 (N_3007,N_2825,N_2936);
nand U3008 (N_3008,N_2876,N_2981);
nor U3009 (N_3009,N_2974,N_2806);
and U3010 (N_3010,N_2965,N_2823);
nand U3011 (N_3011,N_2831,N_2805);
and U3012 (N_3012,N_2951,N_2957);
or U3013 (N_3013,N_2993,N_2845);
or U3014 (N_3014,N_2873,N_2977);
nor U3015 (N_3015,N_2815,N_2940);
and U3016 (N_3016,N_2880,N_2839);
or U3017 (N_3017,N_2950,N_2955);
nand U3018 (N_3018,N_2907,N_2807);
nor U3019 (N_3019,N_2897,N_2992);
xnor U3020 (N_3020,N_2867,N_2984);
and U3021 (N_3021,N_2924,N_2922);
nor U3022 (N_3022,N_2804,N_2828);
xnor U3023 (N_3023,N_2896,N_2833);
xnor U3024 (N_3024,N_2879,N_2872);
and U3025 (N_3025,N_2826,N_2885);
xor U3026 (N_3026,N_2967,N_2988);
nand U3027 (N_3027,N_2973,N_2817);
and U3028 (N_3028,N_2842,N_2865);
nor U3029 (N_3029,N_2813,N_2997);
nand U3030 (N_3030,N_2811,N_2875);
and U3031 (N_3031,N_2836,N_2821);
xor U3032 (N_3032,N_2800,N_2871);
or U3033 (N_3033,N_2862,N_2844);
or U3034 (N_3034,N_2902,N_2878);
nand U3035 (N_3035,N_2818,N_2966);
nand U3036 (N_3036,N_2830,N_2888);
or U3037 (N_3037,N_2855,N_2814);
nor U3038 (N_3038,N_2998,N_2887);
nor U3039 (N_3039,N_2849,N_2891);
xor U3040 (N_3040,N_2954,N_2986);
nor U3041 (N_3041,N_2819,N_2919);
or U3042 (N_3042,N_2802,N_2803);
and U3043 (N_3043,N_2944,N_2914);
nand U3044 (N_3044,N_2937,N_2933);
nor U3045 (N_3045,N_2884,N_2820);
and U3046 (N_3046,N_2829,N_2827);
and U3047 (N_3047,N_2946,N_2971);
or U3048 (N_3048,N_2994,N_2912);
and U3049 (N_3049,N_2964,N_2911);
nand U3050 (N_3050,N_2932,N_2822);
or U3051 (N_3051,N_2941,N_2895);
and U3052 (N_3052,N_2859,N_2846);
xor U3053 (N_3053,N_2906,N_2928);
and U3054 (N_3054,N_2852,N_2898);
and U3055 (N_3055,N_2938,N_2832);
nand U3056 (N_3056,N_2918,N_2935);
xnor U3057 (N_3057,N_2841,N_2857);
nand U3058 (N_3058,N_2969,N_2812);
and U3059 (N_3059,N_2934,N_2910);
and U3060 (N_3060,N_2985,N_2840);
nand U3061 (N_3061,N_2894,N_2908);
xor U3062 (N_3062,N_2980,N_2881);
xnor U3063 (N_3063,N_2877,N_2899);
xor U3064 (N_3064,N_2851,N_2921);
or U3065 (N_3065,N_2853,N_2913);
xor U3066 (N_3066,N_2948,N_2903);
nand U3067 (N_3067,N_2968,N_2975);
nor U3068 (N_3068,N_2837,N_2939);
xor U3069 (N_3069,N_2843,N_2999);
nand U3070 (N_3070,N_2979,N_2945);
or U3071 (N_3071,N_2874,N_2866);
nor U3072 (N_3072,N_2808,N_2916);
xnor U3073 (N_3073,N_2847,N_2848);
or U3074 (N_3074,N_2959,N_2923);
and U3075 (N_3075,N_2892,N_2947);
nor U3076 (N_3076,N_2900,N_2996);
nor U3077 (N_3077,N_2883,N_2890);
nand U3078 (N_3078,N_2886,N_2991);
nand U3079 (N_3079,N_2970,N_2868);
and U3080 (N_3080,N_2893,N_2854);
xnor U3081 (N_3081,N_2809,N_2930);
or U3082 (N_3082,N_2838,N_2901);
and U3083 (N_3083,N_2905,N_2953);
or U3084 (N_3084,N_2961,N_2864);
or U3085 (N_3085,N_2949,N_2835);
xor U3086 (N_3086,N_2889,N_2915);
and U3087 (N_3087,N_2801,N_2858);
xnor U3088 (N_3088,N_2962,N_2925);
nand U3089 (N_3089,N_2982,N_2882);
and U3090 (N_3090,N_2850,N_2870);
or U3091 (N_3091,N_2987,N_2917);
nand U3092 (N_3092,N_2990,N_2931);
nand U3093 (N_3093,N_2904,N_2816);
nor U3094 (N_3094,N_2810,N_2976);
nor U3095 (N_3095,N_2989,N_2958);
xor U3096 (N_3096,N_2963,N_2942);
or U3097 (N_3097,N_2869,N_2856);
xnor U3098 (N_3098,N_2909,N_2927);
nand U3099 (N_3099,N_2952,N_2995);
xnor U3100 (N_3100,N_2875,N_2835);
nand U3101 (N_3101,N_2836,N_2847);
xnor U3102 (N_3102,N_2995,N_2916);
nor U3103 (N_3103,N_2833,N_2870);
nand U3104 (N_3104,N_2908,N_2816);
nor U3105 (N_3105,N_2901,N_2872);
xor U3106 (N_3106,N_2955,N_2878);
nor U3107 (N_3107,N_2973,N_2956);
nand U3108 (N_3108,N_2939,N_2964);
xor U3109 (N_3109,N_2979,N_2856);
or U3110 (N_3110,N_2970,N_2883);
and U3111 (N_3111,N_2886,N_2864);
or U3112 (N_3112,N_2870,N_2943);
and U3113 (N_3113,N_2883,N_2999);
nand U3114 (N_3114,N_2834,N_2886);
or U3115 (N_3115,N_2844,N_2892);
nand U3116 (N_3116,N_2950,N_2927);
nand U3117 (N_3117,N_2955,N_2928);
and U3118 (N_3118,N_2977,N_2895);
and U3119 (N_3119,N_2863,N_2959);
or U3120 (N_3120,N_2904,N_2940);
nor U3121 (N_3121,N_2820,N_2993);
and U3122 (N_3122,N_2885,N_2920);
or U3123 (N_3123,N_2932,N_2878);
xor U3124 (N_3124,N_2838,N_2931);
nand U3125 (N_3125,N_2905,N_2803);
or U3126 (N_3126,N_2953,N_2821);
xor U3127 (N_3127,N_2827,N_2930);
xor U3128 (N_3128,N_2954,N_2845);
nor U3129 (N_3129,N_2949,N_2834);
xor U3130 (N_3130,N_2845,N_2802);
xnor U3131 (N_3131,N_2940,N_2935);
nand U3132 (N_3132,N_2817,N_2940);
xnor U3133 (N_3133,N_2979,N_2968);
nor U3134 (N_3134,N_2845,N_2880);
xor U3135 (N_3135,N_2892,N_2971);
or U3136 (N_3136,N_2828,N_2922);
nor U3137 (N_3137,N_2881,N_2907);
or U3138 (N_3138,N_2949,N_2934);
nor U3139 (N_3139,N_2889,N_2992);
nand U3140 (N_3140,N_2962,N_2845);
nor U3141 (N_3141,N_2864,N_2958);
and U3142 (N_3142,N_2968,N_2851);
and U3143 (N_3143,N_2961,N_2997);
xor U3144 (N_3144,N_2817,N_2831);
nand U3145 (N_3145,N_2941,N_2835);
xor U3146 (N_3146,N_2872,N_2800);
nor U3147 (N_3147,N_2875,N_2845);
and U3148 (N_3148,N_2819,N_2831);
and U3149 (N_3149,N_2860,N_2875);
nor U3150 (N_3150,N_2832,N_2957);
nor U3151 (N_3151,N_2946,N_2976);
nand U3152 (N_3152,N_2963,N_2883);
nor U3153 (N_3153,N_2964,N_2999);
nor U3154 (N_3154,N_2999,N_2935);
and U3155 (N_3155,N_2922,N_2869);
and U3156 (N_3156,N_2856,N_2825);
or U3157 (N_3157,N_2820,N_2937);
nor U3158 (N_3158,N_2913,N_2921);
nor U3159 (N_3159,N_2908,N_2995);
xnor U3160 (N_3160,N_2894,N_2948);
and U3161 (N_3161,N_2853,N_2854);
or U3162 (N_3162,N_2926,N_2917);
or U3163 (N_3163,N_2825,N_2956);
nand U3164 (N_3164,N_2907,N_2836);
nand U3165 (N_3165,N_2961,N_2908);
nand U3166 (N_3166,N_2867,N_2893);
nor U3167 (N_3167,N_2960,N_2841);
or U3168 (N_3168,N_2939,N_2948);
xor U3169 (N_3169,N_2992,N_2804);
and U3170 (N_3170,N_2896,N_2898);
xor U3171 (N_3171,N_2980,N_2943);
xnor U3172 (N_3172,N_2984,N_2879);
or U3173 (N_3173,N_2964,N_2899);
or U3174 (N_3174,N_2879,N_2830);
or U3175 (N_3175,N_2915,N_2922);
nand U3176 (N_3176,N_2976,N_2895);
and U3177 (N_3177,N_2914,N_2929);
nand U3178 (N_3178,N_2959,N_2894);
nand U3179 (N_3179,N_2859,N_2917);
nor U3180 (N_3180,N_2843,N_2819);
xnor U3181 (N_3181,N_2828,N_2971);
or U3182 (N_3182,N_2988,N_2802);
and U3183 (N_3183,N_2812,N_2897);
or U3184 (N_3184,N_2818,N_2905);
or U3185 (N_3185,N_2915,N_2848);
or U3186 (N_3186,N_2983,N_2823);
or U3187 (N_3187,N_2866,N_2823);
or U3188 (N_3188,N_2823,N_2847);
nor U3189 (N_3189,N_2880,N_2965);
and U3190 (N_3190,N_2805,N_2807);
nor U3191 (N_3191,N_2887,N_2839);
nor U3192 (N_3192,N_2839,N_2994);
nor U3193 (N_3193,N_2836,N_2859);
xnor U3194 (N_3194,N_2990,N_2858);
xnor U3195 (N_3195,N_2807,N_2900);
nand U3196 (N_3196,N_2990,N_2876);
nand U3197 (N_3197,N_2856,N_2852);
or U3198 (N_3198,N_2803,N_2834);
or U3199 (N_3199,N_2886,N_2818);
nand U3200 (N_3200,N_3198,N_3043);
nand U3201 (N_3201,N_3091,N_3053);
nor U3202 (N_3202,N_3082,N_3071);
or U3203 (N_3203,N_3182,N_3146);
nand U3204 (N_3204,N_3153,N_3080);
or U3205 (N_3205,N_3065,N_3160);
nand U3206 (N_3206,N_3169,N_3030);
nand U3207 (N_3207,N_3130,N_3180);
nand U3208 (N_3208,N_3084,N_3179);
nand U3209 (N_3209,N_3076,N_3039);
xor U3210 (N_3210,N_3019,N_3097);
nor U3211 (N_3211,N_3199,N_3102);
nor U3212 (N_3212,N_3020,N_3067);
nand U3213 (N_3213,N_3070,N_3123);
nor U3214 (N_3214,N_3178,N_3118);
xnor U3215 (N_3215,N_3167,N_3168);
and U3216 (N_3216,N_3190,N_3108);
nand U3217 (N_3217,N_3023,N_3129);
and U3218 (N_3218,N_3087,N_3104);
nand U3219 (N_3219,N_3176,N_3173);
and U3220 (N_3220,N_3105,N_3092);
and U3221 (N_3221,N_3121,N_3128);
xnor U3222 (N_3222,N_3059,N_3162);
xnor U3223 (N_3223,N_3073,N_3027);
and U3224 (N_3224,N_3103,N_3047);
or U3225 (N_3225,N_3048,N_3191);
nor U3226 (N_3226,N_3037,N_3101);
nor U3227 (N_3227,N_3189,N_3106);
and U3228 (N_3228,N_3116,N_3196);
and U3229 (N_3229,N_3007,N_3188);
and U3230 (N_3230,N_3094,N_3136);
or U3231 (N_3231,N_3197,N_3157);
xnor U3232 (N_3232,N_3117,N_3138);
nand U3233 (N_3233,N_3124,N_3181);
or U3234 (N_3234,N_3046,N_3099);
or U3235 (N_3235,N_3109,N_3171);
xor U3236 (N_3236,N_3166,N_3015);
nor U3237 (N_3237,N_3143,N_3148);
xnor U3238 (N_3238,N_3145,N_3078);
nor U3239 (N_3239,N_3011,N_3120);
and U3240 (N_3240,N_3139,N_3144);
and U3241 (N_3241,N_3086,N_3003);
nor U3242 (N_3242,N_3068,N_3032);
nor U3243 (N_3243,N_3098,N_3049);
or U3244 (N_3244,N_3125,N_3014);
xor U3245 (N_3245,N_3083,N_3149);
nand U3246 (N_3246,N_3147,N_3156);
nand U3247 (N_3247,N_3055,N_3111);
and U3248 (N_3248,N_3085,N_3062);
or U3249 (N_3249,N_3093,N_3172);
xor U3250 (N_3250,N_3018,N_3135);
and U3251 (N_3251,N_3081,N_3077);
nor U3252 (N_3252,N_3122,N_3035);
and U3253 (N_3253,N_3017,N_3194);
or U3254 (N_3254,N_3119,N_3158);
nand U3255 (N_3255,N_3100,N_3064);
nor U3256 (N_3256,N_3132,N_3134);
nand U3257 (N_3257,N_3045,N_3186);
and U3258 (N_3258,N_3074,N_3090);
nand U3259 (N_3259,N_3170,N_3107);
nand U3260 (N_3260,N_3008,N_3110);
nor U3261 (N_3261,N_3133,N_3164);
and U3262 (N_3262,N_3072,N_3060);
or U3263 (N_3263,N_3174,N_3175);
xor U3264 (N_3264,N_3161,N_3012);
and U3265 (N_3265,N_3025,N_3056);
xnor U3266 (N_3266,N_3184,N_3040);
xor U3267 (N_3267,N_3131,N_3154);
nor U3268 (N_3268,N_3038,N_3009);
and U3269 (N_3269,N_3001,N_3137);
xor U3270 (N_3270,N_3028,N_3002);
and U3271 (N_3271,N_3024,N_3041);
xor U3272 (N_3272,N_3061,N_3058);
nand U3273 (N_3273,N_3155,N_3026);
or U3274 (N_3274,N_3033,N_3088);
xor U3275 (N_3275,N_3000,N_3114);
and U3276 (N_3276,N_3079,N_3016);
and U3277 (N_3277,N_3021,N_3152);
nand U3278 (N_3278,N_3031,N_3057);
or U3279 (N_3279,N_3115,N_3034);
nand U3280 (N_3280,N_3177,N_3140);
or U3281 (N_3281,N_3192,N_3163);
nand U3282 (N_3282,N_3142,N_3066);
and U3283 (N_3283,N_3095,N_3042);
xor U3284 (N_3284,N_3063,N_3150);
nand U3285 (N_3285,N_3004,N_3052);
and U3286 (N_3286,N_3195,N_3183);
or U3287 (N_3287,N_3022,N_3193);
or U3288 (N_3288,N_3044,N_3029);
xor U3289 (N_3289,N_3051,N_3089);
nand U3290 (N_3290,N_3010,N_3187);
and U3291 (N_3291,N_3113,N_3127);
and U3292 (N_3292,N_3112,N_3126);
or U3293 (N_3293,N_3075,N_3096);
nor U3294 (N_3294,N_3005,N_3185);
nor U3295 (N_3295,N_3141,N_3036);
and U3296 (N_3296,N_3069,N_3050);
and U3297 (N_3297,N_3054,N_3006);
and U3298 (N_3298,N_3013,N_3159);
and U3299 (N_3299,N_3151,N_3165);
nor U3300 (N_3300,N_3098,N_3138);
nand U3301 (N_3301,N_3139,N_3172);
nand U3302 (N_3302,N_3062,N_3191);
or U3303 (N_3303,N_3026,N_3187);
nor U3304 (N_3304,N_3024,N_3153);
xor U3305 (N_3305,N_3117,N_3058);
xor U3306 (N_3306,N_3173,N_3042);
and U3307 (N_3307,N_3190,N_3067);
xor U3308 (N_3308,N_3188,N_3062);
and U3309 (N_3309,N_3019,N_3152);
and U3310 (N_3310,N_3162,N_3122);
or U3311 (N_3311,N_3191,N_3169);
nand U3312 (N_3312,N_3069,N_3141);
nand U3313 (N_3313,N_3117,N_3047);
nand U3314 (N_3314,N_3003,N_3095);
nand U3315 (N_3315,N_3036,N_3180);
xnor U3316 (N_3316,N_3164,N_3034);
nor U3317 (N_3317,N_3069,N_3042);
xnor U3318 (N_3318,N_3115,N_3159);
nor U3319 (N_3319,N_3161,N_3174);
nor U3320 (N_3320,N_3099,N_3188);
or U3321 (N_3321,N_3073,N_3045);
and U3322 (N_3322,N_3171,N_3060);
xnor U3323 (N_3323,N_3092,N_3094);
nor U3324 (N_3324,N_3095,N_3177);
or U3325 (N_3325,N_3004,N_3103);
xor U3326 (N_3326,N_3195,N_3134);
xor U3327 (N_3327,N_3174,N_3143);
or U3328 (N_3328,N_3045,N_3148);
or U3329 (N_3329,N_3180,N_3083);
and U3330 (N_3330,N_3001,N_3090);
and U3331 (N_3331,N_3161,N_3083);
and U3332 (N_3332,N_3071,N_3016);
nand U3333 (N_3333,N_3054,N_3002);
xnor U3334 (N_3334,N_3069,N_3033);
nor U3335 (N_3335,N_3097,N_3149);
and U3336 (N_3336,N_3032,N_3095);
xor U3337 (N_3337,N_3181,N_3054);
xnor U3338 (N_3338,N_3018,N_3180);
nand U3339 (N_3339,N_3093,N_3185);
and U3340 (N_3340,N_3046,N_3161);
and U3341 (N_3341,N_3115,N_3055);
or U3342 (N_3342,N_3089,N_3128);
xor U3343 (N_3343,N_3144,N_3149);
nand U3344 (N_3344,N_3056,N_3034);
nand U3345 (N_3345,N_3152,N_3087);
or U3346 (N_3346,N_3013,N_3167);
xor U3347 (N_3347,N_3129,N_3108);
and U3348 (N_3348,N_3165,N_3128);
xor U3349 (N_3349,N_3036,N_3116);
nor U3350 (N_3350,N_3130,N_3179);
nand U3351 (N_3351,N_3061,N_3016);
nand U3352 (N_3352,N_3074,N_3039);
or U3353 (N_3353,N_3004,N_3130);
or U3354 (N_3354,N_3170,N_3149);
and U3355 (N_3355,N_3077,N_3030);
nor U3356 (N_3356,N_3028,N_3181);
or U3357 (N_3357,N_3140,N_3165);
or U3358 (N_3358,N_3129,N_3126);
nor U3359 (N_3359,N_3004,N_3015);
nor U3360 (N_3360,N_3185,N_3030);
xnor U3361 (N_3361,N_3121,N_3167);
xor U3362 (N_3362,N_3114,N_3022);
or U3363 (N_3363,N_3173,N_3061);
xor U3364 (N_3364,N_3045,N_3007);
or U3365 (N_3365,N_3039,N_3047);
nor U3366 (N_3366,N_3116,N_3176);
nor U3367 (N_3367,N_3111,N_3057);
and U3368 (N_3368,N_3002,N_3125);
xnor U3369 (N_3369,N_3168,N_3032);
xor U3370 (N_3370,N_3060,N_3001);
nand U3371 (N_3371,N_3114,N_3152);
nor U3372 (N_3372,N_3074,N_3080);
nor U3373 (N_3373,N_3047,N_3138);
xnor U3374 (N_3374,N_3000,N_3155);
nor U3375 (N_3375,N_3080,N_3169);
nand U3376 (N_3376,N_3097,N_3034);
and U3377 (N_3377,N_3156,N_3178);
nand U3378 (N_3378,N_3105,N_3067);
nand U3379 (N_3379,N_3159,N_3005);
xor U3380 (N_3380,N_3081,N_3147);
xor U3381 (N_3381,N_3157,N_3076);
nor U3382 (N_3382,N_3115,N_3099);
nor U3383 (N_3383,N_3108,N_3182);
nand U3384 (N_3384,N_3160,N_3128);
nor U3385 (N_3385,N_3033,N_3012);
xor U3386 (N_3386,N_3169,N_3099);
nand U3387 (N_3387,N_3059,N_3139);
and U3388 (N_3388,N_3038,N_3010);
nand U3389 (N_3389,N_3068,N_3132);
and U3390 (N_3390,N_3095,N_3094);
nor U3391 (N_3391,N_3129,N_3027);
or U3392 (N_3392,N_3012,N_3019);
and U3393 (N_3393,N_3142,N_3121);
xnor U3394 (N_3394,N_3062,N_3081);
xnor U3395 (N_3395,N_3071,N_3072);
nand U3396 (N_3396,N_3190,N_3193);
nand U3397 (N_3397,N_3067,N_3068);
or U3398 (N_3398,N_3080,N_3000);
nand U3399 (N_3399,N_3020,N_3108);
and U3400 (N_3400,N_3236,N_3241);
nor U3401 (N_3401,N_3279,N_3367);
and U3402 (N_3402,N_3266,N_3334);
nor U3403 (N_3403,N_3206,N_3210);
and U3404 (N_3404,N_3298,N_3360);
and U3405 (N_3405,N_3253,N_3313);
and U3406 (N_3406,N_3387,N_3354);
nor U3407 (N_3407,N_3342,N_3363);
nor U3408 (N_3408,N_3211,N_3378);
nor U3409 (N_3409,N_3300,N_3208);
xor U3410 (N_3410,N_3307,N_3349);
nand U3411 (N_3411,N_3333,N_3290);
and U3412 (N_3412,N_3393,N_3287);
xor U3413 (N_3413,N_3324,N_3277);
xor U3414 (N_3414,N_3250,N_3251);
or U3415 (N_3415,N_3375,N_3291);
xor U3416 (N_3416,N_3325,N_3285);
xnor U3417 (N_3417,N_3351,N_3205);
xnor U3418 (N_3418,N_3339,N_3226);
or U3419 (N_3419,N_3332,N_3284);
and U3420 (N_3420,N_3366,N_3269);
xor U3421 (N_3421,N_3383,N_3293);
xnor U3422 (N_3422,N_3306,N_3305);
xnor U3423 (N_3423,N_3243,N_3316);
and U3424 (N_3424,N_3303,N_3249);
xor U3425 (N_3425,N_3213,N_3372);
nor U3426 (N_3426,N_3386,N_3323);
nand U3427 (N_3427,N_3331,N_3273);
or U3428 (N_3428,N_3352,N_3374);
nor U3429 (N_3429,N_3228,N_3280);
xnor U3430 (N_3430,N_3376,N_3289);
or U3431 (N_3431,N_3286,N_3330);
and U3432 (N_3432,N_3319,N_3265);
nand U3433 (N_3433,N_3314,N_3288);
and U3434 (N_3434,N_3384,N_3338);
or U3435 (N_3435,N_3381,N_3394);
and U3436 (N_3436,N_3294,N_3309);
nand U3437 (N_3437,N_3204,N_3245);
nand U3438 (N_3438,N_3242,N_3297);
nor U3439 (N_3439,N_3234,N_3377);
nor U3440 (N_3440,N_3399,N_3256);
nand U3441 (N_3441,N_3322,N_3304);
or U3442 (N_3442,N_3357,N_3396);
xor U3443 (N_3443,N_3281,N_3203);
and U3444 (N_3444,N_3356,N_3235);
nand U3445 (N_3445,N_3246,N_3276);
nor U3446 (N_3446,N_3373,N_3260);
xnor U3447 (N_3447,N_3364,N_3327);
xor U3448 (N_3448,N_3207,N_3318);
nor U3449 (N_3449,N_3222,N_3248);
and U3450 (N_3450,N_3218,N_3344);
nor U3451 (N_3451,N_3310,N_3238);
nand U3452 (N_3452,N_3335,N_3302);
xor U3453 (N_3453,N_3379,N_3247);
xor U3454 (N_3454,N_3295,N_3398);
nor U3455 (N_3455,N_3296,N_3370);
nor U3456 (N_3456,N_3326,N_3261);
or U3457 (N_3457,N_3255,N_3231);
xnor U3458 (N_3458,N_3240,N_3224);
nand U3459 (N_3459,N_3259,N_3233);
and U3460 (N_3460,N_3275,N_3216);
xor U3461 (N_3461,N_3321,N_3353);
xnor U3462 (N_3462,N_3262,N_3345);
nand U3463 (N_3463,N_3312,N_3348);
or U3464 (N_3464,N_3346,N_3272);
xnor U3465 (N_3465,N_3257,N_3308);
and U3466 (N_3466,N_3355,N_3225);
nand U3467 (N_3467,N_3268,N_3221);
xor U3468 (N_3468,N_3336,N_3392);
nor U3469 (N_3469,N_3278,N_3315);
nor U3470 (N_3470,N_3229,N_3350);
nor U3471 (N_3471,N_3270,N_3209);
or U3472 (N_3472,N_3282,N_3232);
nor U3473 (N_3473,N_3397,N_3359);
nand U3474 (N_3474,N_3317,N_3337);
xor U3475 (N_3475,N_3395,N_3219);
and U3476 (N_3476,N_3217,N_3202);
nor U3477 (N_3477,N_3388,N_3299);
xnor U3478 (N_3478,N_3200,N_3369);
xnor U3479 (N_3479,N_3254,N_3358);
or U3480 (N_3480,N_3311,N_3227);
nand U3481 (N_3481,N_3328,N_3362);
nand U3482 (N_3482,N_3292,N_3252);
xnor U3483 (N_3483,N_3271,N_3391);
or U3484 (N_3484,N_3215,N_3274);
or U3485 (N_3485,N_3343,N_3365);
or U3486 (N_3486,N_3220,N_3329);
and U3487 (N_3487,N_3214,N_3389);
nand U3488 (N_3488,N_3267,N_3201);
xor U3489 (N_3489,N_3341,N_3283);
nand U3490 (N_3490,N_3347,N_3239);
nor U3491 (N_3491,N_3237,N_3244);
nor U3492 (N_3492,N_3258,N_3301);
or U3493 (N_3493,N_3385,N_3223);
xnor U3494 (N_3494,N_3212,N_3263);
xnor U3495 (N_3495,N_3340,N_3320);
or U3496 (N_3496,N_3371,N_3380);
or U3497 (N_3497,N_3390,N_3368);
nor U3498 (N_3498,N_3264,N_3382);
nand U3499 (N_3499,N_3230,N_3361);
xor U3500 (N_3500,N_3264,N_3337);
and U3501 (N_3501,N_3296,N_3326);
xor U3502 (N_3502,N_3273,N_3292);
and U3503 (N_3503,N_3308,N_3368);
nand U3504 (N_3504,N_3351,N_3299);
nor U3505 (N_3505,N_3268,N_3232);
or U3506 (N_3506,N_3228,N_3238);
or U3507 (N_3507,N_3342,N_3231);
and U3508 (N_3508,N_3304,N_3372);
xnor U3509 (N_3509,N_3320,N_3353);
nand U3510 (N_3510,N_3343,N_3296);
xnor U3511 (N_3511,N_3325,N_3367);
xor U3512 (N_3512,N_3211,N_3352);
nand U3513 (N_3513,N_3392,N_3227);
xnor U3514 (N_3514,N_3318,N_3295);
xor U3515 (N_3515,N_3308,N_3216);
xor U3516 (N_3516,N_3305,N_3386);
and U3517 (N_3517,N_3224,N_3245);
nor U3518 (N_3518,N_3222,N_3219);
nor U3519 (N_3519,N_3367,N_3370);
nor U3520 (N_3520,N_3240,N_3290);
xor U3521 (N_3521,N_3299,N_3236);
or U3522 (N_3522,N_3309,N_3241);
or U3523 (N_3523,N_3254,N_3269);
nand U3524 (N_3524,N_3331,N_3238);
xnor U3525 (N_3525,N_3234,N_3208);
xnor U3526 (N_3526,N_3210,N_3289);
and U3527 (N_3527,N_3356,N_3328);
xnor U3528 (N_3528,N_3397,N_3330);
nand U3529 (N_3529,N_3347,N_3304);
and U3530 (N_3530,N_3254,N_3247);
nand U3531 (N_3531,N_3218,N_3214);
and U3532 (N_3532,N_3322,N_3309);
nor U3533 (N_3533,N_3389,N_3348);
xor U3534 (N_3534,N_3317,N_3282);
or U3535 (N_3535,N_3207,N_3282);
xor U3536 (N_3536,N_3356,N_3345);
nor U3537 (N_3537,N_3314,N_3371);
or U3538 (N_3538,N_3374,N_3225);
xnor U3539 (N_3539,N_3396,N_3300);
nand U3540 (N_3540,N_3251,N_3327);
or U3541 (N_3541,N_3396,N_3327);
nand U3542 (N_3542,N_3319,N_3325);
xor U3543 (N_3543,N_3232,N_3315);
and U3544 (N_3544,N_3283,N_3347);
nand U3545 (N_3545,N_3215,N_3306);
nor U3546 (N_3546,N_3343,N_3398);
and U3547 (N_3547,N_3342,N_3386);
xor U3548 (N_3548,N_3225,N_3399);
or U3549 (N_3549,N_3304,N_3326);
or U3550 (N_3550,N_3366,N_3331);
and U3551 (N_3551,N_3246,N_3215);
nor U3552 (N_3552,N_3283,N_3356);
xnor U3553 (N_3553,N_3296,N_3257);
nor U3554 (N_3554,N_3359,N_3315);
nor U3555 (N_3555,N_3220,N_3322);
nand U3556 (N_3556,N_3254,N_3282);
and U3557 (N_3557,N_3249,N_3349);
and U3558 (N_3558,N_3261,N_3252);
or U3559 (N_3559,N_3399,N_3259);
or U3560 (N_3560,N_3386,N_3375);
and U3561 (N_3561,N_3202,N_3201);
nor U3562 (N_3562,N_3379,N_3296);
or U3563 (N_3563,N_3313,N_3292);
and U3564 (N_3564,N_3242,N_3263);
or U3565 (N_3565,N_3264,N_3345);
and U3566 (N_3566,N_3354,N_3215);
or U3567 (N_3567,N_3361,N_3318);
nand U3568 (N_3568,N_3299,N_3248);
nand U3569 (N_3569,N_3229,N_3251);
nand U3570 (N_3570,N_3316,N_3294);
and U3571 (N_3571,N_3208,N_3272);
or U3572 (N_3572,N_3232,N_3250);
or U3573 (N_3573,N_3391,N_3353);
xnor U3574 (N_3574,N_3384,N_3276);
and U3575 (N_3575,N_3237,N_3398);
nor U3576 (N_3576,N_3264,N_3371);
and U3577 (N_3577,N_3240,N_3392);
xnor U3578 (N_3578,N_3354,N_3288);
nand U3579 (N_3579,N_3335,N_3215);
or U3580 (N_3580,N_3330,N_3253);
nand U3581 (N_3581,N_3281,N_3272);
or U3582 (N_3582,N_3310,N_3247);
xnor U3583 (N_3583,N_3334,N_3253);
and U3584 (N_3584,N_3202,N_3313);
or U3585 (N_3585,N_3382,N_3365);
nand U3586 (N_3586,N_3284,N_3262);
or U3587 (N_3587,N_3352,N_3236);
and U3588 (N_3588,N_3320,N_3397);
or U3589 (N_3589,N_3308,N_3392);
nor U3590 (N_3590,N_3292,N_3296);
nor U3591 (N_3591,N_3292,N_3250);
nand U3592 (N_3592,N_3216,N_3392);
nand U3593 (N_3593,N_3344,N_3396);
or U3594 (N_3594,N_3287,N_3326);
nor U3595 (N_3595,N_3247,N_3381);
nor U3596 (N_3596,N_3202,N_3225);
nand U3597 (N_3597,N_3243,N_3278);
nor U3598 (N_3598,N_3307,N_3340);
nor U3599 (N_3599,N_3325,N_3334);
nor U3600 (N_3600,N_3462,N_3589);
and U3601 (N_3601,N_3550,N_3562);
or U3602 (N_3602,N_3539,N_3416);
xor U3603 (N_3603,N_3472,N_3590);
xor U3604 (N_3604,N_3512,N_3584);
nor U3605 (N_3605,N_3548,N_3460);
nand U3606 (N_3606,N_3498,N_3510);
nand U3607 (N_3607,N_3575,N_3466);
nand U3608 (N_3608,N_3522,N_3563);
and U3609 (N_3609,N_3429,N_3424);
nor U3610 (N_3610,N_3506,N_3482);
nand U3611 (N_3611,N_3493,N_3565);
nand U3612 (N_3612,N_3552,N_3536);
or U3613 (N_3613,N_3587,N_3530);
or U3614 (N_3614,N_3595,N_3568);
nor U3615 (N_3615,N_3458,N_3592);
nor U3616 (N_3616,N_3526,N_3495);
xnor U3617 (N_3617,N_3447,N_3453);
and U3618 (N_3618,N_3467,N_3491);
nor U3619 (N_3619,N_3564,N_3596);
nor U3620 (N_3620,N_3555,N_3463);
and U3621 (N_3621,N_3483,N_3407);
nor U3622 (N_3622,N_3557,N_3514);
or U3623 (N_3623,N_3410,N_3579);
nor U3624 (N_3624,N_3473,N_3593);
nor U3625 (N_3625,N_3487,N_3569);
nor U3626 (N_3626,N_3537,N_3481);
xor U3627 (N_3627,N_3438,N_3505);
nor U3628 (N_3628,N_3439,N_3449);
nand U3629 (N_3629,N_3413,N_3553);
and U3630 (N_3630,N_3582,N_3515);
and U3631 (N_3631,N_3419,N_3507);
and U3632 (N_3632,N_3422,N_3556);
xor U3633 (N_3633,N_3542,N_3432);
xor U3634 (N_3634,N_3508,N_3509);
or U3635 (N_3635,N_3517,N_3516);
or U3636 (N_3636,N_3459,N_3519);
xnor U3637 (N_3637,N_3561,N_3435);
nor U3638 (N_3638,N_3478,N_3402);
or U3639 (N_3639,N_3475,N_3477);
or U3640 (N_3640,N_3408,N_3543);
or U3641 (N_3641,N_3479,N_3431);
and U3642 (N_3642,N_3457,N_3406);
xor U3643 (N_3643,N_3474,N_3436);
or U3644 (N_3644,N_3502,N_3559);
and U3645 (N_3645,N_3454,N_3573);
and U3646 (N_3646,N_3403,N_3594);
and U3647 (N_3647,N_3588,N_3488);
and U3648 (N_3648,N_3523,N_3534);
or U3649 (N_3649,N_3578,N_3581);
or U3650 (N_3650,N_3411,N_3577);
nand U3651 (N_3651,N_3426,N_3518);
or U3652 (N_3652,N_3598,N_3531);
nor U3653 (N_3653,N_3574,N_3428);
and U3654 (N_3654,N_3485,N_3430);
xor U3655 (N_3655,N_3451,N_3476);
xor U3656 (N_3656,N_3469,N_3455);
or U3657 (N_3657,N_3546,N_3504);
nand U3658 (N_3658,N_3484,N_3586);
nand U3659 (N_3659,N_3520,N_3480);
nand U3660 (N_3660,N_3401,N_3452);
nand U3661 (N_3661,N_3521,N_3461);
nand U3662 (N_3662,N_3541,N_3583);
and U3663 (N_3663,N_3551,N_3427);
nor U3664 (N_3664,N_3404,N_3423);
nand U3665 (N_3665,N_3425,N_3471);
or U3666 (N_3666,N_3448,N_3549);
xor U3667 (N_3667,N_3492,N_3576);
xnor U3668 (N_3668,N_3489,N_3566);
and U3669 (N_3669,N_3544,N_3490);
nand U3670 (N_3670,N_3417,N_3567);
nor U3671 (N_3671,N_3547,N_3456);
nor U3672 (N_3672,N_3444,N_3599);
nand U3673 (N_3673,N_3597,N_3414);
and U3674 (N_3674,N_3524,N_3533);
and U3675 (N_3675,N_3440,N_3418);
and U3676 (N_3676,N_3532,N_3421);
xor U3677 (N_3677,N_3442,N_3571);
nor U3678 (N_3678,N_3409,N_3420);
nand U3679 (N_3679,N_3585,N_3497);
xnor U3680 (N_3680,N_3529,N_3415);
nand U3681 (N_3681,N_3545,N_3496);
nand U3682 (N_3682,N_3412,N_3446);
nand U3683 (N_3683,N_3572,N_3525);
nor U3684 (N_3684,N_3527,N_3434);
and U3685 (N_3685,N_3528,N_3405);
or U3686 (N_3686,N_3511,N_3501);
or U3687 (N_3687,N_3450,N_3464);
nor U3688 (N_3688,N_3486,N_3494);
xnor U3689 (N_3689,N_3570,N_3580);
nor U3690 (N_3690,N_3441,N_3554);
nor U3691 (N_3691,N_3470,N_3465);
xor U3692 (N_3692,N_3400,N_3503);
or U3693 (N_3693,N_3540,N_3538);
nor U3694 (N_3694,N_3499,N_3443);
nor U3695 (N_3695,N_3535,N_3500);
nor U3696 (N_3696,N_3560,N_3468);
or U3697 (N_3697,N_3591,N_3433);
xor U3698 (N_3698,N_3558,N_3437);
xor U3699 (N_3699,N_3513,N_3445);
nand U3700 (N_3700,N_3431,N_3515);
xnor U3701 (N_3701,N_3586,N_3590);
nand U3702 (N_3702,N_3562,N_3469);
or U3703 (N_3703,N_3416,N_3514);
xor U3704 (N_3704,N_3479,N_3550);
nand U3705 (N_3705,N_3403,N_3496);
xor U3706 (N_3706,N_3459,N_3523);
nand U3707 (N_3707,N_3507,N_3574);
nand U3708 (N_3708,N_3546,N_3515);
and U3709 (N_3709,N_3453,N_3498);
or U3710 (N_3710,N_3572,N_3529);
nand U3711 (N_3711,N_3587,N_3430);
xor U3712 (N_3712,N_3482,N_3474);
nor U3713 (N_3713,N_3487,N_3456);
nand U3714 (N_3714,N_3460,N_3594);
xor U3715 (N_3715,N_3556,N_3494);
or U3716 (N_3716,N_3494,N_3411);
xnor U3717 (N_3717,N_3532,N_3458);
nor U3718 (N_3718,N_3587,N_3598);
xnor U3719 (N_3719,N_3518,N_3457);
nand U3720 (N_3720,N_3411,N_3464);
nand U3721 (N_3721,N_3408,N_3531);
nor U3722 (N_3722,N_3433,N_3567);
or U3723 (N_3723,N_3547,N_3580);
nor U3724 (N_3724,N_3426,N_3507);
or U3725 (N_3725,N_3448,N_3414);
nand U3726 (N_3726,N_3546,N_3507);
nor U3727 (N_3727,N_3444,N_3512);
xor U3728 (N_3728,N_3561,N_3422);
or U3729 (N_3729,N_3587,N_3476);
nor U3730 (N_3730,N_3590,N_3435);
and U3731 (N_3731,N_3481,N_3589);
or U3732 (N_3732,N_3576,N_3586);
nor U3733 (N_3733,N_3536,N_3523);
nand U3734 (N_3734,N_3485,N_3537);
or U3735 (N_3735,N_3471,N_3463);
and U3736 (N_3736,N_3486,N_3400);
and U3737 (N_3737,N_3515,N_3592);
nor U3738 (N_3738,N_3505,N_3568);
and U3739 (N_3739,N_3546,N_3526);
and U3740 (N_3740,N_3554,N_3483);
xnor U3741 (N_3741,N_3523,N_3589);
and U3742 (N_3742,N_3597,N_3503);
nand U3743 (N_3743,N_3400,N_3587);
or U3744 (N_3744,N_3537,N_3489);
nor U3745 (N_3745,N_3476,N_3456);
nand U3746 (N_3746,N_3550,N_3410);
or U3747 (N_3747,N_3582,N_3406);
and U3748 (N_3748,N_3517,N_3508);
and U3749 (N_3749,N_3568,N_3574);
xor U3750 (N_3750,N_3507,N_3482);
or U3751 (N_3751,N_3488,N_3403);
or U3752 (N_3752,N_3504,N_3552);
nor U3753 (N_3753,N_3502,N_3441);
or U3754 (N_3754,N_3465,N_3498);
or U3755 (N_3755,N_3478,N_3592);
xnor U3756 (N_3756,N_3406,N_3586);
and U3757 (N_3757,N_3447,N_3528);
and U3758 (N_3758,N_3427,N_3494);
xor U3759 (N_3759,N_3540,N_3443);
nand U3760 (N_3760,N_3533,N_3435);
or U3761 (N_3761,N_3502,N_3407);
xnor U3762 (N_3762,N_3424,N_3404);
nand U3763 (N_3763,N_3410,N_3488);
nand U3764 (N_3764,N_3449,N_3510);
or U3765 (N_3765,N_3429,N_3405);
nand U3766 (N_3766,N_3492,N_3516);
nand U3767 (N_3767,N_3451,N_3559);
and U3768 (N_3768,N_3516,N_3449);
nor U3769 (N_3769,N_3528,N_3556);
and U3770 (N_3770,N_3515,N_3489);
nand U3771 (N_3771,N_3401,N_3547);
xnor U3772 (N_3772,N_3557,N_3472);
or U3773 (N_3773,N_3518,N_3481);
and U3774 (N_3774,N_3480,N_3414);
and U3775 (N_3775,N_3455,N_3520);
and U3776 (N_3776,N_3450,N_3536);
or U3777 (N_3777,N_3497,N_3472);
and U3778 (N_3778,N_3429,N_3511);
or U3779 (N_3779,N_3402,N_3582);
or U3780 (N_3780,N_3452,N_3521);
nand U3781 (N_3781,N_3410,N_3553);
and U3782 (N_3782,N_3570,N_3521);
nand U3783 (N_3783,N_3415,N_3411);
xnor U3784 (N_3784,N_3587,N_3552);
and U3785 (N_3785,N_3597,N_3415);
nand U3786 (N_3786,N_3406,N_3551);
nand U3787 (N_3787,N_3564,N_3476);
and U3788 (N_3788,N_3590,N_3417);
or U3789 (N_3789,N_3465,N_3594);
or U3790 (N_3790,N_3459,N_3478);
nand U3791 (N_3791,N_3544,N_3469);
or U3792 (N_3792,N_3578,N_3430);
nand U3793 (N_3793,N_3497,N_3440);
and U3794 (N_3794,N_3426,N_3443);
and U3795 (N_3795,N_3561,N_3473);
nor U3796 (N_3796,N_3453,N_3417);
nor U3797 (N_3797,N_3416,N_3594);
nor U3798 (N_3798,N_3413,N_3552);
xnor U3799 (N_3799,N_3419,N_3576);
nor U3800 (N_3800,N_3763,N_3605);
and U3801 (N_3801,N_3772,N_3620);
or U3802 (N_3802,N_3780,N_3695);
xor U3803 (N_3803,N_3650,N_3731);
and U3804 (N_3804,N_3746,N_3729);
or U3805 (N_3805,N_3697,N_3642);
and U3806 (N_3806,N_3770,N_3724);
and U3807 (N_3807,N_3687,N_3730);
nor U3808 (N_3808,N_3779,N_3749);
and U3809 (N_3809,N_3771,N_3716);
or U3810 (N_3810,N_3703,N_3758);
or U3811 (N_3811,N_3723,N_3691);
or U3812 (N_3812,N_3663,N_3639);
nor U3813 (N_3813,N_3741,N_3698);
nor U3814 (N_3814,N_3757,N_3707);
xnor U3815 (N_3815,N_3641,N_3640);
xnor U3816 (N_3816,N_3683,N_3789);
xnor U3817 (N_3817,N_3783,N_3680);
nor U3818 (N_3818,N_3700,N_3765);
and U3819 (N_3819,N_3651,N_3662);
xnor U3820 (N_3820,N_3674,N_3714);
or U3821 (N_3821,N_3632,N_3617);
and U3822 (N_3822,N_3743,N_3769);
and U3823 (N_3823,N_3767,N_3694);
nand U3824 (N_3824,N_3709,N_3600);
or U3825 (N_3825,N_3619,N_3701);
nand U3826 (N_3826,N_3616,N_3615);
xor U3827 (N_3827,N_3720,N_3692);
or U3828 (N_3828,N_3686,N_3682);
or U3829 (N_3829,N_3670,N_3705);
and U3830 (N_3830,N_3602,N_3627);
xor U3831 (N_3831,N_3622,N_3603);
nor U3832 (N_3832,N_3638,N_3601);
xor U3833 (N_3833,N_3669,N_3630);
xor U3834 (N_3834,N_3702,N_3735);
and U3835 (N_3835,N_3634,N_3618);
xnor U3836 (N_3836,N_3665,N_3645);
or U3837 (N_3837,N_3752,N_3727);
nand U3838 (N_3838,N_3791,N_3636);
xor U3839 (N_3839,N_3678,N_3613);
nand U3840 (N_3840,N_3737,N_3748);
nor U3841 (N_3841,N_3629,N_3784);
xor U3842 (N_3842,N_3710,N_3736);
and U3843 (N_3843,N_3637,N_3732);
or U3844 (N_3844,N_3668,N_3607);
nor U3845 (N_3845,N_3631,N_3609);
or U3846 (N_3846,N_3798,N_3685);
nor U3847 (N_3847,N_3759,N_3704);
and U3848 (N_3848,N_3675,N_3681);
nor U3849 (N_3849,N_3679,N_3658);
nand U3850 (N_3850,N_3728,N_3734);
and U3851 (N_3851,N_3790,N_3725);
nor U3852 (N_3852,N_3676,N_3761);
xnor U3853 (N_3853,N_3626,N_3777);
and U3854 (N_3854,N_3795,N_3738);
nand U3855 (N_3855,N_3604,N_3797);
nor U3856 (N_3856,N_3677,N_3739);
and U3857 (N_3857,N_3733,N_3745);
xnor U3858 (N_3858,N_3712,N_3754);
xnor U3859 (N_3859,N_3690,N_3715);
nor U3860 (N_3860,N_3606,N_3778);
nor U3861 (N_3861,N_3646,N_3793);
nand U3862 (N_3862,N_3751,N_3661);
xor U3863 (N_3863,N_3711,N_3787);
or U3864 (N_3864,N_3647,N_3718);
nand U3865 (N_3865,N_3671,N_3689);
xnor U3866 (N_3866,N_3708,N_3699);
and U3867 (N_3867,N_3664,N_3776);
nor U3868 (N_3868,N_3688,N_3799);
and U3869 (N_3869,N_3696,N_3786);
xnor U3870 (N_3870,N_3717,N_3781);
or U3871 (N_3871,N_3766,N_3611);
nor U3872 (N_3872,N_3726,N_3623);
nand U3873 (N_3873,N_3653,N_3740);
or U3874 (N_3874,N_3614,N_3713);
nand U3875 (N_3875,N_3655,N_3764);
nand U3876 (N_3876,N_3782,N_3747);
and U3877 (N_3877,N_3672,N_3621);
nand U3878 (N_3878,N_3648,N_3649);
nor U3879 (N_3879,N_3744,N_3625);
nor U3880 (N_3880,N_3643,N_3721);
nand U3881 (N_3881,N_3775,N_3644);
nor U3882 (N_3882,N_3667,N_3773);
xnor U3883 (N_3883,N_3768,N_3755);
and U3884 (N_3884,N_3760,N_3774);
and U3885 (N_3885,N_3788,N_3666);
or U3886 (N_3886,N_3608,N_3656);
nand U3887 (N_3887,N_3753,N_3693);
and U3888 (N_3888,N_3610,N_3673);
nor U3889 (N_3889,N_3659,N_3796);
or U3890 (N_3890,N_3660,N_3794);
and U3891 (N_3891,N_3628,N_3654);
nand U3892 (N_3892,N_3792,N_3612);
or U3893 (N_3893,N_3742,N_3750);
nor U3894 (N_3894,N_3756,N_3652);
and U3895 (N_3895,N_3633,N_3635);
and U3896 (N_3896,N_3719,N_3762);
nor U3897 (N_3897,N_3706,N_3657);
nor U3898 (N_3898,N_3684,N_3722);
or U3899 (N_3899,N_3624,N_3785);
and U3900 (N_3900,N_3626,N_3779);
nor U3901 (N_3901,N_3783,N_3797);
nand U3902 (N_3902,N_3735,N_3757);
nor U3903 (N_3903,N_3695,N_3619);
nand U3904 (N_3904,N_3768,N_3641);
nand U3905 (N_3905,N_3737,N_3712);
xnor U3906 (N_3906,N_3706,N_3680);
or U3907 (N_3907,N_3656,N_3772);
and U3908 (N_3908,N_3726,N_3770);
and U3909 (N_3909,N_3642,N_3675);
nand U3910 (N_3910,N_3618,N_3636);
xnor U3911 (N_3911,N_3649,N_3797);
nand U3912 (N_3912,N_3682,N_3779);
and U3913 (N_3913,N_3711,N_3625);
xnor U3914 (N_3914,N_3624,N_3799);
or U3915 (N_3915,N_3797,N_3794);
xnor U3916 (N_3916,N_3616,N_3707);
nor U3917 (N_3917,N_3673,N_3686);
nor U3918 (N_3918,N_3660,N_3627);
nor U3919 (N_3919,N_3743,N_3710);
nand U3920 (N_3920,N_3690,N_3726);
nor U3921 (N_3921,N_3740,N_3619);
and U3922 (N_3922,N_3693,N_3610);
nand U3923 (N_3923,N_3640,N_3704);
and U3924 (N_3924,N_3717,N_3633);
and U3925 (N_3925,N_3733,N_3782);
and U3926 (N_3926,N_3774,N_3753);
and U3927 (N_3927,N_3698,N_3699);
and U3928 (N_3928,N_3756,N_3696);
and U3929 (N_3929,N_3686,N_3789);
and U3930 (N_3930,N_3690,N_3714);
nand U3931 (N_3931,N_3703,N_3685);
and U3932 (N_3932,N_3612,N_3774);
and U3933 (N_3933,N_3715,N_3684);
nand U3934 (N_3934,N_3773,N_3611);
xnor U3935 (N_3935,N_3697,N_3774);
nor U3936 (N_3936,N_3666,N_3613);
and U3937 (N_3937,N_3654,N_3620);
nor U3938 (N_3938,N_3693,N_3616);
nor U3939 (N_3939,N_3608,N_3612);
or U3940 (N_3940,N_3750,N_3743);
xor U3941 (N_3941,N_3717,N_3798);
nor U3942 (N_3942,N_3757,N_3625);
or U3943 (N_3943,N_3648,N_3792);
or U3944 (N_3944,N_3736,N_3739);
nand U3945 (N_3945,N_3747,N_3660);
xor U3946 (N_3946,N_3772,N_3609);
nand U3947 (N_3947,N_3660,N_3664);
and U3948 (N_3948,N_3635,N_3723);
or U3949 (N_3949,N_3727,N_3662);
and U3950 (N_3950,N_3789,N_3750);
or U3951 (N_3951,N_3690,N_3629);
or U3952 (N_3952,N_3691,N_3626);
and U3953 (N_3953,N_3697,N_3669);
and U3954 (N_3954,N_3633,N_3655);
or U3955 (N_3955,N_3692,N_3661);
and U3956 (N_3956,N_3730,N_3799);
nand U3957 (N_3957,N_3735,N_3732);
and U3958 (N_3958,N_3656,N_3723);
xor U3959 (N_3959,N_3763,N_3786);
nand U3960 (N_3960,N_3728,N_3604);
nor U3961 (N_3961,N_3696,N_3627);
xor U3962 (N_3962,N_3744,N_3707);
or U3963 (N_3963,N_3600,N_3719);
xnor U3964 (N_3964,N_3618,N_3752);
nor U3965 (N_3965,N_3746,N_3764);
xnor U3966 (N_3966,N_3755,N_3756);
or U3967 (N_3967,N_3633,N_3705);
or U3968 (N_3968,N_3755,N_3600);
nand U3969 (N_3969,N_3682,N_3790);
nand U3970 (N_3970,N_3792,N_3650);
or U3971 (N_3971,N_3714,N_3744);
or U3972 (N_3972,N_3683,N_3643);
or U3973 (N_3973,N_3614,N_3628);
and U3974 (N_3974,N_3785,N_3659);
nand U3975 (N_3975,N_3658,N_3718);
xor U3976 (N_3976,N_3607,N_3679);
nor U3977 (N_3977,N_3614,N_3601);
and U3978 (N_3978,N_3781,N_3687);
nand U3979 (N_3979,N_3608,N_3730);
or U3980 (N_3980,N_3773,N_3706);
nor U3981 (N_3981,N_3675,N_3672);
nand U3982 (N_3982,N_3653,N_3776);
nand U3983 (N_3983,N_3721,N_3750);
or U3984 (N_3984,N_3780,N_3685);
nand U3985 (N_3985,N_3764,N_3637);
nor U3986 (N_3986,N_3776,N_3651);
or U3987 (N_3987,N_3613,N_3749);
or U3988 (N_3988,N_3764,N_3653);
or U3989 (N_3989,N_3774,N_3729);
xnor U3990 (N_3990,N_3634,N_3685);
or U3991 (N_3991,N_3746,N_3618);
nand U3992 (N_3992,N_3795,N_3653);
xnor U3993 (N_3993,N_3623,N_3776);
or U3994 (N_3994,N_3701,N_3680);
nor U3995 (N_3995,N_3631,N_3708);
nor U3996 (N_3996,N_3730,N_3781);
or U3997 (N_3997,N_3611,N_3616);
nor U3998 (N_3998,N_3621,N_3766);
nand U3999 (N_3999,N_3611,N_3730);
xor U4000 (N_4000,N_3997,N_3948);
xnor U4001 (N_4001,N_3952,N_3837);
xor U4002 (N_4002,N_3895,N_3930);
nand U4003 (N_4003,N_3898,N_3935);
nand U4004 (N_4004,N_3867,N_3822);
and U4005 (N_4005,N_3974,N_3914);
and U4006 (N_4006,N_3820,N_3893);
nand U4007 (N_4007,N_3847,N_3912);
nand U4008 (N_4008,N_3814,N_3917);
xnor U4009 (N_4009,N_3943,N_3916);
nor U4010 (N_4010,N_3833,N_3955);
or U4011 (N_4011,N_3869,N_3828);
and U4012 (N_4012,N_3849,N_3964);
nor U4013 (N_4013,N_3963,N_3881);
nor U4014 (N_4014,N_3860,N_3823);
or U4015 (N_4015,N_3827,N_3976);
nand U4016 (N_4016,N_3989,N_3942);
nor U4017 (N_4017,N_3947,N_3929);
nand U4018 (N_4018,N_3959,N_3824);
xor U4019 (N_4019,N_3812,N_3938);
or U4020 (N_4020,N_3857,N_3856);
xnor U4021 (N_4021,N_3801,N_3834);
nand U4022 (N_4022,N_3874,N_3825);
xor U4023 (N_4023,N_3884,N_3858);
and U4024 (N_4024,N_3882,N_3870);
and U4025 (N_4025,N_3979,N_3831);
nor U4026 (N_4026,N_3971,N_3946);
and U4027 (N_4027,N_3954,N_3850);
nor U4028 (N_4028,N_3993,N_3908);
nor U4029 (N_4029,N_3889,N_3862);
xor U4030 (N_4030,N_3933,N_3809);
nor U4031 (N_4031,N_3965,N_3808);
xor U4032 (N_4032,N_3949,N_3939);
nand U4033 (N_4033,N_3996,N_3885);
nand U4034 (N_4034,N_3909,N_3932);
or U4035 (N_4035,N_3991,N_3977);
or U4036 (N_4036,N_3957,N_3852);
or U4037 (N_4037,N_3944,N_3805);
or U4038 (N_4038,N_3816,N_3998);
xor U4039 (N_4039,N_3980,N_3992);
or U4040 (N_4040,N_3941,N_3800);
nand U4041 (N_4041,N_3906,N_3864);
or U4042 (N_4042,N_3907,N_3928);
xnor U4043 (N_4043,N_3925,N_3960);
and U4044 (N_4044,N_3975,N_3888);
or U4045 (N_4045,N_3918,N_3830);
and U4046 (N_4046,N_3890,N_3863);
nand U4047 (N_4047,N_3972,N_3842);
xor U4048 (N_4048,N_3926,N_3902);
xnor U4049 (N_4049,N_3844,N_3995);
nand U4050 (N_4050,N_3877,N_3913);
xnor U4051 (N_4051,N_3923,N_3961);
xnor U4052 (N_4052,N_3802,N_3940);
and U4053 (N_4053,N_3845,N_3840);
and U4054 (N_4054,N_3866,N_3892);
or U4055 (N_4055,N_3900,N_3810);
nor U4056 (N_4056,N_3854,N_3829);
xnor U4057 (N_4057,N_3868,N_3910);
xnor U4058 (N_4058,N_3899,N_3851);
xor U4059 (N_4059,N_3886,N_3872);
and U4060 (N_4060,N_3966,N_3817);
nor U4061 (N_4061,N_3873,N_3968);
nor U4062 (N_4062,N_3970,N_3953);
or U4063 (N_4063,N_3988,N_3958);
and U4064 (N_4064,N_3861,N_3839);
or U4065 (N_4065,N_3818,N_3811);
or U4066 (N_4066,N_3876,N_3878);
and U4067 (N_4067,N_3990,N_3835);
or U4068 (N_4068,N_3894,N_3879);
or U4069 (N_4069,N_3813,N_3848);
nor U4070 (N_4070,N_3901,N_3987);
xnor U4071 (N_4071,N_3804,N_3821);
and U4072 (N_4072,N_3887,N_3999);
xor U4073 (N_4073,N_3846,N_3875);
nor U4074 (N_4074,N_3945,N_3956);
xnor U4075 (N_4075,N_3937,N_3896);
nand U4076 (N_4076,N_3982,N_3919);
xor U4077 (N_4077,N_3880,N_3826);
nor U4078 (N_4078,N_3819,N_3815);
or U4079 (N_4079,N_3934,N_3843);
xnor U4080 (N_4080,N_3859,N_3950);
nor U4081 (N_4081,N_3985,N_3903);
and U4082 (N_4082,N_3967,N_3951);
and U4083 (N_4083,N_3936,N_3883);
nand U4084 (N_4084,N_3891,N_3962);
nand U4085 (N_4085,N_3806,N_3986);
xnor U4086 (N_4086,N_3911,N_3920);
nand U4087 (N_4087,N_3807,N_3994);
or U4088 (N_4088,N_3855,N_3969);
and U4089 (N_4089,N_3921,N_3931);
or U4090 (N_4090,N_3897,N_3981);
nand U4091 (N_4091,N_3927,N_3871);
xor U4092 (N_4092,N_3841,N_3924);
nor U4093 (N_4093,N_3983,N_3984);
and U4094 (N_4094,N_3915,N_3905);
nand U4095 (N_4095,N_3838,N_3832);
xor U4096 (N_4096,N_3803,N_3973);
nand U4097 (N_4097,N_3836,N_3904);
xor U4098 (N_4098,N_3853,N_3978);
or U4099 (N_4099,N_3865,N_3922);
xnor U4100 (N_4100,N_3803,N_3820);
or U4101 (N_4101,N_3848,N_3923);
nor U4102 (N_4102,N_3905,N_3950);
xor U4103 (N_4103,N_3813,N_3840);
or U4104 (N_4104,N_3998,N_3897);
nor U4105 (N_4105,N_3836,N_3897);
nand U4106 (N_4106,N_3935,N_3881);
nand U4107 (N_4107,N_3889,N_3903);
or U4108 (N_4108,N_3887,N_3818);
nand U4109 (N_4109,N_3854,N_3922);
xor U4110 (N_4110,N_3920,N_3881);
xor U4111 (N_4111,N_3998,N_3874);
or U4112 (N_4112,N_3900,N_3928);
nand U4113 (N_4113,N_3831,N_3924);
or U4114 (N_4114,N_3970,N_3853);
xnor U4115 (N_4115,N_3826,N_3857);
xor U4116 (N_4116,N_3974,N_3998);
nor U4117 (N_4117,N_3971,N_3898);
xnor U4118 (N_4118,N_3897,N_3838);
or U4119 (N_4119,N_3859,N_3873);
nand U4120 (N_4120,N_3808,N_3921);
nor U4121 (N_4121,N_3800,N_3968);
or U4122 (N_4122,N_3871,N_3899);
or U4123 (N_4123,N_3929,N_3828);
nor U4124 (N_4124,N_3872,N_3826);
nor U4125 (N_4125,N_3824,N_3834);
and U4126 (N_4126,N_3859,N_3830);
and U4127 (N_4127,N_3893,N_3941);
or U4128 (N_4128,N_3839,N_3939);
or U4129 (N_4129,N_3943,N_3870);
nor U4130 (N_4130,N_3911,N_3824);
xnor U4131 (N_4131,N_3838,N_3805);
xor U4132 (N_4132,N_3934,N_3990);
and U4133 (N_4133,N_3993,N_3906);
xor U4134 (N_4134,N_3919,N_3966);
and U4135 (N_4135,N_3882,N_3872);
nor U4136 (N_4136,N_3904,N_3913);
or U4137 (N_4137,N_3976,N_3934);
or U4138 (N_4138,N_3934,N_3879);
or U4139 (N_4139,N_3948,N_3916);
xor U4140 (N_4140,N_3988,N_3836);
nand U4141 (N_4141,N_3961,N_3936);
nand U4142 (N_4142,N_3877,N_3959);
or U4143 (N_4143,N_3839,N_3871);
xor U4144 (N_4144,N_3903,N_3947);
and U4145 (N_4145,N_3852,N_3806);
or U4146 (N_4146,N_3980,N_3943);
xor U4147 (N_4147,N_3855,N_3833);
xnor U4148 (N_4148,N_3933,N_3930);
nor U4149 (N_4149,N_3853,N_3955);
or U4150 (N_4150,N_3855,N_3989);
xnor U4151 (N_4151,N_3902,N_3952);
nor U4152 (N_4152,N_3840,N_3981);
nor U4153 (N_4153,N_3999,N_3959);
or U4154 (N_4154,N_3975,N_3900);
xor U4155 (N_4155,N_3861,N_3918);
xnor U4156 (N_4156,N_3995,N_3892);
nand U4157 (N_4157,N_3941,N_3872);
xnor U4158 (N_4158,N_3874,N_3965);
xnor U4159 (N_4159,N_3909,N_3810);
nand U4160 (N_4160,N_3831,N_3871);
nor U4161 (N_4161,N_3871,N_3954);
nor U4162 (N_4162,N_3942,N_3918);
xnor U4163 (N_4163,N_3884,N_3894);
nor U4164 (N_4164,N_3824,N_3907);
nor U4165 (N_4165,N_3856,N_3940);
or U4166 (N_4166,N_3931,N_3981);
nor U4167 (N_4167,N_3953,N_3976);
nand U4168 (N_4168,N_3983,N_3877);
and U4169 (N_4169,N_3942,N_3827);
and U4170 (N_4170,N_3816,N_3899);
nor U4171 (N_4171,N_3990,N_3949);
or U4172 (N_4172,N_3823,N_3979);
nand U4173 (N_4173,N_3961,N_3972);
xnor U4174 (N_4174,N_3946,N_3814);
and U4175 (N_4175,N_3952,N_3944);
nor U4176 (N_4176,N_3891,N_3887);
xnor U4177 (N_4177,N_3858,N_3817);
nand U4178 (N_4178,N_3848,N_3945);
nor U4179 (N_4179,N_3826,N_3998);
xor U4180 (N_4180,N_3923,N_3972);
nand U4181 (N_4181,N_3991,N_3872);
xor U4182 (N_4182,N_3960,N_3974);
nand U4183 (N_4183,N_3984,N_3804);
nand U4184 (N_4184,N_3831,N_3884);
xnor U4185 (N_4185,N_3839,N_3980);
and U4186 (N_4186,N_3807,N_3804);
or U4187 (N_4187,N_3980,N_3901);
or U4188 (N_4188,N_3950,N_3866);
or U4189 (N_4189,N_3960,N_3800);
nor U4190 (N_4190,N_3987,N_3846);
and U4191 (N_4191,N_3839,N_3944);
xor U4192 (N_4192,N_3934,N_3956);
or U4193 (N_4193,N_3837,N_3980);
nor U4194 (N_4194,N_3985,N_3896);
nand U4195 (N_4195,N_3830,N_3974);
or U4196 (N_4196,N_3898,N_3881);
and U4197 (N_4197,N_3932,N_3929);
nor U4198 (N_4198,N_3982,N_3980);
and U4199 (N_4199,N_3850,N_3918);
nand U4200 (N_4200,N_4038,N_4137);
and U4201 (N_4201,N_4000,N_4189);
nor U4202 (N_4202,N_4020,N_4160);
xnor U4203 (N_4203,N_4106,N_4123);
nor U4204 (N_4204,N_4105,N_4126);
nor U4205 (N_4205,N_4179,N_4024);
xor U4206 (N_4206,N_4102,N_4018);
or U4207 (N_4207,N_4121,N_4188);
and U4208 (N_4208,N_4065,N_4031);
nand U4209 (N_4209,N_4153,N_4009);
or U4210 (N_4210,N_4028,N_4082);
xor U4211 (N_4211,N_4086,N_4149);
and U4212 (N_4212,N_4050,N_4130);
or U4213 (N_4213,N_4129,N_4017);
or U4214 (N_4214,N_4140,N_4139);
nand U4215 (N_4215,N_4035,N_4113);
nand U4216 (N_4216,N_4156,N_4045);
or U4217 (N_4217,N_4011,N_4055);
and U4218 (N_4218,N_4125,N_4063);
nor U4219 (N_4219,N_4138,N_4169);
and U4220 (N_4220,N_4044,N_4079);
xor U4221 (N_4221,N_4054,N_4145);
xor U4222 (N_4222,N_4144,N_4053);
nor U4223 (N_4223,N_4108,N_4095);
xor U4224 (N_4224,N_4034,N_4117);
and U4225 (N_4225,N_4192,N_4096);
nand U4226 (N_4226,N_4152,N_4157);
nand U4227 (N_4227,N_4074,N_4119);
or U4228 (N_4228,N_4143,N_4109);
or U4229 (N_4229,N_4110,N_4136);
nor U4230 (N_4230,N_4151,N_4097);
and U4231 (N_4231,N_4127,N_4042);
nor U4232 (N_4232,N_4002,N_4186);
or U4233 (N_4233,N_4070,N_4163);
and U4234 (N_4234,N_4159,N_4092);
and U4235 (N_4235,N_4003,N_4090);
and U4236 (N_4236,N_4041,N_4183);
nor U4237 (N_4237,N_4062,N_4164);
nand U4238 (N_4238,N_4019,N_4115);
xor U4239 (N_4239,N_4193,N_4030);
or U4240 (N_4240,N_4077,N_4036);
nor U4241 (N_4241,N_4161,N_4081);
and U4242 (N_4242,N_4158,N_4026);
xnor U4243 (N_4243,N_4133,N_4071);
xor U4244 (N_4244,N_4072,N_4083);
xnor U4245 (N_4245,N_4001,N_4069);
or U4246 (N_4246,N_4182,N_4124);
nand U4247 (N_4247,N_4175,N_4148);
xor U4248 (N_4248,N_4184,N_4104);
and U4249 (N_4249,N_4013,N_4005);
xnor U4250 (N_4250,N_4112,N_4174);
or U4251 (N_4251,N_4048,N_4196);
nor U4252 (N_4252,N_4191,N_4032);
nor U4253 (N_4253,N_4085,N_4103);
xor U4254 (N_4254,N_4190,N_4098);
xnor U4255 (N_4255,N_4194,N_4128);
or U4256 (N_4256,N_4195,N_4142);
nor U4257 (N_4257,N_4067,N_4166);
and U4258 (N_4258,N_4016,N_4116);
nand U4259 (N_4259,N_4014,N_4120);
xor U4260 (N_4260,N_4172,N_4033);
and U4261 (N_4261,N_4114,N_4150);
and U4262 (N_4262,N_4198,N_4061);
nand U4263 (N_4263,N_4073,N_4088);
nand U4264 (N_4264,N_4146,N_4049);
nor U4265 (N_4265,N_4084,N_4047);
nand U4266 (N_4266,N_4197,N_4165);
nor U4267 (N_4267,N_4135,N_4021);
and U4268 (N_4268,N_4051,N_4099);
and U4269 (N_4269,N_4122,N_4043);
and U4270 (N_4270,N_4101,N_4180);
and U4271 (N_4271,N_4037,N_4046);
nor U4272 (N_4272,N_4134,N_4171);
nor U4273 (N_4273,N_4176,N_4022);
and U4274 (N_4274,N_4181,N_4015);
nor U4275 (N_4275,N_4111,N_4170);
xor U4276 (N_4276,N_4004,N_4052);
nand U4277 (N_4277,N_4177,N_4199);
nand U4278 (N_4278,N_4185,N_4012);
nor U4279 (N_4279,N_4007,N_4080);
or U4280 (N_4280,N_4068,N_4039);
or U4281 (N_4281,N_4057,N_4075);
or U4282 (N_4282,N_4094,N_4078);
nand U4283 (N_4283,N_4155,N_4107);
xor U4284 (N_4284,N_4173,N_4187);
or U4285 (N_4285,N_4027,N_4132);
nor U4286 (N_4286,N_4006,N_4141);
and U4287 (N_4287,N_4058,N_4008);
nor U4288 (N_4288,N_4056,N_4089);
xnor U4289 (N_4289,N_4066,N_4059);
nor U4290 (N_4290,N_4162,N_4029);
xor U4291 (N_4291,N_4060,N_4167);
xor U4292 (N_4292,N_4023,N_4093);
nand U4293 (N_4293,N_4087,N_4091);
nand U4294 (N_4294,N_4147,N_4118);
nor U4295 (N_4295,N_4040,N_4154);
xor U4296 (N_4296,N_4168,N_4076);
nor U4297 (N_4297,N_4025,N_4131);
or U4298 (N_4298,N_4064,N_4010);
and U4299 (N_4299,N_4100,N_4178);
nor U4300 (N_4300,N_4159,N_4065);
nand U4301 (N_4301,N_4137,N_4019);
and U4302 (N_4302,N_4185,N_4001);
and U4303 (N_4303,N_4135,N_4070);
or U4304 (N_4304,N_4072,N_4146);
and U4305 (N_4305,N_4017,N_4059);
nand U4306 (N_4306,N_4174,N_4097);
nand U4307 (N_4307,N_4154,N_4043);
nand U4308 (N_4308,N_4025,N_4189);
nand U4309 (N_4309,N_4113,N_4178);
nor U4310 (N_4310,N_4140,N_4143);
or U4311 (N_4311,N_4019,N_4070);
or U4312 (N_4312,N_4115,N_4183);
nand U4313 (N_4313,N_4060,N_4048);
xnor U4314 (N_4314,N_4150,N_4052);
xnor U4315 (N_4315,N_4032,N_4124);
nand U4316 (N_4316,N_4159,N_4087);
or U4317 (N_4317,N_4148,N_4059);
xor U4318 (N_4318,N_4142,N_4166);
and U4319 (N_4319,N_4103,N_4041);
or U4320 (N_4320,N_4144,N_4011);
or U4321 (N_4321,N_4182,N_4078);
and U4322 (N_4322,N_4160,N_4041);
and U4323 (N_4323,N_4006,N_4014);
xor U4324 (N_4324,N_4156,N_4039);
or U4325 (N_4325,N_4049,N_4180);
and U4326 (N_4326,N_4199,N_4043);
and U4327 (N_4327,N_4018,N_4177);
nand U4328 (N_4328,N_4181,N_4079);
xnor U4329 (N_4329,N_4050,N_4196);
nor U4330 (N_4330,N_4070,N_4085);
nor U4331 (N_4331,N_4163,N_4011);
and U4332 (N_4332,N_4199,N_4082);
and U4333 (N_4333,N_4127,N_4031);
or U4334 (N_4334,N_4079,N_4025);
and U4335 (N_4335,N_4124,N_4081);
xnor U4336 (N_4336,N_4027,N_4119);
and U4337 (N_4337,N_4192,N_4060);
and U4338 (N_4338,N_4071,N_4140);
xor U4339 (N_4339,N_4142,N_4126);
or U4340 (N_4340,N_4173,N_4109);
xor U4341 (N_4341,N_4004,N_4046);
or U4342 (N_4342,N_4056,N_4117);
nor U4343 (N_4343,N_4037,N_4064);
xnor U4344 (N_4344,N_4026,N_4025);
xnor U4345 (N_4345,N_4100,N_4120);
and U4346 (N_4346,N_4090,N_4068);
xnor U4347 (N_4347,N_4155,N_4197);
nand U4348 (N_4348,N_4074,N_4123);
and U4349 (N_4349,N_4048,N_4132);
nor U4350 (N_4350,N_4033,N_4006);
xor U4351 (N_4351,N_4096,N_4113);
or U4352 (N_4352,N_4169,N_4146);
or U4353 (N_4353,N_4065,N_4035);
or U4354 (N_4354,N_4047,N_4128);
xnor U4355 (N_4355,N_4157,N_4175);
nor U4356 (N_4356,N_4125,N_4008);
nand U4357 (N_4357,N_4174,N_4188);
or U4358 (N_4358,N_4020,N_4055);
xnor U4359 (N_4359,N_4031,N_4039);
and U4360 (N_4360,N_4088,N_4009);
nand U4361 (N_4361,N_4133,N_4139);
and U4362 (N_4362,N_4049,N_4059);
and U4363 (N_4363,N_4008,N_4087);
nor U4364 (N_4364,N_4189,N_4039);
xnor U4365 (N_4365,N_4036,N_4149);
and U4366 (N_4366,N_4090,N_4010);
and U4367 (N_4367,N_4043,N_4170);
xor U4368 (N_4368,N_4011,N_4080);
nand U4369 (N_4369,N_4179,N_4118);
and U4370 (N_4370,N_4185,N_4122);
or U4371 (N_4371,N_4005,N_4199);
or U4372 (N_4372,N_4046,N_4103);
nor U4373 (N_4373,N_4175,N_4173);
and U4374 (N_4374,N_4028,N_4088);
and U4375 (N_4375,N_4070,N_4130);
and U4376 (N_4376,N_4118,N_4026);
or U4377 (N_4377,N_4190,N_4113);
and U4378 (N_4378,N_4144,N_4063);
nand U4379 (N_4379,N_4055,N_4015);
nand U4380 (N_4380,N_4002,N_4160);
or U4381 (N_4381,N_4004,N_4169);
and U4382 (N_4382,N_4047,N_4163);
xor U4383 (N_4383,N_4037,N_4051);
xnor U4384 (N_4384,N_4172,N_4023);
and U4385 (N_4385,N_4048,N_4186);
nor U4386 (N_4386,N_4015,N_4060);
and U4387 (N_4387,N_4169,N_4103);
nor U4388 (N_4388,N_4139,N_4149);
or U4389 (N_4389,N_4006,N_4068);
nand U4390 (N_4390,N_4060,N_4145);
and U4391 (N_4391,N_4040,N_4079);
or U4392 (N_4392,N_4053,N_4076);
or U4393 (N_4393,N_4046,N_4100);
nand U4394 (N_4394,N_4033,N_4191);
nor U4395 (N_4395,N_4150,N_4105);
or U4396 (N_4396,N_4157,N_4102);
nand U4397 (N_4397,N_4178,N_4032);
nor U4398 (N_4398,N_4086,N_4073);
nand U4399 (N_4399,N_4011,N_4082);
and U4400 (N_4400,N_4387,N_4353);
nor U4401 (N_4401,N_4279,N_4288);
and U4402 (N_4402,N_4377,N_4350);
and U4403 (N_4403,N_4366,N_4388);
or U4404 (N_4404,N_4363,N_4303);
nor U4405 (N_4405,N_4324,N_4310);
nand U4406 (N_4406,N_4392,N_4307);
xor U4407 (N_4407,N_4300,N_4340);
and U4408 (N_4408,N_4356,N_4370);
nand U4409 (N_4409,N_4260,N_4311);
nor U4410 (N_4410,N_4206,N_4229);
nand U4411 (N_4411,N_4373,N_4225);
xor U4412 (N_4412,N_4375,N_4272);
and U4413 (N_4413,N_4302,N_4331);
nand U4414 (N_4414,N_4251,N_4265);
and U4415 (N_4415,N_4298,N_4322);
nand U4416 (N_4416,N_4306,N_4355);
nand U4417 (N_4417,N_4367,N_4269);
nor U4418 (N_4418,N_4283,N_4284);
nor U4419 (N_4419,N_4320,N_4201);
and U4420 (N_4420,N_4282,N_4274);
and U4421 (N_4421,N_4285,N_4236);
and U4422 (N_4422,N_4220,N_4389);
nand U4423 (N_4423,N_4261,N_4250);
xor U4424 (N_4424,N_4384,N_4270);
nand U4425 (N_4425,N_4328,N_4200);
or U4426 (N_4426,N_4238,N_4278);
xnor U4427 (N_4427,N_4276,N_4266);
nor U4428 (N_4428,N_4241,N_4335);
and U4429 (N_4429,N_4309,N_4218);
nor U4430 (N_4430,N_4378,N_4330);
or U4431 (N_4431,N_4386,N_4286);
or U4432 (N_4432,N_4232,N_4348);
xnor U4433 (N_4433,N_4243,N_4374);
nand U4434 (N_4434,N_4334,N_4364);
xnor U4435 (N_4435,N_4227,N_4344);
nand U4436 (N_4436,N_4259,N_4319);
or U4437 (N_4437,N_4214,N_4228);
and U4438 (N_4438,N_4380,N_4358);
or U4439 (N_4439,N_4365,N_4290);
nand U4440 (N_4440,N_4346,N_4233);
or U4441 (N_4441,N_4394,N_4264);
or U4442 (N_4442,N_4297,N_4205);
and U4443 (N_4443,N_4219,N_4230);
or U4444 (N_4444,N_4313,N_4254);
and U4445 (N_4445,N_4361,N_4369);
or U4446 (N_4446,N_4224,N_4234);
or U4447 (N_4447,N_4291,N_4372);
and U4448 (N_4448,N_4376,N_4294);
and U4449 (N_4449,N_4256,N_4336);
and U4450 (N_4450,N_4247,N_4327);
xor U4451 (N_4451,N_4223,N_4204);
and U4452 (N_4452,N_4292,N_4257);
nor U4453 (N_4453,N_4317,N_4221);
or U4454 (N_4454,N_4397,N_4385);
nand U4455 (N_4455,N_4301,N_4337);
nor U4456 (N_4456,N_4249,N_4399);
or U4457 (N_4457,N_4347,N_4333);
nand U4458 (N_4458,N_4314,N_4202);
and U4459 (N_4459,N_4352,N_4273);
and U4460 (N_4460,N_4326,N_4289);
nor U4461 (N_4461,N_4296,N_4240);
xor U4462 (N_4462,N_4357,N_4210);
nor U4463 (N_4463,N_4381,N_4299);
nand U4464 (N_4464,N_4354,N_4262);
and U4465 (N_4465,N_4245,N_4360);
or U4466 (N_4466,N_4237,N_4242);
xor U4467 (N_4467,N_4305,N_4208);
or U4468 (N_4468,N_4382,N_4213);
nand U4469 (N_4469,N_4215,N_4255);
xnor U4470 (N_4470,N_4342,N_4258);
or U4471 (N_4471,N_4235,N_4246);
nand U4472 (N_4472,N_4339,N_4281);
or U4473 (N_4473,N_4318,N_4398);
xnor U4474 (N_4474,N_4287,N_4226);
or U4475 (N_4475,N_4304,N_4351);
xor U4476 (N_4476,N_4393,N_4308);
nor U4477 (N_4477,N_4341,N_4280);
nor U4478 (N_4478,N_4332,N_4212);
nand U4479 (N_4479,N_4203,N_4277);
nor U4480 (N_4480,N_4343,N_4396);
or U4481 (N_4481,N_4263,N_4345);
nor U4482 (N_4482,N_4252,N_4222);
and U4483 (N_4483,N_4329,N_4391);
and U4484 (N_4484,N_4248,N_4379);
xnor U4485 (N_4485,N_4268,N_4209);
nor U4486 (N_4486,N_4368,N_4216);
and U4487 (N_4487,N_4315,N_4349);
xnor U4488 (N_4488,N_4275,N_4323);
nor U4489 (N_4489,N_4207,N_4316);
xor U4490 (N_4490,N_4211,N_4395);
xnor U4491 (N_4491,N_4362,N_4371);
nor U4492 (N_4492,N_4321,N_4295);
nor U4493 (N_4493,N_4244,N_4217);
xnor U4494 (N_4494,N_4312,N_4338);
and U4495 (N_4495,N_4383,N_4239);
nand U4496 (N_4496,N_4325,N_4267);
nand U4497 (N_4497,N_4359,N_4253);
and U4498 (N_4498,N_4231,N_4390);
xnor U4499 (N_4499,N_4293,N_4271);
or U4500 (N_4500,N_4294,N_4387);
xnor U4501 (N_4501,N_4200,N_4319);
xor U4502 (N_4502,N_4210,N_4380);
or U4503 (N_4503,N_4356,N_4345);
xor U4504 (N_4504,N_4332,N_4243);
or U4505 (N_4505,N_4300,N_4374);
nand U4506 (N_4506,N_4294,N_4370);
xnor U4507 (N_4507,N_4279,N_4224);
and U4508 (N_4508,N_4346,N_4272);
xnor U4509 (N_4509,N_4294,N_4286);
nand U4510 (N_4510,N_4360,N_4288);
or U4511 (N_4511,N_4379,N_4241);
and U4512 (N_4512,N_4261,N_4236);
or U4513 (N_4513,N_4369,N_4315);
xnor U4514 (N_4514,N_4258,N_4398);
xnor U4515 (N_4515,N_4321,N_4350);
xnor U4516 (N_4516,N_4368,N_4221);
xor U4517 (N_4517,N_4355,N_4246);
nand U4518 (N_4518,N_4374,N_4224);
and U4519 (N_4519,N_4208,N_4337);
nor U4520 (N_4520,N_4396,N_4304);
or U4521 (N_4521,N_4218,N_4302);
nand U4522 (N_4522,N_4394,N_4274);
nand U4523 (N_4523,N_4299,N_4217);
nor U4524 (N_4524,N_4286,N_4367);
and U4525 (N_4525,N_4282,N_4359);
or U4526 (N_4526,N_4313,N_4293);
nand U4527 (N_4527,N_4313,N_4227);
and U4528 (N_4528,N_4399,N_4346);
or U4529 (N_4529,N_4327,N_4293);
xnor U4530 (N_4530,N_4305,N_4304);
and U4531 (N_4531,N_4392,N_4267);
xor U4532 (N_4532,N_4209,N_4262);
nand U4533 (N_4533,N_4207,N_4332);
xor U4534 (N_4534,N_4238,N_4208);
and U4535 (N_4535,N_4351,N_4355);
or U4536 (N_4536,N_4278,N_4269);
nand U4537 (N_4537,N_4329,N_4335);
nor U4538 (N_4538,N_4204,N_4239);
nand U4539 (N_4539,N_4371,N_4304);
or U4540 (N_4540,N_4313,N_4392);
xor U4541 (N_4541,N_4266,N_4296);
nand U4542 (N_4542,N_4228,N_4394);
xor U4543 (N_4543,N_4238,N_4324);
nor U4544 (N_4544,N_4280,N_4316);
and U4545 (N_4545,N_4219,N_4319);
nand U4546 (N_4546,N_4360,N_4228);
xor U4547 (N_4547,N_4213,N_4229);
or U4548 (N_4548,N_4313,N_4217);
and U4549 (N_4549,N_4338,N_4319);
nand U4550 (N_4550,N_4275,N_4353);
xor U4551 (N_4551,N_4286,N_4353);
nand U4552 (N_4552,N_4299,N_4294);
nand U4553 (N_4553,N_4379,N_4362);
xnor U4554 (N_4554,N_4295,N_4297);
xnor U4555 (N_4555,N_4258,N_4338);
xor U4556 (N_4556,N_4315,N_4338);
nand U4557 (N_4557,N_4393,N_4218);
and U4558 (N_4558,N_4389,N_4207);
and U4559 (N_4559,N_4361,N_4237);
or U4560 (N_4560,N_4289,N_4355);
and U4561 (N_4561,N_4224,N_4325);
xor U4562 (N_4562,N_4392,N_4360);
or U4563 (N_4563,N_4342,N_4395);
xor U4564 (N_4564,N_4269,N_4284);
nand U4565 (N_4565,N_4276,N_4330);
nand U4566 (N_4566,N_4372,N_4348);
or U4567 (N_4567,N_4269,N_4245);
nand U4568 (N_4568,N_4393,N_4256);
xnor U4569 (N_4569,N_4360,N_4223);
nor U4570 (N_4570,N_4324,N_4239);
or U4571 (N_4571,N_4334,N_4213);
nand U4572 (N_4572,N_4312,N_4226);
or U4573 (N_4573,N_4340,N_4362);
xor U4574 (N_4574,N_4327,N_4364);
xnor U4575 (N_4575,N_4305,N_4219);
nor U4576 (N_4576,N_4224,N_4343);
nor U4577 (N_4577,N_4305,N_4294);
or U4578 (N_4578,N_4307,N_4364);
or U4579 (N_4579,N_4262,N_4359);
nand U4580 (N_4580,N_4306,N_4282);
nor U4581 (N_4581,N_4330,N_4312);
or U4582 (N_4582,N_4327,N_4357);
nand U4583 (N_4583,N_4251,N_4349);
xnor U4584 (N_4584,N_4378,N_4286);
or U4585 (N_4585,N_4348,N_4362);
and U4586 (N_4586,N_4238,N_4382);
xnor U4587 (N_4587,N_4307,N_4315);
and U4588 (N_4588,N_4271,N_4316);
xnor U4589 (N_4589,N_4386,N_4394);
nand U4590 (N_4590,N_4262,N_4232);
nand U4591 (N_4591,N_4359,N_4387);
and U4592 (N_4592,N_4264,N_4382);
and U4593 (N_4593,N_4235,N_4252);
nor U4594 (N_4594,N_4340,N_4399);
and U4595 (N_4595,N_4353,N_4346);
or U4596 (N_4596,N_4312,N_4306);
xor U4597 (N_4597,N_4391,N_4285);
nand U4598 (N_4598,N_4394,N_4381);
xor U4599 (N_4599,N_4284,N_4361);
xor U4600 (N_4600,N_4517,N_4552);
nor U4601 (N_4601,N_4476,N_4420);
and U4602 (N_4602,N_4512,N_4563);
or U4603 (N_4603,N_4482,N_4421);
and U4604 (N_4604,N_4477,N_4435);
xor U4605 (N_4605,N_4429,N_4442);
or U4606 (N_4606,N_4572,N_4496);
nor U4607 (N_4607,N_4515,N_4587);
or U4608 (N_4608,N_4493,N_4440);
or U4609 (N_4609,N_4504,N_4510);
nand U4610 (N_4610,N_4549,N_4413);
and U4611 (N_4611,N_4414,N_4540);
nand U4612 (N_4612,N_4415,N_4447);
nor U4613 (N_4613,N_4561,N_4526);
nor U4614 (N_4614,N_4524,N_4509);
xor U4615 (N_4615,N_4468,N_4424);
and U4616 (N_4616,N_4588,N_4575);
nor U4617 (N_4617,N_4412,N_4558);
and U4618 (N_4618,N_4450,N_4426);
and U4619 (N_4619,N_4556,N_4436);
nand U4620 (N_4620,N_4446,N_4590);
nand U4621 (N_4621,N_4551,N_4580);
and U4622 (N_4622,N_4569,N_4539);
and U4623 (N_4623,N_4579,N_4439);
xnor U4624 (N_4624,N_4488,N_4459);
xnor U4625 (N_4625,N_4487,N_4423);
nand U4626 (N_4626,N_4438,N_4567);
nand U4627 (N_4627,N_4576,N_4529);
nor U4628 (N_4628,N_4547,N_4598);
and U4629 (N_4629,N_4416,N_4407);
or U4630 (N_4630,N_4503,N_4479);
nor U4631 (N_4631,N_4577,N_4400);
xor U4632 (N_4632,N_4462,N_4451);
nand U4633 (N_4633,N_4571,N_4536);
and U4634 (N_4634,N_4546,N_4570);
nand U4635 (N_4635,N_4521,N_4453);
xor U4636 (N_4636,N_4417,N_4403);
and U4637 (N_4637,N_4454,N_4508);
or U4638 (N_4638,N_4537,N_4593);
and U4639 (N_4639,N_4452,N_4455);
xor U4640 (N_4640,N_4486,N_4520);
and U4641 (N_4641,N_4485,N_4513);
nor U4642 (N_4642,N_4554,N_4463);
nor U4643 (N_4643,N_4557,N_4464);
xnor U4644 (N_4644,N_4528,N_4499);
xor U4645 (N_4645,N_4497,N_4523);
nand U4646 (N_4646,N_4469,N_4430);
or U4647 (N_4647,N_4568,N_4583);
nand U4648 (N_4648,N_4458,N_4530);
nand U4649 (N_4649,N_4475,N_4449);
or U4650 (N_4650,N_4507,N_4465);
xor U4651 (N_4651,N_4408,N_4585);
xor U4652 (N_4652,N_4544,N_4481);
nand U4653 (N_4653,N_4584,N_4592);
or U4654 (N_4654,N_4518,N_4428);
xnor U4655 (N_4655,N_4589,N_4532);
nand U4656 (N_4656,N_4514,N_4456);
and U4657 (N_4657,N_4472,N_4595);
xnor U4658 (N_4658,N_4578,N_4427);
nor U4659 (N_4659,N_4445,N_4555);
or U4660 (N_4660,N_4506,N_4565);
xor U4661 (N_4661,N_4574,N_4418);
or U4662 (N_4662,N_4527,N_4550);
and U4663 (N_4663,N_4591,N_4562);
or U4664 (N_4664,N_4419,N_4534);
nor U4665 (N_4665,N_4564,N_4502);
or U4666 (N_4666,N_4494,N_4525);
or U4667 (N_4667,N_4483,N_4522);
nand U4668 (N_4668,N_4448,N_4410);
xnor U4669 (N_4669,N_4501,N_4582);
nand U4670 (N_4670,N_4489,N_4581);
nor U4671 (N_4671,N_4535,N_4531);
nor U4672 (N_4672,N_4441,N_4559);
xor U4673 (N_4673,N_4470,N_4492);
nor U4674 (N_4674,N_4480,N_4511);
nand U4675 (N_4675,N_4533,N_4437);
nand U4676 (N_4676,N_4457,N_4586);
xor U4677 (N_4677,N_4432,N_4594);
and U4678 (N_4678,N_4573,N_4484);
xor U4679 (N_4679,N_4466,N_4471);
xor U4680 (N_4680,N_4596,N_4473);
nand U4681 (N_4681,N_4434,N_4411);
nor U4682 (N_4682,N_4505,N_4566);
xor U4683 (N_4683,N_4542,N_4498);
xnor U4684 (N_4684,N_4545,N_4516);
or U4685 (N_4685,N_4560,N_4405);
or U4686 (N_4686,N_4543,N_4460);
xnor U4687 (N_4687,N_4425,N_4433);
or U4688 (N_4688,N_4553,N_4597);
and U4689 (N_4689,N_4548,N_4431);
or U4690 (N_4690,N_4599,N_4500);
nor U4691 (N_4691,N_4406,N_4519);
nor U4692 (N_4692,N_4478,N_4409);
xor U4693 (N_4693,N_4444,N_4461);
and U4694 (N_4694,N_4491,N_4474);
nor U4695 (N_4695,N_4422,N_4467);
xor U4696 (N_4696,N_4541,N_4495);
xnor U4697 (N_4697,N_4443,N_4538);
nand U4698 (N_4698,N_4490,N_4404);
nand U4699 (N_4699,N_4401,N_4402);
and U4700 (N_4700,N_4501,N_4424);
and U4701 (N_4701,N_4549,N_4425);
nand U4702 (N_4702,N_4511,N_4433);
nand U4703 (N_4703,N_4491,N_4413);
and U4704 (N_4704,N_4459,N_4482);
and U4705 (N_4705,N_4478,N_4437);
nor U4706 (N_4706,N_4524,N_4528);
or U4707 (N_4707,N_4543,N_4482);
and U4708 (N_4708,N_4542,N_4483);
nand U4709 (N_4709,N_4449,N_4458);
xor U4710 (N_4710,N_4582,N_4439);
nand U4711 (N_4711,N_4530,N_4459);
and U4712 (N_4712,N_4555,N_4573);
nor U4713 (N_4713,N_4497,N_4495);
or U4714 (N_4714,N_4402,N_4482);
nor U4715 (N_4715,N_4439,N_4577);
or U4716 (N_4716,N_4441,N_4452);
and U4717 (N_4717,N_4426,N_4563);
nand U4718 (N_4718,N_4548,N_4580);
nand U4719 (N_4719,N_4494,N_4582);
xnor U4720 (N_4720,N_4529,N_4557);
xnor U4721 (N_4721,N_4410,N_4521);
xor U4722 (N_4722,N_4435,N_4580);
and U4723 (N_4723,N_4572,N_4481);
and U4724 (N_4724,N_4599,N_4403);
nor U4725 (N_4725,N_4501,N_4503);
nor U4726 (N_4726,N_4591,N_4467);
and U4727 (N_4727,N_4415,N_4503);
nand U4728 (N_4728,N_4558,N_4500);
and U4729 (N_4729,N_4404,N_4546);
or U4730 (N_4730,N_4524,N_4551);
and U4731 (N_4731,N_4553,N_4473);
or U4732 (N_4732,N_4451,N_4535);
xor U4733 (N_4733,N_4596,N_4494);
nand U4734 (N_4734,N_4549,N_4566);
or U4735 (N_4735,N_4513,N_4571);
or U4736 (N_4736,N_4410,N_4458);
nor U4737 (N_4737,N_4499,N_4410);
xnor U4738 (N_4738,N_4514,N_4482);
nand U4739 (N_4739,N_4585,N_4544);
nor U4740 (N_4740,N_4433,N_4447);
xor U4741 (N_4741,N_4576,N_4481);
and U4742 (N_4742,N_4477,N_4462);
or U4743 (N_4743,N_4432,N_4463);
nor U4744 (N_4744,N_4492,N_4457);
nand U4745 (N_4745,N_4584,N_4567);
xnor U4746 (N_4746,N_4517,N_4509);
xor U4747 (N_4747,N_4515,N_4439);
or U4748 (N_4748,N_4428,N_4412);
and U4749 (N_4749,N_4427,N_4505);
nor U4750 (N_4750,N_4411,N_4527);
nor U4751 (N_4751,N_4428,N_4413);
or U4752 (N_4752,N_4550,N_4535);
and U4753 (N_4753,N_4573,N_4496);
nand U4754 (N_4754,N_4533,N_4491);
nand U4755 (N_4755,N_4591,N_4597);
nand U4756 (N_4756,N_4565,N_4454);
and U4757 (N_4757,N_4561,N_4592);
nor U4758 (N_4758,N_4493,N_4425);
nand U4759 (N_4759,N_4584,N_4501);
xor U4760 (N_4760,N_4441,N_4567);
nand U4761 (N_4761,N_4548,N_4516);
nand U4762 (N_4762,N_4581,N_4593);
or U4763 (N_4763,N_4456,N_4528);
nand U4764 (N_4764,N_4506,N_4521);
xnor U4765 (N_4765,N_4542,N_4475);
nand U4766 (N_4766,N_4455,N_4456);
and U4767 (N_4767,N_4432,N_4514);
nor U4768 (N_4768,N_4526,N_4551);
nor U4769 (N_4769,N_4435,N_4450);
nand U4770 (N_4770,N_4411,N_4460);
and U4771 (N_4771,N_4572,N_4415);
nand U4772 (N_4772,N_4473,N_4545);
or U4773 (N_4773,N_4586,N_4437);
nand U4774 (N_4774,N_4442,N_4443);
and U4775 (N_4775,N_4556,N_4552);
nor U4776 (N_4776,N_4508,N_4588);
and U4777 (N_4777,N_4461,N_4449);
nor U4778 (N_4778,N_4512,N_4427);
or U4779 (N_4779,N_4521,N_4447);
or U4780 (N_4780,N_4515,N_4412);
and U4781 (N_4781,N_4530,N_4543);
xor U4782 (N_4782,N_4462,N_4510);
and U4783 (N_4783,N_4575,N_4538);
and U4784 (N_4784,N_4594,N_4542);
nand U4785 (N_4785,N_4543,N_4559);
and U4786 (N_4786,N_4575,N_4531);
xnor U4787 (N_4787,N_4594,N_4497);
nor U4788 (N_4788,N_4452,N_4410);
nand U4789 (N_4789,N_4533,N_4451);
or U4790 (N_4790,N_4591,N_4519);
or U4791 (N_4791,N_4480,N_4477);
xnor U4792 (N_4792,N_4429,N_4515);
or U4793 (N_4793,N_4504,N_4568);
and U4794 (N_4794,N_4459,N_4479);
and U4795 (N_4795,N_4487,N_4559);
xor U4796 (N_4796,N_4510,N_4446);
and U4797 (N_4797,N_4505,N_4548);
xnor U4798 (N_4798,N_4515,N_4516);
nor U4799 (N_4799,N_4593,N_4559);
nor U4800 (N_4800,N_4749,N_4693);
xor U4801 (N_4801,N_4682,N_4611);
nand U4802 (N_4802,N_4788,N_4783);
and U4803 (N_4803,N_4677,N_4624);
or U4804 (N_4804,N_4644,N_4623);
xnor U4805 (N_4805,N_4640,N_4722);
and U4806 (N_4806,N_4610,N_4637);
nor U4807 (N_4807,N_4731,N_4621);
nor U4808 (N_4808,N_4703,N_4650);
nor U4809 (N_4809,N_4771,N_4684);
and U4810 (N_4810,N_4665,N_4736);
nor U4811 (N_4811,N_4674,N_4725);
or U4812 (N_4812,N_4666,N_4799);
and U4813 (N_4813,N_4638,N_4766);
nor U4814 (N_4814,N_4661,N_4676);
or U4815 (N_4815,N_4795,N_4695);
and U4816 (N_4816,N_4601,N_4648);
or U4817 (N_4817,N_4691,N_4656);
nand U4818 (N_4818,N_4748,N_4777);
nand U4819 (N_4819,N_4701,N_4641);
or U4820 (N_4820,N_4635,N_4616);
or U4821 (N_4821,N_4762,N_4719);
and U4822 (N_4822,N_4600,N_4755);
nor U4823 (N_4823,N_4752,N_4697);
and U4824 (N_4824,N_4655,N_4652);
xor U4825 (N_4825,N_4653,N_4796);
xnor U4826 (N_4826,N_4679,N_4759);
xnor U4827 (N_4827,N_4617,N_4761);
nand U4828 (N_4828,N_4706,N_4729);
nor U4829 (N_4829,N_4605,N_4692);
nor U4830 (N_4830,N_4724,N_4780);
or U4831 (N_4831,N_4782,N_4757);
or U4832 (N_4832,N_4734,N_4769);
xnor U4833 (N_4833,N_4668,N_4713);
xnor U4834 (N_4834,N_4707,N_4768);
and U4835 (N_4835,N_4700,N_4794);
nor U4836 (N_4836,N_4797,N_4791);
and U4837 (N_4837,N_4711,N_4717);
nand U4838 (N_4838,N_4720,N_4699);
or U4839 (N_4839,N_4739,N_4613);
nand U4840 (N_4840,N_4745,N_4727);
or U4841 (N_4841,N_4747,N_4758);
or U4842 (N_4842,N_4680,N_4667);
or U4843 (N_4843,N_4726,N_4615);
or U4844 (N_4844,N_4781,N_4715);
xor U4845 (N_4845,N_4733,N_4678);
or U4846 (N_4846,N_4741,N_4622);
nand U4847 (N_4847,N_4658,N_4612);
xnor U4848 (N_4848,N_4772,N_4645);
or U4849 (N_4849,N_4790,N_4639);
or U4850 (N_4850,N_4643,N_4633);
xor U4851 (N_4851,N_4778,N_4606);
nand U4852 (N_4852,N_4642,N_4628);
or U4853 (N_4853,N_4764,N_4798);
and U4854 (N_4854,N_4709,N_4705);
nor U4855 (N_4855,N_4664,N_4785);
xnor U4856 (N_4856,N_4730,N_4632);
xor U4857 (N_4857,N_4685,N_4634);
and U4858 (N_4858,N_4604,N_4723);
xnor U4859 (N_4859,N_4689,N_4753);
nand U4860 (N_4860,N_4712,N_4620);
nor U4861 (N_4861,N_4649,N_4625);
nor U4862 (N_4862,N_4735,N_4698);
nand U4863 (N_4863,N_4763,N_4728);
xnor U4864 (N_4864,N_4789,N_4609);
nor U4865 (N_4865,N_4631,N_4687);
nor U4866 (N_4866,N_4629,N_4646);
and U4867 (N_4867,N_4660,N_4688);
and U4868 (N_4868,N_4746,N_4710);
and U4869 (N_4869,N_4670,N_4740);
or U4870 (N_4870,N_4792,N_4770);
and U4871 (N_4871,N_4627,N_4702);
or U4872 (N_4872,N_4614,N_4742);
nor U4873 (N_4873,N_4737,N_4651);
nor U4874 (N_4874,N_4662,N_4619);
and U4875 (N_4875,N_4750,N_4767);
xor U4876 (N_4876,N_4659,N_4779);
and U4877 (N_4877,N_4793,N_4681);
nand U4878 (N_4878,N_4671,N_4602);
or U4879 (N_4879,N_4683,N_4760);
nor U4880 (N_4880,N_4672,N_4721);
nand U4881 (N_4881,N_4751,N_4608);
nor U4882 (N_4882,N_4776,N_4630);
xor U4883 (N_4883,N_4716,N_4773);
or U4884 (N_4884,N_4765,N_4690);
or U4885 (N_4885,N_4756,N_4626);
nand U4886 (N_4886,N_4675,N_4663);
nor U4887 (N_4887,N_4714,N_4673);
nand U4888 (N_4888,N_4607,N_4718);
xnor U4889 (N_4889,N_4786,N_4775);
nand U4890 (N_4890,N_4738,N_4603);
nor U4891 (N_4891,N_4744,N_4636);
nand U4892 (N_4892,N_4654,N_4787);
xor U4893 (N_4893,N_4618,N_4696);
nand U4894 (N_4894,N_4784,N_4754);
xnor U4895 (N_4895,N_4647,N_4732);
or U4896 (N_4896,N_4657,N_4743);
nand U4897 (N_4897,N_4708,N_4686);
nor U4898 (N_4898,N_4669,N_4774);
or U4899 (N_4899,N_4704,N_4694);
or U4900 (N_4900,N_4747,N_4725);
or U4901 (N_4901,N_4660,N_4715);
or U4902 (N_4902,N_4736,N_4776);
and U4903 (N_4903,N_4699,N_4746);
nand U4904 (N_4904,N_4768,N_4794);
nand U4905 (N_4905,N_4744,N_4622);
and U4906 (N_4906,N_4695,N_4771);
nor U4907 (N_4907,N_4768,N_4618);
or U4908 (N_4908,N_4645,N_4749);
nand U4909 (N_4909,N_4601,N_4765);
or U4910 (N_4910,N_4763,N_4766);
nor U4911 (N_4911,N_4757,N_4610);
nand U4912 (N_4912,N_4666,N_4797);
nor U4913 (N_4913,N_4654,N_4698);
or U4914 (N_4914,N_4760,N_4609);
nor U4915 (N_4915,N_4711,N_4691);
or U4916 (N_4916,N_4737,N_4706);
xnor U4917 (N_4917,N_4664,N_4681);
and U4918 (N_4918,N_4742,N_4679);
and U4919 (N_4919,N_4657,N_4642);
nor U4920 (N_4920,N_4683,N_4654);
nand U4921 (N_4921,N_4769,N_4612);
xnor U4922 (N_4922,N_4784,N_4636);
nor U4923 (N_4923,N_4693,N_4700);
or U4924 (N_4924,N_4672,N_4768);
xor U4925 (N_4925,N_4617,N_4647);
xnor U4926 (N_4926,N_4789,N_4734);
xnor U4927 (N_4927,N_4677,N_4763);
nor U4928 (N_4928,N_4703,N_4765);
nor U4929 (N_4929,N_4677,N_4686);
xor U4930 (N_4930,N_4708,N_4795);
or U4931 (N_4931,N_4607,N_4747);
nand U4932 (N_4932,N_4741,N_4736);
nand U4933 (N_4933,N_4715,N_4699);
and U4934 (N_4934,N_4693,N_4629);
or U4935 (N_4935,N_4788,N_4647);
nand U4936 (N_4936,N_4739,N_4797);
or U4937 (N_4937,N_4693,N_4762);
and U4938 (N_4938,N_4775,N_4746);
or U4939 (N_4939,N_4759,N_4671);
nand U4940 (N_4940,N_4798,N_4684);
and U4941 (N_4941,N_4754,N_4687);
nand U4942 (N_4942,N_4699,N_4791);
nor U4943 (N_4943,N_4679,N_4733);
xor U4944 (N_4944,N_4796,N_4656);
nand U4945 (N_4945,N_4735,N_4605);
and U4946 (N_4946,N_4647,N_4630);
and U4947 (N_4947,N_4685,N_4728);
or U4948 (N_4948,N_4611,N_4767);
nor U4949 (N_4949,N_4755,N_4729);
nand U4950 (N_4950,N_4657,N_4777);
or U4951 (N_4951,N_4707,N_4673);
or U4952 (N_4952,N_4679,N_4746);
nand U4953 (N_4953,N_4727,N_4671);
nand U4954 (N_4954,N_4641,N_4620);
xor U4955 (N_4955,N_4680,N_4689);
nor U4956 (N_4956,N_4674,N_4658);
and U4957 (N_4957,N_4700,N_4630);
xnor U4958 (N_4958,N_4693,N_4784);
xor U4959 (N_4959,N_4634,N_4795);
xor U4960 (N_4960,N_4655,N_4725);
xor U4961 (N_4961,N_4706,N_4718);
nand U4962 (N_4962,N_4696,N_4656);
and U4963 (N_4963,N_4638,N_4719);
and U4964 (N_4964,N_4625,N_4787);
nand U4965 (N_4965,N_4767,N_4704);
nor U4966 (N_4966,N_4729,N_4633);
or U4967 (N_4967,N_4795,N_4799);
or U4968 (N_4968,N_4781,N_4734);
xnor U4969 (N_4969,N_4674,N_4693);
xor U4970 (N_4970,N_4756,N_4753);
nor U4971 (N_4971,N_4779,N_4791);
and U4972 (N_4972,N_4643,N_4708);
and U4973 (N_4973,N_4634,N_4741);
or U4974 (N_4974,N_4686,N_4745);
nand U4975 (N_4975,N_4646,N_4692);
xnor U4976 (N_4976,N_4698,N_4633);
xor U4977 (N_4977,N_4799,N_4697);
xnor U4978 (N_4978,N_4741,N_4632);
nor U4979 (N_4979,N_4629,N_4668);
nor U4980 (N_4980,N_4639,N_4716);
or U4981 (N_4981,N_4730,N_4759);
nand U4982 (N_4982,N_4648,N_4627);
nand U4983 (N_4983,N_4627,N_4703);
xnor U4984 (N_4984,N_4679,N_4617);
xor U4985 (N_4985,N_4656,N_4737);
nor U4986 (N_4986,N_4627,N_4754);
nand U4987 (N_4987,N_4749,N_4608);
or U4988 (N_4988,N_4625,N_4690);
xor U4989 (N_4989,N_4778,N_4790);
xnor U4990 (N_4990,N_4619,N_4699);
or U4991 (N_4991,N_4673,N_4688);
nor U4992 (N_4992,N_4660,N_4784);
xor U4993 (N_4993,N_4788,N_4760);
and U4994 (N_4994,N_4626,N_4628);
xor U4995 (N_4995,N_4734,N_4693);
nand U4996 (N_4996,N_4626,N_4670);
xnor U4997 (N_4997,N_4738,N_4678);
nor U4998 (N_4998,N_4640,N_4774);
nor U4999 (N_4999,N_4681,N_4669);
nor U5000 (N_5000,N_4891,N_4809);
xnor U5001 (N_5001,N_4877,N_4912);
and U5002 (N_5002,N_4827,N_4951);
nor U5003 (N_5003,N_4844,N_4833);
or U5004 (N_5004,N_4954,N_4848);
and U5005 (N_5005,N_4858,N_4886);
and U5006 (N_5006,N_4871,N_4842);
and U5007 (N_5007,N_4883,N_4958);
or U5008 (N_5008,N_4935,N_4806);
nor U5009 (N_5009,N_4804,N_4860);
nand U5010 (N_5010,N_4926,N_4993);
nor U5011 (N_5011,N_4838,N_4850);
nor U5012 (N_5012,N_4929,N_4965);
nand U5013 (N_5013,N_4879,N_4889);
nand U5014 (N_5014,N_4897,N_4953);
and U5015 (N_5015,N_4909,N_4852);
or U5016 (N_5016,N_4825,N_4876);
or U5017 (N_5017,N_4990,N_4800);
or U5018 (N_5018,N_4963,N_4836);
nor U5019 (N_5019,N_4974,N_4944);
or U5020 (N_5020,N_4859,N_4808);
and U5021 (N_5021,N_4816,N_4950);
xnor U5022 (N_5022,N_4835,N_4843);
or U5023 (N_5023,N_4933,N_4872);
or U5024 (N_5024,N_4811,N_4986);
and U5025 (N_5025,N_4875,N_4815);
xor U5026 (N_5026,N_4854,N_4878);
xnor U5027 (N_5027,N_4861,N_4928);
nand U5028 (N_5028,N_4812,N_4964);
xnor U5029 (N_5029,N_4866,N_4801);
or U5030 (N_5030,N_4830,N_4895);
and U5031 (N_5031,N_4985,N_4952);
or U5032 (N_5032,N_4956,N_4810);
xor U5033 (N_5033,N_4864,N_4969);
nor U5034 (N_5034,N_4826,N_4820);
xnor U5035 (N_5035,N_4994,N_4885);
nand U5036 (N_5036,N_4960,N_4847);
and U5037 (N_5037,N_4803,N_4892);
nand U5038 (N_5038,N_4906,N_4888);
xnor U5039 (N_5039,N_4957,N_4919);
or U5040 (N_5040,N_4831,N_4939);
xnor U5041 (N_5041,N_4938,N_4870);
and U5042 (N_5042,N_4855,N_4961);
and U5043 (N_5043,N_4997,N_4902);
nor U5044 (N_5044,N_4977,N_4999);
xnor U5045 (N_5045,N_4884,N_4840);
or U5046 (N_5046,N_4887,N_4893);
xnor U5047 (N_5047,N_4823,N_4874);
or U5048 (N_5048,N_4923,N_4834);
and U5049 (N_5049,N_4862,N_4959);
nor U5050 (N_5050,N_4813,N_4921);
nor U5051 (N_5051,N_4970,N_4925);
or U5052 (N_5052,N_4980,N_4818);
nand U5053 (N_5053,N_4942,N_4821);
or U5054 (N_5054,N_4948,N_4920);
and U5055 (N_5055,N_4996,N_4868);
xor U5056 (N_5056,N_4962,N_4863);
nand U5057 (N_5057,N_4901,N_4988);
and U5058 (N_5058,N_4880,N_4869);
xor U5059 (N_5059,N_4890,N_4903);
nand U5060 (N_5060,N_4898,N_4992);
nor U5061 (N_5061,N_4849,N_4937);
nor U5062 (N_5062,N_4913,N_4998);
nor U5063 (N_5063,N_4976,N_4851);
and U5064 (N_5064,N_4949,N_4932);
nor U5065 (N_5065,N_4873,N_4822);
nor U5066 (N_5066,N_4845,N_4911);
xor U5067 (N_5067,N_4967,N_4908);
or U5068 (N_5068,N_4896,N_4857);
or U5069 (N_5069,N_4907,N_4979);
and U5070 (N_5070,N_4915,N_4805);
nor U5071 (N_5071,N_4922,N_4941);
or U5072 (N_5072,N_4945,N_4991);
xnor U5073 (N_5073,N_4802,N_4807);
nor U5074 (N_5074,N_4828,N_4899);
and U5075 (N_5075,N_4978,N_4966);
and U5076 (N_5076,N_4934,N_4927);
nand U5077 (N_5077,N_4841,N_4824);
nor U5078 (N_5078,N_4981,N_4910);
nand U5079 (N_5079,N_4856,N_4817);
xor U5080 (N_5080,N_4881,N_4955);
or U5081 (N_5081,N_4904,N_4914);
nand U5082 (N_5082,N_4853,N_4867);
xor U5083 (N_5083,N_4829,N_4865);
and U5084 (N_5084,N_4984,N_4973);
nand U5085 (N_5085,N_4819,N_4989);
and U5086 (N_5086,N_4936,N_4900);
nor U5087 (N_5087,N_4943,N_4987);
or U5088 (N_5088,N_4814,N_4916);
or U5089 (N_5089,N_4968,N_4972);
xor U5090 (N_5090,N_4982,N_4846);
xnor U5091 (N_5091,N_4946,N_4947);
xor U5092 (N_5092,N_4940,N_4931);
or U5093 (N_5093,N_4839,N_4930);
and U5094 (N_5094,N_4918,N_4995);
and U5095 (N_5095,N_4894,N_4983);
nor U5096 (N_5096,N_4837,N_4832);
nor U5097 (N_5097,N_4905,N_4924);
or U5098 (N_5098,N_4917,N_4882);
and U5099 (N_5099,N_4971,N_4975);
and U5100 (N_5100,N_4979,N_4989);
xnor U5101 (N_5101,N_4832,N_4922);
nor U5102 (N_5102,N_4974,N_4942);
xnor U5103 (N_5103,N_4824,N_4819);
or U5104 (N_5104,N_4812,N_4953);
or U5105 (N_5105,N_4961,N_4829);
xor U5106 (N_5106,N_4867,N_4994);
nand U5107 (N_5107,N_4926,N_4919);
or U5108 (N_5108,N_4892,N_4819);
xor U5109 (N_5109,N_4812,N_4921);
xor U5110 (N_5110,N_4978,N_4920);
or U5111 (N_5111,N_4852,N_4972);
xnor U5112 (N_5112,N_4888,N_4864);
or U5113 (N_5113,N_4887,N_4906);
xnor U5114 (N_5114,N_4947,N_4909);
xnor U5115 (N_5115,N_4929,N_4904);
nand U5116 (N_5116,N_4964,N_4874);
and U5117 (N_5117,N_4967,N_4839);
or U5118 (N_5118,N_4934,N_4963);
xor U5119 (N_5119,N_4925,N_4879);
and U5120 (N_5120,N_4934,N_4877);
xnor U5121 (N_5121,N_4946,N_4820);
or U5122 (N_5122,N_4967,N_4988);
nand U5123 (N_5123,N_4900,N_4896);
or U5124 (N_5124,N_4878,N_4831);
or U5125 (N_5125,N_4932,N_4805);
nor U5126 (N_5126,N_4829,N_4970);
and U5127 (N_5127,N_4943,N_4885);
nor U5128 (N_5128,N_4936,N_4825);
xor U5129 (N_5129,N_4886,N_4996);
or U5130 (N_5130,N_4808,N_4887);
nor U5131 (N_5131,N_4972,N_4821);
xnor U5132 (N_5132,N_4891,N_4928);
nand U5133 (N_5133,N_4950,N_4818);
nand U5134 (N_5134,N_4800,N_4956);
nor U5135 (N_5135,N_4955,N_4827);
nor U5136 (N_5136,N_4872,N_4816);
nand U5137 (N_5137,N_4809,N_4855);
or U5138 (N_5138,N_4956,N_4817);
nand U5139 (N_5139,N_4993,N_4853);
xor U5140 (N_5140,N_4831,N_4819);
xnor U5141 (N_5141,N_4914,N_4864);
nand U5142 (N_5142,N_4837,N_4842);
nand U5143 (N_5143,N_4863,N_4953);
nand U5144 (N_5144,N_4937,N_4826);
xor U5145 (N_5145,N_4831,N_4841);
nand U5146 (N_5146,N_4913,N_4889);
and U5147 (N_5147,N_4851,N_4921);
or U5148 (N_5148,N_4986,N_4926);
xnor U5149 (N_5149,N_4966,N_4831);
nand U5150 (N_5150,N_4994,N_4957);
and U5151 (N_5151,N_4850,N_4980);
nand U5152 (N_5152,N_4838,N_4981);
and U5153 (N_5153,N_4888,N_4984);
nor U5154 (N_5154,N_4825,N_4881);
xnor U5155 (N_5155,N_4954,N_4853);
xnor U5156 (N_5156,N_4954,N_4884);
or U5157 (N_5157,N_4939,N_4979);
or U5158 (N_5158,N_4889,N_4900);
nor U5159 (N_5159,N_4971,N_4909);
or U5160 (N_5160,N_4906,N_4978);
nand U5161 (N_5161,N_4910,N_4953);
nor U5162 (N_5162,N_4965,N_4857);
nand U5163 (N_5163,N_4969,N_4822);
xnor U5164 (N_5164,N_4936,N_4928);
nor U5165 (N_5165,N_4892,N_4994);
nand U5166 (N_5166,N_4943,N_4815);
nand U5167 (N_5167,N_4816,N_4871);
and U5168 (N_5168,N_4829,N_4934);
and U5169 (N_5169,N_4878,N_4913);
and U5170 (N_5170,N_4929,N_4835);
xnor U5171 (N_5171,N_4830,N_4967);
xor U5172 (N_5172,N_4993,N_4850);
or U5173 (N_5173,N_4909,N_4930);
xnor U5174 (N_5174,N_4987,N_4975);
and U5175 (N_5175,N_4951,N_4826);
and U5176 (N_5176,N_4860,N_4918);
and U5177 (N_5177,N_4847,N_4954);
xnor U5178 (N_5178,N_4937,N_4888);
xnor U5179 (N_5179,N_4901,N_4870);
xor U5180 (N_5180,N_4988,N_4958);
xnor U5181 (N_5181,N_4988,N_4882);
or U5182 (N_5182,N_4883,N_4848);
nand U5183 (N_5183,N_4919,N_4955);
nor U5184 (N_5184,N_4807,N_4854);
or U5185 (N_5185,N_4928,N_4818);
xor U5186 (N_5186,N_4963,N_4819);
and U5187 (N_5187,N_4832,N_4951);
xnor U5188 (N_5188,N_4991,N_4811);
and U5189 (N_5189,N_4984,N_4834);
nor U5190 (N_5190,N_4856,N_4963);
and U5191 (N_5191,N_4879,N_4995);
nand U5192 (N_5192,N_4859,N_4999);
or U5193 (N_5193,N_4978,N_4958);
xor U5194 (N_5194,N_4878,N_4861);
or U5195 (N_5195,N_4925,N_4815);
or U5196 (N_5196,N_4984,N_4983);
and U5197 (N_5197,N_4902,N_4883);
nor U5198 (N_5198,N_4993,N_4895);
or U5199 (N_5199,N_4927,N_4971);
xor U5200 (N_5200,N_5135,N_5164);
nor U5201 (N_5201,N_5064,N_5020);
nor U5202 (N_5202,N_5075,N_5196);
nand U5203 (N_5203,N_5179,N_5198);
and U5204 (N_5204,N_5077,N_5141);
xor U5205 (N_5205,N_5058,N_5142);
nor U5206 (N_5206,N_5188,N_5004);
nor U5207 (N_5207,N_5091,N_5008);
xor U5208 (N_5208,N_5090,N_5013);
nor U5209 (N_5209,N_5103,N_5043);
nor U5210 (N_5210,N_5134,N_5145);
xnor U5211 (N_5211,N_5026,N_5067);
xnor U5212 (N_5212,N_5060,N_5106);
nor U5213 (N_5213,N_5037,N_5139);
xnor U5214 (N_5214,N_5088,N_5187);
xor U5215 (N_5215,N_5017,N_5158);
nand U5216 (N_5216,N_5167,N_5076);
and U5217 (N_5217,N_5030,N_5149);
and U5218 (N_5218,N_5104,N_5194);
xnor U5219 (N_5219,N_5022,N_5125);
nor U5220 (N_5220,N_5178,N_5101);
xor U5221 (N_5221,N_5019,N_5078);
nor U5222 (N_5222,N_5097,N_5162);
nand U5223 (N_5223,N_5113,N_5137);
nor U5224 (N_5224,N_5074,N_5199);
and U5225 (N_5225,N_5082,N_5025);
and U5226 (N_5226,N_5061,N_5140);
xor U5227 (N_5227,N_5131,N_5041);
nor U5228 (N_5228,N_5068,N_5072);
xnor U5229 (N_5229,N_5001,N_5053);
xnor U5230 (N_5230,N_5089,N_5123);
xnor U5231 (N_5231,N_5007,N_5021);
xnor U5232 (N_5232,N_5024,N_5111);
or U5233 (N_5233,N_5011,N_5154);
nor U5234 (N_5234,N_5130,N_5047);
nand U5235 (N_5235,N_5031,N_5120);
or U5236 (N_5236,N_5143,N_5056);
nor U5237 (N_5237,N_5049,N_5052);
xnor U5238 (N_5238,N_5093,N_5040);
or U5239 (N_5239,N_5159,N_5084);
nor U5240 (N_5240,N_5034,N_5127);
nand U5241 (N_5241,N_5118,N_5085);
nand U5242 (N_5242,N_5071,N_5027);
nor U5243 (N_5243,N_5128,N_5109);
nor U5244 (N_5244,N_5044,N_5192);
or U5245 (N_5245,N_5069,N_5108);
nand U5246 (N_5246,N_5114,N_5045);
nand U5247 (N_5247,N_5197,N_5018);
or U5248 (N_5248,N_5136,N_5148);
nor U5249 (N_5249,N_5156,N_5023);
nor U5250 (N_5250,N_5070,N_5033);
and U5251 (N_5251,N_5099,N_5190);
or U5252 (N_5252,N_5012,N_5079);
nor U5253 (N_5253,N_5092,N_5186);
and U5254 (N_5254,N_5124,N_5121);
nand U5255 (N_5255,N_5193,N_5096);
nand U5256 (N_5256,N_5161,N_5029);
or U5257 (N_5257,N_5174,N_5042);
or U5258 (N_5258,N_5151,N_5003);
xor U5259 (N_5259,N_5132,N_5184);
and U5260 (N_5260,N_5080,N_5173);
or U5261 (N_5261,N_5165,N_5098);
nor U5262 (N_5262,N_5095,N_5175);
or U5263 (N_5263,N_5189,N_5176);
nor U5264 (N_5264,N_5063,N_5065);
or U5265 (N_5265,N_5153,N_5005);
or U5266 (N_5266,N_5046,N_5144);
xnor U5267 (N_5267,N_5122,N_5002);
and U5268 (N_5268,N_5180,N_5038);
and U5269 (N_5269,N_5073,N_5087);
and U5270 (N_5270,N_5000,N_5166);
nor U5271 (N_5271,N_5185,N_5050);
nor U5272 (N_5272,N_5182,N_5171);
xor U5273 (N_5273,N_5035,N_5009);
nor U5274 (N_5274,N_5015,N_5146);
nand U5275 (N_5275,N_5183,N_5055);
nor U5276 (N_5276,N_5094,N_5032);
and U5277 (N_5277,N_5150,N_5152);
or U5278 (N_5278,N_5119,N_5006);
nand U5279 (N_5279,N_5191,N_5016);
and U5280 (N_5280,N_5014,N_5110);
or U5281 (N_5281,N_5138,N_5181);
or U5282 (N_5282,N_5107,N_5129);
or U5283 (N_5283,N_5133,N_5066);
nor U5284 (N_5284,N_5169,N_5062);
and U5285 (N_5285,N_5195,N_5054);
nand U5286 (N_5286,N_5010,N_5100);
nor U5287 (N_5287,N_5172,N_5115);
nor U5288 (N_5288,N_5168,N_5039);
and U5289 (N_5289,N_5117,N_5147);
xor U5290 (N_5290,N_5102,N_5086);
and U5291 (N_5291,N_5177,N_5059);
xnor U5292 (N_5292,N_5157,N_5048);
or U5293 (N_5293,N_5160,N_5155);
or U5294 (N_5294,N_5083,N_5051);
or U5295 (N_5295,N_5170,N_5105);
and U5296 (N_5296,N_5163,N_5112);
xor U5297 (N_5297,N_5036,N_5057);
nand U5298 (N_5298,N_5116,N_5126);
or U5299 (N_5299,N_5028,N_5081);
nand U5300 (N_5300,N_5185,N_5173);
and U5301 (N_5301,N_5099,N_5042);
or U5302 (N_5302,N_5179,N_5109);
xor U5303 (N_5303,N_5163,N_5152);
xnor U5304 (N_5304,N_5109,N_5198);
nand U5305 (N_5305,N_5001,N_5137);
nor U5306 (N_5306,N_5169,N_5034);
and U5307 (N_5307,N_5131,N_5021);
and U5308 (N_5308,N_5105,N_5050);
nor U5309 (N_5309,N_5056,N_5036);
or U5310 (N_5310,N_5022,N_5008);
nor U5311 (N_5311,N_5066,N_5015);
and U5312 (N_5312,N_5106,N_5132);
nor U5313 (N_5313,N_5151,N_5125);
and U5314 (N_5314,N_5079,N_5161);
xor U5315 (N_5315,N_5185,N_5132);
and U5316 (N_5316,N_5056,N_5004);
nand U5317 (N_5317,N_5085,N_5134);
nand U5318 (N_5318,N_5029,N_5131);
nand U5319 (N_5319,N_5075,N_5043);
or U5320 (N_5320,N_5035,N_5147);
nand U5321 (N_5321,N_5189,N_5043);
or U5322 (N_5322,N_5195,N_5045);
nand U5323 (N_5323,N_5039,N_5051);
nand U5324 (N_5324,N_5179,N_5140);
or U5325 (N_5325,N_5138,N_5172);
xnor U5326 (N_5326,N_5066,N_5121);
or U5327 (N_5327,N_5001,N_5094);
nor U5328 (N_5328,N_5055,N_5192);
and U5329 (N_5329,N_5097,N_5194);
or U5330 (N_5330,N_5038,N_5111);
xor U5331 (N_5331,N_5169,N_5167);
and U5332 (N_5332,N_5191,N_5057);
and U5333 (N_5333,N_5170,N_5048);
xnor U5334 (N_5334,N_5011,N_5023);
and U5335 (N_5335,N_5152,N_5101);
and U5336 (N_5336,N_5147,N_5087);
and U5337 (N_5337,N_5153,N_5129);
xor U5338 (N_5338,N_5053,N_5000);
nor U5339 (N_5339,N_5152,N_5184);
or U5340 (N_5340,N_5149,N_5156);
or U5341 (N_5341,N_5073,N_5118);
or U5342 (N_5342,N_5006,N_5185);
nand U5343 (N_5343,N_5181,N_5149);
nand U5344 (N_5344,N_5072,N_5086);
and U5345 (N_5345,N_5193,N_5057);
nor U5346 (N_5346,N_5128,N_5063);
xnor U5347 (N_5347,N_5145,N_5164);
xnor U5348 (N_5348,N_5012,N_5072);
and U5349 (N_5349,N_5019,N_5168);
xor U5350 (N_5350,N_5029,N_5058);
and U5351 (N_5351,N_5064,N_5071);
and U5352 (N_5352,N_5122,N_5121);
or U5353 (N_5353,N_5014,N_5102);
nand U5354 (N_5354,N_5127,N_5079);
nor U5355 (N_5355,N_5008,N_5192);
nor U5356 (N_5356,N_5079,N_5105);
nand U5357 (N_5357,N_5162,N_5047);
and U5358 (N_5358,N_5074,N_5001);
and U5359 (N_5359,N_5025,N_5102);
xor U5360 (N_5360,N_5049,N_5158);
or U5361 (N_5361,N_5054,N_5151);
nor U5362 (N_5362,N_5191,N_5096);
and U5363 (N_5363,N_5003,N_5120);
nor U5364 (N_5364,N_5137,N_5006);
nand U5365 (N_5365,N_5196,N_5072);
or U5366 (N_5366,N_5144,N_5019);
xor U5367 (N_5367,N_5197,N_5191);
nand U5368 (N_5368,N_5115,N_5029);
nand U5369 (N_5369,N_5072,N_5076);
or U5370 (N_5370,N_5102,N_5002);
nor U5371 (N_5371,N_5103,N_5153);
and U5372 (N_5372,N_5013,N_5157);
or U5373 (N_5373,N_5164,N_5151);
and U5374 (N_5374,N_5100,N_5146);
xnor U5375 (N_5375,N_5190,N_5192);
nor U5376 (N_5376,N_5121,N_5076);
nor U5377 (N_5377,N_5032,N_5118);
xnor U5378 (N_5378,N_5064,N_5161);
and U5379 (N_5379,N_5014,N_5036);
or U5380 (N_5380,N_5067,N_5171);
xor U5381 (N_5381,N_5186,N_5199);
or U5382 (N_5382,N_5161,N_5091);
or U5383 (N_5383,N_5141,N_5112);
or U5384 (N_5384,N_5190,N_5023);
nor U5385 (N_5385,N_5028,N_5080);
nand U5386 (N_5386,N_5176,N_5096);
nor U5387 (N_5387,N_5109,N_5105);
and U5388 (N_5388,N_5076,N_5065);
and U5389 (N_5389,N_5006,N_5087);
nor U5390 (N_5390,N_5169,N_5072);
and U5391 (N_5391,N_5138,N_5022);
xnor U5392 (N_5392,N_5086,N_5061);
or U5393 (N_5393,N_5101,N_5064);
or U5394 (N_5394,N_5089,N_5181);
nand U5395 (N_5395,N_5081,N_5182);
nand U5396 (N_5396,N_5060,N_5149);
xnor U5397 (N_5397,N_5171,N_5180);
nor U5398 (N_5398,N_5157,N_5084);
or U5399 (N_5399,N_5077,N_5060);
and U5400 (N_5400,N_5223,N_5225);
nor U5401 (N_5401,N_5222,N_5205);
xnor U5402 (N_5402,N_5287,N_5296);
nand U5403 (N_5403,N_5389,N_5221);
nand U5404 (N_5404,N_5201,N_5206);
or U5405 (N_5405,N_5233,N_5254);
or U5406 (N_5406,N_5327,N_5330);
or U5407 (N_5407,N_5209,N_5391);
nand U5408 (N_5408,N_5299,N_5235);
nor U5409 (N_5409,N_5231,N_5390);
nor U5410 (N_5410,N_5349,N_5288);
nand U5411 (N_5411,N_5291,N_5274);
nor U5412 (N_5412,N_5310,N_5289);
nand U5413 (N_5413,N_5252,N_5256);
and U5414 (N_5414,N_5344,N_5361);
xnor U5415 (N_5415,N_5238,N_5202);
and U5416 (N_5416,N_5338,N_5328);
or U5417 (N_5417,N_5309,N_5297);
and U5418 (N_5418,N_5216,N_5226);
nand U5419 (N_5419,N_5373,N_5399);
nor U5420 (N_5420,N_5304,N_5245);
nor U5421 (N_5421,N_5294,N_5323);
or U5422 (N_5422,N_5230,N_5321);
nand U5423 (N_5423,N_5394,N_5302);
xnor U5424 (N_5424,N_5290,N_5237);
xor U5425 (N_5425,N_5278,N_5265);
nor U5426 (N_5426,N_5397,N_5312);
or U5427 (N_5427,N_5259,N_5261);
xnor U5428 (N_5428,N_5364,N_5282);
xnor U5429 (N_5429,N_5374,N_5352);
nand U5430 (N_5430,N_5375,N_5348);
nand U5431 (N_5431,N_5317,N_5212);
or U5432 (N_5432,N_5305,N_5244);
or U5433 (N_5433,N_5204,N_5396);
or U5434 (N_5434,N_5283,N_5377);
nor U5435 (N_5435,N_5332,N_5350);
nor U5436 (N_5436,N_5342,N_5219);
and U5437 (N_5437,N_5379,N_5251);
and U5438 (N_5438,N_5372,N_5276);
nand U5439 (N_5439,N_5293,N_5228);
xor U5440 (N_5440,N_5311,N_5346);
nor U5441 (N_5441,N_5383,N_5232);
nand U5442 (N_5442,N_5218,N_5203);
nor U5443 (N_5443,N_5266,N_5267);
or U5444 (N_5444,N_5368,N_5308);
xnor U5445 (N_5445,N_5331,N_5355);
xnor U5446 (N_5446,N_5365,N_5339);
xor U5447 (N_5447,N_5246,N_5381);
nand U5448 (N_5448,N_5363,N_5285);
nor U5449 (N_5449,N_5281,N_5306);
xor U5450 (N_5450,N_5382,N_5277);
or U5451 (N_5451,N_5329,N_5320);
and U5452 (N_5452,N_5298,N_5211);
nand U5453 (N_5453,N_5217,N_5270);
nor U5454 (N_5454,N_5334,N_5242);
or U5455 (N_5455,N_5371,N_5250);
and U5456 (N_5456,N_5347,N_5393);
or U5457 (N_5457,N_5395,N_5257);
nand U5458 (N_5458,N_5241,N_5325);
nand U5459 (N_5459,N_5253,N_5369);
nor U5460 (N_5460,N_5263,N_5353);
nor U5461 (N_5461,N_5258,N_5326);
xnor U5462 (N_5462,N_5380,N_5300);
nor U5463 (N_5463,N_5248,N_5280);
nor U5464 (N_5464,N_5301,N_5319);
and U5465 (N_5465,N_5224,N_5208);
or U5466 (N_5466,N_5357,N_5275);
nand U5467 (N_5467,N_5234,N_5284);
and U5468 (N_5468,N_5214,N_5354);
and U5469 (N_5469,N_5247,N_5240);
nor U5470 (N_5470,N_5316,N_5360);
or U5471 (N_5471,N_5273,N_5269);
nand U5472 (N_5472,N_5335,N_5243);
or U5473 (N_5473,N_5398,N_5314);
or U5474 (N_5474,N_5264,N_5336);
nand U5475 (N_5475,N_5236,N_5286);
xnor U5476 (N_5476,N_5370,N_5313);
or U5477 (N_5477,N_5324,N_5272);
xor U5478 (N_5478,N_5359,N_5322);
or U5479 (N_5479,N_5387,N_5213);
nand U5480 (N_5480,N_5366,N_5333);
and U5481 (N_5481,N_5385,N_5279);
nor U5482 (N_5482,N_5367,N_5337);
and U5483 (N_5483,N_5351,N_5220);
or U5484 (N_5484,N_5229,N_5386);
nor U5485 (N_5485,N_5356,N_5239);
xor U5486 (N_5486,N_5268,N_5255);
or U5487 (N_5487,N_5378,N_5200);
or U5488 (N_5488,N_5215,N_5388);
nand U5489 (N_5489,N_5295,N_5318);
xnor U5490 (N_5490,N_5358,N_5271);
nand U5491 (N_5491,N_5362,N_5343);
and U5492 (N_5492,N_5392,N_5292);
nor U5493 (N_5493,N_5227,N_5345);
or U5494 (N_5494,N_5307,N_5376);
nor U5495 (N_5495,N_5340,N_5384);
and U5496 (N_5496,N_5207,N_5262);
xnor U5497 (N_5497,N_5315,N_5341);
or U5498 (N_5498,N_5249,N_5303);
and U5499 (N_5499,N_5260,N_5210);
or U5500 (N_5500,N_5356,N_5277);
nand U5501 (N_5501,N_5244,N_5266);
or U5502 (N_5502,N_5238,N_5257);
or U5503 (N_5503,N_5292,N_5235);
and U5504 (N_5504,N_5262,N_5224);
nand U5505 (N_5505,N_5355,N_5359);
and U5506 (N_5506,N_5203,N_5371);
and U5507 (N_5507,N_5345,N_5320);
xor U5508 (N_5508,N_5326,N_5200);
nor U5509 (N_5509,N_5317,N_5307);
nand U5510 (N_5510,N_5257,N_5218);
nor U5511 (N_5511,N_5224,N_5211);
or U5512 (N_5512,N_5237,N_5260);
nand U5513 (N_5513,N_5230,N_5315);
or U5514 (N_5514,N_5339,N_5258);
nand U5515 (N_5515,N_5366,N_5254);
nor U5516 (N_5516,N_5300,N_5216);
or U5517 (N_5517,N_5369,N_5304);
xor U5518 (N_5518,N_5283,N_5239);
nand U5519 (N_5519,N_5242,N_5350);
or U5520 (N_5520,N_5327,N_5398);
and U5521 (N_5521,N_5216,N_5273);
nand U5522 (N_5522,N_5325,N_5275);
nand U5523 (N_5523,N_5306,N_5339);
nand U5524 (N_5524,N_5378,N_5266);
and U5525 (N_5525,N_5249,N_5246);
and U5526 (N_5526,N_5303,N_5248);
xnor U5527 (N_5527,N_5244,N_5282);
nand U5528 (N_5528,N_5314,N_5332);
or U5529 (N_5529,N_5280,N_5391);
or U5530 (N_5530,N_5243,N_5366);
and U5531 (N_5531,N_5377,N_5328);
nand U5532 (N_5532,N_5346,N_5370);
xnor U5533 (N_5533,N_5348,N_5323);
nand U5534 (N_5534,N_5374,N_5219);
and U5535 (N_5535,N_5282,N_5356);
and U5536 (N_5536,N_5369,N_5244);
nor U5537 (N_5537,N_5227,N_5294);
nor U5538 (N_5538,N_5224,N_5316);
and U5539 (N_5539,N_5363,N_5326);
or U5540 (N_5540,N_5227,N_5337);
nand U5541 (N_5541,N_5376,N_5333);
and U5542 (N_5542,N_5392,N_5226);
xnor U5543 (N_5543,N_5357,N_5288);
nand U5544 (N_5544,N_5380,N_5348);
nor U5545 (N_5545,N_5268,N_5223);
or U5546 (N_5546,N_5271,N_5297);
and U5547 (N_5547,N_5272,N_5341);
nor U5548 (N_5548,N_5324,N_5397);
and U5549 (N_5549,N_5274,N_5328);
or U5550 (N_5550,N_5217,N_5257);
nor U5551 (N_5551,N_5218,N_5295);
xor U5552 (N_5552,N_5320,N_5272);
and U5553 (N_5553,N_5364,N_5387);
or U5554 (N_5554,N_5291,N_5368);
or U5555 (N_5555,N_5320,N_5211);
or U5556 (N_5556,N_5269,N_5382);
or U5557 (N_5557,N_5339,N_5224);
and U5558 (N_5558,N_5387,N_5245);
nor U5559 (N_5559,N_5225,N_5335);
and U5560 (N_5560,N_5222,N_5319);
nand U5561 (N_5561,N_5205,N_5357);
and U5562 (N_5562,N_5206,N_5293);
or U5563 (N_5563,N_5205,N_5239);
nand U5564 (N_5564,N_5353,N_5340);
and U5565 (N_5565,N_5282,N_5390);
and U5566 (N_5566,N_5310,N_5381);
or U5567 (N_5567,N_5388,N_5205);
nor U5568 (N_5568,N_5311,N_5347);
nor U5569 (N_5569,N_5268,N_5208);
nor U5570 (N_5570,N_5398,N_5365);
and U5571 (N_5571,N_5264,N_5283);
and U5572 (N_5572,N_5203,N_5315);
and U5573 (N_5573,N_5292,N_5274);
xor U5574 (N_5574,N_5331,N_5295);
nand U5575 (N_5575,N_5375,N_5245);
and U5576 (N_5576,N_5294,N_5361);
xnor U5577 (N_5577,N_5247,N_5328);
and U5578 (N_5578,N_5229,N_5247);
nor U5579 (N_5579,N_5219,N_5360);
xor U5580 (N_5580,N_5215,N_5229);
nand U5581 (N_5581,N_5234,N_5211);
nor U5582 (N_5582,N_5205,N_5315);
and U5583 (N_5583,N_5335,N_5250);
nand U5584 (N_5584,N_5354,N_5228);
and U5585 (N_5585,N_5313,N_5215);
or U5586 (N_5586,N_5206,N_5291);
nor U5587 (N_5587,N_5270,N_5200);
or U5588 (N_5588,N_5376,N_5276);
xor U5589 (N_5589,N_5394,N_5241);
xor U5590 (N_5590,N_5236,N_5284);
nor U5591 (N_5591,N_5383,N_5241);
and U5592 (N_5592,N_5360,N_5285);
nand U5593 (N_5593,N_5274,N_5308);
or U5594 (N_5594,N_5312,N_5362);
nor U5595 (N_5595,N_5330,N_5235);
nor U5596 (N_5596,N_5208,N_5306);
xor U5597 (N_5597,N_5343,N_5271);
xnor U5598 (N_5598,N_5202,N_5280);
or U5599 (N_5599,N_5375,N_5231);
and U5600 (N_5600,N_5468,N_5486);
and U5601 (N_5601,N_5418,N_5440);
nand U5602 (N_5602,N_5548,N_5515);
or U5603 (N_5603,N_5441,N_5439);
or U5604 (N_5604,N_5442,N_5529);
nor U5605 (N_5605,N_5541,N_5527);
nand U5606 (N_5606,N_5554,N_5511);
or U5607 (N_5607,N_5449,N_5482);
or U5608 (N_5608,N_5487,N_5467);
and U5609 (N_5609,N_5498,N_5517);
or U5610 (N_5610,N_5577,N_5438);
xor U5611 (N_5611,N_5443,N_5450);
and U5612 (N_5612,N_5580,N_5532);
and U5613 (N_5613,N_5568,N_5586);
nor U5614 (N_5614,N_5534,N_5563);
nand U5615 (N_5615,N_5574,N_5473);
xnor U5616 (N_5616,N_5564,N_5459);
and U5617 (N_5617,N_5591,N_5552);
nor U5618 (N_5618,N_5412,N_5537);
nor U5619 (N_5619,N_5583,N_5495);
xnor U5620 (N_5620,N_5525,N_5557);
and U5621 (N_5621,N_5451,N_5488);
nor U5622 (N_5622,N_5429,N_5403);
and U5623 (N_5623,N_5445,N_5544);
nand U5624 (N_5624,N_5526,N_5565);
nor U5625 (N_5625,N_5542,N_5481);
and U5626 (N_5626,N_5535,N_5489);
or U5627 (N_5627,N_5472,N_5444);
nand U5628 (N_5628,N_5431,N_5496);
and U5629 (N_5629,N_5503,N_5452);
or U5630 (N_5630,N_5499,N_5436);
nand U5631 (N_5631,N_5420,N_5522);
or U5632 (N_5632,N_5582,N_5536);
nor U5633 (N_5633,N_5528,N_5415);
xnor U5634 (N_5634,N_5424,N_5479);
or U5635 (N_5635,N_5587,N_5546);
xor U5636 (N_5636,N_5400,N_5520);
nor U5637 (N_5637,N_5593,N_5437);
nor U5638 (N_5638,N_5426,N_5455);
xor U5639 (N_5639,N_5549,N_5463);
nor U5640 (N_5640,N_5555,N_5456);
xor U5641 (N_5641,N_5471,N_5405);
nor U5642 (N_5642,N_5599,N_5490);
and U5643 (N_5643,N_5576,N_5572);
nor U5644 (N_5644,N_5447,N_5427);
nor U5645 (N_5645,N_5454,N_5598);
and U5646 (N_5646,N_5510,N_5474);
nor U5647 (N_5647,N_5457,N_5562);
nor U5648 (N_5648,N_5566,N_5446);
xnor U5649 (N_5649,N_5584,N_5417);
and U5650 (N_5650,N_5423,N_5575);
nand U5651 (N_5651,N_5458,N_5469);
and U5652 (N_5652,N_5500,N_5569);
and U5653 (N_5653,N_5408,N_5514);
and U5654 (N_5654,N_5533,N_5513);
nand U5655 (N_5655,N_5595,N_5590);
or U5656 (N_5656,N_5494,N_5462);
and U5657 (N_5657,N_5556,N_5540);
or U5658 (N_5658,N_5589,N_5461);
xnor U5659 (N_5659,N_5553,N_5509);
and U5660 (N_5660,N_5402,N_5521);
nor U5661 (N_5661,N_5570,N_5421);
and U5662 (N_5662,N_5428,N_5401);
xnor U5663 (N_5663,N_5413,N_5406);
nand U5664 (N_5664,N_5476,N_5508);
or U5665 (N_5665,N_5484,N_5519);
nand U5666 (N_5666,N_5573,N_5504);
nor U5667 (N_5667,N_5581,N_5594);
nor U5668 (N_5668,N_5571,N_5430);
or U5669 (N_5669,N_5560,N_5578);
and U5670 (N_5670,N_5466,N_5523);
and U5671 (N_5671,N_5547,N_5491);
or U5672 (N_5672,N_5518,N_5502);
nand U5673 (N_5673,N_5470,N_5512);
nor U5674 (N_5674,N_5433,N_5425);
nor U5675 (N_5675,N_5460,N_5539);
nand U5676 (N_5676,N_5465,N_5432);
or U5677 (N_5677,N_5493,N_5464);
and U5678 (N_5678,N_5448,N_5588);
and U5679 (N_5679,N_5411,N_5585);
nor U5680 (N_5680,N_5507,N_5478);
nor U5681 (N_5681,N_5409,N_5559);
nor U5682 (N_5682,N_5480,N_5545);
xor U5683 (N_5683,N_5551,N_5434);
nor U5684 (N_5684,N_5485,N_5530);
xor U5685 (N_5685,N_5501,N_5524);
nand U5686 (N_5686,N_5422,N_5597);
nand U5687 (N_5687,N_5543,N_5419);
or U5688 (N_5688,N_5506,N_5567);
or U5689 (N_5689,N_5477,N_5550);
nand U5690 (N_5690,N_5516,N_5538);
nand U5691 (N_5691,N_5505,N_5558);
xnor U5692 (N_5692,N_5414,N_5483);
and U5693 (N_5693,N_5453,N_5410);
or U5694 (N_5694,N_5475,N_5407);
or U5695 (N_5695,N_5435,N_5416);
xnor U5696 (N_5696,N_5492,N_5592);
nand U5697 (N_5697,N_5497,N_5561);
xor U5698 (N_5698,N_5579,N_5596);
or U5699 (N_5699,N_5531,N_5404);
and U5700 (N_5700,N_5559,N_5439);
nor U5701 (N_5701,N_5530,N_5537);
nand U5702 (N_5702,N_5523,N_5536);
and U5703 (N_5703,N_5550,N_5488);
or U5704 (N_5704,N_5462,N_5421);
xnor U5705 (N_5705,N_5562,N_5573);
or U5706 (N_5706,N_5409,N_5569);
xor U5707 (N_5707,N_5451,N_5490);
and U5708 (N_5708,N_5414,N_5481);
and U5709 (N_5709,N_5537,N_5575);
nand U5710 (N_5710,N_5595,N_5441);
nand U5711 (N_5711,N_5543,N_5544);
xor U5712 (N_5712,N_5509,N_5514);
nand U5713 (N_5713,N_5408,N_5405);
or U5714 (N_5714,N_5599,N_5459);
nand U5715 (N_5715,N_5489,N_5497);
or U5716 (N_5716,N_5587,N_5581);
nor U5717 (N_5717,N_5401,N_5515);
xnor U5718 (N_5718,N_5518,N_5456);
xnor U5719 (N_5719,N_5522,N_5537);
and U5720 (N_5720,N_5410,N_5583);
or U5721 (N_5721,N_5450,N_5448);
or U5722 (N_5722,N_5558,N_5544);
xor U5723 (N_5723,N_5481,N_5426);
nand U5724 (N_5724,N_5554,N_5535);
nor U5725 (N_5725,N_5464,N_5518);
and U5726 (N_5726,N_5537,N_5503);
or U5727 (N_5727,N_5415,N_5555);
and U5728 (N_5728,N_5415,N_5499);
and U5729 (N_5729,N_5426,N_5475);
xor U5730 (N_5730,N_5532,N_5539);
and U5731 (N_5731,N_5525,N_5402);
and U5732 (N_5732,N_5563,N_5455);
and U5733 (N_5733,N_5497,N_5595);
nor U5734 (N_5734,N_5464,N_5432);
xor U5735 (N_5735,N_5408,N_5598);
or U5736 (N_5736,N_5573,N_5526);
or U5737 (N_5737,N_5436,N_5498);
and U5738 (N_5738,N_5410,N_5474);
xnor U5739 (N_5739,N_5469,N_5550);
or U5740 (N_5740,N_5471,N_5455);
and U5741 (N_5741,N_5410,N_5482);
nand U5742 (N_5742,N_5442,N_5568);
or U5743 (N_5743,N_5591,N_5472);
or U5744 (N_5744,N_5419,N_5572);
xor U5745 (N_5745,N_5510,N_5537);
nand U5746 (N_5746,N_5453,N_5530);
and U5747 (N_5747,N_5409,N_5550);
and U5748 (N_5748,N_5529,N_5400);
nand U5749 (N_5749,N_5462,N_5474);
or U5750 (N_5750,N_5575,N_5567);
nand U5751 (N_5751,N_5458,N_5511);
nor U5752 (N_5752,N_5514,N_5489);
nand U5753 (N_5753,N_5554,N_5520);
or U5754 (N_5754,N_5429,N_5443);
xor U5755 (N_5755,N_5557,N_5496);
nand U5756 (N_5756,N_5411,N_5469);
nand U5757 (N_5757,N_5503,N_5532);
nand U5758 (N_5758,N_5558,N_5476);
and U5759 (N_5759,N_5569,N_5468);
and U5760 (N_5760,N_5419,N_5432);
nand U5761 (N_5761,N_5539,N_5475);
xor U5762 (N_5762,N_5526,N_5498);
and U5763 (N_5763,N_5460,N_5484);
and U5764 (N_5764,N_5516,N_5407);
and U5765 (N_5765,N_5476,N_5557);
and U5766 (N_5766,N_5555,N_5417);
nor U5767 (N_5767,N_5487,N_5466);
xnor U5768 (N_5768,N_5426,N_5458);
and U5769 (N_5769,N_5442,N_5567);
nand U5770 (N_5770,N_5579,N_5409);
and U5771 (N_5771,N_5490,N_5567);
or U5772 (N_5772,N_5452,N_5416);
or U5773 (N_5773,N_5566,N_5586);
and U5774 (N_5774,N_5525,N_5407);
and U5775 (N_5775,N_5417,N_5572);
nand U5776 (N_5776,N_5435,N_5519);
nand U5777 (N_5777,N_5487,N_5534);
or U5778 (N_5778,N_5443,N_5409);
nand U5779 (N_5779,N_5518,N_5417);
and U5780 (N_5780,N_5576,N_5594);
nand U5781 (N_5781,N_5468,N_5414);
xnor U5782 (N_5782,N_5400,N_5467);
and U5783 (N_5783,N_5467,N_5406);
or U5784 (N_5784,N_5433,N_5409);
and U5785 (N_5785,N_5469,N_5502);
nor U5786 (N_5786,N_5407,N_5479);
xnor U5787 (N_5787,N_5444,N_5579);
and U5788 (N_5788,N_5537,N_5592);
and U5789 (N_5789,N_5596,N_5408);
nand U5790 (N_5790,N_5536,N_5537);
nand U5791 (N_5791,N_5564,N_5401);
nor U5792 (N_5792,N_5570,N_5469);
xor U5793 (N_5793,N_5539,N_5493);
nand U5794 (N_5794,N_5572,N_5533);
or U5795 (N_5795,N_5498,N_5521);
or U5796 (N_5796,N_5474,N_5452);
nand U5797 (N_5797,N_5504,N_5548);
nor U5798 (N_5798,N_5559,N_5428);
nand U5799 (N_5799,N_5421,N_5418);
nor U5800 (N_5800,N_5676,N_5694);
and U5801 (N_5801,N_5791,N_5734);
xor U5802 (N_5802,N_5765,N_5624);
nor U5803 (N_5803,N_5639,N_5682);
nand U5804 (N_5804,N_5784,N_5608);
and U5805 (N_5805,N_5645,N_5602);
nor U5806 (N_5806,N_5771,N_5697);
nand U5807 (N_5807,N_5668,N_5736);
or U5808 (N_5808,N_5640,N_5794);
xor U5809 (N_5809,N_5774,N_5610);
nand U5810 (N_5810,N_5604,N_5683);
or U5811 (N_5811,N_5621,N_5628);
and U5812 (N_5812,N_5790,N_5754);
and U5813 (N_5813,N_5696,N_5607);
nand U5814 (N_5814,N_5709,N_5631);
and U5815 (N_5815,N_5735,N_5693);
xor U5816 (N_5816,N_5678,N_5638);
nor U5817 (N_5817,N_5724,N_5740);
and U5818 (N_5818,N_5657,N_5633);
nand U5819 (N_5819,N_5727,N_5636);
xnor U5820 (N_5820,N_5691,N_5775);
or U5821 (N_5821,N_5711,N_5647);
nand U5822 (N_5822,N_5772,N_5706);
xor U5823 (N_5823,N_5689,N_5746);
nand U5824 (N_5824,N_5619,N_5778);
nor U5825 (N_5825,N_5725,N_5749);
and U5826 (N_5826,N_5672,N_5704);
nor U5827 (N_5827,N_5719,N_5798);
or U5828 (N_5828,N_5635,N_5732);
or U5829 (N_5829,N_5769,N_5674);
and U5830 (N_5830,N_5653,N_5605);
nand U5831 (N_5831,N_5649,N_5708);
nand U5832 (N_5832,N_5616,N_5690);
nand U5833 (N_5833,N_5726,N_5627);
or U5834 (N_5834,N_5644,N_5703);
and U5835 (N_5835,N_5779,N_5789);
and U5836 (N_5836,N_5656,N_5667);
nand U5837 (N_5837,N_5767,N_5687);
or U5838 (N_5838,N_5669,N_5731);
or U5839 (N_5839,N_5782,N_5629);
xor U5840 (N_5840,N_5614,N_5759);
xor U5841 (N_5841,N_5753,N_5751);
nor U5842 (N_5842,N_5646,N_5793);
nor U5843 (N_5843,N_5603,N_5673);
nand U5844 (N_5844,N_5768,N_5728);
or U5845 (N_5845,N_5617,N_5671);
and U5846 (N_5846,N_5660,N_5714);
or U5847 (N_5847,N_5651,N_5688);
or U5848 (N_5848,N_5670,N_5700);
or U5849 (N_5849,N_5684,N_5659);
and U5850 (N_5850,N_5623,N_5750);
xnor U5851 (N_5851,N_5757,N_5620);
nand U5852 (N_5852,N_5641,N_5622);
nor U5853 (N_5853,N_5763,N_5634);
and U5854 (N_5854,N_5630,N_5625);
nor U5855 (N_5855,N_5786,N_5783);
xor U5856 (N_5856,N_5797,N_5755);
and U5857 (N_5857,N_5681,N_5717);
nand U5858 (N_5858,N_5666,N_5730);
or U5859 (N_5859,N_5760,N_5748);
nor U5860 (N_5860,N_5761,N_5662);
nor U5861 (N_5861,N_5729,N_5716);
nor U5862 (N_5862,N_5737,N_5781);
xor U5863 (N_5863,N_5615,N_5770);
nor U5864 (N_5864,N_5648,N_5664);
or U5865 (N_5865,N_5692,N_5773);
nor U5866 (N_5866,N_5787,N_5720);
and U5867 (N_5867,N_5642,N_5695);
nor U5868 (N_5868,N_5702,N_5698);
xor U5869 (N_5869,N_5766,N_5710);
nor U5870 (N_5870,N_5762,N_5788);
xor U5871 (N_5871,N_5613,N_5758);
nand U5872 (N_5872,N_5744,N_5712);
xnor U5873 (N_5873,N_5685,N_5679);
nand U5874 (N_5874,N_5677,N_5699);
xnor U5875 (N_5875,N_5752,N_5675);
or U5876 (N_5876,N_5600,N_5643);
xnor U5877 (N_5877,N_5743,N_5721);
and U5878 (N_5878,N_5785,N_5652);
xor U5879 (N_5879,N_5738,N_5745);
xnor U5880 (N_5880,N_5780,N_5637);
nand U5881 (N_5881,N_5707,N_5609);
xor U5882 (N_5882,N_5655,N_5739);
nand U5883 (N_5883,N_5665,N_5733);
xor U5884 (N_5884,N_5723,N_5601);
nand U5885 (N_5885,N_5764,N_5606);
or U5886 (N_5886,N_5663,N_5799);
nor U5887 (N_5887,N_5618,N_5713);
or U5888 (N_5888,N_5792,N_5705);
or U5889 (N_5889,N_5777,N_5756);
and U5890 (N_5890,N_5747,N_5715);
or U5891 (N_5891,N_5795,N_5742);
nand U5892 (N_5892,N_5661,N_5776);
xor U5893 (N_5893,N_5612,N_5654);
nor U5894 (N_5894,N_5796,N_5632);
nor U5895 (N_5895,N_5650,N_5686);
xor U5896 (N_5896,N_5718,N_5626);
nand U5897 (N_5897,N_5658,N_5611);
nand U5898 (N_5898,N_5741,N_5680);
or U5899 (N_5899,N_5701,N_5722);
or U5900 (N_5900,N_5743,N_5775);
and U5901 (N_5901,N_5789,N_5690);
or U5902 (N_5902,N_5732,N_5708);
xnor U5903 (N_5903,N_5614,N_5640);
nand U5904 (N_5904,N_5666,N_5731);
nand U5905 (N_5905,N_5785,N_5761);
nand U5906 (N_5906,N_5623,N_5655);
and U5907 (N_5907,N_5763,N_5663);
nor U5908 (N_5908,N_5758,N_5626);
nand U5909 (N_5909,N_5683,N_5649);
nor U5910 (N_5910,N_5684,N_5791);
nor U5911 (N_5911,N_5685,N_5609);
nor U5912 (N_5912,N_5647,N_5694);
or U5913 (N_5913,N_5765,N_5652);
xnor U5914 (N_5914,N_5790,N_5605);
xor U5915 (N_5915,N_5782,N_5640);
nor U5916 (N_5916,N_5681,N_5725);
or U5917 (N_5917,N_5728,N_5735);
and U5918 (N_5918,N_5745,N_5621);
nand U5919 (N_5919,N_5630,N_5613);
and U5920 (N_5920,N_5728,N_5774);
nor U5921 (N_5921,N_5734,N_5726);
nand U5922 (N_5922,N_5783,N_5642);
nor U5923 (N_5923,N_5757,N_5648);
nand U5924 (N_5924,N_5745,N_5680);
or U5925 (N_5925,N_5643,N_5751);
or U5926 (N_5926,N_5758,N_5737);
xnor U5927 (N_5927,N_5654,N_5775);
nand U5928 (N_5928,N_5679,N_5687);
nand U5929 (N_5929,N_5722,N_5751);
or U5930 (N_5930,N_5648,N_5717);
or U5931 (N_5931,N_5761,N_5715);
or U5932 (N_5932,N_5602,N_5631);
nand U5933 (N_5933,N_5770,N_5655);
or U5934 (N_5934,N_5690,N_5635);
xor U5935 (N_5935,N_5692,N_5634);
or U5936 (N_5936,N_5718,N_5639);
nand U5937 (N_5937,N_5663,N_5749);
or U5938 (N_5938,N_5612,N_5787);
or U5939 (N_5939,N_5788,N_5777);
and U5940 (N_5940,N_5698,N_5632);
xor U5941 (N_5941,N_5618,N_5631);
or U5942 (N_5942,N_5643,N_5773);
and U5943 (N_5943,N_5606,N_5708);
xor U5944 (N_5944,N_5698,N_5769);
or U5945 (N_5945,N_5794,N_5758);
and U5946 (N_5946,N_5771,N_5605);
and U5947 (N_5947,N_5626,N_5792);
and U5948 (N_5948,N_5638,N_5762);
nor U5949 (N_5949,N_5738,N_5674);
or U5950 (N_5950,N_5614,N_5744);
nor U5951 (N_5951,N_5698,N_5617);
xnor U5952 (N_5952,N_5601,N_5633);
nand U5953 (N_5953,N_5779,N_5643);
and U5954 (N_5954,N_5754,N_5642);
and U5955 (N_5955,N_5696,N_5710);
nor U5956 (N_5956,N_5751,N_5677);
nor U5957 (N_5957,N_5650,N_5761);
xor U5958 (N_5958,N_5651,N_5684);
xnor U5959 (N_5959,N_5788,N_5716);
nor U5960 (N_5960,N_5665,N_5649);
xor U5961 (N_5961,N_5791,N_5696);
xor U5962 (N_5962,N_5664,N_5602);
xnor U5963 (N_5963,N_5627,N_5693);
and U5964 (N_5964,N_5684,N_5746);
xor U5965 (N_5965,N_5612,N_5775);
xor U5966 (N_5966,N_5706,N_5719);
xor U5967 (N_5967,N_5663,N_5715);
nand U5968 (N_5968,N_5683,N_5643);
nor U5969 (N_5969,N_5645,N_5724);
or U5970 (N_5970,N_5693,N_5738);
and U5971 (N_5971,N_5704,N_5750);
xor U5972 (N_5972,N_5619,N_5767);
and U5973 (N_5973,N_5736,N_5618);
xor U5974 (N_5974,N_5698,N_5600);
nand U5975 (N_5975,N_5743,N_5645);
nand U5976 (N_5976,N_5733,N_5684);
nor U5977 (N_5977,N_5620,N_5709);
nand U5978 (N_5978,N_5778,N_5687);
nand U5979 (N_5979,N_5766,N_5748);
nor U5980 (N_5980,N_5629,N_5780);
nand U5981 (N_5981,N_5798,N_5710);
or U5982 (N_5982,N_5746,N_5615);
nor U5983 (N_5983,N_5767,N_5749);
and U5984 (N_5984,N_5675,N_5633);
or U5985 (N_5985,N_5768,N_5658);
nor U5986 (N_5986,N_5614,N_5706);
nand U5987 (N_5987,N_5781,N_5796);
xor U5988 (N_5988,N_5748,N_5687);
or U5989 (N_5989,N_5716,N_5757);
nor U5990 (N_5990,N_5775,N_5709);
nand U5991 (N_5991,N_5755,N_5641);
or U5992 (N_5992,N_5652,N_5704);
and U5993 (N_5993,N_5612,N_5681);
or U5994 (N_5994,N_5775,N_5630);
nor U5995 (N_5995,N_5741,N_5697);
nand U5996 (N_5996,N_5615,N_5735);
and U5997 (N_5997,N_5692,N_5640);
nor U5998 (N_5998,N_5658,N_5613);
or U5999 (N_5999,N_5602,N_5610);
xnor U6000 (N_6000,N_5825,N_5941);
or U6001 (N_6001,N_5861,N_5939);
xor U6002 (N_6002,N_5838,N_5874);
nand U6003 (N_6003,N_5928,N_5977);
nand U6004 (N_6004,N_5884,N_5994);
xnor U6005 (N_6005,N_5819,N_5975);
or U6006 (N_6006,N_5964,N_5910);
xor U6007 (N_6007,N_5998,N_5892);
and U6008 (N_6008,N_5925,N_5803);
xor U6009 (N_6009,N_5967,N_5801);
or U6010 (N_6010,N_5866,N_5909);
nor U6011 (N_6011,N_5934,N_5856);
and U6012 (N_6012,N_5913,N_5822);
nor U6013 (N_6013,N_5915,N_5860);
nand U6014 (N_6014,N_5824,N_5896);
xnor U6015 (N_6015,N_5827,N_5908);
or U6016 (N_6016,N_5886,N_5836);
or U6017 (N_6017,N_5995,N_5880);
nand U6018 (N_6018,N_5963,N_5806);
xnor U6019 (N_6019,N_5931,N_5805);
nand U6020 (N_6020,N_5834,N_5976);
nand U6021 (N_6021,N_5988,N_5848);
nand U6022 (N_6022,N_5813,N_5877);
xnor U6023 (N_6023,N_5942,N_5949);
nor U6024 (N_6024,N_5843,N_5876);
xnor U6025 (N_6025,N_5930,N_5833);
xnor U6026 (N_6026,N_5887,N_5905);
nand U6027 (N_6027,N_5815,N_5804);
nor U6028 (N_6028,N_5849,N_5923);
and U6029 (N_6029,N_5831,N_5951);
nor U6030 (N_6030,N_5844,N_5904);
nor U6031 (N_6031,N_5889,N_5885);
nand U6032 (N_6032,N_5947,N_5900);
or U6033 (N_6033,N_5956,N_5914);
xor U6034 (N_6034,N_5881,N_5907);
nand U6035 (N_6035,N_5837,N_5997);
nand U6036 (N_6036,N_5882,N_5946);
or U6037 (N_6037,N_5992,N_5868);
nand U6038 (N_6038,N_5828,N_5937);
nor U6039 (N_6039,N_5812,N_5961);
xor U6040 (N_6040,N_5854,N_5902);
or U6041 (N_6041,N_5807,N_5971);
nor U6042 (N_6042,N_5936,N_5983);
or U6043 (N_6043,N_5873,N_5818);
nor U6044 (N_6044,N_5832,N_5845);
nor U6045 (N_6045,N_5809,N_5972);
and U6046 (N_6046,N_5888,N_5968);
or U6047 (N_6047,N_5962,N_5829);
or U6048 (N_6048,N_5916,N_5823);
nor U6049 (N_6049,N_5955,N_5986);
xor U6050 (N_6050,N_5872,N_5852);
nor U6051 (N_6051,N_5974,N_5863);
nand U6052 (N_6052,N_5816,N_5864);
or U6053 (N_6053,N_5959,N_5969);
and U6054 (N_6054,N_5957,N_5938);
and U6055 (N_6055,N_5912,N_5865);
nand U6056 (N_6056,N_5922,N_5891);
nand U6057 (N_6057,N_5841,N_5858);
and U6058 (N_6058,N_5929,N_5862);
nor U6059 (N_6059,N_5999,N_5878);
xnor U6060 (N_6060,N_5820,N_5993);
and U6061 (N_6061,N_5978,N_5933);
nand U6062 (N_6062,N_5871,N_5927);
nand U6063 (N_6063,N_5996,N_5945);
or U6064 (N_6064,N_5965,N_5917);
nor U6065 (N_6065,N_5835,N_5921);
and U6066 (N_6066,N_5966,N_5879);
xnor U6067 (N_6067,N_5973,N_5898);
nor U6068 (N_6068,N_5895,N_5846);
or U6069 (N_6069,N_5826,N_5958);
or U6070 (N_6070,N_5830,N_5883);
nand U6071 (N_6071,N_5919,N_5901);
nor U6072 (N_6072,N_5991,N_5897);
nand U6073 (N_6073,N_5859,N_5855);
nor U6074 (N_6074,N_5911,N_5839);
or U6075 (N_6075,N_5800,N_5875);
or U6076 (N_6076,N_5808,N_5851);
or U6077 (N_6077,N_5950,N_5980);
nand U6078 (N_6078,N_5810,N_5985);
and U6079 (N_6079,N_5948,N_5847);
xor U6080 (N_6080,N_5840,N_5867);
nand U6081 (N_6081,N_5853,N_5811);
and U6082 (N_6082,N_5920,N_5984);
nand U6083 (N_6083,N_5918,N_5926);
and U6084 (N_6084,N_5814,N_5932);
xnor U6085 (N_6085,N_5869,N_5924);
nor U6086 (N_6086,N_5987,N_5960);
or U6087 (N_6087,N_5940,N_5821);
or U6088 (N_6088,N_5990,N_5952);
or U6089 (N_6089,N_5899,N_5954);
and U6090 (N_6090,N_5842,N_5944);
or U6091 (N_6091,N_5893,N_5943);
nand U6092 (N_6092,N_5817,N_5981);
or U6093 (N_6093,N_5989,N_5870);
nand U6094 (N_6094,N_5850,N_5970);
xnor U6095 (N_6095,N_5906,N_5935);
nor U6096 (N_6096,N_5953,N_5894);
and U6097 (N_6097,N_5857,N_5979);
nor U6098 (N_6098,N_5982,N_5903);
xnor U6099 (N_6099,N_5802,N_5890);
nand U6100 (N_6100,N_5813,N_5955);
nor U6101 (N_6101,N_5894,N_5932);
nand U6102 (N_6102,N_5827,N_5899);
nor U6103 (N_6103,N_5976,N_5913);
xor U6104 (N_6104,N_5923,N_5999);
xnor U6105 (N_6105,N_5922,N_5843);
and U6106 (N_6106,N_5916,N_5826);
nor U6107 (N_6107,N_5815,N_5876);
or U6108 (N_6108,N_5991,N_5941);
nor U6109 (N_6109,N_5805,N_5927);
nor U6110 (N_6110,N_5810,N_5874);
or U6111 (N_6111,N_5962,N_5918);
xor U6112 (N_6112,N_5854,N_5807);
or U6113 (N_6113,N_5947,N_5987);
xor U6114 (N_6114,N_5962,N_5983);
and U6115 (N_6115,N_5941,N_5979);
xor U6116 (N_6116,N_5915,N_5887);
nand U6117 (N_6117,N_5974,N_5897);
and U6118 (N_6118,N_5805,N_5923);
nor U6119 (N_6119,N_5979,N_5871);
xnor U6120 (N_6120,N_5876,N_5812);
nand U6121 (N_6121,N_5956,N_5877);
nor U6122 (N_6122,N_5953,N_5979);
xnor U6123 (N_6123,N_5834,N_5988);
or U6124 (N_6124,N_5936,N_5926);
or U6125 (N_6125,N_5952,N_5920);
nor U6126 (N_6126,N_5960,N_5942);
nand U6127 (N_6127,N_5993,N_5946);
or U6128 (N_6128,N_5826,N_5860);
and U6129 (N_6129,N_5985,N_5874);
nand U6130 (N_6130,N_5925,N_5970);
nor U6131 (N_6131,N_5841,N_5998);
xor U6132 (N_6132,N_5947,N_5827);
or U6133 (N_6133,N_5894,N_5910);
nor U6134 (N_6134,N_5844,N_5916);
xnor U6135 (N_6135,N_5966,N_5953);
nor U6136 (N_6136,N_5907,N_5882);
xor U6137 (N_6137,N_5957,N_5857);
nor U6138 (N_6138,N_5835,N_5815);
xor U6139 (N_6139,N_5809,N_5874);
or U6140 (N_6140,N_5984,N_5831);
nand U6141 (N_6141,N_5804,N_5984);
and U6142 (N_6142,N_5833,N_5953);
nand U6143 (N_6143,N_5862,N_5926);
and U6144 (N_6144,N_5932,N_5819);
or U6145 (N_6145,N_5977,N_5997);
nor U6146 (N_6146,N_5932,N_5972);
nor U6147 (N_6147,N_5820,N_5995);
xnor U6148 (N_6148,N_5826,N_5854);
or U6149 (N_6149,N_5898,N_5816);
xor U6150 (N_6150,N_5977,N_5908);
or U6151 (N_6151,N_5861,N_5947);
xor U6152 (N_6152,N_5922,N_5986);
nor U6153 (N_6153,N_5866,N_5949);
nand U6154 (N_6154,N_5936,N_5817);
or U6155 (N_6155,N_5921,N_5984);
or U6156 (N_6156,N_5811,N_5932);
nor U6157 (N_6157,N_5990,N_5827);
or U6158 (N_6158,N_5973,N_5993);
nor U6159 (N_6159,N_5984,N_5904);
nor U6160 (N_6160,N_5804,N_5880);
and U6161 (N_6161,N_5806,N_5915);
and U6162 (N_6162,N_5920,N_5944);
and U6163 (N_6163,N_5878,N_5828);
or U6164 (N_6164,N_5966,N_5918);
nor U6165 (N_6165,N_5852,N_5880);
xnor U6166 (N_6166,N_5872,N_5988);
nand U6167 (N_6167,N_5935,N_5890);
xnor U6168 (N_6168,N_5998,N_5833);
and U6169 (N_6169,N_5949,N_5847);
nor U6170 (N_6170,N_5823,N_5910);
and U6171 (N_6171,N_5881,N_5887);
nand U6172 (N_6172,N_5872,N_5945);
xor U6173 (N_6173,N_5867,N_5914);
or U6174 (N_6174,N_5932,N_5984);
and U6175 (N_6175,N_5918,N_5984);
or U6176 (N_6176,N_5804,N_5844);
and U6177 (N_6177,N_5961,N_5886);
xor U6178 (N_6178,N_5949,N_5981);
nor U6179 (N_6179,N_5997,N_5990);
xnor U6180 (N_6180,N_5982,N_5812);
nor U6181 (N_6181,N_5927,N_5843);
or U6182 (N_6182,N_5937,N_5834);
or U6183 (N_6183,N_5912,N_5812);
or U6184 (N_6184,N_5905,N_5917);
and U6185 (N_6185,N_5863,N_5981);
or U6186 (N_6186,N_5816,N_5876);
nor U6187 (N_6187,N_5947,N_5876);
nor U6188 (N_6188,N_5865,N_5866);
xnor U6189 (N_6189,N_5806,N_5828);
or U6190 (N_6190,N_5874,N_5964);
or U6191 (N_6191,N_5991,N_5844);
nor U6192 (N_6192,N_5939,N_5975);
or U6193 (N_6193,N_5862,N_5880);
or U6194 (N_6194,N_5842,N_5814);
xnor U6195 (N_6195,N_5951,N_5934);
or U6196 (N_6196,N_5961,N_5811);
and U6197 (N_6197,N_5875,N_5803);
nand U6198 (N_6198,N_5981,N_5997);
nor U6199 (N_6199,N_5843,N_5874);
nor U6200 (N_6200,N_6025,N_6087);
and U6201 (N_6201,N_6072,N_6041);
xnor U6202 (N_6202,N_6058,N_6015);
and U6203 (N_6203,N_6088,N_6126);
nand U6204 (N_6204,N_6181,N_6066);
and U6205 (N_6205,N_6130,N_6115);
or U6206 (N_6206,N_6076,N_6166);
or U6207 (N_6207,N_6197,N_6174);
xor U6208 (N_6208,N_6049,N_6082);
nand U6209 (N_6209,N_6112,N_6105);
nor U6210 (N_6210,N_6110,N_6162);
xor U6211 (N_6211,N_6196,N_6185);
and U6212 (N_6212,N_6155,N_6093);
nand U6213 (N_6213,N_6172,N_6096);
or U6214 (N_6214,N_6099,N_6012);
nor U6215 (N_6215,N_6075,N_6055);
xnor U6216 (N_6216,N_6123,N_6167);
nand U6217 (N_6217,N_6141,N_6160);
xor U6218 (N_6218,N_6006,N_6031);
or U6219 (N_6219,N_6040,N_6122);
nand U6220 (N_6220,N_6084,N_6065);
and U6221 (N_6221,N_6038,N_6039);
or U6222 (N_6222,N_6043,N_6153);
or U6223 (N_6223,N_6154,N_6178);
xnor U6224 (N_6224,N_6173,N_6077);
nand U6225 (N_6225,N_6125,N_6023);
or U6226 (N_6226,N_6029,N_6177);
xor U6227 (N_6227,N_6060,N_6113);
nor U6228 (N_6228,N_6131,N_6189);
nand U6229 (N_6229,N_6182,N_6199);
or U6230 (N_6230,N_6079,N_6083);
xor U6231 (N_6231,N_6195,N_6149);
xor U6232 (N_6232,N_6192,N_6059);
nand U6233 (N_6233,N_6108,N_6033);
or U6234 (N_6234,N_6070,N_6078);
and U6235 (N_6235,N_6168,N_6103);
or U6236 (N_6236,N_6044,N_6014);
nor U6237 (N_6237,N_6135,N_6098);
or U6238 (N_6238,N_6143,N_6151);
and U6239 (N_6239,N_6089,N_6030);
nor U6240 (N_6240,N_6095,N_6045);
xnor U6241 (N_6241,N_6117,N_6063);
and U6242 (N_6242,N_6094,N_6109);
and U6243 (N_6243,N_6008,N_6165);
nor U6244 (N_6244,N_6042,N_6119);
xnor U6245 (N_6245,N_6037,N_6010);
nor U6246 (N_6246,N_6001,N_6053);
xor U6247 (N_6247,N_6187,N_6107);
or U6248 (N_6248,N_6188,N_6163);
nor U6249 (N_6249,N_6152,N_6138);
and U6250 (N_6250,N_6158,N_6056);
nand U6251 (N_6251,N_6022,N_6133);
nor U6252 (N_6252,N_6017,N_6120);
nor U6253 (N_6253,N_6136,N_6111);
or U6254 (N_6254,N_6020,N_6193);
or U6255 (N_6255,N_6074,N_6026);
xor U6256 (N_6256,N_6068,N_6027);
or U6257 (N_6257,N_6106,N_6071);
nor U6258 (N_6258,N_6144,N_6054);
or U6259 (N_6259,N_6090,N_6013);
nand U6260 (N_6260,N_6134,N_6016);
xor U6261 (N_6261,N_6018,N_6179);
and U6262 (N_6262,N_6161,N_6116);
and U6263 (N_6263,N_6190,N_6118);
or U6264 (N_6264,N_6170,N_6091);
and U6265 (N_6265,N_6024,N_6121);
or U6266 (N_6266,N_6062,N_6132);
xor U6267 (N_6267,N_6198,N_6191);
or U6268 (N_6268,N_6007,N_6028);
nor U6269 (N_6269,N_6176,N_6061);
nand U6270 (N_6270,N_6159,N_6003);
nand U6271 (N_6271,N_6036,N_6019);
and U6272 (N_6272,N_6035,N_6032);
nand U6273 (N_6273,N_6104,N_6150);
xnor U6274 (N_6274,N_6127,N_6051);
and U6275 (N_6275,N_6147,N_6085);
and U6276 (N_6276,N_6009,N_6156);
or U6277 (N_6277,N_6142,N_6048);
and U6278 (N_6278,N_6100,N_6184);
xor U6279 (N_6279,N_6157,N_6194);
or U6280 (N_6280,N_6140,N_6081);
nand U6281 (N_6281,N_6046,N_6139);
nor U6282 (N_6282,N_6097,N_6064);
or U6283 (N_6283,N_6034,N_6129);
nor U6284 (N_6284,N_6114,N_6183);
and U6285 (N_6285,N_6057,N_6002);
nor U6286 (N_6286,N_6092,N_6052);
and U6287 (N_6287,N_6080,N_6145);
nor U6288 (N_6288,N_6073,N_6086);
or U6289 (N_6289,N_6171,N_6137);
xnor U6290 (N_6290,N_6124,N_6000);
nor U6291 (N_6291,N_6186,N_6175);
or U6292 (N_6292,N_6005,N_6047);
and U6293 (N_6293,N_6004,N_6146);
or U6294 (N_6294,N_6128,N_6069);
nand U6295 (N_6295,N_6148,N_6102);
xor U6296 (N_6296,N_6101,N_6180);
and U6297 (N_6297,N_6169,N_6164);
nand U6298 (N_6298,N_6011,N_6050);
nand U6299 (N_6299,N_6067,N_6021);
xnor U6300 (N_6300,N_6050,N_6187);
nor U6301 (N_6301,N_6116,N_6042);
or U6302 (N_6302,N_6064,N_6063);
nand U6303 (N_6303,N_6143,N_6044);
nor U6304 (N_6304,N_6113,N_6083);
nor U6305 (N_6305,N_6015,N_6002);
nor U6306 (N_6306,N_6083,N_6141);
nand U6307 (N_6307,N_6060,N_6131);
nand U6308 (N_6308,N_6010,N_6019);
xor U6309 (N_6309,N_6061,N_6131);
nor U6310 (N_6310,N_6008,N_6153);
and U6311 (N_6311,N_6090,N_6132);
or U6312 (N_6312,N_6109,N_6028);
xor U6313 (N_6313,N_6083,N_6018);
and U6314 (N_6314,N_6164,N_6007);
nor U6315 (N_6315,N_6122,N_6008);
xnor U6316 (N_6316,N_6138,N_6177);
nor U6317 (N_6317,N_6002,N_6178);
xor U6318 (N_6318,N_6187,N_6015);
or U6319 (N_6319,N_6015,N_6044);
nor U6320 (N_6320,N_6168,N_6044);
and U6321 (N_6321,N_6173,N_6145);
and U6322 (N_6322,N_6019,N_6027);
nor U6323 (N_6323,N_6166,N_6193);
nor U6324 (N_6324,N_6124,N_6108);
nand U6325 (N_6325,N_6088,N_6189);
or U6326 (N_6326,N_6040,N_6185);
xor U6327 (N_6327,N_6035,N_6040);
and U6328 (N_6328,N_6100,N_6012);
nand U6329 (N_6329,N_6034,N_6098);
or U6330 (N_6330,N_6100,N_6056);
or U6331 (N_6331,N_6052,N_6145);
xnor U6332 (N_6332,N_6111,N_6157);
nand U6333 (N_6333,N_6090,N_6063);
nor U6334 (N_6334,N_6146,N_6061);
or U6335 (N_6335,N_6137,N_6036);
and U6336 (N_6336,N_6179,N_6139);
nor U6337 (N_6337,N_6000,N_6095);
or U6338 (N_6338,N_6084,N_6000);
nor U6339 (N_6339,N_6168,N_6113);
or U6340 (N_6340,N_6114,N_6123);
nand U6341 (N_6341,N_6095,N_6102);
xnor U6342 (N_6342,N_6122,N_6099);
nor U6343 (N_6343,N_6068,N_6014);
xnor U6344 (N_6344,N_6192,N_6100);
xor U6345 (N_6345,N_6191,N_6141);
nand U6346 (N_6346,N_6077,N_6192);
nand U6347 (N_6347,N_6062,N_6089);
xnor U6348 (N_6348,N_6031,N_6182);
xnor U6349 (N_6349,N_6048,N_6066);
nand U6350 (N_6350,N_6165,N_6164);
or U6351 (N_6351,N_6006,N_6085);
xor U6352 (N_6352,N_6084,N_6194);
or U6353 (N_6353,N_6085,N_6056);
or U6354 (N_6354,N_6067,N_6007);
or U6355 (N_6355,N_6175,N_6004);
xor U6356 (N_6356,N_6185,N_6152);
nand U6357 (N_6357,N_6073,N_6004);
and U6358 (N_6358,N_6070,N_6172);
nor U6359 (N_6359,N_6161,N_6107);
or U6360 (N_6360,N_6105,N_6143);
xor U6361 (N_6361,N_6183,N_6001);
or U6362 (N_6362,N_6114,N_6095);
and U6363 (N_6363,N_6027,N_6083);
nor U6364 (N_6364,N_6164,N_6124);
nor U6365 (N_6365,N_6139,N_6186);
nand U6366 (N_6366,N_6042,N_6189);
xor U6367 (N_6367,N_6023,N_6167);
and U6368 (N_6368,N_6064,N_6141);
and U6369 (N_6369,N_6108,N_6176);
nor U6370 (N_6370,N_6198,N_6097);
xnor U6371 (N_6371,N_6119,N_6036);
nor U6372 (N_6372,N_6151,N_6054);
xnor U6373 (N_6373,N_6022,N_6006);
xnor U6374 (N_6374,N_6007,N_6195);
xnor U6375 (N_6375,N_6120,N_6155);
nand U6376 (N_6376,N_6109,N_6155);
nand U6377 (N_6377,N_6070,N_6155);
nor U6378 (N_6378,N_6041,N_6088);
xor U6379 (N_6379,N_6091,N_6009);
xor U6380 (N_6380,N_6145,N_6113);
nand U6381 (N_6381,N_6167,N_6095);
nand U6382 (N_6382,N_6149,N_6075);
or U6383 (N_6383,N_6119,N_6022);
or U6384 (N_6384,N_6055,N_6130);
and U6385 (N_6385,N_6117,N_6151);
nand U6386 (N_6386,N_6126,N_6173);
xor U6387 (N_6387,N_6162,N_6144);
xor U6388 (N_6388,N_6019,N_6176);
xnor U6389 (N_6389,N_6137,N_6061);
or U6390 (N_6390,N_6022,N_6168);
nand U6391 (N_6391,N_6014,N_6015);
nor U6392 (N_6392,N_6018,N_6021);
and U6393 (N_6393,N_6057,N_6186);
and U6394 (N_6394,N_6164,N_6128);
and U6395 (N_6395,N_6195,N_6031);
or U6396 (N_6396,N_6076,N_6074);
xnor U6397 (N_6397,N_6077,N_6045);
and U6398 (N_6398,N_6094,N_6195);
nor U6399 (N_6399,N_6087,N_6054);
nand U6400 (N_6400,N_6295,N_6391);
xor U6401 (N_6401,N_6233,N_6296);
nor U6402 (N_6402,N_6349,N_6331);
or U6403 (N_6403,N_6356,N_6247);
nor U6404 (N_6404,N_6362,N_6286);
xnor U6405 (N_6405,N_6281,N_6334);
nor U6406 (N_6406,N_6360,N_6323);
nor U6407 (N_6407,N_6346,N_6377);
or U6408 (N_6408,N_6292,N_6317);
or U6409 (N_6409,N_6273,N_6359);
nand U6410 (N_6410,N_6228,N_6226);
nor U6411 (N_6411,N_6297,N_6245);
nand U6412 (N_6412,N_6382,N_6255);
or U6413 (N_6413,N_6305,N_6222);
nand U6414 (N_6414,N_6306,N_6395);
nand U6415 (N_6415,N_6278,N_6336);
xnor U6416 (N_6416,N_6361,N_6376);
or U6417 (N_6417,N_6308,N_6341);
nor U6418 (N_6418,N_6223,N_6230);
nand U6419 (N_6419,N_6280,N_6271);
nand U6420 (N_6420,N_6327,N_6358);
or U6421 (N_6421,N_6350,N_6256);
nand U6422 (N_6422,N_6248,N_6348);
xnor U6423 (N_6423,N_6347,N_6259);
and U6424 (N_6424,N_6231,N_6343);
nand U6425 (N_6425,N_6284,N_6329);
or U6426 (N_6426,N_6367,N_6325);
nand U6427 (N_6427,N_6312,N_6219);
nand U6428 (N_6428,N_6290,N_6342);
and U6429 (N_6429,N_6217,N_6332);
nand U6430 (N_6430,N_6270,N_6241);
or U6431 (N_6431,N_6339,N_6394);
or U6432 (N_6432,N_6242,N_6236);
or U6433 (N_6433,N_6299,N_6243);
nand U6434 (N_6434,N_6276,N_6269);
xnor U6435 (N_6435,N_6303,N_6211);
nand U6436 (N_6436,N_6294,N_6310);
or U6437 (N_6437,N_6291,N_6220);
xnor U6438 (N_6438,N_6352,N_6216);
xor U6439 (N_6439,N_6316,N_6390);
and U6440 (N_6440,N_6239,N_6398);
nand U6441 (N_6441,N_6311,N_6357);
nand U6442 (N_6442,N_6205,N_6285);
or U6443 (N_6443,N_6372,N_6373);
nand U6444 (N_6444,N_6232,N_6214);
nand U6445 (N_6445,N_6335,N_6399);
or U6446 (N_6446,N_6246,N_6202);
nor U6447 (N_6447,N_6293,N_6266);
or U6448 (N_6448,N_6338,N_6340);
nor U6449 (N_6449,N_6314,N_6386);
and U6450 (N_6450,N_6392,N_6279);
nor U6451 (N_6451,N_6227,N_6326);
or U6452 (N_6452,N_6218,N_6258);
nand U6453 (N_6453,N_6207,N_6371);
nand U6454 (N_6454,N_6263,N_6221);
nor U6455 (N_6455,N_6261,N_6368);
or U6456 (N_6456,N_6351,N_6240);
or U6457 (N_6457,N_6389,N_6337);
or U6458 (N_6458,N_6387,N_6262);
xnor U6459 (N_6459,N_6253,N_6330);
nor U6460 (N_6460,N_6324,N_6288);
and U6461 (N_6461,N_6363,N_6210);
xnor U6462 (N_6462,N_6328,N_6287);
xor U6463 (N_6463,N_6215,N_6260);
nand U6464 (N_6464,N_6378,N_6275);
nor U6465 (N_6465,N_6204,N_6282);
or U6466 (N_6466,N_6397,N_6251);
and U6467 (N_6467,N_6267,N_6315);
or U6468 (N_6468,N_6307,N_6318);
nor U6469 (N_6469,N_6224,N_6381);
nor U6470 (N_6470,N_6298,N_6369);
xnor U6471 (N_6471,N_6244,N_6237);
xor U6472 (N_6472,N_6268,N_6383);
and U6473 (N_6473,N_6225,N_6200);
and U6474 (N_6474,N_6264,N_6379);
and U6475 (N_6475,N_6234,N_6322);
xnor U6476 (N_6476,N_6374,N_6353);
nor U6477 (N_6477,N_6208,N_6364);
nand U6478 (N_6478,N_6254,N_6355);
nand U6479 (N_6479,N_6229,N_6283);
or U6480 (N_6480,N_6345,N_6252);
nor U6481 (N_6481,N_6313,N_6212);
and U6482 (N_6482,N_6272,N_6302);
nand U6483 (N_6483,N_6300,N_6344);
nor U6484 (N_6484,N_6309,N_6321);
nor U6485 (N_6485,N_6304,N_6289);
xnor U6486 (N_6486,N_6274,N_6396);
xor U6487 (N_6487,N_6380,N_6388);
nor U6488 (N_6488,N_6250,N_6319);
nor U6489 (N_6489,N_6370,N_6365);
xnor U6490 (N_6490,N_6375,N_6238);
nand U6491 (N_6491,N_6209,N_6333);
and U6492 (N_6492,N_6213,N_6354);
xnor U6493 (N_6493,N_6320,N_6257);
and U6494 (N_6494,N_6206,N_6384);
nand U6495 (N_6495,N_6277,N_6203);
or U6496 (N_6496,N_6249,N_6201);
nor U6497 (N_6497,N_6366,N_6393);
or U6498 (N_6498,N_6301,N_6385);
or U6499 (N_6499,N_6265,N_6235);
nor U6500 (N_6500,N_6357,N_6285);
and U6501 (N_6501,N_6399,N_6382);
xnor U6502 (N_6502,N_6331,N_6346);
or U6503 (N_6503,N_6385,N_6353);
xnor U6504 (N_6504,N_6305,N_6231);
nor U6505 (N_6505,N_6372,N_6385);
or U6506 (N_6506,N_6205,N_6226);
or U6507 (N_6507,N_6349,N_6259);
or U6508 (N_6508,N_6388,N_6384);
or U6509 (N_6509,N_6381,N_6341);
nand U6510 (N_6510,N_6371,N_6348);
or U6511 (N_6511,N_6272,N_6340);
xnor U6512 (N_6512,N_6258,N_6394);
and U6513 (N_6513,N_6308,N_6241);
xor U6514 (N_6514,N_6247,N_6314);
xor U6515 (N_6515,N_6399,N_6312);
xnor U6516 (N_6516,N_6305,N_6314);
or U6517 (N_6517,N_6259,N_6278);
or U6518 (N_6518,N_6328,N_6311);
nor U6519 (N_6519,N_6360,N_6320);
xor U6520 (N_6520,N_6367,N_6362);
nor U6521 (N_6521,N_6257,N_6364);
nand U6522 (N_6522,N_6388,N_6210);
and U6523 (N_6523,N_6301,N_6341);
and U6524 (N_6524,N_6214,N_6386);
nor U6525 (N_6525,N_6215,N_6347);
nor U6526 (N_6526,N_6327,N_6378);
nand U6527 (N_6527,N_6380,N_6283);
nor U6528 (N_6528,N_6241,N_6234);
xnor U6529 (N_6529,N_6245,N_6349);
nand U6530 (N_6530,N_6290,N_6258);
nor U6531 (N_6531,N_6322,N_6377);
and U6532 (N_6532,N_6238,N_6327);
or U6533 (N_6533,N_6367,N_6392);
or U6534 (N_6534,N_6243,N_6291);
and U6535 (N_6535,N_6250,N_6313);
or U6536 (N_6536,N_6219,N_6290);
xor U6537 (N_6537,N_6267,N_6206);
nand U6538 (N_6538,N_6356,N_6323);
xnor U6539 (N_6539,N_6304,N_6361);
nor U6540 (N_6540,N_6235,N_6328);
nand U6541 (N_6541,N_6289,N_6393);
and U6542 (N_6542,N_6327,N_6207);
or U6543 (N_6543,N_6200,N_6354);
nor U6544 (N_6544,N_6304,N_6238);
nand U6545 (N_6545,N_6357,N_6389);
xor U6546 (N_6546,N_6389,N_6246);
nand U6547 (N_6547,N_6393,N_6358);
nand U6548 (N_6548,N_6227,N_6300);
or U6549 (N_6549,N_6261,N_6255);
and U6550 (N_6550,N_6270,N_6303);
or U6551 (N_6551,N_6209,N_6385);
nand U6552 (N_6552,N_6352,N_6329);
nand U6553 (N_6553,N_6332,N_6387);
nor U6554 (N_6554,N_6271,N_6337);
or U6555 (N_6555,N_6283,N_6255);
nor U6556 (N_6556,N_6353,N_6340);
nand U6557 (N_6557,N_6220,N_6292);
nand U6558 (N_6558,N_6293,N_6327);
and U6559 (N_6559,N_6286,N_6221);
xnor U6560 (N_6560,N_6238,N_6305);
and U6561 (N_6561,N_6300,N_6334);
and U6562 (N_6562,N_6280,N_6320);
nand U6563 (N_6563,N_6237,N_6391);
or U6564 (N_6564,N_6341,N_6270);
nor U6565 (N_6565,N_6228,N_6381);
nor U6566 (N_6566,N_6201,N_6236);
nand U6567 (N_6567,N_6208,N_6391);
or U6568 (N_6568,N_6261,N_6349);
nand U6569 (N_6569,N_6232,N_6315);
and U6570 (N_6570,N_6355,N_6368);
and U6571 (N_6571,N_6251,N_6320);
nand U6572 (N_6572,N_6292,N_6287);
nor U6573 (N_6573,N_6399,N_6329);
xor U6574 (N_6574,N_6247,N_6380);
or U6575 (N_6575,N_6394,N_6328);
or U6576 (N_6576,N_6316,N_6374);
nand U6577 (N_6577,N_6386,N_6341);
and U6578 (N_6578,N_6317,N_6229);
and U6579 (N_6579,N_6342,N_6373);
nor U6580 (N_6580,N_6291,N_6202);
and U6581 (N_6581,N_6278,N_6333);
and U6582 (N_6582,N_6340,N_6365);
or U6583 (N_6583,N_6224,N_6263);
nor U6584 (N_6584,N_6326,N_6344);
nor U6585 (N_6585,N_6310,N_6362);
or U6586 (N_6586,N_6244,N_6362);
nor U6587 (N_6587,N_6389,N_6262);
or U6588 (N_6588,N_6311,N_6321);
and U6589 (N_6589,N_6289,N_6239);
xor U6590 (N_6590,N_6317,N_6214);
or U6591 (N_6591,N_6381,N_6258);
and U6592 (N_6592,N_6250,N_6393);
nand U6593 (N_6593,N_6219,N_6272);
nand U6594 (N_6594,N_6208,N_6206);
nor U6595 (N_6595,N_6240,N_6273);
and U6596 (N_6596,N_6252,N_6304);
or U6597 (N_6597,N_6295,N_6399);
and U6598 (N_6598,N_6394,N_6273);
or U6599 (N_6599,N_6343,N_6364);
and U6600 (N_6600,N_6500,N_6538);
xnor U6601 (N_6601,N_6571,N_6592);
nor U6602 (N_6602,N_6595,N_6404);
nor U6603 (N_6603,N_6587,N_6578);
or U6604 (N_6604,N_6575,N_6461);
xnor U6605 (N_6605,N_6525,N_6492);
or U6606 (N_6606,N_6511,N_6517);
and U6607 (N_6607,N_6530,N_6545);
nand U6608 (N_6608,N_6574,N_6512);
nor U6609 (N_6609,N_6408,N_6467);
nor U6610 (N_6610,N_6481,N_6491);
nor U6611 (N_6611,N_6564,N_6448);
nor U6612 (N_6612,N_6583,N_6487);
and U6613 (N_6613,N_6597,N_6421);
nor U6614 (N_6614,N_6485,N_6503);
nor U6615 (N_6615,N_6432,N_6430);
nand U6616 (N_6616,N_6419,N_6572);
nor U6617 (N_6617,N_6405,N_6560);
nand U6618 (N_6618,N_6537,N_6407);
or U6619 (N_6619,N_6562,N_6541);
and U6620 (N_6620,N_6457,N_6468);
and U6621 (N_6621,N_6593,N_6454);
or U6622 (N_6622,N_6518,N_6416);
and U6623 (N_6623,N_6473,N_6488);
xnor U6624 (N_6624,N_6435,N_6453);
nand U6625 (N_6625,N_6523,N_6563);
or U6626 (N_6626,N_6411,N_6544);
nand U6627 (N_6627,N_6459,N_6504);
nor U6628 (N_6628,N_6494,N_6480);
and U6629 (N_6629,N_6402,N_6521);
nand U6630 (N_6630,N_6425,N_6472);
nand U6631 (N_6631,N_6596,N_6479);
and U6632 (N_6632,N_6505,N_6489);
or U6633 (N_6633,N_6499,N_6447);
nand U6634 (N_6634,N_6599,N_6566);
and U6635 (N_6635,N_6428,N_6438);
xnor U6636 (N_6636,N_6460,N_6439);
nand U6637 (N_6637,N_6547,N_6510);
xnor U6638 (N_6638,N_6549,N_6466);
or U6639 (N_6639,N_6420,N_6514);
xnor U6640 (N_6640,N_6444,N_6427);
nand U6641 (N_6641,N_6590,N_6410);
nor U6642 (N_6642,N_6539,N_6450);
xnor U6643 (N_6643,N_6565,N_6497);
nand U6644 (N_6644,N_6508,N_6550);
nor U6645 (N_6645,N_6465,N_6553);
xnor U6646 (N_6646,N_6559,N_6464);
nor U6647 (N_6647,N_6422,N_6556);
nor U6648 (N_6648,N_6406,N_6548);
or U6649 (N_6649,N_6570,N_6569);
nor U6650 (N_6650,N_6433,N_6412);
xor U6651 (N_6651,N_6598,N_6482);
or U6652 (N_6652,N_6436,N_6437);
nand U6653 (N_6653,N_6582,N_6469);
and U6654 (N_6654,N_6452,N_6451);
xor U6655 (N_6655,N_6536,N_6568);
nand U6656 (N_6656,N_6576,N_6535);
xnor U6657 (N_6657,N_6413,N_6417);
nand U6658 (N_6658,N_6506,N_6586);
and U6659 (N_6659,N_6594,N_6400);
xnor U6660 (N_6660,N_6414,N_6580);
and U6661 (N_6661,N_6552,N_6584);
nand U6662 (N_6662,N_6484,N_6534);
xnor U6663 (N_6663,N_6458,N_6516);
nand U6664 (N_6664,N_6585,N_6532);
xor U6665 (N_6665,N_6507,N_6475);
xor U6666 (N_6666,N_6431,N_6558);
nor U6667 (N_6667,N_6526,N_6401);
nand U6668 (N_6668,N_6557,N_6409);
and U6669 (N_6669,N_6529,N_6490);
and U6670 (N_6670,N_6415,N_6522);
nor U6671 (N_6671,N_6561,N_6513);
or U6672 (N_6672,N_6471,N_6577);
nand U6673 (N_6673,N_6495,N_6589);
xnor U6674 (N_6674,N_6446,N_6524);
xor U6675 (N_6675,N_6515,N_6493);
xor U6676 (N_6676,N_6442,N_6477);
nand U6677 (N_6677,N_6527,N_6474);
and U6678 (N_6678,N_6486,N_6456);
nand U6679 (N_6679,N_6551,N_6573);
nand U6680 (N_6680,N_6403,N_6581);
or U6681 (N_6681,N_6449,N_6445);
and U6682 (N_6682,N_6455,N_6426);
and U6683 (N_6683,N_6509,N_6498);
nand U6684 (N_6684,N_6443,N_6520);
or U6685 (N_6685,N_6418,N_6519);
xor U6686 (N_6686,N_6476,N_6554);
nor U6687 (N_6687,N_6546,N_6543);
nand U6688 (N_6688,N_6528,N_6591);
or U6689 (N_6689,N_6542,N_6424);
xor U6690 (N_6690,N_6531,N_6501);
and U6691 (N_6691,N_6567,N_6429);
xnor U6692 (N_6692,N_6502,N_6555);
xor U6693 (N_6693,N_6496,N_6533);
nor U6694 (N_6694,N_6483,N_6478);
nand U6695 (N_6695,N_6588,N_6423);
and U6696 (N_6696,N_6540,N_6434);
nor U6697 (N_6697,N_6463,N_6440);
xor U6698 (N_6698,N_6579,N_6441);
and U6699 (N_6699,N_6470,N_6462);
or U6700 (N_6700,N_6493,N_6475);
and U6701 (N_6701,N_6564,N_6466);
nor U6702 (N_6702,N_6534,N_6424);
xnor U6703 (N_6703,N_6486,N_6409);
nand U6704 (N_6704,N_6482,N_6597);
nor U6705 (N_6705,N_6500,N_6435);
nor U6706 (N_6706,N_6579,N_6566);
or U6707 (N_6707,N_6541,N_6494);
nor U6708 (N_6708,N_6438,N_6539);
and U6709 (N_6709,N_6477,N_6502);
or U6710 (N_6710,N_6530,N_6473);
nand U6711 (N_6711,N_6435,N_6422);
or U6712 (N_6712,N_6498,N_6468);
and U6713 (N_6713,N_6404,N_6555);
nor U6714 (N_6714,N_6556,N_6406);
nand U6715 (N_6715,N_6558,N_6482);
and U6716 (N_6716,N_6526,N_6427);
xor U6717 (N_6717,N_6427,N_6572);
or U6718 (N_6718,N_6473,N_6449);
and U6719 (N_6719,N_6587,N_6424);
nor U6720 (N_6720,N_6598,N_6578);
and U6721 (N_6721,N_6475,N_6426);
or U6722 (N_6722,N_6562,N_6522);
nand U6723 (N_6723,N_6425,N_6565);
and U6724 (N_6724,N_6581,N_6479);
nand U6725 (N_6725,N_6459,N_6518);
and U6726 (N_6726,N_6461,N_6570);
or U6727 (N_6727,N_6442,N_6569);
nand U6728 (N_6728,N_6475,N_6584);
or U6729 (N_6729,N_6408,N_6400);
nor U6730 (N_6730,N_6567,N_6495);
nor U6731 (N_6731,N_6450,N_6525);
xor U6732 (N_6732,N_6511,N_6580);
nor U6733 (N_6733,N_6409,N_6584);
and U6734 (N_6734,N_6477,N_6562);
or U6735 (N_6735,N_6444,N_6469);
nand U6736 (N_6736,N_6555,N_6486);
and U6737 (N_6737,N_6530,N_6586);
nor U6738 (N_6738,N_6410,N_6534);
and U6739 (N_6739,N_6400,N_6526);
nor U6740 (N_6740,N_6593,N_6519);
xnor U6741 (N_6741,N_6421,N_6573);
nor U6742 (N_6742,N_6470,N_6550);
xnor U6743 (N_6743,N_6408,N_6495);
and U6744 (N_6744,N_6508,N_6462);
or U6745 (N_6745,N_6467,N_6537);
nor U6746 (N_6746,N_6458,N_6582);
nand U6747 (N_6747,N_6412,N_6565);
and U6748 (N_6748,N_6529,N_6407);
and U6749 (N_6749,N_6413,N_6450);
nor U6750 (N_6750,N_6547,N_6500);
nand U6751 (N_6751,N_6424,N_6523);
nand U6752 (N_6752,N_6409,N_6441);
xnor U6753 (N_6753,N_6588,N_6413);
and U6754 (N_6754,N_6493,N_6531);
nand U6755 (N_6755,N_6583,N_6466);
or U6756 (N_6756,N_6496,N_6553);
or U6757 (N_6757,N_6563,N_6448);
and U6758 (N_6758,N_6569,N_6417);
and U6759 (N_6759,N_6544,N_6583);
nand U6760 (N_6760,N_6570,N_6536);
nor U6761 (N_6761,N_6478,N_6554);
or U6762 (N_6762,N_6583,N_6467);
nand U6763 (N_6763,N_6503,N_6450);
xor U6764 (N_6764,N_6453,N_6458);
nand U6765 (N_6765,N_6439,N_6591);
xor U6766 (N_6766,N_6427,N_6551);
xor U6767 (N_6767,N_6435,N_6498);
or U6768 (N_6768,N_6441,N_6596);
and U6769 (N_6769,N_6426,N_6555);
nor U6770 (N_6770,N_6511,N_6565);
or U6771 (N_6771,N_6585,N_6492);
nand U6772 (N_6772,N_6415,N_6449);
and U6773 (N_6773,N_6446,N_6506);
xnor U6774 (N_6774,N_6564,N_6522);
or U6775 (N_6775,N_6546,N_6577);
nor U6776 (N_6776,N_6449,N_6513);
or U6777 (N_6777,N_6540,N_6474);
xnor U6778 (N_6778,N_6428,N_6448);
nor U6779 (N_6779,N_6457,N_6589);
xnor U6780 (N_6780,N_6448,N_6538);
nor U6781 (N_6781,N_6456,N_6549);
or U6782 (N_6782,N_6593,N_6493);
xor U6783 (N_6783,N_6595,N_6564);
and U6784 (N_6784,N_6444,N_6461);
and U6785 (N_6785,N_6591,N_6477);
nor U6786 (N_6786,N_6562,N_6594);
or U6787 (N_6787,N_6474,N_6430);
xor U6788 (N_6788,N_6451,N_6465);
nor U6789 (N_6789,N_6546,N_6568);
or U6790 (N_6790,N_6515,N_6441);
xnor U6791 (N_6791,N_6562,N_6427);
and U6792 (N_6792,N_6477,N_6538);
nor U6793 (N_6793,N_6402,N_6474);
xnor U6794 (N_6794,N_6453,N_6529);
nor U6795 (N_6795,N_6485,N_6501);
nand U6796 (N_6796,N_6413,N_6425);
and U6797 (N_6797,N_6414,N_6547);
and U6798 (N_6798,N_6560,N_6411);
and U6799 (N_6799,N_6458,N_6520);
and U6800 (N_6800,N_6721,N_6765);
xor U6801 (N_6801,N_6688,N_6604);
nand U6802 (N_6802,N_6775,N_6681);
xor U6803 (N_6803,N_6719,N_6639);
and U6804 (N_6804,N_6735,N_6726);
or U6805 (N_6805,N_6745,N_6792);
xor U6806 (N_6806,N_6715,N_6614);
and U6807 (N_6807,N_6632,N_6606);
or U6808 (N_6808,N_6679,N_6694);
and U6809 (N_6809,N_6706,N_6737);
nor U6810 (N_6810,N_6654,N_6616);
and U6811 (N_6811,N_6796,N_6750);
nand U6812 (N_6812,N_6778,N_6731);
or U6813 (N_6813,N_6710,N_6633);
and U6814 (N_6814,N_6774,N_6655);
nand U6815 (N_6815,N_6732,N_6790);
xor U6816 (N_6816,N_6742,N_6646);
or U6817 (N_6817,N_6755,N_6684);
or U6818 (N_6818,N_6608,N_6667);
or U6819 (N_6819,N_6747,N_6795);
xor U6820 (N_6820,N_6611,N_6758);
or U6821 (N_6821,N_6787,N_6615);
or U6822 (N_6822,N_6709,N_6723);
or U6823 (N_6823,N_6617,N_6762);
nand U6824 (N_6824,N_6648,N_6776);
nor U6825 (N_6825,N_6720,N_6647);
nand U6826 (N_6826,N_6707,N_6601);
and U6827 (N_6827,N_6618,N_6786);
nor U6828 (N_6828,N_6751,N_6634);
or U6829 (N_6829,N_6749,N_6711);
and U6830 (N_6830,N_6718,N_6635);
xor U6831 (N_6831,N_6703,N_6780);
and U6832 (N_6832,N_6739,N_6753);
nand U6833 (N_6833,N_6650,N_6717);
or U6834 (N_6834,N_6702,N_6638);
and U6835 (N_6835,N_6769,N_6607);
xnor U6836 (N_6836,N_6657,N_6603);
and U6837 (N_6837,N_6687,N_6701);
nor U6838 (N_6838,N_6783,N_6675);
xor U6839 (N_6839,N_6788,N_6757);
or U6840 (N_6840,N_6649,N_6628);
and U6841 (N_6841,N_6665,N_6724);
xor U6842 (N_6842,N_6690,N_6798);
nor U6843 (N_6843,N_6602,N_6626);
nor U6844 (N_6844,N_6645,N_6781);
or U6845 (N_6845,N_6669,N_6754);
or U6846 (N_6846,N_6704,N_6637);
xnor U6847 (N_6847,N_6625,N_6727);
and U6848 (N_6848,N_6664,N_6714);
and U6849 (N_6849,N_6764,N_6784);
or U6850 (N_6850,N_6746,N_6643);
or U6851 (N_6851,N_6629,N_6779);
or U6852 (N_6852,N_6676,N_6729);
nor U6853 (N_6853,N_6712,N_6767);
and U6854 (N_6854,N_6600,N_6619);
xnor U6855 (N_6855,N_6682,N_6656);
and U6856 (N_6856,N_6631,N_6785);
or U6857 (N_6857,N_6661,N_6700);
or U6858 (N_6858,N_6685,N_6695);
or U6859 (N_6859,N_6692,N_6741);
and U6860 (N_6860,N_6678,N_6623);
nand U6861 (N_6861,N_6662,N_6761);
nor U6862 (N_6862,N_6760,N_6734);
xnor U6863 (N_6863,N_6738,N_6689);
nand U6864 (N_6864,N_6708,N_6653);
or U6865 (N_6865,N_6728,N_6713);
xnor U6866 (N_6866,N_6644,N_6716);
nand U6867 (N_6867,N_6686,N_6766);
nor U6868 (N_6868,N_6797,N_6612);
xnor U6869 (N_6869,N_6671,N_6770);
nand U6870 (N_6870,N_6620,N_6759);
and U6871 (N_6871,N_6773,N_6693);
and U6872 (N_6872,N_6677,N_6610);
nor U6873 (N_6873,N_6722,N_6641);
nor U6874 (N_6874,N_6672,N_6642);
nand U6875 (N_6875,N_6621,N_6670);
xnor U6876 (N_6876,N_6697,N_6624);
or U6877 (N_6877,N_6660,N_6699);
xnor U6878 (N_6878,N_6789,N_6768);
xnor U6879 (N_6879,N_6622,N_6705);
and U6880 (N_6880,N_6748,N_6791);
xnor U6881 (N_6881,N_6782,N_6733);
or U6882 (N_6882,N_6794,N_6627);
nor U6883 (N_6883,N_6652,N_6609);
nand U6884 (N_6884,N_6698,N_6613);
and U6885 (N_6885,N_6658,N_6752);
or U6886 (N_6886,N_6763,N_6605);
and U6887 (N_6887,N_6696,N_6744);
or U6888 (N_6888,N_6691,N_6771);
nand U6889 (N_6889,N_6651,N_6683);
xor U6890 (N_6890,N_6736,N_6756);
or U6891 (N_6891,N_6743,N_6725);
or U6892 (N_6892,N_6674,N_6777);
xor U6893 (N_6893,N_6740,N_6673);
or U6894 (N_6894,N_6730,N_6666);
and U6895 (N_6895,N_6772,N_6636);
nor U6896 (N_6896,N_6799,N_6659);
nor U6897 (N_6897,N_6640,N_6630);
xnor U6898 (N_6898,N_6680,N_6793);
xnor U6899 (N_6899,N_6663,N_6668);
nand U6900 (N_6900,N_6737,N_6783);
nor U6901 (N_6901,N_6613,N_6673);
and U6902 (N_6902,N_6685,N_6621);
and U6903 (N_6903,N_6755,N_6780);
nor U6904 (N_6904,N_6665,N_6691);
xor U6905 (N_6905,N_6701,N_6714);
nand U6906 (N_6906,N_6616,N_6657);
nand U6907 (N_6907,N_6660,N_6784);
and U6908 (N_6908,N_6737,N_6666);
and U6909 (N_6909,N_6666,N_6600);
nand U6910 (N_6910,N_6687,N_6798);
nor U6911 (N_6911,N_6720,N_6668);
nor U6912 (N_6912,N_6731,N_6716);
xor U6913 (N_6913,N_6649,N_6637);
xnor U6914 (N_6914,N_6650,N_6777);
xor U6915 (N_6915,N_6780,N_6685);
xnor U6916 (N_6916,N_6680,N_6611);
xnor U6917 (N_6917,N_6770,N_6661);
xnor U6918 (N_6918,N_6611,N_6695);
xor U6919 (N_6919,N_6752,N_6664);
nor U6920 (N_6920,N_6708,N_6788);
nor U6921 (N_6921,N_6643,N_6644);
nand U6922 (N_6922,N_6704,N_6699);
xor U6923 (N_6923,N_6675,N_6781);
and U6924 (N_6924,N_6648,N_6691);
and U6925 (N_6925,N_6663,N_6635);
xor U6926 (N_6926,N_6600,N_6616);
nor U6927 (N_6927,N_6652,N_6698);
nand U6928 (N_6928,N_6601,N_6672);
and U6929 (N_6929,N_6625,N_6698);
nand U6930 (N_6930,N_6792,N_6701);
nor U6931 (N_6931,N_6631,N_6676);
or U6932 (N_6932,N_6776,N_6671);
or U6933 (N_6933,N_6611,N_6731);
nor U6934 (N_6934,N_6724,N_6678);
xor U6935 (N_6935,N_6766,N_6746);
xor U6936 (N_6936,N_6719,N_6760);
xor U6937 (N_6937,N_6730,N_6698);
nor U6938 (N_6938,N_6614,N_6646);
xnor U6939 (N_6939,N_6713,N_6798);
or U6940 (N_6940,N_6640,N_6787);
nand U6941 (N_6941,N_6765,N_6720);
nand U6942 (N_6942,N_6602,N_6638);
xnor U6943 (N_6943,N_6746,N_6690);
or U6944 (N_6944,N_6640,N_6613);
nor U6945 (N_6945,N_6646,N_6706);
and U6946 (N_6946,N_6653,N_6784);
nor U6947 (N_6947,N_6683,N_6795);
nand U6948 (N_6948,N_6624,N_6728);
or U6949 (N_6949,N_6674,N_6753);
xor U6950 (N_6950,N_6761,N_6700);
or U6951 (N_6951,N_6719,N_6739);
nor U6952 (N_6952,N_6616,N_6620);
nor U6953 (N_6953,N_6638,N_6615);
xnor U6954 (N_6954,N_6788,N_6681);
nor U6955 (N_6955,N_6701,N_6618);
and U6956 (N_6956,N_6681,N_6743);
or U6957 (N_6957,N_6779,N_6721);
nand U6958 (N_6958,N_6666,N_6718);
or U6959 (N_6959,N_6771,N_6715);
or U6960 (N_6960,N_6783,N_6784);
nand U6961 (N_6961,N_6747,N_6791);
nor U6962 (N_6962,N_6690,N_6770);
nand U6963 (N_6963,N_6608,N_6617);
nand U6964 (N_6964,N_6739,N_6625);
or U6965 (N_6965,N_6798,N_6602);
or U6966 (N_6966,N_6664,N_6704);
and U6967 (N_6967,N_6684,N_6664);
or U6968 (N_6968,N_6640,N_6718);
xor U6969 (N_6969,N_6734,N_6668);
and U6970 (N_6970,N_6786,N_6757);
xnor U6971 (N_6971,N_6729,N_6670);
xnor U6972 (N_6972,N_6758,N_6711);
or U6973 (N_6973,N_6768,N_6782);
xnor U6974 (N_6974,N_6656,N_6783);
or U6975 (N_6975,N_6654,N_6752);
and U6976 (N_6976,N_6692,N_6667);
or U6977 (N_6977,N_6724,N_6712);
or U6978 (N_6978,N_6648,N_6773);
xnor U6979 (N_6979,N_6682,N_6766);
nand U6980 (N_6980,N_6716,N_6791);
and U6981 (N_6981,N_6614,N_6659);
and U6982 (N_6982,N_6673,N_6663);
nor U6983 (N_6983,N_6695,N_6762);
or U6984 (N_6984,N_6735,N_6796);
and U6985 (N_6985,N_6671,N_6733);
nor U6986 (N_6986,N_6747,N_6669);
nor U6987 (N_6987,N_6698,N_6740);
xnor U6988 (N_6988,N_6723,N_6699);
or U6989 (N_6989,N_6642,N_6710);
xor U6990 (N_6990,N_6730,N_6778);
xnor U6991 (N_6991,N_6660,N_6600);
xnor U6992 (N_6992,N_6709,N_6694);
and U6993 (N_6993,N_6755,N_6636);
and U6994 (N_6994,N_6723,N_6712);
nor U6995 (N_6995,N_6730,N_6717);
and U6996 (N_6996,N_6701,N_6754);
or U6997 (N_6997,N_6645,N_6630);
nand U6998 (N_6998,N_6620,N_6732);
nand U6999 (N_6999,N_6725,N_6789);
xnor U7000 (N_7000,N_6983,N_6989);
xor U7001 (N_7001,N_6963,N_6978);
xnor U7002 (N_7002,N_6845,N_6887);
xnor U7003 (N_7003,N_6830,N_6891);
nand U7004 (N_7004,N_6976,N_6907);
xor U7005 (N_7005,N_6831,N_6829);
or U7006 (N_7006,N_6881,N_6902);
nand U7007 (N_7007,N_6997,N_6851);
nor U7008 (N_7008,N_6872,N_6812);
or U7009 (N_7009,N_6802,N_6888);
or U7010 (N_7010,N_6856,N_6846);
or U7011 (N_7011,N_6909,N_6984);
nor U7012 (N_7012,N_6925,N_6981);
nor U7013 (N_7013,N_6901,N_6826);
xnor U7014 (N_7014,N_6899,N_6823);
and U7015 (N_7015,N_6889,N_6906);
or U7016 (N_7016,N_6842,N_6999);
nand U7017 (N_7017,N_6897,N_6835);
xor U7018 (N_7018,N_6828,N_6915);
nor U7019 (N_7019,N_6886,N_6844);
nor U7020 (N_7020,N_6814,N_6863);
and U7021 (N_7021,N_6813,N_6838);
and U7022 (N_7022,N_6900,N_6904);
xor U7023 (N_7023,N_6993,N_6950);
xnor U7024 (N_7024,N_6815,N_6956);
nor U7025 (N_7025,N_6874,N_6849);
xnor U7026 (N_7026,N_6917,N_6857);
nand U7027 (N_7027,N_6967,N_6810);
and U7028 (N_7028,N_6855,N_6940);
and U7029 (N_7029,N_6873,N_6858);
xor U7030 (N_7030,N_6961,N_6820);
nand U7031 (N_7031,N_6946,N_6987);
nand U7032 (N_7032,N_6949,N_6818);
or U7033 (N_7033,N_6988,N_6916);
nand U7034 (N_7034,N_6803,N_6893);
xor U7035 (N_7035,N_6951,N_6982);
nand U7036 (N_7036,N_6912,N_6825);
or U7037 (N_7037,N_6832,N_6840);
or U7038 (N_7038,N_6952,N_6927);
xnor U7039 (N_7039,N_6892,N_6990);
nand U7040 (N_7040,N_6938,N_6965);
xnor U7041 (N_7041,N_6998,N_6853);
or U7042 (N_7042,N_6816,N_6977);
and U7043 (N_7043,N_6948,N_6931);
and U7044 (N_7044,N_6876,N_6861);
and U7045 (N_7045,N_6864,N_6975);
or U7046 (N_7046,N_6996,N_6910);
nor U7047 (N_7047,N_6834,N_6937);
nand U7048 (N_7048,N_6800,N_6954);
or U7049 (N_7049,N_6896,N_6885);
or U7050 (N_7050,N_6843,N_6811);
or U7051 (N_7051,N_6809,N_6939);
nor U7052 (N_7052,N_6991,N_6824);
nor U7053 (N_7053,N_6936,N_6877);
or U7054 (N_7054,N_6979,N_6985);
and U7055 (N_7055,N_6808,N_6908);
xor U7056 (N_7056,N_6862,N_6923);
and U7057 (N_7057,N_6913,N_6958);
nor U7058 (N_7058,N_6941,N_6932);
nand U7059 (N_7059,N_6928,N_6964);
xnor U7060 (N_7060,N_6890,N_6879);
xor U7061 (N_7061,N_6960,N_6992);
or U7062 (N_7062,N_6994,N_6870);
or U7063 (N_7063,N_6953,N_6922);
or U7064 (N_7064,N_6866,N_6919);
xnor U7065 (N_7065,N_6929,N_6942);
or U7066 (N_7066,N_6945,N_6935);
and U7067 (N_7067,N_6924,N_6943);
or U7068 (N_7068,N_6966,N_6836);
nor U7069 (N_7069,N_6847,N_6934);
or U7070 (N_7070,N_6839,N_6969);
and U7071 (N_7071,N_6805,N_6995);
and U7072 (N_7072,N_6804,N_6868);
nand U7073 (N_7073,N_6947,N_6875);
xnor U7074 (N_7074,N_6973,N_6955);
nand U7075 (N_7075,N_6850,N_6884);
xor U7076 (N_7076,N_6933,N_6914);
nand U7077 (N_7077,N_6959,N_6918);
or U7078 (N_7078,N_6817,N_6903);
nand U7079 (N_7079,N_6859,N_6980);
nor U7080 (N_7080,N_6841,N_6869);
nand U7081 (N_7081,N_6860,N_6819);
nor U7082 (N_7082,N_6827,N_6970);
and U7083 (N_7083,N_6878,N_6968);
or U7084 (N_7084,N_6837,N_6801);
xor U7085 (N_7085,N_6911,N_6822);
or U7086 (N_7086,N_6871,N_6882);
nand U7087 (N_7087,N_6972,N_6880);
nand U7088 (N_7088,N_6854,N_6944);
nor U7089 (N_7089,N_6883,N_6971);
and U7090 (N_7090,N_6806,N_6905);
or U7091 (N_7091,N_6898,N_6894);
or U7092 (N_7092,N_6852,N_6930);
xnor U7093 (N_7093,N_6821,N_6895);
and U7094 (N_7094,N_6865,N_6920);
nor U7095 (N_7095,N_6957,N_6807);
nand U7096 (N_7096,N_6974,N_6833);
and U7097 (N_7097,N_6867,N_6848);
xor U7098 (N_7098,N_6926,N_6921);
nor U7099 (N_7099,N_6962,N_6986);
and U7100 (N_7100,N_6880,N_6858);
xor U7101 (N_7101,N_6968,N_6833);
nand U7102 (N_7102,N_6888,N_6944);
or U7103 (N_7103,N_6961,N_6809);
xor U7104 (N_7104,N_6842,N_6887);
nand U7105 (N_7105,N_6812,N_6965);
and U7106 (N_7106,N_6829,N_6899);
xnor U7107 (N_7107,N_6813,N_6921);
nand U7108 (N_7108,N_6989,N_6805);
nor U7109 (N_7109,N_6891,N_6905);
xor U7110 (N_7110,N_6939,N_6918);
and U7111 (N_7111,N_6973,N_6896);
and U7112 (N_7112,N_6954,N_6909);
and U7113 (N_7113,N_6928,N_6860);
nand U7114 (N_7114,N_6818,N_6959);
nand U7115 (N_7115,N_6866,N_6911);
or U7116 (N_7116,N_6804,N_6990);
and U7117 (N_7117,N_6888,N_6948);
or U7118 (N_7118,N_6836,N_6847);
and U7119 (N_7119,N_6897,N_6866);
and U7120 (N_7120,N_6890,N_6867);
or U7121 (N_7121,N_6971,N_6887);
and U7122 (N_7122,N_6964,N_6833);
or U7123 (N_7123,N_6958,N_6819);
nand U7124 (N_7124,N_6977,N_6825);
nand U7125 (N_7125,N_6838,N_6819);
or U7126 (N_7126,N_6961,N_6845);
nor U7127 (N_7127,N_6851,N_6816);
nand U7128 (N_7128,N_6967,N_6909);
nor U7129 (N_7129,N_6893,N_6831);
nor U7130 (N_7130,N_6905,N_6991);
xor U7131 (N_7131,N_6845,N_6841);
nor U7132 (N_7132,N_6823,N_6907);
or U7133 (N_7133,N_6964,N_6861);
or U7134 (N_7134,N_6964,N_6906);
or U7135 (N_7135,N_6948,N_6849);
and U7136 (N_7136,N_6865,N_6927);
xor U7137 (N_7137,N_6801,N_6910);
nand U7138 (N_7138,N_6962,N_6881);
and U7139 (N_7139,N_6959,N_6823);
and U7140 (N_7140,N_6857,N_6892);
nand U7141 (N_7141,N_6887,N_6995);
or U7142 (N_7142,N_6978,N_6824);
nor U7143 (N_7143,N_6967,N_6825);
or U7144 (N_7144,N_6929,N_6913);
nor U7145 (N_7145,N_6994,N_6968);
or U7146 (N_7146,N_6935,N_6894);
and U7147 (N_7147,N_6888,N_6800);
nand U7148 (N_7148,N_6884,N_6961);
nor U7149 (N_7149,N_6907,N_6810);
nand U7150 (N_7150,N_6972,N_6898);
and U7151 (N_7151,N_6880,N_6898);
nand U7152 (N_7152,N_6872,N_6983);
or U7153 (N_7153,N_6889,N_6846);
and U7154 (N_7154,N_6976,N_6845);
and U7155 (N_7155,N_6805,N_6900);
nand U7156 (N_7156,N_6955,N_6979);
nor U7157 (N_7157,N_6907,N_6846);
nand U7158 (N_7158,N_6974,N_6992);
nor U7159 (N_7159,N_6889,N_6854);
xor U7160 (N_7160,N_6987,N_6957);
nand U7161 (N_7161,N_6847,N_6999);
nor U7162 (N_7162,N_6929,N_6994);
nor U7163 (N_7163,N_6999,N_6861);
and U7164 (N_7164,N_6993,N_6992);
xnor U7165 (N_7165,N_6809,N_6844);
nand U7166 (N_7166,N_6894,N_6997);
xnor U7167 (N_7167,N_6916,N_6840);
or U7168 (N_7168,N_6887,N_6840);
or U7169 (N_7169,N_6896,N_6980);
and U7170 (N_7170,N_6987,N_6806);
and U7171 (N_7171,N_6841,N_6936);
nor U7172 (N_7172,N_6881,N_6912);
or U7173 (N_7173,N_6976,N_6954);
and U7174 (N_7174,N_6965,N_6861);
nand U7175 (N_7175,N_6870,N_6911);
or U7176 (N_7176,N_6814,N_6829);
nand U7177 (N_7177,N_6820,N_6967);
and U7178 (N_7178,N_6846,N_6927);
nand U7179 (N_7179,N_6933,N_6856);
nor U7180 (N_7180,N_6848,N_6906);
xor U7181 (N_7181,N_6826,N_6898);
xor U7182 (N_7182,N_6985,N_6819);
nand U7183 (N_7183,N_6871,N_6857);
nor U7184 (N_7184,N_6992,N_6912);
xor U7185 (N_7185,N_6952,N_6910);
and U7186 (N_7186,N_6989,N_6840);
and U7187 (N_7187,N_6857,N_6855);
nand U7188 (N_7188,N_6978,N_6974);
or U7189 (N_7189,N_6911,N_6815);
nand U7190 (N_7190,N_6997,N_6927);
xnor U7191 (N_7191,N_6800,N_6972);
nand U7192 (N_7192,N_6805,N_6962);
or U7193 (N_7193,N_6879,N_6972);
or U7194 (N_7194,N_6915,N_6858);
nand U7195 (N_7195,N_6853,N_6814);
or U7196 (N_7196,N_6872,N_6920);
nor U7197 (N_7197,N_6946,N_6847);
nor U7198 (N_7198,N_6992,N_6955);
nand U7199 (N_7199,N_6853,N_6848);
nor U7200 (N_7200,N_7016,N_7150);
and U7201 (N_7201,N_7000,N_7189);
and U7202 (N_7202,N_7097,N_7055);
or U7203 (N_7203,N_7138,N_7159);
or U7204 (N_7204,N_7176,N_7013);
nand U7205 (N_7205,N_7009,N_7023);
xor U7206 (N_7206,N_7123,N_7004);
xnor U7207 (N_7207,N_7056,N_7148);
nor U7208 (N_7208,N_7146,N_7114);
nand U7209 (N_7209,N_7128,N_7046);
and U7210 (N_7210,N_7188,N_7132);
nor U7211 (N_7211,N_7116,N_7145);
nand U7212 (N_7212,N_7048,N_7020);
or U7213 (N_7213,N_7126,N_7091);
xnor U7214 (N_7214,N_7036,N_7025);
xnor U7215 (N_7215,N_7119,N_7078);
xnor U7216 (N_7216,N_7038,N_7197);
or U7217 (N_7217,N_7089,N_7002);
nor U7218 (N_7218,N_7053,N_7101);
or U7219 (N_7219,N_7031,N_7037);
nor U7220 (N_7220,N_7198,N_7170);
nand U7221 (N_7221,N_7165,N_7017);
nand U7222 (N_7222,N_7155,N_7152);
nor U7223 (N_7223,N_7065,N_7098);
xor U7224 (N_7224,N_7105,N_7018);
nand U7225 (N_7225,N_7196,N_7158);
and U7226 (N_7226,N_7045,N_7085);
nor U7227 (N_7227,N_7066,N_7072);
and U7228 (N_7228,N_7083,N_7084);
and U7229 (N_7229,N_7094,N_7014);
nor U7230 (N_7230,N_7068,N_7006);
and U7231 (N_7231,N_7003,N_7069);
nand U7232 (N_7232,N_7092,N_7047);
and U7233 (N_7233,N_7051,N_7186);
nand U7234 (N_7234,N_7131,N_7130);
xnor U7235 (N_7235,N_7043,N_7054);
or U7236 (N_7236,N_7129,N_7193);
nor U7237 (N_7237,N_7007,N_7124);
nor U7238 (N_7238,N_7087,N_7040);
xnor U7239 (N_7239,N_7088,N_7133);
or U7240 (N_7240,N_7182,N_7183);
nand U7241 (N_7241,N_7154,N_7173);
xnor U7242 (N_7242,N_7113,N_7191);
nor U7243 (N_7243,N_7166,N_7112);
nor U7244 (N_7244,N_7100,N_7127);
or U7245 (N_7245,N_7027,N_7076);
nand U7246 (N_7246,N_7160,N_7140);
nand U7247 (N_7247,N_7093,N_7057);
and U7248 (N_7248,N_7095,N_7015);
or U7249 (N_7249,N_7174,N_7073);
or U7250 (N_7250,N_7103,N_7163);
nand U7251 (N_7251,N_7121,N_7178);
nor U7252 (N_7252,N_7029,N_7153);
and U7253 (N_7253,N_7010,N_7071);
or U7254 (N_7254,N_7139,N_7052);
nor U7255 (N_7255,N_7115,N_7192);
nand U7256 (N_7256,N_7172,N_7005);
or U7257 (N_7257,N_7134,N_7059);
and U7258 (N_7258,N_7108,N_7190);
nor U7259 (N_7259,N_7096,N_7177);
and U7260 (N_7260,N_7109,N_7110);
and U7261 (N_7261,N_7033,N_7194);
xor U7262 (N_7262,N_7157,N_7044);
and U7263 (N_7263,N_7164,N_7061);
nand U7264 (N_7264,N_7187,N_7080);
and U7265 (N_7265,N_7199,N_7136);
nand U7266 (N_7266,N_7077,N_7001);
nand U7267 (N_7267,N_7074,N_7167);
nor U7268 (N_7268,N_7032,N_7075);
nor U7269 (N_7269,N_7168,N_7070);
and U7270 (N_7270,N_7180,N_7021);
nand U7271 (N_7271,N_7060,N_7142);
and U7272 (N_7272,N_7117,N_7090);
xor U7273 (N_7273,N_7175,N_7034);
nand U7274 (N_7274,N_7049,N_7147);
and U7275 (N_7275,N_7107,N_7120);
xor U7276 (N_7276,N_7058,N_7008);
xnor U7277 (N_7277,N_7030,N_7099);
or U7278 (N_7278,N_7011,N_7185);
nand U7279 (N_7279,N_7019,N_7086);
xnor U7280 (N_7280,N_7028,N_7082);
and U7281 (N_7281,N_7181,N_7171);
and U7282 (N_7282,N_7151,N_7026);
nand U7283 (N_7283,N_7079,N_7122);
nor U7284 (N_7284,N_7039,N_7195);
or U7285 (N_7285,N_7135,N_7156);
nor U7286 (N_7286,N_7144,N_7042);
nor U7287 (N_7287,N_7081,N_7024);
and U7288 (N_7288,N_7067,N_7106);
nand U7289 (N_7289,N_7118,N_7063);
and U7290 (N_7290,N_7141,N_7179);
nor U7291 (N_7291,N_7022,N_7102);
nor U7292 (N_7292,N_7184,N_7050);
nand U7293 (N_7293,N_7035,N_7137);
or U7294 (N_7294,N_7169,N_7143);
and U7295 (N_7295,N_7041,N_7162);
or U7296 (N_7296,N_7104,N_7149);
nor U7297 (N_7297,N_7125,N_7111);
nor U7298 (N_7298,N_7161,N_7012);
or U7299 (N_7299,N_7064,N_7062);
nand U7300 (N_7300,N_7167,N_7020);
xnor U7301 (N_7301,N_7003,N_7031);
nand U7302 (N_7302,N_7144,N_7136);
or U7303 (N_7303,N_7045,N_7016);
nand U7304 (N_7304,N_7172,N_7097);
and U7305 (N_7305,N_7052,N_7101);
and U7306 (N_7306,N_7164,N_7120);
and U7307 (N_7307,N_7102,N_7174);
or U7308 (N_7308,N_7100,N_7168);
and U7309 (N_7309,N_7017,N_7019);
xor U7310 (N_7310,N_7115,N_7152);
nand U7311 (N_7311,N_7081,N_7174);
or U7312 (N_7312,N_7082,N_7177);
nand U7313 (N_7313,N_7118,N_7169);
xor U7314 (N_7314,N_7062,N_7104);
and U7315 (N_7315,N_7033,N_7021);
nand U7316 (N_7316,N_7149,N_7084);
xnor U7317 (N_7317,N_7084,N_7145);
and U7318 (N_7318,N_7189,N_7152);
xnor U7319 (N_7319,N_7166,N_7061);
and U7320 (N_7320,N_7002,N_7061);
nor U7321 (N_7321,N_7100,N_7193);
or U7322 (N_7322,N_7046,N_7103);
nand U7323 (N_7323,N_7145,N_7175);
nand U7324 (N_7324,N_7057,N_7160);
and U7325 (N_7325,N_7058,N_7046);
nor U7326 (N_7326,N_7043,N_7045);
xor U7327 (N_7327,N_7114,N_7095);
xor U7328 (N_7328,N_7079,N_7006);
and U7329 (N_7329,N_7017,N_7104);
xor U7330 (N_7330,N_7028,N_7040);
nor U7331 (N_7331,N_7086,N_7131);
and U7332 (N_7332,N_7003,N_7100);
nor U7333 (N_7333,N_7160,N_7106);
nand U7334 (N_7334,N_7055,N_7194);
xnor U7335 (N_7335,N_7049,N_7175);
or U7336 (N_7336,N_7034,N_7040);
and U7337 (N_7337,N_7120,N_7025);
or U7338 (N_7338,N_7052,N_7034);
nor U7339 (N_7339,N_7176,N_7101);
and U7340 (N_7340,N_7197,N_7099);
and U7341 (N_7341,N_7001,N_7123);
nand U7342 (N_7342,N_7170,N_7086);
or U7343 (N_7343,N_7033,N_7196);
xor U7344 (N_7344,N_7092,N_7124);
and U7345 (N_7345,N_7022,N_7067);
or U7346 (N_7346,N_7107,N_7104);
nor U7347 (N_7347,N_7018,N_7008);
and U7348 (N_7348,N_7056,N_7121);
or U7349 (N_7349,N_7008,N_7075);
nand U7350 (N_7350,N_7199,N_7170);
nor U7351 (N_7351,N_7147,N_7080);
xnor U7352 (N_7352,N_7133,N_7029);
or U7353 (N_7353,N_7104,N_7015);
nor U7354 (N_7354,N_7117,N_7095);
nand U7355 (N_7355,N_7081,N_7047);
and U7356 (N_7356,N_7123,N_7184);
and U7357 (N_7357,N_7186,N_7177);
or U7358 (N_7358,N_7023,N_7074);
xor U7359 (N_7359,N_7175,N_7123);
or U7360 (N_7360,N_7017,N_7103);
nand U7361 (N_7361,N_7190,N_7184);
nand U7362 (N_7362,N_7164,N_7025);
nand U7363 (N_7363,N_7166,N_7092);
nand U7364 (N_7364,N_7159,N_7015);
nand U7365 (N_7365,N_7044,N_7133);
nor U7366 (N_7366,N_7095,N_7059);
and U7367 (N_7367,N_7197,N_7020);
nand U7368 (N_7368,N_7152,N_7120);
and U7369 (N_7369,N_7035,N_7075);
nand U7370 (N_7370,N_7039,N_7084);
nand U7371 (N_7371,N_7028,N_7180);
xor U7372 (N_7372,N_7008,N_7041);
nor U7373 (N_7373,N_7068,N_7173);
xnor U7374 (N_7374,N_7092,N_7031);
nand U7375 (N_7375,N_7199,N_7153);
xor U7376 (N_7376,N_7056,N_7025);
xor U7377 (N_7377,N_7133,N_7061);
nand U7378 (N_7378,N_7073,N_7143);
or U7379 (N_7379,N_7182,N_7185);
nand U7380 (N_7380,N_7169,N_7013);
nand U7381 (N_7381,N_7036,N_7114);
nand U7382 (N_7382,N_7139,N_7189);
and U7383 (N_7383,N_7195,N_7032);
or U7384 (N_7384,N_7125,N_7183);
xnor U7385 (N_7385,N_7173,N_7166);
xnor U7386 (N_7386,N_7079,N_7167);
nand U7387 (N_7387,N_7160,N_7168);
nand U7388 (N_7388,N_7056,N_7125);
nand U7389 (N_7389,N_7022,N_7170);
xnor U7390 (N_7390,N_7073,N_7118);
or U7391 (N_7391,N_7127,N_7105);
nand U7392 (N_7392,N_7009,N_7107);
nor U7393 (N_7393,N_7127,N_7031);
or U7394 (N_7394,N_7001,N_7103);
and U7395 (N_7395,N_7113,N_7099);
xor U7396 (N_7396,N_7115,N_7084);
xnor U7397 (N_7397,N_7169,N_7119);
or U7398 (N_7398,N_7109,N_7160);
nor U7399 (N_7399,N_7148,N_7199);
and U7400 (N_7400,N_7259,N_7345);
and U7401 (N_7401,N_7313,N_7231);
nand U7402 (N_7402,N_7241,N_7206);
xor U7403 (N_7403,N_7242,N_7326);
or U7404 (N_7404,N_7342,N_7220);
nand U7405 (N_7405,N_7325,N_7244);
and U7406 (N_7406,N_7232,N_7217);
nand U7407 (N_7407,N_7224,N_7304);
nor U7408 (N_7408,N_7356,N_7370);
nor U7409 (N_7409,N_7260,N_7350);
or U7410 (N_7410,N_7391,N_7229);
xor U7411 (N_7411,N_7211,N_7362);
nor U7412 (N_7412,N_7389,N_7317);
nand U7413 (N_7413,N_7215,N_7392);
xnor U7414 (N_7414,N_7296,N_7337);
and U7415 (N_7415,N_7385,N_7340);
and U7416 (N_7416,N_7324,N_7344);
or U7417 (N_7417,N_7388,N_7276);
nor U7418 (N_7418,N_7280,N_7249);
and U7419 (N_7419,N_7390,N_7332);
or U7420 (N_7420,N_7357,N_7387);
or U7421 (N_7421,N_7247,N_7334);
xor U7422 (N_7422,N_7222,N_7289);
nand U7423 (N_7423,N_7251,N_7219);
or U7424 (N_7424,N_7310,N_7360);
xor U7425 (N_7425,N_7363,N_7381);
nor U7426 (N_7426,N_7286,N_7393);
nand U7427 (N_7427,N_7268,N_7203);
nand U7428 (N_7428,N_7282,N_7308);
nor U7429 (N_7429,N_7207,N_7369);
and U7430 (N_7430,N_7298,N_7266);
or U7431 (N_7431,N_7278,N_7394);
nand U7432 (N_7432,N_7293,N_7380);
xor U7433 (N_7433,N_7361,N_7399);
nand U7434 (N_7434,N_7300,N_7267);
and U7435 (N_7435,N_7287,N_7255);
and U7436 (N_7436,N_7378,N_7228);
xor U7437 (N_7437,N_7314,N_7398);
nand U7438 (N_7438,N_7281,N_7265);
nand U7439 (N_7439,N_7352,N_7386);
nand U7440 (N_7440,N_7238,N_7351);
nand U7441 (N_7441,N_7234,N_7301);
or U7442 (N_7442,N_7320,N_7239);
nand U7443 (N_7443,N_7226,N_7302);
nand U7444 (N_7444,N_7285,N_7273);
or U7445 (N_7445,N_7376,N_7318);
nand U7446 (N_7446,N_7316,N_7258);
nand U7447 (N_7447,N_7223,N_7240);
nor U7448 (N_7448,N_7327,N_7322);
or U7449 (N_7449,N_7384,N_7292);
xnor U7450 (N_7450,N_7372,N_7303);
or U7451 (N_7451,N_7227,N_7210);
and U7452 (N_7452,N_7323,N_7218);
nand U7453 (N_7453,N_7377,N_7257);
and U7454 (N_7454,N_7395,N_7269);
or U7455 (N_7455,N_7359,N_7338);
and U7456 (N_7456,N_7306,N_7335);
xnor U7457 (N_7457,N_7262,N_7201);
xor U7458 (N_7458,N_7382,N_7353);
or U7459 (N_7459,N_7290,N_7216);
and U7460 (N_7460,N_7274,N_7321);
nor U7461 (N_7461,N_7271,N_7339);
nor U7462 (N_7462,N_7264,N_7270);
xnor U7463 (N_7463,N_7277,N_7250);
and U7464 (N_7464,N_7364,N_7374);
nand U7465 (N_7465,N_7230,N_7295);
nand U7466 (N_7466,N_7346,N_7319);
and U7467 (N_7467,N_7202,N_7371);
nor U7468 (N_7468,N_7213,N_7383);
nor U7469 (N_7469,N_7225,N_7256);
or U7470 (N_7470,N_7365,N_7397);
xnor U7471 (N_7471,N_7212,N_7275);
nor U7472 (N_7472,N_7272,N_7328);
nand U7473 (N_7473,N_7311,N_7243);
and U7474 (N_7474,N_7307,N_7330);
nor U7475 (N_7475,N_7341,N_7348);
and U7476 (N_7476,N_7305,N_7288);
and U7477 (N_7477,N_7373,N_7294);
and U7478 (N_7478,N_7375,N_7245);
nor U7479 (N_7479,N_7253,N_7235);
or U7480 (N_7480,N_7297,N_7208);
nand U7481 (N_7481,N_7236,N_7205);
nor U7482 (N_7482,N_7366,N_7248);
xnor U7483 (N_7483,N_7200,N_7355);
or U7484 (N_7484,N_7261,N_7349);
nand U7485 (N_7485,N_7396,N_7291);
or U7486 (N_7486,N_7263,N_7309);
nor U7487 (N_7487,N_7315,N_7336);
nor U7488 (N_7488,N_7214,N_7368);
and U7489 (N_7489,N_7283,N_7312);
and U7490 (N_7490,N_7299,N_7254);
nor U7491 (N_7491,N_7221,N_7333);
nand U7492 (N_7492,N_7233,N_7252);
nand U7493 (N_7493,N_7284,N_7358);
and U7494 (N_7494,N_7347,N_7354);
and U7495 (N_7495,N_7343,N_7237);
xnor U7496 (N_7496,N_7367,N_7204);
nor U7497 (N_7497,N_7379,N_7329);
or U7498 (N_7498,N_7246,N_7279);
or U7499 (N_7499,N_7331,N_7209);
or U7500 (N_7500,N_7291,N_7387);
nor U7501 (N_7501,N_7369,N_7210);
nor U7502 (N_7502,N_7215,N_7345);
xnor U7503 (N_7503,N_7350,N_7373);
nand U7504 (N_7504,N_7215,N_7393);
or U7505 (N_7505,N_7344,N_7377);
xnor U7506 (N_7506,N_7337,N_7329);
xor U7507 (N_7507,N_7213,N_7275);
and U7508 (N_7508,N_7238,N_7212);
nor U7509 (N_7509,N_7251,N_7241);
and U7510 (N_7510,N_7299,N_7360);
or U7511 (N_7511,N_7266,N_7299);
and U7512 (N_7512,N_7256,N_7279);
nand U7513 (N_7513,N_7320,N_7215);
or U7514 (N_7514,N_7309,N_7240);
xnor U7515 (N_7515,N_7316,N_7383);
nor U7516 (N_7516,N_7247,N_7390);
and U7517 (N_7517,N_7346,N_7241);
or U7518 (N_7518,N_7389,N_7289);
or U7519 (N_7519,N_7269,N_7223);
or U7520 (N_7520,N_7271,N_7231);
xnor U7521 (N_7521,N_7338,N_7304);
nor U7522 (N_7522,N_7345,N_7285);
xnor U7523 (N_7523,N_7314,N_7350);
or U7524 (N_7524,N_7394,N_7214);
or U7525 (N_7525,N_7338,N_7332);
nor U7526 (N_7526,N_7375,N_7324);
xor U7527 (N_7527,N_7336,N_7333);
xnor U7528 (N_7528,N_7375,N_7207);
xor U7529 (N_7529,N_7227,N_7390);
nor U7530 (N_7530,N_7305,N_7345);
nor U7531 (N_7531,N_7317,N_7229);
nor U7532 (N_7532,N_7314,N_7343);
nor U7533 (N_7533,N_7292,N_7259);
nand U7534 (N_7534,N_7362,N_7262);
nand U7535 (N_7535,N_7388,N_7313);
and U7536 (N_7536,N_7339,N_7212);
xor U7537 (N_7537,N_7311,N_7323);
nor U7538 (N_7538,N_7301,N_7342);
and U7539 (N_7539,N_7294,N_7262);
nor U7540 (N_7540,N_7273,N_7342);
nor U7541 (N_7541,N_7341,N_7301);
or U7542 (N_7542,N_7335,N_7290);
nand U7543 (N_7543,N_7360,N_7324);
or U7544 (N_7544,N_7258,N_7238);
nand U7545 (N_7545,N_7223,N_7253);
or U7546 (N_7546,N_7348,N_7227);
nor U7547 (N_7547,N_7388,N_7230);
and U7548 (N_7548,N_7322,N_7285);
nand U7549 (N_7549,N_7256,N_7211);
nand U7550 (N_7550,N_7212,N_7273);
nand U7551 (N_7551,N_7297,N_7364);
and U7552 (N_7552,N_7344,N_7268);
nor U7553 (N_7553,N_7353,N_7296);
xnor U7554 (N_7554,N_7346,N_7234);
nand U7555 (N_7555,N_7359,N_7330);
nand U7556 (N_7556,N_7301,N_7339);
or U7557 (N_7557,N_7258,N_7341);
nand U7558 (N_7558,N_7228,N_7279);
nor U7559 (N_7559,N_7239,N_7280);
or U7560 (N_7560,N_7335,N_7242);
nor U7561 (N_7561,N_7331,N_7346);
nand U7562 (N_7562,N_7204,N_7305);
xor U7563 (N_7563,N_7303,N_7275);
xnor U7564 (N_7564,N_7391,N_7223);
or U7565 (N_7565,N_7239,N_7395);
and U7566 (N_7566,N_7229,N_7319);
and U7567 (N_7567,N_7272,N_7310);
xor U7568 (N_7568,N_7209,N_7213);
and U7569 (N_7569,N_7229,N_7348);
and U7570 (N_7570,N_7238,N_7333);
and U7571 (N_7571,N_7288,N_7314);
nor U7572 (N_7572,N_7348,N_7294);
and U7573 (N_7573,N_7329,N_7384);
xnor U7574 (N_7574,N_7246,N_7234);
or U7575 (N_7575,N_7319,N_7306);
nand U7576 (N_7576,N_7335,N_7337);
xnor U7577 (N_7577,N_7225,N_7317);
nor U7578 (N_7578,N_7299,N_7237);
nand U7579 (N_7579,N_7227,N_7397);
or U7580 (N_7580,N_7290,N_7377);
nand U7581 (N_7581,N_7399,N_7232);
and U7582 (N_7582,N_7205,N_7265);
nor U7583 (N_7583,N_7252,N_7315);
xnor U7584 (N_7584,N_7334,N_7235);
xnor U7585 (N_7585,N_7221,N_7289);
xor U7586 (N_7586,N_7201,N_7270);
nor U7587 (N_7587,N_7374,N_7205);
nand U7588 (N_7588,N_7305,N_7290);
and U7589 (N_7589,N_7259,N_7355);
nand U7590 (N_7590,N_7228,N_7332);
xor U7591 (N_7591,N_7226,N_7368);
and U7592 (N_7592,N_7275,N_7255);
and U7593 (N_7593,N_7236,N_7381);
or U7594 (N_7594,N_7384,N_7217);
nand U7595 (N_7595,N_7275,N_7344);
or U7596 (N_7596,N_7236,N_7347);
xor U7597 (N_7597,N_7340,N_7355);
or U7598 (N_7598,N_7236,N_7340);
xor U7599 (N_7599,N_7379,N_7371);
nor U7600 (N_7600,N_7493,N_7462);
nand U7601 (N_7601,N_7486,N_7439);
xor U7602 (N_7602,N_7430,N_7468);
nand U7603 (N_7603,N_7572,N_7434);
and U7604 (N_7604,N_7504,N_7455);
nor U7605 (N_7605,N_7470,N_7573);
xnor U7606 (N_7606,N_7511,N_7509);
xnor U7607 (N_7607,N_7526,N_7551);
xor U7608 (N_7608,N_7413,N_7458);
nor U7609 (N_7609,N_7409,N_7593);
nand U7610 (N_7610,N_7587,N_7424);
xnor U7611 (N_7611,N_7448,N_7412);
or U7612 (N_7612,N_7549,N_7418);
or U7613 (N_7613,N_7563,N_7422);
xnor U7614 (N_7614,N_7447,N_7483);
nand U7615 (N_7615,N_7508,N_7461);
nand U7616 (N_7616,N_7442,N_7459);
and U7617 (N_7617,N_7568,N_7479);
and U7618 (N_7618,N_7579,N_7474);
and U7619 (N_7619,N_7534,N_7535);
xnor U7620 (N_7620,N_7516,N_7583);
or U7621 (N_7621,N_7471,N_7499);
or U7622 (N_7622,N_7543,N_7564);
nor U7623 (N_7623,N_7469,N_7420);
nand U7624 (N_7624,N_7557,N_7585);
and U7625 (N_7625,N_7419,N_7555);
nor U7626 (N_7626,N_7435,N_7599);
xnor U7627 (N_7627,N_7530,N_7597);
nand U7628 (N_7628,N_7438,N_7408);
or U7629 (N_7629,N_7506,N_7497);
nand U7630 (N_7630,N_7494,N_7488);
xnor U7631 (N_7631,N_7500,N_7533);
and U7632 (N_7632,N_7431,N_7503);
or U7633 (N_7633,N_7580,N_7481);
nor U7634 (N_7634,N_7432,N_7539);
and U7635 (N_7635,N_7528,N_7514);
or U7636 (N_7636,N_7498,N_7417);
nor U7637 (N_7637,N_7510,N_7480);
xor U7638 (N_7638,N_7570,N_7426);
and U7639 (N_7639,N_7571,N_7450);
or U7640 (N_7640,N_7445,N_7490);
nor U7641 (N_7641,N_7589,N_7495);
or U7642 (N_7642,N_7524,N_7505);
nand U7643 (N_7643,N_7519,N_7496);
or U7644 (N_7644,N_7513,N_7405);
nor U7645 (N_7645,N_7478,N_7460);
xnor U7646 (N_7646,N_7556,N_7591);
and U7647 (N_7647,N_7536,N_7598);
nor U7648 (N_7648,N_7404,N_7429);
nor U7649 (N_7649,N_7565,N_7561);
xor U7650 (N_7650,N_7559,N_7440);
or U7651 (N_7651,N_7415,N_7457);
and U7652 (N_7652,N_7521,N_7552);
nand U7653 (N_7653,N_7473,N_7451);
and U7654 (N_7654,N_7428,N_7423);
xor U7655 (N_7655,N_7523,N_7464);
xnor U7656 (N_7656,N_7581,N_7522);
or U7657 (N_7657,N_7548,N_7444);
xor U7658 (N_7658,N_7578,N_7425);
and U7659 (N_7659,N_7406,N_7463);
or U7660 (N_7660,N_7416,N_7537);
nand U7661 (N_7661,N_7436,N_7595);
and U7662 (N_7662,N_7515,N_7437);
and U7663 (N_7663,N_7454,N_7553);
or U7664 (N_7664,N_7512,N_7544);
or U7665 (N_7665,N_7465,N_7575);
xnor U7666 (N_7666,N_7540,N_7421);
or U7667 (N_7667,N_7584,N_7402);
xor U7668 (N_7668,N_7433,N_7401);
nand U7669 (N_7669,N_7586,N_7577);
and U7670 (N_7670,N_7531,N_7485);
xor U7671 (N_7671,N_7476,N_7452);
nor U7672 (N_7672,N_7525,N_7547);
nor U7673 (N_7673,N_7542,N_7492);
nand U7674 (N_7674,N_7567,N_7507);
xor U7675 (N_7675,N_7592,N_7517);
xnor U7676 (N_7676,N_7520,N_7554);
xnor U7677 (N_7677,N_7472,N_7518);
nor U7678 (N_7678,N_7538,N_7594);
xor U7679 (N_7679,N_7569,N_7491);
and U7680 (N_7680,N_7482,N_7501);
nor U7681 (N_7681,N_7456,N_7446);
and U7682 (N_7682,N_7441,N_7414);
or U7683 (N_7683,N_7532,N_7558);
xor U7684 (N_7684,N_7443,N_7582);
xnor U7685 (N_7685,N_7502,N_7562);
or U7686 (N_7686,N_7487,N_7588);
nand U7687 (N_7687,N_7467,N_7576);
xor U7688 (N_7688,N_7560,N_7484);
xor U7689 (N_7689,N_7590,N_7407);
nand U7690 (N_7690,N_7453,N_7477);
and U7691 (N_7691,N_7411,N_7449);
or U7692 (N_7692,N_7489,N_7545);
nor U7693 (N_7693,N_7403,N_7529);
and U7694 (N_7694,N_7541,N_7427);
nand U7695 (N_7695,N_7566,N_7475);
xnor U7696 (N_7696,N_7466,N_7546);
nand U7697 (N_7697,N_7410,N_7527);
and U7698 (N_7698,N_7550,N_7400);
nand U7699 (N_7699,N_7574,N_7596);
xnor U7700 (N_7700,N_7561,N_7440);
xnor U7701 (N_7701,N_7478,N_7518);
nor U7702 (N_7702,N_7584,N_7416);
or U7703 (N_7703,N_7571,N_7471);
or U7704 (N_7704,N_7417,N_7486);
or U7705 (N_7705,N_7524,N_7494);
nor U7706 (N_7706,N_7498,N_7596);
and U7707 (N_7707,N_7527,N_7481);
nor U7708 (N_7708,N_7524,N_7569);
xor U7709 (N_7709,N_7552,N_7537);
nor U7710 (N_7710,N_7406,N_7422);
nor U7711 (N_7711,N_7454,N_7501);
nand U7712 (N_7712,N_7526,N_7527);
xnor U7713 (N_7713,N_7528,N_7497);
nor U7714 (N_7714,N_7546,N_7403);
and U7715 (N_7715,N_7514,N_7429);
and U7716 (N_7716,N_7573,N_7508);
xor U7717 (N_7717,N_7556,N_7453);
nand U7718 (N_7718,N_7587,N_7446);
and U7719 (N_7719,N_7550,N_7590);
and U7720 (N_7720,N_7538,N_7540);
nor U7721 (N_7721,N_7543,N_7516);
or U7722 (N_7722,N_7469,N_7514);
nor U7723 (N_7723,N_7480,N_7573);
nor U7724 (N_7724,N_7500,N_7420);
xor U7725 (N_7725,N_7500,N_7547);
or U7726 (N_7726,N_7526,N_7508);
and U7727 (N_7727,N_7599,N_7433);
nor U7728 (N_7728,N_7452,N_7403);
and U7729 (N_7729,N_7584,N_7510);
and U7730 (N_7730,N_7542,N_7543);
xnor U7731 (N_7731,N_7449,N_7513);
nor U7732 (N_7732,N_7465,N_7419);
and U7733 (N_7733,N_7453,N_7504);
xor U7734 (N_7734,N_7437,N_7596);
and U7735 (N_7735,N_7466,N_7428);
and U7736 (N_7736,N_7495,N_7574);
nand U7737 (N_7737,N_7550,N_7527);
xnor U7738 (N_7738,N_7475,N_7560);
nand U7739 (N_7739,N_7555,N_7553);
nor U7740 (N_7740,N_7505,N_7514);
and U7741 (N_7741,N_7561,N_7539);
xnor U7742 (N_7742,N_7527,N_7596);
nand U7743 (N_7743,N_7454,N_7477);
and U7744 (N_7744,N_7599,N_7441);
or U7745 (N_7745,N_7496,N_7557);
nand U7746 (N_7746,N_7596,N_7416);
xor U7747 (N_7747,N_7419,N_7550);
or U7748 (N_7748,N_7436,N_7501);
nand U7749 (N_7749,N_7551,N_7566);
and U7750 (N_7750,N_7495,N_7448);
nor U7751 (N_7751,N_7411,N_7557);
nand U7752 (N_7752,N_7437,N_7426);
nor U7753 (N_7753,N_7421,N_7483);
and U7754 (N_7754,N_7508,N_7547);
nor U7755 (N_7755,N_7498,N_7582);
or U7756 (N_7756,N_7405,N_7467);
or U7757 (N_7757,N_7531,N_7522);
and U7758 (N_7758,N_7531,N_7464);
or U7759 (N_7759,N_7436,N_7442);
nand U7760 (N_7760,N_7518,N_7591);
xor U7761 (N_7761,N_7499,N_7567);
nor U7762 (N_7762,N_7561,N_7568);
nor U7763 (N_7763,N_7523,N_7447);
and U7764 (N_7764,N_7444,N_7457);
nand U7765 (N_7765,N_7456,N_7408);
or U7766 (N_7766,N_7590,N_7483);
nor U7767 (N_7767,N_7433,N_7499);
nor U7768 (N_7768,N_7479,N_7592);
xnor U7769 (N_7769,N_7428,N_7554);
or U7770 (N_7770,N_7563,N_7455);
nor U7771 (N_7771,N_7500,N_7540);
and U7772 (N_7772,N_7554,N_7513);
xnor U7773 (N_7773,N_7439,N_7459);
nor U7774 (N_7774,N_7401,N_7563);
or U7775 (N_7775,N_7567,N_7446);
or U7776 (N_7776,N_7591,N_7499);
and U7777 (N_7777,N_7590,N_7463);
nand U7778 (N_7778,N_7538,N_7544);
nand U7779 (N_7779,N_7435,N_7560);
and U7780 (N_7780,N_7532,N_7501);
nor U7781 (N_7781,N_7499,N_7490);
nor U7782 (N_7782,N_7593,N_7535);
nand U7783 (N_7783,N_7536,N_7447);
nor U7784 (N_7784,N_7437,N_7471);
nand U7785 (N_7785,N_7545,N_7566);
nor U7786 (N_7786,N_7405,N_7484);
nor U7787 (N_7787,N_7585,N_7590);
and U7788 (N_7788,N_7565,N_7513);
or U7789 (N_7789,N_7564,N_7460);
and U7790 (N_7790,N_7489,N_7512);
nor U7791 (N_7791,N_7581,N_7420);
nor U7792 (N_7792,N_7411,N_7474);
or U7793 (N_7793,N_7420,N_7463);
and U7794 (N_7794,N_7435,N_7497);
and U7795 (N_7795,N_7557,N_7433);
nand U7796 (N_7796,N_7457,N_7423);
nor U7797 (N_7797,N_7424,N_7533);
nand U7798 (N_7798,N_7470,N_7405);
or U7799 (N_7799,N_7548,N_7578);
and U7800 (N_7800,N_7626,N_7632);
or U7801 (N_7801,N_7610,N_7756);
nand U7802 (N_7802,N_7717,N_7712);
nand U7803 (N_7803,N_7676,N_7746);
or U7804 (N_7804,N_7662,N_7609);
xnor U7805 (N_7805,N_7741,N_7691);
nand U7806 (N_7806,N_7702,N_7661);
nand U7807 (N_7807,N_7674,N_7792);
xor U7808 (N_7808,N_7638,N_7736);
or U7809 (N_7809,N_7726,N_7605);
or U7810 (N_7810,N_7640,N_7666);
nand U7811 (N_7811,N_7635,N_7724);
xor U7812 (N_7812,N_7625,N_7647);
xnor U7813 (N_7813,N_7716,N_7754);
or U7814 (N_7814,N_7630,N_7644);
or U7815 (N_7815,N_7789,N_7732);
and U7816 (N_7816,N_7657,N_7782);
and U7817 (N_7817,N_7739,N_7688);
nor U7818 (N_7818,N_7650,N_7779);
or U7819 (N_7819,N_7670,N_7759);
or U7820 (N_7820,N_7672,N_7678);
nand U7821 (N_7821,N_7682,N_7614);
nand U7822 (N_7822,N_7667,N_7668);
nand U7823 (N_7823,N_7757,N_7663);
nand U7824 (N_7824,N_7737,N_7633);
and U7825 (N_7825,N_7745,N_7677);
nand U7826 (N_7826,N_7786,N_7752);
nor U7827 (N_7827,N_7761,N_7783);
or U7828 (N_7828,N_7725,N_7748);
and U7829 (N_7829,N_7671,N_7664);
xnor U7830 (N_7830,N_7606,N_7619);
xnor U7831 (N_7831,N_7784,N_7623);
xor U7832 (N_7832,N_7794,N_7721);
or U7833 (N_7833,N_7781,N_7772);
or U7834 (N_7834,N_7639,N_7718);
or U7835 (N_7835,N_7695,N_7699);
nand U7836 (N_7836,N_7648,N_7613);
or U7837 (N_7837,N_7627,N_7715);
or U7838 (N_7838,N_7618,N_7655);
nor U7839 (N_7839,N_7747,N_7774);
and U7840 (N_7840,N_7649,N_7767);
xnor U7841 (N_7841,N_7766,N_7637);
and U7842 (N_7842,N_7730,N_7686);
and U7843 (N_7843,N_7628,N_7771);
nand U7844 (N_7844,N_7673,N_7773);
xor U7845 (N_7845,N_7685,N_7616);
nand U7846 (N_7846,N_7742,N_7777);
nand U7847 (N_7847,N_7796,N_7762);
nand U7848 (N_7848,N_7753,N_7793);
and U7849 (N_7849,N_7653,N_7645);
or U7850 (N_7850,N_7646,N_7621);
nor U7851 (N_7851,N_7642,N_7634);
nor U7852 (N_7852,N_7776,N_7780);
xor U7853 (N_7853,N_7778,N_7760);
nand U7854 (N_7854,N_7681,N_7768);
nand U7855 (N_7855,N_7751,N_7624);
and U7856 (N_7856,N_7602,N_7683);
and U7857 (N_7857,N_7693,N_7600);
nand U7858 (N_7858,N_7641,N_7790);
and U7859 (N_7859,N_7675,N_7797);
nor U7860 (N_7860,N_7665,N_7728);
and U7861 (N_7861,N_7679,N_7798);
nor U7862 (N_7862,N_7744,N_7651);
or U7863 (N_7863,N_7775,N_7604);
xor U7864 (N_7864,N_7740,N_7722);
nand U7865 (N_7865,N_7710,N_7701);
nand U7866 (N_7866,N_7692,N_7622);
and U7867 (N_7867,N_7659,N_7652);
and U7868 (N_7868,N_7603,N_7601);
nand U7869 (N_7869,N_7731,N_7631);
and U7870 (N_7870,N_7764,N_7755);
and U7871 (N_7871,N_7660,N_7749);
xor U7872 (N_7872,N_7763,N_7611);
xnor U7873 (N_7873,N_7629,N_7791);
xnor U7874 (N_7874,N_7709,N_7788);
and U7875 (N_7875,N_7708,N_7696);
nor U7876 (N_7876,N_7656,N_7758);
or U7877 (N_7877,N_7711,N_7684);
nor U7878 (N_7878,N_7694,N_7615);
or U7879 (N_7879,N_7727,N_7795);
nor U7880 (N_7880,N_7735,N_7607);
and U7881 (N_7881,N_7706,N_7720);
and U7882 (N_7882,N_7680,N_7643);
xor U7883 (N_7883,N_7698,N_7787);
nand U7884 (N_7884,N_7707,N_7719);
nor U7885 (N_7885,N_7723,N_7705);
nand U7886 (N_7886,N_7750,N_7769);
nor U7887 (N_7887,N_7765,N_7697);
nor U7888 (N_7888,N_7617,N_7669);
nor U7889 (N_7889,N_7714,N_7636);
xnor U7890 (N_7890,N_7654,N_7785);
or U7891 (N_7891,N_7704,N_7687);
xor U7892 (N_7892,N_7658,N_7700);
or U7893 (N_7893,N_7612,N_7608);
or U7894 (N_7894,N_7689,N_7743);
or U7895 (N_7895,N_7713,N_7703);
or U7896 (N_7896,N_7729,N_7733);
nand U7897 (N_7897,N_7799,N_7690);
or U7898 (N_7898,N_7738,N_7770);
and U7899 (N_7899,N_7734,N_7620);
or U7900 (N_7900,N_7645,N_7765);
nor U7901 (N_7901,N_7648,N_7787);
xnor U7902 (N_7902,N_7671,N_7772);
nor U7903 (N_7903,N_7703,N_7643);
and U7904 (N_7904,N_7730,N_7618);
nand U7905 (N_7905,N_7743,N_7710);
nand U7906 (N_7906,N_7763,N_7653);
nand U7907 (N_7907,N_7780,N_7721);
or U7908 (N_7908,N_7768,N_7773);
nand U7909 (N_7909,N_7737,N_7724);
xnor U7910 (N_7910,N_7622,N_7752);
nor U7911 (N_7911,N_7609,N_7685);
nand U7912 (N_7912,N_7619,N_7784);
nand U7913 (N_7913,N_7796,N_7696);
nor U7914 (N_7914,N_7724,N_7758);
nand U7915 (N_7915,N_7605,N_7759);
nor U7916 (N_7916,N_7709,N_7658);
nand U7917 (N_7917,N_7797,N_7677);
xor U7918 (N_7918,N_7677,N_7641);
xor U7919 (N_7919,N_7703,N_7756);
nor U7920 (N_7920,N_7687,N_7660);
nor U7921 (N_7921,N_7723,N_7751);
nand U7922 (N_7922,N_7675,N_7763);
xnor U7923 (N_7923,N_7784,N_7728);
nand U7924 (N_7924,N_7726,N_7724);
nand U7925 (N_7925,N_7752,N_7669);
or U7926 (N_7926,N_7783,N_7615);
xnor U7927 (N_7927,N_7668,N_7739);
and U7928 (N_7928,N_7629,N_7755);
xnor U7929 (N_7929,N_7795,N_7758);
nand U7930 (N_7930,N_7719,N_7717);
nand U7931 (N_7931,N_7652,N_7727);
xnor U7932 (N_7932,N_7633,N_7729);
or U7933 (N_7933,N_7612,N_7722);
or U7934 (N_7934,N_7794,N_7684);
nor U7935 (N_7935,N_7776,N_7797);
nand U7936 (N_7936,N_7715,N_7757);
or U7937 (N_7937,N_7645,N_7710);
xnor U7938 (N_7938,N_7684,N_7657);
and U7939 (N_7939,N_7744,N_7720);
nor U7940 (N_7940,N_7613,N_7684);
or U7941 (N_7941,N_7786,N_7612);
or U7942 (N_7942,N_7755,N_7643);
nor U7943 (N_7943,N_7646,N_7716);
and U7944 (N_7944,N_7765,N_7647);
nor U7945 (N_7945,N_7762,N_7637);
or U7946 (N_7946,N_7743,N_7693);
nor U7947 (N_7947,N_7615,N_7794);
nor U7948 (N_7948,N_7769,N_7694);
and U7949 (N_7949,N_7607,N_7689);
or U7950 (N_7950,N_7613,N_7612);
and U7951 (N_7951,N_7798,N_7623);
xor U7952 (N_7952,N_7606,N_7616);
and U7953 (N_7953,N_7769,N_7737);
and U7954 (N_7954,N_7788,N_7658);
xnor U7955 (N_7955,N_7614,N_7635);
nand U7956 (N_7956,N_7796,N_7667);
nor U7957 (N_7957,N_7783,N_7792);
or U7958 (N_7958,N_7609,N_7767);
and U7959 (N_7959,N_7675,N_7695);
and U7960 (N_7960,N_7702,N_7724);
or U7961 (N_7961,N_7775,N_7722);
xnor U7962 (N_7962,N_7626,N_7735);
nand U7963 (N_7963,N_7740,N_7668);
and U7964 (N_7964,N_7735,N_7707);
nor U7965 (N_7965,N_7721,N_7759);
xor U7966 (N_7966,N_7607,N_7708);
nand U7967 (N_7967,N_7671,N_7773);
nand U7968 (N_7968,N_7710,N_7630);
and U7969 (N_7969,N_7627,N_7764);
nand U7970 (N_7970,N_7619,N_7670);
xnor U7971 (N_7971,N_7646,N_7713);
nor U7972 (N_7972,N_7624,N_7705);
nor U7973 (N_7973,N_7679,N_7685);
and U7974 (N_7974,N_7663,N_7629);
nand U7975 (N_7975,N_7764,N_7651);
nor U7976 (N_7976,N_7611,N_7610);
xnor U7977 (N_7977,N_7756,N_7715);
xor U7978 (N_7978,N_7798,N_7783);
and U7979 (N_7979,N_7669,N_7693);
and U7980 (N_7980,N_7659,N_7779);
xor U7981 (N_7981,N_7661,N_7603);
nand U7982 (N_7982,N_7724,N_7625);
nand U7983 (N_7983,N_7622,N_7779);
and U7984 (N_7984,N_7751,N_7773);
xor U7985 (N_7985,N_7786,N_7747);
or U7986 (N_7986,N_7663,N_7606);
nand U7987 (N_7987,N_7669,N_7738);
or U7988 (N_7988,N_7666,N_7685);
nor U7989 (N_7989,N_7745,N_7736);
and U7990 (N_7990,N_7626,N_7775);
and U7991 (N_7991,N_7628,N_7682);
and U7992 (N_7992,N_7724,N_7794);
and U7993 (N_7993,N_7720,N_7607);
nor U7994 (N_7994,N_7666,N_7699);
nand U7995 (N_7995,N_7678,N_7702);
nor U7996 (N_7996,N_7704,N_7692);
xor U7997 (N_7997,N_7694,N_7793);
nand U7998 (N_7998,N_7690,N_7706);
nand U7999 (N_7999,N_7714,N_7678);
and U8000 (N_8000,N_7801,N_7852);
or U8001 (N_8001,N_7856,N_7827);
nand U8002 (N_8002,N_7883,N_7966);
or U8003 (N_8003,N_7938,N_7984);
xnor U8004 (N_8004,N_7952,N_7957);
and U8005 (N_8005,N_7832,N_7875);
nor U8006 (N_8006,N_7840,N_7997);
or U8007 (N_8007,N_7820,N_7853);
or U8008 (N_8008,N_7915,N_7859);
nor U8009 (N_8009,N_7896,N_7826);
or U8010 (N_8010,N_7964,N_7973);
and U8011 (N_8011,N_7877,N_7812);
xor U8012 (N_8012,N_7946,N_7879);
xnor U8013 (N_8013,N_7903,N_7970);
nand U8014 (N_8014,N_7891,N_7987);
nand U8015 (N_8015,N_7981,N_7871);
xor U8016 (N_8016,N_7948,N_7963);
nand U8017 (N_8017,N_7874,N_7988);
xnor U8018 (N_8018,N_7803,N_7928);
or U8019 (N_8019,N_7895,N_7847);
and U8020 (N_8020,N_7909,N_7993);
nand U8021 (N_8021,N_7890,N_7887);
nand U8022 (N_8022,N_7880,N_7841);
nand U8023 (N_8023,N_7986,N_7810);
nor U8024 (N_8024,N_7975,N_7829);
nor U8025 (N_8025,N_7956,N_7935);
nand U8026 (N_8026,N_7980,N_7907);
or U8027 (N_8027,N_7889,N_7888);
nand U8028 (N_8028,N_7804,N_7991);
nor U8029 (N_8029,N_7979,N_7947);
nand U8030 (N_8030,N_7802,N_7843);
nand U8031 (N_8031,N_7822,N_7912);
xor U8032 (N_8032,N_7916,N_7908);
and U8033 (N_8033,N_7905,N_7958);
or U8034 (N_8034,N_7818,N_7815);
and U8035 (N_8035,N_7985,N_7924);
nand U8036 (N_8036,N_7950,N_7886);
xnor U8037 (N_8037,N_7869,N_7811);
or U8038 (N_8038,N_7837,N_7994);
nand U8039 (N_8039,N_7816,N_7844);
xnor U8040 (N_8040,N_7982,N_7959);
and U8041 (N_8041,N_7855,N_7940);
nor U8042 (N_8042,N_7944,N_7817);
nand U8043 (N_8043,N_7989,N_7901);
xor U8044 (N_8044,N_7834,N_7998);
xor U8045 (N_8045,N_7922,N_7990);
xnor U8046 (N_8046,N_7842,N_7846);
or U8047 (N_8047,N_7858,N_7845);
nand U8048 (N_8048,N_7942,N_7862);
xnor U8049 (N_8049,N_7867,N_7870);
nand U8050 (N_8050,N_7921,N_7839);
or U8051 (N_8051,N_7939,N_7974);
nor U8052 (N_8052,N_7899,N_7932);
xor U8053 (N_8053,N_7807,N_7865);
nand U8054 (N_8054,N_7849,N_7969);
xor U8055 (N_8055,N_7873,N_7960);
xnor U8056 (N_8056,N_7920,N_7930);
nand U8057 (N_8057,N_7983,N_7805);
and U8058 (N_8058,N_7996,N_7949);
and U8059 (N_8059,N_7897,N_7961);
xnor U8060 (N_8060,N_7941,N_7876);
or U8061 (N_8061,N_7819,N_7925);
and U8062 (N_8062,N_7923,N_7830);
and U8063 (N_8063,N_7913,N_7892);
xnor U8064 (N_8064,N_7850,N_7809);
nand U8065 (N_8065,N_7848,N_7934);
or U8066 (N_8066,N_7933,N_7972);
nand U8067 (N_8067,N_7945,N_7831);
and U8068 (N_8068,N_7868,N_7999);
nand U8069 (N_8069,N_7813,N_7833);
nand U8070 (N_8070,N_7835,N_7926);
or U8071 (N_8071,N_7954,N_7976);
nor U8072 (N_8072,N_7860,N_7825);
nor U8073 (N_8073,N_7894,N_7882);
xor U8074 (N_8074,N_7861,N_7823);
nand U8075 (N_8075,N_7902,N_7854);
or U8076 (N_8076,N_7851,N_7808);
or U8077 (N_8077,N_7943,N_7955);
or U8078 (N_8078,N_7857,N_7864);
xor U8079 (N_8079,N_7814,N_7929);
nor U8080 (N_8080,N_7995,N_7904);
nand U8081 (N_8081,N_7893,N_7918);
nand U8082 (N_8082,N_7936,N_7977);
xor U8083 (N_8083,N_7971,N_7967);
or U8084 (N_8084,N_7919,N_7917);
and U8085 (N_8085,N_7906,N_7821);
and U8086 (N_8086,N_7878,N_7872);
nor U8087 (N_8087,N_7968,N_7927);
and U8088 (N_8088,N_7910,N_7800);
nand U8089 (N_8089,N_7866,N_7937);
and U8090 (N_8090,N_7965,N_7885);
nor U8091 (N_8091,N_7931,N_7824);
xor U8092 (N_8092,N_7838,N_7806);
and U8093 (N_8093,N_7951,N_7898);
or U8094 (N_8094,N_7953,N_7863);
and U8095 (N_8095,N_7881,N_7884);
and U8096 (N_8096,N_7914,N_7911);
or U8097 (N_8097,N_7900,N_7992);
or U8098 (N_8098,N_7978,N_7836);
and U8099 (N_8099,N_7962,N_7828);
nand U8100 (N_8100,N_7998,N_7994);
xnor U8101 (N_8101,N_7891,N_7824);
and U8102 (N_8102,N_7838,N_7904);
xnor U8103 (N_8103,N_7814,N_7852);
nor U8104 (N_8104,N_7849,N_7808);
and U8105 (N_8105,N_7958,N_7969);
and U8106 (N_8106,N_7920,N_7944);
or U8107 (N_8107,N_7812,N_7935);
and U8108 (N_8108,N_7954,N_7809);
and U8109 (N_8109,N_7873,N_7947);
nor U8110 (N_8110,N_7800,N_7860);
nor U8111 (N_8111,N_7944,N_7956);
and U8112 (N_8112,N_7932,N_7931);
or U8113 (N_8113,N_7938,N_7851);
nor U8114 (N_8114,N_7825,N_7819);
nand U8115 (N_8115,N_7885,N_7977);
xor U8116 (N_8116,N_7962,N_7989);
nor U8117 (N_8117,N_7866,N_7890);
or U8118 (N_8118,N_7869,N_7956);
nand U8119 (N_8119,N_7897,N_7842);
xnor U8120 (N_8120,N_7962,N_7993);
nor U8121 (N_8121,N_7962,N_7966);
and U8122 (N_8122,N_7849,N_7999);
xnor U8123 (N_8123,N_7867,N_7840);
nand U8124 (N_8124,N_7818,N_7991);
xor U8125 (N_8125,N_7829,N_7889);
nor U8126 (N_8126,N_7981,N_7824);
or U8127 (N_8127,N_7870,N_7830);
or U8128 (N_8128,N_7999,N_7840);
or U8129 (N_8129,N_7991,N_7882);
xor U8130 (N_8130,N_7888,N_7860);
xnor U8131 (N_8131,N_7837,N_7981);
nand U8132 (N_8132,N_7916,N_7954);
nor U8133 (N_8133,N_7969,N_7887);
nor U8134 (N_8134,N_7805,N_7971);
nor U8135 (N_8135,N_7937,N_7811);
nor U8136 (N_8136,N_7850,N_7865);
and U8137 (N_8137,N_7960,N_7965);
and U8138 (N_8138,N_7972,N_7976);
or U8139 (N_8139,N_7801,N_7931);
or U8140 (N_8140,N_7970,N_7982);
or U8141 (N_8141,N_7883,N_7809);
or U8142 (N_8142,N_7866,N_7942);
and U8143 (N_8143,N_7909,N_7805);
nand U8144 (N_8144,N_7822,N_7837);
and U8145 (N_8145,N_7930,N_7875);
or U8146 (N_8146,N_7828,N_7802);
nand U8147 (N_8147,N_7868,N_7888);
nor U8148 (N_8148,N_7933,N_7999);
and U8149 (N_8149,N_7863,N_7914);
and U8150 (N_8150,N_7846,N_7911);
nor U8151 (N_8151,N_7917,N_7871);
xor U8152 (N_8152,N_7958,N_7908);
or U8153 (N_8153,N_7849,N_7942);
xnor U8154 (N_8154,N_7974,N_7892);
or U8155 (N_8155,N_7938,N_7848);
xnor U8156 (N_8156,N_7994,N_7805);
nand U8157 (N_8157,N_7895,N_7973);
nand U8158 (N_8158,N_7878,N_7866);
or U8159 (N_8159,N_7857,N_7908);
or U8160 (N_8160,N_7974,N_7879);
xor U8161 (N_8161,N_7865,N_7857);
or U8162 (N_8162,N_7976,N_7909);
nand U8163 (N_8163,N_7832,N_7952);
xor U8164 (N_8164,N_7993,N_7928);
xnor U8165 (N_8165,N_7846,N_7802);
nand U8166 (N_8166,N_7948,N_7983);
nand U8167 (N_8167,N_7804,N_7892);
nor U8168 (N_8168,N_7880,N_7901);
nand U8169 (N_8169,N_7859,N_7953);
nor U8170 (N_8170,N_7982,N_7803);
nor U8171 (N_8171,N_7821,N_7973);
xnor U8172 (N_8172,N_7813,N_7946);
nand U8173 (N_8173,N_7998,N_7949);
or U8174 (N_8174,N_7988,N_7887);
nand U8175 (N_8175,N_7823,N_7927);
xnor U8176 (N_8176,N_7872,N_7913);
xor U8177 (N_8177,N_7945,N_7824);
nand U8178 (N_8178,N_7842,N_7982);
nand U8179 (N_8179,N_7936,N_7808);
xnor U8180 (N_8180,N_7846,N_7943);
nand U8181 (N_8181,N_7819,N_7928);
xnor U8182 (N_8182,N_7977,N_7888);
nor U8183 (N_8183,N_7860,N_7820);
nand U8184 (N_8184,N_7913,N_7880);
and U8185 (N_8185,N_7926,N_7975);
nor U8186 (N_8186,N_7918,N_7913);
and U8187 (N_8187,N_7952,N_7817);
xnor U8188 (N_8188,N_7908,N_7992);
and U8189 (N_8189,N_7866,N_7857);
nand U8190 (N_8190,N_7864,N_7979);
nor U8191 (N_8191,N_7969,N_7840);
nand U8192 (N_8192,N_7932,N_7914);
nor U8193 (N_8193,N_7941,N_7892);
or U8194 (N_8194,N_7914,N_7881);
nand U8195 (N_8195,N_7826,N_7865);
xnor U8196 (N_8196,N_7920,N_7976);
and U8197 (N_8197,N_7976,N_7872);
xnor U8198 (N_8198,N_7871,N_7838);
nor U8199 (N_8199,N_7945,N_7814);
and U8200 (N_8200,N_8146,N_8099);
nand U8201 (N_8201,N_8023,N_8083);
nand U8202 (N_8202,N_8059,N_8121);
nor U8203 (N_8203,N_8001,N_8073);
and U8204 (N_8204,N_8141,N_8060);
xor U8205 (N_8205,N_8105,N_8123);
or U8206 (N_8206,N_8101,N_8176);
or U8207 (N_8207,N_8010,N_8040);
or U8208 (N_8208,N_8072,N_8156);
or U8209 (N_8209,N_8033,N_8122);
xor U8210 (N_8210,N_8140,N_8197);
and U8211 (N_8211,N_8104,N_8064);
nor U8212 (N_8212,N_8149,N_8017);
or U8213 (N_8213,N_8186,N_8002);
or U8214 (N_8214,N_8160,N_8182);
and U8215 (N_8215,N_8139,N_8069);
nor U8216 (N_8216,N_8047,N_8046);
and U8217 (N_8217,N_8056,N_8092);
nand U8218 (N_8218,N_8079,N_8096);
or U8219 (N_8219,N_8021,N_8129);
nand U8220 (N_8220,N_8116,N_8095);
nand U8221 (N_8221,N_8189,N_8000);
or U8222 (N_8222,N_8067,N_8034);
and U8223 (N_8223,N_8026,N_8113);
nor U8224 (N_8224,N_8037,N_8147);
xor U8225 (N_8225,N_8175,N_8075);
xnor U8226 (N_8226,N_8117,N_8103);
xor U8227 (N_8227,N_8100,N_8187);
nor U8228 (N_8228,N_8198,N_8162);
nand U8229 (N_8229,N_8039,N_8024);
nand U8230 (N_8230,N_8041,N_8020);
xnor U8231 (N_8231,N_8038,N_8136);
nand U8232 (N_8232,N_8170,N_8199);
or U8233 (N_8233,N_8012,N_8159);
or U8234 (N_8234,N_8089,N_8131);
and U8235 (N_8235,N_8157,N_8152);
xnor U8236 (N_8236,N_8062,N_8077);
nand U8237 (N_8237,N_8155,N_8044);
and U8238 (N_8238,N_8030,N_8018);
and U8239 (N_8239,N_8063,N_8013);
xor U8240 (N_8240,N_8179,N_8008);
or U8241 (N_8241,N_8087,N_8066);
xor U8242 (N_8242,N_8164,N_8082);
nor U8243 (N_8243,N_8184,N_8188);
nor U8244 (N_8244,N_8055,N_8169);
nand U8245 (N_8245,N_8015,N_8108);
nor U8246 (N_8246,N_8126,N_8115);
xor U8247 (N_8247,N_8093,N_8194);
xor U8248 (N_8248,N_8135,N_8045);
nand U8249 (N_8249,N_8120,N_8050);
and U8250 (N_8250,N_8193,N_8009);
nand U8251 (N_8251,N_8004,N_8029);
nand U8252 (N_8252,N_8031,N_8173);
nand U8253 (N_8253,N_8074,N_8130);
nor U8254 (N_8254,N_8181,N_8058);
xor U8255 (N_8255,N_8167,N_8097);
and U8256 (N_8256,N_8014,N_8042);
nand U8257 (N_8257,N_8165,N_8106);
nor U8258 (N_8258,N_8027,N_8016);
nor U8259 (N_8259,N_8051,N_8171);
xor U8260 (N_8260,N_8161,N_8005);
nand U8261 (N_8261,N_8142,N_8007);
and U8262 (N_8262,N_8022,N_8057);
nand U8263 (N_8263,N_8118,N_8134);
nor U8264 (N_8264,N_8081,N_8191);
xnor U8265 (N_8265,N_8195,N_8091);
nand U8266 (N_8266,N_8019,N_8185);
or U8267 (N_8267,N_8085,N_8144);
and U8268 (N_8268,N_8084,N_8110);
xnor U8269 (N_8269,N_8048,N_8168);
xnor U8270 (N_8270,N_8124,N_8070);
and U8271 (N_8271,N_8192,N_8065);
nor U8272 (N_8272,N_8076,N_8052);
nor U8273 (N_8273,N_8011,N_8025);
and U8274 (N_8274,N_8196,N_8154);
nand U8275 (N_8275,N_8107,N_8138);
nor U8276 (N_8276,N_8190,N_8049);
nand U8277 (N_8277,N_8178,N_8132);
or U8278 (N_8278,N_8163,N_8028);
nor U8279 (N_8279,N_8153,N_8158);
nand U8280 (N_8280,N_8111,N_8151);
or U8281 (N_8281,N_8090,N_8166);
or U8282 (N_8282,N_8102,N_8109);
nand U8283 (N_8283,N_8180,N_8174);
nor U8284 (N_8284,N_8148,N_8061);
nor U8285 (N_8285,N_8125,N_8003);
and U8286 (N_8286,N_8172,N_8006);
nor U8287 (N_8287,N_8183,N_8098);
or U8288 (N_8288,N_8054,N_8094);
xor U8289 (N_8289,N_8128,N_8119);
xor U8290 (N_8290,N_8053,N_8133);
xor U8291 (N_8291,N_8112,N_8150);
or U8292 (N_8292,N_8036,N_8032);
and U8293 (N_8293,N_8114,N_8086);
xnor U8294 (N_8294,N_8177,N_8088);
or U8295 (N_8295,N_8078,N_8145);
xnor U8296 (N_8296,N_8071,N_8068);
nand U8297 (N_8297,N_8137,N_8127);
or U8298 (N_8298,N_8043,N_8143);
and U8299 (N_8299,N_8080,N_8035);
nand U8300 (N_8300,N_8010,N_8035);
xnor U8301 (N_8301,N_8029,N_8112);
nand U8302 (N_8302,N_8180,N_8158);
or U8303 (N_8303,N_8110,N_8129);
nand U8304 (N_8304,N_8099,N_8106);
and U8305 (N_8305,N_8176,N_8005);
nor U8306 (N_8306,N_8169,N_8071);
xor U8307 (N_8307,N_8190,N_8165);
nor U8308 (N_8308,N_8188,N_8138);
nor U8309 (N_8309,N_8191,N_8106);
nor U8310 (N_8310,N_8111,N_8084);
nor U8311 (N_8311,N_8155,N_8007);
or U8312 (N_8312,N_8069,N_8160);
and U8313 (N_8313,N_8026,N_8126);
nand U8314 (N_8314,N_8140,N_8150);
nand U8315 (N_8315,N_8109,N_8030);
nand U8316 (N_8316,N_8004,N_8156);
nor U8317 (N_8317,N_8126,N_8165);
and U8318 (N_8318,N_8183,N_8144);
nand U8319 (N_8319,N_8104,N_8084);
and U8320 (N_8320,N_8161,N_8085);
and U8321 (N_8321,N_8122,N_8183);
nor U8322 (N_8322,N_8010,N_8007);
nand U8323 (N_8323,N_8048,N_8101);
nand U8324 (N_8324,N_8050,N_8000);
or U8325 (N_8325,N_8087,N_8068);
and U8326 (N_8326,N_8064,N_8173);
nor U8327 (N_8327,N_8082,N_8084);
nor U8328 (N_8328,N_8073,N_8033);
xor U8329 (N_8329,N_8161,N_8067);
or U8330 (N_8330,N_8110,N_8031);
and U8331 (N_8331,N_8143,N_8112);
or U8332 (N_8332,N_8196,N_8028);
xor U8333 (N_8333,N_8032,N_8150);
xor U8334 (N_8334,N_8100,N_8181);
and U8335 (N_8335,N_8177,N_8024);
xor U8336 (N_8336,N_8150,N_8124);
or U8337 (N_8337,N_8013,N_8110);
nand U8338 (N_8338,N_8021,N_8052);
or U8339 (N_8339,N_8123,N_8112);
or U8340 (N_8340,N_8194,N_8197);
and U8341 (N_8341,N_8071,N_8073);
or U8342 (N_8342,N_8154,N_8097);
or U8343 (N_8343,N_8081,N_8158);
or U8344 (N_8344,N_8084,N_8060);
xor U8345 (N_8345,N_8077,N_8046);
xor U8346 (N_8346,N_8039,N_8128);
and U8347 (N_8347,N_8110,N_8142);
and U8348 (N_8348,N_8139,N_8153);
nand U8349 (N_8349,N_8126,N_8091);
and U8350 (N_8350,N_8159,N_8080);
xnor U8351 (N_8351,N_8064,N_8176);
nor U8352 (N_8352,N_8073,N_8128);
nand U8353 (N_8353,N_8036,N_8131);
xnor U8354 (N_8354,N_8153,N_8065);
and U8355 (N_8355,N_8160,N_8118);
nor U8356 (N_8356,N_8014,N_8187);
and U8357 (N_8357,N_8019,N_8087);
and U8358 (N_8358,N_8077,N_8070);
nand U8359 (N_8359,N_8130,N_8085);
nor U8360 (N_8360,N_8168,N_8137);
xnor U8361 (N_8361,N_8079,N_8107);
nor U8362 (N_8362,N_8070,N_8130);
nand U8363 (N_8363,N_8191,N_8099);
nor U8364 (N_8364,N_8038,N_8117);
or U8365 (N_8365,N_8105,N_8161);
nand U8366 (N_8366,N_8130,N_8051);
nor U8367 (N_8367,N_8034,N_8152);
xnor U8368 (N_8368,N_8180,N_8098);
and U8369 (N_8369,N_8011,N_8142);
and U8370 (N_8370,N_8146,N_8121);
and U8371 (N_8371,N_8115,N_8068);
or U8372 (N_8372,N_8049,N_8034);
nand U8373 (N_8373,N_8170,N_8185);
and U8374 (N_8374,N_8070,N_8047);
nand U8375 (N_8375,N_8154,N_8099);
xor U8376 (N_8376,N_8006,N_8053);
xnor U8377 (N_8377,N_8061,N_8165);
and U8378 (N_8378,N_8180,N_8083);
nor U8379 (N_8379,N_8010,N_8185);
nor U8380 (N_8380,N_8136,N_8174);
nor U8381 (N_8381,N_8159,N_8092);
nand U8382 (N_8382,N_8132,N_8067);
or U8383 (N_8383,N_8174,N_8070);
or U8384 (N_8384,N_8040,N_8098);
nor U8385 (N_8385,N_8107,N_8136);
nor U8386 (N_8386,N_8016,N_8031);
nand U8387 (N_8387,N_8095,N_8064);
and U8388 (N_8388,N_8137,N_8054);
xor U8389 (N_8389,N_8049,N_8150);
xnor U8390 (N_8390,N_8140,N_8023);
xor U8391 (N_8391,N_8007,N_8098);
and U8392 (N_8392,N_8039,N_8086);
and U8393 (N_8393,N_8162,N_8061);
nand U8394 (N_8394,N_8036,N_8098);
and U8395 (N_8395,N_8131,N_8190);
and U8396 (N_8396,N_8167,N_8067);
or U8397 (N_8397,N_8185,N_8138);
or U8398 (N_8398,N_8055,N_8144);
or U8399 (N_8399,N_8191,N_8171);
or U8400 (N_8400,N_8322,N_8353);
nor U8401 (N_8401,N_8313,N_8342);
xnor U8402 (N_8402,N_8293,N_8294);
and U8403 (N_8403,N_8200,N_8378);
nor U8404 (N_8404,N_8235,N_8239);
nor U8405 (N_8405,N_8201,N_8391);
nor U8406 (N_8406,N_8269,N_8381);
or U8407 (N_8407,N_8278,N_8373);
nor U8408 (N_8408,N_8386,N_8286);
and U8409 (N_8409,N_8205,N_8334);
and U8410 (N_8410,N_8291,N_8399);
or U8411 (N_8411,N_8394,N_8232);
and U8412 (N_8412,N_8243,N_8330);
xnor U8413 (N_8413,N_8241,N_8212);
and U8414 (N_8414,N_8204,N_8288);
nand U8415 (N_8415,N_8385,N_8344);
and U8416 (N_8416,N_8206,N_8244);
or U8417 (N_8417,N_8375,N_8215);
xor U8418 (N_8418,N_8257,N_8304);
or U8419 (N_8419,N_8301,N_8335);
nor U8420 (N_8420,N_8372,N_8229);
nor U8421 (N_8421,N_8316,N_8392);
nand U8422 (N_8422,N_8389,N_8209);
xor U8423 (N_8423,N_8282,N_8332);
and U8424 (N_8424,N_8219,N_8213);
nor U8425 (N_8425,N_8302,N_8327);
xnor U8426 (N_8426,N_8208,N_8211);
or U8427 (N_8427,N_8272,N_8258);
xnor U8428 (N_8428,N_8326,N_8336);
nor U8429 (N_8429,N_8298,N_8317);
nand U8430 (N_8430,N_8305,N_8383);
nand U8431 (N_8431,N_8210,N_8311);
or U8432 (N_8432,N_8279,N_8397);
or U8433 (N_8433,N_8221,N_8228);
nand U8434 (N_8434,N_8380,N_8226);
xnor U8435 (N_8435,N_8325,N_8339);
xnor U8436 (N_8436,N_8249,N_8275);
nand U8437 (N_8437,N_8233,N_8214);
nand U8438 (N_8438,N_8358,N_8237);
xor U8439 (N_8439,N_8216,N_8289);
or U8440 (N_8440,N_8370,N_8267);
and U8441 (N_8441,N_8250,N_8341);
and U8442 (N_8442,N_8276,N_8247);
xnor U8443 (N_8443,N_8309,N_8310);
and U8444 (N_8444,N_8382,N_8281);
xnor U8445 (N_8445,N_8352,N_8356);
nand U8446 (N_8446,N_8395,N_8285);
or U8447 (N_8447,N_8300,N_8396);
and U8448 (N_8448,N_8303,N_8355);
or U8449 (N_8449,N_8263,N_8217);
nand U8450 (N_8450,N_8331,N_8369);
nor U8451 (N_8451,N_8277,N_8315);
nor U8452 (N_8452,N_8280,N_8230);
xnor U8453 (N_8453,N_8357,N_8371);
nor U8454 (N_8454,N_8318,N_8266);
or U8455 (N_8455,N_8374,N_8359);
and U8456 (N_8456,N_8296,N_8393);
nor U8457 (N_8457,N_8340,N_8225);
or U8458 (N_8458,N_8207,N_8361);
nand U8459 (N_8459,N_8248,N_8268);
or U8460 (N_8460,N_8240,N_8324);
nor U8461 (N_8461,N_8387,N_8284);
or U8462 (N_8462,N_8314,N_8377);
xor U8463 (N_8463,N_8349,N_8218);
nor U8464 (N_8464,N_8319,N_8320);
xor U8465 (N_8465,N_8222,N_8271);
nor U8466 (N_8466,N_8307,N_8236);
xnor U8467 (N_8467,N_8295,N_8368);
xnor U8468 (N_8468,N_8363,N_8347);
and U8469 (N_8469,N_8252,N_8246);
or U8470 (N_8470,N_8220,N_8343);
nor U8471 (N_8471,N_8260,N_8287);
xnor U8472 (N_8472,N_8367,N_8338);
nand U8473 (N_8473,N_8264,N_8306);
nor U8474 (N_8474,N_8366,N_8231);
nand U8475 (N_8475,N_8362,N_8388);
nor U8476 (N_8476,N_8242,N_8292);
nand U8477 (N_8477,N_8398,N_8234);
nand U8478 (N_8478,N_8360,N_8238);
xnor U8479 (N_8479,N_8376,N_8346);
and U8480 (N_8480,N_8348,N_8329);
or U8481 (N_8481,N_8227,N_8251);
nand U8482 (N_8482,N_8333,N_8202);
xnor U8483 (N_8483,N_8351,N_8223);
nor U8484 (N_8484,N_8254,N_8274);
nand U8485 (N_8485,N_8384,N_8245);
and U8486 (N_8486,N_8364,N_8203);
or U8487 (N_8487,N_8350,N_8297);
xor U8488 (N_8488,N_8273,N_8255);
and U8489 (N_8489,N_8345,N_8312);
and U8490 (N_8490,N_8259,N_8256);
nor U8491 (N_8491,N_8308,N_8262);
and U8492 (N_8492,N_8253,N_8283);
xnor U8493 (N_8493,N_8321,N_8390);
nor U8494 (N_8494,N_8261,N_8337);
and U8495 (N_8495,N_8265,N_8224);
and U8496 (N_8496,N_8270,N_8354);
nor U8497 (N_8497,N_8323,N_8299);
or U8498 (N_8498,N_8365,N_8328);
nor U8499 (N_8499,N_8379,N_8290);
or U8500 (N_8500,N_8356,N_8270);
nor U8501 (N_8501,N_8322,N_8212);
nor U8502 (N_8502,N_8264,N_8274);
xnor U8503 (N_8503,N_8291,N_8206);
and U8504 (N_8504,N_8372,N_8260);
nor U8505 (N_8505,N_8391,N_8226);
nand U8506 (N_8506,N_8275,N_8361);
nand U8507 (N_8507,N_8304,N_8284);
nand U8508 (N_8508,N_8224,N_8233);
and U8509 (N_8509,N_8315,N_8309);
nor U8510 (N_8510,N_8386,N_8332);
and U8511 (N_8511,N_8388,N_8231);
nand U8512 (N_8512,N_8371,N_8300);
nand U8513 (N_8513,N_8241,N_8233);
nand U8514 (N_8514,N_8265,N_8253);
and U8515 (N_8515,N_8216,N_8239);
and U8516 (N_8516,N_8363,N_8279);
nor U8517 (N_8517,N_8279,N_8261);
or U8518 (N_8518,N_8266,N_8395);
or U8519 (N_8519,N_8343,N_8314);
xor U8520 (N_8520,N_8326,N_8244);
nand U8521 (N_8521,N_8392,N_8264);
nor U8522 (N_8522,N_8337,N_8329);
and U8523 (N_8523,N_8250,N_8315);
or U8524 (N_8524,N_8276,N_8222);
or U8525 (N_8525,N_8229,N_8269);
xor U8526 (N_8526,N_8303,N_8315);
nor U8527 (N_8527,N_8346,N_8271);
nor U8528 (N_8528,N_8375,N_8333);
or U8529 (N_8529,N_8377,N_8380);
or U8530 (N_8530,N_8382,N_8311);
and U8531 (N_8531,N_8386,N_8255);
nand U8532 (N_8532,N_8305,N_8220);
and U8533 (N_8533,N_8375,N_8237);
or U8534 (N_8534,N_8320,N_8263);
and U8535 (N_8535,N_8372,N_8303);
nor U8536 (N_8536,N_8208,N_8331);
xnor U8537 (N_8537,N_8243,N_8377);
or U8538 (N_8538,N_8232,N_8300);
xor U8539 (N_8539,N_8224,N_8241);
or U8540 (N_8540,N_8203,N_8200);
nor U8541 (N_8541,N_8233,N_8277);
nor U8542 (N_8542,N_8307,N_8381);
xnor U8543 (N_8543,N_8385,N_8388);
or U8544 (N_8544,N_8343,N_8392);
and U8545 (N_8545,N_8351,N_8306);
nor U8546 (N_8546,N_8296,N_8261);
and U8547 (N_8547,N_8331,N_8264);
xnor U8548 (N_8548,N_8268,N_8355);
nand U8549 (N_8549,N_8327,N_8358);
and U8550 (N_8550,N_8388,N_8264);
nand U8551 (N_8551,N_8277,N_8226);
or U8552 (N_8552,N_8308,N_8340);
nand U8553 (N_8553,N_8396,N_8257);
or U8554 (N_8554,N_8271,N_8372);
and U8555 (N_8555,N_8219,N_8370);
or U8556 (N_8556,N_8305,N_8303);
nor U8557 (N_8557,N_8221,N_8284);
xnor U8558 (N_8558,N_8290,N_8215);
nand U8559 (N_8559,N_8205,N_8372);
and U8560 (N_8560,N_8347,N_8329);
xor U8561 (N_8561,N_8306,N_8347);
nor U8562 (N_8562,N_8213,N_8268);
nand U8563 (N_8563,N_8372,N_8343);
nand U8564 (N_8564,N_8395,N_8280);
nand U8565 (N_8565,N_8212,N_8262);
xor U8566 (N_8566,N_8200,N_8318);
xnor U8567 (N_8567,N_8261,N_8225);
nand U8568 (N_8568,N_8397,N_8388);
xor U8569 (N_8569,N_8287,N_8315);
nand U8570 (N_8570,N_8225,N_8347);
or U8571 (N_8571,N_8382,N_8394);
nor U8572 (N_8572,N_8374,N_8200);
and U8573 (N_8573,N_8271,N_8219);
and U8574 (N_8574,N_8209,N_8324);
xor U8575 (N_8575,N_8319,N_8204);
nand U8576 (N_8576,N_8253,N_8233);
and U8577 (N_8577,N_8293,N_8304);
nand U8578 (N_8578,N_8353,N_8371);
and U8579 (N_8579,N_8228,N_8255);
nand U8580 (N_8580,N_8317,N_8213);
nor U8581 (N_8581,N_8243,N_8287);
or U8582 (N_8582,N_8264,N_8252);
nor U8583 (N_8583,N_8354,N_8295);
xnor U8584 (N_8584,N_8200,N_8376);
or U8585 (N_8585,N_8395,N_8236);
nand U8586 (N_8586,N_8206,N_8377);
or U8587 (N_8587,N_8354,N_8378);
nand U8588 (N_8588,N_8343,N_8270);
nand U8589 (N_8589,N_8200,N_8309);
xor U8590 (N_8590,N_8256,N_8366);
xor U8591 (N_8591,N_8333,N_8261);
or U8592 (N_8592,N_8390,N_8250);
nor U8593 (N_8593,N_8206,N_8381);
nor U8594 (N_8594,N_8355,N_8292);
xnor U8595 (N_8595,N_8340,N_8256);
and U8596 (N_8596,N_8342,N_8247);
or U8597 (N_8597,N_8234,N_8341);
and U8598 (N_8598,N_8339,N_8251);
and U8599 (N_8599,N_8272,N_8331);
xor U8600 (N_8600,N_8530,N_8455);
or U8601 (N_8601,N_8417,N_8432);
nand U8602 (N_8602,N_8471,N_8409);
nor U8603 (N_8603,N_8588,N_8434);
xnor U8604 (N_8604,N_8597,N_8454);
xnor U8605 (N_8605,N_8436,N_8502);
or U8606 (N_8606,N_8523,N_8441);
and U8607 (N_8607,N_8499,N_8426);
nor U8608 (N_8608,N_8488,N_8570);
nand U8609 (N_8609,N_8572,N_8527);
xnor U8610 (N_8610,N_8549,N_8560);
xor U8611 (N_8611,N_8403,N_8518);
or U8612 (N_8612,N_8489,N_8457);
nor U8613 (N_8613,N_8438,N_8575);
or U8614 (N_8614,N_8483,N_8507);
or U8615 (N_8615,N_8584,N_8578);
nand U8616 (N_8616,N_8559,N_8539);
nor U8617 (N_8617,N_8558,N_8585);
nor U8618 (N_8618,N_8520,N_8464);
and U8619 (N_8619,N_8477,N_8592);
or U8620 (N_8620,N_8583,N_8548);
nand U8621 (N_8621,N_8472,N_8406);
nand U8622 (N_8622,N_8431,N_8571);
and U8623 (N_8623,N_8561,N_8490);
nand U8624 (N_8624,N_8435,N_8555);
or U8625 (N_8625,N_8475,N_8513);
or U8626 (N_8626,N_8460,N_8508);
xor U8627 (N_8627,N_8517,N_8594);
or U8628 (N_8628,N_8566,N_8540);
or U8629 (N_8629,N_8416,N_8481);
xnor U8630 (N_8630,N_8595,N_8497);
nand U8631 (N_8631,N_8532,N_8545);
or U8632 (N_8632,N_8451,N_8596);
or U8633 (N_8633,N_8599,N_8402);
nand U8634 (N_8634,N_8466,N_8452);
or U8635 (N_8635,N_8492,N_8414);
or U8636 (N_8636,N_8524,N_8569);
xnor U8637 (N_8637,N_8498,N_8586);
and U8638 (N_8638,N_8427,N_8410);
and U8639 (N_8639,N_8456,N_8542);
nor U8640 (N_8640,N_8593,N_8430);
nand U8641 (N_8641,N_8554,N_8538);
xor U8642 (N_8642,N_8400,N_8485);
xor U8643 (N_8643,N_8501,N_8467);
and U8644 (N_8644,N_8437,N_8468);
or U8645 (N_8645,N_8550,N_8557);
or U8646 (N_8646,N_8473,N_8506);
xnor U8647 (N_8647,N_8465,N_8478);
or U8648 (N_8648,N_8419,N_8421);
or U8649 (N_8649,N_8500,N_8579);
or U8650 (N_8650,N_8553,N_8444);
nand U8651 (N_8651,N_8496,N_8439);
nand U8652 (N_8652,N_8440,N_8546);
nor U8653 (N_8653,N_8474,N_8521);
xnor U8654 (N_8654,N_8535,N_8459);
or U8655 (N_8655,N_8494,N_8528);
xnor U8656 (N_8656,N_8526,N_8408);
and U8657 (N_8657,N_8525,N_8505);
and U8658 (N_8658,N_8536,N_8581);
nor U8659 (N_8659,N_8568,N_8482);
and U8660 (N_8660,N_8458,N_8531);
nand U8661 (N_8661,N_8407,N_8463);
nor U8662 (N_8662,N_8551,N_8495);
and U8663 (N_8663,N_8470,N_8462);
or U8664 (N_8664,N_8418,N_8552);
xnor U8665 (N_8665,N_8533,N_8447);
nand U8666 (N_8666,N_8519,N_8428);
nand U8667 (N_8667,N_8476,N_8514);
and U8668 (N_8668,N_8547,N_8405);
xnor U8669 (N_8669,N_8541,N_8504);
and U8670 (N_8670,N_8404,N_8537);
xor U8671 (N_8671,N_8587,N_8484);
nor U8672 (N_8672,N_8577,N_8576);
or U8673 (N_8673,N_8590,N_8574);
xor U8674 (N_8674,N_8442,N_8516);
nor U8675 (N_8675,N_8573,N_8429);
xor U8676 (N_8676,N_8512,N_8461);
nand U8677 (N_8677,N_8509,N_8445);
xnor U8678 (N_8678,N_8591,N_8423);
nand U8679 (N_8679,N_8589,N_8479);
nor U8680 (N_8680,N_8480,N_8487);
xor U8681 (N_8681,N_8510,N_8401);
nor U8682 (N_8682,N_8453,N_8515);
xnor U8683 (N_8683,N_8582,N_8493);
and U8684 (N_8684,N_8446,N_8448);
or U8685 (N_8685,N_8424,N_8562);
nor U8686 (N_8686,N_8425,N_8522);
and U8687 (N_8687,N_8564,N_8443);
nor U8688 (N_8688,N_8580,N_8411);
or U8689 (N_8689,N_8529,N_8433);
nand U8690 (N_8690,N_8449,N_8469);
or U8691 (N_8691,N_8420,N_8563);
and U8692 (N_8692,N_8413,N_8511);
nand U8693 (N_8693,N_8556,N_8503);
nand U8694 (N_8694,N_8450,N_8565);
xor U8695 (N_8695,N_8544,N_8491);
nor U8696 (N_8696,N_8486,N_8415);
and U8697 (N_8697,N_8422,N_8567);
or U8698 (N_8698,N_8598,N_8534);
nand U8699 (N_8699,N_8412,N_8543);
or U8700 (N_8700,N_8552,N_8589);
nand U8701 (N_8701,N_8586,N_8431);
and U8702 (N_8702,N_8404,N_8494);
or U8703 (N_8703,N_8598,N_8473);
nand U8704 (N_8704,N_8497,N_8531);
xor U8705 (N_8705,N_8502,N_8520);
or U8706 (N_8706,N_8504,N_8563);
nand U8707 (N_8707,N_8406,N_8436);
and U8708 (N_8708,N_8444,N_8588);
xor U8709 (N_8709,N_8497,N_8579);
nand U8710 (N_8710,N_8444,N_8468);
nor U8711 (N_8711,N_8433,N_8509);
nor U8712 (N_8712,N_8526,N_8520);
and U8713 (N_8713,N_8428,N_8524);
and U8714 (N_8714,N_8550,N_8587);
xor U8715 (N_8715,N_8422,N_8593);
nand U8716 (N_8716,N_8409,N_8460);
and U8717 (N_8717,N_8443,N_8420);
xor U8718 (N_8718,N_8445,N_8532);
nor U8719 (N_8719,N_8428,N_8419);
or U8720 (N_8720,N_8476,N_8502);
and U8721 (N_8721,N_8560,N_8442);
or U8722 (N_8722,N_8559,N_8585);
and U8723 (N_8723,N_8424,N_8417);
and U8724 (N_8724,N_8401,N_8430);
xor U8725 (N_8725,N_8411,N_8494);
and U8726 (N_8726,N_8503,N_8432);
or U8727 (N_8727,N_8483,N_8481);
or U8728 (N_8728,N_8465,N_8476);
nand U8729 (N_8729,N_8541,N_8473);
nor U8730 (N_8730,N_8561,N_8550);
nor U8731 (N_8731,N_8506,N_8417);
or U8732 (N_8732,N_8580,N_8572);
nor U8733 (N_8733,N_8519,N_8503);
or U8734 (N_8734,N_8547,N_8505);
nor U8735 (N_8735,N_8530,N_8474);
nor U8736 (N_8736,N_8573,N_8422);
nor U8737 (N_8737,N_8510,N_8413);
xor U8738 (N_8738,N_8578,N_8519);
nand U8739 (N_8739,N_8426,N_8585);
and U8740 (N_8740,N_8459,N_8416);
nor U8741 (N_8741,N_8568,N_8571);
xnor U8742 (N_8742,N_8525,N_8555);
or U8743 (N_8743,N_8501,N_8469);
and U8744 (N_8744,N_8469,N_8442);
xnor U8745 (N_8745,N_8592,N_8432);
or U8746 (N_8746,N_8403,N_8504);
nand U8747 (N_8747,N_8581,N_8414);
or U8748 (N_8748,N_8590,N_8594);
xnor U8749 (N_8749,N_8534,N_8559);
or U8750 (N_8750,N_8401,N_8427);
or U8751 (N_8751,N_8573,N_8412);
xnor U8752 (N_8752,N_8533,N_8453);
nor U8753 (N_8753,N_8498,N_8518);
nor U8754 (N_8754,N_8576,N_8471);
and U8755 (N_8755,N_8450,N_8490);
and U8756 (N_8756,N_8504,N_8503);
nand U8757 (N_8757,N_8519,N_8481);
or U8758 (N_8758,N_8483,N_8474);
and U8759 (N_8759,N_8520,N_8555);
nor U8760 (N_8760,N_8400,N_8442);
nor U8761 (N_8761,N_8426,N_8497);
nor U8762 (N_8762,N_8460,N_8585);
xor U8763 (N_8763,N_8550,N_8492);
nand U8764 (N_8764,N_8493,N_8470);
and U8765 (N_8765,N_8445,N_8403);
and U8766 (N_8766,N_8546,N_8426);
nor U8767 (N_8767,N_8404,N_8531);
or U8768 (N_8768,N_8529,N_8432);
or U8769 (N_8769,N_8516,N_8473);
and U8770 (N_8770,N_8492,N_8535);
nor U8771 (N_8771,N_8435,N_8598);
xor U8772 (N_8772,N_8400,N_8467);
and U8773 (N_8773,N_8436,N_8525);
nor U8774 (N_8774,N_8580,N_8402);
and U8775 (N_8775,N_8483,N_8449);
xor U8776 (N_8776,N_8418,N_8583);
xor U8777 (N_8777,N_8524,N_8422);
and U8778 (N_8778,N_8541,N_8435);
and U8779 (N_8779,N_8462,N_8472);
and U8780 (N_8780,N_8407,N_8578);
and U8781 (N_8781,N_8436,N_8540);
nor U8782 (N_8782,N_8570,N_8504);
nor U8783 (N_8783,N_8582,N_8418);
or U8784 (N_8784,N_8417,N_8484);
nor U8785 (N_8785,N_8536,N_8524);
nand U8786 (N_8786,N_8544,N_8463);
or U8787 (N_8787,N_8508,N_8496);
and U8788 (N_8788,N_8401,N_8468);
nor U8789 (N_8789,N_8430,N_8461);
xor U8790 (N_8790,N_8466,N_8548);
and U8791 (N_8791,N_8440,N_8589);
xor U8792 (N_8792,N_8472,N_8570);
nand U8793 (N_8793,N_8415,N_8593);
nor U8794 (N_8794,N_8585,N_8528);
nand U8795 (N_8795,N_8400,N_8542);
nor U8796 (N_8796,N_8434,N_8444);
xor U8797 (N_8797,N_8596,N_8508);
xor U8798 (N_8798,N_8443,N_8504);
nand U8799 (N_8799,N_8446,N_8441);
and U8800 (N_8800,N_8716,N_8622);
or U8801 (N_8801,N_8761,N_8726);
or U8802 (N_8802,N_8668,N_8678);
nor U8803 (N_8803,N_8680,N_8626);
nor U8804 (N_8804,N_8607,N_8650);
or U8805 (N_8805,N_8682,N_8690);
nand U8806 (N_8806,N_8773,N_8713);
and U8807 (N_8807,N_8608,N_8776);
nand U8808 (N_8808,N_8791,N_8747);
nand U8809 (N_8809,N_8621,N_8685);
nand U8810 (N_8810,N_8649,N_8697);
and U8811 (N_8811,N_8752,N_8722);
xnor U8812 (N_8812,N_8727,N_8788);
nor U8813 (N_8813,N_8627,N_8715);
and U8814 (N_8814,N_8798,N_8757);
or U8815 (N_8815,N_8696,N_8655);
xnor U8816 (N_8816,N_8644,N_8744);
nand U8817 (N_8817,N_8783,N_8781);
and U8818 (N_8818,N_8742,N_8725);
nor U8819 (N_8819,N_8611,N_8692);
nand U8820 (N_8820,N_8703,N_8641);
nand U8821 (N_8821,N_8784,N_8698);
or U8822 (N_8822,N_8648,N_8671);
xor U8823 (N_8823,N_8700,N_8669);
and U8824 (N_8824,N_8616,N_8699);
xor U8825 (N_8825,N_8664,N_8777);
nand U8826 (N_8826,N_8701,N_8720);
nor U8827 (N_8827,N_8619,N_8746);
and U8828 (N_8828,N_8656,N_8758);
or U8829 (N_8829,N_8755,N_8740);
xor U8830 (N_8830,N_8736,N_8728);
or U8831 (N_8831,N_8799,N_8674);
nor U8832 (N_8832,N_8617,N_8710);
or U8833 (N_8833,N_8687,N_8652);
or U8834 (N_8834,N_8646,N_8661);
nor U8835 (N_8835,N_8704,N_8603);
nand U8836 (N_8836,N_8675,N_8709);
and U8837 (N_8837,N_8748,N_8794);
xnor U8838 (N_8838,N_8733,N_8637);
nand U8839 (N_8839,N_8775,N_8711);
nand U8840 (N_8840,N_8787,N_8706);
nand U8841 (N_8841,N_8778,N_8763);
nand U8842 (N_8842,N_8705,N_8718);
xnor U8843 (N_8843,N_8750,N_8660);
xor U8844 (N_8844,N_8738,N_8719);
or U8845 (N_8845,N_8647,N_8795);
and U8846 (N_8846,N_8737,N_8691);
and U8847 (N_8847,N_8632,N_8640);
or U8848 (N_8848,N_8739,N_8677);
and U8849 (N_8849,N_8639,N_8673);
xor U8850 (N_8850,N_8731,N_8724);
or U8851 (N_8851,N_8765,N_8768);
or U8852 (N_8852,N_8645,N_8658);
nand U8853 (N_8853,N_8779,N_8628);
nand U8854 (N_8854,N_8624,N_8723);
xnor U8855 (N_8855,N_8657,N_8741);
nand U8856 (N_8856,N_8662,N_8756);
nor U8857 (N_8857,N_8633,N_8614);
nor U8858 (N_8858,N_8659,N_8688);
nand U8859 (N_8859,N_8749,N_8714);
xor U8860 (N_8860,N_8605,N_8672);
or U8861 (N_8861,N_8623,N_8625);
and U8862 (N_8862,N_8681,N_8631);
xnor U8863 (N_8863,N_8789,N_8670);
nand U8864 (N_8864,N_8643,N_8676);
nand U8865 (N_8865,N_8730,N_8707);
xor U8866 (N_8866,N_8782,N_8620);
nor U8867 (N_8867,N_8769,N_8612);
nand U8868 (N_8868,N_8774,N_8721);
nand U8869 (N_8869,N_8604,N_8679);
xnor U8870 (N_8870,N_8729,N_8735);
xnor U8871 (N_8871,N_8792,N_8665);
or U8872 (N_8872,N_8754,N_8642);
or U8873 (N_8873,N_8638,N_8797);
xnor U8874 (N_8874,N_8772,N_8651);
or U8875 (N_8875,N_8654,N_8686);
nand U8876 (N_8876,N_8602,N_8732);
nor U8877 (N_8877,N_8694,N_8667);
xor U8878 (N_8878,N_8663,N_8745);
xnor U8879 (N_8879,N_8712,N_8770);
xor U8880 (N_8880,N_8793,N_8635);
nor U8881 (N_8881,N_8708,N_8609);
and U8882 (N_8882,N_8689,N_8610);
nand U8883 (N_8883,N_8618,N_8759);
xnor U8884 (N_8884,N_8630,N_8767);
nor U8885 (N_8885,N_8780,N_8785);
nor U8886 (N_8886,N_8786,N_8751);
or U8887 (N_8887,N_8613,N_8790);
nand U8888 (N_8888,N_8634,N_8717);
nand U8889 (N_8889,N_8601,N_8743);
or U8890 (N_8890,N_8766,N_8734);
nor U8891 (N_8891,N_8796,N_8683);
nand U8892 (N_8892,N_8771,N_8606);
and U8893 (N_8893,N_8629,N_8615);
nor U8894 (N_8894,N_8760,N_8666);
or U8895 (N_8895,N_8695,N_8684);
xnor U8896 (N_8896,N_8600,N_8762);
nor U8897 (N_8897,N_8653,N_8753);
xor U8898 (N_8898,N_8693,N_8702);
and U8899 (N_8899,N_8636,N_8764);
and U8900 (N_8900,N_8767,N_8723);
xnor U8901 (N_8901,N_8614,N_8768);
nor U8902 (N_8902,N_8711,N_8699);
and U8903 (N_8903,N_8634,N_8631);
xor U8904 (N_8904,N_8749,N_8777);
and U8905 (N_8905,N_8615,N_8778);
nand U8906 (N_8906,N_8607,N_8773);
nand U8907 (N_8907,N_8706,N_8612);
nand U8908 (N_8908,N_8620,N_8759);
or U8909 (N_8909,N_8775,N_8695);
nor U8910 (N_8910,N_8773,N_8620);
or U8911 (N_8911,N_8662,N_8619);
nor U8912 (N_8912,N_8737,N_8640);
and U8913 (N_8913,N_8749,N_8707);
and U8914 (N_8914,N_8654,N_8758);
nor U8915 (N_8915,N_8603,N_8765);
nand U8916 (N_8916,N_8747,N_8786);
nor U8917 (N_8917,N_8781,N_8738);
or U8918 (N_8918,N_8694,N_8715);
xnor U8919 (N_8919,N_8687,N_8682);
or U8920 (N_8920,N_8616,N_8657);
xor U8921 (N_8921,N_8624,N_8772);
xnor U8922 (N_8922,N_8764,N_8768);
xor U8923 (N_8923,N_8764,N_8661);
nand U8924 (N_8924,N_8699,N_8685);
and U8925 (N_8925,N_8728,N_8609);
nor U8926 (N_8926,N_8619,N_8737);
nand U8927 (N_8927,N_8783,N_8797);
or U8928 (N_8928,N_8663,N_8765);
and U8929 (N_8929,N_8789,N_8685);
nor U8930 (N_8930,N_8713,N_8621);
and U8931 (N_8931,N_8775,N_8717);
nor U8932 (N_8932,N_8773,N_8775);
or U8933 (N_8933,N_8791,N_8634);
or U8934 (N_8934,N_8707,N_8754);
and U8935 (N_8935,N_8744,N_8733);
nand U8936 (N_8936,N_8795,N_8783);
nand U8937 (N_8937,N_8650,N_8759);
and U8938 (N_8938,N_8727,N_8627);
nor U8939 (N_8939,N_8741,N_8659);
and U8940 (N_8940,N_8792,N_8744);
or U8941 (N_8941,N_8606,N_8717);
nand U8942 (N_8942,N_8736,N_8758);
nor U8943 (N_8943,N_8667,N_8793);
nor U8944 (N_8944,N_8635,N_8733);
and U8945 (N_8945,N_8713,N_8706);
or U8946 (N_8946,N_8621,N_8684);
and U8947 (N_8947,N_8714,N_8665);
and U8948 (N_8948,N_8653,N_8742);
or U8949 (N_8949,N_8679,N_8769);
xor U8950 (N_8950,N_8654,N_8775);
or U8951 (N_8951,N_8684,N_8641);
nand U8952 (N_8952,N_8616,N_8682);
or U8953 (N_8953,N_8780,N_8611);
xnor U8954 (N_8954,N_8768,N_8694);
and U8955 (N_8955,N_8799,N_8652);
nor U8956 (N_8956,N_8712,N_8648);
and U8957 (N_8957,N_8637,N_8687);
nand U8958 (N_8958,N_8602,N_8779);
and U8959 (N_8959,N_8782,N_8621);
and U8960 (N_8960,N_8752,N_8668);
xnor U8961 (N_8961,N_8623,N_8720);
nor U8962 (N_8962,N_8733,N_8756);
nand U8963 (N_8963,N_8774,N_8717);
and U8964 (N_8964,N_8769,N_8798);
xnor U8965 (N_8965,N_8661,N_8666);
nor U8966 (N_8966,N_8697,N_8606);
and U8967 (N_8967,N_8609,N_8658);
nor U8968 (N_8968,N_8724,N_8707);
xnor U8969 (N_8969,N_8784,N_8666);
nand U8970 (N_8970,N_8631,N_8644);
and U8971 (N_8971,N_8643,N_8690);
nor U8972 (N_8972,N_8685,N_8710);
and U8973 (N_8973,N_8782,N_8647);
or U8974 (N_8974,N_8718,N_8782);
nor U8975 (N_8975,N_8678,N_8613);
or U8976 (N_8976,N_8622,N_8759);
or U8977 (N_8977,N_8796,N_8627);
nor U8978 (N_8978,N_8686,N_8727);
or U8979 (N_8979,N_8721,N_8748);
nand U8980 (N_8980,N_8748,N_8706);
nand U8981 (N_8981,N_8703,N_8727);
and U8982 (N_8982,N_8778,N_8798);
xnor U8983 (N_8983,N_8720,N_8677);
and U8984 (N_8984,N_8654,N_8607);
or U8985 (N_8985,N_8677,N_8606);
nand U8986 (N_8986,N_8618,N_8728);
xnor U8987 (N_8987,N_8784,N_8660);
and U8988 (N_8988,N_8725,N_8644);
xnor U8989 (N_8989,N_8680,N_8620);
and U8990 (N_8990,N_8761,N_8788);
and U8991 (N_8991,N_8625,N_8658);
or U8992 (N_8992,N_8638,N_8627);
and U8993 (N_8993,N_8796,N_8649);
and U8994 (N_8994,N_8687,N_8677);
nor U8995 (N_8995,N_8771,N_8693);
xnor U8996 (N_8996,N_8661,N_8656);
nor U8997 (N_8997,N_8783,N_8784);
or U8998 (N_8998,N_8628,N_8719);
nand U8999 (N_8999,N_8671,N_8709);
nor U9000 (N_9000,N_8863,N_8854);
nor U9001 (N_9001,N_8913,N_8933);
xor U9002 (N_9002,N_8949,N_8941);
xor U9003 (N_9003,N_8864,N_8812);
or U9004 (N_9004,N_8881,N_8829);
and U9005 (N_9005,N_8845,N_8905);
or U9006 (N_9006,N_8887,N_8877);
nor U9007 (N_9007,N_8936,N_8960);
and U9008 (N_9008,N_8934,N_8873);
xnor U9009 (N_9009,N_8850,N_8879);
xnor U9010 (N_9010,N_8954,N_8899);
and U9011 (N_9011,N_8971,N_8807);
xnor U9012 (N_9012,N_8825,N_8875);
and U9013 (N_9013,N_8912,N_8952);
and U9014 (N_9014,N_8803,N_8974);
xor U9015 (N_9015,N_8802,N_8922);
or U9016 (N_9016,N_8862,N_8946);
and U9017 (N_9017,N_8820,N_8921);
nand U9018 (N_9018,N_8866,N_8896);
nand U9019 (N_9019,N_8898,N_8958);
and U9020 (N_9020,N_8824,N_8888);
nor U9021 (N_9021,N_8830,N_8837);
nor U9022 (N_9022,N_8851,N_8943);
xnor U9023 (N_9023,N_8973,N_8843);
xor U9024 (N_9024,N_8935,N_8998);
xor U9025 (N_9025,N_8925,N_8930);
and U9026 (N_9026,N_8882,N_8852);
and U9027 (N_9027,N_8840,N_8844);
and U9028 (N_9028,N_8932,N_8969);
or U9029 (N_9029,N_8906,N_8948);
or U9030 (N_9030,N_8815,N_8811);
nand U9031 (N_9031,N_8865,N_8848);
xnor U9032 (N_9032,N_8907,N_8931);
xnor U9033 (N_9033,N_8904,N_8956);
nand U9034 (N_9034,N_8859,N_8939);
or U9035 (N_9035,N_8834,N_8983);
nand U9036 (N_9036,N_8991,N_8858);
nand U9037 (N_9037,N_8953,N_8918);
or U9038 (N_9038,N_8981,N_8989);
and U9039 (N_9039,N_8914,N_8984);
and U9040 (N_9040,N_8919,N_8846);
xor U9041 (N_9041,N_8920,N_8823);
nand U9042 (N_9042,N_8996,N_8808);
nand U9043 (N_9043,N_8909,N_8861);
nor U9044 (N_9044,N_8841,N_8857);
nor U9045 (N_9045,N_8885,N_8988);
nand U9046 (N_9046,N_8810,N_8992);
nor U9047 (N_9047,N_8869,N_8979);
and U9048 (N_9048,N_8833,N_8860);
and U9049 (N_9049,N_8929,N_8978);
and U9050 (N_9050,N_8839,N_8901);
or U9051 (N_9051,N_8876,N_8892);
nand U9052 (N_9052,N_8856,N_8938);
xor U9053 (N_9053,N_8995,N_8801);
xor U9054 (N_9054,N_8962,N_8911);
nor U9055 (N_9055,N_8997,N_8975);
xnor U9056 (N_9056,N_8924,N_8902);
and U9057 (N_9057,N_8928,N_8970);
xor U9058 (N_9058,N_8806,N_8940);
and U9059 (N_9059,N_8822,N_8951);
and U9060 (N_9060,N_8836,N_8847);
nor U9061 (N_9061,N_8886,N_8985);
nor U9062 (N_9062,N_8967,N_8884);
nand U9063 (N_9063,N_8916,N_8966);
nor U9064 (N_9064,N_8872,N_8893);
or U9065 (N_9065,N_8923,N_8993);
xor U9066 (N_9066,N_8831,N_8900);
and U9067 (N_9067,N_8849,N_8968);
and U9068 (N_9068,N_8926,N_8957);
or U9069 (N_9069,N_8961,N_8842);
xor U9070 (N_9070,N_8999,N_8927);
nor U9071 (N_9071,N_8959,N_8963);
nor U9072 (N_9072,N_8838,N_8871);
nor U9073 (N_9073,N_8990,N_8942);
xnor U9074 (N_9074,N_8818,N_8878);
nand U9075 (N_9075,N_8821,N_8819);
xnor U9076 (N_9076,N_8870,N_8944);
nor U9077 (N_9077,N_8827,N_8977);
xor U9078 (N_9078,N_8835,N_8874);
nand U9079 (N_9079,N_8965,N_8800);
nor U9080 (N_9080,N_8950,N_8855);
nand U9081 (N_9081,N_8889,N_8964);
xor U9082 (N_9082,N_8814,N_8832);
or U9083 (N_9083,N_8982,N_8895);
nand U9084 (N_9084,N_8817,N_8890);
nor U9085 (N_9085,N_8937,N_8945);
and U9086 (N_9086,N_8880,N_8908);
xor U9087 (N_9087,N_8805,N_8903);
or U9088 (N_9088,N_8980,N_8994);
xnor U9089 (N_9089,N_8816,N_8976);
or U9090 (N_9090,N_8867,N_8809);
and U9091 (N_9091,N_8915,N_8987);
and U9092 (N_9092,N_8910,N_8986);
xnor U9093 (N_9093,N_8813,N_8883);
nand U9094 (N_9094,N_8868,N_8917);
xor U9095 (N_9095,N_8947,N_8853);
xor U9096 (N_9096,N_8955,N_8804);
xor U9097 (N_9097,N_8828,N_8972);
or U9098 (N_9098,N_8894,N_8891);
or U9099 (N_9099,N_8826,N_8897);
and U9100 (N_9100,N_8979,N_8834);
or U9101 (N_9101,N_8891,N_8908);
xnor U9102 (N_9102,N_8984,N_8943);
or U9103 (N_9103,N_8884,N_8929);
nor U9104 (N_9104,N_8966,N_8969);
nor U9105 (N_9105,N_8919,N_8840);
and U9106 (N_9106,N_8846,N_8941);
or U9107 (N_9107,N_8927,N_8923);
nand U9108 (N_9108,N_8924,N_8961);
nand U9109 (N_9109,N_8905,N_8968);
xnor U9110 (N_9110,N_8837,N_8937);
or U9111 (N_9111,N_8868,N_8878);
xor U9112 (N_9112,N_8970,N_8915);
or U9113 (N_9113,N_8823,N_8948);
nor U9114 (N_9114,N_8848,N_8962);
xor U9115 (N_9115,N_8927,N_8863);
or U9116 (N_9116,N_8911,N_8840);
and U9117 (N_9117,N_8855,N_8952);
nor U9118 (N_9118,N_8836,N_8880);
nor U9119 (N_9119,N_8938,N_8817);
xnor U9120 (N_9120,N_8864,N_8908);
nor U9121 (N_9121,N_8930,N_8938);
nor U9122 (N_9122,N_8922,N_8908);
or U9123 (N_9123,N_8915,N_8980);
or U9124 (N_9124,N_8935,N_8938);
xnor U9125 (N_9125,N_8903,N_8801);
xor U9126 (N_9126,N_8956,N_8984);
nor U9127 (N_9127,N_8976,N_8918);
xor U9128 (N_9128,N_8904,N_8995);
and U9129 (N_9129,N_8934,N_8870);
xnor U9130 (N_9130,N_8871,N_8978);
and U9131 (N_9131,N_8825,N_8814);
nor U9132 (N_9132,N_8903,N_8893);
nor U9133 (N_9133,N_8846,N_8910);
nand U9134 (N_9134,N_8991,N_8860);
nand U9135 (N_9135,N_8853,N_8907);
nand U9136 (N_9136,N_8822,N_8856);
nor U9137 (N_9137,N_8850,N_8939);
and U9138 (N_9138,N_8912,N_8905);
and U9139 (N_9139,N_8983,N_8838);
xnor U9140 (N_9140,N_8953,N_8920);
and U9141 (N_9141,N_8872,N_8982);
and U9142 (N_9142,N_8820,N_8851);
or U9143 (N_9143,N_8946,N_8823);
and U9144 (N_9144,N_8840,N_8855);
or U9145 (N_9145,N_8806,N_8980);
xor U9146 (N_9146,N_8880,N_8817);
nand U9147 (N_9147,N_8865,N_8887);
or U9148 (N_9148,N_8901,N_8902);
nand U9149 (N_9149,N_8829,N_8879);
xnor U9150 (N_9150,N_8921,N_8868);
nor U9151 (N_9151,N_8914,N_8826);
or U9152 (N_9152,N_8920,N_8892);
and U9153 (N_9153,N_8957,N_8959);
nor U9154 (N_9154,N_8810,N_8873);
or U9155 (N_9155,N_8945,N_8917);
and U9156 (N_9156,N_8842,N_8845);
nor U9157 (N_9157,N_8941,N_8936);
nand U9158 (N_9158,N_8996,N_8986);
nor U9159 (N_9159,N_8943,N_8964);
nand U9160 (N_9160,N_8946,N_8856);
or U9161 (N_9161,N_8952,N_8887);
and U9162 (N_9162,N_8911,N_8944);
or U9163 (N_9163,N_8961,N_8824);
nor U9164 (N_9164,N_8864,N_8961);
xor U9165 (N_9165,N_8904,N_8862);
xnor U9166 (N_9166,N_8961,N_8815);
nand U9167 (N_9167,N_8889,N_8824);
or U9168 (N_9168,N_8876,N_8812);
nor U9169 (N_9169,N_8952,N_8876);
and U9170 (N_9170,N_8881,N_8918);
and U9171 (N_9171,N_8907,N_8976);
and U9172 (N_9172,N_8862,N_8986);
and U9173 (N_9173,N_8901,N_8897);
and U9174 (N_9174,N_8911,N_8971);
nand U9175 (N_9175,N_8888,N_8918);
nand U9176 (N_9176,N_8830,N_8963);
and U9177 (N_9177,N_8955,N_8998);
nor U9178 (N_9178,N_8830,N_8992);
and U9179 (N_9179,N_8980,N_8981);
xnor U9180 (N_9180,N_8868,N_8823);
or U9181 (N_9181,N_8938,N_8975);
or U9182 (N_9182,N_8846,N_8804);
and U9183 (N_9183,N_8847,N_8920);
or U9184 (N_9184,N_8955,N_8841);
and U9185 (N_9185,N_8862,N_8811);
nand U9186 (N_9186,N_8979,N_8941);
xor U9187 (N_9187,N_8941,N_8851);
nor U9188 (N_9188,N_8824,N_8823);
xor U9189 (N_9189,N_8911,N_8844);
nor U9190 (N_9190,N_8906,N_8802);
or U9191 (N_9191,N_8999,N_8826);
nand U9192 (N_9192,N_8844,N_8908);
xor U9193 (N_9193,N_8800,N_8814);
nor U9194 (N_9194,N_8943,N_8959);
or U9195 (N_9195,N_8907,N_8868);
nand U9196 (N_9196,N_8861,N_8851);
nor U9197 (N_9197,N_8833,N_8847);
xnor U9198 (N_9198,N_8978,N_8889);
or U9199 (N_9199,N_8874,N_8879);
xor U9200 (N_9200,N_9092,N_9187);
and U9201 (N_9201,N_9188,N_9090);
and U9202 (N_9202,N_9064,N_9134);
or U9203 (N_9203,N_9095,N_9145);
and U9204 (N_9204,N_9127,N_9091);
or U9205 (N_9205,N_9070,N_9108);
nor U9206 (N_9206,N_9129,N_9085);
or U9207 (N_9207,N_9196,N_9055);
and U9208 (N_9208,N_9184,N_9030);
nand U9209 (N_9209,N_9123,N_9191);
or U9210 (N_9210,N_9156,N_9050);
or U9211 (N_9211,N_9083,N_9101);
and U9212 (N_9212,N_9149,N_9186);
xor U9213 (N_9213,N_9107,N_9160);
nand U9214 (N_9214,N_9148,N_9049);
nor U9215 (N_9215,N_9036,N_9109);
nand U9216 (N_9216,N_9125,N_9044);
and U9217 (N_9217,N_9040,N_9023);
nor U9218 (N_9218,N_9166,N_9118);
and U9219 (N_9219,N_9024,N_9111);
and U9220 (N_9220,N_9000,N_9150);
nand U9221 (N_9221,N_9185,N_9079);
and U9222 (N_9222,N_9112,N_9159);
nand U9223 (N_9223,N_9088,N_9133);
or U9224 (N_9224,N_9047,N_9193);
and U9225 (N_9225,N_9154,N_9042);
nand U9226 (N_9226,N_9155,N_9096);
xor U9227 (N_9227,N_9157,N_9067);
or U9228 (N_9228,N_9080,N_9099);
nor U9229 (N_9229,N_9132,N_9197);
or U9230 (N_9230,N_9128,N_9152);
or U9231 (N_9231,N_9183,N_9025);
or U9232 (N_9232,N_9177,N_9068);
xnor U9233 (N_9233,N_9169,N_9075);
nor U9234 (N_9234,N_9175,N_9142);
nand U9235 (N_9235,N_9027,N_9006);
nand U9236 (N_9236,N_9003,N_9009);
nor U9237 (N_9237,N_9114,N_9135);
nand U9238 (N_9238,N_9051,N_9190);
xor U9239 (N_9239,N_9063,N_9181);
and U9240 (N_9240,N_9043,N_9174);
nor U9241 (N_9241,N_9102,N_9141);
xor U9242 (N_9242,N_9052,N_9192);
and U9243 (N_9243,N_9117,N_9165);
or U9244 (N_9244,N_9057,N_9097);
or U9245 (N_9245,N_9062,N_9010);
xor U9246 (N_9246,N_9153,N_9119);
nand U9247 (N_9247,N_9140,N_9147);
nor U9248 (N_9248,N_9176,N_9124);
and U9249 (N_9249,N_9126,N_9167);
xnor U9250 (N_9250,N_9198,N_9113);
xor U9251 (N_9251,N_9131,N_9069);
and U9252 (N_9252,N_9066,N_9029);
and U9253 (N_9253,N_9077,N_9081);
nor U9254 (N_9254,N_9172,N_9094);
or U9255 (N_9255,N_9106,N_9104);
nor U9256 (N_9256,N_9001,N_9026);
nor U9257 (N_9257,N_9121,N_9005);
nor U9258 (N_9258,N_9138,N_9046);
and U9259 (N_9259,N_9008,N_9130);
and U9260 (N_9260,N_9110,N_9098);
xnor U9261 (N_9261,N_9054,N_9011);
and U9262 (N_9262,N_9059,N_9189);
or U9263 (N_9263,N_9161,N_9032);
nor U9264 (N_9264,N_9137,N_9194);
and U9265 (N_9265,N_9122,N_9093);
or U9266 (N_9266,N_9028,N_9073);
or U9267 (N_9267,N_9017,N_9022);
xnor U9268 (N_9268,N_9144,N_9173);
xor U9269 (N_9269,N_9164,N_9171);
xor U9270 (N_9270,N_9021,N_9012);
nor U9271 (N_9271,N_9045,N_9072);
xnor U9272 (N_9272,N_9058,N_9105);
nand U9273 (N_9273,N_9016,N_9163);
nand U9274 (N_9274,N_9020,N_9084);
xor U9275 (N_9275,N_9041,N_9078);
and U9276 (N_9276,N_9004,N_9116);
or U9277 (N_9277,N_9033,N_9007);
nand U9278 (N_9278,N_9162,N_9031);
xor U9279 (N_9279,N_9087,N_9076);
and U9280 (N_9280,N_9139,N_9086);
nand U9281 (N_9281,N_9168,N_9143);
and U9282 (N_9282,N_9089,N_9179);
nor U9283 (N_9283,N_9019,N_9074);
and U9284 (N_9284,N_9199,N_9120);
and U9285 (N_9285,N_9180,N_9034);
and U9286 (N_9286,N_9048,N_9061);
nand U9287 (N_9287,N_9035,N_9018);
xor U9288 (N_9288,N_9170,N_9065);
and U9289 (N_9289,N_9002,N_9053);
and U9290 (N_9290,N_9136,N_9014);
nand U9291 (N_9291,N_9013,N_9037);
xnor U9292 (N_9292,N_9056,N_9158);
or U9293 (N_9293,N_9146,N_9103);
xor U9294 (N_9294,N_9071,N_9038);
or U9295 (N_9295,N_9115,N_9060);
and U9296 (N_9296,N_9039,N_9182);
or U9297 (N_9297,N_9178,N_9082);
nand U9298 (N_9298,N_9015,N_9151);
nor U9299 (N_9299,N_9100,N_9195);
xor U9300 (N_9300,N_9037,N_9003);
and U9301 (N_9301,N_9197,N_9050);
and U9302 (N_9302,N_9000,N_9066);
and U9303 (N_9303,N_9180,N_9130);
xnor U9304 (N_9304,N_9128,N_9090);
or U9305 (N_9305,N_9118,N_9058);
and U9306 (N_9306,N_9143,N_9163);
nor U9307 (N_9307,N_9082,N_9087);
or U9308 (N_9308,N_9109,N_9078);
or U9309 (N_9309,N_9071,N_9150);
nor U9310 (N_9310,N_9027,N_9064);
nand U9311 (N_9311,N_9104,N_9035);
xnor U9312 (N_9312,N_9036,N_9072);
or U9313 (N_9313,N_9161,N_9196);
or U9314 (N_9314,N_9191,N_9050);
or U9315 (N_9315,N_9032,N_9084);
nand U9316 (N_9316,N_9056,N_9101);
and U9317 (N_9317,N_9011,N_9159);
nand U9318 (N_9318,N_9168,N_9014);
nor U9319 (N_9319,N_9097,N_9151);
nor U9320 (N_9320,N_9189,N_9076);
nor U9321 (N_9321,N_9122,N_9143);
nand U9322 (N_9322,N_9144,N_9131);
nand U9323 (N_9323,N_9020,N_9111);
nor U9324 (N_9324,N_9079,N_9093);
or U9325 (N_9325,N_9043,N_9178);
xor U9326 (N_9326,N_9115,N_9185);
xnor U9327 (N_9327,N_9192,N_9181);
xor U9328 (N_9328,N_9078,N_9108);
nor U9329 (N_9329,N_9132,N_9150);
or U9330 (N_9330,N_9094,N_9045);
and U9331 (N_9331,N_9045,N_9195);
or U9332 (N_9332,N_9160,N_9045);
nor U9333 (N_9333,N_9094,N_9000);
nand U9334 (N_9334,N_9093,N_9130);
and U9335 (N_9335,N_9133,N_9161);
and U9336 (N_9336,N_9094,N_9153);
nor U9337 (N_9337,N_9137,N_9125);
nor U9338 (N_9338,N_9038,N_9065);
nand U9339 (N_9339,N_9038,N_9102);
and U9340 (N_9340,N_9069,N_9038);
nor U9341 (N_9341,N_9020,N_9058);
xnor U9342 (N_9342,N_9035,N_9134);
nand U9343 (N_9343,N_9102,N_9136);
or U9344 (N_9344,N_9075,N_9104);
or U9345 (N_9345,N_9095,N_9049);
and U9346 (N_9346,N_9162,N_9112);
nor U9347 (N_9347,N_9143,N_9018);
nor U9348 (N_9348,N_9026,N_9150);
or U9349 (N_9349,N_9192,N_9167);
xor U9350 (N_9350,N_9046,N_9126);
or U9351 (N_9351,N_9126,N_9069);
and U9352 (N_9352,N_9179,N_9083);
or U9353 (N_9353,N_9126,N_9128);
or U9354 (N_9354,N_9092,N_9058);
and U9355 (N_9355,N_9195,N_9161);
or U9356 (N_9356,N_9079,N_9125);
xor U9357 (N_9357,N_9186,N_9038);
or U9358 (N_9358,N_9008,N_9136);
and U9359 (N_9359,N_9185,N_9114);
nor U9360 (N_9360,N_9183,N_9017);
or U9361 (N_9361,N_9183,N_9152);
xor U9362 (N_9362,N_9199,N_9093);
nand U9363 (N_9363,N_9170,N_9097);
nand U9364 (N_9364,N_9145,N_9137);
or U9365 (N_9365,N_9119,N_9089);
nor U9366 (N_9366,N_9177,N_9171);
nand U9367 (N_9367,N_9158,N_9123);
xnor U9368 (N_9368,N_9009,N_9126);
xor U9369 (N_9369,N_9065,N_9067);
nor U9370 (N_9370,N_9047,N_9060);
and U9371 (N_9371,N_9061,N_9080);
nand U9372 (N_9372,N_9147,N_9199);
or U9373 (N_9373,N_9107,N_9010);
nor U9374 (N_9374,N_9007,N_9081);
nand U9375 (N_9375,N_9110,N_9118);
and U9376 (N_9376,N_9124,N_9054);
xor U9377 (N_9377,N_9105,N_9149);
or U9378 (N_9378,N_9005,N_9031);
or U9379 (N_9379,N_9038,N_9131);
nand U9380 (N_9380,N_9136,N_9164);
or U9381 (N_9381,N_9193,N_9014);
nor U9382 (N_9382,N_9168,N_9179);
xnor U9383 (N_9383,N_9058,N_9010);
nor U9384 (N_9384,N_9042,N_9007);
or U9385 (N_9385,N_9104,N_9082);
or U9386 (N_9386,N_9086,N_9020);
nor U9387 (N_9387,N_9128,N_9191);
nand U9388 (N_9388,N_9042,N_9108);
xor U9389 (N_9389,N_9073,N_9022);
xnor U9390 (N_9390,N_9057,N_9104);
and U9391 (N_9391,N_9048,N_9169);
nor U9392 (N_9392,N_9164,N_9078);
xor U9393 (N_9393,N_9172,N_9052);
nand U9394 (N_9394,N_9128,N_9147);
nor U9395 (N_9395,N_9172,N_9169);
and U9396 (N_9396,N_9008,N_9070);
or U9397 (N_9397,N_9115,N_9148);
xnor U9398 (N_9398,N_9090,N_9110);
or U9399 (N_9399,N_9148,N_9067);
and U9400 (N_9400,N_9208,N_9283);
nand U9401 (N_9401,N_9348,N_9275);
nor U9402 (N_9402,N_9399,N_9333);
nand U9403 (N_9403,N_9280,N_9382);
nand U9404 (N_9404,N_9244,N_9386);
nor U9405 (N_9405,N_9373,N_9293);
nor U9406 (N_9406,N_9320,N_9344);
nor U9407 (N_9407,N_9288,N_9314);
or U9408 (N_9408,N_9266,N_9286);
or U9409 (N_9409,N_9254,N_9218);
nor U9410 (N_9410,N_9287,N_9379);
nor U9411 (N_9411,N_9250,N_9271);
nand U9412 (N_9412,N_9398,N_9324);
or U9413 (N_9413,N_9229,N_9204);
xnor U9414 (N_9414,N_9256,N_9307);
or U9415 (N_9415,N_9397,N_9313);
nor U9416 (N_9416,N_9247,N_9265);
or U9417 (N_9417,N_9235,N_9294);
xor U9418 (N_9418,N_9239,N_9316);
and U9419 (N_9419,N_9301,N_9270);
nor U9420 (N_9420,N_9248,N_9345);
nand U9421 (N_9421,N_9268,N_9364);
and U9422 (N_9422,N_9396,N_9310);
or U9423 (N_9423,N_9380,N_9299);
or U9424 (N_9424,N_9363,N_9231);
nor U9425 (N_9425,N_9371,N_9361);
xor U9426 (N_9426,N_9355,N_9356);
nor U9427 (N_9427,N_9298,N_9216);
nand U9428 (N_9428,N_9325,N_9230);
nand U9429 (N_9429,N_9335,N_9260);
or U9430 (N_9430,N_9261,N_9330);
or U9431 (N_9431,N_9353,N_9370);
or U9432 (N_9432,N_9360,N_9336);
nand U9433 (N_9433,N_9352,N_9211);
and U9434 (N_9434,N_9362,N_9385);
nand U9435 (N_9435,N_9341,N_9289);
xor U9436 (N_9436,N_9224,N_9205);
nor U9437 (N_9437,N_9296,N_9255);
nand U9438 (N_9438,N_9259,N_9291);
or U9439 (N_9439,N_9308,N_9232);
nor U9440 (N_9440,N_9372,N_9359);
nor U9441 (N_9441,N_9318,N_9309);
xor U9442 (N_9442,N_9358,N_9241);
xnor U9443 (N_9443,N_9262,N_9213);
nor U9444 (N_9444,N_9392,N_9311);
nor U9445 (N_9445,N_9393,N_9267);
nand U9446 (N_9446,N_9389,N_9217);
nand U9447 (N_9447,N_9367,N_9365);
nand U9448 (N_9448,N_9338,N_9391);
or U9449 (N_9449,N_9209,N_9378);
xor U9450 (N_9450,N_9278,N_9273);
xor U9451 (N_9451,N_9376,N_9321);
nand U9452 (N_9452,N_9395,N_9282);
nand U9453 (N_9453,N_9292,N_9245);
xor U9454 (N_9454,N_9253,N_9374);
nand U9455 (N_9455,N_9305,N_9368);
or U9456 (N_9456,N_9334,N_9219);
nand U9457 (N_9457,N_9203,N_9236);
nor U9458 (N_9458,N_9349,N_9327);
nand U9459 (N_9459,N_9332,N_9306);
or U9460 (N_9460,N_9300,N_9221);
and U9461 (N_9461,N_9212,N_9234);
nand U9462 (N_9462,N_9274,N_9206);
and U9463 (N_9463,N_9243,N_9375);
or U9464 (N_9464,N_9202,N_9295);
xor U9465 (N_9465,N_9329,N_9228);
and U9466 (N_9466,N_9388,N_9328);
and U9467 (N_9467,N_9279,N_9331);
nor U9468 (N_9468,N_9264,N_9277);
and U9469 (N_9469,N_9233,N_9290);
xor U9470 (N_9470,N_9366,N_9215);
or U9471 (N_9471,N_9201,N_9227);
nand U9472 (N_9472,N_9257,N_9303);
or U9473 (N_9473,N_9323,N_9226);
xor U9474 (N_9474,N_9272,N_9276);
xnor U9475 (N_9475,N_9357,N_9319);
and U9476 (N_9476,N_9258,N_9214);
or U9477 (N_9477,N_9346,N_9390);
nor U9478 (N_9478,N_9238,N_9284);
and U9479 (N_9479,N_9285,N_9315);
nor U9480 (N_9480,N_9322,N_9312);
or U9481 (N_9481,N_9377,N_9225);
and U9482 (N_9482,N_9246,N_9297);
nand U9483 (N_9483,N_9317,N_9340);
xnor U9484 (N_9484,N_9251,N_9351);
or U9485 (N_9485,N_9347,N_9339);
xnor U9486 (N_9486,N_9343,N_9207);
xnor U9487 (N_9487,N_9383,N_9220);
or U9488 (N_9488,N_9242,N_9249);
or U9489 (N_9489,N_9237,N_9394);
nand U9490 (N_9490,N_9387,N_9200);
xnor U9491 (N_9491,N_9222,N_9223);
and U9492 (N_9492,N_9302,N_9281);
or U9493 (N_9493,N_9384,N_9210);
nor U9494 (N_9494,N_9326,N_9337);
nor U9495 (N_9495,N_9269,N_9381);
and U9496 (N_9496,N_9369,N_9342);
nor U9497 (N_9497,N_9240,N_9252);
nor U9498 (N_9498,N_9350,N_9304);
nand U9499 (N_9499,N_9263,N_9354);
nor U9500 (N_9500,N_9319,N_9236);
or U9501 (N_9501,N_9389,N_9224);
and U9502 (N_9502,N_9231,N_9225);
or U9503 (N_9503,N_9294,N_9253);
nand U9504 (N_9504,N_9213,N_9258);
nand U9505 (N_9505,N_9251,N_9332);
xor U9506 (N_9506,N_9256,N_9285);
or U9507 (N_9507,N_9240,N_9320);
xnor U9508 (N_9508,N_9224,N_9346);
nor U9509 (N_9509,N_9214,N_9320);
and U9510 (N_9510,N_9324,N_9314);
xnor U9511 (N_9511,N_9210,N_9325);
xnor U9512 (N_9512,N_9347,N_9271);
nor U9513 (N_9513,N_9355,N_9344);
nand U9514 (N_9514,N_9291,N_9344);
nor U9515 (N_9515,N_9333,N_9238);
nand U9516 (N_9516,N_9266,N_9378);
and U9517 (N_9517,N_9219,N_9200);
xor U9518 (N_9518,N_9358,N_9202);
nor U9519 (N_9519,N_9288,N_9315);
nand U9520 (N_9520,N_9372,N_9237);
nor U9521 (N_9521,N_9256,N_9316);
or U9522 (N_9522,N_9345,N_9227);
or U9523 (N_9523,N_9385,N_9228);
xnor U9524 (N_9524,N_9373,N_9205);
xor U9525 (N_9525,N_9223,N_9309);
or U9526 (N_9526,N_9344,N_9324);
or U9527 (N_9527,N_9312,N_9243);
nor U9528 (N_9528,N_9304,N_9255);
and U9529 (N_9529,N_9369,N_9284);
xnor U9530 (N_9530,N_9366,N_9290);
or U9531 (N_9531,N_9336,N_9242);
nand U9532 (N_9532,N_9371,N_9379);
or U9533 (N_9533,N_9364,N_9223);
or U9534 (N_9534,N_9211,N_9267);
nand U9535 (N_9535,N_9221,N_9261);
or U9536 (N_9536,N_9344,N_9257);
xnor U9537 (N_9537,N_9220,N_9238);
nor U9538 (N_9538,N_9202,N_9336);
and U9539 (N_9539,N_9393,N_9264);
and U9540 (N_9540,N_9359,N_9284);
nand U9541 (N_9541,N_9270,N_9380);
nand U9542 (N_9542,N_9353,N_9364);
and U9543 (N_9543,N_9223,N_9285);
xor U9544 (N_9544,N_9275,N_9305);
nor U9545 (N_9545,N_9359,N_9304);
and U9546 (N_9546,N_9385,N_9235);
and U9547 (N_9547,N_9223,N_9270);
nand U9548 (N_9548,N_9341,N_9316);
nand U9549 (N_9549,N_9384,N_9325);
or U9550 (N_9550,N_9334,N_9341);
or U9551 (N_9551,N_9389,N_9386);
nor U9552 (N_9552,N_9276,N_9234);
or U9553 (N_9553,N_9212,N_9368);
nor U9554 (N_9554,N_9210,N_9394);
nor U9555 (N_9555,N_9268,N_9231);
nor U9556 (N_9556,N_9339,N_9295);
nand U9557 (N_9557,N_9339,N_9374);
or U9558 (N_9558,N_9250,N_9368);
nor U9559 (N_9559,N_9243,N_9322);
and U9560 (N_9560,N_9261,N_9306);
or U9561 (N_9561,N_9206,N_9397);
and U9562 (N_9562,N_9371,N_9261);
nor U9563 (N_9563,N_9330,N_9347);
or U9564 (N_9564,N_9241,N_9305);
nand U9565 (N_9565,N_9395,N_9271);
nand U9566 (N_9566,N_9243,N_9291);
xnor U9567 (N_9567,N_9309,N_9225);
and U9568 (N_9568,N_9271,N_9233);
or U9569 (N_9569,N_9344,N_9249);
and U9570 (N_9570,N_9253,N_9248);
nor U9571 (N_9571,N_9215,N_9208);
nand U9572 (N_9572,N_9246,N_9307);
and U9573 (N_9573,N_9384,N_9324);
and U9574 (N_9574,N_9308,N_9215);
and U9575 (N_9575,N_9320,N_9298);
nor U9576 (N_9576,N_9303,N_9282);
nand U9577 (N_9577,N_9276,N_9285);
nand U9578 (N_9578,N_9355,N_9308);
xor U9579 (N_9579,N_9351,N_9338);
xor U9580 (N_9580,N_9307,N_9226);
and U9581 (N_9581,N_9223,N_9322);
nand U9582 (N_9582,N_9279,N_9205);
nor U9583 (N_9583,N_9309,N_9342);
xnor U9584 (N_9584,N_9393,N_9271);
nor U9585 (N_9585,N_9273,N_9330);
and U9586 (N_9586,N_9298,N_9277);
or U9587 (N_9587,N_9349,N_9215);
nand U9588 (N_9588,N_9298,N_9212);
and U9589 (N_9589,N_9331,N_9249);
nand U9590 (N_9590,N_9221,N_9280);
xor U9591 (N_9591,N_9319,N_9358);
or U9592 (N_9592,N_9284,N_9389);
or U9593 (N_9593,N_9230,N_9338);
nand U9594 (N_9594,N_9374,N_9231);
nor U9595 (N_9595,N_9259,N_9211);
and U9596 (N_9596,N_9362,N_9349);
xnor U9597 (N_9597,N_9391,N_9273);
nand U9598 (N_9598,N_9247,N_9390);
nor U9599 (N_9599,N_9247,N_9248);
nand U9600 (N_9600,N_9561,N_9531);
nand U9601 (N_9601,N_9405,N_9578);
xnor U9602 (N_9602,N_9476,N_9463);
or U9603 (N_9603,N_9492,N_9552);
xnor U9604 (N_9604,N_9536,N_9553);
xnor U9605 (N_9605,N_9439,N_9477);
or U9606 (N_9606,N_9440,N_9436);
or U9607 (N_9607,N_9462,N_9438);
and U9608 (N_9608,N_9448,N_9538);
nor U9609 (N_9609,N_9425,N_9426);
nor U9610 (N_9610,N_9489,N_9595);
xor U9611 (N_9611,N_9550,N_9482);
nand U9612 (N_9612,N_9430,N_9415);
nand U9613 (N_9613,N_9576,N_9461);
or U9614 (N_9614,N_9521,N_9442);
xnor U9615 (N_9615,N_9484,N_9500);
and U9616 (N_9616,N_9487,N_9472);
nand U9617 (N_9617,N_9534,N_9403);
xor U9618 (N_9618,N_9475,N_9429);
nor U9619 (N_9619,N_9474,N_9456);
nand U9620 (N_9620,N_9517,N_9596);
or U9621 (N_9621,N_9404,N_9557);
nor U9622 (N_9622,N_9478,N_9593);
xor U9623 (N_9623,N_9573,N_9453);
xor U9624 (N_9624,N_9490,N_9541);
and U9625 (N_9625,N_9530,N_9514);
nand U9626 (N_9626,N_9592,N_9413);
or U9627 (N_9627,N_9410,N_9519);
and U9628 (N_9628,N_9409,N_9591);
or U9629 (N_9629,N_9495,N_9582);
nand U9630 (N_9630,N_9427,N_9537);
nor U9631 (N_9631,N_9516,N_9542);
nand U9632 (N_9632,N_9509,N_9549);
and U9633 (N_9633,N_9400,N_9451);
xnor U9634 (N_9634,N_9527,N_9547);
nor U9635 (N_9635,N_9554,N_9486);
xnor U9636 (N_9636,N_9572,N_9424);
or U9637 (N_9637,N_9444,N_9598);
nand U9638 (N_9638,N_9523,N_9544);
xor U9639 (N_9639,N_9433,N_9597);
nor U9640 (N_9640,N_9567,N_9432);
xor U9641 (N_9641,N_9466,N_9590);
nand U9642 (N_9642,N_9491,N_9445);
or U9643 (N_9643,N_9513,N_9459);
nor U9644 (N_9644,N_9434,N_9471);
and U9645 (N_9645,N_9498,N_9455);
nand U9646 (N_9646,N_9412,N_9418);
xor U9647 (N_9647,N_9570,N_9589);
xor U9648 (N_9648,N_9422,N_9574);
nor U9649 (N_9649,N_9560,N_9460);
or U9650 (N_9650,N_9506,N_9511);
or U9651 (N_9651,N_9454,N_9581);
and U9652 (N_9652,N_9555,N_9556);
or U9653 (N_9653,N_9579,N_9497);
nand U9654 (N_9654,N_9473,N_9571);
or U9655 (N_9655,N_9449,N_9457);
xor U9656 (N_9656,N_9407,N_9564);
xor U9657 (N_9657,N_9479,N_9435);
nor U9658 (N_9658,N_9488,N_9518);
nor U9659 (N_9659,N_9577,N_9529);
xnor U9660 (N_9660,N_9452,N_9522);
nor U9661 (N_9661,N_9599,N_9526);
or U9662 (N_9662,N_9512,N_9467);
nand U9663 (N_9663,N_9481,N_9569);
nand U9664 (N_9664,N_9594,N_9406);
xnor U9665 (N_9665,N_9525,N_9414);
nor U9666 (N_9666,N_9416,N_9545);
xnor U9667 (N_9667,N_9551,N_9539);
nand U9668 (N_9668,N_9411,N_9507);
and U9669 (N_9669,N_9535,N_9493);
xnor U9670 (N_9670,N_9408,N_9533);
xnor U9671 (N_9671,N_9505,N_9515);
and U9672 (N_9672,N_9401,N_9421);
xor U9673 (N_9673,N_9524,N_9588);
nor U9674 (N_9674,N_9447,N_9568);
xor U9675 (N_9675,N_9584,N_9562);
nor U9676 (N_9676,N_9502,N_9464);
xor U9677 (N_9677,N_9465,N_9528);
or U9678 (N_9678,N_9504,N_9483);
nor U9679 (N_9679,N_9508,N_9458);
nor U9680 (N_9680,N_9469,N_9419);
nand U9681 (N_9681,N_9503,N_9417);
or U9682 (N_9682,N_9437,N_9428);
nor U9683 (N_9683,N_9559,N_9420);
and U9684 (N_9684,N_9510,N_9563);
nand U9685 (N_9685,N_9431,N_9499);
or U9686 (N_9686,N_9546,N_9587);
xnor U9687 (N_9687,N_9566,N_9468);
nor U9688 (N_9688,N_9402,N_9520);
or U9689 (N_9689,N_9532,N_9543);
or U9690 (N_9690,N_9496,N_9494);
and U9691 (N_9691,N_9423,N_9443);
and U9692 (N_9692,N_9558,N_9548);
nand U9693 (N_9693,N_9540,N_9580);
nor U9694 (N_9694,N_9501,N_9575);
nor U9695 (N_9695,N_9585,N_9470);
nor U9696 (N_9696,N_9480,N_9446);
or U9697 (N_9697,N_9565,N_9583);
nand U9698 (N_9698,N_9441,N_9485);
nor U9699 (N_9699,N_9586,N_9450);
nor U9700 (N_9700,N_9457,N_9492);
or U9701 (N_9701,N_9451,N_9510);
xnor U9702 (N_9702,N_9428,N_9578);
nand U9703 (N_9703,N_9595,N_9524);
and U9704 (N_9704,N_9463,N_9559);
nor U9705 (N_9705,N_9572,N_9466);
nor U9706 (N_9706,N_9531,N_9482);
and U9707 (N_9707,N_9517,N_9401);
or U9708 (N_9708,N_9445,N_9584);
and U9709 (N_9709,N_9474,N_9470);
nor U9710 (N_9710,N_9422,N_9478);
nor U9711 (N_9711,N_9550,N_9453);
xnor U9712 (N_9712,N_9547,N_9461);
xnor U9713 (N_9713,N_9428,N_9585);
nor U9714 (N_9714,N_9479,N_9516);
nand U9715 (N_9715,N_9529,N_9580);
or U9716 (N_9716,N_9433,N_9536);
nor U9717 (N_9717,N_9511,N_9568);
and U9718 (N_9718,N_9594,N_9460);
nand U9719 (N_9719,N_9502,N_9524);
nor U9720 (N_9720,N_9532,N_9555);
or U9721 (N_9721,N_9553,N_9434);
nor U9722 (N_9722,N_9573,N_9560);
and U9723 (N_9723,N_9598,N_9540);
xor U9724 (N_9724,N_9471,N_9436);
nand U9725 (N_9725,N_9452,N_9575);
or U9726 (N_9726,N_9437,N_9599);
xnor U9727 (N_9727,N_9587,N_9490);
or U9728 (N_9728,N_9424,N_9477);
and U9729 (N_9729,N_9494,N_9468);
or U9730 (N_9730,N_9475,N_9556);
or U9731 (N_9731,N_9562,N_9411);
nor U9732 (N_9732,N_9584,N_9567);
and U9733 (N_9733,N_9488,N_9545);
nand U9734 (N_9734,N_9567,N_9436);
xor U9735 (N_9735,N_9571,N_9565);
nor U9736 (N_9736,N_9409,N_9440);
and U9737 (N_9737,N_9438,N_9509);
and U9738 (N_9738,N_9450,N_9572);
nand U9739 (N_9739,N_9560,N_9455);
nor U9740 (N_9740,N_9508,N_9572);
nand U9741 (N_9741,N_9574,N_9434);
nand U9742 (N_9742,N_9489,N_9596);
nand U9743 (N_9743,N_9435,N_9586);
nor U9744 (N_9744,N_9423,N_9576);
xor U9745 (N_9745,N_9579,N_9406);
nand U9746 (N_9746,N_9559,N_9434);
and U9747 (N_9747,N_9446,N_9570);
xnor U9748 (N_9748,N_9503,N_9546);
nor U9749 (N_9749,N_9540,N_9409);
or U9750 (N_9750,N_9555,N_9591);
or U9751 (N_9751,N_9401,N_9409);
or U9752 (N_9752,N_9456,N_9516);
and U9753 (N_9753,N_9500,N_9565);
or U9754 (N_9754,N_9519,N_9506);
nor U9755 (N_9755,N_9433,N_9426);
and U9756 (N_9756,N_9470,N_9451);
and U9757 (N_9757,N_9524,N_9521);
and U9758 (N_9758,N_9437,N_9488);
xnor U9759 (N_9759,N_9469,N_9588);
or U9760 (N_9760,N_9467,N_9584);
and U9761 (N_9761,N_9454,N_9569);
or U9762 (N_9762,N_9564,N_9473);
and U9763 (N_9763,N_9573,N_9542);
nor U9764 (N_9764,N_9506,N_9515);
nand U9765 (N_9765,N_9429,N_9496);
xnor U9766 (N_9766,N_9456,N_9565);
nand U9767 (N_9767,N_9596,N_9590);
and U9768 (N_9768,N_9529,N_9483);
or U9769 (N_9769,N_9570,N_9554);
and U9770 (N_9770,N_9403,N_9457);
or U9771 (N_9771,N_9478,N_9466);
or U9772 (N_9772,N_9500,N_9508);
and U9773 (N_9773,N_9466,N_9557);
xnor U9774 (N_9774,N_9552,N_9567);
or U9775 (N_9775,N_9565,N_9498);
nor U9776 (N_9776,N_9557,N_9509);
or U9777 (N_9777,N_9428,N_9497);
xor U9778 (N_9778,N_9432,N_9425);
nor U9779 (N_9779,N_9439,N_9509);
xor U9780 (N_9780,N_9581,N_9466);
or U9781 (N_9781,N_9452,N_9500);
nor U9782 (N_9782,N_9439,N_9516);
and U9783 (N_9783,N_9587,N_9509);
or U9784 (N_9784,N_9588,N_9547);
xnor U9785 (N_9785,N_9436,N_9553);
or U9786 (N_9786,N_9561,N_9438);
xor U9787 (N_9787,N_9443,N_9515);
nor U9788 (N_9788,N_9430,N_9597);
and U9789 (N_9789,N_9476,N_9535);
nor U9790 (N_9790,N_9444,N_9503);
xor U9791 (N_9791,N_9528,N_9438);
xnor U9792 (N_9792,N_9536,N_9463);
nor U9793 (N_9793,N_9578,N_9596);
nor U9794 (N_9794,N_9531,N_9599);
nand U9795 (N_9795,N_9576,N_9570);
nor U9796 (N_9796,N_9469,N_9429);
nor U9797 (N_9797,N_9437,N_9596);
nor U9798 (N_9798,N_9567,N_9496);
or U9799 (N_9799,N_9533,N_9546);
or U9800 (N_9800,N_9681,N_9673);
and U9801 (N_9801,N_9716,N_9755);
xnor U9802 (N_9802,N_9618,N_9626);
and U9803 (N_9803,N_9744,N_9692);
or U9804 (N_9804,N_9739,N_9699);
nor U9805 (N_9805,N_9713,N_9728);
nand U9806 (N_9806,N_9703,N_9748);
and U9807 (N_9807,N_9746,N_9658);
and U9808 (N_9808,N_9687,N_9765);
nor U9809 (N_9809,N_9677,N_9791);
nor U9810 (N_9810,N_9619,N_9641);
or U9811 (N_9811,N_9645,N_9731);
nor U9812 (N_9812,N_9711,N_9768);
nand U9813 (N_9813,N_9644,N_9732);
xor U9814 (N_9814,N_9643,N_9693);
or U9815 (N_9815,N_9774,N_9617);
xnor U9816 (N_9816,N_9763,N_9624);
nand U9817 (N_9817,N_9614,N_9648);
and U9818 (N_9818,N_9789,N_9625);
and U9819 (N_9819,N_9621,N_9636);
xor U9820 (N_9820,N_9653,N_9610);
or U9821 (N_9821,N_9717,N_9706);
xor U9822 (N_9822,N_9678,N_9766);
and U9823 (N_9823,N_9737,N_9776);
nor U9824 (N_9824,N_9724,N_9627);
or U9825 (N_9825,N_9657,N_9727);
nand U9826 (N_9826,N_9694,N_9609);
nand U9827 (N_9827,N_9730,N_9661);
xnor U9828 (N_9828,N_9785,N_9634);
nor U9829 (N_9829,N_9775,N_9611);
nand U9830 (N_9830,N_9721,N_9684);
nor U9831 (N_9831,N_9719,N_9762);
nand U9832 (N_9832,N_9720,N_9722);
and U9833 (N_9833,N_9675,N_9697);
nand U9834 (N_9834,N_9790,N_9650);
xor U9835 (N_9835,N_9740,N_9689);
and U9836 (N_9836,N_9602,N_9769);
xor U9837 (N_9837,N_9799,N_9639);
xor U9838 (N_9838,N_9665,N_9761);
and U9839 (N_9839,N_9705,N_9660);
or U9840 (N_9840,N_9671,N_9793);
nand U9841 (N_9841,N_9628,N_9736);
nor U9842 (N_9842,N_9726,N_9795);
or U9843 (N_9843,N_9608,N_9751);
or U9844 (N_9844,N_9707,N_9710);
nand U9845 (N_9845,N_9637,N_9778);
and U9846 (N_9846,N_9758,N_9753);
and U9847 (N_9847,N_9756,N_9620);
nor U9848 (N_9848,N_9612,N_9742);
xor U9849 (N_9849,N_9784,N_9714);
nor U9850 (N_9850,N_9672,N_9649);
or U9851 (N_9851,N_9603,N_9704);
xor U9852 (N_9852,N_9787,N_9767);
nand U9853 (N_9853,N_9600,N_9601);
and U9854 (N_9854,N_9683,N_9680);
and U9855 (N_9855,N_9685,N_9696);
or U9856 (N_9856,N_9663,N_9733);
or U9857 (N_9857,N_9741,N_9632);
xor U9858 (N_9858,N_9715,N_9613);
or U9859 (N_9859,N_9779,N_9629);
and U9860 (N_9860,N_9666,N_9651);
nand U9861 (N_9861,N_9615,N_9690);
nand U9862 (N_9862,N_9670,N_9788);
nand U9863 (N_9863,N_9664,N_9780);
or U9864 (N_9864,N_9735,N_9708);
nor U9865 (N_9865,N_9630,N_9638);
xnor U9866 (N_9866,N_9764,N_9676);
nor U9867 (N_9867,N_9798,N_9674);
or U9868 (N_9868,N_9659,N_9796);
nand U9869 (N_9869,N_9723,N_9605);
xnor U9870 (N_9870,N_9747,N_9702);
or U9871 (N_9871,N_9667,N_9750);
and U9872 (N_9872,N_9752,N_9772);
or U9873 (N_9873,N_9698,N_9682);
nor U9874 (N_9874,N_9771,N_9631);
and U9875 (N_9875,N_9729,N_9782);
xnor U9876 (N_9876,N_9781,N_9718);
and U9877 (N_9877,N_9760,N_9633);
xnor U9878 (N_9878,N_9646,N_9607);
or U9879 (N_9879,N_9734,N_9712);
nor U9880 (N_9880,N_9773,N_9695);
nor U9881 (N_9881,N_9642,N_9662);
nand U9882 (N_9882,N_9616,N_9759);
nand U9883 (N_9883,N_9743,N_9691);
xor U9884 (N_9884,N_9623,N_9777);
nand U9885 (N_9885,N_9688,N_9754);
or U9886 (N_9886,N_9725,N_9668);
xnor U9887 (N_9887,N_9792,N_9738);
xor U9888 (N_9888,N_9606,N_9647);
nor U9889 (N_9889,N_9770,N_9686);
or U9890 (N_9890,N_9749,N_9786);
nor U9891 (N_9891,N_9797,N_9757);
or U9892 (N_9892,N_9709,N_9652);
nand U9893 (N_9893,N_9700,N_9679);
and U9894 (N_9894,N_9654,N_9783);
and U9895 (N_9895,N_9794,N_9745);
and U9896 (N_9896,N_9656,N_9640);
or U9897 (N_9897,N_9622,N_9701);
nor U9898 (N_9898,N_9635,N_9655);
and U9899 (N_9899,N_9604,N_9669);
and U9900 (N_9900,N_9713,N_9672);
nor U9901 (N_9901,N_9634,N_9767);
xor U9902 (N_9902,N_9732,N_9755);
and U9903 (N_9903,N_9741,N_9767);
and U9904 (N_9904,N_9775,N_9699);
and U9905 (N_9905,N_9761,N_9688);
nand U9906 (N_9906,N_9607,N_9790);
and U9907 (N_9907,N_9687,N_9674);
or U9908 (N_9908,N_9764,N_9724);
nor U9909 (N_9909,N_9752,N_9737);
or U9910 (N_9910,N_9666,N_9768);
and U9911 (N_9911,N_9736,N_9658);
xor U9912 (N_9912,N_9708,N_9749);
or U9913 (N_9913,N_9639,N_9760);
nand U9914 (N_9914,N_9744,N_9642);
and U9915 (N_9915,N_9707,N_9708);
and U9916 (N_9916,N_9615,N_9762);
nand U9917 (N_9917,N_9712,N_9628);
nor U9918 (N_9918,N_9667,N_9725);
xnor U9919 (N_9919,N_9698,N_9636);
nand U9920 (N_9920,N_9628,N_9730);
or U9921 (N_9921,N_9616,N_9727);
or U9922 (N_9922,N_9753,N_9672);
nor U9923 (N_9923,N_9665,N_9601);
nand U9924 (N_9924,N_9797,N_9633);
or U9925 (N_9925,N_9782,N_9665);
xnor U9926 (N_9926,N_9754,N_9736);
and U9927 (N_9927,N_9688,N_9687);
nor U9928 (N_9928,N_9658,N_9735);
xor U9929 (N_9929,N_9656,N_9671);
or U9930 (N_9930,N_9641,N_9683);
and U9931 (N_9931,N_9777,N_9722);
nand U9932 (N_9932,N_9670,N_9638);
nor U9933 (N_9933,N_9775,N_9715);
nand U9934 (N_9934,N_9746,N_9702);
nor U9935 (N_9935,N_9624,N_9670);
and U9936 (N_9936,N_9795,N_9711);
nand U9937 (N_9937,N_9684,N_9776);
nor U9938 (N_9938,N_9714,N_9628);
nor U9939 (N_9939,N_9613,N_9768);
and U9940 (N_9940,N_9610,N_9797);
xor U9941 (N_9941,N_9685,N_9699);
or U9942 (N_9942,N_9784,N_9728);
and U9943 (N_9943,N_9703,N_9674);
nor U9944 (N_9944,N_9758,N_9676);
and U9945 (N_9945,N_9775,N_9671);
nor U9946 (N_9946,N_9658,N_9708);
xor U9947 (N_9947,N_9634,N_9775);
and U9948 (N_9948,N_9619,N_9693);
or U9949 (N_9949,N_9610,N_9729);
nor U9950 (N_9950,N_9675,N_9733);
and U9951 (N_9951,N_9680,N_9632);
nor U9952 (N_9952,N_9679,N_9670);
xor U9953 (N_9953,N_9743,N_9686);
nand U9954 (N_9954,N_9618,N_9782);
and U9955 (N_9955,N_9772,N_9625);
or U9956 (N_9956,N_9766,N_9620);
and U9957 (N_9957,N_9685,N_9619);
xnor U9958 (N_9958,N_9625,N_9649);
nor U9959 (N_9959,N_9677,N_9609);
nand U9960 (N_9960,N_9756,N_9649);
and U9961 (N_9961,N_9780,N_9792);
nand U9962 (N_9962,N_9749,N_9742);
or U9963 (N_9963,N_9610,N_9718);
nor U9964 (N_9964,N_9686,N_9772);
and U9965 (N_9965,N_9680,N_9738);
xnor U9966 (N_9966,N_9655,N_9719);
nand U9967 (N_9967,N_9677,N_9632);
nand U9968 (N_9968,N_9787,N_9796);
or U9969 (N_9969,N_9722,N_9727);
and U9970 (N_9970,N_9738,N_9605);
nand U9971 (N_9971,N_9678,N_9771);
nand U9972 (N_9972,N_9791,N_9712);
xnor U9973 (N_9973,N_9748,N_9635);
nor U9974 (N_9974,N_9733,N_9680);
nor U9975 (N_9975,N_9645,N_9663);
nor U9976 (N_9976,N_9739,N_9660);
nand U9977 (N_9977,N_9605,N_9781);
or U9978 (N_9978,N_9799,N_9635);
or U9979 (N_9979,N_9716,N_9763);
or U9980 (N_9980,N_9732,N_9719);
or U9981 (N_9981,N_9658,N_9765);
and U9982 (N_9982,N_9782,N_9773);
nor U9983 (N_9983,N_9734,N_9773);
and U9984 (N_9984,N_9675,N_9777);
nand U9985 (N_9985,N_9643,N_9771);
or U9986 (N_9986,N_9763,N_9682);
or U9987 (N_9987,N_9626,N_9681);
and U9988 (N_9988,N_9748,N_9618);
and U9989 (N_9989,N_9723,N_9774);
nand U9990 (N_9990,N_9759,N_9668);
or U9991 (N_9991,N_9775,N_9761);
or U9992 (N_9992,N_9683,N_9698);
nand U9993 (N_9993,N_9700,N_9705);
or U9994 (N_9994,N_9785,N_9751);
and U9995 (N_9995,N_9700,N_9746);
or U9996 (N_9996,N_9633,N_9623);
or U9997 (N_9997,N_9703,N_9659);
and U9998 (N_9998,N_9601,N_9607);
nor U9999 (N_9999,N_9650,N_9672);
nand U10000 (N_10000,N_9878,N_9931);
nand U10001 (N_10001,N_9943,N_9914);
nor U10002 (N_10002,N_9990,N_9872);
xnor U10003 (N_10003,N_9918,N_9857);
xnor U10004 (N_10004,N_9836,N_9939);
xnor U10005 (N_10005,N_9913,N_9838);
and U10006 (N_10006,N_9861,N_9889);
or U10007 (N_10007,N_9858,N_9806);
and U10008 (N_10008,N_9803,N_9811);
nor U10009 (N_10009,N_9810,N_9978);
nand U10010 (N_10010,N_9804,N_9988);
and U10011 (N_10011,N_9897,N_9971);
or U10012 (N_10012,N_9921,N_9922);
nand U10013 (N_10013,N_9963,N_9905);
nand U10014 (N_10014,N_9821,N_9852);
or U10015 (N_10015,N_9969,N_9959);
nor U10016 (N_10016,N_9917,N_9866);
nand U10017 (N_10017,N_9805,N_9983);
nor U10018 (N_10018,N_9892,N_9887);
xnor U10019 (N_10019,N_9832,N_9946);
nor U10020 (N_10020,N_9894,N_9885);
nor U10021 (N_10021,N_9947,N_9835);
nor U10022 (N_10022,N_9809,N_9989);
and U10023 (N_10023,N_9953,N_9871);
xor U10024 (N_10024,N_9860,N_9833);
and U10025 (N_10025,N_9954,N_9879);
or U10026 (N_10026,N_9945,N_9813);
and U10027 (N_10027,N_9816,N_9968);
xor U10028 (N_10028,N_9856,N_9976);
nand U10029 (N_10029,N_9823,N_9937);
and U10030 (N_10030,N_9962,N_9824);
nand U10031 (N_10031,N_9848,N_9987);
xor U10032 (N_10032,N_9958,N_9847);
nand U10033 (N_10033,N_9808,N_9955);
and U10034 (N_10034,N_9851,N_9825);
nor U10035 (N_10035,N_9967,N_9814);
or U10036 (N_10036,N_9891,N_9901);
and U10037 (N_10037,N_9993,N_9843);
xor U10038 (N_10038,N_9915,N_9839);
nand U10039 (N_10039,N_9850,N_9819);
nor U10040 (N_10040,N_9882,N_9842);
and U10041 (N_10041,N_9920,N_9979);
xnor U10042 (N_10042,N_9909,N_9986);
and U10043 (N_10043,N_9883,N_9916);
or U10044 (N_10044,N_9985,N_9898);
and U10045 (N_10045,N_9815,N_9965);
nand U10046 (N_10046,N_9975,N_9957);
nor U10047 (N_10047,N_9876,N_9938);
or U10048 (N_10048,N_9831,N_9977);
nor U10049 (N_10049,N_9994,N_9849);
or U10050 (N_10050,N_9929,N_9801);
and U10051 (N_10051,N_9927,N_9999);
nor U10052 (N_10052,N_9951,N_9972);
nor U10053 (N_10053,N_9822,N_9865);
nand U10054 (N_10054,N_9826,N_9888);
or U10055 (N_10055,N_9868,N_9830);
nand U10056 (N_10056,N_9991,N_9974);
or U10057 (N_10057,N_9854,N_9899);
xor U10058 (N_10058,N_9829,N_9893);
nor U10059 (N_10059,N_9934,N_9944);
and U10060 (N_10060,N_9924,N_9923);
nand U10061 (N_10061,N_9911,N_9880);
and U10062 (N_10062,N_9853,N_9904);
nor U10063 (N_10063,N_9964,N_9981);
nor U10064 (N_10064,N_9807,N_9817);
nor U10065 (N_10065,N_9828,N_9942);
xnor U10066 (N_10066,N_9925,N_9940);
nand U10067 (N_10067,N_9903,N_9956);
and U10068 (N_10068,N_9966,N_9812);
xor U10069 (N_10069,N_9970,N_9802);
nor U10070 (N_10070,N_9919,N_9926);
or U10071 (N_10071,N_9930,N_9961);
nand U10072 (N_10072,N_9960,N_9906);
nand U10073 (N_10073,N_9855,N_9874);
nor U10074 (N_10074,N_9984,N_9834);
xor U10075 (N_10075,N_9928,N_9840);
or U10076 (N_10076,N_9935,N_9932);
and U10077 (N_10077,N_9973,N_9863);
nand U10078 (N_10078,N_9859,N_9941);
or U10079 (N_10079,N_9950,N_9948);
nor U10080 (N_10080,N_9936,N_9837);
and U10081 (N_10081,N_9867,N_9869);
xnor U10082 (N_10082,N_9846,N_9884);
nand U10083 (N_10083,N_9895,N_9907);
nand U10084 (N_10084,N_9877,N_9881);
nand U10085 (N_10085,N_9827,N_9864);
and U10086 (N_10086,N_9982,N_9873);
nor U10087 (N_10087,N_9818,N_9841);
nor U10088 (N_10088,N_9902,N_9912);
or U10089 (N_10089,N_9949,N_9870);
xnor U10090 (N_10090,N_9910,N_9890);
and U10091 (N_10091,N_9900,N_9862);
nor U10092 (N_10092,N_9933,N_9992);
nand U10093 (N_10093,N_9998,N_9896);
and U10094 (N_10094,N_9997,N_9844);
or U10095 (N_10095,N_9995,N_9908);
or U10096 (N_10096,N_9875,N_9952);
or U10097 (N_10097,N_9845,N_9800);
xor U10098 (N_10098,N_9820,N_9996);
or U10099 (N_10099,N_9886,N_9980);
nand U10100 (N_10100,N_9872,N_9876);
nand U10101 (N_10101,N_9863,N_9946);
and U10102 (N_10102,N_9826,N_9993);
nand U10103 (N_10103,N_9899,N_9855);
and U10104 (N_10104,N_9991,N_9948);
nand U10105 (N_10105,N_9805,N_9841);
and U10106 (N_10106,N_9966,N_9909);
nor U10107 (N_10107,N_9926,N_9823);
nor U10108 (N_10108,N_9885,N_9893);
nand U10109 (N_10109,N_9987,N_9890);
nor U10110 (N_10110,N_9803,N_9856);
xor U10111 (N_10111,N_9936,N_9908);
and U10112 (N_10112,N_9901,N_9976);
and U10113 (N_10113,N_9866,N_9994);
nor U10114 (N_10114,N_9813,N_9948);
and U10115 (N_10115,N_9968,N_9850);
or U10116 (N_10116,N_9832,N_9839);
nor U10117 (N_10117,N_9889,N_9970);
nor U10118 (N_10118,N_9930,N_9800);
xnor U10119 (N_10119,N_9818,N_9930);
nand U10120 (N_10120,N_9878,N_9991);
nand U10121 (N_10121,N_9934,N_9967);
xnor U10122 (N_10122,N_9929,N_9874);
nand U10123 (N_10123,N_9947,N_9824);
nor U10124 (N_10124,N_9945,N_9906);
nand U10125 (N_10125,N_9825,N_9893);
or U10126 (N_10126,N_9963,N_9851);
nor U10127 (N_10127,N_9946,N_9973);
nand U10128 (N_10128,N_9861,N_9800);
nand U10129 (N_10129,N_9839,N_9852);
and U10130 (N_10130,N_9830,N_9990);
nand U10131 (N_10131,N_9967,N_9838);
nor U10132 (N_10132,N_9907,N_9939);
xor U10133 (N_10133,N_9833,N_9845);
nand U10134 (N_10134,N_9913,N_9890);
nor U10135 (N_10135,N_9958,N_9886);
and U10136 (N_10136,N_9885,N_9837);
nor U10137 (N_10137,N_9914,N_9987);
nand U10138 (N_10138,N_9977,N_9835);
nand U10139 (N_10139,N_9952,N_9953);
xnor U10140 (N_10140,N_9871,N_9907);
nor U10141 (N_10141,N_9907,N_9906);
xor U10142 (N_10142,N_9980,N_9978);
nor U10143 (N_10143,N_9831,N_9903);
and U10144 (N_10144,N_9852,N_9861);
nor U10145 (N_10145,N_9972,N_9999);
and U10146 (N_10146,N_9949,N_9974);
and U10147 (N_10147,N_9995,N_9973);
nor U10148 (N_10148,N_9831,N_9835);
nand U10149 (N_10149,N_9977,N_9974);
xnor U10150 (N_10150,N_9816,N_9966);
nand U10151 (N_10151,N_9950,N_9954);
nor U10152 (N_10152,N_9986,N_9876);
nand U10153 (N_10153,N_9874,N_9935);
nor U10154 (N_10154,N_9804,N_9952);
nand U10155 (N_10155,N_9878,N_9915);
nor U10156 (N_10156,N_9897,N_9998);
nor U10157 (N_10157,N_9940,N_9822);
or U10158 (N_10158,N_9856,N_9937);
nor U10159 (N_10159,N_9892,N_9873);
xnor U10160 (N_10160,N_9823,N_9836);
and U10161 (N_10161,N_9948,N_9972);
nand U10162 (N_10162,N_9874,N_9905);
and U10163 (N_10163,N_9879,N_9882);
xnor U10164 (N_10164,N_9836,N_9978);
or U10165 (N_10165,N_9872,N_9989);
and U10166 (N_10166,N_9897,N_9992);
or U10167 (N_10167,N_9961,N_9896);
nor U10168 (N_10168,N_9847,N_9888);
or U10169 (N_10169,N_9863,N_9993);
and U10170 (N_10170,N_9818,N_9872);
xor U10171 (N_10171,N_9831,N_9978);
and U10172 (N_10172,N_9911,N_9973);
or U10173 (N_10173,N_9990,N_9910);
xnor U10174 (N_10174,N_9889,N_9939);
and U10175 (N_10175,N_9875,N_9877);
and U10176 (N_10176,N_9964,N_9944);
and U10177 (N_10177,N_9942,N_9937);
and U10178 (N_10178,N_9811,N_9938);
nand U10179 (N_10179,N_9946,N_9966);
xnor U10180 (N_10180,N_9864,N_9939);
nor U10181 (N_10181,N_9848,N_9982);
xor U10182 (N_10182,N_9989,N_9953);
and U10183 (N_10183,N_9932,N_9996);
xnor U10184 (N_10184,N_9939,N_9931);
nor U10185 (N_10185,N_9907,N_9822);
xnor U10186 (N_10186,N_9921,N_9975);
xor U10187 (N_10187,N_9956,N_9908);
nand U10188 (N_10188,N_9801,N_9872);
nand U10189 (N_10189,N_9862,N_9864);
nor U10190 (N_10190,N_9961,N_9911);
nand U10191 (N_10191,N_9956,N_9829);
nor U10192 (N_10192,N_9815,N_9975);
xnor U10193 (N_10193,N_9960,N_9866);
and U10194 (N_10194,N_9816,N_9977);
and U10195 (N_10195,N_9975,N_9983);
nand U10196 (N_10196,N_9921,N_9898);
and U10197 (N_10197,N_9812,N_9983);
nor U10198 (N_10198,N_9979,N_9923);
xnor U10199 (N_10199,N_9842,N_9952);
or U10200 (N_10200,N_10005,N_10139);
xor U10201 (N_10201,N_10001,N_10138);
or U10202 (N_10202,N_10037,N_10034);
and U10203 (N_10203,N_10130,N_10192);
nor U10204 (N_10204,N_10155,N_10093);
nor U10205 (N_10205,N_10025,N_10014);
nor U10206 (N_10206,N_10178,N_10193);
or U10207 (N_10207,N_10082,N_10111);
and U10208 (N_10208,N_10194,N_10048);
nand U10209 (N_10209,N_10117,N_10099);
and U10210 (N_10210,N_10079,N_10113);
xor U10211 (N_10211,N_10181,N_10183);
xnor U10212 (N_10212,N_10032,N_10105);
xnor U10213 (N_10213,N_10051,N_10120);
or U10214 (N_10214,N_10008,N_10011);
or U10215 (N_10215,N_10028,N_10062);
nand U10216 (N_10216,N_10163,N_10075);
or U10217 (N_10217,N_10076,N_10080);
nand U10218 (N_10218,N_10009,N_10021);
nand U10219 (N_10219,N_10161,N_10086);
and U10220 (N_10220,N_10114,N_10043);
xnor U10221 (N_10221,N_10084,N_10019);
nor U10222 (N_10222,N_10189,N_10151);
or U10223 (N_10223,N_10018,N_10053);
nand U10224 (N_10224,N_10169,N_10085);
xnor U10225 (N_10225,N_10179,N_10195);
or U10226 (N_10226,N_10087,N_10174);
and U10227 (N_10227,N_10003,N_10126);
nor U10228 (N_10228,N_10102,N_10110);
or U10229 (N_10229,N_10175,N_10128);
and U10230 (N_10230,N_10020,N_10007);
nand U10231 (N_10231,N_10198,N_10153);
nand U10232 (N_10232,N_10177,N_10088);
nand U10233 (N_10233,N_10013,N_10044);
nand U10234 (N_10234,N_10004,N_10171);
nand U10235 (N_10235,N_10060,N_10184);
xor U10236 (N_10236,N_10131,N_10083);
or U10237 (N_10237,N_10038,N_10058);
xor U10238 (N_10238,N_10107,N_10096);
nand U10239 (N_10239,N_10190,N_10010);
and U10240 (N_10240,N_10137,N_10045);
and U10241 (N_10241,N_10109,N_10006);
nand U10242 (N_10242,N_10050,N_10112);
nor U10243 (N_10243,N_10168,N_10191);
xnor U10244 (N_10244,N_10148,N_10152);
nand U10245 (N_10245,N_10091,N_10154);
nor U10246 (N_10246,N_10156,N_10090);
nand U10247 (N_10247,N_10027,N_10125);
or U10248 (N_10248,N_10182,N_10035);
xor U10249 (N_10249,N_10170,N_10040);
xnor U10250 (N_10250,N_10165,N_10104);
xor U10251 (N_10251,N_10015,N_10002);
or U10252 (N_10252,N_10095,N_10036);
and U10253 (N_10253,N_10049,N_10135);
and U10254 (N_10254,N_10068,N_10103);
xor U10255 (N_10255,N_10078,N_10101);
nand U10256 (N_10256,N_10158,N_10066);
and U10257 (N_10257,N_10022,N_10063);
or U10258 (N_10258,N_10186,N_10041);
or U10259 (N_10259,N_10072,N_10132);
or U10260 (N_10260,N_10061,N_10012);
nor U10261 (N_10261,N_10150,N_10094);
xnor U10262 (N_10262,N_10000,N_10092);
nor U10263 (N_10263,N_10054,N_10077);
nor U10264 (N_10264,N_10100,N_10167);
or U10265 (N_10265,N_10134,N_10081);
xor U10266 (N_10266,N_10119,N_10056);
and U10267 (N_10267,N_10157,N_10147);
xor U10268 (N_10268,N_10065,N_10121);
nor U10269 (N_10269,N_10122,N_10055);
or U10270 (N_10270,N_10159,N_10059);
xnor U10271 (N_10271,N_10173,N_10162);
nor U10272 (N_10272,N_10047,N_10188);
or U10273 (N_10273,N_10039,N_10097);
nor U10274 (N_10274,N_10067,N_10064);
xnor U10275 (N_10275,N_10146,N_10166);
nor U10276 (N_10276,N_10098,N_10071);
or U10277 (N_10277,N_10106,N_10164);
nor U10278 (N_10278,N_10026,N_10115);
xnor U10279 (N_10279,N_10160,N_10042);
or U10280 (N_10280,N_10017,N_10185);
nand U10281 (N_10281,N_10172,N_10016);
xnor U10282 (N_10282,N_10127,N_10136);
nand U10283 (N_10283,N_10145,N_10129);
xnor U10284 (N_10284,N_10057,N_10141);
xnor U10285 (N_10285,N_10031,N_10142);
and U10286 (N_10286,N_10133,N_10180);
nand U10287 (N_10287,N_10187,N_10108);
nor U10288 (N_10288,N_10089,N_10046);
xnor U10289 (N_10289,N_10149,N_10176);
xnor U10290 (N_10290,N_10196,N_10143);
and U10291 (N_10291,N_10030,N_10070);
nor U10292 (N_10292,N_10052,N_10073);
xnor U10293 (N_10293,N_10033,N_10118);
and U10294 (N_10294,N_10197,N_10074);
nor U10295 (N_10295,N_10024,N_10029);
and U10296 (N_10296,N_10123,N_10199);
nor U10297 (N_10297,N_10023,N_10069);
nand U10298 (N_10298,N_10140,N_10144);
nand U10299 (N_10299,N_10116,N_10124);
nand U10300 (N_10300,N_10178,N_10087);
nand U10301 (N_10301,N_10142,N_10109);
nor U10302 (N_10302,N_10053,N_10113);
nor U10303 (N_10303,N_10005,N_10079);
nand U10304 (N_10304,N_10161,N_10106);
nor U10305 (N_10305,N_10059,N_10173);
nor U10306 (N_10306,N_10170,N_10050);
nand U10307 (N_10307,N_10072,N_10180);
xor U10308 (N_10308,N_10058,N_10127);
xnor U10309 (N_10309,N_10099,N_10186);
nor U10310 (N_10310,N_10018,N_10106);
or U10311 (N_10311,N_10184,N_10143);
xor U10312 (N_10312,N_10000,N_10026);
or U10313 (N_10313,N_10180,N_10027);
or U10314 (N_10314,N_10167,N_10030);
nand U10315 (N_10315,N_10132,N_10079);
nand U10316 (N_10316,N_10036,N_10023);
nor U10317 (N_10317,N_10118,N_10178);
and U10318 (N_10318,N_10157,N_10141);
nand U10319 (N_10319,N_10083,N_10090);
and U10320 (N_10320,N_10092,N_10101);
and U10321 (N_10321,N_10170,N_10036);
or U10322 (N_10322,N_10007,N_10069);
or U10323 (N_10323,N_10053,N_10058);
or U10324 (N_10324,N_10012,N_10118);
or U10325 (N_10325,N_10142,N_10175);
nor U10326 (N_10326,N_10002,N_10037);
xor U10327 (N_10327,N_10166,N_10037);
xnor U10328 (N_10328,N_10152,N_10142);
or U10329 (N_10329,N_10060,N_10168);
nor U10330 (N_10330,N_10147,N_10161);
nand U10331 (N_10331,N_10008,N_10068);
nor U10332 (N_10332,N_10087,N_10015);
xnor U10333 (N_10333,N_10068,N_10085);
nand U10334 (N_10334,N_10134,N_10024);
nand U10335 (N_10335,N_10008,N_10062);
nand U10336 (N_10336,N_10134,N_10165);
xnor U10337 (N_10337,N_10023,N_10180);
xnor U10338 (N_10338,N_10101,N_10123);
nand U10339 (N_10339,N_10035,N_10177);
nor U10340 (N_10340,N_10030,N_10007);
nor U10341 (N_10341,N_10083,N_10080);
xnor U10342 (N_10342,N_10040,N_10029);
nor U10343 (N_10343,N_10027,N_10028);
nand U10344 (N_10344,N_10081,N_10011);
nand U10345 (N_10345,N_10143,N_10080);
nor U10346 (N_10346,N_10169,N_10097);
nor U10347 (N_10347,N_10068,N_10088);
and U10348 (N_10348,N_10174,N_10015);
xor U10349 (N_10349,N_10025,N_10069);
and U10350 (N_10350,N_10040,N_10146);
nand U10351 (N_10351,N_10185,N_10011);
nand U10352 (N_10352,N_10075,N_10171);
or U10353 (N_10353,N_10167,N_10051);
xor U10354 (N_10354,N_10002,N_10008);
and U10355 (N_10355,N_10072,N_10149);
nand U10356 (N_10356,N_10032,N_10183);
xor U10357 (N_10357,N_10061,N_10018);
xnor U10358 (N_10358,N_10128,N_10157);
and U10359 (N_10359,N_10044,N_10011);
xor U10360 (N_10360,N_10185,N_10121);
and U10361 (N_10361,N_10006,N_10070);
nand U10362 (N_10362,N_10179,N_10153);
nor U10363 (N_10363,N_10087,N_10026);
or U10364 (N_10364,N_10039,N_10009);
and U10365 (N_10365,N_10187,N_10011);
and U10366 (N_10366,N_10124,N_10189);
and U10367 (N_10367,N_10052,N_10123);
and U10368 (N_10368,N_10165,N_10057);
nor U10369 (N_10369,N_10019,N_10025);
nor U10370 (N_10370,N_10043,N_10004);
nand U10371 (N_10371,N_10073,N_10045);
and U10372 (N_10372,N_10001,N_10049);
nor U10373 (N_10373,N_10041,N_10111);
and U10374 (N_10374,N_10109,N_10154);
nor U10375 (N_10375,N_10083,N_10165);
xor U10376 (N_10376,N_10161,N_10083);
or U10377 (N_10377,N_10129,N_10012);
and U10378 (N_10378,N_10136,N_10037);
nor U10379 (N_10379,N_10198,N_10178);
and U10380 (N_10380,N_10122,N_10024);
and U10381 (N_10381,N_10141,N_10154);
nor U10382 (N_10382,N_10170,N_10144);
nor U10383 (N_10383,N_10102,N_10086);
nand U10384 (N_10384,N_10004,N_10035);
nand U10385 (N_10385,N_10009,N_10112);
or U10386 (N_10386,N_10149,N_10157);
or U10387 (N_10387,N_10050,N_10000);
nor U10388 (N_10388,N_10152,N_10129);
nor U10389 (N_10389,N_10053,N_10174);
nor U10390 (N_10390,N_10144,N_10129);
nand U10391 (N_10391,N_10105,N_10138);
nand U10392 (N_10392,N_10050,N_10033);
xnor U10393 (N_10393,N_10025,N_10149);
nor U10394 (N_10394,N_10116,N_10123);
xnor U10395 (N_10395,N_10137,N_10197);
nor U10396 (N_10396,N_10018,N_10014);
or U10397 (N_10397,N_10174,N_10048);
and U10398 (N_10398,N_10061,N_10088);
nand U10399 (N_10399,N_10157,N_10187);
or U10400 (N_10400,N_10264,N_10241);
or U10401 (N_10401,N_10268,N_10360);
nand U10402 (N_10402,N_10259,N_10387);
or U10403 (N_10403,N_10321,N_10316);
xor U10404 (N_10404,N_10248,N_10256);
nand U10405 (N_10405,N_10263,N_10266);
nand U10406 (N_10406,N_10227,N_10231);
xor U10407 (N_10407,N_10285,N_10297);
and U10408 (N_10408,N_10385,N_10291);
nor U10409 (N_10409,N_10375,N_10280);
and U10410 (N_10410,N_10324,N_10255);
or U10411 (N_10411,N_10254,N_10382);
or U10412 (N_10412,N_10222,N_10223);
xnor U10413 (N_10413,N_10214,N_10358);
or U10414 (N_10414,N_10395,N_10299);
or U10415 (N_10415,N_10328,N_10335);
and U10416 (N_10416,N_10312,N_10247);
and U10417 (N_10417,N_10219,N_10287);
and U10418 (N_10418,N_10230,N_10202);
nand U10419 (N_10419,N_10218,N_10304);
xnor U10420 (N_10420,N_10277,N_10210);
nand U10421 (N_10421,N_10365,N_10322);
or U10422 (N_10422,N_10346,N_10340);
and U10423 (N_10423,N_10323,N_10331);
xnor U10424 (N_10424,N_10349,N_10279);
and U10425 (N_10425,N_10267,N_10374);
xor U10426 (N_10426,N_10251,N_10298);
nand U10427 (N_10427,N_10302,N_10221);
nand U10428 (N_10428,N_10327,N_10276);
nor U10429 (N_10429,N_10239,N_10284);
nand U10430 (N_10430,N_10208,N_10288);
or U10431 (N_10431,N_10369,N_10399);
or U10432 (N_10432,N_10319,N_10381);
nand U10433 (N_10433,N_10228,N_10206);
nand U10434 (N_10434,N_10253,N_10378);
nor U10435 (N_10435,N_10326,N_10308);
nand U10436 (N_10436,N_10330,N_10238);
xnor U10437 (N_10437,N_10334,N_10359);
xnor U10438 (N_10438,N_10215,N_10213);
nor U10439 (N_10439,N_10220,N_10361);
nand U10440 (N_10440,N_10234,N_10217);
nand U10441 (N_10441,N_10292,N_10366);
or U10442 (N_10442,N_10394,N_10211);
and U10443 (N_10443,N_10337,N_10318);
nand U10444 (N_10444,N_10362,N_10354);
nand U10445 (N_10445,N_10351,N_10353);
nand U10446 (N_10446,N_10301,N_10283);
xnor U10447 (N_10447,N_10286,N_10314);
xor U10448 (N_10448,N_10204,N_10348);
xor U10449 (N_10449,N_10244,N_10329);
nor U10450 (N_10450,N_10376,N_10236);
nand U10451 (N_10451,N_10303,N_10282);
nor U10452 (N_10452,N_10216,N_10293);
and U10453 (N_10453,N_10281,N_10245);
and U10454 (N_10454,N_10391,N_10235);
or U10455 (N_10455,N_10300,N_10257);
xnor U10456 (N_10456,N_10270,N_10367);
nor U10457 (N_10457,N_10273,N_10243);
or U10458 (N_10458,N_10242,N_10379);
and U10459 (N_10459,N_10290,N_10311);
nand U10460 (N_10460,N_10246,N_10389);
or U10461 (N_10461,N_10224,N_10237);
and U10462 (N_10462,N_10294,N_10262);
xnor U10463 (N_10463,N_10345,N_10357);
xnor U10464 (N_10464,N_10317,N_10332);
nand U10465 (N_10465,N_10258,N_10372);
or U10466 (N_10466,N_10229,N_10364);
nand U10467 (N_10467,N_10265,N_10203);
xor U10468 (N_10468,N_10380,N_10212);
or U10469 (N_10469,N_10201,N_10252);
nor U10470 (N_10470,N_10383,N_10232);
and U10471 (N_10471,N_10355,N_10272);
and U10472 (N_10472,N_10205,N_10356);
nand U10473 (N_10473,N_10295,N_10344);
nor U10474 (N_10474,N_10305,N_10397);
and U10475 (N_10475,N_10352,N_10342);
or U10476 (N_10476,N_10390,N_10278);
xnor U10477 (N_10477,N_10274,N_10240);
nand U10478 (N_10478,N_10275,N_10377);
or U10479 (N_10479,N_10269,N_10386);
or U10480 (N_10480,N_10370,N_10373);
or U10481 (N_10481,N_10336,N_10271);
nor U10482 (N_10482,N_10325,N_10261);
nand U10483 (N_10483,N_10398,N_10233);
nor U10484 (N_10484,N_10388,N_10384);
or U10485 (N_10485,N_10249,N_10320);
nor U10486 (N_10486,N_10371,N_10309);
or U10487 (N_10487,N_10200,N_10307);
xor U10488 (N_10488,N_10368,N_10393);
xor U10489 (N_10489,N_10296,N_10350);
nand U10490 (N_10490,N_10396,N_10260);
xor U10491 (N_10491,N_10313,N_10333);
nor U10492 (N_10492,N_10392,N_10315);
and U10493 (N_10493,N_10341,N_10310);
nor U10494 (N_10494,N_10347,N_10306);
xnor U10495 (N_10495,N_10339,N_10289);
or U10496 (N_10496,N_10226,N_10225);
nor U10497 (N_10497,N_10207,N_10209);
xnor U10498 (N_10498,N_10363,N_10343);
xnor U10499 (N_10499,N_10338,N_10250);
nor U10500 (N_10500,N_10258,N_10329);
and U10501 (N_10501,N_10329,N_10387);
xor U10502 (N_10502,N_10209,N_10202);
nand U10503 (N_10503,N_10389,N_10338);
xor U10504 (N_10504,N_10368,N_10334);
or U10505 (N_10505,N_10375,N_10376);
nor U10506 (N_10506,N_10348,N_10220);
nor U10507 (N_10507,N_10286,N_10334);
nand U10508 (N_10508,N_10318,N_10307);
and U10509 (N_10509,N_10399,N_10290);
nand U10510 (N_10510,N_10211,N_10312);
xor U10511 (N_10511,N_10391,N_10218);
nor U10512 (N_10512,N_10318,N_10355);
and U10513 (N_10513,N_10370,N_10308);
nand U10514 (N_10514,N_10376,N_10361);
or U10515 (N_10515,N_10251,N_10343);
xor U10516 (N_10516,N_10255,N_10219);
or U10517 (N_10517,N_10350,N_10249);
nand U10518 (N_10518,N_10263,N_10245);
nand U10519 (N_10519,N_10262,N_10374);
nor U10520 (N_10520,N_10369,N_10365);
xnor U10521 (N_10521,N_10384,N_10235);
xnor U10522 (N_10522,N_10374,N_10355);
or U10523 (N_10523,N_10350,N_10344);
and U10524 (N_10524,N_10294,N_10349);
xnor U10525 (N_10525,N_10317,N_10211);
xor U10526 (N_10526,N_10266,N_10356);
xnor U10527 (N_10527,N_10235,N_10360);
xor U10528 (N_10528,N_10233,N_10393);
and U10529 (N_10529,N_10388,N_10258);
xnor U10530 (N_10530,N_10311,N_10213);
and U10531 (N_10531,N_10334,N_10304);
nand U10532 (N_10532,N_10304,N_10254);
nand U10533 (N_10533,N_10265,N_10258);
or U10534 (N_10534,N_10351,N_10399);
nand U10535 (N_10535,N_10307,N_10366);
nand U10536 (N_10536,N_10274,N_10261);
nand U10537 (N_10537,N_10296,N_10330);
or U10538 (N_10538,N_10290,N_10298);
xor U10539 (N_10539,N_10231,N_10240);
nand U10540 (N_10540,N_10345,N_10363);
and U10541 (N_10541,N_10238,N_10380);
xor U10542 (N_10542,N_10251,N_10351);
and U10543 (N_10543,N_10325,N_10339);
nand U10544 (N_10544,N_10336,N_10387);
nand U10545 (N_10545,N_10312,N_10300);
nor U10546 (N_10546,N_10206,N_10317);
and U10547 (N_10547,N_10243,N_10206);
or U10548 (N_10548,N_10258,N_10207);
nand U10549 (N_10549,N_10229,N_10265);
xor U10550 (N_10550,N_10200,N_10371);
and U10551 (N_10551,N_10220,N_10203);
nand U10552 (N_10552,N_10343,N_10356);
nand U10553 (N_10553,N_10227,N_10310);
nand U10554 (N_10554,N_10292,N_10293);
nand U10555 (N_10555,N_10304,N_10282);
nand U10556 (N_10556,N_10272,N_10255);
xor U10557 (N_10557,N_10236,N_10396);
nand U10558 (N_10558,N_10296,N_10251);
nor U10559 (N_10559,N_10385,N_10240);
and U10560 (N_10560,N_10361,N_10333);
xor U10561 (N_10561,N_10321,N_10273);
nor U10562 (N_10562,N_10297,N_10395);
nand U10563 (N_10563,N_10276,N_10314);
xnor U10564 (N_10564,N_10287,N_10361);
or U10565 (N_10565,N_10351,N_10349);
nand U10566 (N_10566,N_10232,N_10247);
or U10567 (N_10567,N_10349,N_10243);
or U10568 (N_10568,N_10240,N_10202);
or U10569 (N_10569,N_10330,N_10247);
nor U10570 (N_10570,N_10371,N_10242);
or U10571 (N_10571,N_10393,N_10262);
and U10572 (N_10572,N_10256,N_10245);
or U10573 (N_10573,N_10247,N_10238);
and U10574 (N_10574,N_10303,N_10220);
and U10575 (N_10575,N_10226,N_10332);
nand U10576 (N_10576,N_10263,N_10360);
xnor U10577 (N_10577,N_10325,N_10226);
or U10578 (N_10578,N_10294,N_10322);
or U10579 (N_10579,N_10357,N_10312);
nand U10580 (N_10580,N_10349,N_10281);
and U10581 (N_10581,N_10333,N_10310);
or U10582 (N_10582,N_10226,N_10259);
xor U10583 (N_10583,N_10377,N_10214);
or U10584 (N_10584,N_10201,N_10239);
nor U10585 (N_10585,N_10362,N_10383);
xor U10586 (N_10586,N_10203,N_10262);
xor U10587 (N_10587,N_10237,N_10355);
nand U10588 (N_10588,N_10393,N_10397);
or U10589 (N_10589,N_10225,N_10286);
nand U10590 (N_10590,N_10246,N_10264);
or U10591 (N_10591,N_10286,N_10274);
nand U10592 (N_10592,N_10301,N_10243);
nand U10593 (N_10593,N_10271,N_10329);
xnor U10594 (N_10594,N_10313,N_10297);
nand U10595 (N_10595,N_10273,N_10228);
xnor U10596 (N_10596,N_10340,N_10324);
nor U10597 (N_10597,N_10317,N_10386);
nor U10598 (N_10598,N_10249,N_10279);
nand U10599 (N_10599,N_10374,N_10341);
xor U10600 (N_10600,N_10476,N_10543);
or U10601 (N_10601,N_10449,N_10445);
nand U10602 (N_10602,N_10450,N_10436);
nor U10603 (N_10603,N_10552,N_10422);
nor U10604 (N_10604,N_10410,N_10592);
xnor U10605 (N_10605,N_10475,N_10578);
and U10606 (N_10606,N_10582,N_10457);
and U10607 (N_10607,N_10570,N_10426);
and U10608 (N_10608,N_10580,N_10485);
xor U10609 (N_10609,N_10462,N_10429);
or U10610 (N_10610,N_10527,N_10589);
xor U10611 (N_10611,N_10486,N_10507);
nand U10612 (N_10612,N_10521,N_10510);
and U10613 (N_10613,N_10432,N_10553);
and U10614 (N_10614,N_10407,N_10522);
nand U10615 (N_10615,N_10406,N_10467);
nor U10616 (N_10616,N_10425,N_10549);
and U10617 (N_10617,N_10459,N_10433);
and U10618 (N_10618,N_10488,N_10538);
nor U10619 (N_10619,N_10454,N_10595);
nor U10620 (N_10620,N_10421,N_10484);
or U10621 (N_10621,N_10472,N_10474);
xor U10622 (N_10622,N_10572,N_10588);
xor U10623 (N_10623,N_10428,N_10435);
nand U10624 (N_10624,N_10573,N_10593);
nand U10625 (N_10625,N_10417,N_10400);
or U10626 (N_10626,N_10530,N_10402);
xor U10627 (N_10627,N_10496,N_10565);
nand U10628 (N_10628,N_10430,N_10556);
or U10629 (N_10629,N_10513,N_10451);
or U10630 (N_10630,N_10514,N_10498);
and U10631 (N_10631,N_10517,N_10456);
or U10632 (N_10632,N_10438,N_10569);
xor U10633 (N_10633,N_10544,N_10523);
and U10634 (N_10634,N_10585,N_10473);
and U10635 (N_10635,N_10586,N_10405);
xor U10636 (N_10636,N_10542,N_10529);
xor U10637 (N_10637,N_10443,N_10493);
and U10638 (N_10638,N_10536,N_10494);
and U10639 (N_10639,N_10453,N_10557);
xnor U10640 (N_10640,N_10520,N_10558);
or U10641 (N_10641,N_10584,N_10455);
nand U10642 (N_10642,N_10534,N_10408);
nor U10643 (N_10643,N_10574,N_10568);
nand U10644 (N_10644,N_10541,N_10576);
nand U10645 (N_10645,N_10489,N_10562);
nand U10646 (N_10646,N_10499,N_10437);
nand U10647 (N_10647,N_10590,N_10471);
or U10648 (N_10648,N_10444,N_10434);
or U10649 (N_10649,N_10504,N_10581);
nor U10650 (N_10650,N_10497,N_10579);
or U10651 (N_10651,N_10566,N_10539);
nand U10652 (N_10652,N_10412,N_10446);
nor U10653 (N_10653,N_10519,N_10452);
nor U10654 (N_10654,N_10464,N_10501);
nand U10655 (N_10655,N_10414,N_10509);
nand U10656 (N_10656,N_10526,N_10401);
and U10657 (N_10657,N_10487,N_10439);
nor U10658 (N_10658,N_10516,N_10528);
nand U10659 (N_10659,N_10481,N_10468);
or U10660 (N_10660,N_10477,N_10466);
and U10661 (N_10661,N_10492,N_10448);
xor U10662 (N_10662,N_10518,N_10535);
xor U10663 (N_10663,N_10548,N_10483);
xnor U10664 (N_10664,N_10463,N_10503);
and U10665 (N_10665,N_10480,N_10418);
xnor U10666 (N_10666,N_10469,N_10571);
and U10667 (N_10667,N_10482,N_10419);
or U10668 (N_10668,N_10490,N_10560);
and U10669 (N_10669,N_10403,N_10575);
and U10670 (N_10670,N_10596,N_10547);
nand U10671 (N_10671,N_10404,N_10413);
nor U10672 (N_10672,N_10460,N_10531);
nand U10673 (N_10673,N_10411,N_10461);
xor U10674 (N_10674,N_10440,N_10506);
nand U10675 (N_10675,N_10591,N_10416);
nand U10676 (N_10676,N_10511,N_10508);
nor U10677 (N_10677,N_10423,N_10540);
nand U10678 (N_10678,N_10525,N_10599);
nor U10679 (N_10679,N_10491,N_10597);
or U10680 (N_10680,N_10577,N_10563);
xnor U10681 (N_10681,N_10559,N_10537);
or U10682 (N_10682,N_10447,N_10587);
nand U10683 (N_10683,N_10441,N_10546);
nand U10684 (N_10684,N_10550,N_10533);
xnor U10685 (N_10685,N_10567,N_10561);
nor U10686 (N_10686,N_10409,N_10555);
or U10687 (N_10687,N_10500,N_10598);
and U10688 (N_10688,N_10427,N_10442);
nor U10689 (N_10689,N_10524,N_10583);
nand U10690 (N_10690,N_10424,N_10532);
and U10691 (N_10691,N_10431,N_10564);
nand U10692 (N_10692,N_10545,N_10465);
nand U10693 (N_10693,N_10415,N_10554);
or U10694 (N_10694,N_10458,N_10551);
nand U10695 (N_10695,N_10512,N_10470);
or U10696 (N_10696,N_10502,N_10594);
nand U10697 (N_10697,N_10420,N_10515);
and U10698 (N_10698,N_10505,N_10479);
and U10699 (N_10699,N_10495,N_10478);
nand U10700 (N_10700,N_10589,N_10447);
or U10701 (N_10701,N_10549,N_10518);
and U10702 (N_10702,N_10422,N_10556);
nand U10703 (N_10703,N_10467,N_10452);
nand U10704 (N_10704,N_10561,N_10511);
nand U10705 (N_10705,N_10534,N_10528);
or U10706 (N_10706,N_10449,N_10557);
nor U10707 (N_10707,N_10560,N_10580);
xor U10708 (N_10708,N_10450,N_10547);
xor U10709 (N_10709,N_10568,N_10539);
xor U10710 (N_10710,N_10553,N_10445);
nand U10711 (N_10711,N_10538,N_10536);
nor U10712 (N_10712,N_10470,N_10550);
or U10713 (N_10713,N_10595,N_10447);
and U10714 (N_10714,N_10576,N_10477);
or U10715 (N_10715,N_10579,N_10436);
or U10716 (N_10716,N_10410,N_10491);
xnor U10717 (N_10717,N_10554,N_10483);
xor U10718 (N_10718,N_10472,N_10574);
or U10719 (N_10719,N_10427,N_10502);
and U10720 (N_10720,N_10541,N_10418);
nand U10721 (N_10721,N_10541,N_10565);
xnor U10722 (N_10722,N_10405,N_10597);
or U10723 (N_10723,N_10593,N_10433);
xnor U10724 (N_10724,N_10416,N_10561);
nand U10725 (N_10725,N_10567,N_10572);
and U10726 (N_10726,N_10426,N_10441);
or U10727 (N_10727,N_10528,N_10583);
or U10728 (N_10728,N_10434,N_10424);
or U10729 (N_10729,N_10545,N_10469);
and U10730 (N_10730,N_10503,N_10558);
or U10731 (N_10731,N_10525,N_10532);
nor U10732 (N_10732,N_10551,N_10561);
nand U10733 (N_10733,N_10541,N_10506);
and U10734 (N_10734,N_10455,N_10486);
or U10735 (N_10735,N_10441,N_10548);
xor U10736 (N_10736,N_10504,N_10411);
nor U10737 (N_10737,N_10428,N_10409);
xor U10738 (N_10738,N_10458,N_10453);
and U10739 (N_10739,N_10445,N_10474);
nor U10740 (N_10740,N_10504,N_10593);
or U10741 (N_10741,N_10436,N_10428);
and U10742 (N_10742,N_10422,N_10573);
and U10743 (N_10743,N_10420,N_10563);
and U10744 (N_10744,N_10487,N_10596);
or U10745 (N_10745,N_10521,N_10591);
nand U10746 (N_10746,N_10548,N_10574);
and U10747 (N_10747,N_10504,N_10565);
or U10748 (N_10748,N_10439,N_10452);
nor U10749 (N_10749,N_10575,N_10565);
nor U10750 (N_10750,N_10599,N_10462);
or U10751 (N_10751,N_10543,N_10531);
nand U10752 (N_10752,N_10595,N_10430);
or U10753 (N_10753,N_10595,N_10520);
and U10754 (N_10754,N_10545,N_10567);
nor U10755 (N_10755,N_10577,N_10486);
nor U10756 (N_10756,N_10582,N_10596);
nand U10757 (N_10757,N_10576,N_10590);
or U10758 (N_10758,N_10515,N_10430);
xor U10759 (N_10759,N_10462,N_10479);
nand U10760 (N_10760,N_10517,N_10512);
nand U10761 (N_10761,N_10541,N_10406);
xor U10762 (N_10762,N_10559,N_10543);
xor U10763 (N_10763,N_10503,N_10514);
nor U10764 (N_10764,N_10463,N_10584);
and U10765 (N_10765,N_10453,N_10530);
and U10766 (N_10766,N_10563,N_10494);
xnor U10767 (N_10767,N_10496,N_10559);
and U10768 (N_10768,N_10403,N_10541);
nor U10769 (N_10769,N_10535,N_10512);
or U10770 (N_10770,N_10586,N_10498);
or U10771 (N_10771,N_10580,N_10557);
xor U10772 (N_10772,N_10515,N_10517);
nor U10773 (N_10773,N_10543,N_10435);
xor U10774 (N_10774,N_10414,N_10467);
nand U10775 (N_10775,N_10529,N_10585);
xor U10776 (N_10776,N_10465,N_10487);
nand U10777 (N_10777,N_10494,N_10547);
nand U10778 (N_10778,N_10470,N_10426);
nand U10779 (N_10779,N_10512,N_10525);
xnor U10780 (N_10780,N_10546,N_10471);
xnor U10781 (N_10781,N_10488,N_10571);
xnor U10782 (N_10782,N_10402,N_10488);
xnor U10783 (N_10783,N_10446,N_10486);
xor U10784 (N_10784,N_10517,N_10511);
nand U10785 (N_10785,N_10412,N_10443);
nor U10786 (N_10786,N_10498,N_10577);
xnor U10787 (N_10787,N_10567,N_10513);
nand U10788 (N_10788,N_10449,N_10535);
nor U10789 (N_10789,N_10452,N_10426);
xnor U10790 (N_10790,N_10414,N_10496);
xor U10791 (N_10791,N_10472,N_10528);
nand U10792 (N_10792,N_10490,N_10518);
nand U10793 (N_10793,N_10595,N_10492);
nand U10794 (N_10794,N_10597,N_10553);
xnor U10795 (N_10795,N_10476,N_10562);
nand U10796 (N_10796,N_10582,N_10573);
or U10797 (N_10797,N_10562,N_10441);
xor U10798 (N_10798,N_10573,N_10407);
nor U10799 (N_10799,N_10530,N_10595);
nor U10800 (N_10800,N_10734,N_10714);
xnor U10801 (N_10801,N_10660,N_10699);
and U10802 (N_10802,N_10764,N_10792);
nand U10803 (N_10803,N_10669,N_10719);
nand U10804 (N_10804,N_10642,N_10743);
nor U10805 (N_10805,N_10671,N_10615);
nand U10806 (N_10806,N_10709,N_10613);
and U10807 (N_10807,N_10609,N_10696);
and U10808 (N_10808,N_10747,N_10630);
and U10809 (N_10809,N_10623,N_10791);
and U10810 (N_10810,N_10746,N_10620);
nand U10811 (N_10811,N_10658,N_10700);
nor U10812 (N_10812,N_10664,N_10775);
and U10813 (N_10813,N_10657,N_10683);
and U10814 (N_10814,N_10752,N_10766);
xnor U10815 (N_10815,N_10781,N_10799);
and U10816 (N_10816,N_10785,N_10693);
nor U10817 (N_10817,N_10684,N_10653);
nor U10818 (N_10818,N_10690,N_10685);
and U10819 (N_10819,N_10698,N_10726);
and U10820 (N_10820,N_10647,N_10728);
or U10821 (N_10821,N_10662,N_10672);
nor U10822 (N_10822,N_10617,N_10761);
nand U10823 (N_10823,N_10720,N_10749);
nand U10824 (N_10824,N_10605,N_10654);
or U10825 (N_10825,N_10704,N_10638);
nand U10826 (N_10826,N_10782,N_10784);
or U10827 (N_10827,N_10722,N_10602);
xnor U10828 (N_10828,N_10795,N_10649);
or U10829 (N_10829,N_10745,N_10670);
xnor U10830 (N_10830,N_10681,N_10675);
xnor U10831 (N_10831,N_10631,N_10611);
nor U10832 (N_10832,N_10629,N_10732);
xor U10833 (N_10833,N_10778,N_10652);
nand U10834 (N_10834,N_10679,N_10788);
and U10835 (N_10835,N_10773,N_10691);
and U10836 (N_10836,N_10783,N_10621);
or U10837 (N_10837,N_10689,N_10622);
nand U10838 (N_10838,N_10619,N_10637);
nor U10839 (N_10839,N_10707,N_10706);
nand U10840 (N_10840,N_10608,N_10759);
or U10841 (N_10841,N_10731,N_10600);
nor U10842 (N_10842,N_10760,N_10744);
and U10843 (N_10843,N_10718,N_10786);
or U10844 (N_10844,N_10686,N_10632);
and U10845 (N_10845,N_10741,N_10641);
nor U10846 (N_10846,N_10774,N_10651);
or U10847 (N_10847,N_10694,N_10695);
xor U10848 (N_10848,N_10659,N_10606);
xor U10849 (N_10849,N_10703,N_10650);
or U10850 (N_10850,N_10725,N_10762);
nor U10851 (N_10851,N_10750,N_10702);
and U10852 (N_10852,N_10771,N_10713);
and U10853 (N_10853,N_10717,N_10628);
and U10854 (N_10854,N_10798,N_10610);
nand U10855 (N_10855,N_10633,N_10757);
or U10856 (N_10856,N_10748,N_10730);
xor U10857 (N_10857,N_10680,N_10770);
or U10858 (N_10858,N_10627,N_10635);
nand U10859 (N_10859,N_10682,N_10779);
nand U10860 (N_10860,N_10678,N_10673);
nand U10861 (N_10861,N_10692,N_10655);
or U10862 (N_10862,N_10688,N_10789);
or U10863 (N_10863,N_10607,N_10667);
and U10864 (N_10864,N_10661,N_10735);
nor U10865 (N_10865,N_10636,N_10708);
and U10866 (N_10866,N_10776,N_10711);
or U10867 (N_10867,N_10705,N_10618);
or U10868 (N_10868,N_10780,N_10604);
xnor U10869 (N_10869,N_10674,N_10790);
nor U10870 (N_10870,N_10763,N_10616);
or U10871 (N_10871,N_10656,N_10754);
and U10872 (N_10872,N_10729,N_10742);
and U10873 (N_10873,N_10765,N_10710);
and U10874 (N_10874,N_10755,N_10665);
xor U10875 (N_10875,N_10666,N_10723);
xnor U10876 (N_10876,N_10612,N_10793);
and U10877 (N_10877,N_10769,N_10639);
or U10878 (N_10878,N_10756,N_10721);
xnor U10879 (N_10879,N_10668,N_10768);
and U10880 (N_10880,N_10626,N_10736);
nor U10881 (N_10881,N_10646,N_10663);
and U10882 (N_10882,N_10716,N_10727);
or U10883 (N_10883,N_10644,N_10740);
and U10884 (N_10884,N_10724,N_10625);
or U10885 (N_10885,N_10603,N_10751);
and U10886 (N_10886,N_10648,N_10738);
or U10887 (N_10887,N_10677,N_10733);
nand U10888 (N_10888,N_10697,N_10737);
or U10889 (N_10889,N_10777,N_10643);
xor U10890 (N_10890,N_10634,N_10712);
and U10891 (N_10891,N_10614,N_10715);
nand U10892 (N_10892,N_10645,N_10676);
nor U10893 (N_10893,N_10796,N_10767);
nand U10894 (N_10894,N_10624,N_10794);
nor U10895 (N_10895,N_10753,N_10687);
nor U10896 (N_10896,N_10701,N_10758);
nor U10897 (N_10897,N_10601,N_10739);
and U10898 (N_10898,N_10797,N_10787);
and U10899 (N_10899,N_10772,N_10640);
xnor U10900 (N_10900,N_10786,N_10661);
and U10901 (N_10901,N_10629,N_10640);
or U10902 (N_10902,N_10650,N_10620);
nand U10903 (N_10903,N_10613,N_10794);
nor U10904 (N_10904,N_10745,N_10638);
xor U10905 (N_10905,N_10713,N_10780);
and U10906 (N_10906,N_10632,N_10694);
nand U10907 (N_10907,N_10662,N_10708);
nand U10908 (N_10908,N_10691,N_10798);
nor U10909 (N_10909,N_10693,N_10658);
nor U10910 (N_10910,N_10725,N_10629);
nand U10911 (N_10911,N_10746,N_10608);
xnor U10912 (N_10912,N_10718,N_10753);
nor U10913 (N_10913,N_10650,N_10666);
nand U10914 (N_10914,N_10709,N_10610);
or U10915 (N_10915,N_10787,N_10786);
and U10916 (N_10916,N_10685,N_10710);
or U10917 (N_10917,N_10724,N_10612);
nor U10918 (N_10918,N_10714,N_10712);
nand U10919 (N_10919,N_10767,N_10768);
xnor U10920 (N_10920,N_10743,N_10694);
nor U10921 (N_10921,N_10715,N_10748);
or U10922 (N_10922,N_10663,N_10608);
xor U10923 (N_10923,N_10608,N_10789);
or U10924 (N_10924,N_10630,N_10727);
xnor U10925 (N_10925,N_10782,N_10689);
and U10926 (N_10926,N_10783,N_10735);
nor U10927 (N_10927,N_10794,N_10741);
or U10928 (N_10928,N_10783,N_10761);
nand U10929 (N_10929,N_10751,N_10621);
nand U10930 (N_10930,N_10651,N_10635);
xnor U10931 (N_10931,N_10651,N_10729);
nand U10932 (N_10932,N_10614,N_10781);
or U10933 (N_10933,N_10640,N_10799);
nor U10934 (N_10934,N_10755,N_10725);
nand U10935 (N_10935,N_10732,N_10675);
or U10936 (N_10936,N_10664,N_10653);
and U10937 (N_10937,N_10741,N_10740);
and U10938 (N_10938,N_10766,N_10682);
and U10939 (N_10939,N_10661,N_10643);
and U10940 (N_10940,N_10700,N_10639);
nor U10941 (N_10941,N_10667,N_10657);
nand U10942 (N_10942,N_10765,N_10609);
nand U10943 (N_10943,N_10628,N_10782);
or U10944 (N_10944,N_10627,N_10602);
or U10945 (N_10945,N_10695,N_10709);
or U10946 (N_10946,N_10788,N_10758);
or U10947 (N_10947,N_10676,N_10650);
nor U10948 (N_10948,N_10675,N_10637);
and U10949 (N_10949,N_10619,N_10785);
or U10950 (N_10950,N_10737,N_10760);
and U10951 (N_10951,N_10700,N_10600);
or U10952 (N_10952,N_10630,N_10784);
nand U10953 (N_10953,N_10654,N_10601);
xor U10954 (N_10954,N_10664,N_10643);
xnor U10955 (N_10955,N_10776,N_10757);
or U10956 (N_10956,N_10773,N_10795);
xor U10957 (N_10957,N_10667,N_10630);
or U10958 (N_10958,N_10623,N_10777);
nand U10959 (N_10959,N_10762,N_10794);
xnor U10960 (N_10960,N_10658,N_10614);
and U10961 (N_10961,N_10689,N_10662);
and U10962 (N_10962,N_10621,N_10731);
nand U10963 (N_10963,N_10791,N_10620);
xor U10964 (N_10964,N_10755,N_10739);
or U10965 (N_10965,N_10766,N_10750);
nor U10966 (N_10966,N_10652,N_10782);
xnor U10967 (N_10967,N_10613,N_10730);
xnor U10968 (N_10968,N_10638,N_10749);
xnor U10969 (N_10969,N_10740,N_10767);
nand U10970 (N_10970,N_10687,N_10615);
and U10971 (N_10971,N_10747,N_10752);
nor U10972 (N_10972,N_10632,N_10643);
xnor U10973 (N_10973,N_10663,N_10603);
nand U10974 (N_10974,N_10762,N_10644);
nor U10975 (N_10975,N_10619,N_10697);
xor U10976 (N_10976,N_10727,N_10745);
xor U10977 (N_10977,N_10748,N_10779);
and U10978 (N_10978,N_10681,N_10783);
nand U10979 (N_10979,N_10627,N_10696);
nand U10980 (N_10980,N_10634,N_10683);
and U10981 (N_10981,N_10785,N_10762);
xor U10982 (N_10982,N_10775,N_10767);
xnor U10983 (N_10983,N_10666,N_10685);
nor U10984 (N_10984,N_10655,N_10710);
and U10985 (N_10985,N_10672,N_10777);
xnor U10986 (N_10986,N_10698,N_10780);
nor U10987 (N_10987,N_10747,N_10772);
nor U10988 (N_10988,N_10728,N_10638);
nor U10989 (N_10989,N_10700,N_10777);
and U10990 (N_10990,N_10619,N_10620);
nor U10991 (N_10991,N_10739,N_10771);
nand U10992 (N_10992,N_10669,N_10759);
xor U10993 (N_10993,N_10607,N_10605);
xor U10994 (N_10994,N_10751,N_10706);
nor U10995 (N_10995,N_10792,N_10675);
and U10996 (N_10996,N_10645,N_10791);
nand U10997 (N_10997,N_10709,N_10664);
xnor U10998 (N_10998,N_10632,N_10708);
and U10999 (N_10999,N_10685,N_10606);
xor U11000 (N_11000,N_10853,N_10940);
or U11001 (N_11001,N_10991,N_10984);
or U11002 (N_11002,N_10909,N_10929);
and U11003 (N_11003,N_10855,N_10832);
nor U11004 (N_11004,N_10903,N_10948);
or U11005 (N_11005,N_10838,N_10992);
nand U11006 (N_11006,N_10931,N_10938);
nand U11007 (N_11007,N_10824,N_10939);
or U11008 (N_11008,N_10820,N_10881);
or U11009 (N_11009,N_10955,N_10959);
xor U11010 (N_11010,N_10864,N_10927);
and U11011 (N_11011,N_10829,N_10869);
nand U11012 (N_11012,N_10941,N_10932);
nor U11013 (N_11013,N_10949,N_10906);
nor U11014 (N_11014,N_10848,N_10995);
or U11015 (N_11015,N_10800,N_10850);
nor U11016 (N_11016,N_10930,N_10996);
or U11017 (N_11017,N_10997,N_10803);
or U11018 (N_11018,N_10828,N_10957);
or U11019 (N_11019,N_10841,N_10871);
nand U11020 (N_11020,N_10990,N_10918);
nand U11021 (N_11021,N_10920,N_10859);
or U11022 (N_11022,N_10845,N_10890);
nand U11023 (N_11023,N_10877,N_10846);
or U11024 (N_11024,N_10891,N_10862);
or U11025 (N_11025,N_10937,N_10925);
nand U11026 (N_11026,N_10809,N_10969);
and U11027 (N_11027,N_10921,N_10895);
nor U11028 (N_11028,N_10954,N_10886);
nand U11029 (N_11029,N_10880,N_10946);
nand U11030 (N_11030,N_10973,N_10870);
nor U11031 (N_11031,N_10802,N_10807);
xnor U11032 (N_11032,N_10847,N_10953);
and U11033 (N_11033,N_10823,N_10804);
nand U11034 (N_11034,N_10867,N_10858);
and U11035 (N_11035,N_10952,N_10956);
xor U11036 (N_11036,N_10908,N_10876);
xnor U11037 (N_11037,N_10968,N_10960);
xnor U11038 (N_11038,N_10900,N_10801);
nor U11039 (N_11039,N_10888,N_10872);
or U11040 (N_11040,N_10989,N_10983);
xnor U11041 (N_11041,N_10819,N_10981);
nand U11042 (N_11042,N_10893,N_10896);
and U11043 (N_11043,N_10982,N_10905);
xor U11044 (N_11044,N_10844,N_10854);
nor U11045 (N_11045,N_10993,N_10882);
and U11046 (N_11046,N_10833,N_10928);
or U11047 (N_11047,N_10813,N_10810);
or U11048 (N_11048,N_10985,N_10977);
nand U11049 (N_11049,N_10874,N_10868);
and U11050 (N_11050,N_10904,N_10966);
xor U11051 (N_11051,N_10889,N_10816);
and U11052 (N_11052,N_10971,N_10916);
xor U11053 (N_11053,N_10808,N_10933);
or U11054 (N_11054,N_10897,N_10923);
and U11055 (N_11055,N_10978,N_10894);
or U11056 (N_11056,N_10986,N_10914);
nand U11057 (N_11057,N_10972,N_10861);
and U11058 (N_11058,N_10962,N_10822);
xor U11059 (N_11059,N_10851,N_10965);
or U11060 (N_11060,N_10817,N_10950);
and U11061 (N_11061,N_10866,N_10961);
nand U11062 (N_11062,N_10849,N_10924);
xnor U11063 (N_11063,N_10998,N_10834);
xnor U11064 (N_11064,N_10852,N_10974);
nand U11065 (N_11065,N_10907,N_10839);
nand U11066 (N_11066,N_10976,N_10860);
xnor U11067 (N_11067,N_10910,N_10901);
and U11068 (N_11068,N_10935,N_10856);
xnor U11069 (N_11069,N_10915,N_10942);
nand U11070 (N_11070,N_10963,N_10875);
nand U11071 (N_11071,N_10812,N_10944);
and U11072 (N_11072,N_10934,N_10936);
xnor U11073 (N_11073,N_10919,N_10964);
nor U11074 (N_11074,N_10979,N_10887);
nor U11075 (N_11075,N_10951,N_10912);
and U11076 (N_11076,N_10994,N_10857);
nor U11077 (N_11077,N_10999,N_10873);
or U11078 (N_11078,N_10945,N_10902);
nor U11079 (N_11079,N_10892,N_10913);
xor U11080 (N_11080,N_10884,N_10814);
or U11081 (N_11081,N_10885,N_10899);
and U11082 (N_11082,N_10883,N_10922);
or U11083 (N_11083,N_10825,N_10826);
nand U11084 (N_11084,N_10911,N_10821);
nor U11085 (N_11085,N_10836,N_10827);
or U11086 (N_11086,N_10811,N_10878);
and U11087 (N_11087,N_10898,N_10818);
and U11088 (N_11088,N_10842,N_10970);
nor U11089 (N_11089,N_10947,N_10863);
xnor U11090 (N_11090,N_10943,N_10987);
nand U11091 (N_11091,N_10835,N_10967);
nor U11092 (N_11092,N_10815,N_10879);
nor U11093 (N_11093,N_10837,N_10975);
xor U11094 (N_11094,N_10865,N_10830);
nor U11095 (N_11095,N_10958,N_10805);
nor U11096 (N_11096,N_10843,N_10980);
nor U11097 (N_11097,N_10988,N_10840);
nor U11098 (N_11098,N_10806,N_10926);
xnor U11099 (N_11099,N_10831,N_10917);
nor U11100 (N_11100,N_10830,N_10892);
nand U11101 (N_11101,N_10926,N_10850);
xor U11102 (N_11102,N_10916,N_10816);
xor U11103 (N_11103,N_10861,N_10988);
xor U11104 (N_11104,N_10913,N_10808);
or U11105 (N_11105,N_10957,N_10934);
nor U11106 (N_11106,N_10887,N_10813);
nor U11107 (N_11107,N_10954,N_10943);
nand U11108 (N_11108,N_10891,N_10976);
nand U11109 (N_11109,N_10998,N_10876);
xor U11110 (N_11110,N_10940,N_10813);
xor U11111 (N_11111,N_10917,N_10815);
or U11112 (N_11112,N_10863,N_10896);
nor U11113 (N_11113,N_10999,N_10816);
nor U11114 (N_11114,N_10818,N_10944);
nand U11115 (N_11115,N_10842,N_10909);
and U11116 (N_11116,N_10827,N_10897);
xor U11117 (N_11117,N_10846,N_10872);
nor U11118 (N_11118,N_10819,N_10976);
nor U11119 (N_11119,N_10841,N_10992);
nor U11120 (N_11120,N_10994,N_10966);
and U11121 (N_11121,N_10889,N_10838);
xnor U11122 (N_11122,N_10802,N_10961);
and U11123 (N_11123,N_10977,N_10860);
xor U11124 (N_11124,N_10845,N_10963);
or U11125 (N_11125,N_10897,N_10949);
nand U11126 (N_11126,N_10926,N_10942);
and U11127 (N_11127,N_10801,N_10881);
and U11128 (N_11128,N_10930,N_10843);
and U11129 (N_11129,N_10820,N_10897);
xnor U11130 (N_11130,N_10905,N_10964);
nand U11131 (N_11131,N_10868,N_10811);
or U11132 (N_11132,N_10811,N_10841);
nor U11133 (N_11133,N_10880,N_10974);
xor U11134 (N_11134,N_10811,N_10942);
nor U11135 (N_11135,N_10887,N_10825);
xnor U11136 (N_11136,N_10916,N_10974);
or U11137 (N_11137,N_10874,N_10987);
xnor U11138 (N_11138,N_10810,N_10824);
nor U11139 (N_11139,N_10901,N_10952);
nand U11140 (N_11140,N_10806,N_10936);
nor U11141 (N_11141,N_10963,N_10825);
nand U11142 (N_11142,N_10966,N_10894);
and U11143 (N_11143,N_10974,N_10957);
nand U11144 (N_11144,N_10960,N_10839);
nor U11145 (N_11145,N_10811,N_10994);
nor U11146 (N_11146,N_10919,N_10873);
nand U11147 (N_11147,N_10847,N_10886);
and U11148 (N_11148,N_10947,N_10973);
xnor U11149 (N_11149,N_10901,N_10935);
nor U11150 (N_11150,N_10857,N_10989);
and U11151 (N_11151,N_10987,N_10903);
xor U11152 (N_11152,N_10901,N_10960);
xnor U11153 (N_11153,N_10902,N_10833);
nand U11154 (N_11154,N_10864,N_10815);
nand U11155 (N_11155,N_10839,N_10946);
nor U11156 (N_11156,N_10964,N_10915);
xor U11157 (N_11157,N_10846,N_10863);
nor U11158 (N_11158,N_10949,N_10852);
xnor U11159 (N_11159,N_10898,N_10812);
nand U11160 (N_11160,N_10805,N_10982);
xor U11161 (N_11161,N_10851,N_10897);
and U11162 (N_11162,N_10852,N_10903);
and U11163 (N_11163,N_10981,N_10841);
and U11164 (N_11164,N_10903,N_10980);
nor U11165 (N_11165,N_10841,N_10822);
xnor U11166 (N_11166,N_10978,N_10895);
or U11167 (N_11167,N_10947,N_10930);
nand U11168 (N_11168,N_10905,N_10830);
xor U11169 (N_11169,N_10956,N_10836);
xnor U11170 (N_11170,N_10927,N_10976);
and U11171 (N_11171,N_10892,N_10983);
xnor U11172 (N_11172,N_10878,N_10940);
and U11173 (N_11173,N_10800,N_10852);
nor U11174 (N_11174,N_10902,N_10856);
nand U11175 (N_11175,N_10921,N_10869);
xnor U11176 (N_11176,N_10989,N_10827);
or U11177 (N_11177,N_10992,N_10984);
nor U11178 (N_11178,N_10874,N_10811);
nor U11179 (N_11179,N_10808,N_10971);
xor U11180 (N_11180,N_10997,N_10861);
nor U11181 (N_11181,N_10949,N_10826);
or U11182 (N_11182,N_10871,N_10853);
or U11183 (N_11183,N_10908,N_10814);
nor U11184 (N_11184,N_10887,N_10837);
nand U11185 (N_11185,N_10984,N_10902);
or U11186 (N_11186,N_10809,N_10859);
xor U11187 (N_11187,N_10839,N_10994);
and U11188 (N_11188,N_10983,N_10925);
or U11189 (N_11189,N_10852,N_10893);
nor U11190 (N_11190,N_10899,N_10815);
nand U11191 (N_11191,N_10998,N_10978);
or U11192 (N_11192,N_10818,N_10975);
or U11193 (N_11193,N_10876,N_10890);
xnor U11194 (N_11194,N_10929,N_10990);
nand U11195 (N_11195,N_10950,N_10972);
and U11196 (N_11196,N_10804,N_10957);
xnor U11197 (N_11197,N_10887,N_10991);
or U11198 (N_11198,N_10931,N_10961);
nand U11199 (N_11199,N_10870,N_10902);
or U11200 (N_11200,N_11149,N_11132);
and U11201 (N_11201,N_11113,N_11161);
nor U11202 (N_11202,N_11034,N_11114);
xnor U11203 (N_11203,N_11062,N_11061);
and U11204 (N_11204,N_11126,N_11127);
nor U11205 (N_11205,N_11013,N_11072);
nand U11206 (N_11206,N_11028,N_11185);
or U11207 (N_11207,N_11170,N_11165);
or U11208 (N_11208,N_11036,N_11105);
nor U11209 (N_11209,N_11043,N_11085);
xnor U11210 (N_11210,N_11003,N_11002);
xor U11211 (N_11211,N_11092,N_11186);
nor U11212 (N_11212,N_11141,N_11096);
nor U11213 (N_11213,N_11053,N_11175);
or U11214 (N_11214,N_11071,N_11176);
or U11215 (N_11215,N_11146,N_11029);
xnor U11216 (N_11216,N_11007,N_11156);
xnor U11217 (N_11217,N_11058,N_11065);
and U11218 (N_11218,N_11172,N_11129);
and U11219 (N_11219,N_11154,N_11081);
and U11220 (N_11220,N_11000,N_11120);
nand U11221 (N_11221,N_11138,N_11038);
xnor U11222 (N_11222,N_11106,N_11198);
xor U11223 (N_11223,N_11192,N_11004);
nand U11224 (N_11224,N_11168,N_11103);
and U11225 (N_11225,N_11150,N_11164);
nor U11226 (N_11226,N_11181,N_11073);
nor U11227 (N_11227,N_11115,N_11193);
nor U11228 (N_11228,N_11083,N_11032);
and U11229 (N_11229,N_11035,N_11143);
xnor U11230 (N_11230,N_11060,N_11112);
xor U11231 (N_11231,N_11148,N_11130);
or U11232 (N_11232,N_11079,N_11180);
and U11233 (N_11233,N_11151,N_11191);
nand U11234 (N_11234,N_11009,N_11091);
and U11235 (N_11235,N_11031,N_11016);
xnor U11236 (N_11236,N_11160,N_11006);
nor U11237 (N_11237,N_11040,N_11090);
and U11238 (N_11238,N_11021,N_11199);
and U11239 (N_11239,N_11057,N_11102);
or U11240 (N_11240,N_11158,N_11042);
nand U11241 (N_11241,N_11144,N_11179);
or U11242 (N_11242,N_11069,N_11037);
and U11243 (N_11243,N_11008,N_11015);
xor U11244 (N_11244,N_11173,N_11124);
nand U11245 (N_11245,N_11135,N_11030);
nor U11246 (N_11246,N_11068,N_11117);
and U11247 (N_11247,N_11195,N_11022);
or U11248 (N_11248,N_11104,N_11194);
and U11249 (N_11249,N_11190,N_11100);
nor U11250 (N_11250,N_11084,N_11018);
or U11251 (N_11251,N_11070,N_11041);
or U11252 (N_11252,N_11145,N_11111);
nand U11253 (N_11253,N_11188,N_11098);
nand U11254 (N_11254,N_11128,N_11086);
nor U11255 (N_11255,N_11174,N_11152);
and U11256 (N_11256,N_11052,N_11118);
and U11257 (N_11257,N_11046,N_11163);
nand U11258 (N_11258,N_11121,N_11045);
or U11259 (N_11259,N_11082,N_11020);
xor U11260 (N_11260,N_11099,N_11122);
or U11261 (N_11261,N_11159,N_11017);
and U11262 (N_11262,N_11044,N_11177);
nor U11263 (N_11263,N_11183,N_11169);
nor U11264 (N_11264,N_11184,N_11134);
nor U11265 (N_11265,N_11139,N_11049);
or U11266 (N_11266,N_11131,N_11064);
nand U11267 (N_11267,N_11095,N_11024);
nand U11268 (N_11268,N_11012,N_11087);
and U11269 (N_11269,N_11182,N_11050);
or U11270 (N_11270,N_11055,N_11110);
or U11271 (N_11271,N_11067,N_11014);
nor U11272 (N_11272,N_11054,N_11048);
or U11273 (N_11273,N_11094,N_11047);
xor U11274 (N_11274,N_11051,N_11140);
xnor U11275 (N_11275,N_11116,N_11019);
nor U11276 (N_11276,N_11167,N_11033);
nor U11277 (N_11277,N_11137,N_11189);
nand U11278 (N_11278,N_11166,N_11025);
or U11279 (N_11279,N_11107,N_11101);
or U11280 (N_11280,N_11001,N_11056);
nand U11281 (N_11281,N_11157,N_11026);
nor U11282 (N_11282,N_11027,N_11023);
xor U11283 (N_11283,N_11077,N_11142);
and U11284 (N_11284,N_11136,N_11178);
or U11285 (N_11285,N_11187,N_11125);
nor U11286 (N_11286,N_11133,N_11011);
nand U11287 (N_11287,N_11153,N_11080);
nor U11288 (N_11288,N_11063,N_11162);
and U11289 (N_11289,N_11089,N_11066);
and U11290 (N_11290,N_11088,N_11123);
nand U11291 (N_11291,N_11119,N_11093);
and U11292 (N_11292,N_11097,N_11039);
nand U11293 (N_11293,N_11075,N_11074);
nand U11294 (N_11294,N_11197,N_11155);
nand U11295 (N_11295,N_11147,N_11010);
xnor U11296 (N_11296,N_11078,N_11005);
nor U11297 (N_11297,N_11109,N_11196);
and U11298 (N_11298,N_11076,N_11108);
nor U11299 (N_11299,N_11059,N_11171);
nor U11300 (N_11300,N_11107,N_11124);
nor U11301 (N_11301,N_11061,N_11122);
nor U11302 (N_11302,N_11045,N_11153);
or U11303 (N_11303,N_11137,N_11026);
nor U11304 (N_11304,N_11162,N_11155);
or U11305 (N_11305,N_11064,N_11031);
nor U11306 (N_11306,N_11040,N_11096);
nand U11307 (N_11307,N_11177,N_11191);
xnor U11308 (N_11308,N_11141,N_11153);
xor U11309 (N_11309,N_11146,N_11187);
xnor U11310 (N_11310,N_11005,N_11037);
nand U11311 (N_11311,N_11043,N_11106);
nand U11312 (N_11312,N_11152,N_11060);
and U11313 (N_11313,N_11130,N_11035);
and U11314 (N_11314,N_11072,N_11095);
and U11315 (N_11315,N_11047,N_11171);
or U11316 (N_11316,N_11121,N_11095);
nand U11317 (N_11317,N_11058,N_11038);
and U11318 (N_11318,N_11121,N_11186);
xnor U11319 (N_11319,N_11019,N_11107);
or U11320 (N_11320,N_11009,N_11092);
xnor U11321 (N_11321,N_11126,N_11062);
or U11322 (N_11322,N_11007,N_11197);
nor U11323 (N_11323,N_11166,N_11030);
and U11324 (N_11324,N_11055,N_11163);
and U11325 (N_11325,N_11061,N_11030);
nand U11326 (N_11326,N_11153,N_11046);
xor U11327 (N_11327,N_11089,N_11183);
or U11328 (N_11328,N_11109,N_11064);
nand U11329 (N_11329,N_11066,N_11044);
xnor U11330 (N_11330,N_11180,N_11148);
and U11331 (N_11331,N_11025,N_11014);
and U11332 (N_11332,N_11194,N_11195);
xnor U11333 (N_11333,N_11152,N_11139);
and U11334 (N_11334,N_11081,N_11107);
nor U11335 (N_11335,N_11167,N_11149);
and U11336 (N_11336,N_11098,N_11067);
nor U11337 (N_11337,N_11181,N_11000);
nor U11338 (N_11338,N_11033,N_11173);
nand U11339 (N_11339,N_11144,N_11113);
xor U11340 (N_11340,N_11014,N_11125);
nor U11341 (N_11341,N_11065,N_11134);
or U11342 (N_11342,N_11004,N_11038);
and U11343 (N_11343,N_11153,N_11169);
nand U11344 (N_11344,N_11036,N_11149);
or U11345 (N_11345,N_11011,N_11114);
or U11346 (N_11346,N_11134,N_11164);
and U11347 (N_11347,N_11148,N_11085);
nand U11348 (N_11348,N_11133,N_11068);
xnor U11349 (N_11349,N_11014,N_11147);
or U11350 (N_11350,N_11139,N_11165);
and U11351 (N_11351,N_11061,N_11054);
nand U11352 (N_11352,N_11178,N_11094);
nand U11353 (N_11353,N_11173,N_11152);
and U11354 (N_11354,N_11120,N_11039);
nor U11355 (N_11355,N_11196,N_11057);
nor U11356 (N_11356,N_11151,N_11072);
nand U11357 (N_11357,N_11132,N_11162);
nor U11358 (N_11358,N_11105,N_11183);
and U11359 (N_11359,N_11135,N_11059);
and U11360 (N_11360,N_11020,N_11038);
xor U11361 (N_11361,N_11033,N_11150);
nor U11362 (N_11362,N_11119,N_11154);
xor U11363 (N_11363,N_11007,N_11152);
nand U11364 (N_11364,N_11121,N_11181);
nand U11365 (N_11365,N_11156,N_11111);
nor U11366 (N_11366,N_11110,N_11180);
and U11367 (N_11367,N_11023,N_11143);
or U11368 (N_11368,N_11005,N_11084);
or U11369 (N_11369,N_11001,N_11009);
or U11370 (N_11370,N_11181,N_11103);
or U11371 (N_11371,N_11174,N_11093);
or U11372 (N_11372,N_11018,N_11080);
xor U11373 (N_11373,N_11141,N_11071);
xor U11374 (N_11374,N_11155,N_11032);
xor U11375 (N_11375,N_11013,N_11066);
xnor U11376 (N_11376,N_11051,N_11154);
and U11377 (N_11377,N_11054,N_11186);
xnor U11378 (N_11378,N_11023,N_11138);
xor U11379 (N_11379,N_11176,N_11010);
nor U11380 (N_11380,N_11115,N_11070);
nor U11381 (N_11381,N_11134,N_11077);
or U11382 (N_11382,N_11164,N_11075);
nor U11383 (N_11383,N_11112,N_11147);
nor U11384 (N_11384,N_11134,N_11005);
or U11385 (N_11385,N_11031,N_11090);
xor U11386 (N_11386,N_11165,N_11120);
or U11387 (N_11387,N_11192,N_11117);
and U11388 (N_11388,N_11171,N_11076);
and U11389 (N_11389,N_11155,N_11075);
and U11390 (N_11390,N_11167,N_11067);
and U11391 (N_11391,N_11198,N_11044);
or U11392 (N_11392,N_11082,N_11100);
nor U11393 (N_11393,N_11064,N_11169);
and U11394 (N_11394,N_11032,N_11059);
or U11395 (N_11395,N_11007,N_11097);
xor U11396 (N_11396,N_11111,N_11050);
or U11397 (N_11397,N_11170,N_11195);
xor U11398 (N_11398,N_11055,N_11182);
nand U11399 (N_11399,N_11032,N_11006);
or U11400 (N_11400,N_11260,N_11209);
or U11401 (N_11401,N_11397,N_11263);
nor U11402 (N_11402,N_11319,N_11269);
nand U11403 (N_11403,N_11289,N_11308);
and U11404 (N_11404,N_11213,N_11382);
nand U11405 (N_11405,N_11371,N_11241);
and U11406 (N_11406,N_11337,N_11349);
nor U11407 (N_11407,N_11265,N_11375);
xnor U11408 (N_11408,N_11376,N_11232);
nor U11409 (N_11409,N_11240,N_11330);
xor U11410 (N_11410,N_11243,N_11219);
xnor U11411 (N_11411,N_11208,N_11212);
xnor U11412 (N_11412,N_11314,N_11234);
and U11413 (N_11413,N_11246,N_11211);
xnor U11414 (N_11414,N_11281,N_11248);
nor U11415 (N_11415,N_11298,N_11293);
xnor U11416 (N_11416,N_11365,N_11249);
nor U11417 (N_11417,N_11292,N_11318);
or U11418 (N_11418,N_11374,N_11291);
nand U11419 (N_11419,N_11242,N_11313);
nor U11420 (N_11420,N_11282,N_11297);
nor U11421 (N_11421,N_11202,N_11331);
or U11422 (N_11422,N_11384,N_11256);
xnor U11423 (N_11423,N_11381,N_11316);
and U11424 (N_11424,N_11327,N_11227);
nand U11425 (N_11425,N_11245,N_11262);
xnor U11426 (N_11426,N_11205,N_11317);
xor U11427 (N_11427,N_11323,N_11224);
xor U11428 (N_11428,N_11367,N_11343);
or U11429 (N_11429,N_11392,N_11206);
or U11430 (N_11430,N_11273,N_11370);
and U11431 (N_11431,N_11286,N_11362);
or U11432 (N_11432,N_11244,N_11250);
nand U11433 (N_11433,N_11388,N_11237);
nand U11434 (N_11434,N_11259,N_11257);
nand U11435 (N_11435,N_11334,N_11336);
and U11436 (N_11436,N_11261,N_11214);
nand U11437 (N_11437,N_11275,N_11210);
and U11438 (N_11438,N_11307,N_11268);
or U11439 (N_11439,N_11270,N_11215);
and U11440 (N_11440,N_11221,N_11277);
nand U11441 (N_11441,N_11220,N_11312);
nand U11442 (N_11442,N_11225,N_11355);
nand U11443 (N_11443,N_11373,N_11357);
xor U11444 (N_11444,N_11352,N_11372);
and U11445 (N_11445,N_11368,N_11235);
or U11446 (N_11446,N_11299,N_11229);
nor U11447 (N_11447,N_11353,N_11287);
and U11448 (N_11448,N_11283,N_11267);
xor U11449 (N_11449,N_11254,N_11333);
nor U11450 (N_11450,N_11358,N_11394);
and U11451 (N_11451,N_11340,N_11217);
nand U11452 (N_11452,N_11395,N_11332);
nand U11453 (N_11453,N_11320,N_11310);
nand U11454 (N_11454,N_11284,N_11276);
and U11455 (N_11455,N_11347,N_11322);
and U11456 (N_11456,N_11363,N_11338);
xnor U11457 (N_11457,N_11218,N_11354);
and U11458 (N_11458,N_11345,N_11369);
and U11459 (N_11459,N_11390,N_11290);
xor U11460 (N_11460,N_11328,N_11296);
nand U11461 (N_11461,N_11251,N_11207);
and U11462 (N_11462,N_11315,N_11351);
or U11463 (N_11463,N_11386,N_11383);
nor U11464 (N_11464,N_11366,N_11360);
or U11465 (N_11465,N_11342,N_11398);
and U11466 (N_11466,N_11385,N_11396);
nand U11467 (N_11467,N_11377,N_11200);
or U11468 (N_11468,N_11272,N_11239);
and U11469 (N_11469,N_11359,N_11387);
or U11470 (N_11470,N_11231,N_11285);
and U11471 (N_11471,N_11238,N_11203);
nor U11472 (N_11472,N_11216,N_11223);
nor U11473 (N_11473,N_11258,N_11339);
and U11474 (N_11474,N_11230,N_11306);
nand U11475 (N_11475,N_11378,N_11393);
and U11476 (N_11476,N_11391,N_11271);
and U11477 (N_11477,N_11288,N_11350);
nand U11478 (N_11478,N_11348,N_11255);
nand U11479 (N_11479,N_11356,N_11300);
nor U11480 (N_11480,N_11329,N_11321);
nor U11481 (N_11481,N_11253,N_11311);
nor U11482 (N_11482,N_11264,N_11326);
nor U11483 (N_11483,N_11201,N_11204);
xnor U11484 (N_11484,N_11304,N_11274);
nor U11485 (N_11485,N_11361,N_11278);
xor U11486 (N_11486,N_11309,N_11341);
nor U11487 (N_11487,N_11302,N_11233);
or U11488 (N_11488,N_11226,N_11379);
or U11489 (N_11489,N_11305,N_11279);
xor U11490 (N_11490,N_11364,N_11325);
nor U11491 (N_11491,N_11252,N_11344);
or U11492 (N_11492,N_11301,N_11294);
or U11493 (N_11493,N_11266,N_11389);
nand U11494 (N_11494,N_11247,N_11399);
nand U11495 (N_11495,N_11324,N_11335);
nor U11496 (N_11496,N_11236,N_11380);
nand U11497 (N_11497,N_11295,N_11222);
xor U11498 (N_11498,N_11280,N_11346);
nand U11499 (N_11499,N_11303,N_11228);
nor U11500 (N_11500,N_11214,N_11354);
nand U11501 (N_11501,N_11312,N_11329);
or U11502 (N_11502,N_11298,N_11255);
xor U11503 (N_11503,N_11270,N_11235);
and U11504 (N_11504,N_11362,N_11208);
xnor U11505 (N_11505,N_11373,N_11331);
xnor U11506 (N_11506,N_11355,N_11269);
and U11507 (N_11507,N_11259,N_11226);
or U11508 (N_11508,N_11242,N_11376);
nor U11509 (N_11509,N_11351,N_11288);
nor U11510 (N_11510,N_11373,N_11339);
xor U11511 (N_11511,N_11327,N_11387);
nor U11512 (N_11512,N_11371,N_11216);
xor U11513 (N_11513,N_11336,N_11331);
or U11514 (N_11514,N_11213,N_11298);
nor U11515 (N_11515,N_11233,N_11386);
nor U11516 (N_11516,N_11269,N_11341);
nor U11517 (N_11517,N_11250,N_11201);
nor U11518 (N_11518,N_11391,N_11390);
nand U11519 (N_11519,N_11379,N_11219);
nand U11520 (N_11520,N_11287,N_11348);
nor U11521 (N_11521,N_11203,N_11353);
xor U11522 (N_11522,N_11390,N_11269);
or U11523 (N_11523,N_11357,N_11361);
xor U11524 (N_11524,N_11272,N_11352);
xor U11525 (N_11525,N_11251,N_11264);
xnor U11526 (N_11526,N_11330,N_11229);
or U11527 (N_11527,N_11263,N_11326);
and U11528 (N_11528,N_11373,N_11316);
or U11529 (N_11529,N_11345,N_11328);
nand U11530 (N_11530,N_11320,N_11324);
xnor U11531 (N_11531,N_11305,N_11295);
nor U11532 (N_11532,N_11327,N_11261);
nor U11533 (N_11533,N_11344,N_11330);
xor U11534 (N_11534,N_11208,N_11395);
or U11535 (N_11535,N_11306,N_11239);
and U11536 (N_11536,N_11398,N_11264);
nand U11537 (N_11537,N_11248,N_11213);
nor U11538 (N_11538,N_11222,N_11234);
or U11539 (N_11539,N_11264,N_11374);
or U11540 (N_11540,N_11237,N_11233);
nand U11541 (N_11541,N_11263,N_11324);
nor U11542 (N_11542,N_11330,N_11273);
and U11543 (N_11543,N_11258,N_11200);
and U11544 (N_11544,N_11251,N_11218);
or U11545 (N_11545,N_11293,N_11249);
and U11546 (N_11546,N_11205,N_11241);
and U11547 (N_11547,N_11295,N_11313);
or U11548 (N_11548,N_11275,N_11334);
and U11549 (N_11549,N_11279,N_11320);
nor U11550 (N_11550,N_11221,N_11357);
nor U11551 (N_11551,N_11248,N_11336);
xnor U11552 (N_11552,N_11276,N_11237);
nor U11553 (N_11553,N_11239,N_11215);
nor U11554 (N_11554,N_11244,N_11376);
xnor U11555 (N_11555,N_11206,N_11357);
or U11556 (N_11556,N_11213,N_11376);
nor U11557 (N_11557,N_11300,N_11396);
and U11558 (N_11558,N_11202,N_11394);
or U11559 (N_11559,N_11377,N_11364);
and U11560 (N_11560,N_11289,N_11295);
xor U11561 (N_11561,N_11380,N_11338);
and U11562 (N_11562,N_11379,N_11209);
nor U11563 (N_11563,N_11314,N_11283);
or U11564 (N_11564,N_11349,N_11335);
or U11565 (N_11565,N_11220,N_11302);
and U11566 (N_11566,N_11358,N_11351);
or U11567 (N_11567,N_11253,N_11242);
or U11568 (N_11568,N_11385,N_11217);
xnor U11569 (N_11569,N_11206,N_11255);
nor U11570 (N_11570,N_11255,N_11299);
or U11571 (N_11571,N_11268,N_11377);
nand U11572 (N_11572,N_11379,N_11296);
or U11573 (N_11573,N_11335,N_11392);
and U11574 (N_11574,N_11324,N_11336);
and U11575 (N_11575,N_11332,N_11337);
nor U11576 (N_11576,N_11308,N_11300);
xnor U11577 (N_11577,N_11360,N_11238);
xor U11578 (N_11578,N_11388,N_11251);
nor U11579 (N_11579,N_11395,N_11317);
xor U11580 (N_11580,N_11207,N_11297);
and U11581 (N_11581,N_11375,N_11390);
xnor U11582 (N_11582,N_11321,N_11387);
nand U11583 (N_11583,N_11274,N_11307);
or U11584 (N_11584,N_11210,N_11380);
and U11585 (N_11585,N_11272,N_11274);
or U11586 (N_11586,N_11267,N_11361);
or U11587 (N_11587,N_11393,N_11386);
nand U11588 (N_11588,N_11295,N_11397);
nand U11589 (N_11589,N_11241,N_11254);
and U11590 (N_11590,N_11218,N_11200);
xnor U11591 (N_11591,N_11267,N_11323);
and U11592 (N_11592,N_11239,N_11360);
xor U11593 (N_11593,N_11218,N_11364);
or U11594 (N_11594,N_11376,N_11397);
nand U11595 (N_11595,N_11373,N_11244);
xnor U11596 (N_11596,N_11214,N_11253);
xnor U11597 (N_11597,N_11264,N_11367);
and U11598 (N_11598,N_11223,N_11308);
nand U11599 (N_11599,N_11211,N_11305);
nand U11600 (N_11600,N_11464,N_11462);
xor U11601 (N_11601,N_11515,N_11575);
or U11602 (N_11602,N_11455,N_11514);
nand U11603 (N_11603,N_11457,N_11424);
or U11604 (N_11604,N_11473,N_11489);
xnor U11605 (N_11605,N_11454,N_11491);
nor U11606 (N_11606,N_11484,N_11532);
nand U11607 (N_11607,N_11443,N_11446);
nor U11608 (N_11608,N_11472,N_11400);
nor U11609 (N_11609,N_11411,N_11519);
and U11610 (N_11610,N_11427,N_11414);
nand U11611 (N_11611,N_11487,N_11509);
and U11612 (N_11612,N_11574,N_11564);
and U11613 (N_11613,N_11552,N_11438);
xor U11614 (N_11614,N_11572,N_11577);
nand U11615 (N_11615,N_11520,N_11415);
xnor U11616 (N_11616,N_11579,N_11401);
nand U11617 (N_11617,N_11507,N_11420);
nand U11618 (N_11618,N_11444,N_11486);
and U11619 (N_11619,N_11550,N_11530);
and U11620 (N_11620,N_11566,N_11592);
nand U11621 (N_11621,N_11521,N_11481);
or U11622 (N_11622,N_11527,N_11501);
xor U11623 (N_11623,N_11474,N_11508);
xor U11624 (N_11624,N_11493,N_11593);
nor U11625 (N_11625,N_11548,N_11466);
or U11626 (N_11626,N_11576,N_11429);
nand U11627 (N_11627,N_11560,N_11513);
xor U11628 (N_11628,N_11423,N_11496);
nand U11629 (N_11629,N_11456,N_11459);
nor U11630 (N_11630,N_11436,N_11442);
xor U11631 (N_11631,N_11428,N_11495);
or U11632 (N_11632,N_11525,N_11505);
nand U11633 (N_11633,N_11479,N_11553);
or U11634 (N_11634,N_11555,N_11433);
nor U11635 (N_11635,N_11503,N_11412);
nand U11636 (N_11636,N_11450,N_11586);
or U11637 (N_11637,N_11535,N_11430);
nand U11638 (N_11638,N_11588,N_11598);
and U11639 (N_11639,N_11539,N_11494);
xor U11640 (N_11640,N_11522,N_11589);
or U11641 (N_11641,N_11500,N_11565);
xnor U11642 (N_11642,N_11437,N_11554);
nand U11643 (N_11643,N_11453,N_11562);
or U11644 (N_11644,N_11461,N_11458);
and U11645 (N_11645,N_11528,N_11476);
nand U11646 (N_11646,N_11425,N_11526);
xor U11647 (N_11647,N_11584,N_11595);
or U11648 (N_11648,N_11426,N_11547);
nor U11649 (N_11649,N_11537,N_11490);
nor U11650 (N_11650,N_11523,N_11445);
or U11651 (N_11651,N_11540,N_11568);
or U11652 (N_11652,N_11439,N_11583);
nor U11653 (N_11653,N_11511,N_11417);
nor U11654 (N_11654,N_11483,N_11406);
or U11655 (N_11655,N_11558,N_11416);
nor U11656 (N_11656,N_11549,N_11434);
nand U11657 (N_11657,N_11534,N_11460);
and U11658 (N_11658,N_11512,N_11557);
and U11659 (N_11659,N_11599,N_11573);
nor U11660 (N_11660,N_11402,N_11469);
nand U11661 (N_11661,N_11538,N_11410);
nand U11662 (N_11662,N_11529,N_11404);
nor U11663 (N_11663,N_11421,N_11440);
xnor U11664 (N_11664,N_11435,N_11470);
nand U11665 (N_11665,N_11492,N_11485);
nand U11666 (N_11666,N_11452,N_11488);
xor U11667 (N_11667,N_11546,N_11447);
xor U11668 (N_11668,N_11441,N_11449);
or U11669 (N_11669,N_11597,N_11533);
nand U11670 (N_11670,N_11502,N_11578);
xor U11671 (N_11671,N_11518,N_11563);
or U11672 (N_11672,N_11516,N_11536);
nand U11673 (N_11673,N_11477,N_11585);
nand U11674 (N_11674,N_11497,N_11544);
and U11675 (N_11675,N_11531,N_11506);
or U11676 (N_11676,N_11541,N_11408);
xnor U11677 (N_11677,N_11499,N_11482);
and U11678 (N_11678,N_11475,N_11463);
nand U11679 (N_11679,N_11591,N_11590);
nand U11680 (N_11680,N_11432,N_11465);
and U11681 (N_11681,N_11471,N_11517);
nand U11682 (N_11682,N_11419,N_11407);
nor U11683 (N_11683,N_11431,N_11596);
or U11684 (N_11684,N_11451,N_11504);
nand U11685 (N_11685,N_11418,N_11467);
and U11686 (N_11686,N_11510,N_11478);
nor U11687 (N_11687,N_11524,N_11580);
xnor U11688 (N_11688,N_11570,N_11582);
nor U11689 (N_11689,N_11405,N_11480);
nor U11690 (N_11690,N_11409,N_11556);
nor U11691 (N_11691,N_11422,N_11498);
nor U11692 (N_11692,N_11561,N_11413);
or U11693 (N_11693,N_11594,N_11448);
nand U11694 (N_11694,N_11567,N_11587);
or U11695 (N_11695,N_11468,N_11545);
xor U11696 (N_11696,N_11581,N_11543);
xor U11697 (N_11697,N_11569,N_11403);
and U11698 (N_11698,N_11551,N_11542);
xnor U11699 (N_11699,N_11571,N_11559);
nor U11700 (N_11700,N_11550,N_11495);
nand U11701 (N_11701,N_11544,N_11555);
xor U11702 (N_11702,N_11519,N_11593);
nor U11703 (N_11703,N_11539,N_11563);
xor U11704 (N_11704,N_11546,N_11530);
xnor U11705 (N_11705,N_11412,N_11507);
and U11706 (N_11706,N_11490,N_11492);
and U11707 (N_11707,N_11543,N_11425);
nand U11708 (N_11708,N_11511,N_11512);
and U11709 (N_11709,N_11585,N_11469);
xnor U11710 (N_11710,N_11473,N_11596);
xnor U11711 (N_11711,N_11586,N_11470);
xor U11712 (N_11712,N_11594,N_11414);
and U11713 (N_11713,N_11423,N_11519);
nand U11714 (N_11714,N_11528,N_11437);
nand U11715 (N_11715,N_11500,N_11521);
or U11716 (N_11716,N_11526,N_11521);
and U11717 (N_11717,N_11522,N_11477);
and U11718 (N_11718,N_11417,N_11482);
nand U11719 (N_11719,N_11590,N_11569);
or U11720 (N_11720,N_11447,N_11466);
or U11721 (N_11721,N_11473,N_11597);
or U11722 (N_11722,N_11517,N_11433);
nand U11723 (N_11723,N_11580,N_11459);
xor U11724 (N_11724,N_11534,N_11484);
and U11725 (N_11725,N_11412,N_11597);
nor U11726 (N_11726,N_11532,N_11589);
or U11727 (N_11727,N_11483,N_11548);
nand U11728 (N_11728,N_11485,N_11453);
and U11729 (N_11729,N_11440,N_11589);
nand U11730 (N_11730,N_11444,N_11526);
nand U11731 (N_11731,N_11465,N_11544);
or U11732 (N_11732,N_11484,N_11415);
xnor U11733 (N_11733,N_11531,N_11547);
or U11734 (N_11734,N_11549,N_11577);
or U11735 (N_11735,N_11562,N_11594);
or U11736 (N_11736,N_11456,N_11422);
or U11737 (N_11737,N_11521,N_11517);
or U11738 (N_11738,N_11540,N_11531);
xnor U11739 (N_11739,N_11490,N_11403);
nor U11740 (N_11740,N_11523,N_11560);
nor U11741 (N_11741,N_11438,N_11471);
nor U11742 (N_11742,N_11493,N_11441);
xnor U11743 (N_11743,N_11515,N_11565);
xor U11744 (N_11744,N_11486,N_11581);
and U11745 (N_11745,N_11455,N_11443);
xnor U11746 (N_11746,N_11436,N_11520);
or U11747 (N_11747,N_11557,N_11548);
nor U11748 (N_11748,N_11556,N_11517);
xnor U11749 (N_11749,N_11594,N_11420);
nand U11750 (N_11750,N_11448,N_11524);
nand U11751 (N_11751,N_11513,N_11423);
and U11752 (N_11752,N_11579,N_11478);
and U11753 (N_11753,N_11477,N_11517);
xnor U11754 (N_11754,N_11519,N_11588);
nand U11755 (N_11755,N_11581,N_11549);
xnor U11756 (N_11756,N_11549,N_11524);
xor U11757 (N_11757,N_11457,N_11578);
and U11758 (N_11758,N_11488,N_11548);
nand U11759 (N_11759,N_11547,N_11415);
and U11760 (N_11760,N_11423,N_11506);
and U11761 (N_11761,N_11594,N_11421);
xor U11762 (N_11762,N_11497,N_11487);
nor U11763 (N_11763,N_11465,N_11423);
xnor U11764 (N_11764,N_11500,N_11578);
and U11765 (N_11765,N_11511,N_11424);
and U11766 (N_11766,N_11564,N_11466);
nor U11767 (N_11767,N_11431,N_11550);
nand U11768 (N_11768,N_11434,N_11510);
and U11769 (N_11769,N_11593,N_11586);
and U11770 (N_11770,N_11575,N_11429);
xor U11771 (N_11771,N_11408,N_11585);
and U11772 (N_11772,N_11460,N_11514);
xor U11773 (N_11773,N_11463,N_11551);
and U11774 (N_11774,N_11482,N_11584);
xor U11775 (N_11775,N_11502,N_11467);
nor U11776 (N_11776,N_11407,N_11435);
nor U11777 (N_11777,N_11553,N_11489);
and U11778 (N_11778,N_11588,N_11557);
nand U11779 (N_11779,N_11411,N_11530);
or U11780 (N_11780,N_11434,N_11597);
and U11781 (N_11781,N_11561,N_11429);
and U11782 (N_11782,N_11585,N_11556);
xor U11783 (N_11783,N_11539,N_11521);
nand U11784 (N_11784,N_11571,N_11506);
and U11785 (N_11785,N_11539,N_11530);
nand U11786 (N_11786,N_11598,N_11454);
and U11787 (N_11787,N_11458,N_11427);
xor U11788 (N_11788,N_11517,N_11548);
xnor U11789 (N_11789,N_11437,N_11421);
nor U11790 (N_11790,N_11462,N_11541);
xnor U11791 (N_11791,N_11519,N_11479);
nor U11792 (N_11792,N_11582,N_11448);
xnor U11793 (N_11793,N_11523,N_11535);
nor U11794 (N_11794,N_11508,N_11490);
or U11795 (N_11795,N_11541,N_11481);
or U11796 (N_11796,N_11458,N_11430);
and U11797 (N_11797,N_11541,N_11533);
and U11798 (N_11798,N_11538,N_11527);
nand U11799 (N_11799,N_11583,N_11584);
or U11800 (N_11800,N_11693,N_11793);
xor U11801 (N_11801,N_11734,N_11703);
nand U11802 (N_11802,N_11612,N_11662);
nand U11803 (N_11803,N_11692,N_11778);
or U11804 (N_11804,N_11684,N_11614);
nand U11805 (N_11805,N_11783,N_11636);
and U11806 (N_11806,N_11631,N_11604);
xnor U11807 (N_11807,N_11789,N_11770);
nor U11808 (N_11808,N_11787,N_11706);
xor U11809 (N_11809,N_11796,N_11603);
xnor U11810 (N_11810,N_11715,N_11666);
xor U11811 (N_11811,N_11664,N_11731);
nor U11812 (N_11812,N_11690,N_11699);
xnor U11813 (N_11813,N_11738,N_11680);
xnor U11814 (N_11814,N_11654,N_11663);
nor U11815 (N_11815,N_11764,N_11643);
xnor U11816 (N_11816,N_11766,N_11782);
xor U11817 (N_11817,N_11732,N_11687);
nor U11818 (N_11818,N_11630,N_11747);
nor U11819 (N_11819,N_11682,N_11702);
and U11820 (N_11820,N_11704,N_11722);
nand U11821 (N_11821,N_11611,N_11717);
xnor U11822 (N_11822,N_11619,N_11725);
nand U11823 (N_11823,N_11741,N_11613);
xnor U11824 (N_11824,N_11639,N_11674);
or U11825 (N_11825,N_11786,N_11794);
or U11826 (N_11826,N_11656,N_11625);
nor U11827 (N_11827,N_11675,N_11651);
or U11828 (N_11828,N_11697,N_11665);
nand U11829 (N_11829,N_11755,N_11720);
nor U11830 (N_11830,N_11602,N_11605);
or U11831 (N_11831,N_11678,N_11657);
nor U11832 (N_11832,N_11600,N_11608);
nor U11833 (N_11833,N_11773,N_11750);
or U11834 (N_11834,N_11799,N_11660);
nor U11835 (N_11835,N_11781,N_11744);
and U11836 (N_11836,N_11705,N_11632);
and U11837 (N_11837,N_11752,N_11763);
xor U11838 (N_11838,N_11751,N_11689);
nor U11839 (N_11839,N_11695,N_11749);
and U11840 (N_11840,N_11669,N_11616);
nor U11841 (N_11841,N_11670,N_11607);
xnor U11842 (N_11842,N_11694,N_11658);
and U11843 (N_11843,N_11742,N_11685);
nor U11844 (N_11844,N_11661,N_11753);
nand U11845 (N_11845,N_11677,N_11791);
nand U11846 (N_11846,N_11610,N_11679);
xnor U11847 (N_11847,N_11784,N_11647);
and U11848 (N_11848,N_11748,N_11795);
xor U11849 (N_11849,N_11615,N_11667);
or U11850 (N_11850,N_11760,N_11626);
or U11851 (N_11851,N_11645,N_11730);
xor U11852 (N_11852,N_11727,N_11797);
nand U11853 (N_11853,N_11691,N_11698);
nand U11854 (N_11854,N_11790,N_11642);
or U11855 (N_11855,N_11641,N_11757);
nor U11856 (N_11856,N_11671,N_11673);
nand U11857 (N_11857,N_11686,N_11628);
xnor U11858 (N_11858,N_11627,N_11652);
xnor U11859 (N_11859,N_11609,N_11708);
nand U11860 (N_11860,N_11700,N_11739);
and U11861 (N_11861,N_11754,N_11779);
and U11862 (N_11862,N_11785,N_11758);
xnor U11863 (N_11863,N_11775,N_11601);
nor U11864 (N_11864,N_11756,N_11659);
and U11865 (N_11865,N_11712,N_11723);
nor U11866 (N_11866,N_11746,N_11653);
nor U11867 (N_11867,N_11713,N_11634);
xor U11868 (N_11868,N_11728,N_11638);
or U11869 (N_11869,N_11617,N_11618);
nor U11870 (N_11870,N_11629,N_11759);
nand U11871 (N_11871,N_11798,N_11726);
nand U11872 (N_11872,N_11716,N_11709);
and U11873 (N_11873,N_11765,N_11736);
nand U11874 (N_11874,N_11792,N_11633);
nand U11875 (N_11875,N_11606,N_11701);
and U11876 (N_11876,N_11644,N_11710);
xor U11877 (N_11877,N_11762,N_11721);
or U11878 (N_11878,N_11735,N_11780);
xor U11879 (N_11879,N_11621,N_11622);
or U11880 (N_11880,N_11711,N_11637);
or U11881 (N_11881,N_11777,N_11743);
or U11882 (N_11882,N_11688,N_11655);
or U11883 (N_11883,N_11620,N_11676);
and U11884 (N_11884,N_11672,N_11774);
nand U11885 (N_11885,N_11724,N_11624);
nor U11886 (N_11886,N_11646,N_11649);
nor U11887 (N_11887,N_11683,N_11761);
nor U11888 (N_11888,N_11737,N_11740);
nand U11889 (N_11889,N_11788,N_11640);
or U11890 (N_11890,N_11768,N_11733);
nand U11891 (N_11891,N_11776,N_11771);
xnor U11892 (N_11892,N_11707,N_11635);
or U11893 (N_11893,N_11668,N_11772);
or U11894 (N_11894,N_11714,N_11650);
and U11895 (N_11895,N_11696,N_11729);
nand U11896 (N_11896,N_11681,N_11769);
nor U11897 (N_11897,N_11719,N_11745);
nor U11898 (N_11898,N_11718,N_11623);
and U11899 (N_11899,N_11767,N_11648);
xor U11900 (N_11900,N_11768,N_11638);
xnor U11901 (N_11901,N_11647,N_11635);
or U11902 (N_11902,N_11632,N_11643);
xor U11903 (N_11903,N_11695,N_11639);
or U11904 (N_11904,N_11775,N_11773);
nand U11905 (N_11905,N_11681,N_11748);
and U11906 (N_11906,N_11766,N_11733);
and U11907 (N_11907,N_11603,N_11672);
nand U11908 (N_11908,N_11681,N_11772);
or U11909 (N_11909,N_11778,N_11641);
xnor U11910 (N_11910,N_11600,N_11769);
xor U11911 (N_11911,N_11751,N_11714);
nor U11912 (N_11912,N_11781,N_11772);
and U11913 (N_11913,N_11631,N_11761);
or U11914 (N_11914,N_11654,N_11714);
nand U11915 (N_11915,N_11696,N_11647);
nand U11916 (N_11916,N_11612,N_11681);
and U11917 (N_11917,N_11692,N_11762);
and U11918 (N_11918,N_11745,N_11608);
xnor U11919 (N_11919,N_11644,N_11614);
or U11920 (N_11920,N_11613,N_11797);
nor U11921 (N_11921,N_11694,N_11743);
and U11922 (N_11922,N_11732,N_11719);
xor U11923 (N_11923,N_11619,N_11789);
nand U11924 (N_11924,N_11700,N_11683);
or U11925 (N_11925,N_11698,N_11758);
nor U11926 (N_11926,N_11692,N_11611);
and U11927 (N_11927,N_11744,N_11642);
nand U11928 (N_11928,N_11689,N_11655);
nor U11929 (N_11929,N_11696,N_11721);
nand U11930 (N_11930,N_11727,N_11657);
and U11931 (N_11931,N_11704,N_11672);
nor U11932 (N_11932,N_11602,N_11641);
and U11933 (N_11933,N_11695,N_11756);
nor U11934 (N_11934,N_11790,N_11713);
nand U11935 (N_11935,N_11743,N_11625);
xor U11936 (N_11936,N_11628,N_11738);
and U11937 (N_11937,N_11691,N_11788);
nor U11938 (N_11938,N_11613,N_11631);
and U11939 (N_11939,N_11654,N_11613);
nand U11940 (N_11940,N_11731,N_11743);
nand U11941 (N_11941,N_11683,N_11618);
or U11942 (N_11942,N_11705,N_11703);
and U11943 (N_11943,N_11784,N_11658);
nor U11944 (N_11944,N_11626,N_11766);
nand U11945 (N_11945,N_11615,N_11748);
or U11946 (N_11946,N_11744,N_11793);
and U11947 (N_11947,N_11703,N_11792);
or U11948 (N_11948,N_11601,N_11604);
and U11949 (N_11949,N_11720,N_11624);
or U11950 (N_11950,N_11653,N_11706);
and U11951 (N_11951,N_11701,N_11766);
and U11952 (N_11952,N_11698,N_11766);
xor U11953 (N_11953,N_11788,N_11669);
nand U11954 (N_11954,N_11738,N_11607);
nor U11955 (N_11955,N_11767,N_11740);
nor U11956 (N_11956,N_11694,N_11737);
nor U11957 (N_11957,N_11704,N_11780);
xnor U11958 (N_11958,N_11608,N_11721);
nand U11959 (N_11959,N_11662,N_11698);
and U11960 (N_11960,N_11755,N_11745);
nor U11961 (N_11961,N_11602,N_11764);
and U11962 (N_11962,N_11628,N_11709);
nand U11963 (N_11963,N_11664,N_11677);
xor U11964 (N_11964,N_11693,N_11690);
nand U11965 (N_11965,N_11710,N_11716);
and U11966 (N_11966,N_11680,N_11758);
nor U11967 (N_11967,N_11630,N_11631);
or U11968 (N_11968,N_11759,N_11671);
nand U11969 (N_11969,N_11747,N_11623);
nand U11970 (N_11970,N_11742,N_11641);
nand U11971 (N_11971,N_11612,N_11605);
nand U11972 (N_11972,N_11687,N_11767);
or U11973 (N_11973,N_11648,N_11667);
nand U11974 (N_11974,N_11630,N_11663);
nand U11975 (N_11975,N_11687,N_11713);
and U11976 (N_11976,N_11730,N_11610);
nand U11977 (N_11977,N_11779,N_11727);
xnor U11978 (N_11978,N_11702,N_11736);
nor U11979 (N_11979,N_11607,N_11651);
or U11980 (N_11980,N_11663,N_11795);
or U11981 (N_11981,N_11682,N_11737);
nand U11982 (N_11982,N_11678,N_11634);
xnor U11983 (N_11983,N_11628,N_11654);
nand U11984 (N_11984,N_11723,N_11708);
xnor U11985 (N_11985,N_11776,N_11681);
or U11986 (N_11986,N_11789,N_11678);
xor U11987 (N_11987,N_11638,N_11717);
nor U11988 (N_11988,N_11665,N_11668);
nor U11989 (N_11989,N_11710,N_11791);
xnor U11990 (N_11990,N_11637,N_11786);
nand U11991 (N_11991,N_11683,N_11682);
xor U11992 (N_11992,N_11789,N_11615);
nor U11993 (N_11993,N_11634,N_11619);
xnor U11994 (N_11994,N_11669,N_11683);
or U11995 (N_11995,N_11716,N_11797);
nor U11996 (N_11996,N_11687,N_11711);
nand U11997 (N_11997,N_11753,N_11710);
nand U11998 (N_11998,N_11716,N_11759);
and U11999 (N_11999,N_11604,N_11670);
nor U12000 (N_12000,N_11892,N_11988);
and U12001 (N_12001,N_11804,N_11883);
nor U12002 (N_12002,N_11981,N_11935);
and U12003 (N_12003,N_11984,N_11936);
xor U12004 (N_12004,N_11877,N_11932);
nand U12005 (N_12005,N_11905,N_11881);
and U12006 (N_12006,N_11949,N_11852);
nor U12007 (N_12007,N_11944,N_11957);
nand U12008 (N_12008,N_11912,N_11904);
xor U12009 (N_12009,N_11926,N_11867);
nor U12010 (N_12010,N_11911,N_11996);
nor U12011 (N_12011,N_11816,N_11995);
nand U12012 (N_12012,N_11891,N_11895);
nand U12013 (N_12013,N_11923,N_11908);
nor U12014 (N_12014,N_11898,N_11899);
nor U12015 (N_12015,N_11998,N_11990);
and U12016 (N_12016,N_11919,N_11818);
and U12017 (N_12017,N_11977,N_11834);
nor U12018 (N_12018,N_11888,N_11922);
nand U12019 (N_12019,N_11868,N_11863);
nor U12020 (N_12020,N_11817,N_11800);
nand U12021 (N_12021,N_11857,N_11873);
and U12022 (N_12022,N_11856,N_11841);
xnor U12023 (N_12023,N_11808,N_11987);
and U12024 (N_12024,N_11828,N_11897);
nor U12025 (N_12025,N_11963,N_11941);
and U12026 (N_12026,N_11894,N_11801);
nor U12027 (N_12027,N_11827,N_11844);
nand U12028 (N_12028,N_11915,N_11831);
or U12029 (N_12029,N_11961,N_11855);
and U12030 (N_12030,N_11978,N_11833);
xor U12031 (N_12031,N_11874,N_11980);
and U12032 (N_12032,N_11997,N_11962);
nand U12033 (N_12033,N_11930,N_11969);
nor U12034 (N_12034,N_11982,N_11966);
nand U12035 (N_12035,N_11885,N_11979);
and U12036 (N_12036,N_11843,N_11815);
or U12037 (N_12037,N_11989,N_11983);
nand U12038 (N_12038,N_11967,N_11929);
xor U12039 (N_12039,N_11993,N_11976);
xor U12040 (N_12040,N_11921,N_11946);
nand U12041 (N_12041,N_11851,N_11860);
or U12042 (N_12042,N_11906,N_11973);
xor U12043 (N_12043,N_11928,N_11901);
and U12044 (N_12044,N_11965,N_11854);
and U12045 (N_12045,N_11893,N_11947);
and U12046 (N_12046,N_11880,N_11835);
nor U12047 (N_12047,N_11814,N_11959);
and U12048 (N_12048,N_11845,N_11952);
or U12049 (N_12049,N_11848,N_11825);
xor U12050 (N_12050,N_11991,N_11865);
or U12051 (N_12051,N_11927,N_11972);
nor U12052 (N_12052,N_11836,N_11900);
nand U12053 (N_12053,N_11811,N_11824);
or U12054 (N_12054,N_11840,N_11955);
and U12055 (N_12055,N_11925,N_11896);
and U12056 (N_12056,N_11837,N_11846);
xnor U12057 (N_12057,N_11839,N_11830);
nor U12058 (N_12058,N_11806,N_11933);
xor U12059 (N_12059,N_11872,N_11875);
and U12060 (N_12060,N_11968,N_11913);
xor U12061 (N_12061,N_11975,N_11813);
and U12062 (N_12062,N_11950,N_11999);
nand U12063 (N_12063,N_11938,N_11940);
nor U12064 (N_12064,N_11847,N_11934);
nand U12065 (N_12065,N_11903,N_11809);
xnor U12066 (N_12066,N_11850,N_11864);
or U12067 (N_12067,N_11970,N_11876);
and U12068 (N_12068,N_11939,N_11849);
or U12069 (N_12069,N_11826,N_11971);
or U12070 (N_12070,N_11859,N_11819);
nor U12071 (N_12071,N_11884,N_11964);
and U12072 (N_12072,N_11832,N_11887);
xnor U12073 (N_12073,N_11945,N_11916);
nand U12074 (N_12074,N_11994,N_11879);
xnor U12075 (N_12075,N_11910,N_11948);
xnor U12076 (N_12076,N_11951,N_11853);
and U12077 (N_12077,N_11803,N_11943);
nand U12078 (N_12078,N_11861,N_11866);
nand U12079 (N_12079,N_11937,N_11886);
and U12080 (N_12080,N_11931,N_11924);
nand U12081 (N_12081,N_11822,N_11810);
nor U12082 (N_12082,N_11918,N_11942);
nor U12083 (N_12083,N_11871,N_11878);
xnor U12084 (N_12084,N_11838,N_11992);
xnor U12085 (N_12085,N_11870,N_11820);
and U12086 (N_12086,N_11812,N_11842);
and U12087 (N_12087,N_11917,N_11858);
nor U12088 (N_12088,N_11821,N_11823);
nand U12089 (N_12089,N_11986,N_11805);
or U12090 (N_12090,N_11802,N_11807);
nand U12091 (N_12091,N_11954,N_11829);
xor U12092 (N_12092,N_11890,N_11907);
and U12093 (N_12093,N_11914,N_11882);
and U12094 (N_12094,N_11869,N_11889);
nand U12095 (N_12095,N_11909,N_11974);
nand U12096 (N_12096,N_11956,N_11960);
nand U12097 (N_12097,N_11920,N_11902);
nand U12098 (N_12098,N_11985,N_11953);
or U12099 (N_12099,N_11862,N_11958);
or U12100 (N_12100,N_11911,N_11981);
and U12101 (N_12101,N_11907,N_11840);
nor U12102 (N_12102,N_11990,N_11962);
xor U12103 (N_12103,N_11892,N_11963);
or U12104 (N_12104,N_11892,N_11842);
xor U12105 (N_12105,N_11987,N_11968);
xor U12106 (N_12106,N_11841,N_11901);
or U12107 (N_12107,N_11885,N_11821);
nor U12108 (N_12108,N_11955,N_11906);
and U12109 (N_12109,N_11891,N_11932);
and U12110 (N_12110,N_11840,N_11916);
nand U12111 (N_12111,N_11818,N_11917);
or U12112 (N_12112,N_11885,N_11839);
and U12113 (N_12113,N_11824,N_11903);
nand U12114 (N_12114,N_11949,N_11999);
xnor U12115 (N_12115,N_11846,N_11867);
and U12116 (N_12116,N_11973,N_11893);
nand U12117 (N_12117,N_11867,N_11822);
and U12118 (N_12118,N_11919,N_11868);
xnor U12119 (N_12119,N_11833,N_11891);
nand U12120 (N_12120,N_11863,N_11878);
nor U12121 (N_12121,N_11901,N_11934);
or U12122 (N_12122,N_11819,N_11878);
nand U12123 (N_12123,N_11920,N_11955);
nand U12124 (N_12124,N_11900,N_11811);
nor U12125 (N_12125,N_11829,N_11855);
nand U12126 (N_12126,N_11803,N_11832);
or U12127 (N_12127,N_11934,N_11811);
or U12128 (N_12128,N_11843,N_11964);
nor U12129 (N_12129,N_11986,N_11941);
and U12130 (N_12130,N_11918,N_11954);
or U12131 (N_12131,N_11859,N_11920);
or U12132 (N_12132,N_11834,N_11927);
xnor U12133 (N_12133,N_11897,N_11990);
nand U12134 (N_12134,N_11950,N_11940);
nor U12135 (N_12135,N_11892,N_11819);
and U12136 (N_12136,N_11923,N_11978);
nand U12137 (N_12137,N_11924,N_11939);
nor U12138 (N_12138,N_11935,N_11983);
nor U12139 (N_12139,N_11893,N_11951);
nor U12140 (N_12140,N_11950,N_11914);
nand U12141 (N_12141,N_11981,N_11996);
or U12142 (N_12142,N_11961,N_11963);
or U12143 (N_12143,N_11842,N_11856);
xnor U12144 (N_12144,N_11813,N_11888);
nand U12145 (N_12145,N_11815,N_11997);
or U12146 (N_12146,N_11929,N_11886);
nand U12147 (N_12147,N_11893,N_11868);
xnor U12148 (N_12148,N_11954,N_11997);
and U12149 (N_12149,N_11872,N_11908);
and U12150 (N_12150,N_11982,N_11954);
nand U12151 (N_12151,N_11945,N_11941);
xor U12152 (N_12152,N_11850,N_11821);
and U12153 (N_12153,N_11927,N_11998);
nand U12154 (N_12154,N_11881,N_11893);
xnor U12155 (N_12155,N_11921,N_11809);
nor U12156 (N_12156,N_11906,N_11870);
xor U12157 (N_12157,N_11974,N_11817);
xnor U12158 (N_12158,N_11868,N_11860);
and U12159 (N_12159,N_11962,N_11918);
nand U12160 (N_12160,N_11979,N_11965);
nor U12161 (N_12161,N_11849,N_11811);
nor U12162 (N_12162,N_11838,N_11805);
nor U12163 (N_12163,N_11848,N_11872);
or U12164 (N_12164,N_11920,N_11857);
or U12165 (N_12165,N_11997,N_11841);
nor U12166 (N_12166,N_11858,N_11995);
nand U12167 (N_12167,N_11986,N_11972);
nand U12168 (N_12168,N_11986,N_11999);
and U12169 (N_12169,N_11842,N_11954);
nand U12170 (N_12170,N_11868,N_11932);
or U12171 (N_12171,N_11823,N_11949);
and U12172 (N_12172,N_11911,N_11909);
and U12173 (N_12173,N_11844,N_11865);
and U12174 (N_12174,N_11962,N_11897);
xnor U12175 (N_12175,N_11910,N_11923);
nor U12176 (N_12176,N_11965,N_11841);
xor U12177 (N_12177,N_11837,N_11995);
or U12178 (N_12178,N_11918,N_11912);
xor U12179 (N_12179,N_11964,N_11868);
xnor U12180 (N_12180,N_11938,N_11902);
xor U12181 (N_12181,N_11842,N_11923);
or U12182 (N_12182,N_11847,N_11890);
and U12183 (N_12183,N_11890,N_11933);
nand U12184 (N_12184,N_11837,N_11905);
and U12185 (N_12185,N_11862,N_11951);
or U12186 (N_12186,N_11938,N_11836);
nor U12187 (N_12187,N_11805,N_11890);
xnor U12188 (N_12188,N_11973,N_11927);
or U12189 (N_12189,N_11934,N_11959);
nor U12190 (N_12190,N_11831,N_11948);
and U12191 (N_12191,N_11984,N_11999);
and U12192 (N_12192,N_11810,N_11912);
nor U12193 (N_12193,N_11909,N_11821);
xor U12194 (N_12194,N_11993,N_11847);
or U12195 (N_12195,N_11816,N_11894);
or U12196 (N_12196,N_11847,N_11800);
nor U12197 (N_12197,N_11906,N_11884);
or U12198 (N_12198,N_11976,N_11887);
or U12199 (N_12199,N_11835,N_11924);
nand U12200 (N_12200,N_12127,N_12096);
nor U12201 (N_12201,N_12187,N_12102);
or U12202 (N_12202,N_12014,N_12010);
nor U12203 (N_12203,N_12180,N_12181);
nor U12204 (N_12204,N_12171,N_12122);
nor U12205 (N_12205,N_12182,N_12111);
nand U12206 (N_12206,N_12052,N_12189);
nor U12207 (N_12207,N_12045,N_12057);
or U12208 (N_12208,N_12169,N_12114);
and U12209 (N_12209,N_12011,N_12038);
nand U12210 (N_12210,N_12063,N_12143);
or U12211 (N_12211,N_12138,N_12026);
and U12212 (N_12212,N_12093,N_12148);
nor U12213 (N_12213,N_12040,N_12046);
xnor U12214 (N_12214,N_12083,N_12059);
and U12215 (N_12215,N_12147,N_12061);
xnor U12216 (N_12216,N_12174,N_12141);
nor U12217 (N_12217,N_12088,N_12132);
nand U12218 (N_12218,N_12185,N_12198);
or U12219 (N_12219,N_12023,N_12135);
nor U12220 (N_12220,N_12144,N_12116);
nor U12221 (N_12221,N_12123,N_12074);
nand U12222 (N_12222,N_12033,N_12016);
xnor U12223 (N_12223,N_12175,N_12107);
or U12224 (N_12224,N_12024,N_12190);
or U12225 (N_12225,N_12034,N_12145);
xnor U12226 (N_12226,N_12048,N_12015);
and U12227 (N_12227,N_12091,N_12159);
or U12228 (N_12228,N_12177,N_12100);
nor U12229 (N_12229,N_12153,N_12099);
or U12230 (N_12230,N_12192,N_12004);
or U12231 (N_12231,N_12095,N_12080);
nand U12232 (N_12232,N_12070,N_12071);
nor U12233 (N_12233,N_12008,N_12075);
nand U12234 (N_12234,N_12161,N_12151);
nand U12235 (N_12235,N_12136,N_12030);
and U12236 (N_12236,N_12155,N_12082);
and U12237 (N_12237,N_12098,N_12196);
xor U12238 (N_12238,N_12109,N_12117);
and U12239 (N_12239,N_12101,N_12021);
nand U12240 (N_12240,N_12113,N_12009);
nand U12241 (N_12241,N_12115,N_12125);
nor U12242 (N_12242,N_12168,N_12025);
and U12243 (N_12243,N_12158,N_12022);
and U12244 (N_12244,N_12133,N_12178);
and U12245 (N_12245,N_12050,N_12112);
xnor U12246 (N_12246,N_12058,N_12197);
and U12247 (N_12247,N_12103,N_12126);
nand U12248 (N_12248,N_12186,N_12129);
xnor U12249 (N_12249,N_12157,N_12184);
nor U12250 (N_12250,N_12094,N_12118);
nor U12251 (N_12251,N_12188,N_12119);
and U12252 (N_12252,N_12137,N_12139);
or U12253 (N_12253,N_12064,N_12162);
nand U12254 (N_12254,N_12037,N_12003);
xor U12255 (N_12255,N_12041,N_12069);
or U12256 (N_12256,N_12146,N_12056);
xnor U12257 (N_12257,N_12134,N_12049);
or U12258 (N_12258,N_12047,N_12065);
and U12259 (N_12259,N_12036,N_12097);
or U12260 (N_12260,N_12160,N_12154);
and U12261 (N_12261,N_12077,N_12121);
nor U12262 (N_12262,N_12104,N_12042);
xnor U12263 (N_12263,N_12044,N_12110);
and U12264 (N_12264,N_12076,N_12013);
xnor U12265 (N_12265,N_12128,N_12020);
or U12266 (N_12266,N_12173,N_12150);
and U12267 (N_12267,N_12005,N_12032);
and U12268 (N_12268,N_12176,N_12092);
and U12269 (N_12269,N_12152,N_12028);
nand U12270 (N_12270,N_12199,N_12130);
or U12271 (N_12271,N_12131,N_12170);
and U12272 (N_12272,N_12124,N_12001);
and U12273 (N_12273,N_12039,N_12000);
xor U12274 (N_12274,N_12019,N_12090);
xnor U12275 (N_12275,N_12167,N_12191);
xor U12276 (N_12276,N_12084,N_12120);
and U12277 (N_12277,N_12018,N_12164);
and U12278 (N_12278,N_12054,N_12142);
nor U12279 (N_12279,N_12140,N_12073);
and U12280 (N_12280,N_12031,N_12060);
nor U12281 (N_12281,N_12106,N_12086);
and U12282 (N_12282,N_12165,N_12029);
and U12283 (N_12283,N_12072,N_12085);
nor U12284 (N_12284,N_12194,N_12163);
xor U12285 (N_12285,N_12012,N_12183);
nor U12286 (N_12286,N_12067,N_12053);
or U12287 (N_12287,N_12156,N_12062);
xnor U12288 (N_12288,N_12149,N_12068);
nor U12289 (N_12289,N_12089,N_12035);
and U12290 (N_12290,N_12172,N_12017);
xnor U12291 (N_12291,N_12078,N_12007);
nor U12292 (N_12292,N_12081,N_12195);
nand U12293 (N_12293,N_12027,N_12087);
or U12294 (N_12294,N_12193,N_12055);
and U12295 (N_12295,N_12105,N_12108);
nor U12296 (N_12296,N_12006,N_12079);
or U12297 (N_12297,N_12043,N_12002);
or U12298 (N_12298,N_12051,N_12179);
nor U12299 (N_12299,N_12066,N_12166);
or U12300 (N_12300,N_12006,N_12053);
nor U12301 (N_12301,N_12120,N_12092);
nand U12302 (N_12302,N_12184,N_12117);
or U12303 (N_12303,N_12097,N_12008);
xor U12304 (N_12304,N_12016,N_12111);
and U12305 (N_12305,N_12101,N_12039);
xor U12306 (N_12306,N_12062,N_12107);
or U12307 (N_12307,N_12166,N_12125);
xor U12308 (N_12308,N_12040,N_12088);
xnor U12309 (N_12309,N_12134,N_12030);
nand U12310 (N_12310,N_12111,N_12028);
or U12311 (N_12311,N_12087,N_12050);
and U12312 (N_12312,N_12120,N_12059);
nand U12313 (N_12313,N_12064,N_12180);
nor U12314 (N_12314,N_12087,N_12036);
nand U12315 (N_12315,N_12028,N_12191);
nand U12316 (N_12316,N_12014,N_12012);
and U12317 (N_12317,N_12038,N_12043);
or U12318 (N_12318,N_12112,N_12086);
xor U12319 (N_12319,N_12093,N_12197);
xnor U12320 (N_12320,N_12097,N_12112);
and U12321 (N_12321,N_12048,N_12042);
nor U12322 (N_12322,N_12075,N_12151);
nand U12323 (N_12323,N_12102,N_12018);
nor U12324 (N_12324,N_12009,N_12002);
xnor U12325 (N_12325,N_12178,N_12115);
xor U12326 (N_12326,N_12134,N_12007);
nor U12327 (N_12327,N_12055,N_12107);
nor U12328 (N_12328,N_12009,N_12104);
nor U12329 (N_12329,N_12174,N_12164);
nor U12330 (N_12330,N_12177,N_12096);
or U12331 (N_12331,N_12152,N_12045);
xnor U12332 (N_12332,N_12066,N_12016);
and U12333 (N_12333,N_12131,N_12049);
nand U12334 (N_12334,N_12007,N_12194);
or U12335 (N_12335,N_12053,N_12002);
xor U12336 (N_12336,N_12113,N_12003);
nor U12337 (N_12337,N_12171,N_12142);
or U12338 (N_12338,N_12099,N_12169);
and U12339 (N_12339,N_12040,N_12183);
and U12340 (N_12340,N_12013,N_12143);
xor U12341 (N_12341,N_12044,N_12189);
xor U12342 (N_12342,N_12079,N_12171);
or U12343 (N_12343,N_12140,N_12110);
nand U12344 (N_12344,N_12081,N_12097);
or U12345 (N_12345,N_12174,N_12027);
nand U12346 (N_12346,N_12034,N_12043);
nor U12347 (N_12347,N_12060,N_12004);
or U12348 (N_12348,N_12196,N_12065);
nor U12349 (N_12349,N_12001,N_12155);
and U12350 (N_12350,N_12001,N_12086);
xnor U12351 (N_12351,N_12103,N_12134);
or U12352 (N_12352,N_12067,N_12059);
or U12353 (N_12353,N_12097,N_12177);
nand U12354 (N_12354,N_12158,N_12048);
nor U12355 (N_12355,N_12022,N_12163);
nor U12356 (N_12356,N_12158,N_12108);
xor U12357 (N_12357,N_12006,N_12189);
or U12358 (N_12358,N_12117,N_12195);
nand U12359 (N_12359,N_12182,N_12134);
and U12360 (N_12360,N_12173,N_12062);
xnor U12361 (N_12361,N_12086,N_12182);
and U12362 (N_12362,N_12079,N_12017);
nand U12363 (N_12363,N_12184,N_12030);
xnor U12364 (N_12364,N_12136,N_12145);
xnor U12365 (N_12365,N_12048,N_12070);
nand U12366 (N_12366,N_12154,N_12042);
nor U12367 (N_12367,N_12028,N_12034);
and U12368 (N_12368,N_12099,N_12061);
and U12369 (N_12369,N_12075,N_12066);
and U12370 (N_12370,N_12006,N_12073);
nand U12371 (N_12371,N_12065,N_12164);
xor U12372 (N_12372,N_12123,N_12102);
nor U12373 (N_12373,N_12043,N_12051);
or U12374 (N_12374,N_12048,N_12104);
or U12375 (N_12375,N_12027,N_12172);
nor U12376 (N_12376,N_12002,N_12079);
and U12377 (N_12377,N_12026,N_12074);
and U12378 (N_12378,N_12142,N_12083);
nor U12379 (N_12379,N_12194,N_12199);
xor U12380 (N_12380,N_12111,N_12136);
nand U12381 (N_12381,N_12108,N_12056);
nor U12382 (N_12382,N_12129,N_12085);
nor U12383 (N_12383,N_12006,N_12099);
nor U12384 (N_12384,N_12095,N_12063);
xor U12385 (N_12385,N_12048,N_12188);
nand U12386 (N_12386,N_12105,N_12017);
and U12387 (N_12387,N_12013,N_12094);
xor U12388 (N_12388,N_12035,N_12024);
and U12389 (N_12389,N_12168,N_12148);
nor U12390 (N_12390,N_12150,N_12169);
xnor U12391 (N_12391,N_12195,N_12000);
or U12392 (N_12392,N_12072,N_12069);
nor U12393 (N_12393,N_12154,N_12048);
and U12394 (N_12394,N_12174,N_12186);
and U12395 (N_12395,N_12112,N_12103);
xor U12396 (N_12396,N_12090,N_12198);
and U12397 (N_12397,N_12102,N_12155);
and U12398 (N_12398,N_12085,N_12150);
nor U12399 (N_12399,N_12088,N_12053);
and U12400 (N_12400,N_12396,N_12327);
or U12401 (N_12401,N_12306,N_12208);
nor U12402 (N_12402,N_12316,N_12266);
or U12403 (N_12403,N_12295,N_12210);
or U12404 (N_12404,N_12382,N_12322);
xnor U12405 (N_12405,N_12323,N_12380);
xor U12406 (N_12406,N_12320,N_12237);
and U12407 (N_12407,N_12212,N_12244);
nand U12408 (N_12408,N_12361,N_12368);
nor U12409 (N_12409,N_12261,N_12225);
nor U12410 (N_12410,N_12254,N_12315);
and U12411 (N_12411,N_12355,N_12317);
nand U12412 (N_12412,N_12302,N_12387);
or U12413 (N_12413,N_12239,N_12277);
nand U12414 (N_12414,N_12330,N_12228);
nor U12415 (N_12415,N_12227,N_12359);
or U12416 (N_12416,N_12399,N_12293);
nor U12417 (N_12417,N_12236,N_12220);
and U12418 (N_12418,N_12264,N_12260);
and U12419 (N_12419,N_12258,N_12319);
xnor U12420 (N_12420,N_12267,N_12245);
and U12421 (N_12421,N_12299,N_12204);
xor U12422 (N_12422,N_12218,N_12341);
nand U12423 (N_12423,N_12231,N_12386);
and U12424 (N_12424,N_12262,N_12308);
or U12425 (N_12425,N_12346,N_12242);
nor U12426 (N_12426,N_12339,N_12335);
nand U12427 (N_12427,N_12280,N_12348);
nor U12428 (N_12428,N_12366,N_12294);
nor U12429 (N_12429,N_12363,N_12255);
and U12430 (N_12430,N_12219,N_12376);
xnor U12431 (N_12431,N_12336,N_12373);
and U12432 (N_12432,N_12350,N_12342);
or U12433 (N_12433,N_12321,N_12329);
xnor U12434 (N_12434,N_12392,N_12291);
or U12435 (N_12435,N_12226,N_12233);
nand U12436 (N_12436,N_12313,N_12290);
and U12437 (N_12437,N_12309,N_12285);
nor U12438 (N_12438,N_12334,N_12272);
xor U12439 (N_12439,N_12287,N_12360);
nand U12440 (N_12440,N_12305,N_12282);
nor U12441 (N_12441,N_12249,N_12243);
xnor U12442 (N_12442,N_12263,N_12352);
and U12443 (N_12443,N_12222,N_12358);
or U12444 (N_12444,N_12256,N_12331);
or U12445 (N_12445,N_12279,N_12338);
nand U12446 (N_12446,N_12215,N_12388);
or U12447 (N_12447,N_12292,N_12296);
or U12448 (N_12448,N_12246,N_12398);
or U12449 (N_12449,N_12304,N_12201);
nand U12450 (N_12450,N_12397,N_12247);
nor U12451 (N_12451,N_12209,N_12269);
nor U12452 (N_12452,N_12377,N_12213);
and U12453 (N_12453,N_12325,N_12365);
xor U12454 (N_12454,N_12383,N_12297);
and U12455 (N_12455,N_12337,N_12351);
xnor U12456 (N_12456,N_12253,N_12389);
nor U12457 (N_12457,N_12318,N_12265);
xnor U12458 (N_12458,N_12314,N_12284);
xnor U12459 (N_12459,N_12340,N_12372);
and U12460 (N_12460,N_12235,N_12207);
and U12461 (N_12461,N_12238,N_12278);
or U12462 (N_12462,N_12324,N_12206);
and U12463 (N_12463,N_12353,N_12328);
nor U12464 (N_12464,N_12385,N_12369);
and U12465 (N_12465,N_12300,N_12364);
nor U12466 (N_12466,N_12307,N_12230);
and U12467 (N_12467,N_12223,N_12333);
and U12468 (N_12468,N_12283,N_12381);
nor U12469 (N_12469,N_12273,N_12343);
or U12470 (N_12470,N_12203,N_12374);
nor U12471 (N_12471,N_12221,N_12390);
xor U12472 (N_12472,N_12232,N_12384);
nand U12473 (N_12473,N_12375,N_12240);
nand U12474 (N_12474,N_12301,N_12391);
xor U12475 (N_12475,N_12362,N_12281);
nor U12476 (N_12476,N_12241,N_12354);
nor U12477 (N_12477,N_12257,N_12248);
nand U12478 (N_12478,N_12216,N_12393);
nand U12479 (N_12479,N_12276,N_12250);
nand U12480 (N_12480,N_12252,N_12379);
nor U12481 (N_12481,N_12251,N_12344);
or U12482 (N_12482,N_12395,N_12349);
or U12483 (N_12483,N_12289,N_12347);
xor U12484 (N_12484,N_12332,N_12312);
or U12485 (N_12485,N_12274,N_12370);
or U12486 (N_12486,N_12229,N_12214);
nand U12487 (N_12487,N_12356,N_12394);
xor U12488 (N_12488,N_12378,N_12367);
and U12489 (N_12489,N_12270,N_12202);
nand U12490 (N_12490,N_12311,N_12217);
nor U12491 (N_12491,N_12224,N_12259);
xor U12492 (N_12492,N_12345,N_12211);
nand U12493 (N_12493,N_12200,N_12275);
nand U12494 (N_12494,N_12268,N_12303);
nand U12495 (N_12495,N_12205,N_12271);
and U12496 (N_12496,N_12234,N_12286);
or U12497 (N_12497,N_12357,N_12310);
and U12498 (N_12498,N_12326,N_12298);
nand U12499 (N_12499,N_12288,N_12371);
nand U12500 (N_12500,N_12273,N_12303);
and U12501 (N_12501,N_12290,N_12385);
and U12502 (N_12502,N_12354,N_12358);
nor U12503 (N_12503,N_12207,N_12331);
or U12504 (N_12504,N_12334,N_12296);
or U12505 (N_12505,N_12328,N_12376);
xor U12506 (N_12506,N_12399,N_12262);
nor U12507 (N_12507,N_12291,N_12312);
and U12508 (N_12508,N_12282,N_12307);
nor U12509 (N_12509,N_12291,N_12297);
xnor U12510 (N_12510,N_12399,N_12239);
or U12511 (N_12511,N_12226,N_12356);
and U12512 (N_12512,N_12273,N_12244);
or U12513 (N_12513,N_12338,N_12332);
and U12514 (N_12514,N_12324,N_12208);
nand U12515 (N_12515,N_12259,N_12263);
or U12516 (N_12516,N_12281,N_12317);
xnor U12517 (N_12517,N_12313,N_12234);
nor U12518 (N_12518,N_12212,N_12245);
or U12519 (N_12519,N_12208,N_12289);
or U12520 (N_12520,N_12245,N_12273);
nand U12521 (N_12521,N_12213,N_12274);
nor U12522 (N_12522,N_12386,N_12239);
nor U12523 (N_12523,N_12214,N_12362);
nand U12524 (N_12524,N_12266,N_12374);
nand U12525 (N_12525,N_12252,N_12334);
nand U12526 (N_12526,N_12210,N_12219);
xor U12527 (N_12527,N_12280,N_12241);
xor U12528 (N_12528,N_12226,N_12330);
nand U12529 (N_12529,N_12238,N_12312);
nor U12530 (N_12530,N_12297,N_12216);
nor U12531 (N_12531,N_12289,N_12204);
and U12532 (N_12532,N_12373,N_12222);
or U12533 (N_12533,N_12382,N_12264);
nor U12534 (N_12534,N_12284,N_12303);
or U12535 (N_12535,N_12329,N_12237);
and U12536 (N_12536,N_12257,N_12381);
nand U12537 (N_12537,N_12295,N_12342);
nand U12538 (N_12538,N_12355,N_12288);
xnor U12539 (N_12539,N_12366,N_12242);
and U12540 (N_12540,N_12371,N_12241);
nand U12541 (N_12541,N_12231,N_12352);
or U12542 (N_12542,N_12235,N_12323);
xnor U12543 (N_12543,N_12240,N_12360);
xnor U12544 (N_12544,N_12277,N_12270);
xnor U12545 (N_12545,N_12300,N_12261);
nand U12546 (N_12546,N_12232,N_12347);
xor U12547 (N_12547,N_12340,N_12247);
and U12548 (N_12548,N_12223,N_12388);
nand U12549 (N_12549,N_12384,N_12327);
nand U12550 (N_12550,N_12245,N_12316);
xor U12551 (N_12551,N_12267,N_12274);
and U12552 (N_12552,N_12390,N_12215);
nand U12553 (N_12553,N_12284,N_12392);
nand U12554 (N_12554,N_12310,N_12393);
nand U12555 (N_12555,N_12237,N_12255);
xnor U12556 (N_12556,N_12326,N_12394);
and U12557 (N_12557,N_12312,N_12232);
or U12558 (N_12558,N_12308,N_12224);
nor U12559 (N_12559,N_12337,N_12291);
and U12560 (N_12560,N_12235,N_12371);
or U12561 (N_12561,N_12274,N_12310);
xnor U12562 (N_12562,N_12219,N_12322);
and U12563 (N_12563,N_12265,N_12200);
xor U12564 (N_12564,N_12328,N_12214);
nand U12565 (N_12565,N_12262,N_12367);
nor U12566 (N_12566,N_12372,N_12371);
or U12567 (N_12567,N_12379,N_12257);
or U12568 (N_12568,N_12254,N_12332);
and U12569 (N_12569,N_12347,N_12375);
nand U12570 (N_12570,N_12203,N_12318);
and U12571 (N_12571,N_12270,N_12218);
nor U12572 (N_12572,N_12238,N_12333);
nor U12573 (N_12573,N_12323,N_12300);
nor U12574 (N_12574,N_12316,N_12270);
or U12575 (N_12575,N_12393,N_12345);
nand U12576 (N_12576,N_12254,N_12223);
or U12577 (N_12577,N_12395,N_12371);
or U12578 (N_12578,N_12229,N_12281);
nor U12579 (N_12579,N_12218,N_12316);
nor U12580 (N_12580,N_12205,N_12294);
nand U12581 (N_12581,N_12289,N_12227);
xnor U12582 (N_12582,N_12380,N_12355);
or U12583 (N_12583,N_12377,N_12295);
nand U12584 (N_12584,N_12332,N_12253);
xnor U12585 (N_12585,N_12205,N_12360);
nor U12586 (N_12586,N_12215,N_12394);
and U12587 (N_12587,N_12338,N_12379);
nor U12588 (N_12588,N_12332,N_12229);
nand U12589 (N_12589,N_12322,N_12300);
and U12590 (N_12590,N_12363,N_12242);
nor U12591 (N_12591,N_12236,N_12256);
or U12592 (N_12592,N_12245,N_12284);
nand U12593 (N_12593,N_12297,N_12337);
nand U12594 (N_12594,N_12357,N_12317);
nor U12595 (N_12595,N_12339,N_12212);
or U12596 (N_12596,N_12338,N_12343);
nor U12597 (N_12597,N_12258,N_12243);
and U12598 (N_12598,N_12303,N_12339);
nand U12599 (N_12599,N_12285,N_12284);
or U12600 (N_12600,N_12509,N_12416);
xor U12601 (N_12601,N_12442,N_12516);
or U12602 (N_12602,N_12544,N_12533);
xnor U12603 (N_12603,N_12422,N_12582);
nand U12604 (N_12604,N_12530,N_12431);
or U12605 (N_12605,N_12504,N_12502);
nand U12606 (N_12606,N_12572,N_12465);
xor U12607 (N_12607,N_12491,N_12469);
or U12608 (N_12608,N_12593,N_12458);
nand U12609 (N_12609,N_12576,N_12577);
nand U12610 (N_12610,N_12404,N_12550);
xor U12611 (N_12611,N_12559,N_12457);
xnor U12612 (N_12612,N_12566,N_12489);
nand U12613 (N_12613,N_12432,N_12476);
nand U12614 (N_12614,N_12448,N_12427);
or U12615 (N_12615,N_12505,N_12420);
or U12616 (N_12616,N_12587,N_12490);
nand U12617 (N_12617,N_12400,N_12532);
xor U12618 (N_12618,N_12554,N_12595);
and U12619 (N_12619,N_12545,N_12537);
nand U12620 (N_12620,N_12513,N_12562);
nand U12621 (N_12621,N_12534,N_12402);
or U12622 (N_12622,N_12531,N_12588);
xnor U12623 (N_12623,N_12438,N_12548);
nand U12624 (N_12624,N_12487,N_12565);
xnor U12625 (N_12625,N_12467,N_12441);
and U12626 (N_12626,N_12472,N_12540);
nor U12627 (N_12627,N_12558,N_12560);
nor U12628 (N_12628,N_12453,N_12542);
and U12629 (N_12629,N_12419,N_12498);
or U12630 (N_12630,N_12519,N_12564);
nand U12631 (N_12631,N_12521,N_12483);
xor U12632 (N_12632,N_12401,N_12573);
nand U12633 (N_12633,N_12506,N_12415);
xor U12634 (N_12634,N_12464,N_12597);
nand U12635 (N_12635,N_12446,N_12547);
or U12636 (N_12636,N_12439,N_12523);
and U12637 (N_12637,N_12556,N_12541);
and U12638 (N_12638,N_12425,N_12455);
or U12639 (N_12639,N_12484,N_12557);
or U12640 (N_12640,N_12575,N_12526);
xor U12641 (N_12641,N_12407,N_12580);
nor U12642 (N_12642,N_12410,N_12473);
and U12643 (N_12643,N_12440,N_12459);
nor U12644 (N_12644,N_12585,N_12578);
xor U12645 (N_12645,N_12447,N_12510);
nand U12646 (N_12646,N_12429,N_12437);
xnor U12647 (N_12647,N_12475,N_12503);
nand U12648 (N_12648,N_12553,N_12546);
nor U12649 (N_12649,N_12418,N_12571);
nand U12650 (N_12650,N_12555,N_12549);
xor U12651 (N_12651,N_12449,N_12408);
nand U12652 (N_12652,N_12406,N_12461);
and U12653 (N_12653,N_12488,N_12596);
or U12654 (N_12654,N_12598,N_12589);
nand U12655 (N_12655,N_12450,N_12403);
or U12656 (N_12656,N_12591,N_12581);
and U12657 (N_12657,N_12535,N_12567);
or U12658 (N_12658,N_12486,N_12413);
xnor U12659 (N_12659,N_12500,N_12501);
xnor U12660 (N_12660,N_12417,N_12590);
and U12661 (N_12661,N_12433,N_12574);
nor U12662 (N_12662,N_12552,N_12468);
and U12663 (N_12663,N_12569,N_12543);
nand U12664 (N_12664,N_12480,N_12493);
nand U12665 (N_12665,N_12494,N_12485);
nor U12666 (N_12666,N_12568,N_12583);
and U12667 (N_12667,N_12527,N_12470);
xnor U12668 (N_12668,N_12463,N_12462);
nand U12669 (N_12669,N_12518,N_12508);
and U12670 (N_12670,N_12460,N_12405);
nand U12671 (N_12671,N_12525,N_12421);
or U12672 (N_12672,N_12563,N_12599);
nor U12673 (N_12673,N_12561,N_12512);
nand U12674 (N_12674,N_12496,N_12495);
or U12675 (N_12675,N_12514,N_12570);
or U12676 (N_12676,N_12497,N_12443);
xor U12677 (N_12677,N_12436,N_12538);
or U12678 (N_12678,N_12499,N_12430);
nand U12679 (N_12679,N_12409,N_12492);
nand U12680 (N_12680,N_12529,N_12444);
or U12681 (N_12681,N_12423,N_12594);
and U12682 (N_12682,N_12435,N_12586);
xnor U12683 (N_12683,N_12454,N_12445);
nand U12684 (N_12684,N_12528,N_12517);
xor U12685 (N_12685,N_12456,N_12536);
nand U12686 (N_12686,N_12539,N_12511);
or U12687 (N_12687,N_12579,N_12584);
xor U12688 (N_12688,N_12507,N_12434);
nor U12689 (N_12689,N_12452,N_12524);
or U12690 (N_12690,N_12412,N_12482);
xor U12691 (N_12691,N_12466,N_12515);
nor U12692 (N_12692,N_12478,N_12481);
nand U12693 (N_12693,N_12471,N_12474);
or U12694 (N_12694,N_12520,N_12551);
nand U12695 (N_12695,N_12479,N_12477);
xnor U12696 (N_12696,N_12411,N_12426);
xnor U12697 (N_12697,N_12522,N_12414);
xor U12698 (N_12698,N_12424,N_12451);
and U12699 (N_12699,N_12592,N_12428);
nor U12700 (N_12700,N_12401,N_12524);
nand U12701 (N_12701,N_12592,N_12403);
xnor U12702 (N_12702,N_12459,N_12539);
nand U12703 (N_12703,N_12454,N_12578);
or U12704 (N_12704,N_12526,N_12412);
or U12705 (N_12705,N_12427,N_12460);
and U12706 (N_12706,N_12499,N_12401);
nor U12707 (N_12707,N_12522,N_12442);
and U12708 (N_12708,N_12437,N_12528);
or U12709 (N_12709,N_12537,N_12474);
and U12710 (N_12710,N_12522,N_12571);
xor U12711 (N_12711,N_12563,N_12578);
xor U12712 (N_12712,N_12432,N_12538);
and U12713 (N_12713,N_12494,N_12553);
xor U12714 (N_12714,N_12442,N_12571);
and U12715 (N_12715,N_12475,N_12528);
nand U12716 (N_12716,N_12477,N_12426);
nor U12717 (N_12717,N_12437,N_12408);
nand U12718 (N_12718,N_12560,N_12583);
and U12719 (N_12719,N_12459,N_12491);
or U12720 (N_12720,N_12518,N_12490);
xnor U12721 (N_12721,N_12552,N_12529);
or U12722 (N_12722,N_12483,N_12550);
and U12723 (N_12723,N_12412,N_12465);
and U12724 (N_12724,N_12482,N_12497);
and U12725 (N_12725,N_12548,N_12449);
or U12726 (N_12726,N_12445,N_12568);
xor U12727 (N_12727,N_12515,N_12568);
nand U12728 (N_12728,N_12428,N_12469);
nor U12729 (N_12729,N_12595,N_12566);
xnor U12730 (N_12730,N_12489,N_12596);
nor U12731 (N_12731,N_12571,N_12445);
or U12732 (N_12732,N_12417,N_12517);
nor U12733 (N_12733,N_12545,N_12571);
nor U12734 (N_12734,N_12556,N_12448);
and U12735 (N_12735,N_12518,N_12538);
nor U12736 (N_12736,N_12590,N_12421);
nand U12737 (N_12737,N_12441,N_12484);
nand U12738 (N_12738,N_12555,N_12598);
nand U12739 (N_12739,N_12431,N_12579);
nand U12740 (N_12740,N_12478,N_12564);
nand U12741 (N_12741,N_12451,N_12430);
nor U12742 (N_12742,N_12465,N_12476);
xor U12743 (N_12743,N_12497,N_12544);
nor U12744 (N_12744,N_12579,N_12515);
xor U12745 (N_12745,N_12526,N_12490);
and U12746 (N_12746,N_12512,N_12454);
or U12747 (N_12747,N_12531,N_12560);
nor U12748 (N_12748,N_12424,N_12592);
nand U12749 (N_12749,N_12579,N_12418);
xor U12750 (N_12750,N_12571,N_12518);
and U12751 (N_12751,N_12568,N_12547);
or U12752 (N_12752,N_12436,N_12577);
or U12753 (N_12753,N_12443,N_12523);
nor U12754 (N_12754,N_12509,N_12445);
and U12755 (N_12755,N_12514,N_12452);
xor U12756 (N_12756,N_12527,N_12434);
nor U12757 (N_12757,N_12421,N_12584);
nor U12758 (N_12758,N_12501,N_12422);
nand U12759 (N_12759,N_12433,N_12500);
nand U12760 (N_12760,N_12569,N_12451);
xnor U12761 (N_12761,N_12434,N_12531);
nor U12762 (N_12762,N_12445,N_12407);
or U12763 (N_12763,N_12580,N_12562);
or U12764 (N_12764,N_12434,N_12447);
or U12765 (N_12765,N_12496,N_12576);
nand U12766 (N_12766,N_12529,N_12598);
xnor U12767 (N_12767,N_12589,N_12532);
or U12768 (N_12768,N_12592,N_12554);
and U12769 (N_12769,N_12576,N_12592);
nand U12770 (N_12770,N_12503,N_12489);
nor U12771 (N_12771,N_12461,N_12464);
nand U12772 (N_12772,N_12450,N_12585);
or U12773 (N_12773,N_12421,N_12570);
or U12774 (N_12774,N_12551,N_12594);
or U12775 (N_12775,N_12596,N_12479);
xor U12776 (N_12776,N_12497,N_12501);
nor U12777 (N_12777,N_12587,N_12575);
nand U12778 (N_12778,N_12409,N_12468);
nand U12779 (N_12779,N_12516,N_12476);
or U12780 (N_12780,N_12587,N_12472);
xnor U12781 (N_12781,N_12563,N_12467);
and U12782 (N_12782,N_12444,N_12539);
xor U12783 (N_12783,N_12538,N_12566);
xnor U12784 (N_12784,N_12567,N_12463);
xnor U12785 (N_12785,N_12479,N_12537);
nand U12786 (N_12786,N_12593,N_12589);
nand U12787 (N_12787,N_12512,N_12589);
xnor U12788 (N_12788,N_12422,N_12423);
nor U12789 (N_12789,N_12526,N_12430);
xor U12790 (N_12790,N_12494,N_12503);
nor U12791 (N_12791,N_12497,N_12572);
nor U12792 (N_12792,N_12407,N_12409);
and U12793 (N_12793,N_12598,N_12458);
and U12794 (N_12794,N_12539,N_12493);
and U12795 (N_12795,N_12445,N_12547);
xnor U12796 (N_12796,N_12518,N_12444);
nand U12797 (N_12797,N_12445,N_12455);
and U12798 (N_12798,N_12539,N_12577);
xor U12799 (N_12799,N_12418,N_12439);
and U12800 (N_12800,N_12626,N_12709);
and U12801 (N_12801,N_12720,N_12685);
or U12802 (N_12802,N_12789,N_12634);
xnor U12803 (N_12803,N_12691,N_12764);
nand U12804 (N_12804,N_12786,N_12675);
and U12805 (N_12805,N_12784,N_12790);
xor U12806 (N_12806,N_12735,N_12729);
xnor U12807 (N_12807,N_12683,N_12762);
nand U12808 (N_12808,N_12736,N_12678);
or U12809 (N_12809,N_12738,N_12665);
nor U12810 (N_12810,N_12639,N_12796);
or U12811 (N_12811,N_12636,N_12616);
nand U12812 (N_12812,N_12797,N_12760);
or U12813 (N_12813,N_12656,N_12765);
nor U12814 (N_12814,N_12682,N_12755);
xor U12815 (N_12815,N_12715,N_12707);
nor U12816 (N_12816,N_12652,N_12633);
xor U12817 (N_12817,N_12651,N_12669);
xor U12818 (N_12818,N_12601,N_12664);
xnor U12819 (N_12819,N_12772,N_12611);
xnor U12820 (N_12820,N_12774,N_12734);
nand U12821 (N_12821,N_12702,N_12731);
xnor U12822 (N_12822,N_12699,N_12605);
or U12823 (N_12823,N_12671,N_12647);
and U12824 (N_12824,N_12739,N_12655);
and U12825 (N_12825,N_12712,N_12637);
nand U12826 (N_12826,N_12635,N_12752);
xnor U12827 (N_12827,N_12768,N_12793);
nor U12828 (N_12828,N_12661,N_12770);
and U12829 (N_12829,N_12672,N_12725);
or U12830 (N_12830,N_12619,N_12694);
nor U12831 (N_12831,N_12679,N_12621);
and U12832 (N_12832,N_12604,N_12778);
or U12833 (N_12833,N_12677,N_12719);
nand U12834 (N_12834,N_12761,N_12663);
and U12835 (N_12835,N_12763,N_12613);
xor U12836 (N_12836,N_12713,N_12690);
nor U12837 (N_12837,N_12662,N_12788);
nor U12838 (N_12838,N_12748,N_12706);
or U12839 (N_12839,N_12600,N_12757);
nand U12840 (N_12840,N_12628,N_12723);
nand U12841 (N_12841,N_12703,N_12777);
and U12842 (N_12842,N_12614,N_12782);
nand U12843 (N_12843,N_12629,N_12658);
nor U12844 (N_12844,N_12756,N_12710);
nand U12845 (N_12845,N_12697,N_12620);
and U12846 (N_12846,N_12668,N_12749);
or U12847 (N_12847,N_12769,N_12705);
or U12848 (N_12848,N_12785,N_12631);
or U12849 (N_12849,N_12726,N_12695);
nor U12850 (N_12850,N_12667,N_12698);
nand U12851 (N_12851,N_12745,N_12627);
xnor U12852 (N_12852,N_12794,N_12646);
nor U12853 (N_12853,N_12771,N_12704);
and U12854 (N_12854,N_12746,N_12743);
or U12855 (N_12855,N_12791,N_12798);
nor U12856 (N_12856,N_12700,N_12716);
xnor U12857 (N_12857,N_12741,N_12708);
or U12858 (N_12858,N_12660,N_12692);
xnor U12859 (N_12859,N_12623,N_12758);
and U12860 (N_12860,N_12645,N_12618);
and U12861 (N_12861,N_12670,N_12779);
and U12862 (N_12862,N_12718,N_12632);
or U12863 (N_12863,N_12617,N_12701);
xnor U12864 (N_12864,N_12680,N_12622);
xnor U12865 (N_12865,N_12783,N_12648);
nand U12866 (N_12866,N_12649,N_12747);
and U12867 (N_12867,N_12727,N_12608);
nand U12868 (N_12868,N_12744,N_12781);
nor U12869 (N_12869,N_12740,N_12610);
and U12870 (N_12870,N_12799,N_12717);
or U12871 (N_12871,N_12625,N_12750);
and U12872 (N_12872,N_12780,N_12686);
or U12873 (N_12873,N_12722,N_12615);
and U12874 (N_12874,N_12630,N_12642);
and U12875 (N_12875,N_12641,N_12787);
nand U12876 (N_12876,N_12612,N_12606);
nand U12877 (N_12877,N_12689,N_12792);
or U12878 (N_12878,N_12640,N_12653);
xnor U12879 (N_12879,N_12753,N_12666);
and U12880 (N_12880,N_12603,N_12673);
or U12881 (N_12881,N_12607,N_12732);
or U12882 (N_12882,N_12696,N_12650);
nor U12883 (N_12883,N_12624,N_12693);
nor U12884 (N_12884,N_12674,N_12688);
and U12885 (N_12885,N_12638,N_12775);
nor U12886 (N_12886,N_12759,N_12684);
xor U12887 (N_12887,N_12659,N_12602);
xor U12888 (N_12888,N_12654,N_12766);
nor U12889 (N_12889,N_12721,N_12609);
nand U12890 (N_12890,N_12643,N_12773);
nor U12891 (N_12891,N_12676,N_12724);
nor U12892 (N_12892,N_12728,N_12733);
nand U12893 (N_12893,N_12751,N_12754);
and U12894 (N_12894,N_12644,N_12795);
nand U12895 (N_12895,N_12776,N_12714);
nor U12896 (N_12896,N_12730,N_12767);
nor U12897 (N_12897,N_12711,N_12737);
nand U12898 (N_12898,N_12681,N_12657);
nor U12899 (N_12899,N_12742,N_12687);
or U12900 (N_12900,N_12682,N_12784);
nand U12901 (N_12901,N_12686,N_12696);
and U12902 (N_12902,N_12712,N_12778);
or U12903 (N_12903,N_12780,N_12669);
nor U12904 (N_12904,N_12783,N_12682);
xor U12905 (N_12905,N_12679,N_12638);
nor U12906 (N_12906,N_12770,N_12731);
or U12907 (N_12907,N_12790,N_12779);
or U12908 (N_12908,N_12736,N_12721);
or U12909 (N_12909,N_12798,N_12668);
nor U12910 (N_12910,N_12718,N_12661);
nor U12911 (N_12911,N_12716,N_12685);
nand U12912 (N_12912,N_12781,N_12651);
nand U12913 (N_12913,N_12617,N_12665);
xor U12914 (N_12914,N_12751,N_12629);
nand U12915 (N_12915,N_12742,N_12706);
nor U12916 (N_12916,N_12605,N_12751);
and U12917 (N_12917,N_12684,N_12753);
xnor U12918 (N_12918,N_12701,N_12637);
nor U12919 (N_12919,N_12754,N_12677);
xor U12920 (N_12920,N_12677,N_12736);
or U12921 (N_12921,N_12670,N_12713);
and U12922 (N_12922,N_12677,N_12610);
or U12923 (N_12923,N_12607,N_12664);
xor U12924 (N_12924,N_12669,N_12699);
nor U12925 (N_12925,N_12699,N_12659);
and U12926 (N_12926,N_12641,N_12645);
or U12927 (N_12927,N_12665,N_12684);
nor U12928 (N_12928,N_12789,N_12750);
and U12929 (N_12929,N_12772,N_12628);
or U12930 (N_12930,N_12636,N_12711);
or U12931 (N_12931,N_12793,N_12748);
and U12932 (N_12932,N_12611,N_12791);
nand U12933 (N_12933,N_12792,N_12795);
and U12934 (N_12934,N_12681,N_12700);
xnor U12935 (N_12935,N_12604,N_12632);
nand U12936 (N_12936,N_12618,N_12764);
or U12937 (N_12937,N_12711,N_12656);
nand U12938 (N_12938,N_12710,N_12651);
and U12939 (N_12939,N_12685,N_12649);
nor U12940 (N_12940,N_12657,N_12723);
nand U12941 (N_12941,N_12778,N_12799);
nor U12942 (N_12942,N_12645,N_12690);
and U12943 (N_12943,N_12735,N_12738);
nor U12944 (N_12944,N_12646,N_12658);
nor U12945 (N_12945,N_12769,N_12689);
or U12946 (N_12946,N_12743,N_12636);
xnor U12947 (N_12947,N_12722,N_12641);
nor U12948 (N_12948,N_12710,N_12752);
or U12949 (N_12949,N_12668,N_12615);
nand U12950 (N_12950,N_12687,N_12644);
and U12951 (N_12951,N_12692,N_12613);
nand U12952 (N_12952,N_12684,N_12650);
nor U12953 (N_12953,N_12677,N_12631);
or U12954 (N_12954,N_12630,N_12719);
and U12955 (N_12955,N_12644,N_12602);
nand U12956 (N_12956,N_12791,N_12645);
xor U12957 (N_12957,N_12698,N_12648);
nor U12958 (N_12958,N_12708,N_12785);
nand U12959 (N_12959,N_12662,N_12665);
or U12960 (N_12960,N_12695,N_12723);
xnor U12961 (N_12961,N_12781,N_12618);
xor U12962 (N_12962,N_12651,N_12602);
and U12963 (N_12963,N_12646,N_12662);
xnor U12964 (N_12964,N_12620,N_12792);
nor U12965 (N_12965,N_12734,N_12641);
or U12966 (N_12966,N_12681,N_12697);
nand U12967 (N_12967,N_12651,N_12665);
or U12968 (N_12968,N_12615,N_12794);
nand U12969 (N_12969,N_12790,N_12680);
and U12970 (N_12970,N_12643,N_12673);
xor U12971 (N_12971,N_12695,N_12756);
xnor U12972 (N_12972,N_12741,N_12755);
nor U12973 (N_12973,N_12722,N_12631);
xor U12974 (N_12974,N_12796,N_12799);
nor U12975 (N_12975,N_12616,N_12677);
nand U12976 (N_12976,N_12680,N_12645);
nor U12977 (N_12977,N_12642,N_12683);
and U12978 (N_12978,N_12623,N_12734);
xnor U12979 (N_12979,N_12675,N_12706);
nor U12980 (N_12980,N_12695,N_12753);
and U12981 (N_12981,N_12640,N_12669);
and U12982 (N_12982,N_12766,N_12618);
and U12983 (N_12983,N_12674,N_12617);
and U12984 (N_12984,N_12726,N_12739);
and U12985 (N_12985,N_12690,N_12600);
xnor U12986 (N_12986,N_12750,N_12638);
or U12987 (N_12987,N_12707,N_12633);
nand U12988 (N_12988,N_12779,N_12795);
xnor U12989 (N_12989,N_12721,N_12661);
or U12990 (N_12990,N_12687,N_12749);
nor U12991 (N_12991,N_12755,N_12652);
nand U12992 (N_12992,N_12740,N_12717);
and U12993 (N_12993,N_12772,N_12671);
nor U12994 (N_12994,N_12777,N_12753);
xnor U12995 (N_12995,N_12794,N_12766);
nand U12996 (N_12996,N_12628,N_12781);
xor U12997 (N_12997,N_12764,N_12713);
nand U12998 (N_12998,N_12642,N_12673);
xnor U12999 (N_12999,N_12719,N_12628);
nor U13000 (N_13000,N_12833,N_12926);
nor U13001 (N_13001,N_12805,N_12826);
xnor U13002 (N_13002,N_12888,N_12970);
or U13003 (N_13003,N_12835,N_12823);
and U13004 (N_13004,N_12899,N_12958);
or U13005 (N_13005,N_12868,N_12885);
or U13006 (N_13006,N_12879,N_12822);
nand U13007 (N_13007,N_12815,N_12957);
or U13008 (N_13008,N_12918,N_12900);
nand U13009 (N_13009,N_12865,N_12968);
nor U13010 (N_13010,N_12960,N_12800);
xnor U13011 (N_13011,N_12989,N_12842);
or U13012 (N_13012,N_12961,N_12906);
or U13013 (N_13013,N_12841,N_12983);
and U13014 (N_13014,N_12828,N_12809);
and U13015 (N_13015,N_12866,N_12992);
and U13016 (N_13016,N_12933,N_12880);
and U13017 (N_13017,N_12895,N_12858);
nor U13018 (N_13018,N_12802,N_12945);
nor U13019 (N_13019,N_12901,N_12981);
nor U13020 (N_13020,N_12808,N_12941);
nand U13021 (N_13021,N_12859,N_12829);
xor U13022 (N_13022,N_12988,N_12908);
or U13023 (N_13023,N_12924,N_12942);
nand U13024 (N_13024,N_12979,N_12812);
xnor U13025 (N_13025,N_12964,N_12846);
xnor U13026 (N_13026,N_12915,N_12889);
or U13027 (N_13027,N_12827,N_12905);
nor U13028 (N_13028,N_12814,N_12971);
xor U13029 (N_13029,N_12863,N_12872);
nand U13030 (N_13030,N_12946,N_12925);
nand U13031 (N_13031,N_12876,N_12912);
nor U13032 (N_13032,N_12896,N_12867);
or U13033 (N_13033,N_12874,N_12864);
nor U13034 (N_13034,N_12980,N_12853);
or U13035 (N_13035,N_12848,N_12984);
or U13036 (N_13036,N_12839,N_12855);
xnor U13037 (N_13037,N_12909,N_12999);
nand U13038 (N_13038,N_12852,N_12883);
xnor U13039 (N_13039,N_12840,N_12838);
nand U13040 (N_13040,N_12825,N_12978);
xnor U13041 (N_13041,N_12944,N_12904);
nand U13042 (N_13042,N_12949,N_12870);
nor U13043 (N_13043,N_12894,N_12916);
and U13044 (N_13044,N_12919,N_12920);
and U13045 (N_13045,N_12934,N_12881);
nor U13046 (N_13046,N_12807,N_12854);
xnor U13047 (N_13047,N_12821,N_12976);
or U13048 (N_13048,N_12887,N_12877);
and U13049 (N_13049,N_12950,N_12962);
or U13050 (N_13050,N_12917,N_12910);
or U13051 (N_13051,N_12860,N_12816);
and U13052 (N_13052,N_12834,N_12914);
and U13053 (N_13053,N_12886,N_12851);
or U13054 (N_13054,N_12803,N_12977);
or U13055 (N_13055,N_12813,N_12969);
nand U13056 (N_13056,N_12806,N_12998);
xor U13057 (N_13057,N_12993,N_12811);
xnor U13058 (N_13058,N_12973,N_12975);
and U13059 (N_13059,N_12938,N_12956);
and U13060 (N_13060,N_12990,N_12947);
xnor U13061 (N_13061,N_12804,N_12951);
nor U13062 (N_13062,N_12817,N_12850);
nand U13063 (N_13063,N_12972,N_12985);
nor U13064 (N_13064,N_12974,N_12845);
nor U13065 (N_13065,N_12898,N_12903);
or U13066 (N_13066,N_12922,N_12861);
xnor U13067 (N_13067,N_12818,N_12963);
xnor U13068 (N_13068,N_12953,N_12862);
nand U13069 (N_13069,N_12921,N_12982);
nand U13070 (N_13070,N_12952,N_12892);
nor U13071 (N_13071,N_12897,N_12986);
nand U13072 (N_13072,N_12836,N_12871);
nor U13073 (N_13073,N_12966,N_12890);
xnor U13074 (N_13074,N_12928,N_12955);
nor U13075 (N_13075,N_12967,N_12830);
or U13076 (N_13076,N_12843,N_12857);
nand U13077 (N_13077,N_12837,N_12932);
nor U13078 (N_13078,N_12810,N_12965);
or U13079 (N_13079,N_12873,N_12891);
or U13080 (N_13080,N_12996,N_12923);
or U13081 (N_13081,N_12959,N_12948);
nand U13082 (N_13082,N_12937,N_12875);
xor U13083 (N_13083,N_12893,N_12930);
or U13084 (N_13084,N_12994,N_12939);
nor U13085 (N_13085,N_12940,N_12856);
or U13086 (N_13086,N_12936,N_12931);
xor U13087 (N_13087,N_12847,N_12884);
and U13088 (N_13088,N_12878,N_12844);
and U13089 (N_13089,N_12869,N_12831);
nand U13090 (N_13090,N_12995,N_12902);
nor U13091 (N_13091,N_12929,N_12824);
nand U13092 (N_13092,N_12832,N_12819);
and U13093 (N_13093,N_12997,N_12849);
xnor U13094 (N_13094,N_12943,N_12820);
xor U13095 (N_13095,N_12913,N_12882);
nand U13096 (N_13096,N_12991,N_12927);
and U13097 (N_13097,N_12987,N_12935);
nor U13098 (N_13098,N_12907,N_12911);
nor U13099 (N_13099,N_12954,N_12801);
nand U13100 (N_13100,N_12855,N_12919);
or U13101 (N_13101,N_12930,N_12920);
nor U13102 (N_13102,N_12901,N_12939);
nor U13103 (N_13103,N_12926,N_12976);
xor U13104 (N_13104,N_12881,N_12800);
nor U13105 (N_13105,N_12959,N_12916);
and U13106 (N_13106,N_12918,N_12971);
or U13107 (N_13107,N_12863,N_12835);
nand U13108 (N_13108,N_12843,N_12813);
nand U13109 (N_13109,N_12876,N_12915);
nand U13110 (N_13110,N_12879,N_12818);
xor U13111 (N_13111,N_12987,N_12884);
and U13112 (N_13112,N_12894,N_12837);
xor U13113 (N_13113,N_12879,N_12840);
xor U13114 (N_13114,N_12990,N_12883);
nand U13115 (N_13115,N_12988,N_12897);
nor U13116 (N_13116,N_12908,N_12971);
and U13117 (N_13117,N_12915,N_12920);
and U13118 (N_13118,N_12805,N_12996);
nand U13119 (N_13119,N_12873,N_12954);
nor U13120 (N_13120,N_12872,N_12801);
xor U13121 (N_13121,N_12829,N_12885);
xor U13122 (N_13122,N_12812,N_12806);
nor U13123 (N_13123,N_12835,N_12900);
or U13124 (N_13124,N_12898,N_12886);
nor U13125 (N_13125,N_12941,N_12955);
nand U13126 (N_13126,N_12847,N_12878);
xnor U13127 (N_13127,N_12825,N_12959);
or U13128 (N_13128,N_12895,N_12962);
and U13129 (N_13129,N_12801,N_12852);
nand U13130 (N_13130,N_12914,N_12981);
nor U13131 (N_13131,N_12870,N_12979);
xor U13132 (N_13132,N_12801,N_12975);
and U13133 (N_13133,N_12978,N_12979);
nor U13134 (N_13134,N_12848,N_12853);
nor U13135 (N_13135,N_12808,N_12842);
nand U13136 (N_13136,N_12905,N_12939);
and U13137 (N_13137,N_12988,N_12924);
nor U13138 (N_13138,N_12917,N_12914);
or U13139 (N_13139,N_12828,N_12804);
xor U13140 (N_13140,N_12938,N_12881);
or U13141 (N_13141,N_12865,N_12903);
and U13142 (N_13142,N_12853,N_12970);
nand U13143 (N_13143,N_12800,N_12981);
or U13144 (N_13144,N_12860,N_12906);
nand U13145 (N_13145,N_12858,N_12832);
nand U13146 (N_13146,N_12988,N_12938);
nand U13147 (N_13147,N_12960,N_12932);
or U13148 (N_13148,N_12801,N_12886);
nor U13149 (N_13149,N_12845,N_12982);
and U13150 (N_13150,N_12850,N_12954);
or U13151 (N_13151,N_12907,N_12860);
and U13152 (N_13152,N_12959,N_12999);
and U13153 (N_13153,N_12888,N_12837);
nor U13154 (N_13154,N_12916,N_12817);
nor U13155 (N_13155,N_12858,N_12921);
nor U13156 (N_13156,N_12827,N_12896);
nand U13157 (N_13157,N_12834,N_12974);
xor U13158 (N_13158,N_12863,N_12911);
or U13159 (N_13159,N_12913,N_12993);
and U13160 (N_13160,N_12859,N_12923);
xnor U13161 (N_13161,N_12918,N_12876);
nand U13162 (N_13162,N_12907,N_12802);
nor U13163 (N_13163,N_12820,N_12801);
xor U13164 (N_13164,N_12829,N_12889);
and U13165 (N_13165,N_12814,N_12852);
and U13166 (N_13166,N_12943,N_12918);
nand U13167 (N_13167,N_12949,N_12976);
and U13168 (N_13168,N_12916,N_12831);
nand U13169 (N_13169,N_12898,N_12954);
xnor U13170 (N_13170,N_12909,N_12984);
nand U13171 (N_13171,N_12811,N_12953);
or U13172 (N_13172,N_12969,N_12879);
nor U13173 (N_13173,N_12815,N_12834);
nor U13174 (N_13174,N_12810,N_12993);
xor U13175 (N_13175,N_12870,N_12837);
xor U13176 (N_13176,N_12881,N_12890);
nor U13177 (N_13177,N_12964,N_12872);
nor U13178 (N_13178,N_12916,N_12936);
nand U13179 (N_13179,N_12916,N_12879);
nand U13180 (N_13180,N_12897,N_12916);
nor U13181 (N_13181,N_12969,N_12940);
or U13182 (N_13182,N_12808,N_12815);
xnor U13183 (N_13183,N_12822,N_12908);
nand U13184 (N_13184,N_12937,N_12801);
xor U13185 (N_13185,N_12989,N_12865);
and U13186 (N_13186,N_12947,N_12841);
or U13187 (N_13187,N_12989,N_12808);
or U13188 (N_13188,N_12839,N_12804);
xnor U13189 (N_13189,N_12958,N_12832);
and U13190 (N_13190,N_12875,N_12904);
nor U13191 (N_13191,N_12820,N_12939);
nor U13192 (N_13192,N_12822,N_12994);
or U13193 (N_13193,N_12836,N_12806);
nor U13194 (N_13194,N_12987,N_12894);
or U13195 (N_13195,N_12937,N_12910);
and U13196 (N_13196,N_12987,N_12842);
and U13197 (N_13197,N_12921,N_12903);
xor U13198 (N_13198,N_12848,N_12937);
or U13199 (N_13199,N_12925,N_12816);
nand U13200 (N_13200,N_13000,N_13039);
xor U13201 (N_13201,N_13122,N_13198);
or U13202 (N_13202,N_13157,N_13101);
nor U13203 (N_13203,N_13175,N_13092);
and U13204 (N_13204,N_13158,N_13123);
nand U13205 (N_13205,N_13139,N_13117);
xnor U13206 (N_13206,N_13032,N_13015);
nand U13207 (N_13207,N_13038,N_13180);
xnor U13208 (N_13208,N_13083,N_13024);
xnor U13209 (N_13209,N_13088,N_13150);
nand U13210 (N_13210,N_13067,N_13197);
and U13211 (N_13211,N_13046,N_13146);
xnor U13212 (N_13212,N_13089,N_13086);
xor U13213 (N_13213,N_13087,N_13164);
nor U13214 (N_13214,N_13070,N_13016);
and U13215 (N_13215,N_13134,N_13055);
nor U13216 (N_13216,N_13135,N_13199);
nand U13217 (N_13217,N_13140,N_13188);
nand U13218 (N_13218,N_13163,N_13001);
nor U13219 (N_13219,N_13144,N_13167);
xnor U13220 (N_13220,N_13081,N_13096);
and U13221 (N_13221,N_13011,N_13005);
nor U13222 (N_13222,N_13069,N_13151);
or U13223 (N_13223,N_13100,N_13002);
nor U13224 (N_13224,N_13186,N_13155);
xor U13225 (N_13225,N_13161,N_13022);
xor U13226 (N_13226,N_13078,N_13014);
nand U13227 (N_13227,N_13051,N_13115);
and U13228 (N_13228,N_13165,N_13133);
nand U13229 (N_13229,N_13023,N_13190);
nand U13230 (N_13230,N_13130,N_13107);
xnor U13231 (N_13231,N_13120,N_13154);
nand U13232 (N_13232,N_13181,N_13127);
and U13233 (N_13233,N_13068,N_13017);
nor U13234 (N_13234,N_13152,N_13119);
nor U13235 (N_13235,N_13160,N_13145);
nand U13236 (N_13236,N_13060,N_13042);
and U13237 (N_13237,N_13040,N_13073);
nand U13238 (N_13238,N_13072,N_13148);
and U13239 (N_13239,N_13006,N_13084);
and U13240 (N_13240,N_13065,N_13050);
nand U13241 (N_13241,N_13066,N_13007);
nand U13242 (N_13242,N_13129,N_13108);
and U13243 (N_13243,N_13174,N_13057);
nand U13244 (N_13244,N_13098,N_13193);
or U13245 (N_13245,N_13020,N_13079);
nor U13246 (N_13246,N_13192,N_13106);
nand U13247 (N_13247,N_13026,N_13185);
nor U13248 (N_13248,N_13037,N_13116);
nor U13249 (N_13249,N_13082,N_13137);
nor U13250 (N_13250,N_13169,N_13166);
nand U13251 (N_13251,N_13125,N_13075);
nand U13252 (N_13252,N_13138,N_13184);
nand U13253 (N_13253,N_13187,N_13131);
nor U13254 (N_13254,N_13004,N_13147);
and U13255 (N_13255,N_13010,N_13043);
xnor U13256 (N_13256,N_13177,N_13033);
or U13257 (N_13257,N_13031,N_13071);
and U13258 (N_13258,N_13105,N_13064);
xor U13259 (N_13259,N_13141,N_13091);
nor U13260 (N_13260,N_13030,N_13171);
nand U13261 (N_13261,N_13195,N_13097);
nor U13262 (N_13262,N_13156,N_13128);
and U13263 (N_13263,N_13109,N_13121);
or U13264 (N_13264,N_13085,N_13111);
or U13265 (N_13265,N_13104,N_13189);
or U13266 (N_13266,N_13194,N_13178);
nor U13267 (N_13267,N_13103,N_13142);
xor U13268 (N_13268,N_13153,N_13118);
xor U13269 (N_13269,N_13018,N_13021);
xor U13270 (N_13270,N_13025,N_13102);
and U13271 (N_13271,N_13172,N_13124);
nor U13272 (N_13272,N_13019,N_13059);
nand U13273 (N_13273,N_13036,N_13058);
or U13274 (N_13274,N_13080,N_13056);
xnor U13275 (N_13275,N_13009,N_13041);
xnor U13276 (N_13276,N_13110,N_13029);
nor U13277 (N_13277,N_13093,N_13074);
nor U13278 (N_13278,N_13183,N_13114);
xnor U13279 (N_13279,N_13113,N_13196);
xor U13280 (N_13280,N_13132,N_13034);
and U13281 (N_13281,N_13149,N_13077);
and U13282 (N_13282,N_13012,N_13168);
or U13283 (N_13283,N_13003,N_13047);
nand U13284 (N_13284,N_13126,N_13035);
and U13285 (N_13285,N_13045,N_13008);
nor U13286 (N_13286,N_13049,N_13094);
or U13287 (N_13287,N_13013,N_13143);
and U13288 (N_13288,N_13099,N_13159);
nand U13289 (N_13289,N_13062,N_13054);
and U13290 (N_13290,N_13191,N_13095);
or U13291 (N_13291,N_13182,N_13027);
nand U13292 (N_13292,N_13112,N_13176);
or U13293 (N_13293,N_13162,N_13063);
nand U13294 (N_13294,N_13028,N_13136);
and U13295 (N_13295,N_13053,N_13170);
and U13296 (N_13296,N_13179,N_13173);
and U13297 (N_13297,N_13044,N_13052);
or U13298 (N_13298,N_13076,N_13048);
and U13299 (N_13299,N_13090,N_13061);
nor U13300 (N_13300,N_13112,N_13193);
nand U13301 (N_13301,N_13086,N_13046);
and U13302 (N_13302,N_13034,N_13020);
nand U13303 (N_13303,N_13127,N_13000);
and U13304 (N_13304,N_13194,N_13031);
and U13305 (N_13305,N_13020,N_13059);
xor U13306 (N_13306,N_13088,N_13046);
and U13307 (N_13307,N_13040,N_13198);
xor U13308 (N_13308,N_13106,N_13034);
and U13309 (N_13309,N_13009,N_13083);
nor U13310 (N_13310,N_13080,N_13102);
nand U13311 (N_13311,N_13030,N_13128);
xor U13312 (N_13312,N_13011,N_13186);
xnor U13313 (N_13313,N_13071,N_13168);
or U13314 (N_13314,N_13011,N_13155);
nand U13315 (N_13315,N_13090,N_13101);
nand U13316 (N_13316,N_13110,N_13176);
nor U13317 (N_13317,N_13070,N_13037);
xnor U13318 (N_13318,N_13114,N_13108);
nor U13319 (N_13319,N_13193,N_13140);
and U13320 (N_13320,N_13068,N_13179);
and U13321 (N_13321,N_13015,N_13183);
and U13322 (N_13322,N_13129,N_13072);
nor U13323 (N_13323,N_13186,N_13094);
xor U13324 (N_13324,N_13088,N_13167);
nor U13325 (N_13325,N_13135,N_13035);
xnor U13326 (N_13326,N_13038,N_13112);
nand U13327 (N_13327,N_13175,N_13131);
xnor U13328 (N_13328,N_13173,N_13080);
nor U13329 (N_13329,N_13065,N_13024);
xor U13330 (N_13330,N_13162,N_13005);
or U13331 (N_13331,N_13194,N_13014);
nand U13332 (N_13332,N_13132,N_13062);
or U13333 (N_13333,N_13093,N_13114);
nor U13334 (N_13334,N_13034,N_13198);
xnor U13335 (N_13335,N_13183,N_13121);
and U13336 (N_13336,N_13016,N_13121);
xnor U13337 (N_13337,N_13167,N_13078);
and U13338 (N_13338,N_13186,N_13123);
nor U13339 (N_13339,N_13108,N_13189);
or U13340 (N_13340,N_13057,N_13094);
and U13341 (N_13341,N_13060,N_13059);
and U13342 (N_13342,N_13038,N_13019);
and U13343 (N_13343,N_13081,N_13173);
nand U13344 (N_13344,N_13146,N_13082);
nand U13345 (N_13345,N_13146,N_13152);
and U13346 (N_13346,N_13017,N_13097);
nand U13347 (N_13347,N_13074,N_13035);
nand U13348 (N_13348,N_13194,N_13003);
xor U13349 (N_13349,N_13000,N_13032);
and U13350 (N_13350,N_13144,N_13132);
nand U13351 (N_13351,N_13124,N_13121);
nand U13352 (N_13352,N_13052,N_13003);
nand U13353 (N_13353,N_13075,N_13197);
xnor U13354 (N_13354,N_13142,N_13151);
nor U13355 (N_13355,N_13107,N_13171);
xor U13356 (N_13356,N_13190,N_13024);
or U13357 (N_13357,N_13038,N_13075);
xnor U13358 (N_13358,N_13011,N_13144);
nand U13359 (N_13359,N_13161,N_13050);
xnor U13360 (N_13360,N_13105,N_13047);
and U13361 (N_13361,N_13054,N_13084);
nand U13362 (N_13362,N_13041,N_13195);
nand U13363 (N_13363,N_13133,N_13101);
and U13364 (N_13364,N_13197,N_13155);
nand U13365 (N_13365,N_13015,N_13053);
nor U13366 (N_13366,N_13077,N_13133);
and U13367 (N_13367,N_13085,N_13093);
xor U13368 (N_13368,N_13061,N_13145);
or U13369 (N_13369,N_13190,N_13163);
nand U13370 (N_13370,N_13109,N_13001);
xor U13371 (N_13371,N_13195,N_13029);
nand U13372 (N_13372,N_13006,N_13094);
or U13373 (N_13373,N_13186,N_13093);
nor U13374 (N_13374,N_13053,N_13070);
or U13375 (N_13375,N_13038,N_13174);
or U13376 (N_13376,N_13115,N_13170);
nand U13377 (N_13377,N_13150,N_13152);
and U13378 (N_13378,N_13100,N_13104);
xor U13379 (N_13379,N_13041,N_13001);
nand U13380 (N_13380,N_13171,N_13178);
nor U13381 (N_13381,N_13056,N_13005);
xor U13382 (N_13382,N_13065,N_13144);
xor U13383 (N_13383,N_13188,N_13045);
or U13384 (N_13384,N_13067,N_13161);
or U13385 (N_13385,N_13116,N_13023);
xnor U13386 (N_13386,N_13046,N_13154);
nor U13387 (N_13387,N_13170,N_13178);
xor U13388 (N_13388,N_13137,N_13073);
and U13389 (N_13389,N_13186,N_13054);
nand U13390 (N_13390,N_13017,N_13098);
xnor U13391 (N_13391,N_13193,N_13164);
xnor U13392 (N_13392,N_13071,N_13088);
nor U13393 (N_13393,N_13185,N_13118);
xnor U13394 (N_13394,N_13103,N_13127);
xnor U13395 (N_13395,N_13012,N_13183);
nor U13396 (N_13396,N_13003,N_13045);
or U13397 (N_13397,N_13180,N_13134);
nor U13398 (N_13398,N_13097,N_13159);
xnor U13399 (N_13399,N_13167,N_13068);
xor U13400 (N_13400,N_13288,N_13232);
and U13401 (N_13401,N_13287,N_13271);
nor U13402 (N_13402,N_13234,N_13334);
xnor U13403 (N_13403,N_13318,N_13265);
or U13404 (N_13404,N_13361,N_13391);
nor U13405 (N_13405,N_13349,N_13270);
nor U13406 (N_13406,N_13333,N_13290);
xnor U13407 (N_13407,N_13310,N_13370);
and U13408 (N_13408,N_13252,N_13279);
and U13409 (N_13409,N_13345,N_13217);
and U13410 (N_13410,N_13337,N_13254);
xor U13411 (N_13411,N_13249,N_13202);
nand U13412 (N_13412,N_13352,N_13214);
and U13413 (N_13413,N_13259,N_13253);
nand U13414 (N_13414,N_13387,N_13219);
nand U13415 (N_13415,N_13237,N_13307);
nor U13416 (N_13416,N_13236,N_13289);
or U13417 (N_13417,N_13348,N_13221);
and U13418 (N_13418,N_13229,N_13342);
and U13419 (N_13419,N_13315,N_13274);
or U13420 (N_13420,N_13353,N_13233);
xor U13421 (N_13421,N_13244,N_13346);
or U13422 (N_13422,N_13312,N_13203);
nand U13423 (N_13423,N_13378,N_13360);
nor U13424 (N_13424,N_13322,N_13308);
nand U13425 (N_13425,N_13386,N_13332);
nand U13426 (N_13426,N_13206,N_13328);
or U13427 (N_13427,N_13351,N_13245);
nor U13428 (N_13428,N_13363,N_13235);
and U13429 (N_13429,N_13388,N_13331);
nand U13430 (N_13430,N_13211,N_13220);
xnor U13431 (N_13431,N_13286,N_13281);
nand U13432 (N_13432,N_13303,N_13296);
nand U13433 (N_13433,N_13304,N_13326);
xor U13434 (N_13434,N_13341,N_13263);
or U13435 (N_13435,N_13323,N_13306);
nor U13436 (N_13436,N_13339,N_13284);
xor U13437 (N_13437,N_13314,N_13359);
xnor U13438 (N_13438,N_13273,N_13218);
nand U13439 (N_13439,N_13207,N_13264);
or U13440 (N_13440,N_13258,N_13355);
nor U13441 (N_13441,N_13226,N_13231);
or U13442 (N_13442,N_13397,N_13390);
nor U13443 (N_13443,N_13278,N_13241);
xor U13444 (N_13444,N_13313,N_13301);
nand U13445 (N_13445,N_13392,N_13395);
xnor U13446 (N_13446,N_13257,N_13283);
nor U13447 (N_13447,N_13366,N_13275);
xor U13448 (N_13448,N_13327,N_13210);
and U13449 (N_13449,N_13396,N_13336);
nand U13450 (N_13450,N_13230,N_13381);
nand U13451 (N_13451,N_13223,N_13380);
or U13452 (N_13452,N_13317,N_13276);
xor U13453 (N_13453,N_13347,N_13200);
xnor U13454 (N_13454,N_13238,N_13389);
or U13455 (N_13455,N_13377,N_13399);
xnor U13456 (N_13456,N_13374,N_13269);
nor U13457 (N_13457,N_13225,N_13251);
xor U13458 (N_13458,N_13309,N_13372);
nor U13459 (N_13459,N_13379,N_13209);
nor U13460 (N_13460,N_13268,N_13260);
xor U13461 (N_13461,N_13213,N_13375);
or U13462 (N_13462,N_13205,N_13324);
or U13463 (N_13463,N_13300,N_13291);
nor U13464 (N_13464,N_13297,N_13316);
nor U13465 (N_13465,N_13340,N_13204);
or U13466 (N_13466,N_13295,N_13382);
nor U13467 (N_13467,N_13282,N_13365);
or U13468 (N_13468,N_13299,N_13293);
nor U13469 (N_13469,N_13329,N_13376);
or U13470 (N_13470,N_13247,N_13215);
or U13471 (N_13471,N_13384,N_13227);
nor U13472 (N_13472,N_13261,N_13201);
and U13473 (N_13473,N_13240,N_13311);
and U13474 (N_13474,N_13362,N_13350);
or U13475 (N_13475,N_13364,N_13302);
and U13476 (N_13476,N_13369,N_13367);
or U13477 (N_13477,N_13262,N_13321);
nand U13478 (N_13478,N_13243,N_13280);
and U13479 (N_13479,N_13398,N_13354);
and U13480 (N_13480,N_13298,N_13208);
and U13481 (N_13481,N_13277,N_13272);
nand U13482 (N_13482,N_13325,N_13266);
xor U13483 (N_13483,N_13250,N_13292);
nor U13484 (N_13484,N_13358,N_13338);
nor U13485 (N_13485,N_13385,N_13368);
or U13486 (N_13486,N_13246,N_13343);
nand U13487 (N_13487,N_13267,N_13357);
nor U13488 (N_13488,N_13255,N_13294);
and U13489 (N_13489,N_13239,N_13371);
nor U13490 (N_13490,N_13330,N_13224);
nor U13491 (N_13491,N_13319,N_13356);
nor U13492 (N_13492,N_13212,N_13320);
xnor U13493 (N_13493,N_13373,N_13228);
xnor U13494 (N_13494,N_13344,N_13242);
nand U13495 (N_13495,N_13285,N_13256);
and U13496 (N_13496,N_13335,N_13222);
or U13497 (N_13497,N_13248,N_13394);
nand U13498 (N_13498,N_13305,N_13393);
nand U13499 (N_13499,N_13216,N_13383);
nor U13500 (N_13500,N_13237,N_13303);
and U13501 (N_13501,N_13321,N_13391);
and U13502 (N_13502,N_13302,N_13216);
nor U13503 (N_13503,N_13252,N_13307);
and U13504 (N_13504,N_13318,N_13330);
nand U13505 (N_13505,N_13275,N_13276);
and U13506 (N_13506,N_13301,N_13368);
nor U13507 (N_13507,N_13211,N_13230);
nand U13508 (N_13508,N_13248,N_13327);
xor U13509 (N_13509,N_13383,N_13274);
or U13510 (N_13510,N_13270,N_13214);
and U13511 (N_13511,N_13375,N_13277);
and U13512 (N_13512,N_13264,N_13334);
or U13513 (N_13513,N_13394,N_13202);
xnor U13514 (N_13514,N_13370,N_13213);
and U13515 (N_13515,N_13344,N_13363);
xor U13516 (N_13516,N_13296,N_13275);
nand U13517 (N_13517,N_13353,N_13271);
nor U13518 (N_13518,N_13292,N_13245);
or U13519 (N_13519,N_13336,N_13326);
nor U13520 (N_13520,N_13223,N_13331);
xnor U13521 (N_13521,N_13343,N_13382);
nor U13522 (N_13522,N_13364,N_13366);
xnor U13523 (N_13523,N_13360,N_13301);
nand U13524 (N_13524,N_13389,N_13356);
or U13525 (N_13525,N_13206,N_13236);
and U13526 (N_13526,N_13372,N_13283);
and U13527 (N_13527,N_13357,N_13300);
and U13528 (N_13528,N_13200,N_13264);
xnor U13529 (N_13529,N_13362,N_13353);
or U13530 (N_13530,N_13352,N_13390);
xnor U13531 (N_13531,N_13277,N_13360);
xor U13532 (N_13532,N_13393,N_13309);
and U13533 (N_13533,N_13379,N_13275);
nor U13534 (N_13534,N_13332,N_13226);
and U13535 (N_13535,N_13357,N_13292);
nor U13536 (N_13536,N_13231,N_13295);
nand U13537 (N_13537,N_13224,N_13208);
nor U13538 (N_13538,N_13393,N_13214);
nand U13539 (N_13539,N_13242,N_13346);
and U13540 (N_13540,N_13395,N_13389);
nand U13541 (N_13541,N_13361,N_13297);
nor U13542 (N_13542,N_13345,N_13330);
or U13543 (N_13543,N_13240,N_13339);
or U13544 (N_13544,N_13227,N_13266);
nand U13545 (N_13545,N_13254,N_13295);
nor U13546 (N_13546,N_13383,N_13361);
or U13547 (N_13547,N_13310,N_13224);
nand U13548 (N_13548,N_13350,N_13390);
nor U13549 (N_13549,N_13291,N_13333);
nor U13550 (N_13550,N_13202,N_13339);
and U13551 (N_13551,N_13339,N_13327);
xor U13552 (N_13552,N_13325,N_13366);
xor U13553 (N_13553,N_13212,N_13348);
and U13554 (N_13554,N_13388,N_13247);
or U13555 (N_13555,N_13332,N_13344);
or U13556 (N_13556,N_13372,N_13205);
xor U13557 (N_13557,N_13365,N_13208);
xnor U13558 (N_13558,N_13217,N_13257);
or U13559 (N_13559,N_13326,N_13311);
nor U13560 (N_13560,N_13324,N_13210);
nor U13561 (N_13561,N_13294,N_13326);
xnor U13562 (N_13562,N_13344,N_13309);
nor U13563 (N_13563,N_13208,N_13299);
nand U13564 (N_13564,N_13392,N_13315);
nor U13565 (N_13565,N_13359,N_13363);
xor U13566 (N_13566,N_13240,N_13338);
and U13567 (N_13567,N_13391,N_13202);
xor U13568 (N_13568,N_13280,N_13289);
or U13569 (N_13569,N_13275,N_13278);
xnor U13570 (N_13570,N_13317,N_13371);
nor U13571 (N_13571,N_13223,N_13340);
nor U13572 (N_13572,N_13344,N_13379);
or U13573 (N_13573,N_13247,N_13271);
xor U13574 (N_13574,N_13268,N_13272);
nand U13575 (N_13575,N_13286,N_13324);
and U13576 (N_13576,N_13243,N_13356);
or U13577 (N_13577,N_13237,N_13317);
xnor U13578 (N_13578,N_13212,N_13333);
xnor U13579 (N_13579,N_13355,N_13373);
or U13580 (N_13580,N_13366,N_13322);
and U13581 (N_13581,N_13347,N_13335);
nand U13582 (N_13582,N_13295,N_13283);
and U13583 (N_13583,N_13354,N_13356);
xnor U13584 (N_13584,N_13246,N_13359);
or U13585 (N_13585,N_13331,N_13316);
and U13586 (N_13586,N_13374,N_13341);
and U13587 (N_13587,N_13318,N_13244);
nor U13588 (N_13588,N_13245,N_13251);
nor U13589 (N_13589,N_13312,N_13205);
and U13590 (N_13590,N_13278,N_13377);
and U13591 (N_13591,N_13290,N_13254);
and U13592 (N_13592,N_13222,N_13216);
xnor U13593 (N_13593,N_13365,N_13339);
or U13594 (N_13594,N_13351,N_13318);
or U13595 (N_13595,N_13393,N_13274);
or U13596 (N_13596,N_13217,N_13254);
xor U13597 (N_13597,N_13275,N_13313);
and U13598 (N_13598,N_13376,N_13294);
xnor U13599 (N_13599,N_13309,N_13381);
or U13600 (N_13600,N_13524,N_13558);
xor U13601 (N_13601,N_13571,N_13547);
or U13602 (N_13602,N_13491,N_13508);
xor U13603 (N_13603,N_13507,N_13549);
nand U13604 (N_13604,N_13527,N_13523);
nor U13605 (N_13605,N_13409,N_13461);
nand U13606 (N_13606,N_13484,N_13554);
nor U13607 (N_13607,N_13439,N_13453);
or U13608 (N_13608,N_13522,N_13521);
nor U13609 (N_13609,N_13591,N_13564);
or U13610 (N_13610,N_13586,N_13421);
or U13611 (N_13611,N_13535,N_13451);
and U13612 (N_13612,N_13592,N_13542);
or U13613 (N_13613,N_13427,N_13533);
and U13614 (N_13614,N_13401,N_13477);
nor U13615 (N_13615,N_13436,N_13450);
xor U13616 (N_13616,N_13539,N_13515);
nor U13617 (N_13617,N_13452,N_13541);
or U13618 (N_13618,N_13504,N_13584);
or U13619 (N_13619,N_13486,N_13556);
nor U13620 (N_13620,N_13537,N_13560);
and U13621 (N_13621,N_13438,N_13414);
or U13622 (N_13622,N_13513,N_13440);
xnor U13623 (N_13623,N_13481,N_13526);
or U13624 (N_13624,N_13506,N_13503);
and U13625 (N_13625,N_13550,N_13403);
nand U13626 (N_13626,N_13581,N_13562);
or U13627 (N_13627,N_13411,N_13579);
and U13628 (N_13628,N_13502,N_13434);
nand U13629 (N_13629,N_13566,N_13509);
and U13630 (N_13630,N_13475,N_13531);
nand U13631 (N_13631,N_13460,N_13570);
nor U13632 (N_13632,N_13448,N_13467);
xor U13633 (N_13633,N_13561,N_13543);
nand U13634 (N_13634,N_13407,N_13573);
xor U13635 (N_13635,N_13472,N_13410);
or U13636 (N_13636,N_13424,N_13557);
xnor U13637 (N_13637,N_13446,N_13431);
or U13638 (N_13638,N_13532,N_13488);
nor U13639 (N_13639,N_13490,N_13551);
xor U13640 (N_13640,N_13455,N_13480);
and U13641 (N_13641,N_13470,N_13546);
nor U13642 (N_13642,N_13415,N_13548);
nor U13643 (N_13643,N_13497,N_13516);
nor U13644 (N_13644,N_13514,N_13444);
nor U13645 (N_13645,N_13441,N_13498);
or U13646 (N_13646,N_13593,N_13589);
nand U13647 (N_13647,N_13463,N_13575);
nand U13648 (N_13648,N_13494,N_13572);
xor U13649 (N_13649,N_13587,N_13588);
nor U13650 (N_13650,N_13483,N_13528);
nor U13651 (N_13651,N_13529,N_13469);
or U13652 (N_13652,N_13492,N_13433);
or U13653 (N_13653,N_13555,N_13582);
nor U13654 (N_13654,N_13406,N_13518);
nand U13655 (N_13655,N_13422,N_13519);
nor U13656 (N_13656,N_13417,N_13530);
and U13657 (N_13657,N_13597,N_13520);
nor U13658 (N_13658,N_13496,N_13569);
and U13659 (N_13659,N_13559,N_13493);
nand U13660 (N_13660,N_13479,N_13482);
or U13661 (N_13661,N_13499,N_13456);
nand U13662 (N_13662,N_13487,N_13567);
or U13663 (N_13663,N_13471,N_13576);
nor U13664 (N_13664,N_13580,N_13585);
and U13665 (N_13665,N_13402,N_13512);
xor U13666 (N_13666,N_13423,N_13447);
nand U13667 (N_13667,N_13552,N_13468);
or U13668 (N_13668,N_13544,N_13594);
or U13669 (N_13669,N_13404,N_13525);
xnor U13670 (N_13670,N_13437,N_13599);
or U13671 (N_13671,N_13426,N_13416);
xor U13672 (N_13672,N_13419,N_13459);
nor U13673 (N_13673,N_13553,N_13500);
nand U13674 (N_13674,N_13538,N_13595);
xor U13675 (N_13675,N_13583,N_13545);
or U13676 (N_13676,N_13443,N_13405);
or U13677 (N_13677,N_13485,N_13454);
or U13678 (N_13678,N_13565,N_13430);
nor U13679 (N_13679,N_13501,N_13442);
xnor U13680 (N_13680,N_13429,N_13464);
nand U13681 (N_13681,N_13457,N_13408);
nor U13682 (N_13682,N_13445,N_13536);
or U13683 (N_13683,N_13478,N_13473);
nor U13684 (N_13684,N_13476,N_13425);
nand U13685 (N_13685,N_13596,N_13466);
nand U13686 (N_13686,N_13534,N_13489);
nand U13687 (N_13687,N_13598,N_13458);
nor U13688 (N_13688,N_13568,N_13505);
nor U13689 (N_13689,N_13413,N_13590);
and U13690 (N_13690,N_13428,N_13510);
or U13691 (N_13691,N_13418,N_13578);
xnor U13692 (N_13692,N_13435,N_13540);
nor U13693 (N_13693,N_13517,N_13511);
or U13694 (N_13694,N_13474,N_13449);
and U13695 (N_13695,N_13420,N_13400);
or U13696 (N_13696,N_13432,N_13462);
nand U13697 (N_13697,N_13495,N_13563);
or U13698 (N_13698,N_13574,N_13412);
or U13699 (N_13699,N_13465,N_13577);
and U13700 (N_13700,N_13561,N_13442);
nor U13701 (N_13701,N_13530,N_13579);
nand U13702 (N_13702,N_13552,N_13475);
nand U13703 (N_13703,N_13507,N_13568);
xnor U13704 (N_13704,N_13560,N_13508);
or U13705 (N_13705,N_13441,N_13480);
xor U13706 (N_13706,N_13559,N_13442);
xnor U13707 (N_13707,N_13402,N_13463);
and U13708 (N_13708,N_13502,N_13575);
xnor U13709 (N_13709,N_13584,N_13456);
or U13710 (N_13710,N_13563,N_13506);
nor U13711 (N_13711,N_13528,N_13473);
nor U13712 (N_13712,N_13439,N_13477);
or U13713 (N_13713,N_13401,N_13443);
or U13714 (N_13714,N_13482,N_13464);
xnor U13715 (N_13715,N_13569,N_13497);
xor U13716 (N_13716,N_13544,N_13412);
nand U13717 (N_13717,N_13571,N_13566);
or U13718 (N_13718,N_13414,N_13547);
or U13719 (N_13719,N_13584,N_13487);
and U13720 (N_13720,N_13504,N_13583);
and U13721 (N_13721,N_13508,N_13440);
or U13722 (N_13722,N_13530,N_13542);
nor U13723 (N_13723,N_13491,N_13405);
xor U13724 (N_13724,N_13506,N_13437);
or U13725 (N_13725,N_13484,N_13543);
xnor U13726 (N_13726,N_13418,N_13532);
and U13727 (N_13727,N_13561,N_13569);
nor U13728 (N_13728,N_13475,N_13467);
or U13729 (N_13729,N_13452,N_13498);
and U13730 (N_13730,N_13487,N_13588);
or U13731 (N_13731,N_13564,N_13560);
and U13732 (N_13732,N_13587,N_13466);
nand U13733 (N_13733,N_13521,N_13468);
and U13734 (N_13734,N_13559,N_13405);
xor U13735 (N_13735,N_13488,N_13493);
or U13736 (N_13736,N_13596,N_13579);
nor U13737 (N_13737,N_13511,N_13533);
and U13738 (N_13738,N_13479,N_13545);
nand U13739 (N_13739,N_13462,N_13561);
and U13740 (N_13740,N_13421,N_13455);
and U13741 (N_13741,N_13433,N_13458);
or U13742 (N_13742,N_13497,N_13437);
and U13743 (N_13743,N_13545,N_13438);
and U13744 (N_13744,N_13539,N_13411);
and U13745 (N_13745,N_13408,N_13530);
nor U13746 (N_13746,N_13527,N_13530);
xor U13747 (N_13747,N_13446,N_13453);
and U13748 (N_13748,N_13598,N_13405);
nor U13749 (N_13749,N_13426,N_13404);
nor U13750 (N_13750,N_13414,N_13450);
xnor U13751 (N_13751,N_13597,N_13541);
nor U13752 (N_13752,N_13582,N_13569);
or U13753 (N_13753,N_13566,N_13525);
nor U13754 (N_13754,N_13459,N_13536);
nor U13755 (N_13755,N_13408,N_13445);
nand U13756 (N_13756,N_13485,N_13516);
and U13757 (N_13757,N_13420,N_13498);
or U13758 (N_13758,N_13469,N_13445);
nor U13759 (N_13759,N_13513,N_13520);
and U13760 (N_13760,N_13510,N_13469);
or U13761 (N_13761,N_13501,N_13580);
nand U13762 (N_13762,N_13413,N_13558);
nor U13763 (N_13763,N_13479,N_13594);
nand U13764 (N_13764,N_13565,N_13592);
or U13765 (N_13765,N_13554,N_13570);
and U13766 (N_13766,N_13466,N_13508);
xor U13767 (N_13767,N_13471,N_13418);
nor U13768 (N_13768,N_13405,N_13532);
and U13769 (N_13769,N_13416,N_13492);
and U13770 (N_13770,N_13527,N_13589);
and U13771 (N_13771,N_13544,N_13402);
nand U13772 (N_13772,N_13491,N_13469);
or U13773 (N_13773,N_13510,N_13496);
or U13774 (N_13774,N_13467,N_13472);
xor U13775 (N_13775,N_13592,N_13477);
xnor U13776 (N_13776,N_13406,N_13510);
nand U13777 (N_13777,N_13498,N_13502);
and U13778 (N_13778,N_13413,N_13448);
nor U13779 (N_13779,N_13404,N_13499);
nor U13780 (N_13780,N_13433,N_13479);
nand U13781 (N_13781,N_13462,N_13571);
or U13782 (N_13782,N_13424,N_13475);
nand U13783 (N_13783,N_13479,N_13567);
nor U13784 (N_13784,N_13510,N_13461);
nor U13785 (N_13785,N_13457,N_13591);
nand U13786 (N_13786,N_13453,N_13433);
nor U13787 (N_13787,N_13587,N_13484);
nand U13788 (N_13788,N_13483,N_13543);
nor U13789 (N_13789,N_13413,N_13475);
nor U13790 (N_13790,N_13500,N_13485);
nor U13791 (N_13791,N_13520,N_13599);
and U13792 (N_13792,N_13524,N_13405);
nand U13793 (N_13793,N_13581,N_13589);
xnor U13794 (N_13794,N_13472,N_13491);
or U13795 (N_13795,N_13528,N_13587);
nor U13796 (N_13796,N_13515,N_13543);
or U13797 (N_13797,N_13471,N_13451);
nand U13798 (N_13798,N_13406,N_13598);
nor U13799 (N_13799,N_13553,N_13450);
nand U13800 (N_13800,N_13758,N_13677);
xnor U13801 (N_13801,N_13723,N_13654);
nor U13802 (N_13802,N_13761,N_13688);
nand U13803 (N_13803,N_13691,N_13754);
or U13804 (N_13804,N_13608,N_13774);
xor U13805 (N_13805,N_13744,N_13749);
xor U13806 (N_13806,N_13604,N_13743);
or U13807 (N_13807,N_13724,N_13696);
nand U13808 (N_13808,N_13718,N_13612);
or U13809 (N_13809,N_13660,N_13648);
nand U13810 (N_13810,N_13630,N_13706);
nand U13811 (N_13811,N_13631,N_13759);
xor U13812 (N_13812,N_13610,N_13663);
or U13813 (N_13813,N_13798,N_13791);
xnor U13814 (N_13814,N_13737,N_13679);
nand U13815 (N_13815,N_13767,N_13680);
nor U13816 (N_13816,N_13622,N_13795);
nand U13817 (N_13817,N_13739,N_13678);
nor U13818 (N_13818,N_13632,N_13765);
or U13819 (N_13819,N_13641,N_13670);
or U13820 (N_13820,N_13713,N_13779);
nand U13821 (N_13821,N_13789,N_13689);
nor U13822 (N_13822,N_13729,N_13783);
nor U13823 (N_13823,N_13618,N_13726);
nand U13824 (N_13824,N_13634,N_13674);
and U13825 (N_13825,N_13757,N_13752);
nand U13826 (N_13826,N_13614,N_13609);
and U13827 (N_13827,N_13751,N_13727);
xor U13828 (N_13828,N_13644,N_13709);
or U13829 (N_13829,N_13766,N_13620);
and U13830 (N_13830,N_13717,N_13627);
nor U13831 (N_13831,N_13653,N_13672);
or U13832 (N_13832,N_13658,N_13721);
xnor U13833 (N_13833,N_13719,N_13643);
and U13834 (N_13834,N_13705,N_13628);
nor U13835 (N_13835,N_13728,N_13637);
and U13836 (N_13836,N_13732,N_13683);
nor U13837 (N_13837,N_13745,N_13776);
or U13838 (N_13838,N_13642,N_13699);
xnor U13839 (N_13839,N_13716,N_13623);
or U13840 (N_13840,N_13778,N_13617);
xnor U13841 (N_13841,N_13711,N_13764);
nand U13842 (N_13842,N_13700,N_13746);
nor U13843 (N_13843,N_13686,N_13707);
or U13844 (N_13844,N_13772,N_13602);
nor U13845 (N_13845,N_13792,N_13733);
nand U13846 (N_13846,N_13701,N_13681);
and U13847 (N_13847,N_13742,N_13760);
nand U13848 (N_13848,N_13661,N_13731);
nand U13849 (N_13849,N_13629,N_13646);
and U13850 (N_13850,N_13606,N_13626);
and U13851 (N_13851,N_13712,N_13607);
nor U13852 (N_13852,N_13676,N_13799);
or U13853 (N_13853,N_13753,N_13756);
xor U13854 (N_13854,N_13796,N_13704);
nand U13855 (N_13855,N_13665,N_13673);
xor U13856 (N_13856,N_13695,N_13651);
xor U13857 (N_13857,N_13619,N_13720);
nand U13858 (N_13858,N_13736,N_13730);
xor U13859 (N_13859,N_13750,N_13645);
nor U13860 (N_13860,N_13781,N_13667);
nand U13861 (N_13861,N_13621,N_13762);
and U13862 (N_13862,N_13668,N_13685);
and U13863 (N_13863,N_13664,N_13682);
and U13864 (N_13864,N_13649,N_13636);
nand U13865 (N_13865,N_13611,N_13770);
and U13866 (N_13866,N_13697,N_13755);
xnor U13867 (N_13867,N_13615,N_13777);
nor U13868 (N_13868,N_13793,N_13741);
nor U13869 (N_13869,N_13773,N_13635);
xnor U13870 (N_13870,N_13640,N_13738);
xnor U13871 (N_13871,N_13616,N_13603);
nand U13872 (N_13872,N_13708,N_13784);
nand U13873 (N_13873,N_13652,N_13790);
or U13874 (N_13874,N_13625,N_13671);
and U13875 (N_13875,N_13639,N_13684);
or U13876 (N_13876,N_13692,N_13715);
nand U13877 (N_13877,N_13787,N_13647);
or U13878 (N_13878,N_13771,N_13734);
nand U13879 (N_13879,N_13702,N_13657);
nor U13880 (N_13880,N_13624,N_13633);
nor U13881 (N_13881,N_13788,N_13675);
nor U13882 (N_13882,N_13785,N_13794);
nor U13883 (N_13883,N_13613,N_13735);
nor U13884 (N_13884,N_13725,N_13601);
nor U13885 (N_13885,N_13655,N_13690);
nand U13886 (N_13886,N_13662,N_13782);
or U13887 (N_13887,N_13605,N_13703);
and U13888 (N_13888,N_13786,N_13714);
nand U13889 (N_13889,N_13722,N_13747);
nand U13890 (N_13890,N_13656,N_13659);
or U13891 (N_13891,N_13797,N_13768);
or U13892 (N_13892,N_13740,N_13650);
nand U13893 (N_13893,N_13669,N_13775);
nand U13894 (N_13894,N_13710,N_13763);
nor U13895 (N_13895,N_13600,N_13638);
xor U13896 (N_13896,N_13666,N_13687);
or U13897 (N_13897,N_13769,N_13780);
and U13898 (N_13898,N_13693,N_13698);
and U13899 (N_13899,N_13748,N_13694);
nand U13900 (N_13900,N_13606,N_13650);
and U13901 (N_13901,N_13672,N_13601);
xor U13902 (N_13902,N_13734,N_13606);
and U13903 (N_13903,N_13744,N_13662);
xor U13904 (N_13904,N_13665,N_13611);
nor U13905 (N_13905,N_13632,N_13642);
nor U13906 (N_13906,N_13799,N_13714);
or U13907 (N_13907,N_13748,N_13727);
xor U13908 (N_13908,N_13636,N_13762);
and U13909 (N_13909,N_13653,N_13656);
nor U13910 (N_13910,N_13691,N_13708);
nor U13911 (N_13911,N_13681,N_13709);
xnor U13912 (N_13912,N_13786,N_13621);
nor U13913 (N_13913,N_13739,N_13732);
nand U13914 (N_13914,N_13642,N_13617);
and U13915 (N_13915,N_13701,N_13645);
or U13916 (N_13916,N_13709,N_13609);
and U13917 (N_13917,N_13711,N_13732);
or U13918 (N_13918,N_13787,N_13628);
nor U13919 (N_13919,N_13700,N_13716);
xor U13920 (N_13920,N_13762,N_13742);
and U13921 (N_13921,N_13796,N_13603);
xor U13922 (N_13922,N_13699,N_13723);
xnor U13923 (N_13923,N_13629,N_13665);
xnor U13924 (N_13924,N_13647,N_13712);
xnor U13925 (N_13925,N_13736,N_13729);
xor U13926 (N_13926,N_13749,N_13706);
xor U13927 (N_13927,N_13763,N_13708);
or U13928 (N_13928,N_13655,N_13625);
nand U13929 (N_13929,N_13688,N_13638);
nor U13930 (N_13930,N_13618,N_13793);
nor U13931 (N_13931,N_13649,N_13658);
or U13932 (N_13932,N_13790,N_13653);
or U13933 (N_13933,N_13746,N_13665);
nor U13934 (N_13934,N_13735,N_13660);
xnor U13935 (N_13935,N_13784,N_13732);
nand U13936 (N_13936,N_13795,N_13721);
nand U13937 (N_13937,N_13756,N_13773);
and U13938 (N_13938,N_13646,N_13795);
xor U13939 (N_13939,N_13793,N_13643);
and U13940 (N_13940,N_13693,N_13774);
and U13941 (N_13941,N_13793,N_13711);
and U13942 (N_13942,N_13667,N_13659);
xor U13943 (N_13943,N_13798,N_13650);
or U13944 (N_13944,N_13794,N_13713);
nor U13945 (N_13945,N_13752,N_13764);
and U13946 (N_13946,N_13795,N_13655);
and U13947 (N_13947,N_13753,N_13640);
nand U13948 (N_13948,N_13644,N_13667);
nand U13949 (N_13949,N_13787,N_13775);
nand U13950 (N_13950,N_13722,N_13640);
nand U13951 (N_13951,N_13689,N_13690);
xnor U13952 (N_13952,N_13652,N_13767);
xnor U13953 (N_13953,N_13762,N_13613);
nor U13954 (N_13954,N_13751,N_13664);
and U13955 (N_13955,N_13704,N_13784);
or U13956 (N_13956,N_13728,N_13683);
nor U13957 (N_13957,N_13724,N_13735);
xnor U13958 (N_13958,N_13672,N_13645);
nor U13959 (N_13959,N_13655,N_13710);
and U13960 (N_13960,N_13733,N_13774);
nor U13961 (N_13961,N_13758,N_13620);
nor U13962 (N_13962,N_13712,N_13683);
xnor U13963 (N_13963,N_13782,N_13772);
nor U13964 (N_13964,N_13797,N_13739);
xor U13965 (N_13965,N_13748,N_13654);
xnor U13966 (N_13966,N_13636,N_13686);
and U13967 (N_13967,N_13656,N_13640);
nand U13968 (N_13968,N_13788,N_13781);
or U13969 (N_13969,N_13608,N_13690);
nand U13970 (N_13970,N_13635,N_13769);
and U13971 (N_13971,N_13640,N_13721);
nand U13972 (N_13972,N_13639,N_13653);
nand U13973 (N_13973,N_13752,N_13769);
xnor U13974 (N_13974,N_13655,N_13752);
or U13975 (N_13975,N_13785,N_13766);
nor U13976 (N_13976,N_13740,N_13725);
or U13977 (N_13977,N_13621,N_13770);
or U13978 (N_13978,N_13766,N_13659);
xnor U13979 (N_13979,N_13799,N_13635);
or U13980 (N_13980,N_13680,N_13695);
xor U13981 (N_13981,N_13778,N_13633);
nand U13982 (N_13982,N_13785,N_13682);
nor U13983 (N_13983,N_13775,N_13617);
or U13984 (N_13984,N_13798,N_13723);
xor U13985 (N_13985,N_13668,N_13640);
or U13986 (N_13986,N_13651,N_13745);
xnor U13987 (N_13987,N_13640,N_13607);
nor U13988 (N_13988,N_13704,N_13735);
and U13989 (N_13989,N_13674,N_13746);
nor U13990 (N_13990,N_13640,N_13755);
or U13991 (N_13991,N_13738,N_13778);
nor U13992 (N_13992,N_13724,N_13656);
xnor U13993 (N_13993,N_13787,N_13784);
nor U13994 (N_13994,N_13756,N_13746);
nand U13995 (N_13995,N_13751,N_13763);
xor U13996 (N_13996,N_13718,N_13780);
xnor U13997 (N_13997,N_13698,N_13644);
xor U13998 (N_13998,N_13768,N_13763);
nand U13999 (N_13999,N_13655,N_13618);
or U14000 (N_14000,N_13993,N_13907);
nor U14001 (N_14001,N_13802,N_13990);
and U14002 (N_14002,N_13882,N_13962);
or U14003 (N_14003,N_13933,N_13847);
and U14004 (N_14004,N_13924,N_13816);
and U14005 (N_14005,N_13838,N_13929);
nor U14006 (N_14006,N_13862,N_13869);
nor U14007 (N_14007,N_13958,N_13941);
nor U14008 (N_14008,N_13982,N_13926);
or U14009 (N_14009,N_13983,N_13956);
or U14010 (N_14010,N_13999,N_13881);
and U14011 (N_14011,N_13935,N_13970);
xor U14012 (N_14012,N_13866,N_13953);
or U14013 (N_14013,N_13966,N_13917);
xnor U14014 (N_14014,N_13837,N_13895);
or U14015 (N_14015,N_13844,N_13828);
nand U14016 (N_14016,N_13826,N_13855);
xor U14017 (N_14017,N_13942,N_13850);
xnor U14018 (N_14018,N_13871,N_13987);
or U14019 (N_14019,N_13873,N_13951);
and U14020 (N_14020,N_13812,N_13867);
nor U14021 (N_14021,N_13938,N_13893);
and U14022 (N_14022,N_13872,N_13911);
nand U14023 (N_14023,N_13884,N_13876);
xnor U14024 (N_14024,N_13860,N_13902);
nand U14025 (N_14025,N_13883,N_13868);
xnor U14026 (N_14026,N_13963,N_13814);
and U14027 (N_14027,N_13810,N_13843);
and U14028 (N_14028,N_13848,N_13842);
xor U14029 (N_14029,N_13880,N_13908);
nor U14030 (N_14030,N_13825,N_13940);
or U14031 (N_14031,N_13934,N_13879);
nand U14032 (N_14032,N_13964,N_13813);
nand U14033 (N_14033,N_13968,N_13955);
and U14034 (N_14034,N_13913,N_13853);
xor U14035 (N_14035,N_13833,N_13891);
nand U14036 (N_14036,N_13985,N_13841);
and U14037 (N_14037,N_13887,N_13928);
xor U14038 (N_14038,N_13950,N_13801);
xnor U14039 (N_14039,N_13840,N_13975);
nor U14040 (N_14040,N_13849,N_13910);
xnor U14041 (N_14041,N_13827,N_13889);
or U14042 (N_14042,N_13992,N_13890);
nand U14043 (N_14043,N_13945,N_13896);
nor U14044 (N_14044,N_13846,N_13894);
or U14045 (N_14045,N_13952,N_13998);
nor U14046 (N_14046,N_13888,N_13905);
and U14047 (N_14047,N_13818,N_13996);
and U14048 (N_14048,N_13976,N_13803);
nand U14049 (N_14049,N_13949,N_13925);
nor U14050 (N_14050,N_13892,N_13874);
and U14051 (N_14051,N_13912,N_13977);
or U14052 (N_14052,N_13815,N_13832);
and U14053 (N_14053,N_13967,N_13865);
or U14054 (N_14054,N_13906,N_13973);
nor U14055 (N_14055,N_13984,N_13980);
xnor U14056 (N_14056,N_13918,N_13909);
or U14057 (N_14057,N_13824,N_13919);
or U14058 (N_14058,N_13834,N_13819);
nor U14059 (N_14059,N_13821,N_13947);
nand U14060 (N_14060,N_13800,N_13978);
and U14061 (N_14061,N_13807,N_13948);
nor U14062 (N_14062,N_13930,N_13936);
nand U14063 (N_14063,N_13831,N_13914);
nand U14064 (N_14064,N_13823,N_13878);
xnor U14065 (N_14065,N_13957,N_13989);
xor U14066 (N_14066,N_13870,N_13904);
and U14067 (N_14067,N_13851,N_13817);
xnor U14068 (N_14068,N_13885,N_13994);
nor U14069 (N_14069,N_13971,N_13901);
or U14070 (N_14070,N_13830,N_13820);
or U14071 (N_14071,N_13857,N_13898);
nor U14072 (N_14072,N_13923,N_13986);
xor U14073 (N_14073,N_13959,N_13979);
and U14074 (N_14074,N_13864,N_13916);
and U14075 (N_14075,N_13954,N_13809);
and U14076 (N_14076,N_13939,N_13877);
xor U14077 (N_14077,N_13805,N_13835);
and U14078 (N_14078,N_13981,N_13856);
nand U14079 (N_14079,N_13961,N_13946);
nor U14080 (N_14080,N_13811,N_13969);
nand U14081 (N_14081,N_13858,N_13900);
and U14082 (N_14082,N_13804,N_13927);
nor U14083 (N_14083,N_13995,N_13965);
nor U14084 (N_14084,N_13937,N_13854);
or U14085 (N_14085,N_13931,N_13997);
nor U14086 (N_14086,N_13960,N_13897);
nor U14087 (N_14087,N_13921,N_13899);
nand U14088 (N_14088,N_13922,N_13852);
or U14089 (N_14089,N_13875,N_13836);
nand U14090 (N_14090,N_13863,N_13988);
nor U14091 (N_14091,N_13861,N_13991);
or U14092 (N_14092,N_13829,N_13920);
and U14093 (N_14093,N_13859,N_13932);
xor U14094 (N_14094,N_13806,N_13974);
nor U14095 (N_14095,N_13822,N_13972);
nand U14096 (N_14096,N_13886,N_13839);
nand U14097 (N_14097,N_13915,N_13845);
nor U14098 (N_14098,N_13944,N_13903);
nand U14099 (N_14099,N_13943,N_13808);
nor U14100 (N_14100,N_13954,N_13826);
nor U14101 (N_14101,N_13874,N_13873);
nand U14102 (N_14102,N_13919,N_13855);
nor U14103 (N_14103,N_13812,N_13813);
nand U14104 (N_14104,N_13858,N_13930);
nand U14105 (N_14105,N_13982,N_13875);
nor U14106 (N_14106,N_13971,N_13973);
nor U14107 (N_14107,N_13881,N_13955);
xor U14108 (N_14108,N_13871,N_13957);
nand U14109 (N_14109,N_13857,N_13967);
nand U14110 (N_14110,N_13828,N_13943);
xor U14111 (N_14111,N_13832,N_13897);
xnor U14112 (N_14112,N_13933,N_13915);
or U14113 (N_14113,N_13989,N_13879);
or U14114 (N_14114,N_13958,N_13993);
nor U14115 (N_14115,N_13838,N_13994);
and U14116 (N_14116,N_13961,N_13991);
nand U14117 (N_14117,N_13884,N_13861);
xnor U14118 (N_14118,N_13990,N_13889);
xnor U14119 (N_14119,N_13913,N_13824);
nor U14120 (N_14120,N_13962,N_13983);
xnor U14121 (N_14121,N_13934,N_13935);
nand U14122 (N_14122,N_13856,N_13971);
xnor U14123 (N_14123,N_13807,N_13932);
or U14124 (N_14124,N_13940,N_13934);
xnor U14125 (N_14125,N_13822,N_13919);
nor U14126 (N_14126,N_13846,N_13859);
xor U14127 (N_14127,N_13861,N_13916);
or U14128 (N_14128,N_13921,N_13818);
and U14129 (N_14129,N_13903,N_13864);
nand U14130 (N_14130,N_13891,N_13825);
and U14131 (N_14131,N_13974,N_13926);
nand U14132 (N_14132,N_13866,N_13899);
nand U14133 (N_14133,N_13996,N_13943);
xnor U14134 (N_14134,N_13999,N_13944);
and U14135 (N_14135,N_13939,N_13878);
or U14136 (N_14136,N_13973,N_13845);
and U14137 (N_14137,N_13827,N_13956);
nand U14138 (N_14138,N_13907,N_13895);
nand U14139 (N_14139,N_13895,N_13960);
nand U14140 (N_14140,N_13875,N_13860);
nand U14141 (N_14141,N_13879,N_13811);
and U14142 (N_14142,N_13804,N_13822);
xor U14143 (N_14143,N_13896,N_13881);
and U14144 (N_14144,N_13994,N_13942);
nand U14145 (N_14145,N_13861,N_13879);
xnor U14146 (N_14146,N_13976,N_13808);
and U14147 (N_14147,N_13913,N_13940);
or U14148 (N_14148,N_13944,N_13921);
and U14149 (N_14149,N_13921,N_13923);
nor U14150 (N_14150,N_13928,N_13822);
or U14151 (N_14151,N_13950,N_13884);
xor U14152 (N_14152,N_13994,N_13989);
nor U14153 (N_14153,N_13840,N_13835);
or U14154 (N_14154,N_13881,N_13906);
nand U14155 (N_14155,N_13852,N_13912);
and U14156 (N_14156,N_13900,N_13802);
nand U14157 (N_14157,N_13899,N_13991);
or U14158 (N_14158,N_13853,N_13904);
nand U14159 (N_14159,N_13864,N_13929);
nand U14160 (N_14160,N_13819,N_13961);
xor U14161 (N_14161,N_13824,N_13834);
and U14162 (N_14162,N_13923,N_13822);
nand U14163 (N_14163,N_13878,N_13971);
nor U14164 (N_14164,N_13841,N_13852);
xnor U14165 (N_14165,N_13980,N_13836);
and U14166 (N_14166,N_13896,N_13852);
and U14167 (N_14167,N_13878,N_13956);
and U14168 (N_14168,N_13812,N_13835);
nor U14169 (N_14169,N_13980,N_13867);
and U14170 (N_14170,N_13952,N_13939);
xor U14171 (N_14171,N_13816,N_13995);
nand U14172 (N_14172,N_13917,N_13842);
and U14173 (N_14173,N_13982,N_13909);
nand U14174 (N_14174,N_13998,N_13846);
xnor U14175 (N_14175,N_13954,N_13884);
nor U14176 (N_14176,N_13955,N_13879);
or U14177 (N_14177,N_13833,N_13834);
nor U14178 (N_14178,N_13954,N_13867);
nand U14179 (N_14179,N_13855,N_13969);
nand U14180 (N_14180,N_13983,N_13979);
or U14181 (N_14181,N_13817,N_13821);
xnor U14182 (N_14182,N_13978,N_13864);
xor U14183 (N_14183,N_13936,N_13805);
nand U14184 (N_14184,N_13855,N_13952);
xnor U14185 (N_14185,N_13909,N_13936);
nor U14186 (N_14186,N_13819,N_13892);
nand U14187 (N_14187,N_13926,N_13881);
xnor U14188 (N_14188,N_13967,N_13975);
or U14189 (N_14189,N_13982,N_13968);
nand U14190 (N_14190,N_13988,N_13852);
xor U14191 (N_14191,N_13990,N_13971);
and U14192 (N_14192,N_13815,N_13937);
nand U14193 (N_14193,N_13970,N_13928);
nor U14194 (N_14194,N_13854,N_13848);
xor U14195 (N_14195,N_13919,N_13856);
nor U14196 (N_14196,N_13847,N_13990);
nor U14197 (N_14197,N_13957,N_13975);
and U14198 (N_14198,N_13804,N_13919);
and U14199 (N_14199,N_13978,N_13975);
nor U14200 (N_14200,N_14189,N_14195);
nor U14201 (N_14201,N_14091,N_14060);
and U14202 (N_14202,N_14150,N_14049);
or U14203 (N_14203,N_14088,N_14117);
nor U14204 (N_14204,N_14156,N_14092);
nor U14205 (N_14205,N_14170,N_14187);
nand U14206 (N_14206,N_14120,N_14101);
and U14207 (N_14207,N_14137,N_14163);
or U14208 (N_14208,N_14002,N_14062);
nor U14209 (N_14209,N_14109,N_14198);
nor U14210 (N_14210,N_14035,N_14005);
xnor U14211 (N_14211,N_14197,N_14016);
nand U14212 (N_14212,N_14131,N_14051);
nor U14213 (N_14213,N_14124,N_14040);
xor U14214 (N_14214,N_14143,N_14007);
and U14215 (N_14215,N_14054,N_14075);
nand U14216 (N_14216,N_14173,N_14112);
nor U14217 (N_14217,N_14078,N_14145);
and U14218 (N_14218,N_14100,N_14108);
nor U14219 (N_14219,N_14011,N_14188);
nand U14220 (N_14220,N_14031,N_14154);
xor U14221 (N_14221,N_14063,N_14175);
nand U14222 (N_14222,N_14196,N_14118);
or U14223 (N_14223,N_14190,N_14179);
xor U14224 (N_14224,N_14020,N_14125);
nor U14225 (N_14225,N_14139,N_14013);
or U14226 (N_14226,N_14003,N_14164);
or U14227 (N_14227,N_14015,N_14162);
or U14228 (N_14228,N_14141,N_14183);
and U14229 (N_14229,N_14021,N_14113);
or U14230 (N_14230,N_14089,N_14138);
nor U14231 (N_14231,N_14064,N_14057);
nand U14232 (N_14232,N_14086,N_14014);
nand U14233 (N_14233,N_14025,N_14058);
nand U14234 (N_14234,N_14096,N_14001);
xor U14235 (N_14235,N_14110,N_14043);
xor U14236 (N_14236,N_14192,N_14056);
xor U14237 (N_14237,N_14152,N_14134);
nor U14238 (N_14238,N_14059,N_14023);
xor U14239 (N_14239,N_14099,N_14119);
nor U14240 (N_14240,N_14036,N_14055);
or U14241 (N_14241,N_14050,N_14147);
xnor U14242 (N_14242,N_14038,N_14133);
and U14243 (N_14243,N_14037,N_14144);
xor U14244 (N_14244,N_14066,N_14111);
nor U14245 (N_14245,N_14032,N_14177);
nand U14246 (N_14246,N_14068,N_14114);
or U14247 (N_14247,N_14142,N_14083);
nand U14248 (N_14248,N_14027,N_14082);
nand U14249 (N_14249,N_14130,N_14034);
and U14250 (N_14250,N_14123,N_14052);
nand U14251 (N_14251,N_14107,N_14182);
nand U14252 (N_14252,N_14073,N_14148);
and U14253 (N_14253,N_14181,N_14169);
xor U14254 (N_14254,N_14194,N_14171);
and U14255 (N_14255,N_14061,N_14199);
or U14256 (N_14256,N_14072,N_14185);
nand U14257 (N_14257,N_14071,N_14039);
nand U14258 (N_14258,N_14022,N_14041);
or U14259 (N_14259,N_14077,N_14176);
and U14260 (N_14260,N_14087,N_14172);
nor U14261 (N_14261,N_14004,N_14028);
nand U14262 (N_14262,N_14136,N_14121);
or U14263 (N_14263,N_14030,N_14074);
nand U14264 (N_14264,N_14009,N_14008);
and U14265 (N_14265,N_14157,N_14135);
nand U14266 (N_14266,N_14065,N_14084);
nor U14267 (N_14267,N_14186,N_14159);
nand U14268 (N_14268,N_14127,N_14178);
nand U14269 (N_14269,N_14048,N_14158);
nor U14270 (N_14270,N_14046,N_14006);
nor U14271 (N_14271,N_14151,N_14126);
or U14272 (N_14272,N_14161,N_14067);
nor U14273 (N_14273,N_14167,N_14081);
nor U14274 (N_14274,N_14079,N_14017);
or U14275 (N_14275,N_14069,N_14174);
and U14276 (N_14276,N_14103,N_14090);
or U14277 (N_14277,N_14026,N_14012);
nand U14278 (N_14278,N_14104,N_14033);
and U14279 (N_14279,N_14184,N_14160);
and U14280 (N_14280,N_14166,N_14153);
and U14281 (N_14281,N_14000,N_14149);
nand U14282 (N_14282,N_14047,N_14010);
nor U14283 (N_14283,N_14095,N_14122);
and U14284 (N_14284,N_14116,N_14132);
nand U14285 (N_14285,N_14042,N_14098);
or U14286 (N_14286,N_14094,N_14076);
or U14287 (N_14287,N_14070,N_14097);
xnor U14288 (N_14288,N_14044,N_14165);
xnor U14289 (N_14289,N_14140,N_14146);
and U14290 (N_14290,N_14155,N_14193);
or U14291 (N_14291,N_14024,N_14093);
or U14292 (N_14292,N_14019,N_14128);
xor U14293 (N_14293,N_14045,N_14105);
xor U14294 (N_14294,N_14191,N_14085);
nor U14295 (N_14295,N_14029,N_14102);
or U14296 (N_14296,N_14018,N_14106);
nand U14297 (N_14297,N_14080,N_14168);
nand U14298 (N_14298,N_14129,N_14053);
nand U14299 (N_14299,N_14180,N_14115);
xor U14300 (N_14300,N_14168,N_14102);
or U14301 (N_14301,N_14148,N_14186);
nor U14302 (N_14302,N_14127,N_14166);
xnor U14303 (N_14303,N_14177,N_14055);
nor U14304 (N_14304,N_14118,N_14128);
nand U14305 (N_14305,N_14024,N_14159);
nand U14306 (N_14306,N_14009,N_14138);
nand U14307 (N_14307,N_14097,N_14055);
nand U14308 (N_14308,N_14019,N_14145);
or U14309 (N_14309,N_14046,N_14084);
xnor U14310 (N_14310,N_14175,N_14099);
xor U14311 (N_14311,N_14190,N_14127);
nor U14312 (N_14312,N_14138,N_14155);
and U14313 (N_14313,N_14103,N_14017);
or U14314 (N_14314,N_14143,N_14071);
xor U14315 (N_14315,N_14102,N_14057);
nor U14316 (N_14316,N_14036,N_14019);
nor U14317 (N_14317,N_14056,N_14064);
and U14318 (N_14318,N_14133,N_14112);
nand U14319 (N_14319,N_14026,N_14089);
or U14320 (N_14320,N_14014,N_14005);
and U14321 (N_14321,N_14166,N_14077);
nor U14322 (N_14322,N_14070,N_14030);
nor U14323 (N_14323,N_14180,N_14017);
and U14324 (N_14324,N_14099,N_14036);
nor U14325 (N_14325,N_14095,N_14199);
or U14326 (N_14326,N_14190,N_14065);
nor U14327 (N_14327,N_14000,N_14034);
xnor U14328 (N_14328,N_14022,N_14066);
or U14329 (N_14329,N_14184,N_14194);
nand U14330 (N_14330,N_14090,N_14146);
or U14331 (N_14331,N_14070,N_14023);
xnor U14332 (N_14332,N_14171,N_14196);
nor U14333 (N_14333,N_14160,N_14139);
nor U14334 (N_14334,N_14064,N_14103);
or U14335 (N_14335,N_14171,N_14152);
xnor U14336 (N_14336,N_14183,N_14032);
xnor U14337 (N_14337,N_14163,N_14119);
nor U14338 (N_14338,N_14168,N_14116);
and U14339 (N_14339,N_14090,N_14051);
and U14340 (N_14340,N_14010,N_14039);
or U14341 (N_14341,N_14033,N_14019);
nor U14342 (N_14342,N_14057,N_14137);
xnor U14343 (N_14343,N_14023,N_14179);
nor U14344 (N_14344,N_14145,N_14096);
and U14345 (N_14345,N_14023,N_14143);
or U14346 (N_14346,N_14024,N_14091);
or U14347 (N_14347,N_14074,N_14147);
and U14348 (N_14348,N_14152,N_14088);
nand U14349 (N_14349,N_14030,N_14000);
or U14350 (N_14350,N_14060,N_14150);
and U14351 (N_14351,N_14154,N_14163);
or U14352 (N_14352,N_14084,N_14029);
nand U14353 (N_14353,N_14107,N_14178);
and U14354 (N_14354,N_14079,N_14144);
nor U14355 (N_14355,N_14003,N_14125);
nor U14356 (N_14356,N_14047,N_14060);
xnor U14357 (N_14357,N_14002,N_14109);
and U14358 (N_14358,N_14074,N_14033);
xor U14359 (N_14359,N_14191,N_14196);
xnor U14360 (N_14360,N_14199,N_14193);
nand U14361 (N_14361,N_14076,N_14114);
and U14362 (N_14362,N_14173,N_14168);
nand U14363 (N_14363,N_14119,N_14053);
and U14364 (N_14364,N_14057,N_14007);
or U14365 (N_14365,N_14122,N_14146);
nor U14366 (N_14366,N_14002,N_14003);
or U14367 (N_14367,N_14148,N_14014);
nand U14368 (N_14368,N_14046,N_14197);
or U14369 (N_14369,N_14012,N_14068);
nor U14370 (N_14370,N_14105,N_14138);
nor U14371 (N_14371,N_14190,N_14001);
or U14372 (N_14372,N_14022,N_14142);
and U14373 (N_14373,N_14114,N_14074);
nand U14374 (N_14374,N_14185,N_14006);
xnor U14375 (N_14375,N_14129,N_14094);
nand U14376 (N_14376,N_14085,N_14197);
and U14377 (N_14377,N_14005,N_14033);
nor U14378 (N_14378,N_14037,N_14090);
or U14379 (N_14379,N_14028,N_14129);
nand U14380 (N_14380,N_14061,N_14138);
or U14381 (N_14381,N_14084,N_14144);
and U14382 (N_14382,N_14000,N_14104);
nand U14383 (N_14383,N_14199,N_14136);
nor U14384 (N_14384,N_14046,N_14186);
nor U14385 (N_14385,N_14156,N_14142);
or U14386 (N_14386,N_14162,N_14123);
nor U14387 (N_14387,N_14007,N_14011);
nand U14388 (N_14388,N_14045,N_14168);
nand U14389 (N_14389,N_14166,N_14083);
nor U14390 (N_14390,N_14101,N_14110);
nor U14391 (N_14391,N_14118,N_14121);
nand U14392 (N_14392,N_14129,N_14008);
or U14393 (N_14393,N_14028,N_14157);
nand U14394 (N_14394,N_14167,N_14066);
nand U14395 (N_14395,N_14181,N_14026);
nand U14396 (N_14396,N_14141,N_14123);
and U14397 (N_14397,N_14022,N_14013);
nor U14398 (N_14398,N_14147,N_14076);
nand U14399 (N_14399,N_14052,N_14006);
or U14400 (N_14400,N_14383,N_14298);
and U14401 (N_14401,N_14264,N_14246);
xor U14402 (N_14402,N_14377,N_14206);
and U14403 (N_14403,N_14249,N_14292);
nor U14404 (N_14404,N_14324,N_14222);
nand U14405 (N_14405,N_14336,N_14333);
or U14406 (N_14406,N_14396,N_14301);
or U14407 (N_14407,N_14245,N_14229);
nor U14408 (N_14408,N_14327,N_14265);
nand U14409 (N_14409,N_14274,N_14204);
or U14410 (N_14410,N_14235,N_14314);
xnor U14411 (N_14411,N_14268,N_14275);
or U14412 (N_14412,N_14369,N_14323);
and U14413 (N_14413,N_14375,N_14300);
or U14414 (N_14414,N_14328,N_14390);
nand U14415 (N_14415,N_14283,N_14207);
or U14416 (N_14416,N_14370,N_14242);
xor U14417 (N_14417,N_14337,N_14286);
and U14418 (N_14418,N_14209,N_14287);
and U14419 (N_14419,N_14271,N_14281);
or U14420 (N_14420,N_14344,N_14308);
or U14421 (N_14421,N_14341,N_14355);
nor U14422 (N_14422,N_14272,N_14215);
nor U14423 (N_14423,N_14267,N_14243);
and U14424 (N_14424,N_14358,N_14312);
or U14425 (N_14425,N_14241,N_14247);
xor U14426 (N_14426,N_14213,N_14391);
nand U14427 (N_14427,N_14334,N_14293);
or U14428 (N_14428,N_14397,N_14295);
nand U14429 (N_14429,N_14384,N_14294);
or U14430 (N_14430,N_14342,N_14348);
and U14431 (N_14431,N_14279,N_14262);
and U14432 (N_14432,N_14255,N_14201);
nor U14433 (N_14433,N_14231,N_14357);
or U14434 (N_14434,N_14304,N_14319);
or U14435 (N_14435,N_14368,N_14220);
or U14436 (N_14436,N_14309,N_14311);
nor U14437 (N_14437,N_14261,N_14394);
nor U14438 (N_14438,N_14374,N_14310);
xor U14439 (N_14439,N_14260,N_14343);
and U14440 (N_14440,N_14228,N_14307);
nor U14441 (N_14441,N_14282,N_14366);
nand U14442 (N_14442,N_14296,N_14356);
nand U14443 (N_14443,N_14305,N_14392);
nor U14444 (N_14444,N_14259,N_14339);
nand U14445 (N_14445,N_14338,N_14353);
nor U14446 (N_14446,N_14322,N_14306);
nor U14447 (N_14447,N_14302,N_14257);
and U14448 (N_14448,N_14335,N_14393);
or U14449 (N_14449,N_14297,N_14239);
and U14450 (N_14450,N_14225,N_14252);
or U14451 (N_14451,N_14365,N_14233);
or U14452 (N_14452,N_14250,N_14278);
or U14453 (N_14453,N_14238,N_14321);
xnor U14454 (N_14454,N_14326,N_14237);
or U14455 (N_14455,N_14212,N_14360);
nand U14456 (N_14456,N_14254,N_14329);
and U14457 (N_14457,N_14218,N_14236);
nor U14458 (N_14458,N_14315,N_14253);
nor U14459 (N_14459,N_14219,N_14351);
nor U14460 (N_14460,N_14349,N_14389);
or U14461 (N_14461,N_14270,N_14320);
nor U14462 (N_14462,N_14280,N_14227);
nand U14463 (N_14463,N_14385,N_14291);
nand U14464 (N_14464,N_14203,N_14362);
nor U14465 (N_14465,N_14367,N_14210);
or U14466 (N_14466,N_14202,N_14361);
nand U14467 (N_14467,N_14288,N_14289);
nor U14468 (N_14468,N_14380,N_14224);
xor U14469 (N_14469,N_14216,N_14317);
nand U14470 (N_14470,N_14303,N_14316);
and U14471 (N_14471,N_14232,N_14256);
nand U14472 (N_14472,N_14234,N_14226);
and U14473 (N_14473,N_14251,N_14346);
nand U14474 (N_14474,N_14290,N_14285);
xor U14475 (N_14475,N_14379,N_14387);
and U14476 (N_14476,N_14359,N_14284);
nor U14477 (N_14477,N_14340,N_14350);
nor U14478 (N_14478,N_14221,N_14330);
nand U14479 (N_14479,N_14376,N_14381);
nor U14480 (N_14480,N_14248,N_14208);
nand U14481 (N_14481,N_14354,N_14217);
nor U14482 (N_14482,N_14347,N_14258);
and U14483 (N_14483,N_14230,N_14372);
nand U14484 (N_14484,N_14398,N_14386);
or U14485 (N_14485,N_14378,N_14276);
nor U14486 (N_14486,N_14277,N_14331);
nand U14487 (N_14487,N_14332,N_14299);
or U14488 (N_14488,N_14266,N_14240);
nor U14489 (N_14489,N_14371,N_14244);
or U14490 (N_14490,N_14364,N_14363);
or U14491 (N_14491,N_14214,N_14211);
xor U14492 (N_14492,N_14273,N_14325);
nand U14493 (N_14493,N_14200,N_14345);
nand U14494 (N_14494,N_14373,N_14352);
nand U14495 (N_14495,N_14388,N_14313);
nand U14496 (N_14496,N_14269,N_14223);
and U14497 (N_14497,N_14399,N_14205);
and U14498 (N_14498,N_14382,N_14395);
nand U14499 (N_14499,N_14318,N_14263);
nor U14500 (N_14500,N_14300,N_14322);
and U14501 (N_14501,N_14311,N_14371);
nand U14502 (N_14502,N_14265,N_14237);
nand U14503 (N_14503,N_14212,N_14352);
nor U14504 (N_14504,N_14283,N_14363);
and U14505 (N_14505,N_14262,N_14284);
nor U14506 (N_14506,N_14262,N_14363);
nand U14507 (N_14507,N_14297,N_14290);
nand U14508 (N_14508,N_14381,N_14334);
or U14509 (N_14509,N_14226,N_14374);
or U14510 (N_14510,N_14395,N_14265);
nor U14511 (N_14511,N_14241,N_14328);
xor U14512 (N_14512,N_14319,N_14277);
xnor U14513 (N_14513,N_14309,N_14217);
xnor U14514 (N_14514,N_14329,N_14345);
or U14515 (N_14515,N_14370,N_14258);
and U14516 (N_14516,N_14256,N_14296);
or U14517 (N_14517,N_14272,N_14231);
nand U14518 (N_14518,N_14229,N_14228);
and U14519 (N_14519,N_14210,N_14324);
xor U14520 (N_14520,N_14312,N_14394);
and U14521 (N_14521,N_14307,N_14393);
and U14522 (N_14522,N_14240,N_14249);
nor U14523 (N_14523,N_14375,N_14279);
or U14524 (N_14524,N_14342,N_14384);
xor U14525 (N_14525,N_14395,N_14250);
nand U14526 (N_14526,N_14304,N_14264);
and U14527 (N_14527,N_14343,N_14326);
nand U14528 (N_14528,N_14256,N_14251);
xor U14529 (N_14529,N_14287,N_14343);
nand U14530 (N_14530,N_14308,N_14213);
nor U14531 (N_14531,N_14375,N_14244);
or U14532 (N_14532,N_14338,N_14207);
or U14533 (N_14533,N_14372,N_14215);
nand U14534 (N_14534,N_14228,N_14349);
and U14535 (N_14535,N_14242,N_14336);
or U14536 (N_14536,N_14333,N_14235);
or U14537 (N_14537,N_14265,N_14258);
xor U14538 (N_14538,N_14305,N_14270);
nand U14539 (N_14539,N_14267,N_14384);
xor U14540 (N_14540,N_14291,N_14345);
or U14541 (N_14541,N_14219,N_14229);
nor U14542 (N_14542,N_14260,N_14269);
and U14543 (N_14543,N_14339,N_14242);
xor U14544 (N_14544,N_14236,N_14379);
or U14545 (N_14545,N_14271,N_14251);
or U14546 (N_14546,N_14265,N_14235);
nand U14547 (N_14547,N_14275,N_14317);
nor U14548 (N_14548,N_14238,N_14329);
xnor U14549 (N_14549,N_14392,N_14275);
nand U14550 (N_14550,N_14237,N_14270);
nor U14551 (N_14551,N_14288,N_14279);
or U14552 (N_14552,N_14276,N_14237);
xor U14553 (N_14553,N_14275,N_14339);
nor U14554 (N_14554,N_14371,N_14326);
or U14555 (N_14555,N_14237,N_14325);
nor U14556 (N_14556,N_14343,N_14324);
or U14557 (N_14557,N_14205,N_14204);
or U14558 (N_14558,N_14386,N_14325);
and U14559 (N_14559,N_14360,N_14290);
nor U14560 (N_14560,N_14304,N_14349);
nand U14561 (N_14561,N_14202,N_14284);
and U14562 (N_14562,N_14231,N_14285);
and U14563 (N_14563,N_14369,N_14334);
nor U14564 (N_14564,N_14265,N_14303);
nand U14565 (N_14565,N_14230,N_14277);
nor U14566 (N_14566,N_14371,N_14272);
xnor U14567 (N_14567,N_14216,N_14354);
nand U14568 (N_14568,N_14256,N_14230);
nor U14569 (N_14569,N_14361,N_14311);
xnor U14570 (N_14570,N_14330,N_14309);
nand U14571 (N_14571,N_14213,N_14320);
xor U14572 (N_14572,N_14247,N_14335);
nor U14573 (N_14573,N_14345,N_14365);
or U14574 (N_14574,N_14248,N_14245);
nor U14575 (N_14575,N_14253,N_14356);
xnor U14576 (N_14576,N_14240,N_14229);
or U14577 (N_14577,N_14347,N_14252);
nand U14578 (N_14578,N_14267,N_14263);
or U14579 (N_14579,N_14336,N_14219);
xor U14580 (N_14580,N_14330,N_14286);
and U14581 (N_14581,N_14259,N_14327);
nor U14582 (N_14582,N_14331,N_14286);
or U14583 (N_14583,N_14385,N_14314);
or U14584 (N_14584,N_14226,N_14356);
nand U14585 (N_14585,N_14274,N_14261);
or U14586 (N_14586,N_14201,N_14350);
and U14587 (N_14587,N_14331,N_14363);
and U14588 (N_14588,N_14385,N_14267);
xnor U14589 (N_14589,N_14207,N_14382);
nand U14590 (N_14590,N_14290,N_14316);
nor U14591 (N_14591,N_14354,N_14203);
nor U14592 (N_14592,N_14367,N_14217);
xor U14593 (N_14593,N_14399,N_14336);
or U14594 (N_14594,N_14271,N_14299);
or U14595 (N_14595,N_14282,N_14251);
nor U14596 (N_14596,N_14323,N_14386);
xnor U14597 (N_14597,N_14366,N_14357);
nor U14598 (N_14598,N_14280,N_14233);
or U14599 (N_14599,N_14219,N_14299);
or U14600 (N_14600,N_14428,N_14569);
nand U14601 (N_14601,N_14586,N_14490);
nor U14602 (N_14602,N_14545,N_14474);
xnor U14603 (N_14603,N_14531,N_14424);
nand U14604 (N_14604,N_14447,N_14570);
nand U14605 (N_14605,N_14469,N_14440);
or U14606 (N_14606,N_14519,N_14568);
and U14607 (N_14607,N_14465,N_14438);
or U14608 (N_14608,N_14567,N_14470);
nand U14609 (N_14609,N_14496,N_14429);
nor U14610 (N_14610,N_14425,N_14481);
nand U14611 (N_14611,N_14484,N_14485);
xor U14612 (N_14612,N_14506,N_14525);
nand U14613 (N_14613,N_14450,N_14467);
xnor U14614 (N_14614,N_14599,N_14571);
nor U14615 (N_14615,N_14435,N_14578);
or U14616 (N_14616,N_14463,N_14594);
and U14617 (N_14617,N_14451,N_14493);
or U14618 (N_14618,N_14524,N_14558);
or U14619 (N_14619,N_14588,N_14596);
and U14620 (N_14620,N_14403,N_14529);
and U14621 (N_14621,N_14576,N_14582);
and U14622 (N_14622,N_14457,N_14556);
nor U14623 (N_14623,N_14537,N_14412);
and U14624 (N_14624,N_14411,N_14583);
nor U14625 (N_14625,N_14509,N_14553);
and U14626 (N_14626,N_14595,N_14446);
and U14627 (N_14627,N_14495,N_14400);
nor U14628 (N_14628,N_14422,N_14515);
nand U14629 (N_14629,N_14557,N_14504);
xor U14630 (N_14630,N_14533,N_14540);
and U14631 (N_14631,N_14552,N_14575);
xnor U14632 (N_14632,N_14511,N_14458);
xnor U14633 (N_14633,N_14514,N_14502);
nor U14634 (N_14634,N_14454,N_14407);
nor U14635 (N_14635,N_14418,N_14544);
or U14636 (N_14636,N_14473,N_14536);
nor U14637 (N_14637,N_14518,N_14408);
xnor U14638 (N_14638,N_14406,N_14579);
or U14639 (N_14639,N_14471,N_14449);
nor U14640 (N_14640,N_14409,N_14573);
or U14641 (N_14641,N_14415,N_14443);
and U14642 (N_14642,N_14487,N_14436);
xor U14643 (N_14643,N_14420,N_14431);
nand U14644 (N_14644,N_14483,N_14442);
and U14645 (N_14645,N_14584,N_14534);
nand U14646 (N_14646,N_14563,N_14445);
or U14647 (N_14647,N_14414,N_14572);
xnor U14648 (N_14648,N_14419,N_14551);
nand U14649 (N_14649,N_14426,N_14548);
nand U14650 (N_14650,N_14517,N_14455);
or U14651 (N_14651,N_14591,N_14538);
nor U14652 (N_14652,N_14528,N_14503);
and U14653 (N_14653,N_14423,N_14521);
nor U14654 (N_14654,N_14494,N_14541);
nor U14655 (N_14655,N_14432,N_14546);
nand U14656 (N_14656,N_14460,N_14430);
xnor U14657 (N_14657,N_14456,N_14492);
or U14658 (N_14658,N_14555,N_14535);
nor U14659 (N_14659,N_14489,N_14542);
and U14660 (N_14660,N_14479,N_14421);
xnor U14661 (N_14661,N_14427,N_14439);
xor U14662 (N_14662,N_14527,N_14461);
nor U14663 (N_14663,N_14402,N_14453);
xor U14664 (N_14664,N_14459,N_14561);
nor U14665 (N_14665,N_14480,N_14539);
nand U14666 (N_14666,N_14580,N_14416);
nor U14667 (N_14667,N_14472,N_14543);
nand U14668 (N_14668,N_14434,N_14433);
nand U14669 (N_14669,N_14532,N_14547);
nor U14670 (N_14670,N_14501,N_14452);
nor U14671 (N_14671,N_14565,N_14559);
nor U14672 (N_14672,N_14508,N_14417);
or U14673 (N_14673,N_14513,N_14577);
and U14674 (N_14674,N_14505,N_14500);
or U14675 (N_14675,N_14549,N_14526);
nand U14676 (N_14676,N_14522,N_14478);
or U14677 (N_14677,N_14581,N_14468);
and U14678 (N_14678,N_14585,N_14550);
nand U14679 (N_14679,N_14462,N_14593);
nor U14680 (N_14680,N_14444,N_14592);
xor U14681 (N_14681,N_14589,N_14560);
or U14682 (N_14682,N_14404,N_14523);
xnor U14683 (N_14683,N_14497,N_14564);
or U14684 (N_14684,N_14516,N_14488);
nor U14685 (N_14685,N_14476,N_14510);
nand U14686 (N_14686,N_14499,N_14590);
and U14687 (N_14687,N_14410,N_14498);
or U14688 (N_14688,N_14491,N_14486);
nand U14689 (N_14689,N_14562,N_14405);
nand U14690 (N_14690,N_14554,N_14466);
or U14691 (N_14691,N_14530,N_14441);
nor U14692 (N_14692,N_14574,N_14448);
xor U14693 (N_14693,N_14597,N_14566);
xor U14694 (N_14694,N_14520,N_14401);
or U14695 (N_14695,N_14464,N_14482);
nand U14696 (N_14696,N_14507,N_14413);
nor U14697 (N_14697,N_14437,N_14587);
and U14698 (N_14698,N_14512,N_14598);
or U14699 (N_14699,N_14475,N_14477);
and U14700 (N_14700,N_14574,N_14599);
nor U14701 (N_14701,N_14453,N_14488);
nor U14702 (N_14702,N_14558,N_14585);
nor U14703 (N_14703,N_14562,N_14480);
or U14704 (N_14704,N_14412,N_14465);
nand U14705 (N_14705,N_14437,N_14453);
nand U14706 (N_14706,N_14565,N_14443);
xor U14707 (N_14707,N_14581,N_14405);
or U14708 (N_14708,N_14416,N_14501);
or U14709 (N_14709,N_14443,N_14442);
nand U14710 (N_14710,N_14493,N_14536);
nand U14711 (N_14711,N_14435,N_14480);
and U14712 (N_14712,N_14530,N_14444);
or U14713 (N_14713,N_14530,N_14528);
nand U14714 (N_14714,N_14466,N_14519);
nor U14715 (N_14715,N_14484,N_14403);
xor U14716 (N_14716,N_14597,N_14531);
nor U14717 (N_14717,N_14518,N_14513);
xor U14718 (N_14718,N_14530,N_14404);
and U14719 (N_14719,N_14415,N_14477);
nand U14720 (N_14720,N_14557,N_14573);
nand U14721 (N_14721,N_14557,N_14587);
xor U14722 (N_14722,N_14455,N_14566);
or U14723 (N_14723,N_14529,N_14502);
or U14724 (N_14724,N_14476,N_14451);
nand U14725 (N_14725,N_14527,N_14548);
nand U14726 (N_14726,N_14570,N_14439);
nor U14727 (N_14727,N_14473,N_14582);
nand U14728 (N_14728,N_14559,N_14511);
nor U14729 (N_14729,N_14583,N_14559);
and U14730 (N_14730,N_14501,N_14408);
xnor U14731 (N_14731,N_14403,N_14426);
xor U14732 (N_14732,N_14528,N_14465);
and U14733 (N_14733,N_14511,N_14514);
or U14734 (N_14734,N_14433,N_14412);
xnor U14735 (N_14735,N_14569,N_14563);
nand U14736 (N_14736,N_14567,N_14527);
or U14737 (N_14737,N_14477,N_14554);
nand U14738 (N_14738,N_14512,N_14544);
or U14739 (N_14739,N_14557,N_14482);
nor U14740 (N_14740,N_14497,N_14525);
nand U14741 (N_14741,N_14507,N_14489);
nor U14742 (N_14742,N_14560,N_14590);
or U14743 (N_14743,N_14548,N_14504);
nor U14744 (N_14744,N_14524,N_14581);
nand U14745 (N_14745,N_14488,N_14529);
nor U14746 (N_14746,N_14558,N_14546);
nor U14747 (N_14747,N_14426,N_14493);
xnor U14748 (N_14748,N_14534,N_14538);
xor U14749 (N_14749,N_14467,N_14511);
and U14750 (N_14750,N_14465,N_14546);
nor U14751 (N_14751,N_14554,N_14412);
and U14752 (N_14752,N_14563,N_14586);
or U14753 (N_14753,N_14471,N_14501);
nand U14754 (N_14754,N_14453,N_14438);
nor U14755 (N_14755,N_14485,N_14573);
xor U14756 (N_14756,N_14468,N_14506);
or U14757 (N_14757,N_14470,N_14515);
and U14758 (N_14758,N_14589,N_14412);
or U14759 (N_14759,N_14556,N_14591);
xnor U14760 (N_14760,N_14512,N_14469);
nand U14761 (N_14761,N_14502,N_14518);
nand U14762 (N_14762,N_14592,N_14410);
nor U14763 (N_14763,N_14438,N_14446);
nor U14764 (N_14764,N_14506,N_14549);
xnor U14765 (N_14765,N_14539,N_14534);
and U14766 (N_14766,N_14477,N_14425);
xor U14767 (N_14767,N_14467,N_14413);
nand U14768 (N_14768,N_14507,N_14578);
nor U14769 (N_14769,N_14446,N_14456);
nand U14770 (N_14770,N_14530,N_14473);
and U14771 (N_14771,N_14490,N_14531);
nand U14772 (N_14772,N_14589,N_14463);
and U14773 (N_14773,N_14410,N_14455);
and U14774 (N_14774,N_14428,N_14551);
xor U14775 (N_14775,N_14437,N_14513);
and U14776 (N_14776,N_14572,N_14578);
xor U14777 (N_14777,N_14485,N_14589);
nand U14778 (N_14778,N_14448,N_14597);
xnor U14779 (N_14779,N_14436,N_14503);
xor U14780 (N_14780,N_14430,N_14558);
nor U14781 (N_14781,N_14442,N_14415);
nand U14782 (N_14782,N_14483,N_14446);
nand U14783 (N_14783,N_14491,N_14412);
nor U14784 (N_14784,N_14455,N_14438);
or U14785 (N_14785,N_14463,N_14420);
xnor U14786 (N_14786,N_14599,N_14402);
xnor U14787 (N_14787,N_14447,N_14418);
and U14788 (N_14788,N_14550,N_14423);
nand U14789 (N_14789,N_14418,N_14451);
and U14790 (N_14790,N_14452,N_14498);
and U14791 (N_14791,N_14490,N_14529);
nand U14792 (N_14792,N_14596,N_14531);
nand U14793 (N_14793,N_14515,N_14520);
nand U14794 (N_14794,N_14404,N_14449);
or U14795 (N_14795,N_14555,N_14588);
xnor U14796 (N_14796,N_14517,N_14449);
nor U14797 (N_14797,N_14571,N_14462);
or U14798 (N_14798,N_14490,N_14506);
nor U14799 (N_14799,N_14581,N_14469);
nand U14800 (N_14800,N_14735,N_14763);
nor U14801 (N_14801,N_14682,N_14639);
xnor U14802 (N_14802,N_14786,N_14664);
or U14803 (N_14803,N_14650,N_14680);
nand U14804 (N_14804,N_14630,N_14780);
nand U14805 (N_14805,N_14732,N_14728);
nor U14806 (N_14806,N_14758,N_14666);
and U14807 (N_14807,N_14603,N_14795);
or U14808 (N_14808,N_14742,N_14669);
and U14809 (N_14809,N_14624,N_14750);
xnor U14810 (N_14810,N_14695,N_14738);
nand U14811 (N_14811,N_14674,N_14710);
nand U14812 (N_14812,N_14611,N_14643);
or U14813 (N_14813,N_14770,N_14662);
nor U14814 (N_14814,N_14709,N_14661);
and U14815 (N_14815,N_14693,N_14702);
or U14816 (N_14816,N_14790,N_14657);
and U14817 (N_14817,N_14782,N_14607);
xnor U14818 (N_14818,N_14762,N_14604);
and U14819 (N_14819,N_14736,N_14656);
nor U14820 (N_14820,N_14733,N_14791);
nand U14821 (N_14821,N_14781,N_14606);
and U14822 (N_14822,N_14726,N_14783);
nor U14823 (N_14823,N_14687,N_14755);
nand U14824 (N_14824,N_14718,N_14765);
nor U14825 (N_14825,N_14772,N_14747);
or U14826 (N_14826,N_14760,N_14619);
xnor U14827 (N_14827,N_14794,N_14659);
and U14828 (N_14828,N_14745,N_14644);
xnor U14829 (N_14829,N_14731,N_14752);
and U14830 (N_14830,N_14667,N_14671);
and U14831 (N_14831,N_14730,N_14692);
and U14832 (N_14832,N_14640,N_14793);
nor U14833 (N_14833,N_14697,N_14608);
xor U14834 (N_14834,N_14746,N_14764);
nand U14835 (N_14835,N_14681,N_14645);
xnor U14836 (N_14836,N_14714,N_14668);
xor U14837 (N_14837,N_14642,N_14609);
nand U14838 (N_14838,N_14712,N_14721);
nand U14839 (N_14839,N_14734,N_14722);
nor U14840 (N_14840,N_14796,N_14756);
xor U14841 (N_14841,N_14727,N_14785);
or U14842 (N_14842,N_14672,N_14623);
xnor U14843 (N_14843,N_14663,N_14612);
nand U14844 (N_14844,N_14620,N_14774);
or U14845 (N_14845,N_14618,N_14778);
and U14846 (N_14846,N_14653,N_14789);
nor U14847 (N_14847,N_14696,N_14658);
xnor U14848 (N_14848,N_14632,N_14751);
xnor U14849 (N_14849,N_14629,N_14602);
nand U14850 (N_14850,N_14677,N_14719);
nand U14851 (N_14851,N_14799,N_14627);
and U14852 (N_14852,N_14690,N_14788);
xnor U14853 (N_14853,N_14665,N_14617);
xnor U14854 (N_14854,N_14787,N_14743);
xor U14855 (N_14855,N_14633,N_14683);
xnor U14856 (N_14856,N_14776,N_14757);
nor U14857 (N_14857,N_14647,N_14720);
nor U14858 (N_14858,N_14676,N_14614);
and U14859 (N_14859,N_14717,N_14768);
xnor U14860 (N_14860,N_14775,N_14753);
and U14861 (N_14861,N_14723,N_14626);
nor U14862 (N_14862,N_14673,N_14741);
nor U14863 (N_14863,N_14648,N_14601);
or U14864 (N_14864,N_14637,N_14649);
xor U14865 (N_14865,N_14704,N_14689);
or U14866 (N_14866,N_14740,N_14773);
or U14867 (N_14867,N_14622,N_14797);
xnor U14868 (N_14868,N_14749,N_14759);
nor U14869 (N_14869,N_14646,N_14635);
and U14870 (N_14870,N_14766,N_14685);
nor U14871 (N_14871,N_14655,N_14684);
xnor U14872 (N_14872,N_14703,N_14748);
or U14873 (N_14873,N_14784,N_14700);
or U14874 (N_14874,N_14678,N_14792);
nand U14875 (N_14875,N_14729,N_14701);
nor U14876 (N_14876,N_14725,N_14769);
nor U14877 (N_14877,N_14610,N_14715);
nor U14878 (N_14878,N_14641,N_14686);
and U14879 (N_14879,N_14713,N_14660);
or U14880 (N_14880,N_14698,N_14708);
or U14881 (N_14881,N_14675,N_14679);
and U14882 (N_14882,N_14694,N_14737);
xnor U14883 (N_14883,N_14705,N_14600);
and U14884 (N_14884,N_14754,N_14605);
nor U14885 (N_14885,N_14777,N_14688);
xor U14886 (N_14886,N_14615,N_14767);
nor U14887 (N_14887,N_14654,N_14798);
xor U14888 (N_14888,N_14628,N_14739);
or U14889 (N_14889,N_14652,N_14706);
xnor U14890 (N_14890,N_14638,N_14716);
and U14891 (N_14891,N_14711,N_14771);
nand U14892 (N_14892,N_14761,N_14691);
and U14893 (N_14893,N_14670,N_14724);
nor U14894 (N_14894,N_14636,N_14699);
and U14895 (N_14895,N_14613,N_14631);
nand U14896 (N_14896,N_14651,N_14621);
nand U14897 (N_14897,N_14779,N_14625);
nor U14898 (N_14898,N_14744,N_14707);
xnor U14899 (N_14899,N_14634,N_14616);
xor U14900 (N_14900,N_14604,N_14607);
or U14901 (N_14901,N_14613,N_14645);
nand U14902 (N_14902,N_14697,N_14782);
or U14903 (N_14903,N_14748,N_14765);
nand U14904 (N_14904,N_14614,N_14657);
and U14905 (N_14905,N_14733,N_14741);
nand U14906 (N_14906,N_14625,N_14741);
nor U14907 (N_14907,N_14779,N_14649);
xnor U14908 (N_14908,N_14780,N_14638);
xnor U14909 (N_14909,N_14650,N_14662);
and U14910 (N_14910,N_14708,N_14658);
or U14911 (N_14911,N_14791,N_14685);
xor U14912 (N_14912,N_14775,N_14644);
nand U14913 (N_14913,N_14792,N_14622);
nand U14914 (N_14914,N_14787,N_14760);
or U14915 (N_14915,N_14707,N_14738);
nand U14916 (N_14916,N_14650,N_14655);
xor U14917 (N_14917,N_14773,N_14713);
or U14918 (N_14918,N_14690,N_14738);
nor U14919 (N_14919,N_14693,N_14626);
nand U14920 (N_14920,N_14789,N_14675);
and U14921 (N_14921,N_14643,N_14705);
xor U14922 (N_14922,N_14729,N_14784);
and U14923 (N_14923,N_14648,N_14701);
nand U14924 (N_14924,N_14721,N_14717);
xnor U14925 (N_14925,N_14730,N_14731);
nand U14926 (N_14926,N_14654,N_14650);
nor U14927 (N_14927,N_14604,N_14717);
and U14928 (N_14928,N_14710,N_14614);
nor U14929 (N_14929,N_14601,N_14709);
and U14930 (N_14930,N_14725,N_14632);
nand U14931 (N_14931,N_14691,N_14645);
nor U14932 (N_14932,N_14690,N_14767);
and U14933 (N_14933,N_14730,N_14793);
and U14934 (N_14934,N_14721,N_14728);
xnor U14935 (N_14935,N_14760,N_14628);
nand U14936 (N_14936,N_14618,N_14711);
nor U14937 (N_14937,N_14705,N_14641);
nor U14938 (N_14938,N_14713,N_14671);
and U14939 (N_14939,N_14715,N_14718);
nand U14940 (N_14940,N_14789,N_14647);
xnor U14941 (N_14941,N_14623,N_14733);
nor U14942 (N_14942,N_14692,N_14648);
nor U14943 (N_14943,N_14615,N_14731);
nor U14944 (N_14944,N_14723,N_14620);
or U14945 (N_14945,N_14671,N_14736);
nor U14946 (N_14946,N_14771,N_14794);
or U14947 (N_14947,N_14689,N_14635);
or U14948 (N_14948,N_14776,N_14711);
and U14949 (N_14949,N_14698,N_14605);
nand U14950 (N_14950,N_14739,N_14720);
or U14951 (N_14951,N_14609,N_14772);
xor U14952 (N_14952,N_14721,N_14763);
and U14953 (N_14953,N_14756,N_14626);
nor U14954 (N_14954,N_14685,N_14617);
and U14955 (N_14955,N_14705,N_14635);
nand U14956 (N_14956,N_14646,N_14611);
nand U14957 (N_14957,N_14799,N_14729);
and U14958 (N_14958,N_14725,N_14724);
or U14959 (N_14959,N_14776,N_14742);
or U14960 (N_14960,N_14631,N_14728);
and U14961 (N_14961,N_14793,N_14726);
xor U14962 (N_14962,N_14695,N_14684);
nand U14963 (N_14963,N_14749,N_14786);
nor U14964 (N_14964,N_14681,N_14654);
xnor U14965 (N_14965,N_14750,N_14721);
nand U14966 (N_14966,N_14742,N_14768);
xnor U14967 (N_14967,N_14643,N_14619);
or U14968 (N_14968,N_14656,N_14648);
nor U14969 (N_14969,N_14661,N_14743);
nand U14970 (N_14970,N_14714,N_14789);
nand U14971 (N_14971,N_14791,N_14629);
or U14972 (N_14972,N_14742,N_14687);
xnor U14973 (N_14973,N_14617,N_14633);
nand U14974 (N_14974,N_14762,N_14768);
and U14975 (N_14975,N_14760,N_14653);
or U14976 (N_14976,N_14623,N_14700);
and U14977 (N_14977,N_14759,N_14671);
xor U14978 (N_14978,N_14749,N_14752);
nor U14979 (N_14979,N_14720,N_14740);
and U14980 (N_14980,N_14707,N_14781);
or U14981 (N_14981,N_14786,N_14633);
nand U14982 (N_14982,N_14620,N_14680);
nor U14983 (N_14983,N_14797,N_14779);
xnor U14984 (N_14984,N_14666,N_14772);
nand U14985 (N_14985,N_14731,N_14769);
nand U14986 (N_14986,N_14791,N_14658);
nand U14987 (N_14987,N_14668,N_14711);
xor U14988 (N_14988,N_14722,N_14629);
and U14989 (N_14989,N_14692,N_14717);
nor U14990 (N_14990,N_14799,N_14618);
xnor U14991 (N_14991,N_14785,N_14746);
xnor U14992 (N_14992,N_14719,N_14776);
or U14993 (N_14993,N_14605,N_14635);
xnor U14994 (N_14994,N_14604,N_14661);
xnor U14995 (N_14995,N_14668,N_14684);
or U14996 (N_14996,N_14630,N_14665);
xnor U14997 (N_14997,N_14797,N_14753);
nor U14998 (N_14998,N_14615,N_14792);
nand U14999 (N_14999,N_14646,N_14796);
nand UO_0 (O_0,N_14912,N_14956);
xnor UO_1 (O_1,N_14907,N_14829);
or UO_2 (O_2,N_14849,N_14945);
or UO_3 (O_3,N_14939,N_14835);
or UO_4 (O_4,N_14925,N_14982);
or UO_5 (O_5,N_14926,N_14974);
nor UO_6 (O_6,N_14809,N_14957);
and UO_7 (O_7,N_14811,N_14988);
and UO_8 (O_8,N_14978,N_14864);
nor UO_9 (O_9,N_14966,N_14892);
or UO_10 (O_10,N_14885,N_14842);
xnor UO_11 (O_11,N_14962,N_14946);
xor UO_12 (O_12,N_14879,N_14810);
nor UO_13 (O_13,N_14807,N_14936);
nor UO_14 (O_14,N_14824,N_14823);
nand UO_15 (O_15,N_14803,N_14806);
and UO_16 (O_16,N_14884,N_14913);
and UO_17 (O_17,N_14890,N_14911);
or UO_18 (O_18,N_14960,N_14963);
xor UO_19 (O_19,N_14918,N_14856);
xnor UO_20 (O_20,N_14910,N_14919);
xnor UO_21 (O_21,N_14924,N_14941);
nand UO_22 (O_22,N_14889,N_14942);
nor UO_23 (O_23,N_14985,N_14954);
xor UO_24 (O_24,N_14970,N_14853);
and UO_25 (O_25,N_14801,N_14971);
xnor UO_26 (O_26,N_14851,N_14979);
or UO_27 (O_27,N_14896,N_14815);
or UO_28 (O_28,N_14950,N_14872);
or UO_29 (O_29,N_14871,N_14914);
or UO_30 (O_30,N_14986,N_14969);
xor UO_31 (O_31,N_14862,N_14828);
and UO_32 (O_32,N_14836,N_14876);
or UO_33 (O_33,N_14857,N_14987);
and UO_34 (O_34,N_14874,N_14947);
xor UO_35 (O_35,N_14991,N_14998);
and UO_36 (O_36,N_14819,N_14989);
nor UO_37 (O_37,N_14917,N_14920);
nor UO_38 (O_38,N_14997,N_14983);
nand UO_39 (O_39,N_14882,N_14973);
nor UO_40 (O_40,N_14990,N_14940);
and UO_41 (O_41,N_14886,N_14865);
xor UO_42 (O_42,N_14976,N_14869);
and UO_43 (O_43,N_14933,N_14881);
and UO_44 (O_44,N_14938,N_14800);
xor UO_45 (O_45,N_14814,N_14887);
nand UO_46 (O_46,N_14904,N_14897);
nand UO_47 (O_47,N_14841,N_14980);
nor UO_48 (O_48,N_14880,N_14873);
nor UO_49 (O_49,N_14900,N_14854);
nor UO_50 (O_50,N_14839,N_14894);
or UO_51 (O_51,N_14821,N_14802);
xnor UO_52 (O_52,N_14859,N_14858);
nor UO_53 (O_53,N_14967,N_14943);
xnor UO_54 (O_54,N_14843,N_14826);
and UO_55 (O_55,N_14867,N_14944);
nand UO_56 (O_56,N_14827,N_14955);
and UO_57 (O_57,N_14959,N_14834);
or UO_58 (O_58,N_14916,N_14965);
xnor UO_59 (O_59,N_14994,N_14932);
nor UO_60 (O_60,N_14952,N_14903);
xor UO_61 (O_61,N_14915,N_14968);
and UO_62 (O_62,N_14868,N_14975);
nor UO_63 (O_63,N_14937,N_14804);
or UO_64 (O_64,N_14805,N_14905);
nor UO_65 (O_65,N_14992,N_14995);
nor UO_66 (O_66,N_14877,N_14935);
or UO_67 (O_67,N_14848,N_14844);
and UO_68 (O_68,N_14930,N_14931);
nand UO_69 (O_69,N_14972,N_14822);
nand UO_70 (O_70,N_14934,N_14863);
or UO_71 (O_71,N_14812,N_14830);
nand UO_72 (O_72,N_14977,N_14818);
nor UO_73 (O_73,N_14999,N_14850);
xor UO_74 (O_74,N_14961,N_14866);
nor UO_75 (O_75,N_14908,N_14981);
nand UO_76 (O_76,N_14878,N_14846);
and UO_77 (O_77,N_14899,N_14825);
nor UO_78 (O_78,N_14847,N_14883);
nand UO_79 (O_79,N_14901,N_14928);
xor UO_80 (O_80,N_14845,N_14927);
xnor UO_81 (O_81,N_14808,N_14893);
nor UO_82 (O_82,N_14929,N_14813);
and UO_83 (O_83,N_14816,N_14832);
xnor UO_84 (O_84,N_14993,N_14852);
xnor UO_85 (O_85,N_14948,N_14984);
or UO_86 (O_86,N_14958,N_14895);
and UO_87 (O_87,N_14838,N_14902);
nor UO_88 (O_88,N_14875,N_14888);
or UO_89 (O_89,N_14831,N_14840);
xor UO_90 (O_90,N_14861,N_14922);
xnor UO_91 (O_91,N_14833,N_14949);
xor UO_92 (O_92,N_14837,N_14964);
and UO_93 (O_93,N_14870,N_14906);
nand UO_94 (O_94,N_14996,N_14953);
nand UO_95 (O_95,N_14817,N_14951);
or UO_96 (O_96,N_14898,N_14909);
nand UO_97 (O_97,N_14921,N_14891);
nand UO_98 (O_98,N_14855,N_14923);
nand UO_99 (O_99,N_14860,N_14820);
and UO_100 (O_100,N_14884,N_14915);
xor UO_101 (O_101,N_14873,N_14940);
nand UO_102 (O_102,N_14909,N_14803);
xor UO_103 (O_103,N_14881,N_14804);
xor UO_104 (O_104,N_14913,N_14954);
and UO_105 (O_105,N_14802,N_14931);
xor UO_106 (O_106,N_14807,N_14804);
nor UO_107 (O_107,N_14847,N_14904);
nand UO_108 (O_108,N_14932,N_14857);
nand UO_109 (O_109,N_14948,N_14906);
nor UO_110 (O_110,N_14822,N_14940);
or UO_111 (O_111,N_14957,N_14923);
or UO_112 (O_112,N_14918,N_14852);
xor UO_113 (O_113,N_14927,N_14855);
nor UO_114 (O_114,N_14911,N_14887);
nor UO_115 (O_115,N_14968,N_14824);
xnor UO_116 (O_116,N_14817,N_14903);
or UO_117 (O_117,N_14869,N_14890);
nor UO_118 (O_118,N_14940,N_14914);
or UO_119 (O_119,N_14848,N_14980);
and UO_120 (O_120,N_14934,N_14968);
or UO_121 (O_121,N_14960,N_14981);
nand UO_122 (O_122,N_14916,N_14803);
xor UO_123 (O_123,N_14921,N_14968);
nor UO_124 (O_124,N_14990,N_14897);
and UO_125 (O_125,N_14855,N_14991);
nand UO_126 (O_126,N_14813,N_14939);
nor UO_127 (O_127,N_14883,N_14856);
xnor UO_128 (O_128,N_14816,N_14839);
or UO_129 (O_129,N_14970,N_14920);
or UO_130 (O_130,N_14923,N_14954);
nand UO_131 (O_131,N_14815,N_14818);
or UO_132 (O_132,N_14938,N_14889);
and UO_133 (O_133,N_14834,N_14907);
or UO_134 (O_134,N_14893,N_14870);
or UO_135 (O_135,N_14940,N_14957);
nand UO_136 (O_136,N_14993,N_14959);
or UO_137 (O_137,N_14933,N_14888);
or UO_138 (O_138,N_14973,N_14933);
nor UO_139 (O_139,N_14991,N_14870);
nand UO_140 (O_140,N_14805,N_14885);
nor UO_141 (O_141,N_14951,N_14876);
nor UO_142 (O_142,N_14822,N_14870);
nand UO_143 (O_143,N_14864,N_14986);
xnor UO_144 (O_144,N_14811,N_14850);
nor UO_145 (O_145,N_14827,N_14880);
xor UO_146 (O_146,N_14874,N_14929);
xnor UO_147 (O_147,N_14821,N_14925);
nor UO_148 (O_148,N_14939,N_14846);
nor UO_149 (O_149,N_14946,N_14992);
or UO_150 (O_150,N_14934,N_14950);
nand UO_151 (O_151,N_14991,N_14916);
nor UO_152 (O_152,N_14866,N_14998);
xor UO_153 (O_153,N_14805,N_14976);
nand UO_154 (O_154,N_14931,N_14976);
or UO_155 (O_155,N_14870,N_14856);
xor UO_156 (O_156,N_14988,N_14832);
xor UO_157 (O_157,N_14985,N_14888);
nor UO_158 (O_158,N_14930,N_14915);
nor UO_159 (O_159,N_14946,N_14856);
nand UO_160 (O_160,N_14873,N_14876);
and UO_161 (O_161,N_14826,N_14952);
xnor UO_162 (O_162,N_14885,N_14971);
nor UO_163 (O_163,N_14813,N_14899);
xor UO_164 (O_164,N_14829,N_14924);
nor UO_165 (O_165,N_14854,N_14828);
and UO_166 (O_166,N_14993,N_14932);
and UO_167 (O_167,N_14868,N_14821);
nor UO_168 (O_168,N_14824,N_14839);
xor UO_169 (O_169,N_14995,N_14927);
or UO_170 (O_170,N_14820,N_14808);
nand UO_171 (O_171,N_14950,N_14864);
and UO_172 (O_172,N_14855,N_14856);
xor UO_173 (O_173,N_14994,N_14984);
and UO_174 (O_174,N_14963,N_14970);
nand UO_175 (O_175,N_14934,N_14975);
nand UO_176 (O_176,N_14855,N_14920);
and UO_177 (O_177,N_14841,N_14964);
nand UO_178 (O_178,N_14972,N_14897);
xor UO_179 (O_179,N_14905,N_14840);
xnor UO_180 (O_180,N_14939,N_14871);
nor UO_181 (O_181,N_14932,N_14957);
nand UO_182 (O_182,N_14937,N_14955);
nand UO_183 (O_183,N_14896,N_14936);
xor UO_184 (O_184,N_14894,N_14888);
nor UO_185 (O_185,N_14953,N_14911);
and UO_186 (O_186,N_14984,N_14954);
xnor UO_187 (O_187,N_14922,N_14949);
xor UO_188 (O_188,N_14931,N_14814);
or UO_189 (O_189,N_14862,N_14800);
nand UO_190 (O_190,N_14827,N_14836);
nand UO_191 (O_191,N_14981,N_14896);
and UO_192 (O_192,N_14840,N_14868);
or UO_193 (O_193,N_14992,N_14903);
nor UO_194 (O_194,N_14839,N_14940);
and UO_195 (O_195,N_14859,N_14946);
nand UO_196 (O_196,N_14936,N_14981);
xnor UO_197 (O_197,N_14910,N_14898);
xor UO_198 (O_198,N_14997,N_14965);
nor UO_199 (O_199,N_14927,N_14935);
nor UO_200 (O_200,N_14916,N_14827);
nor UO_201 (O_201,N_14824,N_14920);
and UO_202 (O_202,N_14969,N_14846);
or UO_203 (O_203,N_14978,N_14899);
nand UO_204 (O_204,N_14925,N_14868);
xnor UO_205 (O_205,N_14856,N_14863);
nor UO_206 (O_206,N_14977,N_14855);
or UO_207 (O_207,N_14930,N_14956);
or UO_208 (O_208,N_14878,N_14999);
nand UO_209 (O_209,N_14811,N_14930);
and UO_210 (O_210,N_14988,N_14931);
and UO_211 (O_211,N_14939,N_14920);
nand UO_212 (O_212,N_14855,N_14859);
nand UO_213 (O_213,N_14979,N_14841);
xor UO_214 (O_214,N_14855,N_14964);
nor UO_215 (O_215,N_14826,N_14815);
nor UO_216 (O_216,N_14990,N_14900);
and UO_217 (O_217,N_14851,N_14930);
xnor UO_218 (O_218,N_14933,N_14907);
and UO_219 (O_219,N_14807,N_14864);
nand UO_220 (O_220,N_14991,N_14948);
xor UO_221 (O_221,N_14878,N_14829);
nand UO_222 (O_222,N_14834,N_14823);
xor UO_223 (O_223,N_14844,N_14893);
and UO_224 (O_224,N_14944,N_14866);
xor UO_225 (O_225,N_14840,N_14811);
nand UO_226 (O_226,N_14991,N_14976);
or UO_227 (O_227,N_14974,N_14838);
and UO_228 (O_228,N_14872,N_14919);
xor UO_229 (O_229,N_14965,N_14883);
or UO_230 (O_230,N_14812,N_14874);
xnor UO_231 (O_231,N_14927,N_14980);
or UO_232 (O_232,N_14842,N_14946);
xor UO_233 (O_233,N_14824,N_14881);
xnor UO_234 (O_234,N_14857,N_14994);
and UO_235 (O_235,N_14911,N_14884);
or UO_236 (O_236,N_14904,N_14983);
or UO_237 (O_237,N_14855,N_14904);
nor UO_238 (O_238,N_14800,N_14904);
or UO_239 (O_239,N_14964,N_14822);
and UO_240 (O_240,N_14879,N_14932);
or UO_241 (O_241,N_14963,N_14834);
and UO_242 (O_242,N_14952,N_14923);
nor UO_243 (O_243,N_14920,N_14887);
and UO_244 (O_244,N_14981,N_14879);
or UO_245 (O_245,N_14943,N_14924);
nor UO_246 (O_246,N_14905,N_14800);
xor UO_247 (O_247,N_14863,N_14993);
nand UO_248 (O_248,N_14886,N_14810);
nor UO_249 (O_249,N_14913,N_14858);
xnor UO_250 (O_250,N_14864,N_14852);
nor UO_251 (O_251,N_14827,N_14984);
xor UO_252 (O_252,N_14965,N_14801);
nand UO_253 (O_253,N_14950,N_14916);
xor UO_254 (O_254,N_14851,N_14952);
nor UO_255 (O_255,N_14953,N_14861);
and UO_256 (O_256,N_14990,N_14925);
nand UO_257 (O_257,N_14975,N_14972);
xor UO_258 (O_258,N_14843,N_14923);
or UO_259 (O_259,N_14826,N_14965);
nor UO_260 (O_260,N_14984,N_14851);
nand UO_261 (O_261,N_14845,N_14926);
nand UO_262 (O_262,N_14852,N_14985);
or UO_263 (O_263,N_14932,N_14846);
and UO_264 (O_264,N_14825,N_14800);
or UO_265 (O_265,N_14942,N_14884);
nor UO_266 (O_266,N_14983,N_14849);
or UO_267 (O_267,N_14910,N_14909);
nor UO_268 (O_268,N_14967,N_14932);
and UO_269 (O_269,N_14950,N_14828);
nand UO_270 (O_270,N_14938,N_14853);
nand UO_271 (O_271,N_14857,N_14908);
nor UO_272 (O_272,N_14836,N_14926);
or UO_273 (O_273,N_14930,N_14926);
or UO_274 (O_274,N_14848,N_14988);
or UO_275 (O_275,N_14983,N_14885);
xor UO_276 (O_276,N_14813,N_14831);
nand UO_277 (O_277,N_14985,N_14863);
nand UO_278 (O_278,N_14823,N_14860);
nor UO_279 (O_279,N_14814,N_14963);
nor UO_280 (O_280,N_14916,N_14866);
xnor UO_281 (O_281,N_14897,N_14886);
or UO_282 (O_282,N_14957,N_14838);
nand UO_283 (O_283,N_14891,N_14924);
xor UO_284 (O_284,N_14880,N_14946);
nand UO_285 (O_285,N_14979,N_14948);
and UO_286 (O_286,N_14869,N_14982);
xnor UO_287 (O_287,N_14999,N_14899);
nand UO_288 (O_288,N_14866,N_14877);
and UO_289 (O_289,N_14875,N_14970);
or UO_290 (O_290,N_14928,N_14990);
and UO_291 (O_291,N_14968,N_14919);
nor UO_292 (O_292,N_14826,N_14927);
nor UO_293 (O_293,N_14915,N_14925);
xnor UO_294 (O_294,N_14801,N_14831);
nand UO_295 (O_295,N_14805,N_14917);
xor UO_296 (O_296,N_14914,N_14811);
xor UO_297 (O_297,N_14961,N_14885);
xnor UO_298 (O_298,N_14820,N_14906);
or UO_299 (O_299,N_14911,N_14974);
nand UO_300 (O_300,N_14911,N_14855);
xor UO_301 (O_301,N_14852,N_14851);
nand UO_302 (O_302,N_14890,N_14898);
nand UO_303 (O_303,N_14912,N_14924);
xor UO_304 (O_304,N_14800,N_14869);
and UO_305 (O_305,N_14997,N_14863);
or UO_306 (O_306,N_14998,N_14995);
or UO_307 (O_307,N_14874,N_14955);
nand UO_308 (O_308,N_14928,N_14912);
and UO_309 (O_309,N_14878,N_14983);
and UO_310 (O_310,N_14881,N_14895);
and UO_311 (O_311,N_14860,N_14967);
nor UO_312 (O_312,N_14803,N_14875);
or UO_313 (O_313,N_14983,N_14952);
and UO_314 (O_314,N_14916,N_14829);
and UO_315 (O_315,N_14981,N_14836);
nand UO_316 (O_316,N_14987,N_14896);
xnor UO_317 (O_317,N_14847,N_14874);
and UO_318 (O_318,N_14929,N_14881);
nor UO_319 (O_319,N_14871,N_14953);
or UO_320 (O_320,N_14868,N_14959);
nor UO_321 (O_321,N_14996,N_14969);
nand UO_322 (O_322,N_14816,N_14866);
and UO_323 (O_323,N_14881,N_14803);
and UO_324 (O_324,N_14907,N_14994);
nor UO_325 (O_325,N_14947,N_14914);
nand UO_326 (O_326,N_14865,N_14802);
or UO_327 (O_327,N_14804,N_14854);
and UO_328 (O_328,N_14803,N_14867);
xor UO_329 (O_329,N_14950,N_14998);
and UO_330 (O_330,N_14843,N_14903);
or UO_331 (O_331,N_14912,N_14856);
nand UO_332 (O_332,N_14816,N_14954);
xor UO_333 (O_333,N_14919,N_14908);
or UO_334 (O_334,N_14847,N_14894);
or UO_335 (O_335,N_14862,N_14963);
nand UO_336 (O_336,N_14851,N_14848);
xnor UO_337 (O_337,N_14862,N_14923);
nand UO_338 (O_338,N_14863,N_14922);
and UO_339 (O_339,N_14869,N_14847);
nor UO_340 (O_340,N_14811,N_14837);
nand UO_341 (O_341,N_14932,N_14803);
and UO_342 (O_342,N_14856,N_14859);
xor UO_343 (O_343,N_14915,N_14802);
nand UO_344 (O_344,N_14899,N_14800);
and UO_345 (O_345,N_14949,N_14947);
and UO_346 (O_346,N_14843,N_14851);
nand UO_347 (O_347,N_14894,N_14867);
nor UO_348 (O_348,N_14963,N_14897);
nor UO_349 (O_349,N_14845,N_14897);
and UO_350 (O_350,N_14878,N_14955);
nor UO_351 (O_351,N_14910,N_14953);
and UO_352 (O_352,N_14806,N_14950);
and UO_353 (O_353,N_14996,N_14988);
nor UO_354 (O_354,N_14900,N_14995);
and UO_355 (O_355,N_14928,N_14815);
and UO_356 (O_356,N_14961,N_14849);
xor UO_357 (O_357,N_14905,N_14932);
and UO_358 (O_358,N_14826,N_14947);
xor UO_359 (O_359,N_14912,N_14998);
nand UO_360 (O_360,N_14829,N_14988);
and UO_361 (O_361,N_14890,N_14919);
and UO_362 (O_362,N_14803,N_14868);
and UO_363 (O_363,N_14808,N_14910);
xnor UO_364 (O_364,N_14963,N_14859);
nand UO_365 (O_365,N_14972,N_14824);
nand UO_366 (O_366,N_14831,N_14907);
nand UO_367 (O_367,N_14917,N_14817);
and UO_368 (O_368,N_14976,N_14814);
xor UO_369 (O_369,N_14870,N_14802);
or UO_370 (O_370,N_14933,N_14963);
nor UO_371 (O_371,N_14807,N_14965);
or UO_372 (O_372,N_14915,N_14936);
or UO_373 (O_373,N_14809,N_14916);
or UO_374 (O_374,N_14910,N_14935);
xnor UO_375 (O_375,N_14824,N_14802);
xor UO_376 (O_376,N_14818,N_14854);
or UO_377 (O_377,N_14955,N_14972);
nor UO_378 (O_378,N_14861,N_14878);
nand UO_379 (O_379,N_14855,N_14921);
nor UO_380 (O_380,N_14961,N_14897);
and UO_381 (O_381,N_14835,N_14808);
nand UO_382 (O_382,N_14965,N_14836);
nor UO_383 (O_383,N_14875,N_14879);
xnor UO_384 (O_384,N_14908,N_14872);
nor UO_385 (O_385,N_14921,N_14947);
xnor UO_386 (O_386,N_14907,N_14899);
or UO_387 (O_387,N_14860,N_14812);
nand UO_388 (O_388,N_14859,N_14825);
and UO_389 (O_389,N_14982,N_14886);
xor UO_390 (O_390,N_14903,N_14809);
nand UO_391 (O_391,N_14990,N_14891);
xnor UO_392 (O_392,N_14824,N_14898);
nor UO_393 (O_393,N_14874,N_14914);
xor UO_394 (O_394,N_14962,N_14862);
nor UO_395 (O_395,N_14960,N_14839);
xnor UO_396 (O_396,N_14866,N_14810);
and UO_397 (O_397,N_14893,N_14852);
or UO_398 (O_398,N_14981,N_14811);
or UO_399 (O_399,N_14939,N_14836);
or UO_400 (O_400,N_14871,N_14894);
nand UO_401 (O_401,N_14800,N_14927);
xnor UO_402 (O_402,N_14915,N_14914);
nor UO_403 (O_403,N_14958,N_14862);
and UO_404 (O_404,N_14812,N_14904);
and UO_405 (O_405,N_14941,N_14892);
or UO_406 (O_406,N_14922,N_14830);
and UO_407 (O_407,N_14924,N_14975);
nor UO_408 (O_408,N_14861,N_14841);
nand UO_409 (O_409,N_14930,N_14808);
xnor UO_410 (O_410,N_14951,N_14880);
or UO_411 (O_411,N_14825,N_14836);
and UO_412 (O_412,N_14896,N_14837);
or UO_413 (O_413,N_14975,N_14907);
xnor UO_414 (O_414,N_14826,N_14849);
or UO_415 (O_415,N_14931,N_14821);
or UO_416 (O_416,N_14852,N_14868);
xnor UO_417 (O_417,N_14809,N_14973);
and UO_418 (O_418,N_14954,N_14807);
and UO_419 (O_419,N_14903,N_14882);
nand UO_420 (O_420,N_14979,N_14916);
nand UO_421 (O_421,N_14931,N_14932);
nor UO_422 (O_422,N_14832,N_14922);
and UO_423 (O_423,N_14815,N_14841);
or UO_424 (O_424,N_14806,N_14920);
xnor UO_425 (O_425,N_14944,N_14884);
xor UO_426 (O_426,N_14871,N_14838);
nor UO_427 (O_427,N_14878,N_14812);
or UO_428 (O_428,N_14936,N_14931);
and UO_429 (O_429,N_14995,N_14830);
xnor UO_430 (O_430,N_14840,N_14994);
nand UO_431 (O_431,N_14854,N_14860);
xnor UO_432 (O_432,N_14800,N_14889);
and UO_433 (O_433,N_14861,N_14842);
nand UO_434 (O_434,N_14982,N_14951);
nor UO_435 (O_435,N_14813,N_14912);
and UO_436 (O_436,N_14805,N_14897);
and UO_437 (O_437,N_14930,N_14981);
xnor UO_438 (O_438,N_14800,N_14857);
nor UO_439 (O_439,N_14873,N_14858);
or UO_440 (O_440,N_14945,N_14984);
and UO_441 (O_441,N_14876,N_14831);
nor UO_442 (O_442,N_14875,N_14918);
nand UO_443 (O_443,N_14917,N_14869);
nand UO_444 (O_444,N_14968,N_14825);
nand UO_445 (O_445,N_14891,N_14859);
xnor UO_446 (O_446,N_14808,N_14841);
nand UO_447 (O_447,N_14876,N_14819);
xnor UO_448 (O_448,N_14949,N_14958);
xnor UO_449 (O_449,N_14969,N_14950);
xor UO_450 (O_450,N_14996,N_14805);
nand UO_451 (O_451,N_14958,N_14850);
xnor UO_452 (O_452,N_14863,N_14999);
nand UO_453 (O_453,N_14888,N_14870);
or UO_454 (O_454,N_14948,N_14858);
and UO_455 (O_455,N_14856,N_14887);
and UO_456 (O_456,N_14977,N_14829);
and UO_457 (O_457,N_14931,N_14949);
nand UO_458 (O_458,N_14932,N_14917);
nor UO_459 (O_459,N_14904,N_14861);
nor UO_460 (O_460,N_14880,N_14958);
or UO_461 (O_461,N_14905,N_14897);
nor UO_462 (O_462,N_14985,N_14978);
nand UO_463 (O_463,N_14847,N_14915);
and UO_464 (O_464,N_14997,N_14830);
nand UO_465 (O_465,N_14832,N_14920);
nor UO_466 (O_466,N_14996,N_14951);
xnor UO_467 (O_467,N_14833,N_14837);
and UO_468 (O_468,N_14887,N_14843);
and UO_469 (O_469,N_14946,N_14989);
or UO_470 (O_470,N_14906,N_14953);
nand UO_471 (O_471,N_14870,N_14942);
or UO_472 (O_472,N_14927,N_14824);
nor UO_473 (O_473,N_14975,N_14908);
nand UO_474 (O_474,N_14816,N_14930);
xor UO_475 (O_475,N_14826,N_14879);
nor UO_476 (O_476,N_14828,N_14809);
nand UO_477 (O_477,N_14858,N_14987);
or UO_478 (O_478,N_14818,N_14823);
or UO_479 (O_479,N_14818,N_14968);
nor UO_480 (O_480,N_14909,N_14806);
nor UO_481 (O_481,N_14910,N_14897);
and UO_482 (O_482,N_14892,N_14866);
and UO_483 (O_483,N_14964,N_14895);
and UO_484 (O_484,N_14959,N_14986);
or UO_485 (O_485,N_14893,N_14814);
and UO_486 (O_486,N_14961,N_14901);
xnor UO_487 (O_487,N_14934,N_14839);
nor UO_488 (O_488,N_14862,N_14830);
or UO_489 (O_489,N_14863,N_14870);
and UO_490 (O_490,N_14818,N_14893);
or UO_491 (O_491,N_14937,N_14968);
and UO_492 (O_492,N_14805,N_14863);
nand UO_493 (O_493,N_14866,N_14964);
nand UO_494 (O_494,N_14953,N_14975);
xnor UO_495 (O_495,N_14969,N_14910);
nor UO_496 (O_496,N_14940,N_14851);
or UO_497 (O_497,N_14851,N_14844);
and UO_498 (O_498,N_14980,N_14820);
or UO_499 (O_499,N_14819,N_14908);
nand UO_500 (O_500,N_14959,N_14825);
nand UO_501 (O_501,N_14968,N_14895);
and UO_502 (O_502,N_14991,N_14949);
and UO_503 (O_503,N_14993,N_14971);
nand UO_504 (O_504,N_14889,N_14826);
or UO_505 (O_505,N_14908,N_14896);
xor UO_506 (O_506,N_14983,N_14853);
or UO_507 (O_507,N_14810,N_14850);
and UO_508 (O_508,N_14857,N_14807);
xor UO_509 (O_509,N_14986,N_14927);
nor UO_510 (O_510,N_14991,N_14987);
nand UO_511 (O_511,N_14943,N_14802);
xnor UO_512 (O_512,N_14814,N_14884);
xnor UO_513 (O_513,N_14907,N_14852);
xor UO_514 (O_514,N_14971,N_14986);
nor UO_515 (O_515,N_14842,N_14811);
and UO_516 (O_516,N_14842,N_14894);
and UO_517 (O_517,N_14843,N_14928);
nor UO_518 (O_518,N_14802,N_14830);
xnor UO_519 (O_519,N_14801,N_14803);
xnor UO_520 (O_520,N_14804,N_14801);
and UO_521 (O_521,N_14843,N_14875);
nand UO_522 (O_522,N_14991,N_14964);
and UO_523 (O_523,N_14864,N_14901);
nand UO_524 (O_524,N_14864,N_14889);
nor UO_525 (O_525,N_14948,N_14871);
nand UO_526 (O_526,N_14817,N_14923);
nor UO_527 (O_527,N_14908,N_14932);
nor UO_528 (O_528,N_14969,N_14829);
nor UO_529 (O_529,N_14887,N_14840);
nand UO_530 (O_530,N_14867,N_14883);
nor UO_531 (O_531,N_14867,N_14855);
nor UO_532 (O_532,N_14803,N_14887);
nand UO_533 (O_533,N_14950,N_14845);
nand UO_534 (O_534,N_14992,N_14940);
or UO_535 (O_535,N_14845,N_14979);
nor UO_536 (O_536,N_14840,N_14934);
nand UO_537 (O_537,N_14874,N_14982);
xnor UO_538 (O_538,N_14954,N_14870);
and UO_539 (O_539,N_14825,N_14889);
or UO_540 (O_540,N_14807,N_14944);
and UO_541 (O_541,N_14840,N_14958);
xor UO_542 (O_542,N_14802,N_14833);
and UO_543 (O_543,N_14925,N_14979);
or UO_544 (O_544,N_14837,N_14963);
or UO_545 (O_545,N_14890,N_14861);
or UO_546 (O_546,N_14879,N_14944);
and UO_547 (O_547,N_14970,N_14898);
xnor UO_548 (O_548,N_14933,N_14827);
xnor UO_549 (O_549,N_14832,N_14885);
xor UO_550 (O_550,N_14944,N_14993);
or UO_551 (O_551,N_14943,N_14852);
nor UO_552 (O_552,N_14963,N_14983);
nand UO_553 (O_553,N_14865,N_14951);
and UO_554 (O_554,N_14800,N_14976);
or UO_555 (O_555,N_14978,N_14838);
nor UO_556 (O_556,N_14816,N_14889);
and UO_557 (O_557,N_14912,N_14991);
nor UO_558 (O_558,N_14994,N_14996);
or UO_559 (O_559,N_14955,N_14970);
or UO_560 (O_560,N_14998,N_14888);
nand UO_561 (O_561,N_14961,N_14983);
xor UO_562 (O_562,N_14826,N_14953);
and UO_563 (O_563,N_14986,N_14868);
nor UO_564 (O_564,N_14891,N_14819);
or UO_565 (O_565,N_14810,N_14877);
nand UO_566 (O_566,N_14969,N_14927);
nand UO_567 (O_567,N_14915,N_14991);
or UO_568 (O_568,N_14885,N_14916);
xor UO_569 (O_569,N_14995,N_14873);
xnor UO_570 (O_570,N_14855,N_14955);
xor UO_571 (O_571,N_14836,N_14948);
xor UO_572 (O_572,N_14926,N_14927);
nor UO_573 (O_573,N_14854,N_14889);
xor UO_574 (O_574,N_14807,N_14925);
and UO_575 (O_575,N_14868,N_14871);
and UO_576 (O_576,N_14932,N_14874);
nand UO_577 (O_577,N_14923,N_14927);
nor UO_578 (O_578,N_14804,N_14964);
xor UO_579 (O_579,N_14995,N_14885);
or UO_580 (O_580,N_14999,N_14845);
nand UO_581 (O_581,N_14964,N_14849);
nor UO_582 (O_582,N_14845,N_14904);
xor UO_583 (O_583,N_14822,N_14853);
or UO_584 (O_584,N_14934,N_14965);
nor UO_585 (O_585,N_14907,N_14910);
and UO_586 (O_586,N_14805,N_14910);
xnor UO_587 (O_587,N_14946,N_14930);
nor UO_588 (O_588,N_14925,N_14977);
nor UO_589 (O_589,N_14981,N_14838);
nor UO_590 (O_590,N_14992,N_14986);
or UO_591 (O_591,N_14806,N_14958);
and UO_592 (O_592,N_14968,N_14809);
nor UO_593 (O_593,N_14996,N_14877);
or UO_594 (O_594,N_14854,N_14998);
nand UO_595 (O_595,N_14964,N_14863);
nor UO_596 (O_596,N_14943,N_14951);
or UO_597 (O_597,N_14939,N_14811);
nor UO_598 (O_598,N_14869,N_14979);
xnor UO_599 (O_599,N_14824,N_14919);
and UO_600 (O_600,N_14815,N_14882);
and UO_601 (O_601,N_14979,N_14853);
xor UO_602 (O_602,N_14844,N_14846);
xnor UO_603 (O_603,N_14922,N_14843);
nand UO_604 (O_604,N_14918,N_14945);
nand UO_605 (O_605,N_14840,N_14842);
and UO_606 (O_606,N_14885,N_14993);
nand UO_607 (O_607,N_14864,N_14811);
or UO_608 (O_608,N_14822,N_14851);
nand UO_609 (O_609,N_14990,N_14829);
nand UO_610 (O_610,N_14829,N_14945);
and UO_611 (O_611,N_14998,N_14830);
nand UO_612 (O_612,N_14809,N_14939);
or UO_613 (O_613,N_14887,N_14907);
nand UO_614 (O_614,N_14945,N_14959);
and UO_615 (O_615,N_14943,N_14826);
xnor UO_616 (O_616,N_14864,N_14963);
nor UO_617 (O_617,N_14947,N_14835);
xnor UO_618 (O_618,N_14957,N_14861);
nor UO_619 (O_619,N_14848,N_14866);
nand UO_620 (O_620,N_14918,N_14890);
nor UO_621 (O_621,N_14852,N_14872);
nand UO_622 (O_622,N_14831,N_14851);
nor UO_623 (O_623,N_14903,N_14893);
and UO_624 (O_624,N_14938,N_14810);
nand UO_625 (O_625,N_14979,N_14999);
or UO_626 (O_626,N_14932,N_14929);
xor UO_627 (O_627,N_14878,N_14817);
xnor UO_628 (O_628,N_14882,N_14874);
or UO_629 (O_629,N_14968,N_14812);
or UO_630 (O_630,N_14896,N_14978);
nand UO_631 (O_631,N_14865,N_14926);
or UO_632 (O_632,N_14934,N_14978);
xnor UO_633 (O_633,N_14895,N_14827);
xnor UO_634 (O_634,N_14867,N_14852);
or UO_635 (O_635,N_14947,N_14969);
or UO_636 (O_636,N_14938,N_14884);
nand UO_637 (O_637,N_14981,N_14946);
nand UO_638 (O_638,N_14932,N_14836);
nor UO_639 (O_639,N_14981,N_14825);
nand UO_640 (O_640,N_14816,N_14873);
xor UO_641 (O_641,N_14944,N_14957);
nand UO_642 (O_642,N_14964,N_14853);
nor UO_643 (O_643,N_14935,N_14923);
or UO_644 (O_644,N_14823,N_14963);
or UO_645 (O_645,N_14913,N_14818);
nor UO_646 (O_646,N_14941,N_14849);
and UO_647 (O_647,N_14850,N_14802);
xor UO_648 (O_648,N_14913,N_14829);
nor UO_649 (O_649,N_14863,N_14835);
xnor UO_650 (O_650,N_14810,N_14991);
and UO_651 (O_651,N_14948,N_14819);
and UO_652 (O_652,N_14966,N_14823);
nor UO_653 (O_653,N_14920,N_14909);
and UO_654 (O_654,N_14969,N_14866);
nor UO_655 (O_655,N_14939,N_14878);
and UO_656 (O_656,N_14950,N_14808);
or UO_657 (O_657,N_14904,N_14877);
xnor UO_658 (O_658,N_14870,N_14980);
xor UO_659 (O_659,N_14841,N_14934);
or UO_660 (O_660,N_14954,N_14915);
and UO_661 (O_661,N_14966,N_14938);
nor UO_662 (O_662,N_14833,N_14914);
xor UO_663 (O_663,N_14977,N_14900);
and UO_664 (O_664,N_14958,N_14838);
or UO_665 (O_665,N_14866,N_14960);
and UO_666 (O_666,N_14819,N_14978);
xnor UO_667 (O_667,N_14803,N_14938);
nand UO_668 (O_668,N_14846,N_14824);
xor UO_669 (O_669,N_14918,N_14921);
and UO_670 (O_670,N_14943,N_14906);
and UO_671 (O_671,N_14915,N_14981);
xor UO_672 (O_672,N_14814,N_14933);
nand UO_673 (O_673,N_14939,N_14938);
xor UO_674 (O_674,N_14915,N_14899);
xor UO_675 (O_675,N_14807,N_14964);
nand UO_676 (O_676,N_14809,N_14982);
nor UO_677 (O_677,N_14893,N_14916);
or UO_678 (O_678,N_14816,N_14886);
or UO_679 (O_679,N_14830,N_14810);
or UO_680 (O_680,N_14985,N_14804);
xor UO_681 (O_681,N_14893,N_14802);
and UO_682 (O_682,N_14802,N_14812);
nand UO_683 (O_683,N_14800,N_14895);
and UO_684 (O_684,N_14893,N_14975);
and UO_685 (O_685,N_14887,N_14857);
and UO_686 (O_686,N_14938,N_14957);
nor UO_687 (O_687,N_14863,N_14897);
xnor UO_688 (O_688,N_14931,N_14812);
nor UO_689 (O_689,N_14992,N_14828);
and UO_690 (O_690,N_14909,N_14936);
nor UO_691 (O_691,N_14830,N_14994);
nand UO_692 (O_692,N_14895,N_14938);
nand UO_693 (O_693,N_14881,N_14852);
nand UO_694 (O_694,N_14891,N_14906);
and UO_695 (O_695,N_14841,N_14820);
or UO_696 (O_696,N_14910,N_14833);
nand UO_697 (O_697,N_14970,N_14828);
nor UO_698 (O_698,N_14948,N_14999);
nand UO_699 (O_699,N_14877,N_14970);
nor UO_700 (O_700,N_14896,N_14885);
xor UO_701 (O_701,N_14920,N_14944);
and UO_702 (O_702,N_14970,N_14864);
nor UO_703 (O_703,N_14960,N_14855);
nor UO_704 (O_704,N_14919,N_14813);
nand UO_705 (O_705,N_14841,N_14898);
xor UO_706 (O_706,N_14894,N_14946);
nand UO_707 (O_707,N_14833,N_14819);
xnor UO_708 (O_708,N_14962,N_14859);
nor UO_709 (O_709,N_14819,N_14953);
xor UO_710 (O_710,N_14993,N_14843);
nand UO_711 (O_711,N_14896,N_14934);
xor UO_712 (O_712,N_14963,N_14879);
nor UO_713 (O_713,N_14981,N_14874);
xor UO_714 (O_714,N_14997,N_14891);
nand UO_715 (O_715,N_14806,N_14917);
or UO_716 (O_716,N_14952,N_14854);
and UO_717 (O_717,N_14846,N_14809);
xor UO_718 (O_718,N_14819,N_14866);
and UO_719 (O_719,N_14913,N_14936);
and UO_720 (O_720,N_14906,N_14864);
or UO_721 (O_721,N_14926,N_14966);
nand UO_722 (O_722,N_14954,N_14987);
and UO_723 (O_723,N_14882,N_14998);
or UO_724 (O_724,N_14803,N_14985);
nand UO_725 (O_725,N_14874,N_14863);
and UO_726 (O_726,N_14899,N_14830);
and UO_727 (O_727,N_14851,N_14893);
and UO_728 (O_728,N_14903,N_14838);
or UO_729 (O_729,N_14896,N_14845);
xor UO_730 (O_730,N_14956,N_14870);
or UO_731 (O_731,N_14895,N_14901);
xor UO_732 (O_732,N_14846,N_14811);
or UO_733 (O_733,N_14923,N_14823);
nor UO_734 (O_734,N_14851,N_14939);
xor UO_735 (O_735,N_14898,N_14969);
nand UO_736 (O_736,N_14864,N_14808);
and UO_737 (O_737,N_14832,N_14882);
or UO_738 (O_738,N_14805,N_14836);
xnor UO_739 (O_739,N_14953,N_14851);
nor UO_740 (O_740,N_14886,N_14947);
and UO_741 (O_741,N_14900,N_14817);
or UO_742 (O_742,N_14886,N_14986);
nor UO_743 (O_743,N_14966,N_14999);
nand UO_744 (O_744,N_14942,N_14871);
nand UO_745 (O_745,N_14863,N_14831);
nand UO_746 (O_746,N_14944,N_14990);
or UO_747 (O_747,N_14916,N_14836);
or UO_748 (O_748,N_14811,N_14803);
nand UO_749 (O_749,N_14921,N_14911);
xnor UO_750 (O_750,N_14801,N_14937);
or UO_751 (O_751,N_14851,N_14891);
or UO_752 (O_752,N_14842,N_14957);
nor UO_753 (O_753,N_14989,N_14853);
or UO_754 (O_754,N_14844,N_14956);
nor UO_755 (O_755,N_14983,N_14805);
or UO_756 (O_756,N_14911,N_14815);
nor UO_757 (O_757,N_14914,N_14985);
or UO_758 (O_758,N_14953,N_14864);
nor UO_759 (O_759,N_14910,N_14817);
or UO_760 (O_760,N_14854,N_14905);
or UO_761 (O_761,N_14914,N_14827);
xor UO_762 (O_762,N_14923,N_14933);
and UO_763 (O_763,N_14847,N_14938);
xnor UO_764 (O_764,N_14937,N_14952);
and UO_765 (O_765,N_14864,N_14914);
and UO_766 (O_766,N_14852,N_14947);
or UO_767 (O_767,N_14969,N_14990);
nand UO_768 (O_768,N_14915,N_14943);
or UO_769 (O_769,N_14944,N_14883);
nor UO_770 (O_770,N_14995,N_14820);
nor UO_771 (O_771,N_14830,N_14879);
xnor UO_772 (O_772,N_14873,N_14802);
xor UO_773 (O_773,N_14834,N_14980);
and UO_774 (O_774,N_14945,N_14814);
nor UO_775 (O_775,N_14971,N_14869);
and UO_776 (O_776,N_14812,N_14810);
and UO_777 (O_777,N_14986,N_14950);
nor UO_778 (O_778,N_14837,N_14957);
nor UO_779 (O_779,N_14934,N_14851);
and UO_780 (O_780,N_14812,N_14843);
and UO_781 (O_781,N_14896,N_14953);
nor UO_782 (O_782,N_14915,N_14928);
nand UO_783 (O_783,N_14944,N_14862);
and UO_784 (O_784,N_14988,N_14942);
xnor UO_785 (O_785,N_14942,N_14921);
nor UO_786 (O_786,N_14816,N_14994);
xnor UO_787 (O_787,N_14947,N_14907);
and UO_788 (O_788,N_14918,N_14822);
xnor UO_789 (O_789,N_14822,N_14933);
xnor UO_790 (O_790,N_14992,N_14989);
xor UO_791 (O_791,N_14855,N_14954);
xor UO_792 (O_792,N_14897,N_14992);
or UO_793 (O_793,N_14996,N_14853);
nand UO_794 (O_794,N_14903,N_14801);
nor UO_795 (O_795,N_14963,N_14905);
xnor UO_796 (O_796,N_14988,N_14995);
xor UO_797 (O_797,N_14975,N_14838);
nand UO_798 (O_798,N_14834,N_14865);
and UO_799 (O_799,N_14923,N_14988);
xnor UO_800 (O_800,N_14830,N_14883);
nand UO_801 (O_801,N_14963,N_14811);
xor UO_802 (O_802,N_14890,N_14936);
or UO_803 (O_803,N_14864,N_14858);
nand UO_804 (O_804,N_14976,N_14817);
nor UO_805 (O_805,N_14844,N_14842);
xnor UO_806 (O_806,N_14837,N_14919);
and UO_807 (O_807,N_14956,N_14935);
or UO_808 (O_808,N_14880,N_14832);
nor UO_809 (O_809,N_14987,N_14910);
nor UO_810 (O_810,N_14871,N_14930);
nand UO_811 (O_811,N_14834,N_14827);
xnor UO_812 (O_812,N_14936,N_14929);
nor UO_813 (O_813,N_14874,N_14975);
nor UO_814 (O_814,N_14867,N_14859);
xnor UO_815 (O_815,N_14910,N_14900);
nor UO_816 (O_816,N_14803,N_14805);
nor UO_817 (O_817,N_14866,N_14972);
nand UO_818 (O_818,N_14948,N_14968);
or UO_819 (O_819,N_14843,N_14958);
nor UO_820 (O_820,N_14971,N_14979);
nand UO_821 (O_821,N_14939,N_14890);
or UO_822 (O_822,N_14894,N_14809);
nor UO_823 (O_823,N_14976,N_14881);
and UO_824 (O_824,N_14998,N_14824);
xnor UO_825 (O_825,N_14930,N_14960);
xnor UO_826 (O_826,N_14948,N_14922);
nand UO_827 (O_827,N_14948,N_14891);
nand UO_828 (O_828,N_14925,N_14999);
nand UO_829 (O_829,N_14812,N_14815);
and UO_830 (O_830,N_14815,N_14904);
nand UO_831 (O_831,N_14927,N_14827);
xor UO_832 (O_832,N_14953,N_14867);
nand UO_833 (O_833,N_14880,N_14808);
xor UO_834 (O_834,N_14805,N_14953);
nor UO_835 (O_835,N_14883,N_14815);
nand UO_836 (O_836,N_14961,N_14988);
nand UO_837 (O_837,N_14830,N_14837);
nand UO_838 (O_838,N_14920,N_14943);
nor UO_839 (O_839,N_14972,N_14950);
or UO_840 (O_840,N_14981,N_14970);
nand UO_841 (O_841,N_14831,N_14886);
xor UO_842 (O_842,N_14815,N_14816);
nor UO_843 (O_843,N_14868,N_14854);
and UO_844 (O_844,N_14871,N_14996);
and UO_845 (O_845,N_14829,N_14917);
xor UO_846 (O_846,N_14893,N_14986);
xnor UO_847 (O_847,N_14830,N_14882);
nor UO_848 (O_848,N_14884,N_14833);
and UO_849 (O_849,N_14915,N_14841);
nor UO_850 (O_850,N_14802,N_14974);
nor UO_851 (O_851,N_14859,N_14890);
xnor UO_852 (O_852,N_14938,N_14915);
and UO_853 (O_853,N_14858,N_14956);
nor UO_854 (O_854,N_14857,N_14924);
xor UO_855 (O_855,N_14913,N_14887);
and UO_856 (O_856,N_14847,N_14996);
xor UO_857 (O_857,N_14937,N_14803);
xor UO_858 (O_858,N_14986,N_14908);
nor UO_859 (O_859,N_14825,N_14862);
or UO_860 (O_860,N_14872,N_14938);
and UO_861 (O_861,N_14863,N_14992);
nor UO_862 (O_862,N_14862,N_14959);
xnor UO_863 (O_863,N_14911,N_14897);
nand UO_864 (O_864,N_14884,N_14926);
or UO_865 (O_865,N_14900,N_14885);
xor UO_866 (O_866,N_14875,N_14907);
and UO_867 (O_867,N_14907,N_14968);
and UO_868 (O_868,N_14889,N_14892);
or UO_869 (O_869,N_14870,N_14834);
xor UO_870 (O_870,N_14882,N_14966);
or UO_871 (O_871,N_14893,N_14835);
nand UO_872 (O_872,N_14812,N_14926);
and UO_873 (O_873,N_14946,N_14920);
nor UO_874 (O_874,N_14862,N_14890);
or UO_875 (O_875,N_14896,N_14963);
nor UO_876 (O_876,N_14977,N_14918);
nand UO_877 (O_877,N_14839,N_14828);
or UO_878 (O_878,N_14887,N_14926);
nand UO_879 (O_879,N_14992,N_14883);
xnor UO_880 (O_880,N_14967,N_14908);
nor UO_881 (O_881,N_14841,N_14876);
nand UO_882 (O_882,N_14901,N_14835);
or UO_883 (O_883,N_14959,N_14965);
nor UO_884 (O_884,N_14996,N_14835);
nand UO_885 (O_885,N_14819,N_14824);
nand UO_886 (O_886,N_14802,N_14867);
and UO_887 (O_887,N_14940,N_14924);
nor UO_888 (O_888,N_14931,N_14803);
and UO_889 (O_889,N_14967,N_14821);
and UO_890 (O_890,N_14865,N_14999);
nor UO_891 (O_891,N_14901,N_14886);
xor UO_892 (O_892,N_14948,N_14855);
and UO_893 (O_893,N_14963,N_14914);
or UO_894 (O_894,N_14908,N_14904);
nand UO_895 (O_895,N_14953,N_14966);
nor UO_896 (O_896,N_14800,N_14890);
nand UO_897 (O_897,N_14887,N_14930);
nand UO_898 (O_898,N_14869,N_14868);
nor UO_899 (O_899,N_14943,N_14999);
or UO_900 (O_900,N_14992,N_14895);
or UO_901 (O_901,N_14929,N_14840);
and UO_902 (O_902,N_14859,N_14967);
and UO_903 (O_903,N_14805,N_14874);
and UO_904 (O_904,N_14939,N_14966);
xor UO_905 (O_905,N_14914,N_14916);
nand UO_906 (O_906,N_14839,N_14944);
nor UO_907 (O_907,N_14880,N_14955);
nor UO_908 (O_908,N_14990,N_14816);
or UO_909 (O_909,N_14936,N_14851);
or UO_910 (O_910,N_14878,N_14901);
nor UO_911 (O_911,N_14873,N_14870);
xnor UO_912 (O_912,N_14950,N_14895);
and UO_913 (O_913,N_14976,N_14946);
or UO_914 (O_914,N_14944,N_14923);
or UO_915 (O_915,N_14816,N_14884);
nand UO_916 (O_916,N_14809,N_14980);
nand UO_917 (O_917,N_14815,N_14903);
nor UO_918 (O_918,N_14947,N_14911);
nor UO_919 (O_919,N_14856,N_14916);
and UO_920 (O_920,N_14833,N_14872);
or UO_921 (O_921,N_14859,N_14844);
nand UO_922 (O_922,N_14858,N_14904);
and UO_923 (O_923,N_14815,N_14830);
xnor UO_924 (O_924,N_14896,N_14843);
xor UO_925 (O_925,N_14827,N_14896);
nor UO_926 (O_926,N_14899,N_14868);
or UO_927 (O_927,N_14903,N_14820);
xnor UO_928 (O_928,N_14943,N_14978);
xnor UO_929 (O_929,N_14896,N_14983);
or UO_930 (O_930,N_14942,N_14834);
nor UO_931 (O_931,N_14851,N_14840);
nor UO_932 (O_932,N_14935,N_14929);
xor UO_933 (O_933,N_14990,N_14885);
or UO_934 (O_934,N_14821,N_14920);
and UO_935 (O_935,N_14914,N_14852);
and UO_936 (O_936,N_14990,N_14805);
nand UO_937 (O_937,N_14991,N_14844);
nand UO_938 (O_938,N_14801,N_14861);
nor UO_939 (O_939,N_14893,N_14878);
nand UO_940 (O_940,N_14961,N_14895);
nand UO_941 (O_941,N_14916,N_14837);
and UO_942 (O_942,N_14817,N_14909);
and UO_943 (O_943,N_14808,N_14960);
and UO_944 (O_944,N_14881,N_14998);
nor UO_945 (O_945,N_14951,N_14977);
nor UO_946 (O_946,N_14924,N_14889);
nand UO_947 (O_947,N_14958,N_14893);
xnor UO_948 (O_948,N_14828,N_14960);
nor UO_949 (O_949,N_14901,N_14833);
xnor UO_950 (O_950,N_14816,N_14804);
xor UO_951 (O_951,N_14812,N_14863);
nand UO_952 (O_952,N_14879,N_14850);
and UO_953 (O_953,N_14974,N_14821);
or UO_954 (O_954,N_14939,N_14914);
nand UO_955 (O_955,N_14929,N_14971);
nand UO_956 (O_956,N_14930,N_14802);
and UO_957 (O_957,N_14828,N_14898);
and UO_958 (O_958,N_14843,N_14897);
nor UO_959 (O_959,N_14893,N_14827);
and UO_960 (O_960,N_14891,N_14880);
xor UO_961 (O_961,N_14983,N_14930);
or UO_962 (O_962,N_14986,N_14878);
nand UO_963 (O_963,N_14966,N_14958);
and UO_964 (O_964,N_14923,N_14800);
or UO_965 (O_965,N_14803,N_14878);
nor UO_966 (O_966,N_14920,N_14840);
xor UO_967 (O_967,N_14982,N_14912);
nor UO_968 (O_968,N_14940,N_14872);
nor UO_969 (O_969,N_14994,N_14801);
nor UO_970 (O_970,N_14902,N_14831);
nor UO_971 (O_971,N_14968,N_14956);
nor UO_972 (O_972,N_14816,N_14933);
and UO_973 (O_973,N_14994,N_14912);
nor UO_974 (O_974,N_14918,N_14941);
nand UO_975 (O_975,N_14881,N_14839);
nor UO_976 (O_976,N_14879,N_14801);
nand UO_977 (O_977,N_14906,N_14874);
xnor UO_978 (O_978,N_14807,N_14963);
nand UO_979 (O_979,N_14892,N_14971);
and UO_980 (O_980,N_14923,N_14830);
nand UO_981 (O_981,N_14828,N_14833);
nor UO_982 (O_982,N_14925,N_14962);
or UO_983 (O_983,N_14959,N_14988);
xor UO_984 (O_984,N_14897,N_14875);
and UO_985 (O_985,N_14870,N_14989);
nand UO_986 (O_986,N_14837,N_14874);
xnor UO_987 (O_987,N_14960,N_14967);
xnor UO_988 (O_988,N_14971,N_14903);
nand UO_989 (O_989,N_14956,N_14957);
nand UO_990 (O_990,N_14817,N_14880);
xnor UO_991 (O_991,N_14802,N_14899);
nand UO_992 (O_992,N_14820,N_14855);
or UO_993 (O_993,N_14918,N_14813);
nand UO_994 (O_994,N_14951,N_14967);
and UO_995 (O_995,N_14996,N_14925);
nor UO_996 (O_996,N_14838,N_14904);
and UO_997 (O_997,N_14971,N_14972);
nor UO_998 (O_998,N_14979,N_14806);
and UO_999 (O_999,N_14843,N_14955);
nor UO_1000 (O_1000,N_14969,N_14879);
nand UO_1001 (O_1001,N_14976,N_14877);
xnor UO_1002 (O_1002,N_14970,N_14985);
nand UO_1003 (O_1003,N_14876,N_14960);
nand UO_1004 (O_1004,N_14885,N_14940);
or UO_1005 (O_1005,N_14970,N_14939);
xor UO_1006 (O_1006,N_14920,N_14987);
xor UO_1007 (O_1007,N_14880,N_14915);
nor UO_1008 (O_1008,N_14852,N_14806);
nor UO_1009 (O_1009,N_14898,N_14831);
xnor UO_1010 (O_1010,N_14825,N_14931);
xnor UO_1011 (O_1011,N_14988,N_14872);
nor UO_1012 (O_1012,N_14931,N_14923);
and UO_1013 (O_1013,N_14986,N_14932);
and UO_1014 (O_1014,N_14878,N_14907);
xor UO_1015 (O_1015,N_14849,N_14926);
or UO_1016 (O_1016,N_14936,N_14918);
and UO_1017 (O_1017,N_14810,N_14818);
nor UO_1018 (O_1018,N_14985,N_14893);
nand UO_1019 (O_1019,N_14870,N_14882);
nand UO_1020 (O_1020,N_14832,N_14842);
nor UO_1021 (O_1021,N_14813,N_14926);
xnor UO_1022 (O_1022,N_14925,N_14932);
and UO_1023 (O_1023,N_14839,N_14951);
or UO_1024 (O_1024,N_14929,N_14828);
or UO_1025 (O_1025,N_14816,N_14921);
nor UO_1026 (O_1026,N_14889,N_14908);
or UO_1027 (O_1027,N_14944,N_14900);
nand UO_1028 (O_1028,N_14855,N_14853);
nor UO_1029 (O_1029,N_14842,N_14929);
and UO_1030 (O_1030,N_14935,N_14824);
xnor UO_1031 (O_1031,N_14994,N_14893);
nand UO_1032 (O_1032,N_14853,N_14913);
nor UO_1033 (O_1033,N_14926,N_14806);
or UO_1034 (O_1034,N_14972,N_14907);
or UO_1035 (O_1035,N_14947,N_14819);
xnor UO_1036 (O_1036,N_14841,N_14826);
xnor UO_1037 (O_1037,N_14840,N_14988);
and UO_1038 (O_1038,N_14855,N_14850);
nand UO_1039 (O_1039,N_14904,N_14961);
and UO_1040 (O_1040,N_14964,N_14871);
nor UO_1041 (O_1041,N_14843,N_14846);
xnor UO_1042 (O_1042,N_14935,N_14987);
nand UO_1043 (O_1043,N_14928,N_14910);
nand UO_1044 (O_1044,N_14863,N_14872);
or UO_1045 (O_1045,N_14975,N_14835);
and UO_1046 (O_1046,N_14978,N_14833);
nand UO_1047 (O_1047,N_14872,N_14867);
or UO_1048 (O_1048,N_14882,N_14972);
and UO_1049 (O_1049,N_14840,N_14817);
nor UO_1050 (O_1050,N_14974,N_14809);
xnor UO_1051 (O_1051,N_14877,N_14852);
and UO_1052 (O_1052,N_14849,N_14904);
nor UO_1053 (O_1053,N_14867,N_14980);
xnor UO_1054 (O_1054,N_14967,N_14853);
and UO_1055 (O_1055,N_14904,N_14933);
or UO_1056 (O_1056,N_14896,N_14849);
nand UO_1057 (O_1057,N_14902,N_14990);
and UO_1058 (O_1058,N_14947,N_14840);
and UO_1059 (O_1059,N_14860,N_14887);
nor UO_1060 (O_1060,N_14910,N_14911);
nand UO_1061 (O_1061,N_14940,N_14981);
or UO_1062 (O_1062,N_14909,N_14969);
nand UO_1063 (O_1063,N_14870,N_14946);
or UO_1064 (O_1064,N_14954,N_14956);
nand UO_1065 (O_1065,N_14859,N_14815);
nand UO_1066 (O_1066,N_14875,N_14949);
xor UO_1067 (O_1067,N_14836,N_14960);
xor UO_1068 (O_1068,N_14917,N_14989);
or UO_1069 (O_1069,N_14804,N_14837);
nor UO_1070 (O_1070,N_14876,N_14931);
or UO_1071 (O_1071,N_14892,N_14825);
nor UO_1072 (O_1072,N_14916,N_14909);
and UO_1073 (O_1073,N_14810,N_14853);
xor UO_1074 (O_1074,N_14980,N_14940);
or UO_1075 (O_1075,N_14905,N_14868);
xor UO_1076 (O_1076,N_14901,N_14897);
or UO_1077 (O_1077,N_14921,N_14823);
xnor UO_1078 (O_1078,N_14894,N_14910);
nor UO_1079 (O_1079,N_14851,N_14810);
nor UO_1080 (O_1080,N_14906,N_14947);
nand UO_1081 (O_1081,N_14833,N_14846);
nand UO_1082 (O_1082,N_14992,N_14917);
or UO_1083 (O_1083,N_14972,N_14807);
nor UO_1084 (O_1084,N_14962,N_14887);
xor UO_1085 (O_1085,N_14812,N_14994);
nor UO_1086 (O_1086,N_14873,N_14928);
and UO_1087 (O_1087,N_14945,N_14946);
or UO_1088 (O_1088,N_14978,N_14939);
xnor UO_1089 (O_1089,N_14973,N_14902);
xor UO_1090 (O_1090,N_14818,N_14885);
nand UO_1091 (O_1091,N_14949,N_14905);
nor UO_1092 (O_1092,N_14953,N_14845);
xnor UO_1093 (O_1093,N_14917,N_14980);
nor UO_1094 (O_1094,N_14901,N_14825);
nand UO_1095 (O_1095,N_14953,N_14872);
and UO_1096 (O_1096,N_14936,N_14848);
nor UO_1097 (O_1097,N_14918,N_14968);
nand UO_1098 (O_1098,N_14800,N_14845);
xnor UO_1099 (O_1099,N_14834,N_14976);
or UO_1100 (O_1100,N_14956,N_14993);
nand UO_1101 (O_1101,N_14804,N_14978);
nand UO_1102 (O_1102,N_14925,N_14860);
and UO_1103 (O_1103,N_14865,N_14870);
or UO_1104 (O_1104,N_14888,N_14954);
xnor UO_1105 (O_1105,N_14829,N_14892);
nand UO_1106 (O_1106,N_14864,N_14819);
or UO_1107 (O_1107,N_14845,N_14965);
and UO_1108 (O_1108,N_14933,N_14849);
or UO_1109 (O_1109,N_14959,N_14943);
nand UO_1110 (O_1110,N_14977,N_14850);
nor UO_1111 (O_1111,N_14850,N_14894);
nor UO_1112 (O_1112,N_14910,N_14821);
nor UO_1113 (O_1113,N_14889,N_14840);
xor UO_1114 (O_1114,N_14954,N_14828);
nand UO_1115 (O_1115,N_14946,N_14959);
xnor UO_1116 (O_1116,N_14896,N_14840);
and UO_1117 (O_1117,N_14917,N_14839);
xor UO_1118 (O_1118,N_14851,N_14958);
xor UO_1119 (O_1119,N_14926,N_14854);
and UO_1120 (O_1120,N_14981,N_14869);
or UO_1121 (O_1121,N_14835,N_14832);
or UO_1122 (O_1122,N_14903,N_14874);
xor UO_1123 (O_1123,N_14887,N_14829);
or UO_1124 (O_1124,N_14913,N_14912);
or UO_1125 (O_1125,N_14892,N_14833);
or UO_1126 (O_1126,N_14874,N_14891);
or UO_1127 (O_1127,N_14882,N_14976);
and UO_1128 (O_1128,N_14811,N_14955);
and UO_1129 (O_1129,N_14825,N_14967);
xnor UO_1130 (O_1130,N_14804,N_14905);
or UO_1131 (O_1131,N_14889,N_14824);
or UO_1132 (O_1132,N_14889,N_14967);
and UO_1133 (O_1133,N_14825,N_14813);
and UO_1134 (O_1134,N_14961,N_14842);
or UO_1135 (O_1135,N_14834,N_14973);
xnor UO_1136 (O_1136,N_14915,N_14817);
nor UO_1137 (O_1137,N_14902,N_14985);
nand UO_1138 (O_1138,N_14844,N_14986);
nor UO_1139 (O_1139,N_14807,N_14911);
and UO_1140 (O_1140,N_14930,N_14833);
or UO_1141 (O_1141,N_14876,N_14844);
and UO_1142 (O_1142,N_14971,N_14880);
nand UO_1143 (O_1143,N_14838,N_14801);
nor UO_1144 (O_1144,N_14885,N_14941);
and UO_1145 (O_1145,N_14893,N_14874);
nand UO_1146 (O_1146,N_14930,N_14913);
nor UO_1147 (O_1147,N_14895,N_14828);
or UO_1148 (O_1148,N_14926,N_14998);
and UO_1149 (O_1149,N_14857,N_14817);
or UO_1150 (O_1150,N_14966,N_14857);
nor UO_1151 (O_1151,N_14985,N_14885);
and UO_1152 (O_1152,N_14866,N_14864);
or UO_1153 (O_1153,N_14942,N_14925);
nand UO_1154 (O_1154,N_14926,N_14905);
or UO_1155 (O_1155,N_14971,N_14906);
or UO_1156 (O_1156,N_14877,N_14918);
and UO_1157 (O_1157,N_14819,N_14941);
xor UO_1158 (O_1158,N_14823,N_14884);
nor UO_1159 (O_1159,N_14904,N_14979);
nor UO_1160 (O_1160,N_14994,N_14885);
nor UO_1161 (O_1161,N_14936,N_14935);
and UO_1162 (O_1162,N_14806,N_14809);
xnor UO_1163 (O_1163,N_14996,N_14948);
or UO_1164 (O_1164,N_14987,N_14994);
nor UO_1165 (O_1165,N_14909,N_14930);
and UO_1166 (O_1166,N_14853,N_14939);
or UO_1167 (O_1167,N_14914,N_14804);
nor UO_1168 (O_1168,N_14871,N_14808);
or UO_1169 (O_1169,N_14855,N_14840);
or UO_1170 (O_1170,N_14985,N_14982);
nor UO_1171 (O_1171,N_14950,N_14884);
or UO_1172 (O_1172,N_14986,N_14873);
and UO_1173 (O_1173,N_14908,N_14802);
nor UO_1174 (O_1174,N_14800,N_14906);
xnor UO_1175 (O_1175,N_14999,N_14840);
and UO_1176 (O_1176,N_14823,N_14926);
nand UO_1177 (O_1177,N_14838,N_14808);
nand UO_1178 (O_1178,N_14997,N_14833);
xnor UO_1179 (O_1179,N_14986,N_14831);
xnor UO_1180 (O_1180,N_14810,N_14826);
xnor UO_1181 (O_1181,N_14898,N_14966);
and UO_1182 (O_1182,N_14825,N_14927);
nand UO_1183 (O_1183,N_14926,N_14857);
nand UO_1184 (O_1184,N_14803,N_14951);
and UO_1185 (O_1185,N_14817,N_14930);
nand UO_1186 (O_1186,N_14888,N_14822);
and UO_1187 (O_1187,N_14869,N_14873);
and UO_1188 (O_1188,N_14935,N_14902);
and UO_1189 (O_1189,N_14968,N_14917);
or UO_1190 (O_1190,N_14849,N_14810);
nand UO_1191 (O_1191,N_14849,N_14876);
and UO_1192 (O_1192,N_14844,N_14868);
or UO_1193 (O_1193,N_14877,N_14961);
or UO_1194 (O_1194,N_14979,N_14868);
and UO_1195 (O_1195,N_14844,N_14882);
nor UO_1196 (O_1196,N_14950,N_14963);
nor UO_1197 (O_1197,N_14833,N_14900);
xor UO_1198 (O_1198,N_14924,N_14815);
nor UO_1199 (O_1199,N_14992,N_14854);
nor UO_1200 (O_1200,N_14925,N_14963);
nor UO_1201 (O_1201,N_14945,N_14955);
nor UO_1202 (O_1202,N_14932,N_14818);
xor UO_1203 (O_1203,N_14946,N_14847);
nand UO_1204 (O_1204,N_14925,N_14912);
nor UO_1205 (O_1205,N_14839,N_14859);
nor UO_1206 (O_1206,N_14967,N_14924);
nand UO_1207 (O_1207,N_14824,N_14840);
nor UO_1208 (O_1208,N_14901,N_14965);
nor UO_1209 (O_1209,N_14863,N_14888);
and UO_1210 (O_1210,N_14934,N_14827);
nand UO_1211 (O_1211,N_14917,N_14969);
nor UO_1212 (O_1212,N_14925,N_14843);
and UO_1213 (O_1213,N_14920,N_14834);
nand UO_1214 (O_1214,N_14848,N_14908);
nor UO_1215 (O_1215,N_14966,N_14930);
or UO_1216 (O_1216,N_14957,N_14954);
nor UO_1217 (O_1217,N_14810,N_14935);
xor UO_1218 (O_1218,N_14846,N_14989);
and UO_1219 (O_1219,N_14907,N_14884);
or UO_1220 (O_1220,N_14945,N_14934);
and UO_1221 (O_1221,N_14960,N_14834);
nor UO_1222 (O_1222,N_14954,N_14848);
or UO_1223 (O_1223,N_14820,N_14930);
xnor UO_1224 (O_1224,N_14935,N_14924);
or UO_1225 (O_1225,N_14809,N_14877);
nor UO_1226 (O_1226,N_14950,N_14930);
or UO_1227 (O_1227,N_14823,N_14838);
nor UO_1228 (O_1228,N_14979,N_14861);
xnor UO_1229 (O_1229,N_14882,N_14981);
or UO_1230 (O_1230,N_14837,N_14900);
or UO_1231 (O_1231,N_14877,N_14931);
xor UO_1232 (O_1232,N_14810,N_14860);
xnor UO_1233 (O_1233,N_14813,N_14994);
nor UO_1234 (O_1234,N_14830,N_14874);
nor UO_1235 (O_1235,N_14967,N_14989);
nor UO_1236 (O_1236,N_14997,N_14922);
nand UO_1237 (O_1237,N_14939,N_14983);
nand UO_1238 (O_1238,N_14857,N_14850);
nor UO_1239 (O_1239,N_14928,N_14896);
or UO_1240 (O_1240,N_14831,N_14912);
and UO_1241 (O_1241,N_14928,N_14951);
or UO_1242 (O_1242,N_14970,N_14973);
nand UO_1243 (O_1243,N_14971,N_14805);
xor UO_1244 (O_1244,N_14879,N_14940);
nand UO_1245 (O_1245,N_14817,N_14803);
and UO_1246 (O_1246,N_14902,N_14834);
xor UO_1247 (O_1247,N_14929,N_14862);
or UO_1248 (O_1248,N_14975,N_14875);
nor UO_1249 (O_1249,N_14968,N_14989);
nand UO_1250 (O_1250,N_14820,N_14871);
and UO_1251 (O_1251,N_14871,N_14852);
nand UO_1252 (O_1252,N_14804,N_14809);
nor UO_1253 (O_1253,N_14860,N_14986);
and UO_1254 (O_1254,N_14829,N_14908);
nand UO_1255 (O_1255,N_14965,N_14953);
xnor UO_1256 (O_1256,N_14998,N_14946);
nor UO_1257 (O_1257,N_14977,N_14997);
xor UO_1258 (O_1258,N_14845,N_14901);
and UO_1259 (O_1259,N_14992,N_14872);
nand UO_1260 (O_1260,N_14881,N_14955);
nand UO_1261 (O_1261,N_14980,N_14851);
or UO_1262 (O_1262,N_14927,N_14858);
xor UO_1263 (O_1263,N_14999,N_14986);
and UO_1264 (O_1264,N_14860,N_14997);
and UO_1265 (O_1265,N_14909,N_14836);
or UO_1266 (O_1266,N_14997,N_14882);
or UO_1267 (O_1267,N_14826,N_14848);
or UO_1268 (O_1268,N_14919,N_14893);
or UO_1269 (O_1269,N_14968,N_14969);
nand UO_1270 (O_1270,N_14843,N_14894);
nand UO_1271 (O_1271,N_14823,N_14954);
and UO_1272 (O_1272,N_14950,N_14994);
xnor UO_1273 (O_1273,N_14925,N_14980);
xnor UO_1274 (O_1274,N_14947,N_14990);
or UO_1275 (O_1275,N_14975,N_14992);
nand UO_1276 (O_1276,N_14850,N_14896);
nor UO_1277 (O_1277,N_14867,N_14927);
xnor UO_1278 (O_1278,N_14906,N_14828);
xor UO_1279 (O_1279,N_14925,N_14920);
nor UO_1280 (O_1280,N_14953,N_14919);
nor UO_1281 (O_1281,N_14890,N_14896);
xor UO_1282 (O_1282,N_14967,N_14971);
nor UO_1283 (O_1283,N_14811,N_14959);
or UO_1284 (O_1284,N_14877,N_14965);
xor UO_1285 (O_1285,N_14806,N_14867);
or UO_1286 (O_1286,N_14801,N_14999);
nand UO_1287 (O_1287,N_14835,N_14818);
and UO_1288 (O_1288,N_14872,N_14998);
and UO_1289 (O_1289,N_14816,N_14844);
and UO_1290 (O_1290,N_14894,N_14999);
xor UO_1291 (O_1291,N_14801,N_14809);
or UO_1292 (O_1292,N_14858,N_14906);
xnor UO_1293 (O_1293,N_14942,N_14831);
xor UO_1294 (O_1294,N_14820,N_14966);
and UO_1295 (O_1295,N_14858,N_14806);
and UO_1296 (O_1296,N_14818,N_14881);
xnor UO_1297 (O_1297,N_14913,N_14879);
nor UO_1298 (O_1298,N_14887,N_14972);
or UO_1299 (O_1299,N_14832,N_14957);
or UO_1300 (O_1300,N_14844,N_14950);
nand UO_1301 (O_1301,N_14953,N_14897);
xnor UO_1302 (O_1302,N_14819,N_14884);
nand UO_1303 (O_1303,N_14830,N_14825);
and UO_1304 (O_1304,N_14899,N_14987);
xnor UO_1305 (O_1305,N_14891,N_14804);
and UO_1306 (O_1306,N_14979,N_14938);
nand UO_1307 (O_1307,N_14832,N_14843);
or UO_1308 (O_1308,N_14891,N_14968);
and UO_1309 (O_1309,N_14915,N_14934);
nor UO_1310 (O_1310,N_14943,N_14971);
and UO_1311 (O_1311,N_14960,N_14931);
xor UO_1312 (O_1312,N_14907,N_14946);
xnor UO_1313 (O_1313,N_14981,N_14817);
nor UO_1314 (O_1314,N_14938,N_14953);
nor UO_1315 (O_1315,N_14845,N_14883);
nor UO_1316 (O_1316,N_14936,N_14814);
xor UO_1317 (O_1317,N_14925,N_14907);
and UO_1318 (O_1318,N_14977,N_14917);
nand UO_1319 (O_1319,N_14905,N_14855);
nand UO_1320 (O_1320,N_14858,N_14847);
or UO_1321 (O_1321,N_14803,N_14936);
nor UO_1322 (O_1322,N_14960,N_14976);
xor UO_1323 (O_1323,N_14871,N_14921);
or UO_1324 (O_1324,N_14872,N_14916);
nor UO_1325 (O_1325,N_14901,N_14926);
nor UO_1326 (O_1326,N_14951,N_14918);
xnor UO_1327 (O_1327,N_14904,N_14867);
nor UO_1328 (O_1328,N_14850,N_14898);
xor UO_1329 (O_1329,N_14801,N_14910);
xnor UO_1330 (O_1330,N_14909,N_14813);
nand UO_1331 (O_1331,N_14801,N_14985);
and UO_1332 (O_1332,N_14927,N_14972);
xnor UO_1333 (O_1333,N_14885,N_14860);
nor UO_1334 (O_1334,N_14956,N_14823);
nor UO_1335 (O_1335,N_14965,N_14806);
and UO_1336 (O_1336,N_14896,N_14895);
xnor UO_1337 (O_1337,N_14964,N_14840);
or UO_1338 (O_1338,N_14929,N_14837);
and UO_1339 (O_1339,N_14871,N_14905);
or UO_1340 (O_1340,N_14896,N_14828);
and UO_1341 (O_1341,N_14868,N_14967);
nand UO_1342 (O_1342,N_14857,N_14895);
or UO_1343 (O_1343,N_14986,N_14949);
and UO_1344 (O_1344,N_14869,N_14934);
and UO_1345 (O_1345,N_14912,N_14878);
and UO_1346 (O_1346,N_14916,N_14845);
nand UO_1347 (O_1347,N_14845,N_14920);
nor UO_1348 (O_1348,N_14811,N_14979);
nor UO_1349 (O_1349,N_14807,N_14831);
nor UO_1350 (O_1350,N_14874,N_14887);
xor UO_1351 (O_1351,N_14835,N_14891);
or UO_1352 (O_1352,N_14807,N_14956);
or UO_1353 (O_1353,N_14956,N_14830);
nor UO_1354 (O_1354,N_14815,N_14835);
or UO_1355 (O_1355,N_14906,N_14917);
xnor UO_1356 (O_1356,N_14982,N_14836);
or UO_1357 (O_1357,N_14901,N_14994);
nand UO_1358 (O_1358,N_14906,N_14950);
nand UO_1359 (O_1359,N_14854,N_14817);
or UO_1360 (O_1360,N_14863,N_14821);
nor UO_1361 (O_1361,N_14956,N_14875);
or UO_1362 (O_1362,N_14969,N_14816);
nand UO_1363 (O_1363,N_14931,N_14968);
and UO_1364 (O_1364,N_14966,N_14925);
or UO_1365 (O_1365,N_14884,N_14878);
and UO_1366 (O_1366,N_14904,N_14856);
and UO_1367 (O_1367,N_14994,N_14872);
nor UO_1368 (O_1368,N_14867,N_14821);
and UO_1369 (O_1369,N_14906,N_14954);
xnor UO_1370 (O_1370,N_14853,N_14960);
and UO_1371 (O_1371,N_14801,N_14930);
nor UO_1372 (O_1372,N_14979,N_14823);
nor UO_1373 (O_1373,N_14879,N_14890);
xor UO_1374 (O_1374,N_14875,N_14877);
and UO_1375 (O_1375,N_14817,N_14928);
or UO_1376 (O_1376,N_14849,N_14890);
or UO_1377 (O_1377,N_14849,N_14948);
and UO_1378 (O_1378,N_14967,N_14850);
nand UO_1379 (O_1379,N_14812,N_14936);
xor UO_1380 (O_1380,N_14849,N_14816);
or UO_1381 (O_1381,N_14979,N_14831);
nor UO_1382 (O_1382,N_14933,N_14942);
nand UO_1383 (O_1383,N_14941,N_14895);
and UO_1384 (O_1384,N_14959,N_14895);
and UO_1385 (O_1385,N_14851,N_14836);
nor UO_1386 (O_1386,N_14892,N_14909);
nand UO_1387 (O_1387,N_14964,N_14821);
and UO_1388 (O_1388,N_14937,N_14948);
nand UO_1389 (O_1389,N_14867,N_14801);
nor UO_1390 (O_1390,N_14916,N_14823);
or UO_1391 (O_1391,N_14871,N_14802);
and UO_1392 (O_1392,N_14868,N_14892);
xor UO_1393 (O_1393,N_14893,N_14881);
and UO_1394 (O_1394,N_14985,N_14824);
nor UO_1395 (O_1395,N_14897,N_14858);
xor UO_1396 (O_1396,N_14954,N_14936);
or UO_1397 (O_1397,N_14933,N_14920);
xnor UO_1398 (O_1398,N_14806,N_14857);
nand UO_1399 (O_1399,N_14882,N_14988);
nor UO_1400 (O_1400,N_14972,N_14846);
nor UO_1401 (O_1401,N_14851,N_14895);
nor UO_1402 (O_1402,N_14918,N_14919);
or UO_1403 (O_1403,N_14983,N_14966);
nor UO_1404 (O_1404,N_14842,N_14805);
or UO_1405 (O_1405,N_14905,N_14877);
xor UO_1406 (O_1406,N_14879,N_14952);
nor UO_1407 (O_1407,N_14993,N_14884);
nand UO_1408 (O_1408,N_14969,N_14860);
nand UO_1409 (O_1409,N_14990,N_14830);
and UO_1410 (O_1410,N_14985,N_14977);
nand UO_1411 (O_1411,N_14852,N_14837);
xnor UO_1412 (O_1412,N_14872,N_14943);
and UO_1413 (O_1413,N_14885,N_14964);
or UO_1414 (O_1414,N_14880,N_14945);
and UO_1415 (O_1415,N_14862,N_14870);
nand UO_1416 (O_1416,N_14893,N_14934);
nand UO_1417 (O_1417,N_14897,N_14854);
nor UO_1418 (O_1418,N_14854,N_14872);
nor UO_1419 (O_1419,N_14923,N_14858);
and UO_1420 (O_1420,N_14846,N_14992);
and UO_1421 (O_1421,N_14879,N_14905);
or UO_1422 (O_1422,N_14886,N_14824);
xor UO_1423 (O_1423,N_14917,N_14893);
xor UO_1424 (O_1424,N_14967,N_14931);
or UO_1425 (O_1425,N_14929,N_14961);
nand UO_1426 (O_1426,N_14877,N_14816);
xor UO_1427 (O_1427,N_14946,N_14875);
nand UO_1428 (O_1428,N_14854,N_14885);
nor UO_1429 (O_1429,N_14877,N_14869);
nand UO_1430 (O_1430,N_14953,N_14958);
and UO_1431 (O_1431,N_14900,N_14991);
and UO_1432 (O_1432,N_14819,N_14912);
and UO_1433 (O_1433,N_14844,N_14889);
or UO_1434 (O_1434,N_14843,N_14957);
or UO_1435 (O_1435,N_14828,N_14916);
and UO_1436 (O_1436,N_14939,N_14909);
nand UO_1437 (O_1437,N_14804,N_14916);
nand UO_1438 (O_1438,N_14896,N_14892);
and UO_1439 (O_1439,N_14811,N_14863);
xor UO_1440 (O_1440,N_14869,N_14942);
nand UO_1441 (O_1441,N_14857,N_14931);
nand UO_1442 (O_1442,N_14888,N_14917);
and UO_1443 (O_1443,N_14897,N_14816);
nand UO_1444 (O_1444,N_14970,N_14835);
nand UO_1445 (O_1445,N_14903,N_14987);
nor UO_1446 (O_1446,N_14875,N_14895);
nor UO_1447 (O_1447,N_14892,N_14830);
and UO_1448 (O_1448,N_14834,N_14819);
nand UO_1449 (O_1449,N_14921,N_14900);
nand UO_1450 (O_1450,N_14851,N_14869);
xnor UO_1451 (O_1451,N_14961,N_14896);
or UO_1452 (O_1452,N_14986,N_14888);
or UO_1453 (O_1453,N_14984,N_14908);
and UO_1454 (O_1454,N_14828,N_14915);
nor UO_1455 (O_1455,N_14980,N_14957);
or UO_1456 (O_1456,N_14808,N_14994);
nand UO_1457 (O_1457,N_14803,N_14973);
nor UO_1458 (O_1458,N_14896,N_14911);
or UO_1459 (O_1459,N_14967,N_14906);
and UO_1460 (O_1460,N_14910,N_14825);
xnor UO_1461 (O_1461,N_14962,N_14998);
nor UO_1462 (O_1462,N_14888,N_14997);
or UO_1463 (O_1463,N_14896,N_14834);
xnor UO_1464 (O_1464,N_14897,N_14941);
nand UO_1465 (O_1465,N_14845,N_14894);
and UO_1466 (O_1466,N_14999,N_14874);
and UO_1467 (O_1467,N_14844,N_14905);
xor UO_1468 (O_1468,N_14805,N_14861);
or UO_1469 (O_1469,N_14915,N_14809);
and UO_1470 (O_1470,N_14844,N_14870);
xor UO_1471 (O_1471,N_14865,N_14996);
or UO_1472 (O_1472,N_14936,N_14822);
nand UO_1473 (O_1473,N_14818,N_14806);
and UO_1474 (O_1474,N_14914,N_14856);
and UO_1475 (O_1475,N_14942,N_14801);
nor UO_1476 (O_1476,N_14977,N_14894);
xnor UO_1477 (O_1477,N_14871,N_14908);
and UO_1478 (O_1478,N_14884,N_14834);
and UO_1479 (O_1479,N_14945,N_14928);
and UO_1480 (O_1480,N_14931,N_14830);
nor UO_1481 (O_1481,N_14813,N_14814);
xor UO_1482 (O_1482,N_14943,N_14916);
nand UO_1483 (O_1483,N_14862,N_14883);
or UO_1484 (O_1484,N_14853,N_14952);
nand UO_1485 (O_1485,N_14972,N_14880);
nor UO_1486 (O_1486,N_14946,N_14892);
nor UO_1487 (O_1487,N_14928,N_14954);
nand UO_1488 (O_1488,N_14982,N_14804);
nand UO_1489 (O_1489,N_14931,N_14871);
nand UO_1490 (O_1490,N_14922,N_14947);
nand UO_1491 (O_1491,N_14981,N_14953);
nand UO_1492 (O_1492,N_14992,N_14817);
and UO_1493 (O_1493,N_14893,N_14832);
or UO_1494 (O_1494,N_14908,N_14926);
or UO_1495 (O_1495,N_14863,N_14900);
xor UO_1496 (O_1496,N_14940,N_14991);
xnor UO_1497 (O_1497,N_14850,N_14866);
nor UO_1498 (O_1498,N_14828,N_14910);
nand UO_1499 (O_1499,N_14976,N_14894);
xnor UO_1500 (O_1500,N_14822,N_14912);
or UO_1501 (O_1501,N_14848,N_14853);
nand UO_1502 (O_1502,N_14845,N_14977);
xor UO_1503 (O_1503,N_14929,N_14917);
or UO_1504 (O_1504,N_14909,N_14966);
or UO_1505 (O_1505,N_14912,N_14848);
nand UO_1506 (O_1506,N_14866,N_14949);
and UO_1507 (O_1507,N_14854,N_14831);
nand UO_1508 (O_1508,N_14904,N_14857);
nand UO_1509 (O_1509,N_14948,N_14843);
and UO_1510 (O_1510,N_14889,N_14836);
or UO_1511 (O_1511,N_14891,N_14999);
nor UO_1512 (O_1512,N_14933,N_14960);
nand UO_1513 (O_1513,N_14903,N_14979);
xor UO_1514 (O_1514,N_14949,N_14879);
or UO_1515 (O_1515,N_14849,N_14934);
nand UO_1516 (O_1516,N_14868,N_14874);
xor UO_1517 (O_1517,N_14986,N_14856);
and UO_1518 (O_1518,N_14926,N_14987);
xnor UO_1519 (O_1519,N_14970,N_14855);
or UO_1520 (O_1520,N_14908,N_14992);
xor UO_1521 (O_1521,N_14815,N_14966);
nand UO_1522 (O_1522,N_14866,N_14923);
nand UO_1523 (O_1523,N_14806,N_14930);
xnor UO_1524 (O_1524,N_14989,N_14924);
nor UO_1525 (O_1525,N_14836,N_14995);
and UO_1526 (O_1526,N_14852,N_14827);
and UO_1527 (O_1527,N_14869,N_14927);
and UO_1528 (O_1528,N_14871,N_14943);
or UO_1529 (O_1529,N_14984,N_14836);
and UO_1530 (O_1530,N_14972,N_14961);
nand UO_1531 (O_1531,N_14836,N_14893);
or UO_1532 (O_1532,N_14888,N_14925);
or UO_1533 (O_1533,N_14826,N_14845);
and UO_1534 (O_1534,N_14889,N_14981);
nor UO_1535 (O_1535,N_14915,N_14867);
nand UO_1536 (O_1536,N_14842,N_14927);
xor UO_1537 (O_1537,N_14925,N_14985);
nor UO_1538 (O_1538,N_14873,N_14800);
xnor UO_1539 (O_1539,N_14963,N_14971);
and UO_1540 (O_1540,N_14805,N_14818);
nand UO_1541 (O_1541,N_14828,N_14981);
or UO_1542 (O_1542,N_14805,N_14913);
nor UO_1543 (O_1543,N_14801,N_14826);
or UO_1544 (O_1544,N_14826,N_14918);
or UO_1545 (O_1545,N_14925,N_14917);
nor UO_1546 (O_1546,N_14930,N_14836);
and UO_1547 (O_1547,N_14940,N_14895);
xnor UO_1548 (O_1548,N_14857,N_14922);
or UO_1549 (O_1549,N_14927,N_14971);
xor UO_1550 (O_1550,N_14832,N_14918);
or UO_1551 (O_1551,N_14935,N_14812);
nor UO_1552 (O_1552,N_14997,N_14868);
xor UO_1553 (O_1553,N_14849,N_14939);
xor UO_1554 (O_1554,N_14856,N_14838);
xor UO_1555 (O_1555,N_14925,N_14968);
nand UO_1556 (O_1556,N_14978,N_14917);
nand UO_1557 (O_1557,N_14958,N_14877);
and UO_1558 (O_1558,N_14996,N_14936);
nor UO_1559 (O_1559,N_14859,N_14925);
or UO_1560 (O_1560,N_14811,N_14866);
xnor UO_1561 (O_1561,N_14955,N_14849);
and UO_1562 (O_1562,N_14861,N_14968);
nor UO_1563 (O_1563,N_14965,N_14844);
or UO_1564 (O_1564,N_14808,N_14972);
or UO_1565 (O_1565,N_14971,N_14833);
xnor UO_1566 (O_1566,N_14857,N_14961);
or UO_1567 (O_1567,N_14910,N_14947);
nor UO_1568 (O_1568,N_14858,N_14992);
or UO_1569 (O_1569,N_14999,N_14869);
nand UO_1570 (O_1570,N_14910,N_14926);
xor UO_1571 (O_1571,N_14999,N_14937);
xnor UO_1572 (O_1572,N_14857,N_14892);
and UO_1573 (O_1573,N_14838,N_14992);
and UO_1574 (O_1574,N_14956,N_14828);
nand UO_1575 (O_1575,N_14929,N_14960);
and UO_1576 (O_1576,N_14894,N_14978);
nor UO_1577 (O_1577,N_14857,N_14943);
and UO_1578 (O_1578,N_14871,N_14986);
xnor UO_1579 (O_1579,N_14864,N_14949);
nor UO_1580 (O_1580,N_14912,N_14970);
and UO_1581 (O_1581,N_14887,N_14844);
nor UO_1582 (O_1582,N_14810,N_14987);
nor UO_1583 (O_1583,N_14810,N_14878);
or UO_1584 (O_1584,N_14813,N_14878);
nor UO_1585 (O_1585,N_14951,N_14892);
or UO_1586 (O_1586,N_14845,N_14819);
xnor UO_1587 (O_1587,N_14958,N_14853);
nand UO_1588 (O_1588,N_14838,N_14850);
and UO_1589 (O_1589,N_14994,N_14831);
nor UO_1590 (O_1590,N_14933,N_14810);
or UO_1591 (O_1591,N_14932,N_14979);
nor UO_1592 (O_1592,N_14968,N_14862);
and UO_1593 (O_1593,N_14996,N_14879);
or UO_1594 (O_1594,N_14956,N_14862);
xor UO_1595 (O_1595,N_14934,N_14943);
nor UO_1596 (O_1596,N_14954,N_14935);
and UO_1597 (O_1597,N_14948,N_14802);
nand UO_1598 (O_1598,N_14842,N_14975);
xor UO_1599 (O_1599,N_14987,N_14886);
nand UO_1600 (O_1600,N_14889,N_14961);
xnor UO_1601 (O_1601,N_14907,N_14896);
nand UO_1602 (O_1602,N_14871,N_14982);
and UO_1603 (O_1603,N_14817,N_14801);
or UO_1604 (O_1604,N_14922,N_14817);
or UO_1605 (O_1605,N_14952,N_14990);
nand UO_1606 (O_1606,N_14946,N_14804);
xnor UO_1607 (O_1607,N_14914,N_14896);
and UO_1608 (O_1608,N_14859,N_14929);
nor UO_1609 (O_1609,N_14844,N_14996);
or UO_1610 (O_1610,N_14857,N_14914);
nand UO_1611 (O_1611,N_14888,N_14967);
xnor UO_1612 (O_1612,N_14913,N_14922);
xor UO_1613 (O_1613,N_14950,N_14905);
nand UO_1614 (O_1614,N_14947,N_14970);
or UO_1615 (O_1615,N_14970,N_14862);
or UO_1616 (O_1616,N_14854,N_14917);
and UO_1617 (O_1617,N_14870,N_14815);
or UO_1618 (O_1618,N_14948,N_14814);
and UO_1619 (O_1619,N_14998,N_14885);
or UO_1620 (O_1620,N_14951,N_14902);
nor UO_1621 (O_1621,N_14972,N_14854);
nand UO_1622 (O_1622,N_14907,N_14865);
nand UO_1623 (O_1623,N_14907,N_14850);
xor UO_1624 (O_1624,N_14936,N_14834);
or UO_1625 (O_1625,N_14838,N_14896);
or UO_1626 (O_1626,N_14891,N_14935);
or UO_1627 (O_1627,N_14966,N_14956);
nor UO_1628 (O_1628,N_14924,N_14823);
or UO_1629 (O_1629,N_14941,N_14802);
or UO_1630 (O_1630,N_14948,N_14804);
nand UO_1631 (O_1631,N_14921,N_14890);
nand UO_1632 (O_1632,N_14908,N_14922);
nand UO_1633 (O_1633,N_14845,N_14857);
xor UO_1634 (O_1634,N_14910,N_14902);
and UO_1635 (O_1635,N_14813,N_14971);
or UO_1636 (O_1636,N_14876,N_14812);
nor UO_1637 (O_1637,N_14900,N_14895);
and UO_1638 (O_1638,N_14904,N_14811);
or UO_1639 (O_1639,N_14878,N_14851);
xor UO_1640 (O_1640,N_14881,N_14862);
nand UO_1641 (O_1641,N_14900,N_14826);
nor UO_1642 (O_1642,N_14930,N_14949);
and UO_1643 (O_1643,N_14868,N_14893);
and UO_1644 (O_1644,N_14929,N_14844);
or UO_1645 (O_1645,N_14805,N_14988);
nor UO_1646 (O_1646,N_14907,N_14919);
or UO_1647 (O_1647,N_14853,N_14849);
xnor UO_1648 (O_1648,N_14966,N_14935);
nor UO_1649 (O_1649,N_14976,N_14900);
xor UO_1650 (O_1650,N_14938,N_14929);
nand UO_1651 (O_1651,N_14973,N_14942);
or UO_1652 (O_1652,N_14809,N_14892);
or UO_1653 (O_1653,N_14931,N_14978);
and UO_1654 (O_1654,N_14924,N_14812);
or UO_1655 (O_1655,N_14879,N_14957);
xor UO_1656 (O_1656,N_14876,N_14820);
and UO_1657 (O_1657,N_14939,N_14936);
nand UO_1658 (O_1658,N_14825,N_14928);
or UO_1659 (O_1659,N_14810,N_14840);
or UO_1660 (O_1660,N_14829,N_14845);
nand UO_1661 (O_1661,N_14807,N_14893);
xor UO_1662 (O_1662,N_14966,N_14918);
nor UO_1663 (O_1663,N_14830,N_14977);
and UO_1664 (O_1664,N_14803,N_14892);
xnor UO_1665 (O_1665,N_14826,N_14911);
nor UO_1666 (O_1666,N_14984,N_14881);
or UO_1667 (O_1667,N_14877,N_14979);
xnor UO_1668 (O_1668,N_14883,N_14966);
and UO_1669 (O_1669,N_14899,N_14893);
or UO_1670 (O_1670,N_14917,N_14975);
and UO_1671 (O_1671,N_14993,N_14809);
nor UO_1672 (O_1672,N_14828,N_14952);
nand UO_1673 (O_1673,N_14866,N_14904);
and UO_1674 (O_1674,N_14838,N_14983);
xnor UO_1675 (O_1675,N_14929,N_14868);
or UO_1676 (O_1676,N_14809,N_14814);
and UO_1677 (O_1677,N_14950,N_14801);
or UO_1678 (O_1678,N_14949,N_14920);
or UO_1679 (O_1679,N_14894,N_14815);
or UO_1680 (O_1680,N_14944,N_14870);
nor UO_1681 (O_1681,N_14865,N_14945);
nand UO_1682 (O_1682,N_14983,N_14862);
or UO_1683 (O_1683,N_14827,N_14965);
or UO_1684 (O_1684,N_14970,N_14925);
and UO_1685 (O_1685,N_14824,N_14943);
nor UO_1686 (O_1686,N_14882,N_14989);
nor UO_1687 (O_1687,N_14879,N_14907);
nand UO_1688 (O_1688,N_14954,N_14850);
and UO_1689 (O_1689,N_14950,N_14816);
or UO_1690 (O_1690,N_14840,N_14916);
or UO_1691 (O_1691,N_14856,N_14968);
and UO_1692 (O_1692,N_14851,N_14873);
nand UO_1693 (O_1693,N_14872,N_14989);
or UO_1694 (O_1694,N_14891,N_14939);
xnor UO_1695 (O_1695,N_14942,N_14819);
or UO_1696 (O_1696,N_14828,N_14808);
or UO_1697 (O_1697,N_14859,N_14806);
nor UO_1698 (O_1698,N_14833,N_14911);
nand UO_1699 (O_1699,N_14991,N_14968);
and UO_1700 (O_1700,N_14871,N_14849);
nor UO_1701 (O_1701,N_14895,N_14826);
or UO_1702 (O_1702,N_14852,N_14866);
and UO_1703 (O_1703,N_14849,N_14928);
nor UO_1704 (O_1704,N_14854,N_14842);
or UO_1705 (O_1705,N_14917,N_14891);
xor UO_1706 (O_1706,N_14944,N_14825);
nand UO_1707 (O_1707,N_14935,N_14944);
nand UO_1708 (O_1708,N_14869,N_14889);
and UO_1709 (O_1709,N_14975,N_14949);
xor UO_1710 (O_1710,N_14878,N_14877);
and UO_1711 (O_1711,N_14839,N_14848);
xnor UO_1712 (O_1712,N_14812,N_14803);
nand UO_1713 (O_1713,N_14973,N_14957);
nand UO_1714 (O_1714,N_14822,N_14838);
nor UO_1715 (O_1715,N_14948,N_14864);
and UO_1716 (O_1716,N_14805,N_14969);
xnor UO_1717 (O_1717,N_14871,N_14824);
xor UO_1718 (O_1718,N_14991,N_14980);
and UO_1719 (O_1719,N_14987,N_14894);
and UO_1720 (O_1720,N_14999,N_14825);
nand UO_1721 (O_1721,N_14970,N_14845);
or UO_1722 (O_1722,N_14992,N_14979);
nand UO_1723 (O_1723,N_14824,N_14863);
nand UO_1724 (O_1724,N_14866,N_14869);
nand UO_1725 (O_1725,N_14856,N_14832);
and UO_1726 (O_1726,N_14825,N_14809);
xnor UO_1727 (O_1727,N_14899,N_14887);
nor UO_1728 (O_1728,N_14809,N_14949);
and UO_1729 (O_1729,N_14968,N_14924);
nand UO_1730 (O_1730,N_14923,N_14981);
and UO_1731 (O_1731,N_14817,N_14908);
and UO_1732 (O_1732,N_14962,N_14826);
nor UO_1733 (O_1733,N_14889,N_14849);
nand UO_1734 (O_1734,N_14828,N_14962);
and UO_1735 (O_1735,N_14844,N_14920);
nor UO_1736 (O_1736,N_14909,N_14833);
xnor UO_1737 (O_1737,N_14885,N_14919);
nor UO_1738 (O_1738,N_14859,N_14913);
and UO_1739 (O_1739,N_14874,N_14943);
xor UO_1740 (O_1740,N_14980,N_14969);
xor UO_1741 (O_1741,N_14992,N_14939);
xor UO_1742 (O_1742,N_14999,N_14838);
and UO_1743 (O_1743,N_14889,N_14925);
or UO_1744 (O_1744,N_14830,N_14833);
and UO_1745 (O_1745,N_14883,N_14896);
nand UO_1746 (O_1746,N_14936,N_14949);
nor UO_1747 (O_1747,N_14837,N_14959);
nor UO_1748 (O_1748,N_14901,N_14836);
xnor UO_1749 (O_1749,N_14895,N_14842);
and UO_1750 (O_1750,N_14896,N_14954);
or UO_1751 (O_1751,N_14866,N_14840);
xor UO_1752 (O_1752,N_14806,N_14837);
or UO_1753 (O_1753,N_14843,N_14917);
nand UO_1754 (O_1754,N_14982,N_14847);
xor UO_1755 (O_1755,N_14983,N_14877);
nor UO_1756 (O_1756,N_14964,N_14818);
or UO_1757 (O_1757,N_14957,N_14812);
or UO_1758 (O_1758,N_14868,N_14839);
and UO_1759 (O_1759,N_14817,N_14969);
nor UO_1760 (O_1760,N_14924,N_14830);
nand UO_1761 (O_1761,N_14997,N_14974);
or UO_1762 (O_1762,N_14828,N_14973);
and UO_1763 (O_1763,N_14975,N_14897);
and UO_1764 (O_1764,N_14921,N_14984);
and UO_1765 (O_1765,N_14982,N_14860);
xnor UO_1766 (O_1766,N_14939,N_14927);
nand UO_1767 (O_1767,N_14876,N_14895);
or UO_1768 (O_1768,N_14971,N_14861);
nand UO_1769 (O_1769,N_14802,N_14886);
and UO_1770 (O_1770,N_14993,N_14875);
and UO_1771 (O_1771,N_14863,N_14858);
or UO_1772 (O_1772,N_14843,N_14981);
xor UO_1773 (O_1773,N_14813,N_14877);
nand UO_1774 (O_1774,N_14802,N_14971);
and UO_1775 (O_1775,N_14837,N_14872);
nand UO_1776 (O_1776,N_14978,N_14963);
or UO_1777 (O_1777,N_14965,N_14964);
or UO_1778 (O_1778,N_14817,N_14921);
and UO_1779 (O_1779,N_14833,N_14860);
nor UO_1780 (O_1780,N_14865,N_14868);
and UO_1781 (O_1781,N_14929,N_14916);
xnor UO_1782 (O_1782,N_14866,N_14992);
nor UO_1783 (O_1783,N_14972,N_14997);
nand UO_1784 (O_1784,N_14882,N_14897);
or UO_1785 (O_1785,N_14807,N_14890);
xor UO_1786 (O_1786,N_14874,N_14931);
nand UO_1787 (O_1787,N_14917,N_14866);
or UO_1788 (O_1788,N_14972,N_14859);
and UO_1789 (O_1789,N_14961,N_14997);
nand UO_1790 (O_1790,N_14886,N_14917);
and UO_1791 (O_1791,N_14865,N_14849);
or UO_1792 (O_1792,N_14984,N_14966);
nor UO_1793 (O_1793,N_14888,N_14887);
nor UO_1794 (O_1794,N_14854,N_14936);
nor UO_1795 (O_1795,N_14823,N_14953);
and UO_1796 (O_1796,N_14853,N_14950);
or UO_1797 (O_1797,N_14846,N_14921);
xor UO_1798 (O_1798,N_14943,N_14970);
and UO_1799 (O_1799,N_14929,N_14924);
nand UO_1800 (O_1800,N_14847,N_14944);
nand UO_1801 (O_1801,N_14889,N_14989);
xor UO_1802 (O_1802,N_14964,N_14930);
nor UO_1803 (O_1803,N_14842,N_14807);
nor UO_1804 (O_1804,N_14982,N_14977);
nand UO_1805 (O_1805,N_14946,N_14915);
xor UO_1806 (O_1806,N_14920,N_14945);
nor UO_1807 (O_1807,N_14931,N_14977);
nand UO_1808 (O_1808,N_14971,N_14882);
nand UO_1809 (O_1809,N_14996,N_14801);
nor UO_1810 (O_1810,N_14968,N_14868);
and UO_1811 (O_1811,N_14986,N_14815);
and UO_1812 (O_1812,N_14819,N_14905);
nand UO_1813 (O_1813,N_14810,N_14953);
or UO_1814 (O_1814,N_14939,N_14886);
nor UO_1815 (O_1815,N_14986,N_14809);
or UO_1816 (O_1816,N_14858,N_14854);
and UO_1817 (O_1817,N_14899,N_14845);
nand UO_1818 (O_1818,N_14919,N_14933);
and UO_1819 (O_1819,N_14863,N_14951);
nor UO_1820 (O_1820,N_14800,N_14991);
nor UO_1821 (O_1821,N_14846,N_14813);
xnor UO_1822 (O_1822,N_14882,N_14865);
nand UO_1823 (O_1823,N_14903,N_14842);
nand UO_1824 (O_1824,N_14823,N_14973);
xnor UO_1825 (O_1825,N_14934,N_14876);
nor UO_1826 (O_1826,N_14999,N_14971);
nor UO_1827 (O_1827,N_14860,N_14851);
nand UO_1828 (O_1828,N_14810,N_14962);
nand UO_1829 (O_1829,N_14820,N_14944);
or UO_1830 (O_1830,N_14898,N_14871);
nor UO_1831 (O_1831,N_14928,N_14995);
or UO_1832 (O_1832,N_14865,N_14969);
nand UO_1833 (O_1833,N_14891,N_14978);
or UO_1834 (O_1834,N_14864,N_14912);
nand UO_1835 (O_1835,N_14980,N_14891);
and UO_1836 (O_1836,N_14826,N_14886);
nor UO_1837 (O_1837,N_14959,N_14985);
nor UO_1838 (O_1838,N_14905,N_14841);
nand UO_1839 (O_1839,N_14823,N_14947);
nand UO_1840 (O_1840,N_14869,N_14872);
and UO_1841 (O_1841,N_14917,N_14934);
nor UO_1842 (O_1842,N_14837,N_14913);
xnor UO_1843 (O_1843,N_14909,N_14864);
xnor UO_1844 (O_1844,N_14957,N_14823);
xnor UO_1845 (O_1845,N_14855,N_14831);
and UO_1846 (O_1846,N_14999,N_14853);
and UO_1847 (O_1847,N_14978,N_14841);
xnor UO_1848 (O_1848,N_14826,N_14873);
nand UO_1849 (O_1849,N_14913,N_14952);
nor UO_1850 (O_1850,N_14817,N_14927);
nand UO_1851 (O_1851,N_14913,N_14920);
or UO_1852 (O_1852,N_14914,N_14912);
nand UO_1853 (O_1853,N_14863,N_14829);
and UO_1854 (O_1854,N_14921,N_14985);
xnor UO_1855 (O_1855,N_14902,N_14913);
xnor UO_1856 (O_1856,N_14935,N_14919);
nand UO_1857 (O_1857,N_14816,N_14963);
or UO_1858 (O_1858,N_14973,N_14988);
or UO_1859 (O_1859,N_14826,N_14932);
nand UO_1860 (O_1860,N_14999,N_14892);
or UO_1861 (O_1861,N_14856,N_14810);
or UO_1862 (O_1862,N_14869,N_14954);
nand UO_1863 (O_1863,N_14964,N_14839);
xor UO_1864 (O_1864,N_14992,N_14934);
nand UO_1865 (O_1865,N_14863,N_14850);
nor UO_1866 (O_1866,N_14969,N_14911);
xor UO_1867 (O_1867,N_14801,N_14816);
nand UO_1868 (O_1868,N_14913,N_14899);
or UO_1869 (O_1869,N_14850,N_14944);
nor UO_1870 (O_1870,N_14994,N_14832);
nand UO_1871 (O_1871,N_14924,N_14835);
and UO_1872 (O_1872,N_14960,N_14885);
or UO_1873 (O_1873,N_14826,N_14823);
xor UO_1874 (O_1874,N_14958,N_14822);
xor UO_1875 (O_1875,N_14857,N_14841);
xnor UO_1876 (O_1876,N_14923,N_14941);
and UO_1877 (O_1877,N_14994,N_14891);
nor UO_1878 (O_1878,N_14836,N_14953);
xor UO_1879 (O_1879,N_14893,N_14963);
nand UO_1880 (O_1880,N_14870,N_14951);
and UO_1881 (O_1881,N_14984,N_14844);
xor UO_1882 (O_1882,N_14815,N_14972);
xnor UO_1883 (O_1883,N_14849,N_14978);
nand UO_1884 (O_1884,N_14974,N_14842);
nand UO_1885 (O_1885,N_14946,N_14978);
nor UO_1886 (O_1886,N_14964,N_14905);
xor UO_1887 (O_1887,N_14816,N_14943);
and UO_1888 (O_1888,N_14907,N_14991);
and UO_1889 (O_1889,N_14996,N_14855);
xor UO_1890 (O_1890,N_14952,N_14907);
nand UO_1891 (O_1891,N_14993,N_14913);
or UO_1892 (O_1892,N_14878,N_14880);
and UO_1893 (O_1893,N_14960,N_14904);
xor UO_1894 (O_1894,N_14978,N_14980);
and UO_1895 (O_1895,N_14931,N_14918);
nand UO_1896 (O_1896,N_14959,N_14996);
nand UO_1897 (O_1897,N_14987,N_14973);
nor UO_1898 (O_1898,N_14818,N_14975);
nor UO_1899 (O_1899,N_14880,N_14904);
nand UO_1900 (O_1900,N_14961,N_14956);
nand UO_1901 (O_1901,N_14824,N_14810);
nand UO_1902 (O_1902,N_14835,N_14967);
nor UO_1903 (O_1903,N_14972,N_14913);
xor UO_1904 (O_1904,N_14988,N_14944);
xnor UO_1905 (O_1905,N_14868,N_14976);
or UO_1906 (O_1906,N_14922,N_14959);
xor UO_1907 (O_1907,N_14845,N_14873);
nor UO_1908 (O_1908,N_14899,N_14924);
and UO_1909 (O_1909,N_14953,N_14850);
nor UO_1910 (O_1910,N_14893,N_14871);
nor UO_1911 (O_1911,N_14861,N_14849);
nand UO_1912 (O_1912,N_14906,N_14979);
nand UO_1913 (O_1913,N_14989,N_14800);
xor UO_1914 (O_1914,N_14847,N_14917);
xor UO_1915 (O_1915,N_14879,N_14828);
nand UO_1916 (O_1916,N_14987,N_14997);
xor UO_1917 (O_1917,N_14910,N_14877);
or UO_1918 (O_1918,N_14878,N_14906);
or UO_1919 (O_1919,N_14833,N_14921);
and UO_1920 (O_1920,N_14859,N_14928);
xnor UO_1921 (O_1921,N_14809,N_14924);
nand UO_1922 (O_1922,N_14895,N_14908);
nand UO_1923 (O_1923,N_14996,N_14903);
or UO_1924 (O_1924,N_14878,N_14982);
or UO_1925 (O_1925,N_14981,N_14983);
xor UO_1926 (O_1926,N_14960,N_14832);
nand UO_1927 (O_1927,N_14843,N_14856);
and UO_1928 (O_1928,N_14917,N_14880);
xnor UO_1929 (O_1929,N_14980,N_14935);
nor UO_1930 (O_1930,N_14959,N_14818);
or UO_1931 (O_1931,N_14853,N_14841);
nand UO_1932 (O_1932,N_14943,N_14822);
or UO_1933 (O_1933,N_14977,N_14969);
nand UO_1934 (O_1934,N_14933,N_14983);
and UO_1935 (O_1935,N_14985,N_14827);
nand UO_1936 (O_1936,N_14995,N_14811);
xnor UO_1937 (O_1937,N_14843,N_14999);
and UO_1938 (O_1938,N_14889,N_14855);
xnor UO_1939 (O_1939,N_14843,N_14830);
and UO_1940 (O_1940,N_14847,N_14891);
or UO_1941 (O_1941,N_14826,N_14913);
and UO_1942 (O_1942,N_14882,N_14942);
nand UO_1943 (O_1943,N_14957,N_14854);
xnor UO_1944 (O_1944,N_14958,N_14930);
nor UO_1945 (O_1945,N_14893,N_14913);
nor UO_1946 (O_1946,N_14976,N_14861);
xor UO_1947 (O_1947,N_14824,N_14875);
or UO_1948 (O_1948,N_14857,N_14902);
nand UO_1949 (O_1949,N_14867,N_14837);
xnor UO_1950 (O_1950,N_14912,N_14943);
or UO_1951 (O_1951,N_14826,N_14987);
xor UO_1952 (O_1952,N_14980,N_14973);
nor UO_1953 (O_1953,N_14960,N_14813);
and UO_1954 (O_1954,N_14877,N_14894);
and UO_1955 (O_1955,N_14928,N_14886);
and UO_1956 (O_1956,N_14942,N_14980);
xnor UO_1957 (O_1957,N_14889,N_14894);
nor UO_1958 (O_1958,N_14901,N_14876);
nand UO_1959 (O_1959,N_14999,N_14950);
nand UO_1960 (O_1960,N_14867,N_14800);
nor UO_1961 (O_1961,N_14976,N_14884);
xor UO_1962 (O_1962,N_14860,N_14990);
or UO_1963 (O_1963,N_14822,N_14859);
xor UO_1964 (O_1964,N_14873,N_14882);
or UO_1965 (O_1965,N_14958,N_14811);
nand UO_1966 (O_1966,N_14831,N_14827);
xor UO_1967 (O_1967,N_14984,N_14987);
and UO_1968 (O_1968,N_14846,N_14917);
nand UO_1969 (O_1969,N_14821,N_14897);
and UO_1970 (O_1970,N_14851,N_14804);
nand UO_1971 (O_1971,N_14910,N_14835);
xor UO_1972 (O_1972,N_14948,N_14917);
or UO_1973 (O_1973,N_14822,N_14891);
xor UO_1974 (O_1974,N_14879,N_14998);
and UO_1975 (O_1975,N_14995,N_14845);
nor UO_1976 (O_1976,N_14807,N_14856);
nand UO_1977 (O_1977,N_14923,N_14851);
nand UO_1978 (O_1978,N_14984,N_14956);
nand UO_1979 (O_1979,N_14834,N_14990);
xnor UO_1980 (O_1980,N_14906,N_14896);
nor UO_1981 (O_1981,N_14830,N_14929);
nor UO_1982 (O_1982,N_14988,N_14835);
nand UO_1983 (O_1983,N_14872,N_14945);
nand UO_1984 (O_1984,N_14854,N_14805);
nand UO_1985 (O_1985,N_14801,N_14824);
xor UO_1986 (O_1986,N_14965,N_14998);
nand UO_1987 (O_1987,N_14963,N_14947);
nor UO_1988 (O_1988,N_14839,N_14936);
nor UO_1989 (O_1989,N_14856,N_14862);
nor UO_1990 (O_1990,N_14821,N_14827);
or UO_1991 (O_1991,N_14885,N_14863);
xnor UO_1992 (O_1992,N_14891,N_14987);
nor UO_1993 (O_1993,N_14888,N_14860);
or UO_1994 (O_1994,N_14853,N_14968);
nor UO_1995 (O_1995,N_14932,N_14858);
nor UO_1996 (O_1996,N_14810,N_14918);
nand UO_1997 (O_1997,N_14835,N_14862);
nand UO_1998 (O_1998,N_14980,N_14808);
and UO_1999 (O_1999,N_14957,N_14991);
endmodule