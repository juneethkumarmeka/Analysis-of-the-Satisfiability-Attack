module basic_500_3000_500_5_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_303,In_137);
nand U1 (N_1,In_285,In_11);
and U2 (N_2,In_220,In_152);
nand U3 (N_3,In_49,In_288);
nor U4 (N_4,In_144,In_440);
nand U5 (N_5,In_455,In_432);
and U6 (N_6,In_204,In_9);
nand U7 (N_7,In_145,In_372);
nand U8 (N_8,In_336,In_207);
and U9 (N_9,In_244,In_438);
or U10 (N_10,In_471,In_211);
or U11 (N_11,In_417,In_113);
nor U12 (N_12,In_369,In_305);
nor U13 (N_13,In_361,In_178);
and U14 (N_14,In_194,In_197);
or U15 (N_15,In_87,In_157);
nor U16 (N_16,In_266,In_86);
and U17 (N_17,In_402,In_57);
and U18 (N_18,In_460,In_163);
and U19 (N_19,In_279,In_7);
nor U20 (N_20,In_88,In_2);
nor U21 (N_21,In_184,In_232);
or U22 (N_22,In_387,In_325);
and U23 (N_23,In_381,In_323);
or U24 (N_24,In_100,In_287);
or U25 (N_25,In_248,In_456);
nand U26 (N_26,In_160,In_459);
nor U27 (N_27,In_332,In_185);
or U28 (N_28,In_154,In_312);
and U29 (N_29,In_4,In_403);
or U30 (N_30,In_482,In_379);
or U31 (N_31,In_259,In_40);
and U32 (N_32,In_71,In_498);
and U33 (N_33,In_291,In_179);
and U34 (N_34,In_223,In_231);
or U35 (N_35,In_156,In_173);
nand U36 (N_36,In_245,In_434);
and U37 (N_37,In_127,In_35);
or U38 (N_38,In_356,In_366);
and U39 (N_39,In_239,In_225);
nand U40 (N_40,In_147,In_300);
nand U41 (N_41,In_358,In_265);
and U42 (N_42,In_31,In_364);
nand U43 (N_43,In_380,In_481);
nand U44 (N_44,In_267,In_487);
nand U45 (N_45,In_110,In_66);
nand U46 (N_46,In_187,In_316);
and U47 (N_47,In_18,In_238);
nand U48 (N_48,In_202,In_492);
nor U49 (N_49,In_419,In_105);
nand U50 (N_50,In_52,In_404);
or U51 (N_51,In_335,In_409);
nor U52 (N_52,In_190,In_390);
nand U53 (N_53,In_345,In_118);
nor U54 (N_54,In_457,In_21);
or U55 (N_55,In_470,In_442);
nor U56 (N_56,In_129,In_67);
nand U57 (N_57,In_227,In_111);
nand U58 (N_58,In_472,In_339);
nor U59 (N_59,In_180,In_155);
nor U60 (N_60,In_447,In_191);
and U61 (N_61,In_495,In_75);
and U62 (N_62,In_469,In_277);
nor U63 (N_63,In_255,In_79);
nand U64 (N_64,In_50,In_315);
nor U65 (N_65,In_69,In_397);
and U66 (N_66,In_219,In_406);
nor U67 (N_67,In_450,In_437);
nor U68 (N_68,In_98,In_452);
nand U69 (N_69,In_422,In_47);
nor U70 (N_70,In_92,In_165);
nand U71 (N_71,In_373,In_85);
or U72 (N_72,In_334,In_148);
and U73 (N_73,In_273,In_424);
and U74 (N_74,In_213,In_65);
nor U75 (N_75,In_12,In_297);
nand U76 (N_76,In_443,In_107);
and U77 (N_77,In_410,In_493);
and U78 (N_78,In_427,In_188);
and U79 (N_79,In_269,In_331);
nand U80 (N_80,In_433,In_119);
or U81 (N_81,In_13,In_206);
or U82 (N_82,In_313,In_330);
and U83 (N_83,In_237,In_90);
and U84 (N_84,In_258,In_99);
nand U85 (N_85,In_476,In_264);
nor U86 (N_86,In_276,In_228);
and U87 (N_87,In_307,In_448);
nor U88 (N_88,In_63,In_242);
and U89 (N_89,In_278,In_272);
xor U90 (N_90,In_243,In_226);
nand U91 (N_91,In_172,In_344);
nor U92 (N_92,In_474,In_473);
nor U93 (N_93,In_186,In_169);
and U94 (N_94,In_195,In_193);
or U95 (N_95,In_143,In_435);
and U96 (N_96,In_382,In_221);
nor U97 (N_97,In_412,In_337);
or U98 (N_98,In_353,In_26);
nand U99 (N_99,In_347,In_27);
and U100 (N_100,In_138,In_91);
and U101 (N_101,In_8,In_396);
nand U102 (N_102,In_14,In_196);
or U103 (N_103,In_252,In_484);
nor U104 (N_104,In_109,In_420);
xor U105 (N_105,In_415,In_386);
nor U106 (N_106,In_400,In_200);
and U107 (N_107,In_296,In_384);
nor U108 (N_108,In_385,In_149);
nor U109 (N_109,In_230,In_496);
or U110 (N_110,In_10,In_314);
nor U111 (N_111,In_461,In_439);
nor U112 (N_112,In_399,In_341);
xnor U113 (N_113,In_25,In_262);
nand U114 (N_114,In_311,In_430);
or U115 (N_115,In_17,In_280);
and U116 (N_116,In_120,In_161);
nand U117 (N_117,In_451,In_168);
and U118 (N_118,In_189,In_141);
nand U119 (N_119,In_407,In_383);
or U120 (N_120,In_393,In_37);
nand U121 (N_121,In_458,In_254);
nor U122 (N_122,In_370,In_46);
and U123 (N_123,In_72,In_218);
and U124 (N_124,In_97,In_454);
nor U125 (N_125,In_68,In_104);
nor U126 (N_126,In_103,In_24);
nor U127 (N_127,In_44,In_411);
nor U128 (N_128,In_320,In_294);
nand U129 (N_129,In_449,In_122);
nor U130 (N_130,In_319,In_301);
or U131 (N_131,In_263,In_74);
or U132 (N_132,In_428,In_310);
nand U133 (N_133,In_181,In_249);
or U134 (N_134,In_414,In_233);
nand U135 (N_135,In_367,In_465);
and U136 (N_136,In_462,In_201);
nand U137 (N_137,In_94,In_328);
and U138 (N_138,In_241,In_36);
and U139 (N_139,In_229,In_464);
nand U140 (N_140,In_51,In_136);
nand U141 (N_141,In_253,In_298);
nor U142 (N_142,In_42,In_497);
and U143 (N_143,In_142,In_171);
nor U144 (N_144,In_453,In_81);
and U145 (N_145,In_284,In_56);
or U146 (N_146,In_485,In_215);
nor U147 (N_147,In_394,In_425);
or U148 (N_148,In_174,In_441);
and U149 (N_149,In_401,In_368);
nand U150 (N_150,In_43,In_283);
nand U151 (N_151,In_426,In_346);
or U152 (N_152,In_395,In_126);
or U153 (N_153,In_3,In_123);
nor U154 (N_154,In_96,In_480);
or U155 (N_155,In_479,In_32);
xnor U156 (N_156,In_29,In_256);
and U157 (N_157,In_117,In_392);
or U158 (N_158,In_116,In_159);
nand U159 (N_159,In_106,In_365);
or U160 (N_160,In_359,In_20);
nor U161 (N_161,In_61,In_483);
nand U162 (N_162,In_22,In_318);
or U163 (N_163,In_475,In_134);
nand U164 (N_164,In_349,In_139);
nand U165 (N_165,In_41,In_135);
and U166 (N_166,In_413,In_357);
or U167 (N_167,In_55,In_444);
nand U168 (N_168,In_302,In_342);
nand U169 (N_169,In_251,In_286);
nor U170 (N_170,In_131,In_445);
and U171 (N_171,In_234,In_355);
and U172 (N_172,In_321,In_130);
and U173 (N_173,In_375,In_374);
and U174 (N_174,In_153,In_309);
nand U175 (N_175,In_0,In_93);
nand U176 (N_176,In_6,In_140);
or U177 (N_177,In_33,In_209);
or U178 (N_178,In_16,In_95);
nand U179 (N_179,In_19,In_292);
nor U180 (N_180,In_224,In_102);
or U181 (N_181,In_491,In_377);
and U182 (N_182,In_70,In_360);
and U183 (N_183,In_261,In_468);
nand U184 (N_184,In_274,In_478);
nor U185 (N_185,In_490,In_175);
and U186 (N_186,In_282,In_133);
nor U187 (N_187,In_436,In_351);
and U188 (N_188,In_348,In_121);
or U189 (N_189,In_5,In_322);
xor U190 (N_190,In_371,In_378);
and U191 (N_191,In_376,In_408);
nand U192 (N_192,In_115,In_53);
and U193 (N_193,In_363,In_304);
or U194 (N_194,In_326,In_212);
xnor U195 (N_195,In_151,In_62);
nor U196 (N_196,In_210,In_290);
nand U197 (N_197,In_60,In_166);
nand U198 (N_198,In_317,In_80);
or U199 (N_199,In_340,In_48);
and U200 (N_200,In_329,In_308);
nand U201 (N_201,In_170,In_466);
nand U202 (N_202,In_73,In_240);
or U203 (N_203,In_198,In_34);
and U204 (N_204,In_236,In_362);
and U205 (N_205,In_158,In_306);
and U206 (N_206,In_208,In_418);
or U207 (N_207,In_176,In_352);
and U208 (N_208,In_494,In_271);
nor U209 (N_209,In_28,In_289);
nor U210 (N_210,In_84,In_343);
and U211 (N_211,In_101,In_295);
or U212 (N_212,In_124,In_389);
xor U213 (N_213,In_114,In_182);
and U214 (N_214,In_45,In_486);
nor U215 (N_215,In_112,In_83);
and U216 (N_216,In_78,In_77);
nor U217 (N_217,In_23,In_192);
and U218 (N_218,In_82,In_203);
xnor U219 (N_219,In_281,In_270);
and U220 (N_220,In_429,In_463);
and U221 (N_221,In_58,In_293);
and U222 (N_222,In_299,In_489);
nand U223 (N_223,In_128,In_216);
nand U224 (N_224,In_398,In_416);
xor U225 (N_225,In_132,In_30);
nand U226 (N_226,In_446,In_247);
and U227 (N_227,In_354,In_64);
nand U228 (N_228,In_217,In_327);
and U229 (N_229,In_205,In_214);
nand U230 (N_230,In_150,In_391);
nand U231 (N_231,In_125,In_388);
nand U232 (N_232,In_477,In_59);
nand U233 (N_233,In_235,In_324);
xor U234 (N_234,In_268,In_1);
and U235 (N_235,In_162,In_405);
xnor U236 (N_236,In_38,In_246);
nand U237 (N_237,In_333,In_39);
and U238 (N_238,In_183,In_164);
or U239 (N_239,In_431,In_177);
or U240 (N_240,In_89,In_421);
or U241 (N_241,In_260,In_467);
nor U242 (N_242,In_350,In_76);
nand U243 (N_243,In_250,In_257);
and U244 (N_244,In_338,In_167);
nor U245 (N_245,In_499,In_423);
nand U246 (N_246,In_15,In_108);
and U247 (N_247,In_146,In_54);
or U248 (N_248,In_488,In_222);
or U249 (N_249,In_275,In_199);
nand U250 (N_250,In_361,In_405);
nor U251 (N_251,In_369,In_55);
and U252 (N_252,In_269,In_375);
and U253 (N_253,In_325,In_214);
nor U254 (N_254,In_258,In_191);
or U255 (N_255,In_74,In_224);
or U256 (N_256,In_213,In_253);
nand U257 (N_257,In_309,In_124);
or U258 (N_258,In_356,In_168);
and U259 (N_259,In_445,In_495);
nand U260 (N_260,In_99,In_373);
xnor U261 (N_261,In_187,In_128);
or U262 (N_262,In_428,In_61);
xor U263 (N_263,In_230,In_258);
or U264 (N_264,In_100,In_67);
nand U265 (N_265,In_460,In_415);
nor U266 (N_266,In_197,In_449);
or U267 (N_267,In_45,In_182);
and U268 (N_268,In_147,In_58);
and U269 (N_269,In_56,In_100);
nand U270 (N_270,In_414,In_478);
nor U271 (N_271,In_496,In_167);
nand U272 (N_272,In_396,In_84);
nand U273 (N_273,In_407,In_358);
or U274 (N_274,In_40,In_136);
or U275 (N_275,In_179,In_359);
nand U276 (N_276,In_376,In_405);
or U277 (N_277,In_1,In_334);
nand U278 (N_278,In_318,In_486);
or U279 (N_279,In_275,In_247);
xnor U280 (N_280,In_347,In_344);
xnor U281 (N_281,In_89,In_59);
xor U282 (N_282,In_213,In_44);
and U283 (N_283,In_224,In_445);
nor U284 (N_284,In_168,In_358);
or U285 (N_285,In_267,In_362);
or U286 (N_286,In_119,In_100);
nand U287 (N_287,In_428,In_384);
or U288 (N_288,In_94,In_346);
xnor U289 (N_289,In_109,In_476);
and U290 (N_290,In_213,In_8);
xor U291 (N_291,In_247,In_61);
or U292 (N_292,In_401,In_45);
nand U293 (N_293,In_271,In_106);
nand U294 (N_294,In_209,In_76);
or U295 (N_295,In_292,In_124);
nand U296 (N_296,In_171,In_167);
nor U297 (N_297,In_383,In_227);
nor U298 (N_298,In_289,In_275);
and U299 (N_299,In_35,In_152);
nand U300 (N_300,In_68,In_57);
nor U301 (N_301,In_480,In_123);
or U302 (N_302,In_490,In_326);
or U303 (N_303,In_190,In_125);
or U304 (N_304,In_44,In_458);
nand U305 (N_305,In_85,In_343);
and U306 (N_306,In_51,In_206);
nand U307 (N_307,In_157,In_186);
nor U308 (N_308,In_84,In_196);
or U309 (N_309,In_284,In_137);
or U310 (N_310,In_307,In_46);
and U311 (N_311,In_387,In_155);
and U312 (N_312,In_342,In_314);
and U313 (N_313,In_478,In_190);
nor U314 (N_314,In_497,In_286);
and U315 (N_315,In_351,In_173);
xor U316 (N_316,In_42,In_432);
and U317 (N_317,In_328,In_316);
nor U318 (N_318,In_418,In_51);
nand U319 (N_319,In_270,In_242);
and U320 (N_320,In_295,In_494);
xnor U321 (N_321,In_146,In_265);
xor U322 (N_322,In_482,In_79);
nor U323 (N_323,In_65,In_127);
nor U324 (N_324,In_211,In_194);
xnor U325 (N_325,In_360,In_333);
and U326 (N_326,In_297,In_261);
nor U327 (N_327,In_224,In_85);
and U328 (N_328,In_374,In_350);
or U329 (N_329,In_383,In_304);
and U330 (N_330,In_113,In_316);
xnor U331 (N_331,In_286,In_134);
xnor U332 (N_332,In_209,In_91);
or U333 (N_333,In_364,In_44);
or U334 (N_334,In_367,In_126);
xnor U335 (N_335,In_392,In_443);
or U336 (N_336,In_272,In_416);
or U337 (N_337,In_23,In_14);
and U338 (N_338,In_103,In_360);
or U339 (N_339,In_142,In_228);
nand U340 (N_340,In_177,In_15);
or U341 (N_341,In_498,In_169);
nor U342 (N_342,In_328,In_69);
nor U343 (N_343,In_494,In_209);
or U344 (N_344,In_464,In_211);
nor U345 (N_345,In_307,In_63);
or U346 (N_346,In_456,In_92);
and U347 (N_347,In_437,In_353);
nand U348 (N_348,In_87,In_97);
nor U349 (N_349,In_82,In_311);
nor U350 (N_350,In_314,In_277);
nand U351 (N_351,In_376,In_383);
xor U352 (N_352,In_27,In_223);
nand U353 (N_353,In_36,In_440);
nand U354 (N_354,In_332,In_124);
nor U355 (N_355,In_162,In_20);
nand U356 (N_356,In_307,In_200);
nand U357 (N_357,In_238,In_470);
nor U358 (N_358,In_256,In_416);
and U359 (N_359,In_175,In_346);
or U360 (N_360,In_214,In_428);
and U361 (N_361,In_364,In_218);
nor U362 (N_362,In_355,In_240);
nand U363 (N_363,In_145,In_181);
nor U364 (N_364,In_380,In_311);
nor U365 (N_365,In_57,In_137);
nor U366 (N_366,In_116,In_439);
xor U367 (N_367,In_76,In_328);
and U368 (N_368,In_251,In_456);
or U369 (N_369,In_103,In_460);
or U370 (N_370,In_319,In_88);
and U371 (N_371,In_299,In_105);
and U372 (N_372,In_152,In_374);
or U373 (N_373,In_173,In_471);
xor U374 (N_374,In_121,In_70);
nor U375 (N_375,In_155,In_223);
or U376 (N_376,In_211,In_247);
and U377 (N_377,In_139,In_469);
or U378 (N_378,In_207,In_159);
nor U379 (N_379,In_163,In_357);
and U380 (N_380,In_365,In_471);
and U381 (N_381,In_48,In_216);
and U382 (N_382,In_303,In_256);
and U383 (N_383,In_371,In_62);
nand U384 (N_384,In_247,In_421);
nor U385 (N_385,In_115,In_202);
nor U386 (N_386,In_273,In_420);
nand U387 (N_387,In_330,In_230);
nand U388 (N_388,In_486,In_245);
and U389 (N_389,In_335,In_177);
or U390 (N_390,In_389,In_402);
or U391 (N_391,In_445,In_275);
xnor U392 (N_392,In_60,In_286);
xnor U393 (N_393,In_363,In_450);
and U394 (N_394,In_4,In_7);
nand U395 (N_395,In_313,In_474);
nor U396 (N_396,In_282,In_455);
nor U397 (N_397,In_293,In_454);
and U398 (N_398,In_280,In_51);
or U399 (N_399,In_18,In_42);
nor U400 (N_400,In_398,In_343);
nand U401 (N_401,In_334,In_115);
nor U402 (N_402,In_313,In_310);
xor U403 (N_403,In_396,In_98);
and U404 (N_404,In_205,In_115);
or U405 (N_405,In_256,In_150);
and U406 (N_406,In_472,In_360);
nor U407 (N_407,In_475,In_183);
nand U408 (N_408,In_157,In_478);
nand U409 (N_409,In_269,In_405);
and U410 (N_410,In_244,In_241);
xor U411 (N_411,In_128,In_139);
nand U412 (N_412,In_257,In_267);
or U413 (N_413,In_475,In_80);
nor U414 (N_414,In_292,In_248);
nor U415 (N_415,In_339,In_404);
xor U416 (N_416,In_274,In_179);
and U417 (N_417,In_156,In_77);
nand U418 (N_418,In_78,In_259);
or U419 (N_419,In_340,In_175);
nor U420 (N_420,In_459,In_59);
nand U421 (N_421,In_278,In_214);
nand U422 (N_422,In_34,In_227);
and U423 (N_423,In_396,In_58);
nor U424 (N_424,In_120,In_277);
or U425 (N_425,In_92,In_420);
xnor U426 (N_426,In_197,In_330);
nand U427 (N_427,In_19,In_162);
and U428 (N_428,In_331,In_371);
nand U429 (N_429,In_306,In_266);
nand U430 (N_430,In_208,In_321);
nand U431 (N_431,In_396,In_441);
and U432 (N_432,In_314,In_113);
nand U433 (N_433,In_491,In_494);
or U434 (N_434,In_183,In_303);
or U435 (N_435,In_173,In_324);
nand U436 (N_436,In_440,In_66);
nor U437 (N_437,In_75,In_46);
or U438 (N_438,In_498,In_178);
nor U439 (N_439,In_42,In_115);
nand U440 (N_440,In_227,In_165);
and U441 (N_441,In_82,In_163);
nand U442 (N_442,In_75,In_492);
and U443 (N_443,In_481,In_411);
nor U444 (N_444,In_290,In_77);
xor U445 (N_445,In_133,In_128);
nor U446 (N_446,In_88,In_133);
nor U447 (N_447,In_467,In_475);
or U448 (N_448,In_329,In_169);
and U449 (N_449,In_478,In_471);
nor U450 (N_450,In_170,In_303);
and U451 (N_451,In_57,In_54);
xor U452 (N_452,In_19,In_369);
or U453 (N_453,In_347,In_189);
nand U454 (N_454,In_186,In_223);
nor U455 (N_455,In_378,In_21);
or U456 (N_456,In_145,In_174);
or U457 (N_457,In_236,In_272);
nor U458 (N_458,In_492,In_398);
nor U459 (N_459,In_281,In_278);
nor U460 (N_460,In_260,In_240);
nor U461 (N_461,In_334,In_469);
nand U462 (N_462,In_145,In_84);
and U463 (N_463,In_293,In_328);
and U464 (N_464,In_129,In_76);
xnor U465 (N_465,In_74,In_23);
or U466 (N_466,In_44,In_498);
xor U467 (N_467,In_129,In_333);
xor U468 (N_468,In_27,In_255);
nor U469 (N_469,In_486,In_241);
and U470 (N_470,In_282,In_134);
and U471 (N_471,In_19,In_414);
nor U472 (N_472,In_12,In_258);
and U473 (N_473,In_476,In_283);
nand U474 (N_474,In_55,In_210);
nand U475 (N_475,In_247,In_110);
or U476 (N_476,In_430,In_93);
or U477 (N_477,In_316,In_30);
xor U478 (N_478,In_193,In_348);
nor U479 (N_479,In_265,In_135);
nor U480 (N_480,In_183,In_390);
or U481 (N_481,In_236,In_130);
and U482 (N_482,In_285,In_305);
xnor U483 (N_483,In_224,In_12);
and U484 (N_484,In_153,In_249);
and U485 (N_485,In_210,In_113);
and U486 (N_486,In_165,In_295);
and U487 (N_487,In_291,In_299);
or U488 (N_488,In_424,In_77);
and U489 (N_489,In_270,In_179);
xor U490 (N_490,In_11,In_259);
nor U491 (N_491,In_194,In_359);
and U492 (N_492,In_230,In_30);
nor U493 (N_493,In_128,In_213);
nand U494 (N_494,In_73,In_208);
or U495 (N_495,In_197,In_146);
nand U496 (N_496,In_405,In_462);
nand U497 (N_497,In_466,In_99);
nor U498 (N_498,In_257,In_406);
or U499 (N_499,In_301,In_389);
nor U500 (N_500,In_330,In_278);
nand U501 (N_501,In_463,In_79);
nand U502 (N_502,In_208,In_474);
or U503 (N_503,In_469,In_33);
xor U504 (N_504,In_363,In_327);
xnor U505 (N_505,In_18,In_128);
and U506 (N_506,In_229,In_95);
or U507 (N_507,In_132,In_441);
xnor U508 (N_508,In_6,In_166);
and U509 (N_509,In_391,In_354);
xnor U510 (N_510,In_316,In_396);
or U511 (N_511,In_322,In_331);
or U512 (N_512,In_351,In_175);
nand U513 (N_513,In_396,In_197);
or U514 (N_514,In_399,In_212);
xnor U515 (N_515,In_297,In_412);
and U516 (N_516,In_163,In_259);
nor U517 (N_517,In_179,In_74);
or U518 (N_518,In_162,In_249);
or U519 (N_519,In_302,In_132);
nor U520 (N_520,In_219,In_466);
xor U521 (N_521,In_23,In_153);
xnor U522 (N_522,In_335,In_192);
nor U523 (N_523,In_492,In_136);
nor U524 (N_524,In_31,In_155);
nand U525 (N_525,In_415,In_486);
or U526 (N_526,In_312,In_5);
or U527 (N_527,In_475,In_322);
and U528 (N_528,In_479,In_347);
nand U529 (N_529,In_250,In_215);
xor U530 (N_530,In_154,In_468);
nor U531 (N_531,In_185,In_401);
nor U532 (N_532,In_182,In_488);
and U533 (N_533,In_31,In_470);
xnor U534 (N_534,In_181,In_11);
and U535 (N_535,In_409,In_152);
and U536 (N_536,In_286,In_281);
xor U537 (N_537,In_271,In_91);
or U538 (N_538,In_486,In_224);
nand U539 (N_539,In_68,In_230);
or U540 (N_540,In_11,In_416);
or U541 (N_541,In_125,In_192);
or U542 (N_542,In_360,In_435);
or U543 (N_543,In_271,In_34);
nand U544 (N_544,In_324,In_74);
xor U545 (N_545,In_6,In_489);
or U546 (N_546,In_253,In_249);
and U547 (N_547,In_24,In_325);
or U548 (N_548,In_1,In_98);
nand U549 (N_549,In_30,In_412);
nand U550 (N_550,In_148,In_90);
and U551 (N_551,In_24,In_263);
nor U552 (N_552,In_71,In_377);
nor U553 (N_553,In_292,In_164);
xnor U554 (N_554,In_353,In_4);
and U555 (N_555,In_147,In_399);
xor U556 (N_556,In_278,In_402);
nor U557 (N_557,In_227,In_319);
nor U558 (N_558,In_317,In_130);
and U559 (N_559,In_466,In_387);
xnor U560 (N_560,In_134,In_131);
nor U561 (N_561,In_461,In_427);
or U562 (N_562,In_62,In_301);
nand U563 (N_563,In_11,In_383);
nor U564 (N_564,In_187,In_45);
and U565 (N_565,In_122,In_396);
and U566 (N_566,In_152,In_154);
xnor U567 (N_567,In_253,In_409);
nor U568 (N_568,In_424,In_82);
and U569 (N_569,In_466,In_474);
and U570 (N_570,In_382,In_62);
or U571 (N_571,In_189,In_427);
xor U572 (N_572,In_311,In_158);
nor U573 (N_573,In_452,In_237);
nor U574 (N_574,In_269,In_57);
nand U575 (N_575,In_454,In_206);
and U576 (N_576,In_201,In_90);
nand U577 (N_577,In_250,In_249);
nand U578 (N_578,In_404,In_49);
nand U579 (N_579,In_248,In_371);
nor U580 (N_580,In_182,In_110);
or U581 (N_581,In_238,In_231);
nor U582 (N_582,In_158,In_27);
and U583 (N_583,In_105,In_22);
and U584 (N_584,In_35,In_39);
nand U585 (N_585,In_292,In_170);
or U586 (N_586,In_217,In_143);
nand U587 (N_587,In_100,In_154);
and U588 (N_588,In_450,In_325);
xor U589 (N_589,In_333,In_132);
and U590 (N_590,In_126,In_132);
nor U591 (N_591,In_48,In_211);
nand U592 (N_592,In_467,In_362);
and U593 (N_593,In_430,In_283);
nand U594 (N_594,In_8,In_165);
or U595 (N_595,In_247,In_113);
or U596 (N_596,In_464,In_263);
nor U597 (N_597,In_188,In_63);
and U598 (N_598,In_196,In_432);
or U599 (N_599,In_56,In_237);
or U600 (N_600,N_192,N_230);
or U601 (N_601,N_475,N_105);
nand U602 (N_602,N_289,N_243);
or U603 (N_603,N_519,N_29);
or U604 (N_604,N_435,N_335);
or U605 (N_605,N_8,N_391);
and U606 (N_606,N_222,N_577);
or U607 (N_607,N_494,N_414);
or U608 (N_608,N_210,N_584);
and U609 (N_609,N_256,N_583);
and U610 (N_610,N_66,N_78);
or U611 (N_611,N_20,N_412);
nor U612 (N_612,N_261,N_509);
and U613 (N_613,N_181,N_228);
xnor U614 (N_614,N_407,N_553);
and U615 (N_615,N_572,N_88);
and U616 (N_616,N_429,N_202);
and U617 (N_617,N_346,N_428);
or U618 (N_618,N_305,N_41);
or U619 (N_619,N_340,N_334);
nand U620 (N_620,N_128,N_466);
nor U621 (N_621,N_100,N_488);
xnor U622 (N_622,N_424,N_208);
xnor U623 (N_623,N_381,N_568);
nand U624 (N_624,N_156,N_510);
and U625 (N_625,N_598,N_550);
nand U626 (N_626,N_366,N_361);
xnor U627 (N_627,N_102,N_409);
or U628 (N_628,N_533,N_106);
nor U629 (N_629,N_5,N_59);
nand U630 (N_630,N_524,N_207);
nor U631 (N_631,N_443,N_399);
or U632 (N_632,N_307,N_564);
nand U633 (N_633,N_413,N_125);
nor U634 (N_634,N_427,N_75);
nand U635 (N_635,N_184,N_2);
or U636 (N_636,N_85,N_51);
or U637 (N_637,N_436,N_549);
and U638 (N_638,N_288,N_81);
nand U639 (N_639,N_209,N_594);
nand U640 (N_640,N_4,N_582);
nor U641 (N_641,N_159,N_529);
nand U642 (N_642,N_151,N_500);
nor U643 (N_643,N_87,N_538);
xor U644 (N_644,N_219,N_499);
or U645 (N_645,N_461,N_60);
or U646 (N_646,N_291,N_512);
nor U647 (N_647,N_281,N_345);
nor U648 (N_648,N_503,N_259);
nand U649 (N_649,N_303,N_420);
xnor U650 (N_650,N_489,N_43);
nor U651 (N_651,N_279,N_23);
nand U652 (N_652,N_132,N_507);
nor U653 (N_653,N_387,N_235);
xor U654 (N_654,N_310,N_552);
nor U655 (N_655,N_229,N_473);
and U656 (N_656,N_144,N_203);
xnor U657 (N_657,N_155,N_38);
and U658 (N_658,N_445,N_395);
or U659 (N_659,N_393,N_165);
nand U660 (N_660,N_306,N_188);
nand U661 (N_661,N_397,N_343);
and U662 (N_662,N_506,N_109);
nand U663 (N_663,N_589,N_54);
and U664 (N_664,N_39,N_15);
nor U665 (N_665,N_505,N_196);
nor U666 (N_666,N_250,N_247);
and U667 (N_667,N_540,N_173);
nor U668 (N_668,N_373,N_403);
and U669 (N_669,N_421,N_548);
and U670 (N_670,N_380,N_569);
nand U671 (N_671,N_599,N_455);
nor U672 (N_672,N_73,N_292);
nand U673 (N_673,N_411,N_49);
and U674 (N_674,N_356,N_137);
nor U675 (N_675,N_103,N_270);
and U676 (N_676,N_442,N_378);
or U677 (N_677,N_40,N_493);
and U678 (N_678,N_591,N_131);
nor U679 (N_679,N_471,N_419);
and U680 (N_680,N_171,N_326);
or U681 (N_681,N_178,N_339);
nand U682 (N_682,N_468,N_145);
and U683 (N_683,N_308,N_496);
nor U684 (N_684,N_161,N_501);
nand U685 (N_685,N_3,N_14);
or U686 (N_686,N_104,N_555);
nand U687 (N_687,N_545,N_236);
nand U688 (N_688,N_439,N_86);
nand U689 (N_689,N_441,N_206);
nand U690 (N_690,N_143,N_331);
or U691 (N_691,N_425,N_267);
nand U692 (N_692,N_426,N_398);
or U693 (N_693,N_566,N_33);
nor U694 (N_694,N_392,N_543);
nand U695 (N_695,N_285,N_299);
and U696 (N_696,N_140,N_314);
or U697 (N_697,N_18,N_262);
and U698 (N_698,N_309,N_431);
and U699 (N_699,N_263,N_45);
nand U700 (N_700,N_220,N_576);
and U701 (N_701,N_296,N_417);
nor U702 (N_702,N_320,N_1);
and U703 (N_703,N_469,N_107);
nand U704 (N_704,N_370,N_482);
nor U705 (N_705,N_401,N_573);
or U706 (N_706,N_134,N_304);
and U707 (N_707,N_71,N_255);
and U708 (N_708,N_337,N_347);
and U709 (N_709,N_199,N_251);
and U710 (N_710,N_226,N_447);
nor U711 (N_711,N_28,N_79);
nor U712 (N_712,N_204,N_185);
xor U713 (N_713,N_197,N_115);
and U714 (N_714,N_430,N_191);
and U715 (N_715,N_514,N_215);
and U716 (N_716,N_234,N_32);
nand U717 (N_717,N_176,N_24);
nor U718 (N_718,N_84,N_218);
xor U719 (N_719,N_48,N_82);
or U720 (N_720,N_121,N_96);
and U721 (N_721,N_301,N_362);
nor U722 (N_722,N_574,N_205);
nand U723 (N_723,N_225,N_369);
nor U724 (N_724,N_46,N_77);
and U725 (N_725,N_183,N_186);
or U726 (N_726,N_168,N_67);
xnor U727 (N_727,N_283,N_458);
nor U728 (N_728,N_454,N_223);
nor U729 (N_729,N_195,N_198);
or U730 (N_730,N_333,N_17);
or U731 (N_731,N_123,N_354);
or U732 (N_732,N_565,N_531);
nor U733 (N_733,N_596,N_365);
nor U734 (N_734,N_271,N_98);
nand U735 (N_735,N_47,N_402);
nor U736 (N_736,N_277,N_374);
or U737 (N_737,N_313,N_90);
or U738 (N_738,N_592,N_497);
or U739 (N_739,N_316,N_537);
nand U740 (N_740,N_597,N_26);
and U741 (N_741,N_258,N_534);
xor U742 (N_742,N_53,N_358);
and U743 (N_743,N_118,N_252);
or U744 (N_744,N_302,N_245);
nor U745 (N_745,N_536,N_150);
xor U746 (N_746,N_112,N_216);
nand U747 (N_747,N_492,N_246);
nand U748 (N_748,N_450,N_55);
and U749 (N_749,N_367,N_491);
nand U750 (N_750,N_190,N_227);
and U751 (N_751,N_446,N_76);
and U752 (N_752,N_127,N_511);
or U753 (N_753,N_300,N_169);
xnor U754 (N_754,N_31,N_541);
nand U755 (N_755,N_264,N_554);
nand U756 (N_756,N_37,N_253);
nand U757 (N_757,N_16,N_116);
or U758 (N_758,N_83,N_383);
or U759 (N_759,N_244,N_50);
or U760 (N_760,N_30,N_579);
nor U761 (N_761,N_74,N_516);
or U762 (N_762,N_89,N_360);
or U763 (N_763,N_350,N_551);
or U764 (N_764,N_324,N_194);
nand U765 (N_765,N_422,N_36);
and U766 (N_766,N_415,N_286);
nor U767 (N_767,N_269,N_490);
or U768 (N_768,N_319,N_248);
or U769 (N_769,N_586,N_561);
and U770 (N_770,N_321,N_318);
nor U771 (N_771,N_290,N_472);
or U772 (N_772,N_241,N_539);
or U773 (N_773,N_348,N_390);
and U774 (N_774,N_142,N_344);
and U775 (N_775,N_578,N_135);
and U776 (N_776,N_353,N_462);
and U777 (N_777,N_182,N_265);
and U778 (N_778,N_504,N_213);
nor U779 (N_779,N_357,N_136);
xnor U780 (N_780,N_58,N_352);
and U781 (N_781,N_349,N_117);
nor U782 (N_782,N_560,N_242);
xor U783 (N_783,N_463,N_110);
and U784 (N_784,N_260,N_64);
and U785 (N_785,N_359,N_298);
xnor U786 (N_786,N_526,N_238);
or U787 (N_787,N_101,N_470);
nand U788 (N_788,N_129,N_297);
xor U789 (N_789,N_410,N_61);
xor U790 (N_790,N_523,N_379);
xor U791 (N_791,N_249,N_200);
and U792 (N_792,N_355,N_166);
or U793 (N_793,N_162,N_449);
and U794 (N_794,N_294,N_217);
and U795 (N_795,N_590,N_287);
and U796 (N_796,N_364,N_175);
nor U797 (N_797,N_10,N_556);
xnor U798 (N_798,N_92,N_465);
or U799 (N_799,N_484,N_177);
and U800 (N_800,N_276,N_495);
and U801 (N_801,N_396,N_400);
nor U802 (N_802,N_154,N_438);
nand U803 (N_803,N_328,N_476);
or U804 (N_804,N_385,N_418);
and U805 (N_805,N_240,N_485);
or U806 (N_806,N_315,N_68);
or U807 (N_807,N_487,N_167);
nand U808 (N_808,N_444,N_193);
and U809 (N_809,N_513,N_323);
nor U810 (N_810,N_515,N_464);
or U811 (N_811,N_587,N_327);
or U812 (N_812,N_133,N_224);
and U813 (N_813,N_317,N_557);
nor U814 (N_814,N_80,N_520);
xnor U815 (N_815,N_575,N_581);
or U816 (N_816,N_544,N_474);
nor U817 (N_817,N_93,N_120);
nor U818 (N_818,N_69,N_22);
or U819 (N_819,N_174,N_157);
nor U820 (N_820,N_170,N_280);
and U821 (N_821,N_44,N_152);
and U822 (N_822,N_141,N_522);
xnor U823 (N_823,N_91,N_122);
nand U824 (N_824,N_97,N_457);
or U825 (N_825,N_114,N_19);
or U826 (N_826,N_517,N_201);
nand U827 (N_827,N_570,N_70);
xnor U828 (N_828,N_214,N_486);
nor U829 (N_829,N_521,N_329);
and U830 (N_830,N_336,N_63);
nand U831 (N_831,N_139,N_332);
and U832 (N_832,N_498,N_282);
or U833 (N_833,N_322,N_558);
and U834 (N_834,N_232,N_126);
and U835 (N_835,N_404,N_372);
and U836 (N_836,N_481,N_257);
or U837 (N_837,N_593,N_371);
nand U838 (N_838,N_508,N_478);
nand U839 (N_839,N_147,N_179);
nand U840 (N_840,N_477,N_571);
nand U841 (N_841,N_35,N_562);
nor U842 (N_842,N_164,N_62);
xnor U843 (N_843,N_563,N_460);
or U844 (N_844,N_351,N_254);
nand U845 (N_845,N_416,N_342);
or U846 (N_846,N_432,N_368);
or U847 (N_847,N_448,N_275);
or U848 (N_848,N_211,N_130);
nand U849 (N_849,N_278,N_72);
and U850 (N_850,N_42,N_530);
nor U851 (N_851,N_377,N_233);
or U852 (N_852,N_113,N_108);
and U853 (N_853,N_434,N_479);
nand U854 (N_854,N_527,N_382);
nor U855 (N_855,N_146,N_325);
nor U856 (N_856,N_375,N_386);
and U857 (N_857,N_111,N_559);
nor U858 (N_858,N_212,N_595);
nand U859 (N_859,N_99,N_9);
nor U860 (N_860,N_423,N_363);
nor U861 (N_861,N_65,N_341);
nor U862 (N_862,N_388,N_172);
nand U863 (N_863,N_160,N_535);
and U864 (N_864,N_440,N_163);
nor U865 (N_865,N_119,N_7);
nand U866 (N_866,N_25,N_34);
and U867 (N_867,N_433,N_153);
nor U868 (N_868,N_57,N_542);
and U869 (N_869,N_52,N_405);
nand U870 (N_870,N_467,N_272);
nand U871 (N_871,N_0,N_237);
nor U872 (N_872,N_547,N_588);
nor U873 (N_873,N_124,N_293);
nor U874 (N_874,N_452,N_239);
xnor U875 (N_875,N_311,N_408);
nor U876 (N_876,N_546,N_187);
and U877 (N_877,N_21,N_27);
or U878 (N_878,N_180,N_437);
xor U879 (N_879,N_330,N_406);
nand U880 (N_880,N_394,N_312);
or U881 (N_881,N_273,N_480);
nor U882 (N_882,N_456,N_149);
nand U883 (N_883,N_532,N_56);
nand U884 (N_884,N_268,N_338);
nand U885 (N_885,N_221,N_451);
nor U886 (N_886,N_148,N_12);
xnor U887 (N_887,N_11,N_453);
nor U888 (N_888,N_158,N_567);
or U889 (N_889,N_376,N_525);
nand U890 (N_890,N_502,N_274);
nor U891 (N_891,N_528,N_384);
or U892 (N_892,N_189,N_13);
or U893 (N_893,N_6,N_95);
or U894 (N_894,N_138,N_580);
nand U895 (N_895,N_284,N_295);
nor U896 (N_896,N_389,N_94);
or U897 (N_897,N_585,N_483);
xor U898 (N_898,N_518,N_266);
or U899 (N_899,N_459,N_231);
nand U900 (N_900,N_391,N_472);
xnor U901 (N_901,N_490,N_28);
nand U902 (N_902,N_474,N_87);
nand U903 (N_903,N_501,N_407);
nor U904 (N_904,N_124,N_366);
nand U905 (N_905,N_352,N_34);
nor U906 (N_906,N_178,N_564);
nor U907 (N_907,N_350,N_203);
nor U908 (N_908,N_568,N_581);
nor U909 (N_909,N_242,N_90);
and U910 (N_910,N_428,N_86);
nand U911 (N_911,N_312,N_128);
nor U912 (N_912,N_311,N_88);
nor U913 (N_913,N_407,N_16);
or U914 (N_914,N_556,N_139);
and U915 (N_915,N_132,N_525);
nand U916 (N_916,N_176,N_35);
and U917 (N_917,N_571,N_214);
nor U918 (N_918,N_227,N_565);
and U919 (N_919,N_441,N_496);
or U920 (N_920,N_214,N_488);
xnor U921 (N_921,N_181,N_203);
or U922 (N_922,N_378,N_321);
or U923 (N_923,N_251,N_168);
xor U924 (N_924,N_274,N_367);
nand U925 (N_925,N_165,N_430);
nand U926 (N_926,N_53,N_317);
nand U927 (N_927,N_345,N_359);
nor U928 (N_928,N_207,N_505);
xor U929 (N_929,N_204,N_527);
and U930 (N_930,N_404,N_79);
or U931 (N_931,N_216,N_154);
or U932 (N_932,N_84,N_370);
or U933 (N_933,N_33,N_523);
and U934 (N_934,N_255,N_164);
nand U935 (N_935,N_75,N_589);
nand U936 (N_936,N_251,N_388);
nand U937 (N_937,N_499,N_279);
or U938 (N_938,N_347,N_273);
and U939 (N_939,N_429,N_102);
nor U940 (N_940,N_13,N_200);
or U941 (N_941,N_400,N_413);
and U942 (N_942,N_406,N_452);
nor U943 (N_943,N_401,N_351);
nor U944 (N_944,N_561,N_281);
and U945 (N_945,N_12,N_389);
and U946 (N_946,N_504,N_70);
xor U947 (N_947,N_117,N_250);
and U948 (N_948,N_496,N_492);
xor U949 (N_949,N_267,N_134);
nand U950 (N_950,N_417,N_360);
and U951 (N_951,N_396,N_467);
or U952 (N_952,N_246,N_429);
nor U953 (N_953,N_285,N_19);
nor U954 (N_954,N_208,N_269);
and U955 (N_955,N_521,N_583);
and U956 (N_956,N_378,N_402);
nand U957 (N_957,N_348,N_113);
nor U958 (N_958,N_63,N_345);
and U959 (N_959,N_176,N_117);
nand U960 (N_960,N_398,N_429);
and U961 (N_961,N_413,N_357);
nor U962 (N_962,N_576,N_120);
or U963 (N_963,N_457,N_397);
and U964 (N_964,N_414,N_148);
nand U965 (N_965,N_329,N_424);
nand U966 (N_966,N_241,N_227);
nor U967 (N_967,N_193,N_308);
or U968 (N_968,N_442,N_427);
nor U969 (N_969,N_290,N_226);
and U970 (N_970,N_479,N_369);
nand U971 (N_971,N_453,N_266);
nand U972 (N_972,N_116,N_337);
nand U973 (N_973,N_599,N_365);
and U974 (N_974,N_39,N_422);
nor U975 (N_975,N_145,N_11);
or U976 (N_976,N_414,N_320);
xnor U977 (N_977,N_411,N_555);
nor U978 (N_978,N_403,N_515);
and U979 (N_979,N_56,N_572);
and U980 (N_980,N_5,N_223);
or U981 (N_981,N_122,N_593);
nand U982 (N_982,N_119,N_301);
and U983 (N_983,N_226,N_504);
and U984 (N_984,N_573,N_79);
or U985 (N_985,N_372,N_122);
nand U986 (N_986,N_273,N_41);
nand U987 (N_987,N_453,N_295);
and U988 (N_988,N_103,N_550);
and U989 (N_989,N_238,N_301);
nand U990 (N_990,N_364,N_386);
xnor U991 (N_991,N_430,N_271);
nor U992 (N_992,N_361,N_428);
or U993 (N_993,N_273,N_269);
and U994 (N_994,N_547,N_442);
nor U995 (N_995,N_480,N_410);
nand U996 (N_996,N_217,N_513);
nor U997 (N_997,N_384,N_518);
nand U998 (N_998,N_357,N_450);
nand U999 (N_999,N_511,N_390);
nor U1000 (N_1000,N_344,N_363);
or U1001 (N_1001,N_285,N_78);
or U1002 (N_1002,N_496,N_1);
nand U1003 (N_1003,N_491,N_380);
nor U1004 (N_1004,N_115,N_87);
and U1005 (N_1005,N_231,N_398);
nand U1006 (N_1006,N_521,N_513);
nand U1007 (N_1007,N_175,N_595);
and U1008 (N_1008,N_313,N_260);
nand U1009 (N_1009,N_224,N_65);
nor U1010 (N_1010,N_543,N_56);
xnor U1011 (N_1011,N_246,N_150);
nand U1012 (N_1012,N_349,N_543);
and U1013 (N_1013,N_406,N_160);
nand U1014 (N_1014,N_487,N_344);
or U1015 (N_1015,N_11,N_529);
nor U1016 (N_1016,N_543,N_156);
or U1017 (N_1017,N_513,N_232);
nand U1018 (N_1018,N_416,N_456);
xnor U1019 (N_1019,N_80,N_382);
and U1020 (N_1020,N_128,N_213);
nand U1021 (N_1021,N_47,N_356);
nor U1022 (N_1022,N_440,N_414);
or U1023 (N_1023,N_413,N_17);
nand U1024 (N_1024,N_450,N_558);
or U1025 (N_1025,N_371,N_78);
or U1026 (N_1026,N_469,N_419);
nor U1027 (N_1027,N_281,N_167);
nand U1028 (N_1028,N_123,N_510);
nor U1029 (N_1029,N_185,N_470);
or U1030 (N_1030,N_253,N_94);
or U1031 (N_1031,N_538,N_382);
and U1032 (N_1032,N_64,N_250);
xnor U1033 (N_1033,N_1,N_575);
xnor U1034 (N_1034,N_222,N_483);
nand U1035 (N_1035,N_18,N_514);
nor U1036 (N_1036,N_308,N_124);
nor U1037 (N_1037,N_532,N_407);
or U1038 (N_1038,N_37,N_285);
xor U1039 (N_1039,N_330,N_182);
nor U1040 (N_1040,N_343,N_103);
nand U1041 (N_1041,N_380,N_499);
and U1042 (N_1042,N_305,N_160);
and U1043 (N_1043,N_457,N_442);
nor U1044 (N_1044,N_228,N_299);
nor U1045 (N_1045,N_153,N_311);
and U1046 (N_1046,N_245,N_455);
or U1047 (N_1047,N_230,N_398);
or U1048 (N_1048,N_28,N_238);
nor U1049 (N_1049,N_39,N_115);
nor U1050 (N_1050,N_585,N_425);
and U1051 (N_1051,N_24,N_471);
nand U1052 (N_1052,N_488,N_306);
or U1053 (N_1053,N_82,N_372);
nor U1054 (N_1054,N_463,N_54);
xor U1055 (N_1055,N_380,N_197);
or U1056 (N_1056,N_536,N_489);
or U1057 (N_1057,N_272,N_296);
or U1058 (N_1058,N_88,N_581);
and U1059 (N_1059,N_81,N_64);
or U1060 (N_1060,N_180,N_572);
and U1061 (N_1061,N_248,N_365);
or U1062 (N_1062,N_18,N_273);
or U1063 (N_1063,N_593,N_104);
nand U1064 (N_1064,N_576,N_17);
nand U1065 (N_1065,N_78,N_501);
nor U1066 (N_1066,N_16,N_98);
or U1067 (N_1067,N_220,N_393);
and U1068 (N_1068,N_182,N_212);
nand U1069 (N_1069,N_46,N_491);
or U1070 (N_1070,N_221,N_156);
or U1071 (N_1071,N_479,N_169);
xor U1072 (N_1072,N_493,N_491);
and U1073 (N_1073,N_72,N_446);
xnor U1074 (N_1074,N_383,N_266);
and U1075 (N_1075,N_396,N_137);
nor U1076 (N_1076,N_525,N_515);
and U1077 (N_1077,N_255,N_366);
or U1078 (N_1078,N_161,N_482);
or U1079 (N_1079,N_215,N_122);
and U1080 (N_1080,N_479,N_301);
nor U1081 (N_1081,N_492,N_125);
nor U1082 (N_1082,N_245,N_483);
nor U1083 (N_1083,N_324,N_158);
xnor U1084 (N_1084,N_283,N_285);
nor U1085 (N_1085,N_180,N_198);
nor U1086 (N_1086,N_131,N_344);
and U1087 (N_1087,N_63,N_312);
nor U1088 (N_1088,N_63,N_203);
nand U1089 (N_1089,N_147,N_576);
nor U1090 (N_1090,N_522,N_382);
nand U1091 (N_1091,N_201,N_290);
nor U1092 (N_1092,N_367,N_577);
and U1093 (N_1093,N_579,N_0);
and U1094 (N_1094,N_212,N_384);
nor U1095 (N_1095,N_139,N_230);
and U1096 (N_1096,N_212,N_308);
and U1097 (N_1097,N_494,N_287);
xnor U1098 (N_1098,N_82,N_40);
nor U1099 (N_1099,N_1,N_74);
nand U1100 (N_1100,N_246,N_526);
nor U1101 (N_1101,N_529,N_495);
or U1102 (N_1102,N_275,N_2);
nor U1103 (N_1103,N_208,N_301);
xor U1104 (N_1104,N_225,N_218);
nand U1105 (N_1105,N_533,N_494);
nor U1106 (N_1106,N_463,N_547);
nor U1107 (N_1107,N_312,N_534);
nand U1108 (N_1108,N_525,N_226);
and U1109 (N_1109,N_496,N_364);
nand U1110 (N_1110,N_250,N_55);
nor U1111 (N_1111,N_39,N_367);
and U1112 (N_1112,N_117,N_576);
and U1113 (N_1113,N_591,N_51);
nor U1114 (N_1114,N_328,N_474);
and U1115 (N_1115,N_109,N_269);
or U1116 (N_1116,N_166,N_80);
and U1117 (N_1117,N_399,N_164);
xor U1118 (N_1118,N_586,N_19);
nand U1119 (N_1119,N_257,N_352);
xnor U1120 (N_1120,N_91,N_390);
nand U1121 (N_1121,N_517,N_294);
nand U1122 (N_1122,N_343,N_207);
nor U1123 (N_1123,N_340,N_186);
nand U1124 (N_1124,N_275,N_195);
and U1125 (N_1125,N_126,N_230);
or U1126 (N_1126,N_193,N_79);
and U1127 (N_1127,N_367,N_570);
or U1128 (N_1128,N_178,N_64);
nand U1129 (N_1129,N_225,N_211);
xor U1130 (N_1130,N_428,N_476);
nand U1131 (N_1131,N_66,N_358);
nor U1132 (N_1132,N_402,N_146);
nand U1133 (N_1133,N_266,N_125);
xor U1134 (N_1134,N_385,N_577);
nand U1135 (N_1135,N_417,N_41);
and U1136 (N_1136,N_532,N_198);
and U1137 (N_1137,N_596,N_215);
or U1138 (N_1138,N_47,N_37);
and U1139 (N_1139,N_419,N_71);
nor U1140 (N_1140,N_241,N_122);
or U1141 (N_1141,N_239,N_292);
or U1142 (N_1142,N_392,N_307);
xnor U1143 (N_1143,N_402,N_553);
and U1144 (N_1144,N_242,N_357);
and U1145 (N_1145,N_581,N_240);
nand U1146 (N_1146,N_500,N_588);
and U1147 (N_1147,N_204,N_108);
nand U1148 (N_1148,N_208,N_24);
or U1149 (N_1149,N_93,N_193);
nand U1150 (N_1150,N_591,N_24);
or U1151 (N_1151,N_458,N_499);
nand U1152 (N_1152,N_410,N_9);
nor U1153 (N_1153,N_553,N_81);
and U1154 (N_1154,N_464,N_500);
xor U1155 (N_1155,N_485,N_74);
nand U1156 (N_1156,N_118,N_68);
or U1157 (N_1157,N_405,N_360);
xor U1158 (N_1158,N_529,N_595);
nor U1159 (N_1159,N_440,N_43);
nor U1160 (N_1160,N_10,N_3);
and U1161 (N_1161,N_401,N_285);
or U1162 (N_1162,N_234,N_592);
nand U1163 (N_1163,N_400,N_255);
or U1164 (N_1164,N_451,N_390);
or U1165 (N_1165,N_167,N_574);
xor U1166 (N_1166,N_7,N_219);
nor U1167 (N_1167,N_386,N_275);
and U1168 (N_1168,N_382,N_457);
xor U1169 (N_1169,N_56,N_429);
nor U1170 (N_1170,N_81,N_88);
or U1171 (N_1171,N_272,N_41);
and U1172 (N_1172,N_174,N_343);
nand U1173 (N_1173,N_463,N_369);
and U1174 (N_1174,N_563,N_439);
and U1175 (N_1175,N_444,N_212);
or U1176 (N_1176,N_266,N_163);
and U1177 (N_1177,N_28,N_37);
nor U1178 (N_1178,N_102,N_354);
and U1179 (N_1179,N_376,N_486);
nor U1180 (N_1180,N_296,N_447);
and U1181 (N_1181,N_30,N_450);
nand U1182 (N_1182,N_313,N_41);
and U1183 (N_1183,N_47,N_411);
nor U1184 (N_1184,N_237,N_34);
and U1185 (N_1185,N_460,N_5);
nor U1186 (N_1186,N_183,N_493);
nand U1187 (N_1187,N_126,N_479);
xor U1188 (N_1188,N_283,N_539);
xor U1189 (N_1189,N_201,N_174);
nand U1190 (N_1190,N_371,N_151);
or U1191 (N_1191,N_105,N_321);
and U1192 (N_1192,N_282,N_186);
and U1193 (N_1193,N_216,N_100);
and U1194 (N_1194,N_550,N_186);
or U1195 (N_1195,N_278,N_110);
or U1196 (N_1196,N_241,N_130);
nand U1197 (N_1197,N_111,N_549);
or U1198 (N_1198,N_237,N_303);
and U1199 (N_1199,N_94,N_372);
and U1200 (N_1200,N_843,N_1175);
xnor U1201 (N_1201,N_1079,N_758);
and U1202 (N_1202,N_816,N_1125);
nand U1203 (N_1203,N_1152,N_888);
and U1204 (N_1204,N_842,N_777);
nand U1205 (N_1205,N_1133,N_992);
or U1206 (N_1206,N_608,N_637);
nor U1207 (N_1207,N_771,N_780);
nand U1208 (N_1208,N_1195,N_1070);
nor U1209 (N_1209,N_689,N_1106);
or U1210 (N_1210,N_657,N_703);
or U1211 (N_1211,N_721,N_905);
nand U1212 (N_1212,N_870,N_912);
or U1213 (N_1213,N_834,N_977);
and U1214 (N_1214,N_656,N_1198);
or U1215 (N_1215,N_801,N_981);
nor U1216 (N_1216,N_1132,N_1167);
and U1217 (N_1217,N_916,N_720);
nor U1218 (N_1218,N_1166,N_601);
nand U1219 (N_1219,N_983,N_1112);
nor U1220 (N_1220,N_996,N_701);
and U1221 (N_1221,N_640,N_845);
or U1222 (N_1222,N_957,N_614);
and U1223 (N_1223,N_1055,N_726);
and U1224 (N_1224,N_1134,N_787);
and U1225 (N_1225,N_1072,N_891);
or U1226 (N_1226,N_663,N_1016);
xor U1227 (N_1227,N_974,N_802);
nor U1228 (N_1228,N_664,N_984);
nor U1229 (N_1229,N_788,N_894);
nor U1230 (N_1230,N_826,N_806);
nand U1231 (N_1231,N_918,N_1184);
or U1232 (N_1232,N_669,N_739);
and U1233 (N_1233,N_1093,N_970);
nor U1234 (N_1234,N_849,N_619);
nor U1235 (N_1235,N_1199,N_1110);
or U1236 (N_1236,N_618,N_817);
and U1237 (N_1237,N_973,N_959);
nor U1238 (N_1238,N_877,N_1138);
and U1239 (N_1239,N_807,N_1127);
and U1240 (N_1240,N_1096,N_958);
or U1241 (N_1241,N_860,N_790);
or U1242 (N_1242,N_913,N_990);
and U1243 (N_1243,N_661,N_910);
nor U1244 (N_1244,N_688,N_994);
nand U1245 (N_1245,N_662,N_792);
nand U1246 (N_1246,N_706,N_915);
nand U1247 (N_1247,N_925,N_815);
nor U1248 (N_1248,N_940,N_965);
nor U1249 (N_1249,N_715,N_1118);
nand U1250 (N_1250,N_677,N_969);
and U1251 (N_1251,N_799,N_1062);
nor U1252 (N_1252,N_833,N_865);
nor U1253 (N_1253,N_735,N_961);
nor U1254 (N_1254,N_773,N_675);
and U1255 (N_1255,N_779,N_737);
nand U1256 (N_1256,N_1089,N_821);
or U1257 (N_1257,N_639,N_606);
xor U1258 (N_1258,N_921,N_653);
nand U1259 (N_1259,N_650,N_613);
or U1260 (N_1260,N_927,N_723);
or U1261 (N_1261,N_649,N_698);
and U1262 (N_1262,N_1058,N_1029);
nand U1263 (N_1263,N_630,N_682);
nand U1264 (N_1264,N_690,N_1050);
nor U1265 (N_1265,N_896,N_869);
and U1266 (N_1266,N_738,N_1101);
or U1267 (N_1267,N_725,N_1042);
nand U1268 (N_1268,N_1009,N_1066);
nor U1269 (N_1269,N_864,N_926);
or U1270 (N_1270,N_979,N_665);
or U1271 (N_1271,N_1174,N_644);
nor U1272 (N_1272,N_1035,N_818);
nor U1273 (N_1273,N_786,N_862);
or U1274 (N_1274,N_765,N_700);
nand U1275 (N_1275,N_1038,N_828);
or U1276 (N_1276,N_634,N_945);
nor U1277 (N_1277,N_829,N_646);
nand U1278 (N_1278,N_1154,N_658);
or U1279 (N_1279,N_1027,N_968);
xnor U1280 (N_1280,N_1103,N_673);
xnor U1281 (N_1281,N_1164,N_617);
and U1282 (N_1282,N_1182,N_895);
and U1283 (N_1283,N_1054,N_1030);
and U1284 (N_1284,N_1105,N_728);
nand U1285 (N_1285,N_672,N_1092);
xnor U1286 (N_1286,N_797,N_827);
or U1287 (N_1287,N_727,N_670);
nand U1288 (N_1288,N_1005,N_881);
nand U1289 (N_1289,N_1071,N_948);
nand U1290 (N_1290,N_620,N_1080);
or U1291 (N_1291,N_930,N_755);
nor U1292 (N_1292,N_1033,N_1019);
or U1293 (N_1293,N_1081,N_732);
nand U1294 (N_1294,N_678,N_1015);
nor U1295 (N_1295,N_874,N_1017);
xnor U1296 (N_1296,N_1187,N_1056);
or U1297 (N_1297,N_887,N_847);
nand U1298 (N_1298,N_1122,N_627);
xnor U1299 (N_1299,N_840,N_1143);
and U1300 (N_1300,N_1116,N_685);
and U1301 (N_1301,N_729,N_1082);
nand U1302 (N_1302,N_605,N_623);
nand U1303 (N_1303,N_609,N_772);
and U1304 (N_1304,N_1156,N_784);
nor U1305 (N_1305,N_1045,N_964);
and U1306 (N_1306,N_1057,N_1064);
xor U1307 (N_1307,N_615,N_907);
xor U1308 (N_1308,N_1048,N_804);
nor U1309 (N_1309,N_805,N_632);
and U1310 (N_1310,N_830,N_1136);
or U1311 (N_1311,N_1173,N_971);
nand U1312 (N_1312,N_922,N_1194);
nor U1313 (N_1313,N_743,N_1069);
nor U1314 (N_1314,N_759,N_949);
nor U1315 (N_1315,N_1075,N_684);
nor U1316 (N_1316,N_696,N_796);
nand U1317 (N_1317,N_704,N_782);
nand U1318 (N_1318,N_975,N_951);
and U1319 (N_1319,N_1128,N_836);
nand U1320 (N_1320,N_871,N_686);
and U1321 (N_1321,N_1098,N_624);
nand U1322 (N_1322,N_1003,N_1145);
and U1323 (N_1323,N_603,N_1140);
nor U1324 (N_1324,N_791,N_960);
nand U1325 (N_1325,N_1063,N_1094);
and U1326 (N_1326,N_838,N_941);
nor U1327 (N_1327,N_929,N_846);
nand U1328 (N_1328,N_939,N_955);
and U1329 (N_1329,N_1013,N_919);
and U1330 (N_1330,N_1160,N_946);
nand U1331 (N_1331,N_884,N_1171);
nor U1332 (N_1332,N_962,N_789);
or U1333 (N_1333,N_1020,N_1067);
xnor U1334 (N_1334,N_1120,N_943);
and U1335 (N_1335,N_1124,N_745);
and U1336 (N_1336,N_1170,N_1104);
nor U1337 (N_1337,N_988,N_825);
nor U1338 (N_1338,N_1165,N_1126);
and U1339 (N_1339,N_694,N_692);
xnor U1340 (N_1340,N_610,N_803);
xnor U1341 (N_1341,N_1002,N_991);
and U1342 (N_1342,N_898,N_1014);
or U1343 (N_1343,N_1012,N_892);
nand U1344 (N_1344,N_1037,N_1185);
nor U1345 (N_1345,N_902,N_1053);
nor U1346 (N_1346,N_638,N_1011);
xor U1347 (N_1347,N_911,N_1022);
or U1348 (N_1348,N_1032,N_848);
and U1349 (N_1349,N_748,N_736);
xor U1350 (N_1350,N_839,N_600);
or U1351 (N_1351,N_1169,N_611);
and U1352 (N_1352,N_1028,N_1065);
or U1353 (N_1353,N_820,N_1059);
and U1354 (N_1354,N_747,N_966);
or U1355 (N_1355,N_641,N_770);
or U1356 (N_1356,N_722,N_989);
nor U1357 (N_1357,N_942,N_1180);
nand U1358 (N_1358,N_856,N_740);
xor U1359 (N_1359,N_742,N_1197);
and U1360 (N_1360,N_1129,N_795);
and U1361 (N_1361,N_1010,N_1047);
nor U1362 (N_1362,N_1097,N_668);
nor U1363 (N_1363,N_724,N_1087);
nor U1364 (N_1364,N_1151,N_831);
nor U1365 (N_1365,N_985,N_950);
nand U1366 (N_1366,N_1091,N_978);
or U1367 (N_1367,N_982,N_794);
nor U1368 (N_1368,N_659,N_835);
nand U1369 (N_1369,N_642,N_1141);
nand U1370 (N_1370,N_652,N_878);
nand U1371 (N_1371,N_844,N_1114);
nor U1372 (N_1372,N_868,N_1025);
xor U1373 (N_1373,N_1043,N_1131);
and U1374 (N_1374,N_967,N_876);
nand U1375 (N_1375,N_1108,N_900);
and U1376 (N_1376,N_1026,N_655);
and U1377 (N_1377,N_622,N_1039);
and U1378 (N_1378,N_811,N_651);
and U1379 (N_1379,N_1153,N_762);
nor U1380 (N_1380,N_853,N_956);
and U1381 (N_1381,N_1041,N_1007);
or U1382 (N_1382,N_674,N_1188);
or U1383 (N_1383,N_1192,N_824);
and U1384 (N_1384,N_712,N_719);
and U1385 (N_1385,N_875,N_1190);
or U1386 (N_1386,N_708,N_920);
or U1387 (N_1387,N_1163,N_886);
and U1388 (N_1388,N_681,N_934);
nand U1389 (N_1389,N_947,N_1158);
nand U1390 (N_1390,N_1196,N_936);
or U1391 (N_1391,N_626,N_768);
and U1392 (N_1392,N_1000,N_1083);
nor U1393 (N_1393,N_1102,N_889);
and U1394 (N_1394,N_707,N_1168);
nor U1395 (N_1395,N_1001,N_775);
nand U1396 (N_1396,N_963,N_778);
and U1397 (N_1397,N_935,N_1161);
and U1398 (N_1398,N_858,N_903);
nor U1399 (N_1399,N_1130,N_635);
and U1400 (N_1400,N_810,N_751);
xor U1401 (N_1401,N_883,N_1018);
nand U1402 (N_1402,N_976,N_1149);
or U1403 (N_1403,N_953,N_1176);
and U1404 (N_1404,N_1077,N_741);
or U1405 (N_1405,N_914,N_998);
and U1406 (N_1406,N_800,N_1024);
nor U1407 (N_1407,N_631,N_937);
and U1408 (N_1408,N_753,N_699);
or U1409 (N_1409,N_1086,N_1078);
and U1410 (N_1410,N_628,N_1052);
and U1411 (N_1411,N_890,N_863);
or U1412 (N_1412,N_814,N_711);
or U1413 (N_1413,N_1181,N_1178);
nand U1414 (N_1414,N_687,N_660);
nand U1415 (N_1415,N_1060,N_944);
or U1416 (N_1416,N_746,N_904);
nand U1417 (N_1417,N_972,N_813);
and U1418 (N_1418,N_604,N_679);
nand U1419 (N_1419,N_852,N_676);
nor U1420 (N_1420,N_1109,N_633);
and U1421 (N_1421,N_693,N_757);
nand U1422 (N_1422,N_808,N_931);
and U1423 (N_1423,N_785,N_861);
nor U1424 (N_1424,N_1090,N_809);
xor U1425 (N_1425,N_1147,N_1183);
and U1426 (N_1426,N_885,N_938);
nand U1427 (N_1427,N_1044,N_909);
nor U1428 (N_1428,N_1135,N_1121);
and U1429 (N_1429,N_752,N_616);
and U1430 (N_1430,N_798,N_1117);
nand U1431 (N_1431,N_893,N_749);
and U1432 (N_1432,N_781,N_1021);
or U1433 (N_1433,N_1004,N_837);
nor U1434 (N_1434,N_756,N_841);
nor U1435 (N_1435,N_851,N_691);
or U1436 (N_1436,N_1076,N_629);
and U1437 (N_1437,N_764,N_1088);
or U1438 (N_1438,N_1068,N_709);
nor U1439 (N_1439,N_1074,N_645);
nand U1440 (N_1440,N_647,N_999);
and U1441 (N_1441,N_1095,N_854);
and U1442 (N_1442,N_1100,N_714);
or U1443 (N_1443,N_901,N_1150);
or U1444 (N_1444,N_710,N_1084);
nand U1445 (N_1445,N_1157,N_812);
nor U1446 (N_1446,N_1023,N_872);
nor U1447 (N_1447,N_1115,N_731);
nand U1448 (N_1448,N_1179,N_713);
nand U1449 (N_1449,N_643,N_734);
xor U1450 (N_1450,N_702,N_625);
or U1451 (N_1451,N_1172,N_1036);
nor U1452 (N_1452,N_897,N_857);
nand U1453 (N_1453,N_987,N_1099);
nand U1454 (N_1454,N_733,N_1006);
and U1455 (N_1455,N_680,N_832);
nor U1456 (N_1456,N_683,N_744);
nand U1457 (N_1457,N_1159,N_997);
or U1458 (N_1458,N_774,N_932);
nand U1459 (N_1459,N_636,N_760);
nand U1460 (N_1460,N_750,N_859);
xnor U1461 (N_1461,N_899,N_882);
and U1462 (N_1462,N_697,N_666);
nand U1463 (N_1463,N_1061,N_1191);
nor U1464 (N_1464,N_1142,N_822);
and U1465 (N_1465,N_880,N_1034);
xor U1466 (N_1466,N_823,N_761);
nand U1467 (N_1467,N_924,N_783);
or U1468 (N_1468,N_952,N_1113);
nor U1469 (N_1469,N_1144,N_1193);
nand U1470 (N_1470,N_705,N_1049);
nand U1471 (N_1471,N_763,N_879);
nor U1472 (N_1472,N_1123,N_866);
and U1473 (N_1473,N_1155,N_980);
nand U1474 (N_1474,N_1177,N_1040);
and U1475 (N_1475,N_1111,N_1046);
nand U1476 (N_1476,N_716,N_917);
or U1477 (N_1477,N_1146,N_867);
and U1478 (N_1478,N_621,N_928);
and U1479 (N_1479,N_954,N_1031);
and U1480 (N_1480,N_717,N_1051);
nand U1481 (N_1481,N_995,N_819);
xnor U1482 (N_1482,N_612,N_1186);
nor U1483 (N_1483,N_923,N_776);
nand U1484 (N_1484,N_1139,N_754);
nor U1485 (N_1485,N_986,N_769);
xor U1486 (N_1486,N_767,N_873);
or U1487 (N_1487,N_718,N_906);
xor U1488 (N_1488,N_648,N_695);
nand U1489 (N_1489,N_933,N_1137);
or U1490 (N_1490,N_1085,N_654);
or U1491 (N_1491,N_908,N_793);
nor U1492 (N_1492,N_1119,N_671);
nor U1493 (N_1493,N_607,N_602);
nor U1494 (N_1494,N_1162,N_1107);
nand U1495 (N_1495,N_1073,N_850);
and U1496 (N_1496,N_1148,N_993);
nor U1497 (N_1497,N_667,N_730);
nor U1498 (N_1498,N_855,N_766);
xnor U1499 (N_1499,N_1008,N_1189);
nand U1500 (N_1500,N_1048,N_717);
nor U1501 (N_1501,N_1096,N_1077);
nand U1502 (N_1502,N_1152,N_715);
xor U1503 (N_1503,N_884,N_1131);
and U1504 (N_1504,N_745,N_958);
nor U1505 (N_1505,N_633,N_634);
nor U1506 (N_1506,N_964,N_609);
nor U1507 (N_1507,N_608,N_803);
xor U1508 (N_1508,N_816,N_1170);
nand U1509 (N_1509,N_994,N_979);
and U1510 (N_1510,N_1077,N_710);
and U1511 (N_1511,N_1129,N_1031);
nor U1512 (N_1512,N_899,N_1147);
nor U1513 (N_1513,N_833,N_1090);
nand U1514 (N_1514,N_1043,N_1133);
and U1515 (N_1515,N_603,N_772);
nor U1516 (N_1516,N_1137,N_1048);
or U1517 (N_1517,N_859,N_1071);
nand U1518 (N_1518,N_809,N_1033);
or U1519 (N_1519,N_688,N_945);
nor U1520 (N_1520,N_647,N_1108);
and U1521 (N_1521,N_955,N_889);
nand U1522 (N_1522,N_890,N_1095);
xor U1523 (N_1523,N_992,N_917);
nand U1524 (N_1524,N_1048,N_1169);
or U1525 (N_1525,N_756,N_875);
nand U1526 (N_1526,N_695,N_977);
xnor U1527 (N_1527,N_1014,N_962);
nand U1528 (N_1528,N_1090,N_669);
nand U1529 (N_1529,N_1069,N_627);
and U1530 (N_1530,N_806,N_641);
or U1531 (N_1531,N_728,N_1085);
and U1532 (N_1532,N_1160,N_704);
xnor U1533 (N_1533,N_976,N_1044);
nand U1534 (N_1534,N_1016,N_749);
nor U1535 (N_1535,N_844,N_986);
nand U1536 (N_1536,N_1096,N_1048);
nand U1537 (N_1537,N_865,N_1061);
and U1538 (N_1538,N_1078,N_751);
nand U1539 (N_1539,N_1025,N_1030);
nor U1540 (N_1540,N_623,N_1010);
and U1541 (N_1541,N_973,N_775);
nand U1542 (N_1542,N_1154,N_749);
or U1543 (N_1543,N_655,N_661);
nor U1544 (N_1544,N_626,N_903);
or U1545 (N_1545,N_887,N_1000);
nand U1546 (N_1546,N_670,N_716);
xnor U1547 (N_1547,N_815,N_756);
or U1548 (N_1548,N_870,N_1198);
and U1549 (N_1549,N_1038,N_987);
xor U1550 (N_1550,N_1092,N_728);
nand U1551 (N_1551,N_757,N_711);
nand U1552 (N_1552,N_730,N_1087);
and U1553 (N_1553,N_721,N_1197);
or U1554 (N_1554,N_757,N_784);
or U1555 (N_1555,N_717,N_691);
or U1556 (N_1556,N_1138,N_646);
xnor U1557 (N_1557,N_639,N_673);
nor U1558 (N_1558,N_985,N_933);
nor U1559 (N_1559,N_911,N_1052);
nor U1560 (N_1560,N_1008,N_729);
nand U1561 (N_1561,N_611,N_1146);
nand U1562 (N_1562,N_914,N_830);
and U1563 (N_1563,N_790,N_1168);
xor U1564 (N_1564,N_1073,N_854);
or U1565 (N_1565,N_621,N_828);
xor U1566 (N_1566,N_1172,N_656);
nand U1567 (N_1567,N_1052,N_1126);
or U1568 (N_1568,N_1122,N_1070);
nor U1569 (N_1569,N_753,N_689);
nand U1570 (N_1570,N_820,N_972);
and U1571 (N_1571,N_1013,N_721);
nor U1572 (N_1572,N_1025,N_761);
or U1573 (N_1573,N_796,N_1086);
or U1574 (N_1574,N_1112,N_652);
and U1575 (N_1575,N_656,N_768);
nand U1576 (N_1576,N_992,N_714);
or U1577 (N_1577,N_872,N_914);
or U1578 (N_1578,N_1046,N_628);
and U1579 (N_1579,N_736,N_1082);
and U1580 (N_1580,N_703,N_890);
and U1581 (N_1581,N_1057,N_674);
and U1582 (N_1582,N_870,N_886);
and U1583 (N_1583,N_702,N_1018);
and U1584 (N_1584,N_1103,N_988);
nor U1585 (N_1585,N_1080,N_748);
and U1586 (N_1586,N_736,N_893);
nand U1587 (N_1587,N_945,N_807);
nor U1588 (N_1588,N_656,N_1108);
nor U1589 (N_1589,N_789,N_758);
nor U1590 (N_1590,N_994,N_931);
nor U1591 (N_1591,N_1080,N_670);
nor U1592 (N_1592,N_830,N_1047);
nor U1593 (N_1593,N_1141,N_961);
nor U1594 (N_1594,N_652,N_768);
nand U1595 (N_1595,N_921,N_1146);
and U1596 (N_1596,N_1037,N_995);
or U1597 (N_1597,N_641,N_632);
xnor U1598 (N_1598,N_873,N_775);
or U1599 (N_1599,N_1131,N_971);
or U1600 (N_1600,N_659,N_977);
nand U1601 (N_1601,N_1169,N_1114);
nor U1602 (N_1602,N_1011,N_605);
or U1603 (N_1603,N_1008,N_1113);
nor U1604 (N_1604,N_883,N_614);
nor U1605 (N_1605,N_877,N_956);
nand U1606 (N_1606,N_1195,N_703);
xnor U1607 (N_1607,N_693,N_855);
nor U1608 (N_1608,N_1138,N_1108);
nor U1609 (N_1609,N_808,N_954);
or U1610 (N_1610,N_940,N_755);
nand U1611 (N_1611,N_600,N_1114);
and U1612 (N_1612,N_650,N_1174);
xor U1613 (N_1613,N_1138,N_911);
xor U1614 (N_1614,N_1145,N_1070);
nor U1615 (N_1615,N_692,N_722);
and U1616 (N_1616,N_800,N_641);
nand U1617 (N_1617,N_735,N_1081);
nand U1618 (N_1618,N_989,N_964);
xor U1619 (N_1619,N_640,N_1153);
nor U1620 (N_1620,N_1070,N_876);
nor U1621 (N_1621,N_1150,N_1079);
xnor U1622 (N_1622,N_960,N_913);
or U1623 (N_1623,N_779,N_602);
nor U1624 (N_1624,N_621,N_891);
xnor U1625 (N_1625,N_710,N_737);
and U1626 (N_1626,N_779,N_632);
or U1627 (N_1627,N_1178,N_769);
or U1628 (N_1628,N_648,N_980);
nand U1629 (N_1629,N_1093,N_690);
or U1630 (N_1630,N_827,N_1072);
or U1631 (N_1631,N_807,N_1142);
nor U1632 (N_1632,N_1141,N_1167);
or U1633 (N_1633,N_1152,N_892);
xor U1634 (N_1634,N_1064,N_937);
or U1635 (N_1635,N_764,N_1168);
and U1636 (N_1636,N_952,N_615);
nor U1637 (N_1637,N_1004,N_728);
xnor U1638 (N_1638,N_833,N_1012);
nand U1639 (N_1639,N_999,N_733);
or U1640 (N_1640,N_833,N_853);
nand U1641 (N_1641,N_1043,N_1115);
nand U1642 (N_1642,N_796,N_1187);
and U1643 (N_1643,N_648,N_757);
nand U1644 (N_1644,N_709,N_1146);
or U1645 (N_1645,N_993,N_731);
xor U1646 (N_1646,N_1161,N_875);
nand U1647 (N_1647,N_611,N_883);
nor U1648 (N_1648,N_756,N_739);
nand U1649 (N_1649,N_760,N_728);
or U1650 (N_1650,N_699,N_1003);
nor U1651 (N_1651,N_1059,N_1030);
and U1652 (N_1652,N_914,N_700);
xnor U1653 (N_1653,N_981,N_1025);
and U1654 (N_1654,N_731,N_629);
nand U1655 (N_1655,N_953,N_640);
xnor U1656 (N_1656,N_651,N_667);
and U1657 (N_1657,N_677,N_1155);
nor U1658 (N_1658,N_925,N_754);
nand U1659 (N_1659,N_825,N_605);
nand U1660 (N_1660,N_1119,N_1028);
nor U1661 (N_1661,N_1130,N_1139);
nand U1662 (N_1662,N_717,N_1155);
nor U1663 (N_1663,N_1137,N_622);
or U1664 (N_1664,N_982,N_1036);
or U1665 (N_1665,N_816,N_796);
xnor U1666 (N_1666,N_610,N_1146);
xnor U1667 (N_1667,N_991,N_638);
nand U1668 (N_1668,N_1192,N_902);
nand U1669 (N_1669,N_1164,N_937);
nor U1670 (N_1670,N_1178,N_637);
and U1671 (N_1671,N_825,N_726);
nor U1672 (N_1672,N_641,N_1041);
nand U1673 (N_1673,N_1131,N_1098);
or U1674 (N_1674,N_757,N_1159);
or U1675 (N_1675,N_722,N_923);
and U1676 (N_1676,N_985,N_921);
nor U1677 (N_1677,N_1125,N_846);
nor U1678 (N_1678,N_1033,N_816);
or U1679 (N_1679,N_1118,N_1114);
or U1680 (N_1680,N_697,N_878);
and U1681 (N_1681,N_980,N_635);
or U1682 (N_1682,N_1057,N_800);
nand U1683 (N_1683,N_972,N_1113);
nand U1684 (N_1684,N_895,N_1177);
nor U1685 (N_1685,N_645,N_1105);
nor U1686 (N_1686,N_738,N_974);
and U1687 (N_1687,N_711,N_928);
or U1688 (N_1688,N_1143,N_841);
xnor U1689 (N_1689,N_992,N_680);
and U1690 (N_1690,N_790,N_858);
nor U1691 (N_1691,N_971,N_665);
and U1692 (N_1692,N_891,N_1145);
and U1693 (N_1693,N_1085,N_1009);
or U1694 (N_1694,N_1034,N_1077);
nor U1695 (N_1695,N_980,N_679);
nor U1696 (N_1696,N_612,N_1045);
or U1697 (N_1697,N_1030,N_635);
nand U1698 (N_1698,N_665,N_652);
nor U1699 (N_1699,N_1034,N_1124);
or U1700 (N_1700,N_779,N_886);
nor U1701 (N_1701,N_1032,N_678);
nand U1702 (N_1702,N_677,N_900);
nand U1703 (N_1703,N_888,N_984);
nand U1704 (N_1704,N_1006,N_678);
xnor U1705 (N_1705,N_1179,N_1043);
xnor U1706 (N_1706,N_1180,N_958);
nor U1707 (N_1707,N_1176,N_864);
nand U1708 (N_1708,N_846,N_1179);
nor U1709 (N_1709,N_744,N_1092);
or U1710 (N_1710,N_993,N_605);
nor U1711 (N_1711,N_811,N_918);
xor U1712 (N_1712,N_1066,N_671);
nor U1713 (N_1713,N_1110,N_759);
or U1714 (N_1714,N_905,N_1192);
nand U1715 (N_1715,N_664,N_1187);
or U1716 (N_1716,N_620,N_959);
or U1717 (N_1717,N_1193,N_701);
xnor U1718 (N_1718,N_834,N_617);
and U1719 (N_1719,N_998,N_1192);
nor U1720 (N_1720,N_630,N_934);
xor U1721 (N_1721,N_697,N_976);
nor U1722 (N_1722,N_1186,N_1029);
nor U1723 (N_1723,N_993,N_878);
xor U1724 (N_1724,N_822,N_812);
or U1725 (N_1725,N_690,N_1114);
or U1726 (N_1726,N_704,N_1177);
and U1727 (N_1727,N_725,N_639);
or U1728 (N_1728,N_1167,N_723);
or U1729 (N_1729,N_741,N_941);
nand U1730 (N_1730,N_1072,N_957);
nand U1731 (N_1731,N_740,N_1062);
nor U1732 (N_1732,N_1141,N_1008);
and U1733 (N_1733,N_1196,N_894);
nand U1734 (N_1734,N_874,N_822);
nor U1735 (N_1735,N_708,N_971);
nand U1736 (N_1736,N_938,N_1092);
nand U1737 (N_1737,N_723,N_672);
or U1738 (N_1738,N_786,N_1075);
nand U1739 (N_1739,N_988,N_648);
or U1740 (N_1740,N_843,N_1081);
and U1741 (N_1741,N_699,N_641);
nand U1742 (N_1742,N_748,N_777);
nand U1743 (N_1743,N_859,N_960);
xor U1744 (N_1744,N_1116,N_1087);
nand U1745 (N_1745,N_1011,N_705);
or U1746 (N_1746,N_1199,N_871);
or U1747 (N_1747,N_643,N_773);
nand U1748 (N_1748,N_1043,N_897);
nand U1749 (N_1749,N_635,N_745);
or U1750 (N_1750,N_969,N_1039);
xor U1751 (N_1751,N_917,N_867);
or U1752 (N_1752,N_1058,N_921);
nor U1753 (N_1753,N_951,N_823);
and U1754 (N_1754,N_690,N_958);
and U1755 (N_1755,N_908,N_839);
and U1756 (N_1756,N_913,N_1053);
or U1757 (N_1757,N_771,N_741);
or U1758 (N_1758,N_932,N_623);
xnor U1759 (N_1759,N_1064,N_713);
nor U1760 (N_1760,N_850,N_1100);
nor U1761 (N_1761,N_754,N_848);
xor U1762 (N_1762,N_690,N_1077);
or U1763 (N_1763,N_954,N_828);
nor U1764 (N_1764,N_826,N_1109);
and U1765 (N_1765,N_873,N_629);
xor U1766 (N_1766,N_1090,N_986);
and U1767 (N_1767,N_1024,N_1072);
or U1768 (N_1768,N_791,N_1034);
or U1769 (N_1769,N_854,N_728);
xor U1770 (N_1770,N_666,N_760);
nor U1771 (N_1771,N_733,N_1125);
and U1772 (N_1772,N_790,N_733);
xnor U1773 (N_1773,N_798,N_702);
or U1774 (N_1774,N_865,N_691);
nor U1775 (N_1775,N_883,N_1199);
or U1776 (N_1776,N_682,N_992);
nand U1777 (N_1777,N_1079,N_755);
nor U1778 (N_1778,N_1038,N_1111);
nand U1779 (N_1779,N_871,N_667);
nand U1780 (N_1780,N_712,N_1179);
and U1781 (N_1781,N_646,N_1090);
xnor U1782 (N_1782,N_939,N_1146);
xnor U1783 (N_1783,N_751,N_1005);
or U1784 (N_1784,N_1111,N_1108);
nor U1785 (N_1785,N_908,N_1058);
or U1786 (N_1786,N_1036,N_814);
nand U1787 (N_1787,N_662,N_856);
and U1788 (N_1788,N_665,N_886);
and U1789 (N_1789,N_1038,N_605);
nor U1790 (N_1790,N_886,N_1171);
nor U1791 (N_1791,N_1154,N_852);
and U1792 (N_1792,N_747,N_679);
nor U1793 (N_1793,N_696,N_1016);
xor U1794 (N_1794,N_684,N_1179);
or U1795 (N_1795,N_1078,N_721);
nor U1796 (N_1796,N_603,N_976);
or U1797 (N_1797,N_998,N_794);
nor U1798 (N_1798,N_858,N_925);
nand U1799 (N_1799,N_704,N_1141);
or U1800 (N_1800,N_1767,N_1258);
or U1801 (N_1801,N_1226,N_1592);
nor U1802 (N_1802,N_1380,N_1751);
or U1803 (N_1803,N_1462,N_1401);
or U1804 (N_1804,N_1383,N_1400);
nor U1805 (N_1805,N_1288,N_1270);
and U1806 (N_1806,N_1218,N_1627);
and U1807 (N_1807,N_1696,N_1614);
nor U1808 (N_1808,N_1563,N_1640);
nand U1809 (N_1809,N_1312,N_1345);
and U1810 (N_1810,N_1395,N_1608);
and U1811 (N_1811,N_1513,N_1552);
nor U1812 (N_1812,N_1799,N_1720);
nand U1813 (N_1813,N_1209,N_1330);
nor U1814 (N_1814,N_1570,N_1474);
and U1815 (N_1815,N_1337,N_1680);
nor U1816 (N_1816,N_1564,N_1622);
nor U1817 (N_1817,N_1795,N_1535);
and U1818 (N_1818,N_1568,N_1508);
and U1819 (N_1819,N_1755,N_1675);
nand U1820 (N_1820,N_1211,N_1743);
or U1821 (N_1821,N_1545,N_1710);
or U1822 (N_1822,N_1749,N_1346);
and U1823 (N_1823,N_1398,N_1217);
xor U1824 (N_1824,N_1632,N_1269);
and U1825 (N_1825,N_1382,N_1309);
and U1826 (N_1826,N_1770,N_1559);
and U1827 (N_1827,N_1365,N_1277);
nor U1828 (N_1828,N_1734,N_1514);
nor U1829 (N_1829,N_1452,N_1421);
xor U1830 (N_1830,N_1342,N_1373);
and U1831 (N_1831,N_1348,N_1470);
nor U1832 (N_1832,N_1263,N_1408);
and U1833 (N_1833,N_1260,N_1284);
or U1834 (N_1834,N_1569,N_1688);
nor U1835 (N_1835,N_1293,N_1453);
nor U1836 (N_1836,N_1724,N_1550);
or U1837 (N_1837,N_1325,N_1369);
or U1838 (N_1838,N_1245,N_1281);
or U1839 (N_1839,N_1443,N_1718);
or U1840 (N_1840,N_1643,N_1723);
nor U1841 (N_1841,N_1250,N_1705);
or U1842 (N_1842,N_1339,N_1310);
xnor U1843 (N_1843,N_1684,N_1206);
xor U1844 (N_1844,N_1596,N_1612);
nor U1845 (N_1845,N_1789,N_1754);
or U1846 (N_1846,N_1798,N_1220);
nand U1847 (N_1847,N_1756,N_1660);
xnor U1848 (N_1848,N_1457,N_1690);
or U1849 (N_1849,N_1685,N_1308);
xnor U1850 (N_1850,N_1602,N_1628);
or U1851 (N_1851,N_1529,N_1794);
nor U1852 (N_1852,N_1673,N_1577);
nand U1853 (N_1853,N_1431,N_1573);
and U1854 (N_1854,N_1547,N_1735);
nand U1855 (N_1855,N_1594,N_1322);
xnor U1856 (N_1856,N_1387,N_1674);
and U1857 (N_1857,N_1253,N_1787);
or U1858 (N_1858,N_1448,N_1279);
and U1859 (N_1859,N_1469,N_1423);
or U1860 (N_1860,N_1638,N_1426);
and U1861 (N_1861,N_1571,N_1483);
or U1862 (N_1862,N_1522,N_1273);
nand U1863 (N_1863,N_1721,N_1671);
and U1864 (N_1864,N_1579,N_1344);
and U1865 (N_1865,N_1641,N_1392);
or U1866 (N_1866,N_1587,N_1501);
or U1867 (N_1867,N_1302,N_1733);
nor U1868 (N_1868,N_1444,N_1357);
and U1869 (N_1869,N_1766,N_1757);
nor U1870 (N_1870,N_1677,N_1333);
or U1871 (N_1871,N_1737,N_1617);
xnor U1872 (N_1872,N_1497,N_1630);
xnor U1873 (N_1873,N_1764,N_1238);
or U1874 (N_1874,N_1399,N_1739);
nand U1875 (N_1875,N_1229,N_1374);
and U1876 (N_1876,N_1222,N_1366);
and U1877 (N_1877,N_1326,N_1275);
nor U1878 (N_1878,N_1285,N_1420);
and U1879 (N_1879,N_1347,N_1396);
or U1880 (N_1880,N_1364,N_1416);
and U1881 (N_1881,N_1664,N_1466);
or U1882 (N_1882,N_1580,N_1358);
xnor U1883 (N_1883,N_1318,N_1572);
or U1884 (N_1884,N_1538,N_1693);
nand U1885 (N_1885,N_1615,N_1409);
or U1886 (N_1886,N_1445,N_1338);
and U1887 (N_1887,N_1502,N_1629);
nor U1888 (N_1888,N_1717,N_1781);
and U1889 (N_1889,N_1243,N_1419);
nand U1890 (N_1890,N_1311,N_1565);
and U1891 (N_1891,N_1236,N_1256);
nand U1892 (N_1892,N_1758,N_1642);
xnor U1893 (N_1893,N_1670,N_1556);
xor U1894 (N_1894,N_1598,N_1621);
and U1895 (N_1895,N_1562,N_1210);
and U1896 (N_1896,N_1404,N_1593);
nand U1897 (N_1897,N_1287,N_1410);
or U1898 (N_1898,N_1495,N_1661);
nor U1899 (N_1899,N_1200,N_1653);
nand U1900 (N_1900,N_1438,N_1456);
nor U1901 (N_1901,N_1205,N_1247);
xor U1902 (N_1902,N_1481,N_1519);
and U1903 (N_1903,N_1533,N_1768);
or U1904 (N_1904,N_1613,N_1499);
or U1905 (N_1905,N_1320,N_1707);
and U1906 (N_1906,N_1526,N_1434);
nand U1907 (N_1907,N_1595,N_1397);
xnor U1908 (N_1908,N_1703,N_1729);
nand U1909 (N_1909,N_1271,N_1249);
nand U1910 (N_1910,N_1225,N_1785);
and U1911 (N_1911,N_1738,N_1414);
nand U1912 (N_1912,N_1528,N_1731);
nand U1913 (N_1913,N_1202,N_1566);
xor U1914 (N_1914,N_1272,N_1665);
or U1915 (N_1915,N_1385,N_1510);
or U1916 (N_1916,N_1544,N_1407);
nor U1917 (N_1917,N_1235,N_1644);
and U1918 (N_1918,N_1626,N_1433);
or U1919 (N_1919,N_1760,N_1578);
and U1920 (N_1920,N_1561,N_1694);
nor U1921 (N_1921,N_1553,N_1403);
nor U1922 (N_1922,N_1362,N_1241);
xor U1923 (N_1923,N_1771,N_1582);
nand U1924 (N_1924,N_1511,N_1790);
nor U1925 (N_1925,N_1759,N_1542);
xor U1926 (N_1926,N_1716,N_1478);
nor U1927 (N_1927,N_1278,N_1714);
and U1928 (N_1928,N_1231,N_1482);
nor U1929 (N_1929,N_1777,N_1468);
and U1930 (N_1930,N_1728,N_1605);
nand U1931 (N_1931,N_1585,N_1435);
xnor U1932 (N_1932,N_1662,N_1753);
or U1933 (N_1933,N_1363,N_1681);
or U1934 (N_1934,N_1201,N_1744);
or U1935 (N_1935,N_1389,N_1575);
xnor U1936 (N_1936,N_1543,N_1240);
and U1937 (N_1937,N_1666,N_1750);
nor U1938 (N_1938,N_1207,N_1340);
or U1939 (N_1939,N_1725,N_1336);
nand U1940 (N_1940,N_1541,N_1518);
xor U1941 (N_1941,N_1221,N_1525);
xnor U1942 (N_1942,N_1415,N_1224);
xor U1943 (N_1943,N_1476,N_1442);
or U1944 (N_1944,N_1450,N_1359);
or U1945 (N_1945,N_1252,N_1736);
xor U1946 (N_1946,N_1289,N_1603);
nand U1947 (N_1947,N_1485,N_1449);
and U1948 (N_1948,N_1490,N_1548);
nor U1949 (N_1949,N_1464,N_1496);
xnor U1950 (N_1950,N_1506,N_1687);
nor U1951 (N_1951,N_1554,N_1586);
xnor U1952 (N_1952,N_1583,N_1254);
xor U1953 (N_1953,N_1261,N_1659);
and U1954 (N_1954,N_1712,N_1355);
nor U1955 (N_1955,N_1321,N_1623);
xor U1956 (N_1956,N_1491,N_1237);
and U1957 (N_1957,N_1428,N_1599);
or U1958 (N_1958,N_1708,N_1331);
nand U1959 (N_1959,N_1430,N_1588);
nor U1960 (N_1960,N_1604,N_1391);
nand U1961 (N_1961,N_1276,N_1793);
nand U1962 (N_1962,N_1370,N_1591);
nor U1963 (N_1963,N_1292,N_1779);
nor U1964 (N_1964,N_1204,N_1424);
and U1965 (N_1965,N_1300,N_1551);
xor U1966 (N_1966,N_1504,N_1699);
nor U1967 (N_1967,N_1778,N_1298);
xor U1968 (N_1968,N_1214,N_1780);
xnor U1969 (N_1969,N_1334,N_1763);
or U1970 (N_1970,N_1652,N_1500);
and U1971 (N_1971,N_1650,N_1625);
nor U1972 (N_1972,N_1371,N_1746);
and U1973 (N_1973,N_1631,N_1440);
nor U1974 (N_1974,N_1709,N_1691);
or U1975 (N_1975,N_1676,N_1546);
nand U1976 (N_1976,N_1488,N_1555);
and U1977 (N_1977,N_1507,N_1290);
or U1978 (N_1978,N_1792,N_1411);
nor U1979 (N_1979,N_1557,N_1378);
nand U1980 (N_1980,N_1446,N_1668);
or U1981 (N_1981,N_1259,N_1244);
nor U1982 (N_1982,N_1493,N_1697);
nor U1983 (N_1983,N_1647,N_1698);
xnor U1984 (N_1984,N_1472,N_1447);
nand U1985 (N_1985,N_1796,N_1223);
or U1986 (N_1986,N_1784,N_1576);
and U1987 (N_1987,N_1306,N_1212);
nand U1988 (N_1988,N_1248,N_1748);
and U1989 (N_1989,N_1461,N_1203);
and U1990 (N_1990,N_1667,N_1351);
or U1991 (N_1991,N_1479,N_1618);
nand U1992 (N_1992,N_1327,N_1639);
xor U1993 (N_1993,N_1633,N_1772);
nor U1994 (N_1994,N_1536,N_1295);
nand U1995 (N_1995,N_1460,N_1219);
nor U1996 (N_1996,N_1658,N_1390);
xor U1997 (N_1997,N_1762,N_1689);
nand U1998 (N_1998,N_1524,N_1480);
or U1999 (N_1999,N_1624,N_1422);
nor U2000 (N_2000,N_1268,N_1324);
or U2001 (N_2001,N_1607,N_1727);
and U2002 (N_2002,N_1567,N_1558);
and U2003 (N_2003,N_1636,N_1646);
or U2004 (N_2004,N_1465,N_1341);
nor U2005 (N_2005,N_1280,N_1537);
and U2006 (N_2006,N_1701,N_1797);
or U2007 (N_2007,N_1523,N_1328);
and U2008 (N_2008,N_1406,N_1726);
and U2009 (N_2009,N_1242,N_1706);
and U2010 (N_2010,N_1540,N_1711);
or U2011 (N_2011,N_1264,N_1294);
or U2012 (N_2012,N_1686,N_1305);
nor U2013 (N_2013,N_1314,N_1560);
nor U2014 (N_2014,N_1335,N_1730);
nor U2015 (N_2015,N_1377,N_1429);
and U2016 (N_2016,N_1329,N_1375);
and U2017 (N_2017,N_1776,N_1505);
and U2018 (N_2018,N_1317,N_1427);
nand U2019 (N_2019,N_1682,N_1520);
nor U2020 (N_2020,N_1360,N_1352);
nand U2021 (N_2021,N_1301,N_1274);
or U2022 (N_2022,N_1791,N_1299);
and U2023 (N_2023,N_1255,N_1307);
and U2024 (N_2024,N_1246,N_1788);
and U2025 (N_2025,N_1234,N_1740);
nor U2026 (N_2026,N_1425,N_1637);
or U2027 (N_2027,N_1498,N_1402);
nor U2028 (N_2028,N_1303,N_1475);
nor U2029 (N_2029,N_1531,N_1601);
nor U2030 (N_2030,N_1649,N_1648);
xor U2031 (N_2031,N_1509,N_1645);
nor U2032 (N_2032,N_1609,N_1527);
and U2033 (N_2033,N_1620,N_1319);
and U2034 (N_2034,N_1635,N_1437);
and U2035 (N_2035,N_1678,N_1257);
xnor U2036 (N_2036,N_1775,N_1413);
and U2037 (N_2037,N_1379,N_1741);
nand U2038 (N_2038,N_1417,N_1463);
nand U2039 (N_2039,N_1584,N_1367);
and U2040 (N_2040,N_1765,N_1393);
xnor U2041 (N_2041,N_1655,N_1656);
xor U2042 (N_2042,N_1532,N_1376);
xnor U2043 (N_2043,N_1286,N_1323);
or U2044 (N_2044,N_1215,N_1774);
nand U2045 (N_2045,N_1384,N_1267);
nor U2046 (N_2046,N_1503,N_1669);
nand U2047 (N_2047,N_1683,N_1769);
nor U2048 (N_2048,N_1432,N_1651);
or U2049 (N_2049,N_1233,N_1230);
nor U2050 (N_2050,N_1232,N_1486);
nor U2051 (N_2051,N_1418,N_1386);
or U2052 (N_2052,N_1654,N_1657);
nor U2053 (N_2053,N_1265,N_1606);
and U2054 (N_2054,N_1239,N_1451);
nand U2055 (N_2055,N_1782,N_1549);
nand U2056 (N_2056,N_1719,N_1368);
or U2057 (N_2057,N_1539,N_1467);
or U2058 (N_2058,N_1304,N_1332);
nor U2059 (N_2059,N_1471,N_1732);
or U2060 (N_2060,N_1589,N_1600);
or U2061 (N_2061,N_1313,N_1349);
nand U2062 (N_2062,N_1492,N_1394);
and U2063 (N_2063,N_1356,N_1610);
or U2064 (N_2064,N_1262,N_1745);
nand U2065 (N_2065,N_1679,N_1534);
or U2066 (N_2066,N_1530,N_1619);
nand U2067 (N_2067,N_1405,N_1516);
nor U2068 (N_2068,N_1700,N_1266);
nor U2069 (N_2069,N_1574,N_1590);
nor U2070 (N_2070,N_1512,N_1489);
or U2071 (N_2071,N_1484,N_1350);
or U2072 (N_2072,N_1439,N_1441);
nor U2073 (N_2073,N_1715,N_1455);
or U2074 (N_2074,N_1412,N_1353);
nand U2075 (N_2075,N_1704,N_1316);
nand U2076 (N_2076,N_1722,N_1477);
nor U2077 (N_2077,N_1786,N_1515);
xor U2078 (N_2078,N_1663,N_1283);
or U2079 (N_2079,N_1672,N_1459);
nor U2080 (N_2080,N_1381,N_1747);
nand U2081 (N_2081,N_1361,N_1695);
and U2082 (N_2082,N_1597,N_1692);
nand U2083 (N_2083,N_1291,N_1473);
or U2084 (N_2084,N_1521,N_1783);
nand U2085 (N_2085,N_1494,N_1343);
or U2086 (N_2086,N_1388,N_1436);
nor U2087 (N_2087,N_1216,N_1752);
or U2088 (N_2088,N_1761,N_1208);
nand U2089 (N_2089,N_1581,N_1282);
nor U2090 (N_2090,N_1251,N_1454);
nor U2091 (N_2091,N_1616,N_1372);
xor U2092 (N_2092,N_1634,N_1517);
nor U2093 (N_2093,N_1742,N_1702);
nand U2094 (N_2094,N_1213,N_1297);
and U2095 (N_2095,N_1296,N_1773);
xor U2096 (N_2096,N_1487,N_1228);
and U2097 (N_2097,N_1611,N_1458);
or U2098 (N_2098,N_1315,N_1227);
xor U2099 (N_2099,N_1354,N_1713);
and U2100 (N_2100,N_1354,N_1299);
nor U2101 (N_2101,N_1637,N_1289);
and U2102 (N_2102,N_1348,N_1506);
nor U2103 (N_2103,N_1588,N_1542);
nor U2104 (N_2104,N_1753,N_1777);
xor U2105 (N_2105,N_1350,N_1533);
xnor U2106 (N_2106,N_1536,N_1361);
or U2107 (N_2107,N_1522,N_1470);
or U2108 (N_2108,N_1787,N_1771);
nand U2109 (N_2109,N_1342,N_1671);
nand U2110 (N_2110,N_1257,N_1242);
nor U2111 (N_2111,N_1202,N_1210);
and U2112 (N_2112,N_1492,N_1423);
and U2113 (N_2113,N_1528,N_1589);
and U2114 (N_2114,N_1559,N_1786);
or U2115 (N_2115,N_1643,N_1463);
and U2116 (N_2116,N_1778,N_1564);
and U2117 (N_2117,N_1573,N_1740);
or U2118 (N_2118,N_1767,N_1245);
or U2119 (N_2119,N_1492,N_1757);
and U2120 (N_2120,N_1402,N_1445);
and U2121 (N_2121,N_1212,N_1433);
and U2122 (N_2122,N_1349,N_1546);
xnor U2123 (N_2123,N_1635,N_1628);
or U2124 (N_2124,N_1585,N_1427);
nor U2125 (N_2125,N_1251,N_1465);
and U2126 (N_2126,N_1385,N_1234);
nor U2127 (N_2127,N_1695,N_1579);
and U2128 (N_2128,N_1259,N_1686);
nor U2129 (N_2129,N_1210,N_1509);
nor U2130 (N_2130,N_1303,N_1678);
nor U2131 (N_2131,N_1709,N_1481);
and U2132 (N_2132,N_1628,N_1203);
and U2133 (N_2133,N_1403,N_1308);
or U2134 (N_2134,N_1429,N_1696);
nand U2135 (N_2135,N_1305,N_1479);
nor U2136 (N_2136,N_1484,N_1531);
nand U2137 (N_2137,N_1407,N_1533);
or U2138 (N_2138,N_1661,N_1670);
or U2139 (N_2139,N_1690,N_1754);
nor U2140 (N_2140,N_1513,N_1714);
and U2141 (N_2141,N_1513,N_1309);
and U2142 (N_2142,N_1341,N_1683);
and U2143 (N_2143,N_1645,N_1389);
nor U2144 (N_2144,N_1598,N_1783);
nand U2145 (N_2145,N_1711,N_1776);
nor U2146 (N_2146,N_1330,N_1789);
or U2147 (N_2147,N_1408,N_1443);
nor U2148 (N_2148,N_1604,N_1714);
or U2149 (N_2149,N_1458,N_1389);
and U2150 (N_2150,N_1706,N_1744);
nor U2151 (N_2151,N_1653,N_1502);
nor U2152 (N_2152,N_1233,N_1591);
nand U2153 (N_2153,N_1668,N_1493);
and U2154 (N_2154,N_1423,N_1748);
nor U2155 (N_2155,N_1740,N_1244);
and U2156 (N_2156,N_1407,N_1245);
xnor U2157 (N_2157,N_1738,N_1616);
or U2158 (N_2158,N_1714,N_1659);
nor U2159 (N_2159,N_1445,N_1214);
nand U2160 (N_2160,N_1287,N_1639);
nand U2161 (N_2161,N_1505,N_1278);
nor U2162 (N_2162,N_1224,N_1570);
nand U2163 (N_2163,N_1775,N_1588);
nand U2164 (N_2164,N_1518,N_1741);
nor U2165 (N_2165,N_1656,N_1262);
nor U2166 (N_2166,N_1209,N_1503);
nor U2167 (N_2167,N_1779,N_1498);
and U2168 (N_2168,N_1637,N_1506);
and U2169 (N_2169,N_1545,N_1393);
nand U2170 (N_2170,N_1740,N_1381);
xor U2171 (N_2171,N_1690,N_1328);
nand U2172 (N_2172,N_1790,N_1210);
or U2173 (N_2173,N_1511,N_1449);
nand U2174 (N_2174,N_1709,N_1227);
nor U2175 (N_2175,N_1264,N_1265);
and U2176 (N_2176,N_1272,N_1487);
and U2177 (N_2177,N_1278,N_1792);
and U2178 (N_2178,N_1521,N_1604);
and U2179 (N_2179,N_1733,N_1591);
or U2180 (N_2180,N_1273,N_1227);
nand U2181 (N_2181,N_1394,N_1683);
nand U2182 (N_2182,N_1712,N_1266);
or U2183 (N_2183,N_1281,N_1405);
or U2184 (N_2184,N_1340,N_1494);
nor U2185 (N_2185,N_1790,N_1316);
and U2186 (N_2186,N_1733,N_1553);
nand U2187 (N_2187,N_1716,N_1200);
nor U2188 (N_2188,N_1750,N_1644);
nor U2189 (N_2189,N_1347,N_1261);
nand U2190 (N_2190,N_1220,N_1774);
nand U2191 (N_2191,N_1522,N_1390);
nor U2192 (N_2192,N_1206,N_1609);
nand U2193 (N_2193,N_1795,N_1377);
nand U2194 (N_2194,N_1532,N_1748);
nor U2195 (N_2195,N_1339,N_1480);
or U2196 (N_2196,N_1654,N_1292);
and U2197 (N_2197,N_1504,N_1322);
and U2198 (N_2198,N_1336,N_1239);
nor U2199 (N_2199,N_1615,N_1401);
and U2200 (N_2200,N_1755,N_1727);
and U2201 (N_2201,N_1200,N_1472);
nor U2202 (N_2202,N_1227,N_1735);
nor U2203 (N_2203,N_1715,N_1766);
and U2204 (N_2204,N_1656,N_1298);
xnor U2205 (N_2205,N_1247,N_1307);
or U2206 (N_2206,N_1754,N_1493);
or U2207 (N_2207,N_1272,N_1661);
xnor U2208 (N_2208,N_1631,N_1637);
and U2209 (N_2209,N_1399,N_1758);
nor U2210 (N_2210,N_1510,N_1421);
or U2211 (N_2211,N_1211,N_1559);
nand U2212 (N_2212,N_1255,N_1548);
nor U2213 (N_2213,N_1565,N_1708);
nor U2214 (N_2214,N_1202,N_1442);
xor U2215 (N_2215,N_1477,N_1491);
and U2216 (N_2216,N_1315,N_1770);
nor U2217 (N_2217,N_1399,N_1203);
nand U2218 (N_2218,N_1697,N_1385);
nand U2219 (N_2219,N_1292,N_1466);
or U2220 (N_2220,N_1266,N_1778);
or U2221 (N_2221,N_1377,N_1416);
or U2222 (N_2222,N_1356,N_1785);
and U2223 (N_2223,N_1502,N_1590);
and U2224 (N_2224,N_1668,N_1410);
or U2225 (N_2225,N_1436,N_1260);
or U2226 (N_2226,N_1502,N_1396);
nor U2227 (N_2227,N_1206,N_1463);
nor U2228 (N_2228,N_1302,N_1266);
xnor U2229 (N_2229,N_1539,N_1213);
or U2230 (N_2230,N_1612,N_1276);
or U2231 (N_2231,N_1398,N_1470);
or U2232 (N_2232,N_1618,N_1334);
or U2233 (N_2233,N_1229,N_1485);
nor U2234 (N_2234,N_1402,N_1795);
and U2235 (N_2235,N_1794,N_1448);
nand U2236 (N_2236,N_1524,N_1621);
or U2237 (N_2237,N_1765,N_1731);
and U2238 (N_2238,N_1339,N_1597);
and U2239 (N_2239,N_1289,N_1436);
nand U2240 (N_2240,N_1561,N_1643);
and U2241 (N_2241,N_1457,N_1579);
nor U2242 (N_2242,N_1654,N_1485);
nor U2243 (N_2243,N_1751,N_1298);
and U2244 (N_2244,N_1410,N_1483);
and U2245 (N_2245,N_1388,N_1690);
nand U2246 (N_2246,N_1525,N_1386);
and U2247 (N_2247,N_1581,N_1601);
nand U2248 (N_2248,N_1592,N_1381);
or U2249 (N_2249,N_1200,N_1606);
or U2250 (N_2250,N_1523,N_1792);
nand U2251 (N_2251,N_1257,N_1227);
nand U2252 (N_2252,N_1207,N_1609);
or U2253 (N_2253,N_1518,N_1313);
nor U2254 (N_2254,N_1708,N_1635);
nor U2255 (N_2255,N_1635,N_1363);
and U2256 (N_2256,N_1672,N_1608);
nor U2257 (N_2257,N_1592,N_1555);
nor U2258 (N_2258,N_1630,N_1412);
nand U2259 (N_2259,N_1508,N_1662);
or U2260 (N_2260,N_1619,N_1765);
or U2261 (N_2261,N_1207,N_1725);
or U2262 (N_2262,N_1237,N_1268);
nor U2263 (N_2263,N_1764,N_1560);
and U2264 (N_2264,N_1519,N_1677);
nand U2265 (N_2265,N_1501,N_1395);
xnor U2266 (N_2266,N_1408,N_1466);
and U2267 (N_2267,N_1623,N_1262);
nand U2268 (N_2268,N_1498,N_1610);
nand U2269 (N_2269,N_1448,N_1630);
or U2270 (N_2270,N_1461,N_1650);
and U2271 (N_2271,N_1253,N_1417);
and U2272 (N_2272,N_1501,N_1319);
or U2273 (N_2273,N_1219,N_1353);
or U2274 (N_2274,N_1358,N_1412);
nor U2275 (N_2275,N_1696,N_1431);
and U2276 (N_2276,N_1568,N_1577);
nand U2277 (N_2277,N_1767,N_1377);
and U2278 (N_2278,N_1324,N_1279);
nand U2279 (N_2279,N_1296,N_1765);
nor U2280 (N_2280,N_1789,N_1236);
xnor U2281 (N_2281,N_1535,N_1418);
nor U2282 (N_2282,N_1218,N_1513);
and U2283 (N_2283,N_1292,N_1412);
and U2284 (N_2284,N_1666,N_1691);
xor U2285 (N_2285,N_1320,N_1538);
nor U2286 (N_2286,N_1612,N_1351);
nor U2287 (N_2287,N_1793,N_1374);
nor U2288 (N_2288,N_1462,N_1349);
nand U2289 (N_2289,N_1341,N_1672);
nor U2290 (N_2290,N_1361,N_1459);
and U2291 (N_2291,N_1250,N_1434);
and U2292 (N_2292,N_1783,N_1734);
and U2293 (N_2293,N_1786,N_1531);
or U2294 (N_2294,N_1335,N_1600);
and U2295 (N_2295,N_1533,N_1594);
nor U2296 (N_2296,N_1728,N_1376);
nor U2297 (N_2297,N_1282,N_1672);
nand U2298 (N_2298,N_1294,N_1321);
nor U2299 (N_2299,N_1749,N_1267);
nand U2300 (N_2300,N_1570,N_1458);
nand U2301 (N_2301,N_1445,N_1341);
and U2302 (N_2302,N_1640,N_1326);
nand U2303 (N_2303,N_1245,N_1789);
and U2304 (N_2304,N_1403,N_1633);
xnor U2305 (N_2305,N_1503,N_1274);
nor U2306 (N_2306,N_1288,N_1402);
or U2307 (N_2307,N_1778,N_1588);
xor U2308 (N_2308,N_1349,N_1432);
nor U2309 (N_2309,N_1225,N_1207);
nand U2310 (N_2310,N_1554,N_1331);
and U2311 (N_2311,N_1674,N_1750);
or U2312 (N_2312,N_1399,N_1570);
nor U2313 (N_2313,N_1307,N_1657);
nor U2314 (N_2314,N_1479,N_1668);
nand U2315 (N_2315,N_1430,N_1214);
and U2316 (N_2316,N_1619,N_1605);
nor U2317 (N_2317,N_1508,N_1277);
nor U2318 (N_2318,N_1561,N_1598);
or U2319 (N_2319,N_1530,N_1531);
and U2320 (N_2320,N_1396,N_1666);
nand U2321 (N_2321,N_1761,N_1272);
nand U2322 (N_2322,N_1668,N_1482);
xor U2323 (N_2323,N_1760,N_1507);
xnor U2324 (N_2324,N_1421,N_1263);
nand U2325 (N_2325,N_1355,N_1606);
or U2326 (N_2326,N_1479,N_1771);
nor U2327 (N_2327,N_1485,N_1684);
xor U2328 (N_2328,N_1758,N_1431);
nor U2329 (N_2329,N_1675,N_1301);
and U2330 (N_2330,N_1655,N_1290);
or U2331 (N_2331,N_1588,N_1244);
nand U2332 (N_2332,N_1502,N_1373);
nand U2333 (N_2333,N_1608,N_1425);
and U2334 (N_2334,N_1703,N_1796);
or U2335 (N_2335,N_1426,N_1281);
nor U2336 (N_2336,N_1640,N_1419);
nor U2337 (N_2337,N_1559,N_1634);
or U2338 (N_2338,N_1637,N_1706);
or U2339 (N_2339,N_1366,N_1237);
and U2340 (N_2340,N_1267,N_1210);
and U2341 (N_2341,N_1289,N_1643);
or U2342 (N_2342,N_1277,N_1691);
and U2343 (N_2343,N_1257,N_1367);
nor U2344 (N_2344,N_1696,N_1414);
nor U2345 (N_2345,N_1643,N_1786);
nand U2346 (N_2346,N_1426,N_1405);
nand U2347 (N_2347,N_1300,N_1371);
or U2348 (N_2348,N_1640,N_1569);
nand U2349 (N_2349,N_1365,N_1346);
or U2350 (N_2350,N_1205,N_1581);
nand U2351 (N_2351,N_1746,N_1300);
xor U2352 (N_2352,N_1354,N_1264);
xnor U2353 (N_2353,N_1305,N_1515);
xor U2354 (N_2354,N_1650,N_1688);
nand U2355 (N_2355,N_1340,N_1566);
nand U2356 (N_2356,N_1441,N_1708);
nand U2357 (N_2357,N_1716,N_1702);
and U2358 (N_2358,N_1404,N_1301);
nor U2359 (N_2359,N_1324,N_1486);
or U2360 (N_2360,N_1245,N_1494);
nor U2361 (N_2361,N_1432,N_1463);
nor U2362 (N_2362,N_1765,N_1486);
nor U2363 (N_2363,N_1438,N_1786);
nor U2364 (N_2364,N_1312,N_1786);
and U2365 (N_2365,N_1700,N_1707);
or U2366 (N_2366,N_1500,N_1735);
nand U2367 (N_2367,N_1238,N_1498);
and U2368 (N_2368,N_1479,N_1760);
nor U2369 (N_2369,N_1694,N_1330);
and U2370 (N_2370,N_1465,N_1536);
and U2371 (N_2371,N_1542,N_1492);
nand U2372 (N_2372,N_1626,N_1560);
nand U2373 (N_2373,N_1450,N_1305);
or U2374 (N_2374,N_1237,N_1547);
and U2375 (N_2375,N_1495,N_1739);
nand U2376 (N_2376,N_1763,N_1753);
and U2377 (N_2377,N_1503,N_1373);
or U2378 (N_2378,N_1399,N_1228);
or U2379 (N_2379,N_1775,N_1208);
or U2380 (N_2380,N_1672,N_1614);
nor U2381 (N_2381,N_1630,N_1626);
and U2382 (N_2382,N_1399,N_1225);
nand U2383 (N_2383,N_1267,N_1765);
or U2384 (N_2384,N_1396,N_1337);
nand U2385 (N_2385,N_1773,N_1495);
or U2386 (N_2386,N_1564,N_1656);
xor U2387 (N_2387,N_1436,N_1734);
xnor U2388 (N_2388,N_1546,N_1588);
and U2389 (N_2389,N_1708,N_1660);
and U2390 (N_2390,N_1432,N_1274);
or U2391 (N_2391,N_1400,N_1231);
and U2392 (N_2392,N_1731,N_1359);
and U2393 (N_2393,N_1531,N_1251);
or U2394 (N_2394,N_1436,N_1656);
nor U2395 (N_2395,N_1583,N_1460);
xor U2396 (N_2396,N_1643,N_1313);
nor U2397 (N_2397,N_1534,N_1375);
and U2398 (N_2398,N_1782,N_1504);
and U2399 (N_2399,N_1775,N_1720);
or U2400 (N_2400,N_1954,N_1992);
and U2401 (N_2401,N_2282,N_1867);
nand U2402 (N_2402,N_2091,N_2126);
or U2403 (N_2403,N_2326,N_2379);
nand U2404 (N_2404,N_2382,N_2195);
nor U2405 (N_2405,N_1920,N_2045);
xor U2406 (N_2406,N_2308,N_2303);
xnor U2407 (N_2407,N_2322,N_2048);
nor U2408 (N_2408,N_2294,N_1840);
or U2409 (N_2409,N_2118,N_1806);
and U2410 (N_2410,N_2176,N_2177);
nand U2411 (N_2411,N_1851,N_2287);
nor U2412 (N_2412,N_2312,N_2265);
nor U2413 (N_2413,N_2119,N_2068);
xor U2414 (N_2414,N_2135,N_2384);
or U2415 (N_2415,N_2125,N_1937);
nor U2416 (N_2416,N_1958,N_1823);
nand U2417 (N_2417,N_2112,N_1997);
xnor U2418 (N_2418,N_2277,N_1896);
nand U2419 (N_2419,N_2040,N_2145);
nor U2420 (N_2420,N_1810,N_2107);
nor U2421 (N_2421,N_1816,N_2353);
or U2422 (N_2422,N_1874,N_2229);
nor U2423 (N_2423,N_2319,N_2344);
nand U2424 (N_2424,N_1939,N_2204);
or U2425 (N_2425,N_1809,N_2008);
xnor U2426 (N_2426,N_1802,N_2031);
nand U2427 (N_2427,N_1933,N_2148);
nand U2428 (N_2428,N_2037,N_2222);
and U2429 (N_2429,N_1967,N_2178);
nor U2430 (N_2430,N_1994,N_2210);
nor U2431 (N_2431,N_2216,N_2390);
and U2432 (N_2432,N_2202,N_2200);
or U2433 (N_2433,N_1808,N_2323);
xor U2434 (N_2434,N_1860,N_2170);
and U2435 (N_2435,N_1969,N_1936);
nand U2436 (N_2436,N_2386,N_1906);
and U2437 (N_2437,N_1948,N_2093);
nor U2438 (N_2438,N_1996,N_1966);
or U2439 (N_2439,N_2127,N_2026);
and U2440 (N_2440,N_2317,N_1842);
nor U2441 (N_2441,N_2381,N_2298);
or U2442 (N_2442,N_2044,N_2370);
and U2443 (N_2443,N_1991,N_2023);
nor U2444 (N_2444,N_1905,N_2343);
nand U2445 (N_2445,N_2183,N_1947);
nand U2446 (N_2446,N_2191,N_1854);
nand U2447 (N_2447,N_2376,N_2198);
or U2448 (N_2448,N_2030,N_2062);
and U2449 (N_2449,N_1856,N_2083);
nand U2450 (N_2450,N_1981,N_2258);
nor U2451 (N_2451,N_2077,N_2243);
nor U2452 (N_2452,N_2086,N_2399);
nor U2453 (N_2453,N_1899,N_2297);
nand U2454 (N_2454,N_1927,N_1822);
and U2455 (N_2455,N_2041,N_2288);
nand U2456 (N_2456,N_1878,N_1945);
and U2457 (N_2457,N_1919,N_1862);
nor U2458 (N_2458,N_1889,N_1903);
or U2459 (N_2459,N_2331,N_2306);
nor U2460 (N_2460,N_2096,N_2071);
nand U2461 (N_2461,N_2007,N_1852);
and U2462 (N_2462,N_1864,N_2117);
or U2463 (N_2463,N_1880,N_2133);
or U2464 (N_2464,N_1916,N_1908);
nor U2465 (N_2465,N_2289,N_2389);
nand U2466 (N_2466,N_1817,N_2366);
nor U2467 (N_2467,N_2028,N_1872);
or U2468 (N_2468,N_2113,N_2034);
or U2469 (N_2469,N_1940,N_2168);
nor U2470 (N_2470,N_1891,N_2371);
nor U2471 (N_2471,N_2315,N_2347);
and U2472 (N_2472,N_2035,N_2162);
and U2473 (N_2473,N_2150,N_1941);
nor U2474 (N_2474,N_2260,N_2305);
nand U2475 (N_2475,N_2257,N_1885);
nor U2476 (N_2476,N_2039,N_2348);
nand U2477 (N_2477,N_2249,N_2064);
and U2478 (N_2478,N_2088,N_2182);
nand U2479 (N_2479,N_2055,N_1847);
nor U2480 (N_2480,N_1932,N_2397);
or U2481 (N_2481,N_2380,N_1866);
nand U2482 (N_2482,N_1875,N_2002);
nand U2483 (N_2483,N_1974,N_2017);
and U2484 (N_2484,N_2094,N_2130);
nor U2485 (N_2485,N_2215,N_2301);
nor U2486 (N_2486,N_2074,N_2203);
or U2487 (N_2487,N_2393,N_2066);
or U2488 (N_2488,N_1938,N_2291);
nor U2489 (N_2489,N_2372,N_1826);
nor U2490 (N_2490,N_2223,N_2383);
or U2491 (N_2491,N_2122,N_2010);
and U2492 (N_2492,N_2327,N_1887);
nor U2493 (N_2493,N_1870,N_1993);
and U2494 (N_2494,N_2139,N_1848);
nand U2495 (N_2495,N_1931,N_1883);
nand U2496 (N_2496,N_2085,N_1935);
nor U2497 (N_2497,N_2213,N_1984);
or U2498 (N_2498,N_2226,N_2299);
or U2499 (N_2499,N_2254,N_1979);
or U2500 (N_2500,N_2274,N_1950);
nand U2501 (N_2501,N_2019,N_2328);
and U2502 (N_2502,N_2285,N_2194);
nor U2503 (N_2503,N_2188,N_2240);
and U2504 (N_2504,N_2280,N_2212);
or U2505 (N_2505,N_1913,N_2067);
or U2506 (N_2506,N_2185,N_1825);
nand U2507 (N_2507,N_1934,N_2310);
nand U2508 (N_2508,N_1912,N_1946);
or U2509 (N_2509,N_1815,N_2244);
and U2510 (N_2510,N_2321,N_2275);
and U2511 (N_2511,N_2192,N_2284);
and U2512 (N_2512,N_2043,N_2070);
and U2513 (N_2513,N_2164,N_2346);
nor U2514 (N_2514,N_2264,N_1929);
or U2515 (N_2515,N_2334,N_2167);
nor U2516 (N_2516,N_1973,N_2325);
or U2517 (N_2517,N_2174,N_2106);
or U2518 (N_2518,N_2209,N_2032);
and U2519 (N_2519,N_2109,N_1800);
or U2520 (N_2520,N_1845,N_1917);
nor U2521 (N_2521,N_2314,N_1962);
or U2522 (N_2522,N_1869,N_1944);
xnor U2523 (N_2523,N_2022,N_2263);
xor U2524 (N_2524,N_1855,N_2313);
nand U2525 (N_2525,N_2024,N_1836);
nor U2526 (N_2526,N_2340,N_1890);
nand U2527 (N_2527,N_2193,N_1858);
and U2528 (N_2528,N_2270,N_2214);
and U2529 (N_2529,N_2155,N_2369);
nor U2530 (N_2530,N_1999,N_2387);
nand U2531 (N_2531,N_2360,N_1957);
nand U2532 (N_2532,N_2058,N_2232);
nand U2533 (N_2533,N_1814,N_1915);
nor U2534 (N_2534,N_1820,N_2281);
nor U2535 (N_2535,N_1923,N_2330);
or U2536 (N_2536,N_2042,N_2336);
nand U2537 (N_2537,N_1884,N_2033);
nand U2538 (N_2538,N_2116,N_2374);
nand U2539 (N_2539,N_2175,N_1955);
nand U2540 (N_2540,N_2054,N_2069);
and U2541 (N_2541,N_2092,N_2341);
and U2542 (N_2542,N_2292,N_2025);
nand U2543 (N_2543,N_1983,N_1942);
and U2544 (N_2544,N_1961,N_1871);
or U2545 (N_2545,N_1926,N_2300);
nand U2546 (N_2546,N_2337,N_2159);
xnor U2547 (N_2547,N_2250,N_2283);
nand U2548 (N_2548,N_1907,N_2247);
nand U2549 (N_2549,N_2256,N_1951);
nor U2550 (N_2550,N_1978,N_2108);
nor U2551 (N_2551,N_2158,N_1995);
nor U2552 (N_2552,N_1949,N_2181);
or U2553 (N_2553,N_2267,N_2259);
xor U2554 (N_2554,N_1894,N_2161);
and U2555 (N_2555,N_2377,N_2396);
nor U2556 (N_2556,N_2004,N_1975);
and U2557 (N_2557,N_2166,N_2190);
and U2558 (N_2558,N_1834,N_2103);
or U2559 (N_2559,N_1818,N_2378);
or U2560 (N_2560,N_2047,N_2208);
xnor U2561 (N_2561,N_2349,N_2189);
or U2562 (N_2562,N_2266,N_2234);
or U2563 (N_2563,N_2302,N_2278);
nand U2564 (N_2564,N_2339,N_2012);
nor U2565 (N_2565,N_2335,N_1861);
xnor U2566 (N_2566,N_2036,N_2157);
or U2567 (N_2567,N_1857,N_2354);
nand U2568 (N_2568,N_2398,N_1930);
or U2569 (N_2569,N_1803,N_2027);
and U2570 (N_2570,N_2011,N_1843);
nor U2571 (N_2571,N_2255,N_1897);
nand U2572 (N_2572,N_1819,N_2163);
xnor U2573 (N_2573,N_2051,N_2152);
nand U2574 (N_2574,N_2241,N_1965);
nand U2575 (N_2575,N_2049,N_2143);
and U2576 (N_2576,N_2079,N_1849);
nor U2577 (N_2577,N_2014,N_2217);
or U2578 (N_2578,N_2087,N_1928);
or U2579 (N_2579,N_2197,N_2138);
and U2580 (N_2580,N_2015,N_1990);
nor U2581 (N_2581,N_1838,N_2221);
and U2582 (N_2582,N_1918,N_1953);
and U2583 (N_2583,N_2020,N_2097);
nand U2584 (N_2584,N_1877,N_2123);
xor U2585 (N_2585,N_2385,N_2172);
and U2586 (N_2586,N_2059,N_2149);
or U2587 (N_2587,N_1922,N_2076);
or U2588 (N_2588,N_1964,N_2307);
or U2589 (N_2589,N_2373,N_1886);
or U2590 (N_2590,N_2224,N_1960);
and U2591 (N_2591,N_2338,N_2290);
nor U2592 (N_2592,N_1971,N_1977);
nand U2593 (N_2593,N_2053,N_2359);
or U2594 (N_2594,N_2351,N_2173);
xor U2595 (N_2595,N_2072,N_2375);
nand U2596 (N_2596,N_2352,N_2246);
and U2597 (N_2597,N_1876,N_2364);
and U2598 (N_2598,N_2095,N_2356);
or U2599 (N_2599,N_2388,N_2345);
nor U2600 (N_2600,N_2147,N_2272);
or U2601 (N_2601,N_2239,N_2361);
and U2602 (N_2602,N_2156,N_2233);
xor U2603 (N_2603,N_2251,N_2081);
nor U2604 (N_2604,N_2365,N_1972);
or U2605 (N_2605,N_2237,N_2084);
nand U2606 (N_2606,N_2395,N_1956);
nand U2607 (N_2607,N_1910,N_1925);
xor U2608 (N_2608,N_2052,N_1853);
nand U2609 (N_2609,N_2211,N_1812);
and U2610 (N_2610,N_2114,N_1959);
and U2611 (N_2611,N_2392,N_1873);
nand U2612 (N_2612,N_2279,N_1943);
nor U2613 (N_2613,N_2218,N_2220);
nand U2614 (N_2614,N_1846,N_1811);
xnor U2615 (N_2615,N_1988,N_2179);
and U2616 (N_2616,N_2187,N_2367);
and U2617 (N_2617,N_1980,N_1888);
nand U2618 (N_2618,N_1801,N_2065);
nand U2619 (N_2619,N_2132,N_2286);
or U2620 (N_2620,N_1882,N_1892);
nor U2621 (N_2621,N_2134,N_1833);
xnor U2622 (N_2622,N_1813,N_2089);
nor U2623 (N_2623,N_2080,N_1850);
and U2624 (N_2624,N_1841,N_2018);
nor U2625 (N_2625,N_2180,N_2357);
nor U2626 (N_2626,N_2391,N_2046);
and U2627 (N_2627,N_1881,N_2332);
xor U2628 (N_2628,N_2236,N_2075);
nor U2629 (N_2629,N_1868,N_2329);
or U2630 (N_2630,N_2006,N_2120);
nor U2631 (N_2631,N_2228,N_1898);
or U2632 (N_2632,N_1835,N_2063);
nor U2633 (N_2633,N_2003,N_2219);
nor U2634 (N_2634,N_2005,N_2362);
nand U2635 (N_2635,N_1829,N_2358);
nand U2636 (N_2636,N_1828,N_1987);
xnor U2637 (N_2637,N_2296,N_1901);
nor U2638 (N_2638,N_1821,N_2021);
nand U2639 (N_2639,N_2196,N_2142);
nand U2640 (N_2640,N_2269,N_2057);
nand U2641 (N_2641,N_2154,N_2102);
nor U2642 (N_2642,N_1807,N_2082);
or U2643 (N_2643,N_2252,N_1879);
or U2644 (N_2644,N_1986,N_2311);
nand U2645 (N_2645,N_2098,N_2110);
nor U2646 (N_2646,N_1830,N_1839);
nand U2647 (N_2647,N_2333,N_2128);
nand U2648 (N_2648,N_2276,N_2144);
nor U2649 (N_2649,N_2304,N_2227);
nand U2650 (N_2650,N_2061,N_2293);
or U2651 (N_2651,N_1985,N_1844);
and U2652 (N_2652,N_1865,N_2121);
and U2653 (N_2653,N_2184,N_1859);
nor U2654 (N_2654,N_2029,N_2151);
nor U2655 (N_2655,N_2363,N_2105);
nand U2656 (N_2656,N_2146,N_2160);
or U2657 (N_2657,N_1863,N_1963);
and U2658 (N_2658,N_2394,N_2273);
and U2659 (N_2659,N_2245,N_2000);
or U2660 (N_2660,N_1924,N_2355);
nand U2661 (N_2661,N_2137,N_2207);
or U2662 (N_2662,N_1805,N_2141);
nand U2663 (N_2663,N_1824,N_1909);
nand U2664 (N_2664,N_2090,N_1900);
and U2665 (N_2665,N_2368,N_2115);
nor U2666 (N_2666,N_2099,N_2016);
or U2667 (N_2667,N_2342,N_2124);
nor U2668 (N_2668,N_1968,N_2268);
nand U2669 (N_2669,N_2242,N_2165);
and U2670 (N_2670,N_1921,N_1895);
nand U2671 (N_2671,N_1989,N_1893);
xor U2672 (N_2672,N_1827,N_2253);
nor U2673 (N_2673,N_1976,N_2261);
nand U2674 (N_2674,N_2136,N_2262);
and U2675 (N_2675,N_1831,N_2238);
or U2676 (N_2676,N_2013,N_2295);
nand U2677 (N_2677,N_1837,N_2230);
xnor U2678 (N_2678,N_2153,N_2038);
xor U2679 (N_2679,N_2350,N_2199);
and U2680 (N_2680,N_2231,N_2009);
nor U2681 (N_2681,N_2271,N_2078);
nand U2682 (N_2682,N_1998,N_1902);
nand U2683 (N_2683,N_2318,N_2056);
nand U2684 (N_2684,N_2073,N_2050);
nor U2685 (N_2685,N_2129,N_2100);
xor U2686 (N_2686,N_2101,N_2001);
or U2687 (N_2687,N_2131,N_1911);
nor U2688 (N_2688,N_1952,N_2320);
or U2689 (N_2689,N_2316,N_1904);
or U2690 (N_2690,N_2060,N_2140);
nor U2691 (N_2691,N_2206,N_1804);
nand U2692 (N_2692,N_1982,N_2104);
and U2693 (N_2693,N_2169,N_2309);
nand U2694 (N_2694,N_2201,N_2111);
or U2695 (N_2695,N_2186,N_1970);
nand U2696 (N_2696,N_2324,N_2225);
and U2697 (N_2697,N_2248,N_2205);
nor U2698 (N_2698,N_2235,N_1914);
and U2699 (N_2699,N_2171,N_1832);
and U2700 (N_2700,N_1990,N_1964);
and U2701 (N_2701,N_2369,N_2208);
nand U2702 (N_2702,N_1982,N_2059);
nor U2703 (N_2703,N_2316,N_1879);
xnor U2704 (N_2704,N_2287,N_1881);
and U2705 (N_2705,N_2237,N_2101);
or U2706 (N_2706,N_2143,N_2053);
or U2707 (N_2707,N_2376,N_1805);
nand U2708 (N_2708,N_2138,N_2079);
nand U2709 (N_2709,N_2327,N_2294);
or U2710 (N_2710,N_1832,N_1819);
nand U2711 (N_2711,N_2027,N_1835);
xor U2712 (N_2712,N_2168,N_2319);
xnor U2713 (N_2713,N_2155,N_2105);
xnor U2714 (N_2714,N_2282,N_2069);
nand U2715 (N_2715,N_2189,N_1885);
or U2716 (N_2716,N_2270,N_2021);
or U2717 (N_2717,N_1810,N_1871);
or U2718 (N_2718,N_1899,N_2132);
and U2719 (N_2719,N_1953,N_2026);
nor U2720 (N_2720,N_1967,N_2053);
and U2721 (N_2721,N_2281,N_2120);
and U2722 (N_2722,N_2275,N_2165);
and U2723 (N_2723,N_1823,N_2281);
nor U2724 (N_2724,N_2069,N_2016);
nor U2725 (N_2725,N_2145,N_2155);
xnor U2726 (N_2726,N_2187,N_2123);
xnor U2727 (N_2727,N_2097,N_2393);
and U2728 (N_2728,N_1974,N_2277);
nand U2729 (N_2729,N_2381,N_1989);
or U2730 (N_2730,N_2224,N_2163);
and U2731 (N_2731,N_1962,N_1939);
and U2732 (N_2732,N_2168,N_1891);
xor U2733 (N_2733,N_2090,N_2101);
xnor U2734 (N_2734,N_2257,N_2049);
nand U2735 (N_2735,N_2354,N_2085);
or U2736 (N_2736,N_2377,N_1818);
and U2737 (N_2737,N_1999,N_1803);
or U2738 (N_2738,N_2149,N_2026);
nand U2739 (N_2739,N_2338,N_2061);
nand U2740 (N_2740,N_2265,N_2241);
and U2741 (N_2741,N_2193,N_2108);
or U2742 (N_2742,N_2072,N_2116);
and U2743 (N_2743,N_2348,N_1942);
nor U2744 (N_2744,N_2146,N_2282);
xnor U2745 (N_2745,N_2203,N_1894);
nor U2746 (N_2746,N_1882,N_2373);
or U2747 (N_2747,N_1945,N_2288);
nor U2748 (N_2748,N_1959,N_1936);
or U2749 (N_2749,N_2150,N_2045);
or U2750 (N_2750,N_2067,N_2058);
or U2751 (N_2751,N_2314,N_2389);
and U2752 (N_2752,N_2155,N_2374);
and U2753 (N_2753,N_2326,N_2214);
nor U2754 (N_2754,N_2284,N_2133);
and U2755 (N_2755,N_1991,N_2079);
or U2756 (N_2756,N_2333,N_2284);
nand U2757 (N_2757,N_2111,N_2124);
nor U2758 (N_2758,N_1844,N_2281);
and U2759 (N_2759,N_2036,N_1972);
nand U2760 (N_2760,N_2083,N_1843);
nor U2761 (N_2761,N_1946,N_1899);
nor U2762 (N_2762,N_1983,N_2043);
nor U2763 (N_2763,N_1933,N_1960);
nor U2764 (N_2764,N_2240,N_2017);
nor U2765 (N_2765,N_1802,N_1975);
nor U2766 (N_2766,N_2361,N_1968);
and U2767 (N_2767,N_1884,N_2101);
nand U2768 (N_2768,N_2215,N_2230);
nor U2769 (N_2769,N_1841,N_2213);
or U2770 (N_2770,N_2377,N_1897);
nor U2771 (N_2771,N_2322,N_2282);
and U2772 (N_2772,N_1864,N_2354);
and U2773 (N_2773,N_1920,N_2311);
or U2774 (N_2774,N_2294,N_2045);
xor U2775 (N_2775,N_2248,N_2374);
nor U2776 (N_2776,N_1854,N_2192);
xnor U2777 (N_2777,N_2276,N_2380);
or U2778 (N_2778,N_2376,N_1912);
nor U2779 (N_2779,N_2056,N_2007);
nand U2780 (N_2780,N_2141,N_1829);
nand U2781 (N_2781,N_1985,N_1907);
or U2782 (N_2782,N_1873,N_2359);
or U2783 (N_2783,N_2191,N_1881);
xnor U2784 (N_2784,N_2011,N_2022);
or U2785 (N_2785,N_2290,N_2057);
nor U2786 (N_2786,N_1900,N_2307);
or U2787 (N_2787,N_1971,N_1880);
and U2788 (N_2788,N_1946,N_2105);
nand U2789 (N_2789,N_2027,N_1881);
and U2790 (N_2790,N_2015,N_2266);
or U2791 (N_2791,N_2010,N_1838);
xnor U2792 (N_2792,N_2152,N_2102);
and U2793 (N_2793,N_2277,N_1967);
or U2794 (N_2794,N_2060,N_2216);
xnor U2795 (N_2795,N_1804,N_2329);
nand U2796 (N_2796,N_1848,N_2294);
xor U2797 (N_2797,N_2124,N_1851);
and U2798 (N_2798,N_2059,N_2111);
nor U2799 (N_2799,N_2149,N_2250);
or U2800 (N_2800,N_2231,N_2179);
xor U2801 (N_2801,N_2373,N_1906);
xnor U2802 (N_2802,N_2060,N_1993);
xor U2803 (N_2803,N_1945,N_2207);
and U2804 (N_2804,N_2298,N_2377);
nand U2805 (N_2805,N_2262,N_2377);
nor U2806 (N_2806,N_1867,N_2179);
nor U2807 (N_2807,N_1881,N_2136);
and U2808 (N_2808,N_2170,N_2209);
nor U2809 (N_2809,N_1978,N_1800);
or U2810 (N_2810,N_2285,N_2385);
and U2811 (N_2811,N_1922,N_2279);
and U2812 (N_2812,N_1945,N_2054);
xor U2813 (N_2813,N_2320,N_2103);
or U2814 (N_2814,N_1905,N_2018);
nand U2815 (N_2815,N_1803,N_1934);
or U2816 (N_2816,N_1976,N_2337);
xor U2817 (N_2817,N_2040,N_1804);
or U2818 (N_2818,N_1849,N_2147);
nor U2819 (N_2819,N_1867,N_2306);
nand U2820 (N_2820,N_1940,N_2338);
xor U2821 (N_2821,N_1973,N_2120);
nand U2822 (N_2822,N_2299,N_2088);
or U2823 (N_2823,N_2017,N_2119);
and U2824 (N_2824,N_2165,N_2348);
nand U2825 (N_2825,N_2256,N_2344);
nor U2826 (N_2826,N_2211,N_2255);
nor U2827 (N_2827,N_1946,N_2193);
xnor U2828 (N_2828,N_1983,N_1934);
nand U2829 (N_2829,N_2197,N_2309);
nand U2830 (N_2830,N_2183,N_1962);
or U2831 (N_2831,N_2193,N_2137);
nor U2832 (N_2832,N_1980,N_2139);
nor U2833 (N_2833,N_2289,N_2177);
nor U2834 (N_2834,N_2287,N_1884);
or U2835 (N_2835,N_2055,N_2204);
nor U2836 (N_2836,N_2119,N_2171);
nand U2837 (N_2837,N_2307,N_2209);
nor U2838 (N_2838,N_2308,N_1887);
nand U2839 (N_2839,N_1853,N_2363);
or U2840 (N_2840,N_2211,N_1843);
nor U2841 (N_2841,N_2023,N_2082);
nand U2842 (N_2842,N_2374,N_2327);
and U2843 (N_2843,N_1836,N_1818);
or U2844 (N_2844,N_2082,N_1861);
nor U2845 (N_2845,N_2335,N_1933);
xor U2846 (N_2846,N_1909,N_1852);
nand U2847 (N_2847,N_2163,N_2046);
nor U2848 (N_2848,N_2344,N_2025);
nor U2849 (N_2849,N_1923,N_2327);
or U2850 (N_2850,N_2374,N_2135);
nor U2851 (N_2851,N_1815,N_2269);
and U2852 (N_2852,N_2371,N_2097);
nand U2853 (N_2853,N_1825,N_2371);
nand U2854 (N_2854,N_2115,N_2032);
nand U2855 (N_2855,N_2167,N_2149);
and U2856 (N_2856,N_2338,N_2250);
xor U2857 (N_2857,N_2332,N_2386);
xor U2858 (N_2858,N_2398,N_2112);
and U2859 (N_2859,N_1846,N_2257);
or U2860 (N_2860,N_2306,N_2360);
or U2861 (N_2861,N_2070,N_1955);
nand U2862 (N_2862,N_1915,N_1914);
and U2863 (N_2863,N_1875,N_1992);
or U2864 (N_2864,N_1812,N_1975);
or U2865 (N_2865,N_1991,N_1911);
nor U2866 (N_2866,N_1843,N_2297);
or U2867 (N_2867,N_2043,N_1996);
nor U2868 (N_2868,N_1990,N_2275);
nor U2869 (N_2869,N_1870,N_1895);
or U2870 (N_2870,N_2174,N_1942);
and U2871 (N_2871,N_1954,N_2300);
nand U2872 (N_2872,N_2091,N_1820);
or U2873 (N_2873,N_1830,N_2209);
nand U2874 (N_2874,N_1998,N_1841);
nand U2875 (N_2875,N_1944,N_1918);
nor U2876 (N_2876,N_1878,N_2113);
nor U2877 (N_2877,N_1846,N_2147);
or U2878 (N_2878,N_2052,N_2129);
or U2879 (N_2879,N_2091,N_2283);
nor U2880 (N_2880,N_1857,N_1834);
nor U2881 (N_2881,N_2088,N_2257);
and U2882 (N_2882,N_2247,N_1924);
nand U2883 (N_2883,N_1836,N_2014);
nand U2884 (N_2884,N_1946,N_2259);
and U2885 (N_2885,N_2215,N_2201);
or U2886 (N_2886,N_2051,N_2352);
xor U2887 (N_2887,N_1832,N_2114);
xnor U2888 (N_2888,N_2098,N_2050);
xnor U2889 (N_2889,N_2305,N_2059);
nor U2890 (N_2890,N_2280,N_1876);
xor U2891 (N_2891,N_1992,N_2384);
and U2892 (N_2892,N_2202,N_2007);
or U2893 (N_2893,N_2160,N_2343);
xnor U2894 (N_2894,N_1895,N_2375);
xnor U2895 (N_2895,N_2386,N_1880);
and U2896 (N_2896,N_2188,N_1969);
and U2897 (N_2897,N_2035,N_1958);
nor U2898 (N_2898,N_2099,N_2086);
or U2899 (N_2899,N_2207,N_2162);
nand U2900 (N_2900,N_2337,N_2142);
and U2901 (N_2901,N_2082,N_1965);
nand U2902 (N_2902,N_2142,N_2303);
or U2903 (N_2903,N_2367,N_2053);
and U2904 (N_2904,N_2016,N_2236);
nand U2905 (N_2905,N_1908,N_2232);
nand U2906 (N_2906,N_2091,N_2208);
xnor U2907 (N_2907,N_2182,N_2275);
nand U2908 (N_2908,N_2187,N_2183);
nand U2909 (N_2909,N_2102,N_1845);
xor U2910 (N_2910,N_2194,N_2281);
and U2911 (N_2911,N_1822,N_1964);
nor U2912 (N_2912,N_1968,N_1813);
or U2913 (N_2913,N_2159,N_1882);
or U2914 (N_2914,N_2178,N_2020);
nor U2915 (N_2915,N_1941,N_2395);
xor U2916 (N_2916,N_2244,N_2286);
nor U2917 (N_2917,N_2060,N_1964);
and U2918 (N_2918,N_2316,N_2261);
nand U2919 (N_2919,N_2249,N_1880);
or U2920 (N_2920,N_1870,N_1821);
or U2921 (N_2921,N_2387,N_2214);
and U2922 (N_2922,N_2299,N_2177);
and U2923 (N_2923,N_2153,N_2170);
nor U2924 (N_2924,N_1976,N_2176);
and U2925 (N_2925,N_1808,N_2263);
and U2926 (N_2926,N_2040,N_1829);
xnor U2927 (N_2927,N_2031,N_2280);
nor U2928 (N_2928,N_2293,N_2391);
nand U2929 (N_2929,N_2134,N_2244);
and U2930 (N_2930,N_1896,N_1923);
or U2931 (N_2931,N_2256,N_2234);
or U2932 (N_2932,N_2331,N_2179);
or U2933 (N_2933,N_1966,N_2248);
nor U2934 (N_2934,N_2289,N_2384);
nand U2935 (N_2935,N_2360,N_2004);
nor U2936 (N_2936,N_1824,N_2336);
nand U2937 (N_2937,N_2239,N_1952);
or U2938 (N_2938,N_2058,N_2263);
nand U2939 (N_2939,N_2081,N_1952);
nor U2940 (N_2940,N_1853,N_2381);
or U2941 (N_2941,N_2350,N_2316);
or U2942 (N_2942,N_2383,N_2046);
and U2943 (N_2943,N_2085,N_1966);
and U2944 (N_2944,N_2168,N_2064);
nor U2945 (N_2945,N_2204,N_1843);
and U2946 (N_2946,N_2283,N_2062);
nor U2947 (N_2947,N_2133,N_2264);
nor U2948 (N_2948,N_2075,N_2014);
or U2949 (N_2949,N_2047,N_2325);
nor U2950 (N_2950,N_2236,N_2277);
nor U2951 (N_2951,N_2354,N_2333);
nor U2952 (N_2952,N_2119,N_2148);
nor U2953 (N_2953,N_2285,N_2221);
nor U2954 (N_2954,N_2268,N_2208);
nor U2955 (N_2955,N_2105,N_1815);
or U2956 (N_2956,N_2385,N_1848);
xor U2957 (N_2957,N_1919,N_2035);
nand U2958 (N_2958,N_2330,N_2363);
and U2959 (N_2959,N_1883,N_1909);
nand U2960 (N_2960,N_2279,N_1999);
or U2961 (N_2961,N_2043,N_1805);
nor U2962 (N_2962,N_2129,N_2155);
nor U2963 (N_2963,N_2206,N_2391);
or U2964 (N_2964,N_2174,N_1953);
nor U2965 (N_2965,N_2361,N_2010);
or U2966 (N_2966,N_2189,N_2145);
and U2967 (N_2967,N_1979,N_2184);
nand U2968 (N_2968,N_1855,N_2161);
xor U2969 (N_2969,N_2031,N_2365);
and U2970 (N_2970,N_2187,N_1840);
or U2971 (N_2971,N_1930,N_2160);
and U2972 (N_2972,N_1875,N_1920);
nand U2973 (N_2973,N_2357,N_1905);
nand U2974 (N_2974,N_2252,N_1978);
and U2975 (N_2975,N_2027,N_2282);
nor U2976 (N_2976,N_2161,N_2196);
or U2977 (N_2977,N_2374,N_1919);
nor U2978 (N_2978,N_2011,N_2134);
nand U2979 (N_2979,N_2208,N_2087);
nor U2980 (N_2980,N_1837,N_2127);
nor U2981 (N_2981,N_1968,N_1884);
nor U2982 (N_2982,N_2172,N_2241);
or U2983 (N_2983,N_1850,N_2174);
nand U2984 (N_2984,N_2215,N_1841);
or U2985 (N_2985,N_2385,N_2333);
nand U2986 (N_2986,N_1931,N_1949);
or U2987 (N_2987,N_2288,N_2191);
nand U2988 (N_2988,N_2220,N_1837);
nor U2989 (N_2989,N_2083,N_1928);
nand U2990 (N_2990,N_1928,N_2306);
and U2991 (N_2991,N_2329,N_1875);
and U2992 (N_2992,N_2352,N_2062);
nor U2993 (N_2993,N_2379,N_2010);
or U2994 (N_2994,N_2390,N_1885);
and U2995 (N_2995,N_2076,N_2099);
nor U2996 (N_2996,N_1911,N_2198);
or U2997 (N_2997,N_2124,N_2139);
nor U2998 (N_2998,N_2068,N_2271);
nand U2999 (N_2999,N_2118,N_2167);
and UO_0 (O_0,N_2768,N_2810);
or UO_1 (O_1,N_2727,N_2912);
or UO_2 (O_2,N_2494,N_2421);
or UO_3 (O_3,N_2908,N_2485);
and UO_4 (O_4,N_2698,N_2693);
nand UO_5 (O_5,N_2794,N_2612);
or UO_6 (O_6,N_2564,N_2888);
or UO_7 (O_7,N_2547,N_2932);
or UO_8 (O_8,N_2500,N_2817);
or UO_9 (O_9,N_2882,N_2968);
and UO_10 (O_10,N_2903,N_2654);
xor UO_11 (O_11,N_2592,N_2925);
and UO_12 (O_12,N_2789,N_2900);
and UO_13 (O_13,N_2501,N_2934);
and UO_14 (O_14,N_2548,N_2420);
and UO_15 (O_15,N_2668,N_2555);
or UO_16 (O_16,N_2844,N_2438);
nor UO_17 (O_17,N_2468,N_2920);
nand UO_18 (O_18,N_2804,N_2590);
nand UO_19 (O_19,N_2510,N_2955);
nand UO_20 (O_20,N_2446,N_2574);
or UO_21 (O_21,N_2954,N_2672);
or UO_22 (O_22,N_2509,N_2976);
nor UO_23 (O_23,N_2694,N_2476);
or UO_24 (O_24,N_2498,N_2695);
xnor UO_25 (O_25,N_2481,N_2589);
and UO_26 (O_26,N_2608,N_2958);
nand UO_27 (O_27,N_2667,N_2401);
nor UO_28 (O_28,N_2400,N_2851);
or UO_29 (O_29,N_2896,N_2975);
nand UO_30 (O_30,N_2866,N_2665);
or UO_31 (O_31,N_2834,N_2701);
and UO_32 (O_32,N_2803,N_2953);
and UO_33 (O_33,N_2906,N_2785);
nand UO_34 (O_34,N_2514,N_2604);
xnor UO_35 (O_35,N_2824,N_2875);
xnor UO_36 (O_36,N_2515,N_2483);
nand UO_37 (O_37,N_2477,N_2594);
nor UO_38 (O_38,N_2772,N_2842);
nor UO_39 (O_39,N_2940,N_2791);
and UO_40 (O_40,N_2562,N_2725);
xnor UO_41 (O_41,N_2947,N_2827);
nand UO_42 (O_42,N_2542,N_2459);
nand UO_43 (O_43,N_2469,N_2605);
xnor UO_44 (O_44,N_2664,N_2448);
nand UO_45 (O_45,N_2796,N_2613);
nand UO_46 (O_46,N_2713,N_2656);
nand UO_47 (O_47,N_2849,N_2990);
nand UO_48 (O_48,N_2653,N_2433);
and UO_49 (O_49,N_2516,N_2557);
or UO_50 (O_50,N_2885,N_2543);
nand UO_51 (O_51,N_2938,N_2811);
and UO_52 (O_52,N_2951,N_2863);
nand UO_53 (O_53,N_2445,N_2864);
nand UO_54 (O_54,N_2933,N_2795);
xor UO_55 (O_55,N_2845,N_2606);
xor UO_56 (O_56,N_2731,N_2591);
and UO_57 (O_57,N_2862,N_2859);
and UO_58 (O_58,N_2751,N_2745);
nand UO_59 (O_59,N_2648,N_2831);
nor UO_60 (O_60,N_2490,N_2950);
or UO_61 (O_61,N_2887,N_2684);
nand UO_62 (O_62,N_2517,N_2764);
or UO_63 (O_63,N_2716,N_2414);
and UO_64 (O_64,N_2561,N_2629);
or UO_65 (O_65,N_2584,N_2992);
nor UO_66 (O_66,N_2460,N_2743);
and UO_67 (O_67,N_2999,N_2416);
nor UO_68 (O_68,N_2923,N_2914);
or UO_69 (O_69,N_2565,N_2602);
and UO_70 (O_70,N_2634,N_2986);
and UO_71 (O_71,N_2610,N_2626);
xnor UO_72 (O_72,N_2723,N_2722);
or UO_73 (O_73,N_2640,N_2823);
and UO_74 (O_74,N_2867,N_2969);
nor UO_75 (O_75,N_2440,N_2441);
nand UO_76 (O_76,N_2746,N_2773);
nand UO_77 (O_77,N_2541,N_2577);
nand UO_78 (O_78,N_2686,N_2627);
or UO_79 (O_79,N_2778,N_2918);
and UO_80 (O_80,N_2550,N_2675);
nor UO_81 (O_81,N_2639,N_2611);
nand UO_82 (O_82,N_2585,N_2961);
xor UO_83 (O_83,N_2669,N_2871);
nor UO_84 (O_84,N_2457,N_2595);
nor UO_85 (O_85,N_2527,N_2995);
and UO_86 (O_86,N_2536,N_2878);
nand UO_87 (O_87,N_2832,N_2637);
xor UO_88 (O_88,N_2787,N_2600);
or UO_89 (O_89,N_2593,N_2818);
nand UO_90 (O_90,N_2521,N_2666);
xor UO_91 (O_91,N_2971,N_2911);
xnor UO_92 (O_92,N_2784,N_2852);
xor UO_93 (O_93,N_2437,N_2736);
nand UO_94 (O_94,N_2869,N_2544);
and UO_95 (O_95,N_2614,N_2905);
and UO_96 (O_96,N_2588,N_2926);
and UO_97 (O_97,N_2616,N_2569);
and UO_98 (O_98,N_2529,N_2688);
nor UO_99 (O_99,N_2431,N_2525);
nand UO_100 (O_100,N_2843,N_2705);
or UO_101 (O_101,N_2609,N_2426);
nor UO_102 (O_102,N_2805,N_2897);
or UO_103 (O_103,N_2537,N_2775);
or UO_104 (O_104,N_2967,N_2748);
and UO_105 (O_105,N_2858,N_2812);
nor UO_106 (O_106,N_2676,N_2774);
nand UO_107 (O_107,N_2681,N_2465);
nand UO_108 (O_108,N_2597,N_2993);
nand UO_109 (O_109,N_2755,N_2724);
and UO_110 (O_110,N_2428,N_2628);
or UO_111 (O_111,N_2894,N_2939);
xor UO_112 (O_112,N_2726,N_2522);
nand UO_113 (O_113,N_2470,N_2566);
nor UO_114 (O_114,N_2671,N_2892);
nor UO_115 (O_115,N_2422,N_2449);
or UO_116 (O_116,N_2409,N_2435);
nand UO_117 (O_117,N_2580,N_2413);
and UO_118 (O_118,N_2474,N_2462);
nand UO_119 (O_119,N_2466,N_2645);
nor UO_120 (O_120,N_2982,N_2750);
xnor UO_121 (O_121,N_2677,N_2496);
nand UO_122 (O_122,N_2404,N_2799);
xnor UO_123 (O_123,N_2545,N_2499);
or UO_124 (O_124,N_2425,N_2957);
nand UO_125 (O_125,N_2988,N_2822);
nor UO_126 (O_126,N_2962,N_2747);
or UO_127 (O_127,N_2405,N_2836);
or UO_128 (O_128,N_2786,N_2567);
nand UO_129 (O_129,N_2873,N_2689);
or UO_130 (O_130,N_2769,N_2941);
nor UO_131 (O_131,N_2872,N_2857);
nor UO_132 (O_132,N_2734,N_2635);
nand UO_133 (O_133,N_2929,N_2770);
xnor UO_134 (O_134,N_2556,N_2646);
nor UO_135 (O_135,N_2807,N_2876);
or UO_136 (O_136,N_2512,N_2447);
or UO_137 (O_137,N_2919,N_2412);
nor UO_138 (O_138,N_2758,N_2994);
or UO_139 (O_139,N_2808,N_2733);
or UO_140 (O_140,N_2503,N_2793);
or UO_141 (O_141,N_2586,N_2899);
or UO_142 (O_142,N_2568,N_2402);
nand UO_143 (O_143,N_2697,N_2523);
or UO_144 (O_144,N_2410,N_2598);
and UO_145 (O_145,N_2452,N_2582);
and UO_146 (O_146,N_2717,N_2884);
nor UO_147 (O_147,N_2708,N_2835);
or UO_148 (O_148,N_2901,N_2620);
nand UO_149 (O_149,N_2489,N_2782);
and UO_150 (O_150,N_2524,N_2907);
nand UO_151 (O_151,N_2921,N_2883);
nor UO_152 (O_152,N_2909,N_2936);
or UO_153 (O_153,N_2998,N_2703);
or UO_154 (O_154,N_2777,N_2828);
or UO_155 (O_155,N_2484,N_2513);
nand UO_156 (O_156,N_2752,N_2649);
or UO_157 (O_157,N_2575,N_2935);
and UO_158 (O_158,N_2572,N_2554);
xor UO_159 (O_159,N_2493,N_2928);
nor UO_160 (O_160,N_2607,N_2407);
nand UO_161 (O_161,N_2624,N_2757);
or UO_162 (O_162,N_2690,N_2739);
or UO_163 (O_163,N_2816,N_2488);
and UO_164 (O_164,N_2644,N_2948);
or UO_165 (O_165,N_2619,N_2809);
xor UO_166 (O_166,N_2943,N_2821);
nand UO_167 (O_167,N_2815,N_2464);
nor UO_168 (O_168,N_2472,N_2622);
or UO_169 (O_169,N_2458,N_2443);
xor UO_170 (O_170,N_2406,N_2989);
xor UO_171 (O_171,N_2877,N_2519);
and UO_172 (O_172,N_2670,N_2587);
nor UO_173 (O_173,N_2531,N_2625);
or UO_174 (O_174,N_2732,N_2453);
or UO_175 (O_175,N_2487,N_2738);
or UO_176 (O_176,N_2729,N_2532);
xnor UO_177 (O_177,N_2632,N_2507);
nand UO_178 (O_178,N_2570,N_2661);
nand UO_179 (O_179,N_2418,N_2535);
xnor UO_180 (O_180,N_2802,N_2655);
nand UO_181 (O_181,N_2767,N_2898);
and UO_182 (O_182,N_2825,N_2442);
or UO_183 (O_183,N_2973,N_2800);
nor UO_184 (O_184,N_2946,N_2740);
or UO_185 (O_185,N_2779,N_2930);
or UO_186 (O_186,N_2505,N_2839);
nor UO_187 (O_187,N_2819,N_2826);
or UO_188 (O_188,N_2699,N_2492);
and UO_189 (O_189,N_2444,N_2683);
nand UO_190 (O_190,N_2652,N_2854);
or UO_191 (O_191,N_2599,N_2538);
nand UO_192 (O_192,N_2518,N_2742);
and UO_193 (O_193,N_2874,N_2855);
and UO_194 (O_194,N_2436,N_2497);
nand UO_195 (O_195,N_2636,N_2552);
or UO_196 (O_196,N_2455,N_2830);
nand UO_197 (O_197,N_2643,N_2910);
or UO_198 (O_198,N_2451,N_2571);
nand UO_199 (O_199,N_2415,N_2952);
xor UO_200 (O_200,N_2692,N_2814);
and UO_201 (O_201,N_2707,N_2848);
or UO_202 (O_202,N_2942,N_2944);
nand UO_203 (O_203,N_2980,N_2621);
and UO_204 (O_204,N_2720,N_2482);
nand UO_205 (O_205,N_2801,N_2997);
nand UO_206 (O_206,N_2633,N_2991);
and UO_207 (O_207,N_2924,N_2762);
or UO_208 (O_208,N_2850,N_2647);
nand UO_209 (O_209,N_2847,N_2853);
xnor UO_210 (O_210,N_2837,N_2479);
nor UO_211 (O_211,N_2700,N_2981);
nor UO_212 (O_212,N_2578,N_2454);
or UO_213 (O_213,N_2984,N_2623);
nand UO_214 (O_214,N_2781,N_2660);
nand UO_215 (O_215,N_2411,N_2709);
nand UO_216 (O_216,N_2965,N_2956);
nand UO_217 (O_217,N_2881,N_2949);
nand UO_218 (O_218,N_2495,N_2450);
and UO_219 (O_219,N_2706,N_2429);
nor UO_220 (O_220,N_2502,N_2783);
nand UO_221 (O_221,N_2533,N_2904);
and UO_222 (O_222,N_2662,N_2546);
nor UO_223 (O_223,N_2728,N_2673);
or UO_224 (O_224,N_2846,N_2679);
or UO_225 (O_225,N_2718,N_2797);
or UO_226 (O_226,N_2766,N_2638);
nand UO_227 (O_227,N_2576,N_2558);
nor UO_228 (O_228,N_2735,N_2868);
and UO_229 (O_229,N_2721,N_2579);
and UO_230 (O_230,N_2931,N_2719);
or UO_231 (O_231,N_2461,N_2702);
and UO_232 (O_232,N_2549,N_2715);
and UO_233 (O_233,N_2408,N_2504);
nand UO_234 (O_234,N_2687,N_2927);
and UO_235 (O_235,N_2829,N_2691);
or UO_236 (O_236,N_2419,N_2714);
or UO_237 (O_237,N_2890,N_2473);
nor UO_238 (O_238,N_2583,N_2642);
nand UO_239 (O_239,N_2663,N_2680);
and UO_240 (O_240,N_2551,N_2916);
and UO_241 (O_241,N_2870,N_2651);
nand UO_242 (O_242,N_2741,N_2761);
nand UO_243 (O_243,N_2520,N_2710);
nand UO_244 (O_244,N_2895,N_2573);
xnor UO_245 (O_245,N_2753,N_2760);
xor UO_246 (O_246,N_2749,N_2534);
and UO_247 (O_247,N_2596,N_2902);
nand UO_248 (O_248,N_2838,N_2659);
and UO_249 (O_249,N_2427,N_2430);
or UO_250 (O_250,N_2915,N_2423);
or UO_251 (O_251,N_2560,N_2630);
and UO_252 (O_252,N_2711,N_2641);
nor UO_253 (O_253,N_2985,N_2432);
and UO_254 (O_254,N_2617,N_2879);
nor UO_255 (O_255,N_2539,N_2417);
or UO_256 (O_256,N_2979,N_2553);
and UO_257 (O_257,N_2475,N_2860);
nand UO_258 (O_258,N_2581,N_2511);
and UO_259 (O_259,N_2983,N_2685);
or UO_260 (O_260,N_2917,N_2737);
or UO_261 (O_261,N_2765,N_2792);
xor UO_262 (O_262,N_2922,N_2704);
nand UO_263 (O_263,N_2780,N_2963);
or UO_264 (O_264,N_2977,N_2891);
nand UO_265 (O_265,N_2959,N_2658);
nor UO_266 (O_266,N_2486,N_2601);
nand UO_267 (O_267,N_2841,N_2913);
or UO_268 (O_268,N_2434,N_2754);
or UO_269 (O_269,N_2508,N_2674);
nand UO_270 (O_270,N_2820,N_2833);
or UO_271 (O_271,N_2526,N_2491);
or UO_272 (O_272,N_2467,N_2563);
and UO_273 (O_273,N_2856,N_2528);
and UO_274 (O_274,N_2478,N_2424);
nand UO_275 (O_275,N_2865,N_2756);
and UO_276 (O_276,N_2618,N_2945);
xnor UO_277 (O_277,N_2861,N_2650);
nand UO_278 (O_278,N_2987,N_2978);
and UO_279 (O_279,N_2776,N_2788);
and UO_280 (O_280,N_2763,N_2712);
or UO_281 (O_281,N_2759,N_2889);
and UO_282 (O_282,N_2840,N_2559);
or UO_283 (O_283,N_2972,N_2506);
and UO_284 (O_284,N_2937,N_2615);
nor UO_285 (O_285,N_2970,N_2603);
xnor UO_286 (O_286,N_2974,N_2439);
nor UO_287 (O_287,N_2813,N_2471);
nand UO_288 (O_288,N_2631,N_2678);
nand UO_289 (O_289,N_2540,N_2960);
or UO_290 (O_290,N_2964,N_2463);
nor UO_291 (O_291,N_2806,N_2744);
and UO_292 (O_292,N_2771,N_2480);
nand UO_293 (O_293,N_2886,N_2696);
or UO_294 (O_294,N_2966,N_2403);
xnor UO_295 (O_295,N_2530,N_2682);
nand UO_296 (O_296,N_2893,N_2456);
nand UO_297 (O_297,N_2790,N_2657);
or UO_298 (O_298,N_2730,N_2880);
nand UO_299 (O_299,N_2996,N_2798);
xnor UO_300 (O_300,N_2420,N_2958);
nor UO_301 (O_301,N_2664,N_2473);
nor UO_302 (O_302,N_2815,N_2918);
nand UO_303 (O_303,N_2689,N_2983);
or UO_304 (O_304,N_2684,N_2952);
nand UO_305 (O_305,N_2569,N_2824);
nor UO_306 (O_306,N_2774,N_2713);
and UO_307 (O_307,N_2573,N_2856);
and UO_308 (O_308,N_2985,N_2855);
and UO_309 (O_309,N_2981,N_2493);
and UO_310 (O_310,N_2679,N_2917);
nand UO_311 (O_311,N_2842,N_2684);
nand UO_312 (O_312,N_2617,N_2744);
nor UO_313 (O_313,N_2826,N_2999);
nor UO_314 (O_314,N_2400,N_2475);
nand UO_315 (O_315,N_2763,N_2889);
nand UO_316 (O_316,N_2504,N_2989);
nand UO_317 (O_317,N_2560,N_2406);
nor UO_318 (O_318,N_2665,N_2858);
nand UO_319 (O_319,N_2719,N_2648);
xnor UO_320 (O_320,N_2868,N_2987);
nand UO_321 (O_321,N_2918,N_2581);
and UO_322 (O_322,N_2551,N_2471);
nor UO_323 (O_323,N_2793,N_2830);
and UO_324 (O_324,N_2549,N_2798);
nand UO_325 (O_325,N_2852,N_2833);
and UO_326 (O_326,N_2713,N_2780);
and UO_327 (O_327,N_2411,N_2902);
xnor UO_328 (O_328,N_2954,N_2763);
xor UO_329 (O_329,N_2423,N_2772);
nand UO_330 (O_330,N_2693,N_2449);
and UO_331 (O_331,N_2599,N_2474);
or UO_332 (O_332,N_2827,N_2934);
nand UO_333 (O_333,N_2685,N_2955);
nand UO_334 (O_334,N_2703,N_2905);
nand UO_335 (O_335,N_2435,N_2679);
nor UO_336 (O_336,N_2818,N_2653);
nor UO_337 (O_337,N_2638,N_2450);
xor UO_338 (O_338,N_2478,N_2477);
nor UO_339 (O_339,N_2433,N_2802);
and UO_340 (O_340,N_2413,N_2492);
nand UO_341 (O_341,N_2954,N_2632);
nand UO_342 (O_342,N_2806,N_2827);
xnor UO_343 (O_343,N_2918,N_2743);
nand UO_344 (O_344,N_2401,N_2611);
or UO_345 (O_345,N_2510,N_2631);
or UO_346 (O_346,N_2986,N_2526);
nor UO_347 (O_347,N_2735,N_2643);
or UO_348 (O_348,N_2597,N_2527);
or UO_349 (O_349,N_2909,N_2751);
nand UO_350 (O_350,N_2552,N_2823);
nand UO_351 (O_351,N_2766,N_2823);
nor UO_352 (O_352,N_2557,N_2556);
nand UO_353 (O_353,N_2462,N_2836);
and UO_354 (O_354,N_2419,N_2722);
nand UO_355 (O_355,N_2421,N_2869);
nor UO_356 (O_356,N_2769,N_2669);
and UO_357 (O_357,N_2410,N_2805);
or UO_358 (O_358,N_2658,N_2816);
and UO_359 (O_359,N_2463,N_2460);
and UO_360 (O_360,N_2852,N_2544);
xnor UO_361 (O_361,N_2692,N_2804);
nor UO_362 (O_362,N_2801,N_2887);
or UO_363 (O_363,N_2746,N_2863);
and UO_364 (O_364,N_2956,N_2652);
nand UO_365 (O_365,N_2939,N_2942);
and UO_366 (O_366,N_2736,N_2484);
and UO_367 (O_367,N_2571,N_2626);
and UO_368 (O_368,N_2471,N_2686);
nor UO_369 (O_369,N_2748,N_2981);
and UO_370 (O_370,N_2407,N_2891);
nand UO_371 (O_371,N_2692,N_2744);
and UO_372 (O_372,N_2524,N_2883);
and UO_373 (O_373,N_2701,N_2538);
and UO_374 (O_374,N_2985,N_2722);
nor UO_375 (O_375,N_2680,N_2585);
or UO_376 (O_376,N_2893,N_2583);
nand UO_377 (O_377,N_2761,N_2649);
nand UO_378 (O_378,N_2605,N_2478);
and UO_379 (O_379,N_2875,N_2998);
and UO_380 (O_380,N_2695,N_2459);
nand UO_381 (O_381,N_2524,N_2500);
nand UO_382 (O_382,N_2816,N_2438);
or UO_383 (O_383,N_2575,N_2766);
and UO_384 (O_384,N_2516,N_2987);
nand UO_385 (O_385,N_2616,N_2879);
nand UO_386 (O_386,N_2538,N_2625);
or UO_387 (O_387,N_2705,N_2775);
and UO_388 (O_388,N_2846,N_2699);
nand UO_389 (O_389,N_2511,N_2561);
nor UO_390 (O_390,N_2758,N_2947);
and UO_391 (O_391,N_2439,N_2505);
nand UO_392 (O_392,N_2789,N_2488);
and UO_393 (O_393,N_2981,N_2727);
or UO_394 (O_394,N_2418,N_2799);
nand UO_395 (O_395,N_2436,N_2753);
nand UO_396 (O_396,N_2403,N_2533);
or UO_397 (O_397,N_2432,N_2961);
and UO_398 (O_398,N_2448,N_2721);
nor UO_399 (O_399,N_2673,N_2998);
and UO_400 (O_400,N_2865,N_2704);
or UO_401 (O_401,N_2960,N_2788);
nor UO_402 (O_402,N_2793,N_2936);
nand UO_403 (O_403,N_2524,N_2851);
nand UO_404 (O_404,N_2653,N_2959);
or UO_405 (O_405,N_2404,N_2847);
nor UO_406 (O_406,N_2773,N_2856);
nand UO_407 (O_407,N_2888,N_2807);
and UO_408 (O_408,N_2539,N_2988);
or UO_409 (O_409,N_2637,N_2411);
or UO_410 (O_410,N_2991,N_2899);
nand UO_411 (O_411,N_2623,N_2429);
or UO_412 (O_412,N_2697,N_2630);
xnor UO_413 (O_413,N_2962,N_2707);
or UO_414 (O_414,N_2569,N_2972);
xnor UO_415 (O_415,N_2887,N_2519);
or UO_416 (O_416,N_2895,N_2676);
and UO_417 (O_417,N_2884,N_2462);
nand UO_418 (O_418,N_2458,N_2982);
xor UO_419 (O_419,N_2650,N_2824);
and UO_420 (O_420,N_2611,N_2962);
nand UO_421 (O_421,N_2718,N_2687);
nor UO_422 (O_422,N_2611,N_2698);
and UO_423 (O_423,N_2920,N_2874);
or UO_424 (O_424,N_2444,N_2540);
nor UO_425 (O_425,N_2629,N_2913);
nor UO_426 (O_426,N_2852,N_2648);
nor UO_427 (O_427,N_2986,N_2644);
nand UO_428 (O_428,N_2566,N_2903);
xnor UO_429 (O_429,N_2951,N_2923);
or UO_430 (O_430,N_2659,N_2928);
and UO_431 (O_431,N_2523,N_2563);
and UO_432 (O_432,N_2864,N_2550);
or UO_433 (O_433,N_2437,N_2974);
xnor UO_434 (O_434,N_2566,N_2782);
or UO_435 (O_435,N_2539,N_2467);
or UO_436 (O_436,N_2906,N_2642);
and UO_437 (O_437,N_2587,N_2607);
nor UO_438 (O_438,N_2913,N_2559);
or UO_439 (O_439,N_2992,N_2577);
nand UO_440 (O_440,N_2543,N_2947);
nor UO_441 (O_441,N_2587,N_2405);
nand UO_442 (O_442,N_2614,N_2466);
xnor UO_443 (O_443,N_2668,N_2558);
nor UO_444 (O_444,N_2530,N_2610);
or UO_445 (O_445,N_2747,N_2744);
or UO_446 (O_446,N_2465,N_2525);
nor UO_447 (O_447,N_2810,N_2400);
nand UO_448 (O_448,N_2843,N_2619);
nor UO_449 (O_449,N_2448,N_2976);
or UO_450 (O_450,N_2441,N_2803);
or UO_451 (O_451,N_2687,N_2757);
xnor UO_452 (O_452,N_2561,N_2825);
xor UO_453 (O_453,N_2958,N_2479);
nor UO_454 (O_454,N_2672,N_2702);
and UO_455 (O_455,N_2873,N_2638);
nand UO_456 (O_456,N_2554,N_2565);
xnor UO_457 (O_457,N_2423,N_2932);
xor UO_458 (O_458,N_2763,N_2619);
nor UO_459 (O_459,N_2954,N_2677);
and UO_460 (O_460,N_2779,N_2948);
and UO_461 (O_461,N_2833,N_2708);
and UO_462 (O_462,N_2940,N_2832);
or UO_463 (O_463,N_2494,N_2637);
and UO_464 (O_464,N_2490,N_2430);
nand UO_465 (O_465,N_2453,N_2859);
or UO_466 (O_466,N_2410,N_2466);
nor UO_467 (O_467,N_2761,N_2855);
and UO_468 (O_468,N_2618,N_2494);
nand UO_469 (O_469,N_2800,N_2703);
and UO_470 (O_470,N_2503,N_2510);
xor UO_471 (O_471,N_2947,N_2877);
xnor UO_472 (O_472,N_2576,N_2529);
or UO_473 (O_473,N_2756,N_2696);
and UO_474 (O_474,N_2432,N_2416);
nand UO_475 (O_475,N_2575,N_2629);
nand UO_476 (O_476,N_2539,N_2882);
nand UO_477 (O_477,N_2881,N_2795);
or UO_478 (O_478,N_2574,N_2738);
nand UO_479 (O_479,N_2858,N_2956);
nor UO_480 (O_480,N_2961,N_2986);
nand UO_481 (O_481,N_2930,N_2820);
nand UO_482 (O_482,N_2941,N_2443);
xor UO_483 (O_483,N_2762,N_2664);
nor UO_484 (O_484,N_2860,N_2513);
xnor UO_485 (O_485,N_2598,N_2493);
xnor UO_486 (O_486,N_2550,N_2720);
and UO_487 (O_487,N_2929,N_2972);
or UO_488 (O_488,N_2627,N_2810);
nand UO_489 (O_489,N_2965,N_2566);
nor UO_490 (O_490,N_2911,N_2727);
xor UO_491 (O_491,N_2577,N_2989);
nor UO_492 (O_492,N_2501,N_2741);
xnor UO_493 (O_493,N_2437,N_2659);
and UO_494 (O_494,N_2773,N_2524);
xor UO_495 (O_495,N_2687,N_2612);
nand UO_496 (O_496,N_2993,N_2962);
or UO_497 (O_497,N_2651,N_2741);
or UO_498 (O_498,N_2680,N_2858);
xnor UO_499 (O_499,N_2881,N_2461);
endmodule