module basic_750_5000_1000_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_268,In_438);
nand U1 (N_1,In_383,In_418);
and U2 (N_2,In_247,In_595);
xnor U3 (N_3,In_458,In_87);
and U4 (N_4,In_167,In_539);
xor U5 (N_5,In_544,In_546);
nor U6 (N_6,In_370,In_38);
xnor U7 (N_7,In_697,In_22);
xnor U8 (N_8,In_4,In_447);
and U9 (N_9,In_643,In_580);
xor U10 (N_10,In_675,In_282);
nor U11 (N_11,In_319,In_56);
nor U12 (N_12,In_484,In_355);
xnor U13 (N_13,In_474,In_563);
xnor U14 (N_14,In_227,In_23);
and U15 (N_15,In_210,In_288);
or U16 (N_16,In_341,In_224);
xnor U17 (N_17,In_688,In_242);
nor U18 (N_18,In_535,In_47);
nor U19 (N_19,In_538,In_165);
xor U20 (N_20,In_274,In_482);
and U21 (N_21,In_492,In_453);
nand U22 (N_22,In_521,In_507);
nor U23 (N_23,In_245,In_145);
and U24 (N_24,In_321,In_510);
nor U25 (N_25,In_259,In_333);
or U26 (N_26,In_309,In_327);
or U27 (N_27,In_138,In_515);
nor U28 (N_28,In_212,In_1);
nor U29 (N_29,In_106,In_740);
xor U30 (N_30,In_359,In_394);
xnor U31 (N_31,In_419,In_99);
and U32 (N_32,In_400,In_496);
xor U33 (N_33,In_253,In_69);
and U34 (N_34,In_201,In_631);
and U35 (N_35,In_32,In_91);
nand U36 (N_36,In_218,In_78);
nand U37 (N_37,In_410,In_735);
nor U38 (N_38,In_3,In_293);
xnor U39 (N_39,In_207,In_582);
or U40 (N_40,In_188,In_72);
xor U41 (N_41,In_565,In_96);
xnor U42 (N_42,In_486,In_391);
or U43 (N_43,In_585,In_202);
and U44 (N_44,In_52,In_80);
nand U45 (N_45,In_456,In_665);
or U46 (N_46,In_275,In_471);
xnor U47 (N_47,In_555,In_107);
nand U48 (N_48,In_264,In_360);
or U49 (N_49,In_64,In_708);
and U50 (N_50,In_266,In_386);
nand U51 (N_51,In_426,In_663);
nand U52 (N_52,In_692,In_35);
or U53 (N_53,In_720,In_694);
nand U54 (N_54,In_412,In_377);
nor U55 (N_55,In_34,In_488);
xor U56 (N_56,In_123,In_609);
and U57 (N_57,In_57,In_340);
nand U58 (N_58,In_473,In_173);
nor U59 (N_59,In_304,In_232);
nand U60 (N_60,In_379,In_113);
nor U61 (N_61,In_334,In_706);
nor U62 (N_62,In_598,In_130);
nor U63 (N_63,In_85,In_661);
or U64 (N_64,In_323,In_193);
nand U65 (N_65,In_351,In_660);
or U66 (N_66,In_483,In_635);
and U67 (N_67,In_110,In_448);
nand U68 (N_68,In_166,In_168);
nand U69 (N_69,In_689,In_393);
nand U70 (N_70,In_147,In_435);
nor U71 (N_71,In_623,In_709);
nand U72 (N_72,In_707,In_325);
and U73 (N_73,In_137,In_525);
nor U74 (N_74,In_650,In_672);
nand U75 (N_75,In_701,In_90);
and U76 (N_76,In_656,In_671);
nand U77 (N_77,In_28,In_125);
and U78 (N_78,In_151,In_417);
or U79 (N_79,In_430,In_40);
xnor U80 (N_80,In_208,In_365);
and U81 (N_81,In_249,In_562);
or U82 (N_82,In_378,In_463);
nand U83 (N_83,In_746,In_508);
xnor U84 (N_84,In_577,In_285);
or U85 (N_85,In_454,In_440);
or U86 (N_86,In_5,In_462);
xor U87 (N_87,In_251,In_112);
and U88 (N_88,In_53,In_586);
nand U89 (N_89,In_213,In_558);
xnor U90 (N_90,In_639,In_200);
xor U91 (N_91,In_673,In_33);
or U92 (N_92,In_633,In_556);
xor U93 (N_93,In_342,In_399);
or U94 (N_94,In_315,In_573);
and U95 (N_95,In_127,In_31);
xor U96 (N_96,In_414,In_375);
or U97 (N_97,In_194,In_731);
nand U98 (N_98,In_445,In_286);
or U99 (N_99,In_183,In_551);
nor U100 (N_100,In_144,In_662);
nand U101 (N_101,In_326,In_714);
xor U102 (N_102,In_135,In_49);
and U103 (N_103,In_512,In_14);
xor U104 (N_104,In_12,In_726);
and U105 (N_105,In_362,In_46);
and U106 (N_106,In_613,In_528);
nor U107 (N_107,In_742,In_339);
or U108 (N_108,In_615,In_605);
or U109 (N_109,In_256,In_284);
and U110 (N_110,In_103,In_199);
nand U111 (N_111,In_296,In_710);
and U112 (N_112,In_402,In_429);
xnor U113 (N_113,In_248,In_353);
nand U114 (N_114,In_617,In_713);
and U115 (N_115,In_344,In_600);
or U116 (N_116,In_686,In_197);
xor U117 (N_117,In_612,In_308);
and U118 (N_118,In_126,In_579);
xnor U119 (N_119,In_185,In_277);
and U120 (N_120,In_398,In_36);
or U121 (N_121,In_603,In_316);
nand U122 (N_122,In_132,In_516);
and U123 (N_123,In_567,In_230);
xor U124 (N_124,In_743,In_269);
and U125 (N_125,In_497,In_221);
nor U126 (N_126,In_728,In_470);
xor U127 (N_127,In_206,In_541);
and U128 (N_128,In_225,In_519);
nor U129 (N_129,In_150,In_322);
or U130 (N_130,In_654,In_273);
nor U131 (N_131,In_587,In_629);
or U132 (N_132,In_390,In_244);
nor U133 (N_133,In_217,In_18);
nand U134 (N_134,In_566,In_11);
nand U135 (N_135,In_310,In_718);
nor U136 (N_136,In_174,In_156);
xnor U137 (N_137,In_401,In_680);
nor U138 (N_138,In_608,In_128);
xor U139 (N_139,In_65,In_494);
xnor U140 (N_140,In_659,In_55);
and U141 (N_141,In_161,In_343);
nand U142 (N_142,In_584,In_349);
and U143 (N_143,In_677,In_95);
and U144 (N_144,In_478,In_411);
or U145 (N_145,In_588,In_721);
or U146 (N_146,In_279,In_644);
nand U147 (N_147,In_564,In_203);
and U148 (N_148,In_0,In_108);
and U149 (N_149,In_589,In_278);
and U150 (N_150,In_243,In_198);
or U151 (N_151,In_283,In_58);
or U152 (N_152,In_100,In_569);
nor U153 (N_153,In_744,In_748);
or U154 (N_154,In_502,In_363);
xnor U155 (N_155,In_690,In_485);
xnor U156 (N_156,In_88,In_298);
nor U157 (N_157,In_177,In_531);
or U158 (N_158,In_83,In_517);
nor U159 (N_159,In_254,In_260);
nand U160 (N_160,In_594,In_666);
nand U161 (N_161,In_66,In_336);
nand U162 (N_162,In_468,In_318);
nand U163 (N_163,In_724,In_619);
nand U164 (N_164,In_530,In_543);
or U165 (N_165,In_331,In_387);
nor U166 (N_166,In_547,In_591);
and U167 (N_167,In_117,In_271);
nand U168 (N_168,In_446,In_648);
or U169 (N_169,In_157,In_652);
and U170 (N_170,In_596,In_26);
or U171 (N_171,In_733,In_76);
nand U172 (N_172,In_477,In_114);
and U173 (N_173,In_21,In_30);
or U174 (N_174,In_186,In_634);
or U175 (N_175,In_739,In_373);
xor U176 (N_176,In_719,In_532);
or U177 (N_177,In_730,In_548);
or U178 (N_178,In_441,In_523);
and U179 (N_179,In_736,In_592);
or U180 (N_180,In_493,In_537);
or U181 (N_181,In_314,In_215);
xnor U182 (N_182,In_54,In_44);
and U183 (N_183,In_364,In_664);
nor U184 (N_184,In_101,In_674);
nand U185 (N_185,In_518,In_311);
nand U186 (N_186,In_27,In_272);
and U187 (N_187,In_59,In_382);
or U188 (N_188,In_307,In_653);
and U189 (N_189,In_574,In_153);
nor U190 (N_190,In_433,In_231);
or U191 (N_191,In_550,In_189);
or U192 (N_192,In_306,In_238);
or U193 (N_193,In_667,In_741);
or U194 (N_194,In_214,In_122);
and U195 (N_195,In_646,In_190);
and U196 (N_196,In_368,In_683);
xnor U197 (N_197,In_7,In_571);
nand U198 (N_198,In_301,In_529);
nand U199 (N_199,In_17,In_641);
and U200 (N_200,In_422,In_403);
nand U201 (N_201,In_747,In_389);
nand U202 (N_202,In_261,In_572);
nor U203 (N_203,In_226,In_459);
nand U204 (N_204,In_16,In_159);
nand U205 (N_205,In_599,In_649);
nor U206 (N_206,In_729,In_143);
nor U207 (N_207,In_475,In_223);
nor U208 (N_208,In_449,In_61);
nor U209 (N_209,In_172,In_71);
and U210 (N_210,In_255,In_404);
xnor U211 (N_211,In_732,In_415);
xor U212 (N_212,In_361,In_102);
nand U213 (N_213,In_68,In_104);
nand U214 (N_214,In_263,In_75);
nor U215 (N_215,In_427,In_229);
nor U216 (N_216,In_679,In_469);
and U217 (N_217,In_554,In_703);
or U218 (N_218,In_39,In_366);
or U219 (N_219,In_669,In_237);
nand U220 (N_220,In_116,In_6);
xnor U221 (N_221,In_324,In_372);
and U222 (N_222,In_220,In_424);
xnor U223 (N_223,In_111,In_124);
nor U224 (N_224,In_630,In_678);
nor U225 (N_225,In_380,In_534);
nand U226 (N_226,In_235,In_62);
xnor U227 (N_227,In_495,In_406);
nand U228 (N_228,In_711,In_570);
nor U229 (N_229,In_158,In_487);
nor U230 (N_230,In_70,In_109);
xnor U231 (N_231,In_211,In_60);
xor U232 (N_232,In_347,In_560);
and U233 (N_233,In_628,In_352);
and U234 (N_234,In_503,In_51);
xnor U235 (N_235,In_581,In_506);
nand U236 (N_236,In_489,In_131);
and U237 (N_237,In_722,In_460);
nor U238 (N_238,In_542,In_552);
nor U239 (N_239,In_171,In_413);
or U240 (N_240,In_170,In_627);
and U241 (N_241,In_303,In_191);
or U242 (N_242,In_337,In_696);
nand U243 (N_243,In_294,In_265);
nor U244 (N_244,In_638,In_681);
nor U245 (N_245,In_332,In_312);
nand U246 (N_246,In_329,In_524);
nor U247 (N_247,In_620,In_616);
xor U248 (N_248,In_241,In_50);
or U249 (N_249,In_670,In_610);
and U250 (N_250,In_43,In_444);
nand U251 (N_251,In_118,In_149);
nand U252 (N_252,In_396,In_698);
xor U253 (N_253,In_348,In_395);
xnor U254 (N_254,In_15,In_601);
xnor U255 (N_255,In_734,In_621);
and U256 (N_256,In_511,In_295);
xnor U257 (N_257,In_385,In_490);
nand U258 (N_258,In_257,In_451);
nor U259 (N_259,In_19,In_602);
or U260 (N_260,In_606,In_142);
nand U261 (N_261,In_578,In_749);
nor U262 (N_262,In_704,In_642);
or U263 (N_263,In_42,In_182);
nand U264 (N_264,In_317,In_439);
nor U265 (N_265,In_712,In_45);
nor U266 (N_266,In_67,In_436);
nor U267 (N_267,In_184,In_338);
and U268 (N_268,In_479,In_136);
xor U269 (N_269,In_133,In_155);
or U270 (N_270,In_725,In_236);
and U271 (N_271,In_388,In_354);
and U272 (N_272,In_330,In_509);
and U273 (N_273,In_597,In_205);
or U274 (N_274,In_645,In_514);
and U275 (N_275,In_611,In_723);
or U276 (N_276,In_687,In_357);
nand U277 (N_277,In_452,In_397);
and U278 (N_278,In_501,In_745);
and U279 (N_279,In_121,In_464);
or U280 (N_280,In_63,In_9);
and U281 (N_281,In_302,In_392);
or U282 (N_282,In_89,In_437);
xor U283 (N_283,In_141,In_105);
xnor U284 (N_284,In_407,In_250);
xor U285 (N_285,In_702,In_416);
or U286 (N_286,In_367,In_637);
nor U287 (N_287,In_536,In_222);
nor U288 (N_288,In_561,In_187);
nand U289 (N_289,In_376,In_176);
xor U290 (N_290,In_632,In_162);
nand U291 (N_291,In_239,In_500);
nor U292 (N_292,In_480,In_280);
nor U293 (N_293,In_276,In_540);
and U294 (N_294,In_246,In_358);
or U295 (N_295,In_655,In_119);
or U296 (N_296,In_420,In_291);
nor U297 (N_297,In_262,In_97);
or U298 (N_298,In_685,In_467);
nand U299 (N_299,In_432,In_8);
and U300 (N_300,In_179,In_74);
nand U301 (N_301,In_472,In_73);
nor U302 (N_302,In_727,In_93);
or U303 (N_303,In_614,In_204);
or U304 (N_304,In_527,In_428);
or U305 (N_305,In_216,In_545);
xnor U306 (N_306,In_647,In_25);
nand U307 (N_307,In_526,In_421);
nor U308 (N_308,In_575,In_450);
nand U309 (N_309,In_289,In_181);
nor U310 (N_310,In_651,In_498);
or U311 (N_311,In_593,In_715);
or U312 (N_312,In_693,In_233);
and U313 (N_313,In_115,In_684);
xnor U314 (N_314,In_154,In_270);
xor U315 (N_315,In_499,In_676);
nor U316 (N_316,In_408,In_409);
nand U317 (N_317,In_146,In_625);
nor U318 (N_318,In_129,In_668);
xnor U319 (N_319,In_658,In_24);
or U320 (N_320,In_94,In_37);
and U321 (N_321,In_41,In_20);
and U322 (N_322,In_299,In_576);
nor U323 (N_323,In_82,In_695);
and U324 (N_324,In_2,In_29);
or U325 (N_325,In_369,In_86);
nor U326 (N_326,In_292,In_175);
or U327 (N_327,In_491,In_180);
or U328 (N_328,In_636,In_13);
xnor U329 (N_329,In_196,In_228);
or U330 (N_330,In_140,In_476);
nand U331 (N_331,In_79,In_346);
and U332 (N_332,In_192,In_152);
xor U333 (N_333,In_290,In_10);
nor U334 (N_334,In_305,In_405);
xor U335 (N_335,In_267,In_700);
xnor U336 (N_336,In_705,In_691);
nor U337 (N_337,In_481,In_163);
nand U338 (N_338,In_559,In_504);
nor U339 (N_339,In_657,In_624);
and U340 (N_340,In_92,In_443);
and U341 (N_341,In_622,In_195);
and U342 (N_342,In_520,In_84);
or U343 (N_343,In_465,In_640);
or U344 (N_344,In_607,In_77);
nor U345 (N_345,In_209,In_381);
nor U346 (N_346,In_505,In_350);
xnor U347 (N_347,In_328,In_169);
nand U348 (N_348,In_626,In_583);
and U349 (N_349,In_513,In_604);
or U350 (N_350,In_425,In_618);
nor U351 (N_351,In_219,In_434);
xor U352 (N_352,In_374,In_252);
and U353 (N_353,In_335,In_568);
or U354 (N_354,In_466,In_48);
and U355 (N_355,In_431,In_345);
nor U356 (N_356,In_371,In_590);
nor U357 (N_357,In_81,In_557);
nor U358 (N_358,In_455,In_240);
and U359 (N_359,In_164,In_716);
nor U360 (N_360,In_738,In_533);
nand U361 (N_361,In_297,In_717);
nor U362 (N_362,In_160,In_442);
xnor U363 (N_363,In_178,In_461);
or U364 (N_364,In_522,In_737);
or U365 (N_365,In_313,In_134);
and U366 (N_366,In_457,In_384);
or U367 (N_367,In_120,In_139);
nand U368 (N_368,In_287,In_549);
nand U369 (N_369,In_356,In_234);
xnor U370 (N_370,In_423,In_300);
nand U371 (N_371,In_320,In_682);
nand U372 (N_372,In_148,In_98);
or U373 (N_373,In_553,In_281);
xor U374 (N_374,In_258,In_699);
or U375 (N_375,In_164,In_744);
nor U376 (N_376,In_47,In_615);
nor U377 (N_377,In_421,In_452);
and U378 (N_378,In_44,In_260);
nor U379 (N_379,In_572,In_16);
and U380 (N_380,In_323,In_342);
or U381 (N_381,In_272,In_200);
or U382 (N_382,In_532,In_351);
nor U383 (N_383,In_440,In_301);
or U384 (N_384,In_104,In_710);
nand U385 (N_385,In_538,In_699);
nand U386 (N_386,In_516,In_675);
nand U387 (N_387,In_460,In_586);
xor U388 (N_388,In_449,In_261);
or U389 (N_389,In_341,In_180);
or U390 (N_390,In_366,In_619);
nor U391 (N_391,In_33,In_64);
or U392 (N_392,In_235,In_529);
and U393 (N_393,In_652,In_354);
nor U394 (N_394,In_3,In_506);
xor U395 (N_395,In_331,In_257);
xnor U396 (N_396,In_298,In_544);
or U397 (N_397,In_202,In_579);
xor U398 (N_398,In_495,In_159);
and U399 (N_399,In_95,In_617);
xor U400 (N_400,In_410,In_135);
or U401 (N_401,In_593,In_104);
nand U402 (N_402,In_494,In_141);
and U403 (N_403,In_733,In_379);
or U404 (N_404,In_616,In_717);
nor U405 (N_405,In_654,In_583);
xor U406 (N_406,In_607,In_535);
xnor U407 (N_407,In_156,In_107);
or U408 (N_408,In_30,In_669);
and U409 (N_409,In_39,In_735);
nor U410 (N_410,In_81,In_391);
nor U411 (N_411,In_577,In_3);
nand U412 (N_412,In_301,In_749);
or U413 (N_413,In_671,In_749);
xor U414 (N_414,In_13,In_352);
nor U415 (N_415,In_91,In_472);
and U416 (N_416,In_68,In_698);
xor U417 (N_417,In_106,In_578);
or U418 (N_418,In_396,In_80);
and U419 (N_419,In_135,In_635);
nand U420 (N_420,In_414,In_575);
nand U421 (N_421,In_42,In_193);
and U422 (N_422,In_698,In_323);
nand U423 (N_423,In_435,In_189);
nand U424 (N_424,In_38,In_115);
and U425 (N_425,In_502,In_247);
nand U426 (N_426,In_724,In_650);
xnor U427 (N_427,In_161,In_547);
nor U428 (N_428,In_165,In_49);
and U429 (N_429,In_48,In_419);
and U430 (N_430,In_270,In_66);
nor U431 (N_431,In_732,In_361);
or U432 (N_432,In_497,In_92);
and U433 (N_433,In_10,In_526);
or U434 (N_434,In_161,In_445);
or U435 (N_435,In_582,In_412);
or U436 (N_436,In_351,In_277);
or U437 (N_437,In_476,In_544);
nor U438 (N_438,In_684,In_216);
xor U439 (N_439,In_472,In_151);
nand U440 (N_440,In_734,In_194);
nand U441 (N_441,In_92,In_234);
xnor U442 (N_442,In_363,In_405);
and U443 (N_443,In_35,In_207);
or U444 (N_444,In_52,In_553);
nand U445 (N_445,In_359,In_603);
nand U446 (N_446,In_367,In_22);
nor U447 (N_447,In_336,In_583);
and U448 (N_448,In_85,In_45);
xor U449 (N_449,In_533,In_301);
or U450 (N_450,In_432,In_459);
and U451 (N_451,In_693,In_542);
nand U452 (N_452,In_99,In_393);
xnor U453 (N_453,In_248,In_701);
and U454 (N_454,In_85,In_248);
xnor U455 (N_455,In_75,In_589);
nand U456 (N_456,In_705,In_715);
xor U457 (N_457,In_114,In_299);
or U458 (N_458,In_338,In_188);
nand U459 (N_459,In_2,In_236);
nor U460 (N_460,In_441,In_519);
and U461 (N_461,In_309,In_481);
xnor U462 (N_462,In_573,In_699);
nor U463 (N_463,In_142,In_307);
and U464 (N_464,In_693,In_372);
xor U465 (N_465,In_296,In_176);
and U466 (N_466,In_346,In_16);
or U467 (N_467,In_629,In_446);
or U468 (N_468,In_727,In_446);
nor U469 (N_469,In_289,In_282);
xor U470 (N_470,In_432,In_348);
xnor U471 (N_471,In_467,In_390);
nor U472 (N_472,In_633,In_645);
or U473 (N_473,In_635,In_68);
and U474 (N_474,In_634,In_492);
nor U475 (N_475,In_311,In_654);
xor U476 (N_476,In_329,In_658);
or U477 (N_477,In_540,In_196);
or U478 (N_478,In_437,In_450);
or U479 (N_479,In_104,In_395);
xnor U480 (N_480,In_388,In_651);
nor U481 (N_481,In_45,In_203);
or U482 (N_482,In_387,In_611);
nor U483 (N_483,In_262,In_25);
xnor U484 (N_484,In_89,In_537);
nand U485 (N_485,In_378,In_541);
nand U486 (N_486,In_72,In_710);
xnor U487 (N_487,In_532,In_401);
nand U488 (N_488,In_304,In_89);
and U489 (N_489,In_50,In_555);
and U490 (N_490,In_132,In_219);
and U491 (N_491,In_700,In_153);
or U492 (N_492,In_41,In_377);
and U493 (N_493,In_33,In_309);
and U494 (N_494,In_150,In_400);
or U495 (N_495,In_346,In_140);
xor U496 (N_496,In_145,In_39);
and U497 (N_497,In_679,In_327);
or U498 (N_498,In_647,In_31);
nand U499 (N_499,In_672,In_504);
or U500 (N_500,In_334,In_108);
nand U501 (N_501,In_736,In_729);
xnor U502 (N_502,In_389,In_191);
xnor U503 (N_503,In_486,In_80);
nand U504 (N_504,In_638,In_270);
nor U505 (N_505,In_77,In_736);
nor U506 (N_506,In_68,In_563);
nand U507 (N_507,In_244,In_471);
nand U508 (N_508,In_445,In_7);
or U509 (N_509,In_587,In_502);
nand U510 (N_510,In_316,In_619);
or U511 (N_511,In_321,In_349);
and U512 (N_512,In_393,In_595);
or U513 (N_513,In_97,In_403);
and U514 (N_514,In_559,In_108);
nor U515 (N_515,In_678,In_687);
xnor U516 (N_516,In_70,In_132);
or U517 (N_517,In_527,In_9);
nand U518 (N_518,In_526,In_378);
and U519 (N_519,In_48,In_723);
xnor U520 (N_520,In_398,In_444);
nand U521 (N_521,In_715,In_537);
nand U522 (N_522,In_638,In_125);
or U523 (N_523,In_658,In_190);
xnor U524 (N_524,In_429,In_472);
xor U525 (N_525,In_661,In_486);
or U526 (N_526,In_314,In_595);
nor U527 (N_527,In_30,In_288);
nand U528 (N_528,In_371,In_630);
nand U529 (N_529,In_305,In_24);
nand U530 (N_530,In_250,In_295);
nor U531 (N_531,In_538,In_104);
or U532 (N_532,In_538,In_32);
xnor U533 (N_533,In_426,In_401);
nand U534 (N_534,In_530,In_555);
and U535 (N_535,In_433,In_738);
nand U536 (N_536,In_80,In_724);
nand U537 (N_537,In_453,In_27);
and U538 (N_538,In_621,In_467);
nand U539 (N_539,In_588,In_472);
xnor U540 (N_540,In_556,In_291);
xor U541 (N_541,In_344,In_82);
and U542 (N_542,In_189,In_81);
nor U543 (N_543,In_403,In_456);
and U544 (N_544,In_222,In_165);
xnor U545 (N_545,In_211,In_308);
and U546 (N_546,In_15,In_502);
xor U547 (N_547,In_172,In_30);
xnor U548 (N_548,In_225,In_740);
and U549 (N_549,In_444,In_459);
nand U550 (N_550,In_702,In_372);
nor U551 (N_551,In_137,In_271);
xnor U552 (N_552,In_458,In_487);
nor U553 (N_553,In_258,In_83);
and U554 (N_554,In_659,In_399);
xnor U555 (N_555,In_226,In_296);
nor U556 (N_556,In_191,In_218);
nor U557 (N_557,In_737,In_241);
or U558 (N_558,In_692,In_577);
nand U559 (N_559,In_479,In_428);
and U560 (N_560,In_280,In_323);
xor U561 (N_561,In_704,In_257);
nor U562 (N_562,In_67,In_23);
xnor U563 (N_563,In_394,In_269);
and U564 (N_564,In_453,In_299);
xnor U565 (N_565,In_309,In_490);
and U566 (N_566,In_570,In_478);
nor U567 (N_567,In_213,In_143);
or U568 (N_568,In_271,In_706);
xnor U569 (N_569,In_88,In_653);
and U570 (N_570,In_428,In_408);
and U571 (N_571,In_534,In_526);
or U572 (N_572,In_670,In_17);
and U573 (N_573,In_709,In_215);
nor U574 (N_574,In_486,In_684);
nor U575 (N_575,In_562,In_609);
nor U576 (N_576,In_114,In_536);
xor U577 (N_577,In_694,In_525);
or U578 (N_578,In_181,In_258);
nand U579 (N_579,In_408,In_68);
nor U580 (N_580,In_284,In_320);
nand U581 (N_581,In_411,In_26);
xor U582 (N_582,In_60,In_325);
nand U583 (N_583,In_559,In_463);
nand U584 (N_584,In_153,In_456);
xnor U585 (N_585,In_58,In_171);
nand U586 (N_586,In_620,In_110);
xnor U587 (N_587,In_109,In_33);
nor U588 (N_588,In_351,In_626);
and U589 (N_589,In_115,In_410);
or U590 (N_590,In_439,In_512);
and U591 (N_591,In_130,In_736);
nor U592 (N_592,In_614,In_501);
or U593 (N_593,In_646,In_313);
xor U594 (N_594,In_154,In_555);
nor U595 (N_595,In_583,In_223);
nor U596 (N_596,In_689,In_70);
nor U597 (N_597,In_542,In_667);
xor U598 (N_598,In_86,In_428);
nand U599 (N_599,In_201,In_742);
nand U600 (N_600,In_428,In_373);
and U601 (N_601,In_216,In_560);
nor U602 (N_602,In_171,In_159);
or U603 (N_603,In_149,In_39);
and U604 (N_604,In_251,In_749);
xor U605 (N_605,In_197,In_514);
nor U606 (N_606,In_368,In_6);
xnor U607 (N_607,In_296,In_18);
and U608 (N_608,In_377,In_17);
or U609 (N_609,In_289,In_313);
or U610 (N_610,In_423,In_8);
and U611 (N_611,In_684,In_156);
or U612 (N_612,In_435,In_199);
nand U613 (N_613,In_47,In_685);
nor U614 (N_614,In_151,In_585);
nor U615 (N_615,In_472,In_166);
nand U616 (N_616,In_670,In_136);
nor U617 (N_617,In_21,In_685);
or U618 (N_618,In_457,In_126);
or U619 (N_619,In_61,In_511);
or U620 (N_620,In_509,In_25);
and U621 (N_621,In_452,In_445);
xnor U622 (N_622,In_500,In_735);
nand U623 (N_623,In_255,In_291);
nand U624 (N_624,In_432,In_290);
nand U625 (N_625,In_186,In_725);
nor U626 (N_626,In_356,In_115);
nand U627 (N_627,In_633,In_502);
nand U628 (N_628,In_329,In_83);
xnor U629 (N_629,In_112,In_583);
and U630 (N_630,In_165,In_204);
or U631 (N_631,In_442,In_228);
nor U632 (N_632,In_721,In_344);
or U633 (N_633,In_195,In_444);
nor U634 (N_634,In_165,In_548);
or U635 (N_635,In_633,In_327);
and U636 (N_636,In_620,In_589);
or U637 (N_637,In_289,In_304);
xnor U638 (N_638,In_725,In_164);
xnor U639 (N_639,In_462,In_598);
nor U640 (N_640,In_287,In_208);
and U641 (N_641,In_392,In_673);
xnor U642 (N_642,In_471,In_345);
xnor U643 (N_643,In_35,In_373);
xnor U644 (N_644,In_456,In_334);
xor U645 (N_645,In_79,In_445);
xnor U646 (N_646,In_433,In_104);
or U647 (N_647,In_415,In_446);
or U648 (N_648,In_403,In_270);
xor U649 (N_649,In_437,In_202);
xor U650 (N_650,In_655,In_379);
and U651 (N_651,In_55,In_522);
xor U652 (N_652,In_13,In_21);
nor U653 (N_653,In_145,In_711);
or U654 (N_654,In_289,In_417);
or U655 (N_655,In_499,In_409);
nor U656 (N_656,In_100,In_222);
nand U657 (N_657,In_352,In_427);
xor U658 (N_658,In_123,In_176);
xnor U659 (N_659,In_3,In_150);
nand U660 (N_660,In_338,In_9);
and U661 (N_661,In_345,In_43);
nor U662 (N_662,In_120,In_42);
or U663 (N_663,In_671,In_522);
nor U664 (N_664,In_210,In_299);
nand U665 (N_665,In_200,In_293);
or U666 (N_666,In_613,In_394);
nand U667 (N_667,In_5,In_408);
and U668 (N_668,In_75,In_592);
and U669 (N_669,In_257,In_592);
and U670 (N_670,In_710,In_194);
xor U671 (N_671,In_337,In_524);
nand U672 (N_672,In_90,In_312);
nand U673 (N_673,In_89,In_532);
nand U674 (N_674,In_476,In_451);
or U675 (N_675,In_703,In_325);
and U676 (N_676,In_415,In_51);
nand U677 (N_677,In_308,In_465);
nor U678 (N_678,In_736,In_21);
nor U679 (N_679,In_145,In_588);
and U680 (N_680,In_570,In_471);
nor U681 (N_681,In_409,In_659);
and U682 (N_682,In_507,In_143);
or U683 (N_683,In_221,In_625);
xor U684 (N_684,In_557,In_475);
or U685 (N_685,In_200,In_402);
nand U686 (N_686,In_620,In_515);
and U687 (N_687,In_382,In_331);
nand U688 (N_688,In_554,In_12);
and U689 (N_689,In_56,In_282);
or U690 (N_690,In_327,In_536);
xnor U691 (N_691,In_28,In_305);
and U692 (N_692,In_684,In_347);
xnor U693 (N_693,In_606,In_195);
and U694 (N_694,In_412,In_368);
nor U695 (N_695,In_79,In_728);
nand U696 (N_696,In_189,In_486);
and U697 (N_697,In_388,In_280);
xnor U698 (N_698,In_363,In_585);
or U699 (N_699,In_705,In_603);
or U700 (N_700,In_317,In_726);
and U701 (N_701,In_373,In_675);
nand U702 (N_702,In_172,In_81);
xnor U703 (N_703,In_359,In_238);
xnor U704 (N_704,In_651,In_722);
and U705 (N_705,In_491,In_463);
nand U706 (N_706,In_125,In_51);
nand U707 (N_707,In_554,In_137);
or U708 (N_708,In_136,In_177);
xor U709 (N_709,In_632,In_401);
nor U710 (N_710,In_622,In_391);
xnor U711 (N_711,In_164,In_455);
nand U712 (N_712,In_519,In_64);
nor U713 (N_713,In_392,In_659);
xor U714 (N_714,In_581,In_440);
nand U715 (N_715,In_14,In_192);
nor U716 (N_716,In_657,In_665);
nor U717 (N_717,In_452,In_536);
nor U718 (N_718,In_464,In_589);
nand U719 (N_719,In_443,In_429);
and U720 (N_720,In_54,In_37);
nand U721 (N_721,In_356,In_471);
nor U722 (N_722,In_295,In_325);
xnor U723 (N_723,In_656,In_362);
and U724 (N_724,In_26,In_150);
xor U725 (N_725,In_349,In_41);
nor U726 (N_726,In_155,In_281);
xnor U727 (N_727,In_618,In_240);
nor U728 (N_728,In_129,In_373);
and U729 (N_729,In_635,In_254);
xor U730 (N_730,In_57,In_208);
or U731 (N_731,In_545,In_635);
or U732 (N_732,In_189,In_392);
xnor U733 (N_733,In_145,In_586);
nand U734 (N_734,In_240,In_460);
nand U735 (N_735,In_489,In_150);
nor U736 (N_736,In_74,In_406);
and U737 (N_737,In_189,In_637);
nand U738 (N_738,In_452,In_619);
nor U739 (N_739,In_32,In_486);
or U740 (N_740,In_243,In_162);
and U741 (N_741,In_740,In_86);
xor U742 (N_742,In_325,In_74);
or U743 (N_743,In_3,In_520);
xnor U744 (N_744,In_411,In_351);
xor U745 (N_745,In_436,In_535);
nor U746 (N_746,In_620,In_95);
nor U747 (N_747,In_355,In_509);
and U748 (N_748,In_570,In_73);
nor U749 (N_749,In_99,In_256);
nand U750 (N_750,In_434,In_123);
nor U751 (N_751,In_388,In_525);
or U752 (N_752,In_56,In_89);
xor U753 (N_753,In_551,In_722);
and U754 (N_754,In_679,In_577);
nor U755 (N_755,In_664,In_86);
xor U756 (N_756,In_446,In_425);
xnor U757 (N_757,In_694,In_298);
and U758 (N_758,In_285,In_316);
nand U759 (N_759,In_740,In_9);
or U760 (N_760,In_591,In_535);
nor U761 (N_761,In_436,In_171);
or U762 (N_762,In_107,In_212);
xnor U763 (N_763,In_162,In_184);
nand U764 (N_764,In_326,In_642);
nor U765 (N_765,In_305,In_446);
nor U766 (N_766,In_27,In_281);
xnor U767 (N_767,In_118,In_427);
and U768 (N_768,In_58,In_185);
xnor U769 (N_769,In_245,In_290);
and U770 (N_770,In_478,In_365);
and U771 (N_771,In_290,In_497);
or U772 (N_772,In_526,In_723);
nor U773 (N_773,In_296,In_411);
and U774 (N_774,In_739,In_728);
or U775 (N_775,In_332,In_84);
or U776 (N_776,In_407,In_382);
and U777 (N_777,In_425,In_61);
and U778 (N_778,In_329,In_283);
and U779 (N_779,In_42,In_254);
or U780 (N_780,In_52,In_409);
or U781 (N_781,In_190,In_448);
xor U782 (N_782,In_523,In_171);
or U783 (N_783,In_458,In_647);
and U784 (N_784,In_717,In_12);
nor U785 (N_785,In_582,In_556);
nand U786 (N_786,In_98,In_720);
nand U787 (N_787,In_303,In_405);
and U788 (N_788,In_95,In_267);
nand U789 (N_789,In_321,In_153);
nand U790 (N_790,In_581,In_568);
nor U791 (N_791,In_681,In_708);
and U792 (N_792,In_310,In_10);
nand U793 (N_793,In_694,In_550);
nor U794 (N_794,In_283,In_693);
and U795 (N_795,In_576,In_513);
or U796 (N_796,In_47,In_72);
xor U797 (N_797,In_95,In_695);
nor U798 (N_798,In_265,In_636);
and U799 (N_799,In_29,In_730);
and U800 (N_800,In_523,In_701);
xor U801 (N_801,In_740,In_353);
and U802 (N_802,In_487,In_252);
xnor U803 (N_803,In_694,In_269);
or U804 (N_804,In_267,In_442);
nor U805 (N_805,In_30,In_221);
xnor U806 (N_806,In_497,In_278);
nand U807 (N_807,In_224,In_45);
or U808 (N_808,In_495,In_663);
or U809 (N_809,In_655,In_745);
nor U810 (N_810,In_243,In_275);
xnor U811 (N_811,In_630,In_158);
and U812 (N_812,In_122,In_107);
or U813 (N_813,In_316,In_296);
nand U814 (N_814,In_442,In_139);
nand U815 (N_815,In_533,In_523);
nand U816 (N_816,In_528,In_439);
nor U817 (N_817,In_707,In_33);
or U818 (N_818,In_308,In_130);
or U819 (N_819,In_221,In_204);
nand U820 (N_820,In_186,In_310);
nor U821 (N_821,In_2,In_438);
and U822 (N_822,In_32,In_609);
nand U823 (N_823,In_699,In_391);
xnor U824 (N_824,In_736,In_92);
and U825 (N_825,In_334,In_683);
or U826 (N_826,In_487,In_154);
nor U827 (N_827,In_707,In_284);
nand U828 (N_828,In_381,In_544);
and U829 (N_829,In_732,In_181);
or U830 (N_830,In_1,In_512);
and U831 (N_831,In_562,In_169);
nor U832 (N_832,In_48,In_695);
xnor U833 (N_833,In_582,In_142);
and U834 (N_834,In_415,In_725);
nor U835 (N_835,In_477,In_488);
xor U836 (N_836,In_172,In_530);
xor U837 (N_837,In_451,In_711);
and U838 (N_838,In_194,In_32);
nand U839 (N_839,In_270,In_238);
nand U840 (N_840,In_468,In_663);
nand U841 (N_841,In_303,In_327);
nor U842 (N_842,In_552,In_633);
and U843 (N_843,In_44,In_241);
and U844 (N_844,In_439,In_366);
nor U845 (N_845,In_647,In_425);
xor U846 (N_846,In_275,In_579);
nor U847 (N_847,In_653,In_623);
nor U848 (N_848,In_189,In_214);
or U849 (N_849,In_145,In_736);
and U850 (N_850,In_720,In_730);
nand U851 (N_851,In_593,In_317);
nand U852 (N_852,In_658,In_672);
xnor U853 (N_853,In_716,In_467);
xnor U854 (N_854,In_507,In_623);
nor U855 (N_855,In_262,In_154);
or U856 (N_856,In_448,In_404);
and U857 (N_857,In_122,In_392);
or U858 (N_858,In_147,In_598);
nand U859 (N_859,In_45,In_242);
nor U860 (N_860,In_742,In_418);
and U861 (N_861,In_371,In_330);
nand U862 (N_862,In_136,In_484);
and U863 (N_863,In_565,In_423);
or U864 (N_864,In_286,In_116);
or U865 (N_865,In_337,In_335);
or U866 (N_866,In_294,In_207);
xor U867 (N_867,In_146,In_531);
xor U868 (N_868,In_650,In_71);
or U869 (N_869,In_165,In_22);
nor U870 (N_870,In_67,In_646);
or U871 (N_871,In_21,In_734);
nand U872 (N_872,In_248,In_734);
nor U873 (N_873,In_94,In_202);
and U874 (N_874,In_141,In_43);
and U875 (N_875,In_703,In_380);
and U876 (N_876,In_649,In_91);
nand U877 (N_877,In_147,In_705);
xor U878 (N_878,In_198,In_235);
or U879 (N_879,In_108,In_637);
and U880 (N_880,In_137,In_413);
nand U881 (N_881,In_328,In_576);
xor U882 (N_882,In_190,In_615);
nand U883 (N_883,In_726,In_58);
nand U884 (N_884,In_77,In_635);
nor U885 (N_885,In_423,In_392);
or U886 (N_886,In_318,In_719);
and U887 (N_887,In_124,In_323);
and U888 (N_888,In_469,In_346);
and U889 (N_889,In_17,In_676);
and U890 (N_890,In_298,In_107);
nor U891 (N_891,In_375,In_243);
nor U892 (N_892,In_749,In_480);
or U893 (N_893,In_630,In_514);
nand U894 (N_894,In_28,In_521);
xor U895 (N_895,In_71,In_522);
nand U896 (N_896,In_270,In_622);
xnor U897 (N_897,In_38,In_723);
or U898 (N_898,In_61,In_747);
or U899 (N_899,In_316,In_55);
and U900 (N_900,In_510,In_572);
nor U901 (N_901,In_353,In_718);
and U902 (N_902,In_345,In_274);
or U903 (N_903,In_697,In_691);
xor U904 (N_904,In_732,In_693);
nand U905 (N_905,In_483,In_552);
or U906 (N_906,In_416,In_398);
xnor U907 (N_907,In_587,In_192);
nor U908 (N_908,In_392,In_152);
and U909 (N_909,In_266,In_77);
xnor U910 (N_910,In_341,In_606);
and U911 (N_911,In_413,In_364);
and U912 (N_912,In_205,In_570);
or U913 (N_913,In_47,In_721);
xnor U914 (N_914,In_720,In_401);
and U915 (N_915,In_621,In_432);
and U916 (N_916,In_507,In_299);
or U917 (N_917,In_121,In_581);
nand U918 (N_918,In_625,In_245);
and U919 (N_919,In_36,In_591);
nor U920 (N_920,In_366,In_448);
nand U921 (N_921,In_345,In_647);
nor U922 (N_922,In_341,In_23);
xor U923 (N_923,In_682,In_649);
or U924 (N_924,In_346,In_622);
nand U925 (N_925,In_546,In_358);
and U926 (N_926,In_607,In_278);
or U927 (N_927,In_422,In_328);
nor U928 (N_928,In_366,In_485);
xnor U929 (N_929,In_481,In_231);
or U930 (N_930,In_591,In_202);
nand U931 (N_931,In_126,In_731);
nor U932 (N_932,In_172,In_270);
or U933 (N_933,In_704,In_668);
nand U934 (N_934,In_207,In_494);
or U935 (N_935,In_56,In_66);
nand U936 (N_936,In_468,In_477);
nor U937 (N_937,In_691,In_335);
and U938 (N_938,In_257,In_426);
xor U939 (N_939,In_527,In_706);
or U940 (N_940,In_713,In_685);
nor U941 (N_941,In_258,In_650);
xnor U942 (N_942,In_670,In_315);
nand U943 (N_943,In_340,In_184);
nand U944 (N_944,In_409,In_49);
nor U945 (N_945,In_564,In_563);
or U946 (N_946,In_27,In_531);
nand U947 (N_947,In_492,In_92);
nor U948 (N_948,In_634,In_687);
xnor U949 (N_949,In_345,In_609);
nor U950 (N_950,In_164,In_338);
nand U951 (N_951,In_470,In_729);
and U952 (N_952,In_211,In_231);
nor U953 (N_953,In_142,In_35);
nor U954 (N_954,In_329,In_501);
xnor U955 (N_955,In_427,In_611);
nor U956 (N_956,In_554,In_38);
and U957 (N_957,In_483,In_16);
or U958 (N_958,In_378,In_496);
and U959 (N_959,In_189,In_429);
nor U960 (N_960,In_434,In_721);
or U961 (N_961,In_568,In_723);
nand U962 (N_962,In_248,In_244);
nor U963 (N_963,In_493,In_392);
nor U964 (N_964,In_459,In_52);
or U965 (N_965,In_653,In_116);
nand U966 (N_966,In_399,In_744);
nand U967 (N_967,In_629,In_300);
and U968 (N_968,In_402,In_9);
or U969 (N_969,In_394,In_278);
xnor U970 (N_970,In_560,In_357);
and U971 (N_971,In_516,In_582);
nand U972 (N_972,In_142,In_662);
or U973 (N_973,In_485,In_478);
xnor U974 (N_974,In_179,In_745);
xnor U975 (N_975,In_415,In_613);
and U976 (N_976,In_190,In_495);
or U977 (N_977,In_299,In_394);
xnor U978 (N_978,In_265,In_304);
or U979 (N_979,In_493,In_691);
nor U980 (N_980,In_626,In_108);
xnor U981 (N_981,In_331,In_664);
and U982 (N_982,In_286,In_415);
and U983 (N_983,In_433,In_465);
xor U984 (N_984,In_410,In_194);
nor U985 (N_985,In_655,In_82);
and U986 (N_986,In_416,In_334);
nand U987 (N_987,In_336,In_324);
nand U988 (N_988,In_543,In_568);
xnor U989 (N_989,In_329,In_586);
or U990 (N_990,In_568,In_122);
or U991 (N_991,In_81,In_332);
and U992 (N_992,In_712,In_527);
nand U993 (N_993,In_475,In_697);
or U994 (N_994,In_464,In_44);
nor U995 (N_995,In_166,In_172);
and U996 (N_996,In_737,In_196);
nor U997 (N_997,In_734,In_748);
or U998 (N_998,In_645,In_61);
and U999 (N_999,In_320,In_317);
nor U1000 (N_1000,N_59,N_413);
xnor U1001 (N_1001,N_664,N_426);
nor U1002 (N_1002,N_670,N_706);
nor U1003 (N_1003,N_779,N_209);
nor U1004 (N_1004,N_283,N_720);
nor U1005 (N_1005,N_95,N_963);
and U1006 (N_1006,N_399,N_889);
xor U1007 (N_1007,N_571,N_648);
nand U1008 (N_1008,N_660,N_324);
xnor U1009 (N_1009,N_338,N_469);
nand U1010 (N_1010,N_654,N_38);
nor U1011 (N_1011,N_113,N_255);
and U1012 (N_1012,N_888,N_274);
nand U1013 (N_1013,N_750,N_611);
or U1014 (N_1014,N_176,N_980);
nor U1015 (N_1015,N_277,N_144);
nand U1016 (N_1016,N_60,N_160);
nand U1017 (N_1017,N_441,N_987);
nor U1018 (N_1018,N_314,N_690);
nand U1019 (N_1019,N_710,N_61);
nand U1020 (N_1020,N_813,N_728);
nand U1021 (N_1021,N_610,N_993);
or U1022 (N_1022,N_178,N_18);
xor U1023 (N_1023,N_535,N_336);
xnor U1024 (N_1024,N_492,N_446);
xnor U1025 (N_1025,N_74,N_206);
and U1026 (N_1026,N_186,N_663);
and U1027 (N_1027,N_164,N_444);
nor U1028 (N_1028,N_222,N_879);
nor U1029 (N_1029,N_581,N_536);
and U1030 (N_1030,N_190,N_622);
nor U1031 (N_1031,N_935,N_912);
and U1032 (N_1032,N_604,N_613);
or U1033 (N_1033,N_311,N_133);
nand U1034 (N_1034,N_337,N_383);
xor U1035 (N_1035,N_600,N_135);
or U1036 (N_1036,N_104,N_851);
or U1037 (N_1037,N_293,N_842);
or U1038 (N_1038,N_681,N_325);
xnor U1039 (N_1039,N_515,N_394);
and U1040 (N_1040,N_601,N_758);
or U1041 (N_1041,N_697,N_519);
nand U1042 (N_1042,N_726,N_708);
xor U1043 (N_1043,N_675,N_530);
or U1044 (N_1044,N_19,N_162);
and U1045 (N_1045,N_86,N_915);
or U1046 (N_1046,N_943,N_470);
xnor U1047 (N_1047,N_11,N_953);
or U1048 (N_1048,N_572,N_579);
nand U1049 (N_1049,N_983,N_916);
or U1050 (N_1050,N_696,N_353);
or U1051 (N_1051,N_557,N_478);
xnor U1052 (N_1052,N_339,N_724);
nor U1053 (N_1053,N_958,N_374);
nand U1054 (N_1054,N_440,N_810);
xnor U1055 (N_1055,N_553,N_296);
or U1056 (N_1056,N_34,N_508);
nand U1057 (N_1057,N_168,N_674);
or U1058 (N_1058,N_29,N_84);
xnor U1059 (N_1059,N_533,N_804);
nor U1060 (N_1060,N_518,N_873);
xnor U1061 (N_1061,N_629,N_420);
and U1062 (N_1062,N_619,N_31);
and U1063 (N_1063,N_636,N_850);
nor U1064 (N_1064,N_445,N_678);
nor U1065 (N_1065,N_302,N_717);
and U1066 (N_1066,N_735,N_177);
or U1067 (N_1067,N_20,N_33);
xor U1068 (N_1068,N_925,N_656);
nand U1069 (N_1069,N_514,N_752);
xor U1070 (N_1070,N_2,N_407);
and U1071 (N_1071,N_844,N_884);
nor U1072 (N_1072,N_94,N_303);
or U1073 (N_1073,N_942,N_409);
or U1074 (N_1074,N_560,N_590);
and U1075 (N_1075,N_68,N_385);
or U1076 (N_1076,N_340,N_567);
xor U1077 (N_1077,N_364,N_323);
nand U1078 (N_1078,N_658,N_711);
or U1079 (N_1079,N_1,N_753);
and U1080 (N_1080,N_286,N_791);
or U1081 (N_1081,N_241,N_695);
or U1082 (N_1082,N_300,N_807);
nor U1083 (N_1083,N_513,N_712);
nor U1084 (N_1084,N_173,N_854);
or U1085 (N_1085,N_92,N_734);
nor U1086 (N_1086,N_98,N_891);
nand U1087 (N_1087,N_782,N_527);
xor U1088 (N_1088,N_718,N_580);
and U1089 (N_1089,N_9,N_281);
nor U1090 (N_1090,N_438,N_150);
xor U1091 (N_1091,N_995,N_673);
nand U1092 (N_1092,N_877,N_269);
nor U1093 (N_1093,N_192,N_398);
and U1094 (N_1094,N_827,N_384);
nand U1095 (N_1095,N_974,N_727);
nor U1096 (N_1096,N_745,N_795);
nor U1097 (N_1097,N_459,N_39);
nand U1098 (N_1098,N_465,N_76);
and U1099 (N_1099,N_0,N_165);
or U1100 (N_1100,N_202,N_56);
nor U1101 (N_1101,N_218,N_549);
nor U1102 (N_1102,N_297,N_531);
and U1103 (N_1103,N_126,N_432);
nor U1104 (N_1104,N_411,N_460);
nand U1105 (N_1105,N_332,N_883);
or U1106 (N_1106,N_285,N_327);
and U1107 (N_1107,N_537,N_351);
and U1108 (N_1108,N_331,N_228);
nand U1109 (N_1109,N_627,N_917);
or U1110 (N_1110,N_573,N_748);
and U1111 (N_1111,N_227,N_990);
or U1112 (N_1112,N_387,N_45);
xnor U1113 (N_1113,N_644,N_510);
nor U1114 (N_1114,N_404,N_174);
nand U1115 (N_1115,N_544,N_333);
nand U1116 (N_1116,N_418,N_456);
nand U1117 (N_1117,N_52,N_180);
and U1118 (N_1118,N_668,N_511);
xor U1119 (N_1119,N_941,N_731);
and U1120 (N_1120,N_175,N_947);
xor U1121 (N_1121,N_266,N_365);
or U1122 (N_1122,N_522,N_871);
and U1123 (N_1123,N_170,N_217);
xor U1124 (N_1124,N_908,N_280);
and U1125 (N_1125,N_767,N_632);
or U1126 (N_1126,N_251,N_204);
and U1127 (N_1127,N_761,N_906);
and U1128 (N_1128,N_732,N_262);
and U1129 (N_1129,N_306,N_985);
nor U1130 (N_1130,N_65,N_248);
xnor U1131 (N_1131,N_815,N_652);
xnor U1132 (N_1132,N_903,N_819);
nand U1133 (N_1133,N_959,N_812);
or U1134 (N_1134,N_584,N_477);
nand U1135 (N_1135,N_714,N_754);
or U1136 (N_1136,N_263,N_253);
or U1137 (N_1137,N_7,N_973);
or U1138 (N_1138,N_372,N_642);
and U1139 (N_1139,N_777,N_647);
and U1140 (N_1140,N_319,N_49);
nor U1141 (N_1141,N_99,N_342);
nor U1142 (N_1142,N_450,N_876);
and U1143 (N_1143,N_775,N_747);
and U1144 (N_1144,N_121,N_243);
xor U1145 (N_1145,N_53,N_163);
xnor U1146 (N_1146,N_79,N_833);
nor U1147 (N_1147,N_907,N_811);
or U1148 (N_1148,N_396,N_605);
xor U1149 (N_1149,N_541,N_631);
nor U1150 (N_1150,N_866,N_780);
and U1151 (N_1151,N_785,N_483);
and U1152 (N_1152,N_455,N_984);
or U1153 (N_1153,N_434,N_586);
nand U1154 (N_1154,N_474,N_725);
xnor U1155 (N_1155,N_578,N_181);
or U1156 (N_1156,N_479,N_899);
or U1157 (N_1157,N_591,N_628);
nand U1158 (N_1158,N_85,N_161);
nand U1159 (N_1159,N_298,N_152);
nor U1160 (N_1160,N_41,N_361);
and U1161 (N_1161,N_880,N_901);
or U1162 (N_1162,N_13,N_645);
and U1163 (N_1163,N_881,N_910);
or U1164 (N_1164,N_329,N_313);
nand U1165 (N_1165,N_582,N_288);
xor U1166 (N_1166,N_259,N_921);
nor U1167 (N_1167,N_539,N_26);
and U1168 (N_1168,N_603,N_597);
nor U1169 (N_1169,N_58,N_258);
or U1170 (N_1170,N_97,N_436);
nand U1171 (N_1171,N_719,N_615);
xor U1172 (N_1172,N_207,N_978);
xor U1173 (N_1173,N_198,N_408);
nand U1174 (N_1174,N_229,N_766);
nor U1175 (N_1175,N_834,N_992);
nand U1176 (N_1176,N_713,N_491);
xor U1177 (N_1177,N_828,N_986);
nor U1178 (N_1178,N_989,N_760);
xnor U1179 (N_1179,N_556,N_27);
or U1180 (N_1180,N_278,N_172);
or U1181 (N_1181,N_742,N_158);
xor U1182 (N_1182,N_382,N_471);
and U1183 (N_1183,N_952,N_142);
nand U1184 (N_1184,N_141,N_389);
xor U1185 (N_1185,N_505,N_356);
and U1186 (N_1186,N_183,N_816);
xnor U1187 (N_1187,N_729,N_12);
and U1188 (N_1188,N_516,N_704);
xnor U1189 (N_1189,N_669,N_448);
and U1190 (N_1190,N_683,N_321);
and U1191 (N_1191,N_44,N_151);
xnor U1192 (N_1192,N_830,N_381);
and U1193 (N_1193,N_562,N_215);
and U1194 (N_1194,N_310,N_359);
nand U1195 (N_1195,N_81,N_860);
or U1196 (N_1196,N_265,N_156);
and U1197 (N_1197,N_100,N_929);
nand U1198 (N_1198,N_837,N_651);
or U1199 (N_1199,N_494,N_268);
nand U1200 (N_1200,N_938,N_246);
xor U1201 (N_1201,N_223,N_517);
and U1202 (N_1202,N_132,N_96);
xnor U1203 (N_1203,N_894,N_540);
xnor U1204 (N_1204,N_721,N_368);
and U1205 (N_1205,N_415,N_312);
or U1206 (N_1206,N_657,N_504);
and U1207 (N_1207,N_275,N_946);
nand U1208 (N_1208,N_405,N_352);
nand U1209 (N_1209,N_334,N_525);
or U1210 (N_1210,N_256,N_427);
xnor U1211 (N_1211,N_521,N_898);
or U1212 (N_1212,N_242,N_191);
nand U1213 (N_1213,N_490,N_107);
nand U1214 (N_1214,N_488,N_464);
nor U1215 (N_1215,N_762,N_765);
xnor U1216 (N_1216,N_50,N_808);
nand U1217 (N_1217,N_127,N_451);
and U1218 (N_1218,N_264,N_686);
xor U1219 (N_1219,N_78,N_787);
and U1220 (N_1220,N_634,N_927);
xor U1221 (N_1221,N_252,N_933);
nand U1222 (N_1222,N_185,N_892);
or U1223 (N_1223,N_679,N_838);
xor U1224 (N_1224,N_902,N_140);
or U1225 (N_1225,N_292,N_272);
xor U1226 (N_1226,N_981,N_284);
and U1227 (N_1227,N_260,N_406);
and U1228 (N_1228,N_70,N_937);
nor U1229 (N_1229,N_360,N_424);
or U1230 (N_1230,N_857,N_497);
and U1231 (N_1231,N_672,N_369);
xor U1232 (N_1232,N_769,N_676);
or U1233 (N_1233,N_467,N_211);
xnor U1234 (N_1234,N_196,N_184);
nand U1235 (N_1235,N_3,N_22);
xnor U1236 (N_1236,N_143,N_349);
and U1237 (N_1237,N_994,N_570);
nor U1238 (N_1238,N_370,N_878);
nor U1239 (N_1239,N_410,N_920);
xnor U1240 (N_1240,N_437,N_821);
and U1241 (N_1241,N_130,N_194);
xnor U1242 (N_1242,N_110,N_40);
and U1243 (N_1243,N_738,N_125);
nand U1244 (N_1244,N_435,N_638);
or U1245 (N_1245,N_709,N_646);
or U1246 (N_1246,N_520,N_773);
nand U1247 (N_1247,N_790,N_225);
or U1248 (N_1248,N_57,N_796);
and U1249 (N_1249,N_829,N_179);
xor U1250 (N_1250,N_962,N_749);
nor U1251 (N_1251,N_169,N_805);
xor U1252 (N_1252,N_764,N_118);
or U1253 (N_1253,N_358,N_665);
nand U1254 (N_1254,N_392,N_997);
and U1255 (N_1255,N_393,N_730);
and U1256 (N_1256,N_524,N_171);
or U1257 (N_1257,N_203,N_476);
xor U1258 (N_1258,N_320,N_793);
nor U1259 (N_1259,N_979,N_345);
and U1260 (N_1260,N_37,N_309);
xor U1261 (N_1261,N_220,N_124);
nand U1262 (N_1262,N_378,N_774);
nand U1263 (N_1263,N_969,N_188);
and U1264 (N_1264,N_928,N_823);
nand U1265 (N_1265,N_101,N_803);
or U1266 (N_1266,N_569,N_443);
and U1267 (N_1267,N_403,N_201);
or U1268 (N_1268,N_155,N_367);
and U1269 (N_1269,N_195,N_271);
or U1270 (N_1270,N_700,N_976);
xnor U1271 (N_1271,N_48,N_818);
or U1272 (N_1272,N_341,N_214);
xnor U1273 (N_1273,N_498,N_346);
and U1274 (N_1274,N_301,N_347);
nand U1275 (N_1275,N_452,N_453);
xor U1276 (N_1276,N_481,N_786);
and U1277 (N_1277,N_400,N_131);
xnor U1278 (N_1278,N_391,N_563);
or U1279 (N_1279,N_576,N_28);
nand U1280 (N_1280,N_967,N_14);
nor U1281 (N_1281,N_90,N_166);
and U1282 (N_1282,N_956,N_875);
nor U1283 (N_1283,N_565,N_354);
and U1284 (N_1284,N_972,N_932);
and U1285 (N_1285,N_473,N_957);
or U1286 (N_1286,N_267,N_982);
xnor U1287 (N_1287,N_841,N_955);
and U1288 (N_1288,N_134,N_608);
xnor U1289 (N_1289,N_236,N_197);
nor U1290 (N_1290,N_149,N_858);
xor U1291 (N_1291,N_547,N_468);
xor U1292 (N_1292,N_139,N_503);
nor U1293 (N_1293,N_988,N_970);
nand U1294 (N_1294,N_30,N_315);
nor U1295 (N_1295,N_395,N_111);
nand U1296 (N_1296,N_421,N_254);
and U1297 (N_1297,N_864,N_826);
xnor U1298 (N_1298,N_677,N_751);
nand U1299 (N_1299,N_123,N_89);
or U1300 (N_1300,N_689,N_363);
xnor U1301 (N_1301,N_51,N_47);
and U1302 (N_1302,N_493,N_846);
nor U1303 (N_1303,N_495,N_276);
or U1304 (N_1304,N_950,N_546);
nor U1305 (N_1305,N_755,N_216);
nor U1306 (N_1306,N_845,N_423);
nor U1307 (N_1307,N_335,N_386);
or U1308 (N_1308,N_189,N_430);
or U1309 (N_1309,N_736,N_897);
xor U1310 (N_1310,N_966,N_233);
and U1311 (N_1311,N_120,N_794);
nand U1312 (N_1312,N_602,N_287);
or U1313 (N_1313,N_388,N_317);
xor U1314 (N_1314,N_614,N_523);
xnor U1315 (N_1315,N_832,N_73);
nand U1316 (N_1316,N_620,N_893);
nand U1317 (N_1317,N_77,N_799);
xnor U1318 (N_1318,N_859,N_763);
xnor U1319 (N_1319,N_357,N_487);
and U1320 (N_1320,N_862,N_671);
or U1321 (N_1321,N_716,N_759);
nor U1322 (N_1322,N_931,N_741);
or U1323 (N_1323,N_330,N_270);
and U1324 (N_1324,N_555,N_63);
xnor U1325 (N_1325,N_655,N_653);
nand U1326 (N_1326,N_509,N_737);
nand U1327 (N_1327,N_362,N_699);
and U1328 (N_1328,N_103,N_273);
xor U1329 (N_1329,N_35,N_934);
nand U1330 (N_1330,N_526,N_500);
or U1331 (N_1331,N_853,N_305);
or U1332 (N_1332,N_538,N_688);
or U1333 (N_1333,N_626,N_789);
xnor U1334 (N_1334,N_15,N_756);
and U1335 (N_1335,N_948,N_461);
nand U1336 (N_1336,N_472,N_598);
nand U1337 (N_1337,N_375,N_788);
and U1338 (N_1338,N_219,N_643);
nor U1339 (N_1339,N_114,N_93);
xor U1340 (N_1340,N_776,N_146);
or U1341 (N_1341,N_566,N_801);
nor U1342 (N_1342,N_422,N_109);
or U1343 (N_1343,N_623,N_945);
and U1344 (N_1344,N_824,N_116);
nand U1345 (N_1345,N_744,N_588);
and U1346 (N_1346,N_852,N_739);
and U1347 (N_1347,N_905,N_817);
nand U1348 (N_1348,N_157,N_640);
nand U1349 (N_1349,N_621,N_757);
xnor U1350 (N_1350,N_802,N_25);
or U1351 (N_1351,N_914,N_102);
nor U1352 (N_1352,N_856,N_502);
xor U1353 (N_1353,N_849,N_24);
and U1354 (N_1354,N_691,N_442);
and U1355 (N_1355,N_783,N_507);
nor U1356 (N_1356,N_304,N_199);
and U1357 (N_1357,N_746,N_294);
nor U1358 (N_1358,N_554,N_159);
nor U1359 (N_1359,N_454,N_390);
xnor U1360 (N_1360,N_609,N_182);
nor U1361 (N_1361,N_715,N_904);
xnor U1362 (N_1362,N_639,N_869);
and U1363 (N_1363,N_318,N_863);
and U1364 (N_1364,N_705,N_592);
and U1365 (N_1365,N_698,N_583);
or U1366 (N_1366,N_944,N_212);
nand U1367 (N_1367,N_42,N_112);
xnor U1368 (N_1368,N_213,N_308);
or U1369 (N_1369,N_128,N_900);
xnor U1370 (N_1370,N_193,N_373);
and U1371 (N_1371,N_295,N_496);
and U1372 (N_1372,N_882,N_240);
nand U1373 (N_1373,N_230,N_247);
or U1374 (N_1374,N_564,N_949);
nor U1375 (N_1375,N_326,N_380);
or U1376 (N_1376,N_244,N_599);
and U1377 (N_1377,N_91,N_806);
and U1378 (N_1378,N_210,N_299);
nor U1379 (N_1379,N_624,N_153);
nor U1380 (N_1380,N_106,N_83);
or U1381 (N_1381,N_419,N_350);
or U1382 (N_1382,N_328,N_148);
or U1383 (N_1383,N_659,N_397);
nand U1384 (N_1384,N_772,N_551);
xnor U1385 (N_1385,N_770,N_66);
nor U1386 (N_1386,N_4,N_250);
and U1387 (N_1387,N_625,N_589);
xor U1388 (N_1388,N_23,N_896);
nand U1389 (N_1389,N_552,N_307);
and U1390 (N_1390,N_743,N_482);
nand U1391 (N_1391,N_798,N_200);
nand U1392 (N_1392,N_480,N_80);
and U1393 (N_1393,N_122,N_62);
and U1394 (N_1394,N_475,N_684);
or U1395 (N_1395,N_618,N_996);
xnor U1396 (N_1396,N_371,N_792);
and U1397 (N_1397,N_137,N_72);
nor U1398 (N_1398,N_376,N_800);
nor U1399 (N_1399,N_701,N_617);
nor U1400 (N_1400,N_861,N_187);
xor U1401 (N_1401,N_630,N_88);
xnor U1402 (N_1402,N_208,N_685);
nor U1403 (N_1403,N_936,N_633);
nand U1404 (N_1404,N_797,N_577);
nand U1405 (N_1405,N_587,N_909);
xor U1406 (N_1406,N_105,N_940);
nor U1407 (N_1407,N_666,N_412);
xnor U1408 (N_1408,N_872,N_784);
nor U1409 (N_1409,N_108,N_82);
xor U1410 (N_1410,N_650,N_954);
nor U1411 (N_1411,N_528,N_887);
nand U1412 (N_1412,N_585,N_449);
and U1413 (N_1413,N_291,N_596);
xnor U1414 (N_1414,N_489,N_707);
nand U1415 (N_1415,N_235,N_692);
nand U1416 (N_1416,N_506,N_316);
nor U1417 (N_1417,N_238,N_21);
nand U1418 (N_1418,N_594,N_855);
nand U1419 (N_1419,N_971,N_568);
nor U1420 (N_1420,N_667,N_612);
and U1421 (N_1421,N_550,N_417);
nand U1422 (N_1422,N_17,N_379);
nor U1423 (N_1423,N_64,N_723);
nor U1424 (N_1424,N_54,N_224);
nand U1425 (N_1425,N_843,N_279);
xnor U1426 (N_1426,N_960,N_913);
and U1427 (N_1427,N_43,N_662);
xor U1428 (N_1428,N_534,N_485);
nand U1429 (N_1429,N_433,N_975);
nand U1430 (N_1430,N_693,N_694);
nor U1431 (N_1431,N_484,N_348);
xnor U1432 (N_1432,N_366,N_428);
nand U1433 (N_1433,N_249,N_635);
and U1434 (N_1434,N_138,N_922);
xor U1435 (N_1435,N_847,N_416);
and U1436 (N_1436,N_680,N_814);
xor U1437 (N_1437,N_768,N_414);
nor U1438 (N_1438,N_740,N_778);
nor U1439 (N_1439,N_67,N_8);
nand U1440 (N_1440,N_951,N_835);
or U1441 (N_1441,N_221,N_661);
nand U1442 (N_1442,N_848,N_911);
and U1443 (N_1443,N_607,N_926);
xor U1444 (N_1444,N_239,N_71);
and U1445 (N_1445,N_687,N_559);
nand U1446 (N_1446,N_119,N_574);
nor U1447 (N_1447,N_512,N_5);
xnor U1448 (N_1448,N_10,N_532);
xnor U1449 (N_1449,N_575,N_865);
or U1450 (N_1450,N_542,N_282);
or U1451 (N_1451,N_154,N_839);
nor U1452 (N_1452,N_402,N_377);
or U1453 (N_1453,N_840,N_75);
or U1454 (N_1454,N_289,N_702);
xor U1455 (N_1455,N_447,N_991);
xnor U1456 (N_1456,N_401,N_930);
or U1457 (N_1457,N_939,N_593);
and U1458 (N_1458,N_237,N_595);
and U1459 (N_1459,N_344,N_234);
nor U1460 (N_1460,N_998,N_458);
nor U1461 (N_1461,N_964,N_868);
xor U1462 (N_1462,N_771,N_343);
xor U1463 (N_1463,N_977,N_867);
nor U1464 (N_1464,N_129,N_890);
and U1465 (N_1465,N_809,N_69);
or U1466 (N_1466,N_703,N_147);
or U1467 (N_1467,N_425,N_355);
nor U1468 (N_1468,N_261,N_733);
or U1469 (N_1469,N_36,N_924);
xor U1470 (N_1470,N_722,N_545);
nor U1471 (N_1471,N_486,N_46);
nor U1472 (N_1472,N_463,N_439);
or U1473 (N_1473,N_999,N_637);
nand U1474 (N_1474,N_87,N_895);
or U1475 (N_1475,N_499,N_885);
nand U1476 (N_1476,N_548,N_616);
nand U1477 (N_1477,N_145,N_466);
and U1478 (N_1478,N_961,N_501);
nor U1479 (N_1479,N_918,N_641);
xor U1480 (N_1480,N_886,N_822);
nor U1481 (N_1481,N_781,N_820);
or U1482 (N_1482,N_429,N_55);
or U1483 (N_1483,N_32,N_606);
xor U1484 (N_1484,N_874,N_431);
nor U1485 (N_1485,N_923,N_870);
or U1486 (N_1486,N_919,N_462);
or U1487 (N_1487,N_831,N_167);
or U1488 (N_1488,N_257,N_836);
or U1489 (N_1489,N_205,N_965);
or U1490 (N_1490,N_245,N_322);
nand U1491 (N_1491,N_529,N_457);
or U1492 (N_1492,N_543,N_231);
nor U1493 (N_1493,N_136,N_115);
nand U1494 (N_1494,N_290,N_16);
and U1495 (N_1495,N_226,N_561);
and U1496 (N_1496,N_232,N_682);
and U1497 (N_1497,N_558,N_649);
and U1498 (N_1498,N_117,N_6);
xnor U1499 (N_1499,N_968,N_825);
nor U1500 (N_1500,N_90,N_175);
and U1501 (N_1501,N_36,N_329);
nand U1502 (N_1502,N_715,N_864);
nand U1503 (N_1503,N_632,N_105);
nor U1504 (N_1504,N_378,N_277);
nor U1505 (N_1505,N_94,N_484);
and U1506 (N_1506,N_283,N_934);
xor U1507 (N_1507,N_568,N_694);
nand U1508 (N_1508,N_990,N_353);
xnor U1509 (N_1509,N_37,N_392);
or U1510 (N_1510,N_727,N_754);
nand U1511 (N_1511,N_619,N_230);
xor U1512 (N_1512,N_876,N_702);
and U1513 (N_1513,N_277,N_386);
xor U1514 (N_1514,N_218,N_753);
and U1515 (N_1515,N_377,N_673);
and U1516 (N_1516,N_813,N_460);
nand U1517 (N_1517,N_239,N_8);
xnor U1518 (N_1518,N_433,N_599);
xor U1519 (N_1519,N_726,N_547);
nor U1520 (N_1520,N_649,N_521);
nand U1521 (N_1521,N_721,N_132);
xor U1522 (N_1522,N_109,N_314);
nand U1523 (N_1523,N_942,N_687);
nand U1524 (N_1524,N_952,N_413);
xor U1525 (N_1525,N_539,N_837);
nor U1526 (N_1526,N_271,N_0);
and U1527 (N_1527,N_107,N_278);
nand U1528 (N_1528,N_120,N_733);
nand U1529 (N_1529,N_809,N_422);
and U1530 (N_1530,N_763,N_44);
or U1531 (N_1531,N_867,N_289);
and U1532 (N_1532,N_705,N_570);
xor U1533 (N_1533,N_812,N_45);
nor U1534 (N_1534,N_778,N_972);
nor U1535 (N_1535,N_441,N_742);
nor U1536 (N_1536,N_806,N_140);
nor U1537 (N_1537,N_662,N_524);
or U1538 (N_1538,N_37,N_711);
nor U1539 (N_1539,N_521,N_614);
nor U1540 (N_1540,N_542,N_277);
nor U1541 (N_1541,N_673,N_299);
and U1542 (N_1542,N_590,N_647);
xnor U1543 (N_1543,N_506,N_660);
nand U1544 (N_1544,N_948,N_155);
xnor U1545 (N_1545,N_842,N_9);
and U1546 (N_1546,N_311,N_251);
nor U1547 (N_1547,N_149,N_244);
xnor U1548 (N_1548,N_337,N_94);
or U1549 (N_1549,N_598,N_418);
and U1550 (N_1550,N_780,N_577);
and U1551 (N_1551,N_565,N_834);
nand U1552 (N_1552,N_916,N_566);
nor U1553 (N_1553,N_665,N_2);
nand U1554 (N_1554,N_828,N_899);
nor U1555 (N_1555,N_95,N_329);
nand U1556 (N_1556,N_91,N_327);
nor U1557 (N_1557,N_223,N_892);
nand U1558 (N_1558,N_279,N_656);
xnor U1559 (N_1559,N_964,N_386);
xor U1560 (N_1560,N_551,N_670);
and U1561 (N_1561,N_697,N_487);
nor U1562 (N_1562,N_531,N_728);
nand U1563 (N_1563,N_567,N_732);
nand U1564 (N_1564,N_731,N_945);
or U1565 (N_1565,N_769,N_610);
or U1566 (N_1566,N_483,N_582);
nor U1567 (N_1567,N_98,N_291);
and U1568 (N_1568,N_336,N_55);
and U1569 (N_1569,N_414,N_252);
nand U1570 (N_1570,N_92,N_184);
xnor U1571 (N_1571,N_331,N_397);
or U1572 (N_1572,N_355,N_256);
and U1573 (N_1573,N_88,N_351);
or U1574 (N_1574,N_676,N_44);
nand U1575 (N_1575,N_265,N_253);
or U1576 (N_1576,N_894,N_96);
or U1577 (N_1577,N_575,N_605);
nor U1578 (N_1578,N_38,N_957);
xor U1579 (N_1579,N_609,N_107);
and U1580 (N_1580,N_592,N_579);
nor U1581 (N_1581,N_243,N_804);
and U1582 (N_1582,N_630,N_607);
nand U1583 (N_1583,N_214,N_186);
and U1584 (N_1584,N_39,N_249);
nand U1585 (N_1585,N_245,N_232);
or U1586 (N_1586,N_428,N_520);
and U1587 (N_1587,N_389,N_759);
or U1588 (N_1588,N_1,N_24);
nand U1589 (N_1589,N_255,N_353);
and U1590 (N_1590,N_891,N_798);
nand U1591 (N_1591,N_18,N_25);
nor U1592 (N_1592,N_106,N_909);
nor U1593 (N_1593,N_506,N_552);
or U1594 (N_1594,N_946,N_932);
xnor U1595 (N_1595,N_941,N_825);
xor U1596 (N_1596,N_745,N_220);
or U1597 (N_1597,N_480,N_121);
nor U1598 (N_1598,N_847,N_796);
or U1599 (N_1599,N_476,N_473);
nand U1600 (N_1600,N_267,N_846);
or U1601 (N_1601,N_819,N_127);
or U1602 (N_1602,N_562,N_531);
xor U1603 (N_1603,N_678,N_325);
nand U1604 (N_1604,N_437,N_607);
nor U1605 (N_1605,N_744,N_722);
xnor U1606 (N_1606,N_518,N_729);
nor U1607 (N_1607,N_450,N_394);
xnor U1608 (N_1608,N_197,N_996);
nand U1609 (N_1609,N_253,N_726);
and U1610 (N_1610,N_824,N_633);
nand U1611 (N_1611,N_799,N_566);
and U1612 (N_1612,N_754,N_87);
or U1613 (N_1613,N_61,N_50);
or U1614 (N_1614,N_309,N_442);
or U1615 (N_1615,N_548,N_285);
nor U1616 (N_1616,N_378,N_659);
and U1617 (N_1617,N_327,N_565);
nor U1618 (N_1618,N_645,N_244);
nand U1619 (N_1619,N_980,N_69);
or U1620 (N_1620,N_226,N_710);
xnor U1621 (N_1621,N_894,N_566);
or U1622 (N_1622,N_187,N_868);
xnor U1623 (N_1623,N_11,N_607);
xnor U1624 (N_1624,N_476,N_28);
nor U1625 (N_1625,N_437,N_551);
nand U1626 (N_1626,N_764,N_162);
nor U1627 (N_1627,N_609,N_856);
and U1628 (N_1628,N_46,N_919);
xnor U1629 (N_1629,N_301,N_550);
nand U1630 (N_1630,N_494,N_881);
nand U1631 (N_1631,N_976,N_663);
xnor U1632 (N_1632,N_978,N_786);
nand U1633 (N_1633,N_649,N_940);
nor U1634 (N_1634,N_726,N_959);
nor U1635 (N_1635,N_315,N_80);
or U1636 (N_1636,N_864,N_55);
nor U1637 (N_1637,N_252,N_750);
nor U1638 (N_1638,N_915,N_262);
nand U1639 (N_1639,N_725,N_498);
nor U1640 (N_1640,N_235,N_520);
or U1641 (N_1641,N_690,N_329);
nand U1642 (N_1642,N_901,N_205);
xnor U1643 (N_1643,N_618,N_804);
nand U1644 (N_1644,N_463,N_723);
or U1645 (N_1645,N_164,N_435);
or U1646 (N_1646,N_175,N_654);
nor U1647 (N_1647,N_564,N_958);
xnor U1648 (N_1648,N_633,N_726);
or U1649 (N_1649,N_706,N_820);
xor U1650 (N_1650,N_238,N_990);
nor U1651 (N_1651,N_366,N_224);
xor U1652 (N_1652,N_582,N_151);
xor U1653 (N_1653,N_778,N_575);
nor U1654 (N_1654,N_734,N_10);
or U1655 (N_1655,N_357,N_319);
nor U1656 (N_1656,N_332,N_669);
nand U1657 (N_1657,N_779,N_21);
nor U1658 (N_1658,N_889,N_124);
xor U1659 (N_1659,N_227,N_824);
and U1660 (N_1660,N_754,N_353);
xnor U1661 (N_1661,N_967,N_492);
or U1662 (N_1662,N_101,N_306);
nor U1663 (N_1663,N_842,N_496);
xor U1664 (N_1664,N_212,N_723);
or U1665 (N_1665,N_337,N_603);
xor U1666 (N_1666,N_922,N_891);
or U1667 (N_1667,N_599,N_941);
and U1668 (N_1668,N_577,N_112);
and U1669 (N_1669,N_918,N_388);
nand U1670 (N_1670,N_107,N_529);
and U1671 (N_1671,N_277,N_270);
and U1672 (N_1672,N_190,N_691);
or U1673 (N_1673,N_405,N_578);
and U1674 (N_1674,N_969,N_508);
xor U1675 (N_1675,N_357,N_28);
nor U1676 (N_1676,N_619,N_865);
or U1677 (N_1677,N_563,N_148);
nor U1678 (N_1678,N_493,N_87);
and U1679 (N_1679,N_625,N_559);
nand U1680 (N_1680,N_791,N_649);
nand U1681 (N_1681,N_735,N_876);
and U1682 (N_1682,N_752,N_210);
xor U1683 (N_1683,N_838,N_47);
or U1684 (N_1684,N_731,N_890);
and U1685 (N_1685,N_497,N_738);
nor U1686 (N_1686,N_870,N_67);
nand U1687 (N_1687,N_989,N_786);
xnor U1688 (N_1688,N_47,N_257);
or U1689 (N_1689,N_95,N_289);
or U1690 (N_1690,N_369,N_86);
nand U1691 (N_1691,N_404,N_729);
xnor U1692 (N_1692,N_953,N_791);
and U1693 (N_1693,N_922,N_176);
xnor U1694 (N_1694,N_969,N_968);
or U1695 (N_1695,N_752,N_540);
nor U1696 (N_1696,N_798,N_606);
xor U1697 (N_1697,N_623,N_73);
and U1698 (N_1698,N_834,N_923);
and U1699 (N_1699,N_225,N_603);
or U1700 (N_1700,N_164,N_357);
nand U1701 (N_1701,N_231,N_421);
and U1702 (N_1702,N_449,N_498);
and U1703 (N_1703,N_103,N_381);
or U1704 (N_1704,N_944,N_809);
and U1705 (N_1705,N_30,N_979);
xnor U1706 (N_1706,N_810,N_783);
or U1707 (N_1707,N_408,N_382);
xor U1708 (N_1708,N_382,N_956);
xor U1709 (N_1709,N_530,N_32);
or U1710 (N_1710,N_622,N_304);
xor U1711 (N_1711,N_362,N_502);
nor U1712 (N_1712,N_529,N_915);
xor U1713 (N_1713,N_992,N_491);
nand U1714 (N_1714,N_843,N_235);
xnor U1715 (N_1715,N_966,N_529);
xor U1716 (N_1716,N_763,N_19);
nor U1717 (N_1717,N_670,N_649);
and U1718 (N_1718,N_483,N_154);
and U1719 (N_1719,N_26,N_538);
and U1720 (N_1720,N_697,N_912);
or U1721 (N_1721,N_737,N_806);
nand U1722 (N_1722,N_398,N_447);
xnor U1723 (N_1723,N_420,N_52);
or U1724 (N_1724,N_245,N_893);
xnor U1725 (N_1725,N_804,N_895);
nor U1726 (N_1726,N_357,N_47);
nand U1727 (N_1727,N_244,N_676);
or U1728 (N_1728,N_754,N_10);
xor U1729 (N_1729,N_271,N_788);
xnor U1730 (N_1730,N_261,N_226);
xnor U1731 (N_1731,N_578,N_299);
nand U1732 (N_1732,N_236,N_570);
xnor U1733 (N_1733,N_75,N_744);
nor U1734 (N_1734,N_2,N_76);
nand U1735 (N_1735,N_273,N_81);
nand U1736 (N_1736,N_509,N_139);
xor U1737 (N_1737,N_587,N_185);
or U1738 (N_1738,N_499,N_345);
and U1739 (N_1739,N_702,N_861);
or U1740 (N_1740,N_137,N_275);
or U1741 (N_1741,N_493,N_619);
nor U1742 (N_1742,N_414,N_450);
nand U1743 (N_1743,N_172,N_61);
xor U1744 (N_1744,N_373,N_176);
or U1745 (N_1745,N_569,N_281);
nand U1746 (N_1746,N_245,N_289);
xor U1747 (N_1747,N_327,N_711);
nor U1748 (N_1748,N_821,N_902);
or U1749 (N_1749,N_220,N_981);
nor U1750 (N_1750,N_430,N_301);
or U1751 (N_1751,N_699,N_864);
and U1752 (N_1752,N_236,N_753);
nand U1753 (N_1753,N_51,N_160);
nand U1754 (N_1754,N_519,N_12);
nand U1755 (N_1755,N_74,N_448);
xor U1756 (N_1756,N_912,N_985);
or U1757 (N_1757,N_877,N_87);
nor U1758 (N_1758,N_532,N_940);
nand U1759 (N_1759,N_382,N_799);
or U1760 (N_1760,N_19,N_391);
nor U1761 (N_1761,N_627,N_32);
xor U1762 (N_1762,N_279,N_559);
nand U1763 (N_1763,N_365,N_66);
xnor U1764 (N_1764,N_788,N_551);
or U1765 (N_1765,N_698,N_619);
and U1766 (N_1766,N_75,N_218);
and U1767 (N_1767,N_973,N_879);
nand U1768 (N_1768,N_680,N_963);
xor U1769 (N_1769,N_747,N_612);
nand U1770 (N_1770,N_437,N_459);
or U1771 (N_1771,N_317,N_272);
and U1772 (N_1772,N_696,N_903);
xnor U1773 (N_1773,N_665,N_755);
xnor U1774 (N_1774,N_832,N_908);
or U1775 (N_1775,N_460,N_552);
nand U1776 (N_1776,N_797,N_167);
nor U1777 (N_1777,N_864,N_796);
and U1778 (N_1778,N_735,N_358);
nand U1779 (N_1779,N_37,N_312);
nand U1780 (N_1780,N_916,N_229);
nand U1781 (N_1781,N_830,N_298);
xnor U1782 (N_1782,N_702,N_435);
xor U1783 (N_1783,N_390,N_268);
nor U1784 (N_1784,N_629,N_854);
or U1785 (N_1785,N_275,N_734);
nand U1786 (N_1786,N_503,N_251);
nand U1787 (N_1787,N_873,N_54);
and U1788 (N_1788,N_284,N_726);
and U1789 (N_1789,N_649,N_841);
or U1790 (N_1790,N_212,N_826);
nand U1791 (N_1791,N_47,N_632);
or U1792 (N_1792,N_15,N_445);
and U1793 (N_1793,N_689,N_23);
nand U1794 (N_1794,N_818,N_351);
nor U1795 (N_1795,N_919,N_167);
nand U1796 (N_1796,N_52,N_532);
and U1797 (N_1797,N_358,N_539);
nor U1798 (N_1798,N_923,N_619);
xor U1799 (N_1799,N_48,N_803);
nor U1800 (N_1800,N_414,N_244);
nand U1801 (N_1801,N_703,N_788);
or U1802 (N_1802,N_552,N_190);
xor U1803 (N_1803,N_910,N_363);
nand U1804 (N_1804,N_211,N_266);
nand U1805 (N_1805,N_723,N_433);
or U1806 (N_1806,N_944,N_965);
nor U1807 (N_1807,N_767,N_804);
and U1808 (N_1808,N_676,N_605);
or U1809 (N_1809,N_327,N_649);
nor U1810 (N_1810,N_385,N_749);
and U1811 (N_1811,N_648,N_710);
and U1812 (N_1812,N_756,N_701);
nand U1813 (N_1813,N_372,N_333);
or U1814 (N_1814,N_195,N_714);
nor U1815 (N_1815,N_539,N_492);
xnor U1816 (N_1816,N_687,N_327);
and U1817 (N_1817,N_288,N_897);
nor U1818 (N_1818,N_614,N_525);
nor U1819 (N_1819,N_336,N_784);
or U1820 (N_1820,N_688,N_620);
or U1821 (N_1821,N_246,N_2);
nand U1822 (N_1822,N_621,N_105);
nor U1823 (N_1823,N_833,N_268);
xor U1824 (N_1824,N_99,N_388);
and U1825 (N_1825,N_348,N_906);
nor U1826 (N_1826,N_173,N_665);
and U1827 (N_1827,N_710,N_761);
or U1828 (N_1828,N_709,N_330);
xnor U1829 (N_1829,N_105,N_113);
nand U1830 (N_1830,N_411,N_978);
or U1831 (N_1831,N_596,N_851);
nand U1832 (N_1832,N_712,N_968);
or U1833 (N_1833,N_594,N_457);
xor U1834 (N_1834,N_745,N_193);
and U1835 (N_1835,N_794,N_180);
xor U1836 (N_1836,N_572,N_382);
or U1837 (N_1837,N_220,N_820);
nor U1838 (N_1838,N_100,N_582);
xnor U1839 (N_1839,N_114,N_274);
nor U1840 (N_1840,N_461,N_12);
or U1841 (N_1841,N_587,N_747);
or U1842 (N_1842,N_332,N_597);
or U1843 (N_1843,N_176,N_357);
xor U1844 (N_1844,N_195,N_364);
xnor U1845 (N_1845,N_519,N_272);
and U1846 (N_1846,N_204,N_137);
nor U1847 (N_1847,N_298,N_803);
and U1848 (N_1848,N_626,N_555);
or U1849 (N_1849,N_78,N_545);
nor U1850 (N_1850,N_205,N_5);
nor U1851 (N_1851,N_123,N_673);
nand U1852 (N_1852,N_670,N_179);
nand U1853 (N_1853,N_127,N_823);
nor U1854 (N_1854,N_26,N_675);
and U1855 (N_1855,N_398,N_794);
xnor U1856 (N_1856,N_985,N_814);
nand U1857 (N_1857,N_203,N_357);
or U1858 (N_1858,N_97,N_385);
xnor U1859 (N_1859,N_810,N_101);
nand U1860 (N_1860,N_401,N_345);
and U1861 (N_1861,N_390,N_972);
nand U1862 (N_1862,N_884,N_137);
xnor U1863 (N_1863,N_415,N_177);
xnor U1864 (N_1864,N_131,N_74);
nand U1865 (N_1865,N_46,N_457);
xnor U1866 (N_1866,N_937,N_203);
xor U1867 (N_1867,N_987,N_582);
xnor U1868 (N_1868,N_812,N_477);
xor U1869 (N_1869,N_222,N_654);
or U1870 (N_1870,N_714,N_326);
nand U1871 (N_1871,N_592,N_555);
xor U1872 (N_1872,N_22,N_42);
xnor U1873 (N_1873,N_586,N_622);
nand U1874 (N_1874,N_662,N_706);
and U1875 (N_1875,N_257,N_670);
or U1876 (N_1876,N_744,N_906);
and U1877 (N_1877,N_751,N_173);
nand U1878 (N_1878,N_642,N_758);
and U1879 (N_1879,N_419,N_76);
nor U1880 (N_1880,N_770,N_132);
or U1881 (N_1881,N_186,N_640);
or U1882 (N_1882,N_993,N_518);
xor U1883 (N_1883,N_272,N_19);
or U1884 (N_1884,N_291,N_838);
nor U1885 (N_1885,N_613,N_130);
or U1886 (N_1886,N_48,N_381);
and U1887 (N_1887,N_704,N_923);
nand U1888 (N_1888,N_538,N_400);
nor U1889 (N_1889,N_98,N_631);
nor U1890 (N_1890,N_584,N_272);
or U1891 (N_1891,N_671,N_378);
and U1892 (N_1892,N_156,N_417);
xnor U1893 (N_1893,N_507,N_304);
xnor U1894 (N_1894,N_336,N_936);
or U1895 (N_1895,N_630,N_362);
and U1896 (N_1896,N_39,N_147);
nor U1897 (N_1897,N_537,N_146);
nand U1898 (N_1898,N_289,N_74);
nand U1899 (N_1899,N_779,N_966);
and U1900 (N_1900,N_855,N_701);
xnor U1901 (N_1901,N_26,N_970);
and U1902 (N_1902,N_5,N_439);
nand U1903 (N_1903,N_637,N_360);
xor U1904 (N_1904,N_411,N_230);
xor U1905 (N_1905,N_848,N_481);
and U1906 (N_1906,N_268,N_989);
or U1907 (N_1907,N_795,N_871);
nor U1908 (N_1908,N_532,N_697);
nand U1909 (N_1909,N_560,N_846);
xnor U1910 (N_1910,N_451,N_938);
and U1911 (N_1911,N_84,N_191);
nor U1912 (N_1912,N_480,N_751);
xor U1913 (N_1913,N_329,N_726);
nand U1914 (N_1914,N_624,N_631);
and U1915 (N_1915,N_495,N_675);
and U1916 (N_1916,N_844,N_336);
nand U1917 (N_1917,N_535,N_482);
nor U1918 (N_1918,N_373,N_924);
xnor U1919 (N_1919,N_504,N_815);
or U1920 (N_1920,N_605,N_202);
and U1921 (N_1921,N_689,N_466);
nand U1922 (N_1922,N_739,N_753);
or U1923 (N_1923,N_152,N_61);
and U1924 (N_1924,N_926,N_669);
xor U1925 (N_1925,N_294,N_260);
nor U1926 (N_1926,N_654,N_344);
and U1927 (N_1927,N_910,N_678);
nor U1928 (N_1928,N_45,N_318);
or U1929 (N_1929,N_307,N_150);
or U1930 (N_1930,N_310,N_579);
nor U1931 (N_1931,N_562,N_761);
nand U1932 (N_1932,N_613,N_274);
and U1933 (N_1933,N_497,N_472);
xor U1934 (N_1934,N_467,N_813);
xnor U1935 (N_1935,N_907,N_522);
xnor U1936 (N_1936,N_581,N_673);
or U1937 (N_1937,N_617,N_843);
xnor U1938 (N_1938,N_9,N_931);
or U1939 (N_1939,N_919,N_830);
nor U1940 (N_1940,N_155,N_578);
or U1941 (N_1941,N_895,N_373);
nand U1942 (N_1942,N_259,N_76);
and U1943 (N_1943,N_919,N_853);
or U1944 (N_1944,N_93,N_306);
and U1945 (N_1945,N_124,N_744);
xor U1946 (N_1946,N_124,N_613);
xnor U1947 (N_1947,N_916,N_869);
nor U1948 (N_1948,N_64,N_641);
or U1949 (N_1949,N_674,N_274);
and U1950 (N_1950,N_127,N_685);
xor U1951 (N_1951,N_667,N_732);
xor U1952 (N_1952,N_578,N_998);
or U1953 (N_1953,N_466,N_650);
and U1954 (N_1954,N_147,N_192);
nand U1955 (N_1955,N_143,N_795);
or U1956 (N_1956,N_469,N_453);
nand U1957 (N_1957,N_564,N_49);
nor U1958 (N_1958,N_650,N_759);
nand U1959 (N_1959,N_499,N_124);
and U1960 (N_1960,N_932,N_891);
or U1961 (N_1961,N_223,N_712);
nor U1962 (N_1962,N_222,N_306);
nand U1963 (N_1963,N_973,N_647);
nand U1964 (N_1964,N_526,N_397);
nor U1965 (N_1965,N_335,N_92);
and U1966 (N_1966,N_874,N_477);
nor U1967 (N_1967,N_627,N_231);
xor U1968 (N_1968,N_562,N_732);
and U1969 (N_1969,N_3,N_870);
nor U1970 (N_1970,N_277,N_971);
nand U1971 (N_1971,N_16,N_439);
nor U1972 (N_1972,N_197,N_979);
xnor U1973 (N_1973,N_448,N_665);
xnor U1974 (N_1974,N_86,N_255);
nand U1975 (N_1975,N_642,N_444);
nand U1976 (N_1976,N_491,N_526);
nand U1977 (N_1977,N_16,N_600);
nand U1978 (N_1978,N_466,N_92);
and U1979 (N_1979,N_603,N_760);
and U1980 (N_1980,N_338,N_462);
xnor U1981 (N_1981,N_903,N_6);
xnor U1982 (N_1982,N_816,N_852);
xnor U1983 (N_1983,N_979,N_466);
and U1984 (N_1984,N_34,N_532);
nand U1985 (N_1985,N_73,N_891);
nand U1986 (N_1986,N_490,N_697);
nand U1987 (N_1987,N_549,N_857);
nor U1988 (N_1988,N_464,N_384);
and U1989 (N_1989,N_577,N_571);
nor U1990 (N_1990,N_917,N_361);
nor U1991 (N_1991,N_65,N_973);
and U1992 (N_1992,N_419,N_984);
or U1993 (N_1993,N_163,N_495);
xor U1994 (N_1994,N_925,N_546);
nor U1995 (N_1995,N_384,N_552);
nand U1996 (N_1996,N_2,N_837);
or U1997 (N_1997,N_891,N_472);
nor U1998 (N_1998,N_50,N_52);
or U1999 (N_1999,N_87,N_7);
and U2000 (N_2000,N_1212,N_1515);
nand U2001 (N_2001,N_1111,N_1385);
nor U2002 (N_2002,N_1912,N_1715);
nor U2003 (N_2003,N_1832,N_1195);
nor U2004 (N_2004,N_1357,N_1299);
nand U2005 (N_2005,N_1548,N_1849);
xnor U2006 (N_2006,N_1455,N_1817);
nand U2007 (N_2007,N_1102,N_1061);
nand U2008 (N_2008,N_1313,N_1487);
or U2009 (N_2009,N_1944,N_1230);
or U2010 (N_2010,N_1118,N_1044);
nand U2011 (N_2011,N_1448,N_1622);
xor U2012 (N_2012,N_1200,N_1030);
or U2013 (N_2013,N_1986,N_1175);
or U2014 (N_2014,N_1388,N_1908);
nand U2015 (N_2015,N_1786,N_1462);
or U2016 (N_2016,N_1775,N_1383);
nor U2017 (N_2017,N_1379,N_1966);
xor U2018 (N_2018,N_1626,N_1749);
xnor U2019 (N_2019,N_1063,N_1289);
and U2020 (N_2020,N_1425,N_1885);
nand U2021 (N_2021,N_1856,N_1360);
nor U2022 (N_2022,N_1130,N_1241);
nand U2023 (N_2023,N_1354,N_1311);
xnor U2024 (N_2024,N_1987,N_1623);
or U2025 (N_2025,N_1797,N_1416);
nand U2026 (N_2026,N_1043,N_1516);
and U2027 (N_2027,N_1016,N_1911);
nand U2028 (N_2028,N_1288,N_1024);
xor U2029 (N_2029,N_1133,N_1841);
and U2030 (N_2030,N_1657,N_1082);
xor U2031 (N_2031,N_1605,N_1371);
nand U2032 (N_2032,N_1834,N_1143);
xnor U2033 (N_2033,N_1062,N_1902);
nor U2034 (N_2034,N_1835,N_1337);
nand U2035 (N_2035,N_1333,N_1843);
nor U2036 (N_2036,N_1478,N_1501);
or U2037 (N_2037,N_1847,N_1512);
and U2038 (N_2038,N_1895,N_1837);
and U2039 (N_2039,N_1581,N_1977);
xnor U2040 (N_2040,N_1265,N_1142);
or U2041 (N_2041,N_1056,N_1374);
nand U2042 (N_2042,N_1361,N_1005);
nand U2043 (N_2043,N_1694,N_1316);
nor U2044 (N_2044,N_1092,N_1765);
xnor U2045 (N_2045,N_1366,N_1579);
nor U2046 (N_2046,N_1392,N_1629);
and U2047 (N_2047,N_1536,N_1719);
xnor U2048 (N_2048,N_1875,N_1563);
nor U2049 (N_2049,N_1009,N_1934);
nor U2050 (N_2050,N_1317,N_1370);
nor U2051 (N_2051,N_1463,N_1611);
or U2052 (N_2052,N_1356,N_1459);
nand U2053 (N_2053,N_1336,N_1635);
nand U2054 (N_2054,N_1960,N_1935);
or U2055 (N_2055,N_1739,N_1238);
xor U2056 (N_2056,N_1482,N_1619);
or U2057 (N_2057,N_1653,N_1669);
and U2058 (N_2058,N_1025,N_1612);
or U2059 (N_2059,N_1217,N_1907);
or U2060 (N_2060,N_1465,N_1625);
and U2061 (N_2061,N_1682,N_1822);
or U2062 (N_2062,N_1876,N_1393);
nand U2063 (N_2063,N_1840,N_1312);
and U2064 (N_2064,N_1365,N_1338);
and U2065 (N_2065,N_1162,N_1494);
and U2066 (N_2066,N_1576,N_1945);
nor U2067 (N_2067,N_1546,N_1464);
or U2068 (N_2068,N_1661,N_1387);
nor U2069 (N_2069,N_1743,N_1262);
or U2070 (N_2070,N_1326,N_1714);
and U2071 (N_2071,N_1893,N_1754);
nor U2072 (N_2072,N_1319,N_1003);
xnor U2073 (N_2073,N_1147,N_1483);
and U2074 (N_2074,N_1242,N_1268);
or U2075 (N_2075,N_1011,N_1164);
nor U2076 (N_2076,N_1770,N_1302);
nor U2077 (N_2077,N_1567,N_1584);
and U2078 (N_2078,N_1921,N_1747);
xnor U2079 (N_2079,N_1000,N_1137);
or U2080 (N_2080,N_1931,N_1359);
or U2081 (N_2081,N_1666,N_1367);
xor U2082 (N_2082,N_1826,N_1176);
xnor U2083 (N_2083,N_1368,N_1583);
xnor U2084 (N_2084,N_1178,N_1624);
or U2085 (N_2085,N_1110,N_1794);
nor U2086 (N_2086,N_1260,N_1777);
and U2087 (N_2087,N_1037,N_1404);
xnor U2088 (N_2088,N_1636,N_1245);
nor U2089 (N_2089,N_1124,N_1377);
or U2090 (N_2090,N_1809,N_1943);
xnor U2091 (N_2091,N_1671,N_1812);
nand U2092 (N_2092,N_1693,N_1014);
nor U2093 (N_2093,N_1284,N_1928);
or U2094 (N_2094,N_1120,N_1440);
nor U2095 (N_2095,N_1259,N_1709);
xor U2096 (N_2096,N_1380,N_1559);
or U2097 (N_2097,N_1099,N_1324);
nand U2098 (N_2098,N_1929,N_1270);
xnor U2099 (N_2099,N_1261,N_1329);
or U2100 (N_2100,N_1683,N_1010);
nor U2101 (N_2101,N_1039,N_1664);
and U2102 (N_2102,N_1557,N_1331);
and U2103 (N_2103,N_1112,N_1107);
or U2104 (N_2104,N_1229,N_1086);
and U2105 (N_2105,N_1156,N_1184);
and U2106 (N_2106,N_1988,N_1205);
nand U2107 (N_2107,N_1036,N_1627);
nand U2108 (N_2108,N_1158,N_1924);
nor U2109 (N_2109,N_1364,N_1057);
nand U2110 (N_2110,N_1767,N_1948);
nand U2111 (N_2111,N_1293,N_1613);
nor U2112 (N_2112,N_1077,N_1836);
nand U2113 (N_2113,N_1742,N_1633);
or U2114 (N_2114,N_1867,N_1597);
nor U2115 (N_2115,N_1710,N_1119);
and U2116 (N_2116,N_1760,N_1290);
and U2117 (N_2117,N_1862,N_1582);
nor U2118 (N_2118,N_1444,N_1511);
xor U2119 (N_2119,N_1236,N_1081);
and U2120 (N_2120,N_1746,N_1691);
nand U2121 (N_2121,N_1269,N_1053);
nor U2122 (N_2122,N_1466,N_1655);
or U2123 (N_2123,N_1609,N_1185);
nand U2124 (N_2124,N_1246,N_1071);
xnor U2125 (N_2125,N_1741,N_1266);
xnor U2126 (N_2126,N_1562,N_1221);
xor U2127 (N_2127,N_1272,N_1378);
and U2128 (N_2128,N_1280,N_1806);
or U2129 (N_2129,N_1373,N_1630);
nand U2130 (N_2130,N_1572,N_1493);
nand U2131 (N_2131,N_1752,N_1632);
or U2132 (N_2132,N_1473,N_1985);
nand U2133 (N_2133,N_1731,N_1561);
nand U2134 (N_2134,N_1306,N_1419);
or U2135 (N_2135,N_1698,N_1474);
nand U2136 (N_2136,N_1972,N_1406);
nor U2137 (N_2137,N_1070,N_1638);
and U2138 (N_2138,N_1545,N_1699);
or U2139 (N_2139,N_1964,N_1104);
xnor U2140 (N_2140,N_1244,N_1131);
and U2141 (N_2141,N_1254,N_1642);
or U2142 (N_2142,N_1798,N_1888);
nand U2143 (N_2143,N_1506,N_1873);
nor U2144 (N_2144,N_1762,N_1349);
nor U2145 (N_2145,N_1869,N_1128);
nor U2146 (N_2146,N_1983,N_1432);
and U2147 (N_2147,N_1883,N_1072);
xnor U2148 (N_2148,N_1858,N_1237);
nand U2149 (N_2149,N_1083,N_1891);
nor U2150 (N_2150,N_1517,N_1839);
and U2151 (N_2151,N_1369,N_1938);
nor U2152 (N_2152,N_1066,N_1748);
nor U2153 (N_2153,N_1295,N_1614);
and U2154 (N_2154,N_1541,N_1204);
and U2155 (N_2155,N_1880,N_1397);
nand U2156 (N_2156,N_1136,N_1502);
or U2157 (N_2157,N_1219,N_1159);
and U2158 (N_2158,N_1232,N_1171);
xor U2159 (N_2159,N_1967,N_1304);
or U2160 (N_2160,N_1643,N_1787);
or U2161 (N_2161,N_1507,N_1298);
xnor U2162 (N_2162,N_1441,N_1192);
or U2163 (N_2163,N_1115,N_1227);
xnor U2164 (N_2164,N_1553,N_1210);
or U2165 (N_2165,N_1804,N_1951);
or U2166 (N_2166,N_1410,N_1267);
nand U2167 (N_2167,N_1504,N_1530);
and U2168 (N_2168,N_1716,N_1727);
nor U2169 (N_2169,N_1045,N_1590);
xnor U2170 (N_2170,N_1052,N_1900);
or U2171 (N_2171,N_1776,N_1050);
nand U2172 (N_2172,N_1255,N_1520);
or U2173 (N_2173,N_1347,N_1215);
nor U2174 (N_2174,N_1861,N_1993);
or U2175 (N_2175,N_1384,N_1533);
xnor U2176 (N_2176,N_1292,N_1527);
or U2177 (N_2177,N_1844,N_1424);
xnor U2178 (N_2178,N_1962,N_1346);
nand U2179 (N_2179,N_1577,N_1882);
nor U2180 (N_2180,N_1558,N_1505);
nand U2181 (N_2181,N_1603,N_1477);
xnor U2182 (N_2182,N_1305,N_1447);
or U2183 (N_2183,N_1509,N_1355);
xor U2184 (N_2184,N_1146,N_1897);
xor U2185 (N_2185,N_1223,N_1251);
xnor U2186 (N_2186,N_1824,N_1398);
nand U2187 (N_2187,N_1064,N_1825);
or U2188 (N_2188,N_1264,N_1665);
nor U2189 (N_2189,N_1974,N_1157);
nor U2190 (N_2190,N_1386,N_1508);
and U2191 (N_2191,N_1994,N_1941);
nor U2192 (N_2192,N_1678,N_1495);
and U2193 (N_2193,N_1711,N_1981);
and U2194 (N_2194,N_1303,N_1422);
xor U2195 (N_2195,N_1173,N_1568);
or U2196 (N_2196,N_1889,N_1180);
and U2197 (N_2197,N_1187,N_1018);
and U2198 (N_2198,N_1183,N_1552);
or U2199 (N_2199,N_1046,N_1574);
nor U2200 (N_2200,N_1969,N_1389);
or U2201 (N_2201,N_1274,N_1652);
or U2202 (N_2202,N_1022,N_1729);
or U2203 (N_2203,N_1990,N_1055);
or U2204 (N_2204,N_1421,N_1872);
or U2205 (N_2205,N_1730,N_1013);
and U2206 (N_2206,N_1959,N_1109);
xnor U2207 (N_2207,N_1904,N_1496);
or U2208 (N_2208,N_1409,N_1769);
nor U2209 (N_2209,N_1500,N_1712);
xor U2210 (N_2210,N_1998,N_1756);
nor U2211 (N_2211,N_1203,N_1172);
nand U2212 (N_2212,N_1758,N_1968);
xnor U2213 (N_2213,N_1222,N_1982);
or U2214 (N_2214,N_1917,N_1961);
xor U2215 (N_2215,N_1439,N_1021);
xnor U2216 (N_2216,N_1975,N_1181);
or U2217 (N_2217,N_1795,N_1401);
nand U2218 (N_2218,N_1829,N_1139);
nor U2219 (N_2219,N_1980,N_1953);
and U2220 (N_2220,N_1126,N_1922);
nor U2221 (N_2221,N_1901,N_1855);
xor U2222 (N_2222,N_1191,N_1348);
or U2223 (N_2223,N_1695,N_1048);
or U2224 (N_2224,N_1209,N_1177);
nor U2225 (N_2225,N_1485,N_1282);
and U2226 (N_2226,N_1810,N_1239);
nor U2227 (N_2227,N_1087,N_1028);
nand U2228 (N_2228,N_1674,N_1224);
and U2229 (N_2229,N_1616,N_1454);
nor U2230 (N_2230,N_1101,N_1721);
and U2231 (N_2231,N_1750,N_1116);
or U2232 (N_2232,N_1725,N_1549);
nor U2233 (N_2233,N_1654,N_1755);
or U2234 (N_2234,N_1341,N_1343);
or U2235 (N_2235,N_1182,N_1351);
nor U2236 (N_2236,N_1382,N_1744);
nor U2237 (N_2237,N_1788,N_1012);
nand U2238 (N_2238,N_1098,N_1537);
and U2239 (N_2239,N_1151,N_1813);
nor U2240 (N_2240,N_1811,N_1491);
xnor U2241 (N_2241,N_1249,N_1390);
or U2242 (N_2242,N_1471,N_1723);
nor U2243 (N_2243,N_1641,N_1646);
xnor U2244 (N_2244,N_1503,N_1886);
nand U2245 (N_2245,N_1189,N_1538);
nand U2246 (N_2246,N_1396,N_1412);
nand U2247 (N_2247,N_1395,N_1970);
nor U2248 (N_2248,N_1645,N_1617);
or U2249 (N_2249,N_1342,N_1035);
nand U2250 (N_2250,N_1846,N_1704);
and U2251 (N_2251,N_1575,N_1535);
and U2252 (N_2252,N_1325,N_1958);
nand U2253 (N_2253,N_1615,N_1167);
nor U2254 (N_2254,N_1789,N_1675);
nand U2255 (N_2255,N_1978,N_1936);
nor U2256 (N_2256,N_1816,N_1550);
and U2257 (N_2257,N_1783,N_1257);
xor U2258 (N_2258,N_1468,N_1670);
and U2259 (N_2259,N_1915,N_1218);
or U2260 (N_2260,N_1526,N_1381);
xnor U2261 (N_2261,N_1093,N_1427);
xor U2262 (N_2262,N_1123,N_1054);
xnor U2263 (N_2263,N_1910,N_1141);
xor U2264 (N_2264,N_1854,N_1802);
and U2265 (N_2265,N_1857,N_1573);
or U2266 (N_2266,N_1321,N_1310);
or U2267 (N_2267,N_1275,N_1492);
nor U2268 (N_2268,N_1201,N_1866);
nand U2269 (N_2269,N_1089,N_1706);
nor U2270 (N_2270,N_1831,N_1434);
nand U2271 (N_2271,N_1732,N_1528);
nor U2272 (N_2272,N_1845,N_1091);
xor U2273 (N_2273,N_1997,N_1618);
nor U2274 (N_2274,N_1713,N_1129);
or U2275 (N_2275,N_1407,N_1426);
or U2276 (N_2276,N_1879,N_1593);
and U2277 (N_2277,N_1677,N_1995);
nor U2278 (N_2278,N_1318,N_1436);
or U2279 (N_2279,N_1955,N_1644);
nor U2280 (N_2280,N_1358,N_1808);
or U2281 (N_2281,N_1790,N_1127);
nand U2282 (N_2282,N_1438,N_1589);
and U2283 (N_2283,N_1942,N_1456);
or U2284 (N_2284,N_1247,N_1957);
nand U2285 (N_2285,N_1122,N_1352);
xnor U2286 (N_2286,N_1954,N_1405);
xor U2287 (N_2287,N_1174,N_1768);
nand U2288 (N_2288,N_1565,N_1668);
nor U2289 (N_2289,N_1345,N_1534);
or U2290 (N_2290,N_1340,N_1339);
nand U2291 (N_2291,N_1531,N_1874);
xnor U2292 (N_2292,N_1821,N_1034);
nand U2293 (N_2293,N_1315,N_1937);
nor U2294 (N_2294,N_1307,N_1453);
nor U2295 (N_2295,N_1163,N_1481);
nor U2296 (N_2296,N_1446,N_1460);
nor U2297 (N_2297,N_1042,N_1461);
and U2298 (N_2298,N_1566,N_1898);
nor U2299 (N_2299,N_1198,N_1870);
nor U2300 (N_2300,N_1335,N_1472);
and U2301 (N_2301,N_1068,N_1792);
nor U2302 (N_2302,N_1148,N_1234);
and U2303 (N_2303,N_1963,N_1927);
xnor U2304 (N_2304,N_1196,N_1300);
nand U2305 (N_2305,N_1864,N_1094);
nand U2306 (N_2306,N_1801,N_1051);
and U2307 (N_2307,N_1796,N_1038);
nand U2308 (N_2308,N_1740,N_1871);
nor U2309 (N_2309,N_1610,N_1428);
and U2310 (N_2310,N_1297,N_1031);
nand U2311 (N_2311,N_1235,N_1764);
xor U2312 (N_2312,N_1637,N_1169);
nor U2313 (N_2313,N_1601,N_1686);
and U2314 (N_2314,N_1296,N_1814);
nor U2315 (N_2315,N_1308,N_1585);
xnor U2316 (N_2316,N_1784,N_1728);
nand U2317 (N_2317,N_1006,N_1108);
nand U2318 (N_2318,N_1479,N_1703);
xnor U2319 (N_2319,N_1940,N_1949);
nand U2320 (N_2320,N_1134,N_1853);
xor U2321 (N_2321,N_1277,N_1090);
and U2322 (N_2322,N_1322,N_1569);
nor U2323 (N_2323,N_1604,N_1785);
xnor U2324 (N_2324,N_1400,N_1414);
nor U2325 (N_2325,N_1663,N_1916);
xor U2326 (N_2326,N_1586,N_1914);
nor U2327 (N_2327,N_1435,N_1486);
xor U2328 (N_2328,N_1827,N_1059);
and U2329 (N_2329,N_1078,N_1040);
and U2330 (N_2330,N_1079,N_1206);
or U2331 (N_2331,N_1166,N_1631);
xor U2332 (N_2332,N_1065,N_1830);
nor U2333 (N_2333,N_1376,N_1667);
xor U2334 (N_2334,N_1592,N_1570);
nor U2335 (N_2335,N_1580,N_1165);
xor U2336 (N_2336,N_1015,N_1228);
nand U2337 (N_2337,N_1539,N_1923);
and U2338 (N_2338,N_1620,N_1032);
xor U2339 (N_2339,N_1925,N_1542);
and U2340 (N_2340,N_1689,N_1271);
xnor U2341 (N_2341,N_1722,N_1488);
and U2342 (N_2342,N_1132,N_1168);
nor U2343 (N_2343,N_1708,N_1859);
and U2344 (N_2344,N_1773,N_1278);
or U2345 (N_2345,N_1252,N_1152);
nor U2346 (N_2346,N_1253,N_1469);
nand U2347 (N_2347,N_1639,N_1105);
or U2348 (N_2348,N_1648,N_1328);
nor U2349 (N_2349,N_1805,N_1423);
nor U2350 (N_2350,N_1145,N_1599);
nand U2351 (N_2351,N_1106,N_1170);
nor U2352 (N_2352,N_1403,N_1117);
nor U2353 (N_2353,N_1757,N_1930);
xnor U2354 (N_2354,N_1673,N_1323);
nor U2355 (N_2355,N_1860,N_1628);
nand U2356 (N_2356,N_1903,N_1430);
and U2357 (N_2357,N_1679,N_1362);
nor U2358 (N_2358,N_1096,N_1334);
and U2359 (N_2359,N_1294,N_1939);
or U2360 (N_2360,N_1519,N_1800);
or U2361 (N_2361,N_1417,N_1067);
and U2362 (N_2362,N_1220,N_1918);
nor U2363 (N_2363,N_1594,N_1420);
nand U2364 (N_2364,N_1027,N_1602);
xnor U2365 (N_2365,N_1571,N_1965);
xnor U2366 (N_2366,N_1726,N_1640);
or U2367 (N_2367,N_1480,N_1350);
and U2368 (N_2368,N_1375,N_1681);
or U2369 (N_2369,N_1399,N_1971);
nor U2370 (N_2370,N_1451,N_1705);
or U2371 (N_2371,N_1088,N_1452);
or U2372 (N_2372,N_1256,N_1720);
or U2373 (N_2373,N_1947,N_1233);
nand U2374 (N_2374,N_1084,N_1283);
and U2375 (N_2375,N_1258,N_1838);
or U2376 (N_2376,N_1865,N_1905);
or U2377 (N_2377,N_1819,N_1926);
xor U2378 (N_2378,N_1475,N_1717);
nand U2379 (N_2379,N_1153,N_1114);
xnor U2380 (N_2380,N_1179,N_1291);
xnor U2381 (N_2381,N_1076,N_1587);
and U2382 (N_2382,N_1413,N_1656);
nand U2383 (N_2383,N_1772,N_1216);
and U2384 (N_2384,N_1660,N_1411);
xor U2385 (N_2385,N_1848,N_1029);
xor U2386 (N_2386,N_1842,N_1286);
xnor U2387 (N_2387,N_1588,N_1208);
xor U2388 (N_2388,N_1763,N_1095);
and U2389 (N_2389,N_1608,N_1301);
xnor U2390 (N_2390,N_1909,N_1186);
or U2391 (N_2391,N_1202,N_1372);
xor U2392 (N_2392,N_1946,N_1919);
and U2393 (N_2393,N_1863,N_1884);
nor U2394 (N_2394,N_1135,N_1529);
xnor U2395 (N_2395,N_1598,N_1332);
nand U2396 (N_2396,N_1733,N_1458);
or U2397 (N_2397,N_1887,N_1649);
nor U2398 (N_2398,N_1188,N_1724);
and U2399 (N_2399,N_1578,N_1820);
nand U2400 (N_2400,N_1952,N_1815);
xnor U2401 (N_2401,N_1007,N_1737);
nor U2402 (N_2402,N_1778,N_1696);
and U2403 (N_2403,N_1833,N_1881);
xnor U2404 (N_2404,N_1596,N_1226);
or U2405 (N_2405,N_1155,N_1781);
nor U2406 (N_2406,N_1736,N_1144);
or U2407 (N_2407,N_1906,N_1659);
xnor U2408 (N_2408,N_1634,N_1564);
xor U2409 (N_2409,N_1248,N_1525);
nand U2410 (N_2410,N_1779,N_1522);
and U2411 (N_2411,N_1363,N_1085);
nand U2412 (N_2412,N_1672,N_1950);
or U2413 (N_2413,N_1606,N_1279);
and U2414 (N_2414,N_1433,N_1658);
nand U2415 (N_2415,N_1791,N_1243);
or U2416 (N_2416,N_1753,N_1418);
nand U2417 (N_2417,N_1979,N_1467);
xnor U2418 (N_2418,N_1149,N_1073);
nand U2419 (N_2419,N_1932,N_1676);
xnor U2420 (N_2420,N_1892,N_1484);
xnor U2421 (N_2421,N_1991,N_1999);
xnor U2422 (N_2422,N_1718,N_1852);
nand U2423 (N_2423,N_1514,N_1510);
nor U2424 (N_2424,N_1069,N_1281);
nor U2425 (N_2425,N_1556,N_1457);
nor U2426 (N_2426,N_1470,N_1100);
or U2427 (N_2427,N_1591,N_1896);
nor U2428 (N_2428,N_1276,N_1551);
nor U2429 (N_2429,N_1700,N_1499);
nor U2430 (N_2430,N_1759,N_1019);
and U2431 (N_2431,N_1524,N_1449);
or U2432 (N_2432,N_1913,N_1560);
or U2433 (N_2433,N_1330,N_1554);
and U2434 (N_2434,N_1685,N_1489);
and U2435 (N_2435,N_1097,N_1001);
xor U2436 (N_2436,N_1140,N_1956);
nor U2437 (N_2437,N_1074,N_1850);
nor U2438 (N_2438,N_1738,N_1992);
xor U2439 (N_2439,N_1877,N_1690);
nor U2440 (N_2440,N_1745,N_1799);
nor U2441 (N_2441,N_1075,N_1287);
or U2442 (N_2442,N_1314,N_1701);
and U2443 (N_2443,N_1213,N_1651);
and U2444 (N_2444,N_1734,N_1662);
or U2445 (N_2445,N_1199,N_1761);
or U2446 (N_2446,N_1523,N_1920);
xor U2447 (N_2447,N_1049,N_1450);
or U2448 (N_2448,N_1437,N_1020);
xor U2449 (N_2449,N_1543,N_1008);
or U2450 (N_2450,N_1408,N_1973);
nor U2451 (N_2451,N_1320,N_1415);
nor U2452 (N_2452,N_1544,N_1240);
and U2453 (N_2453,N_1002,N_1976);
xor U2454 (N_2454,N_1692,N_1868);
nor U2455 (N_2455,N_1309,N_1391);
and U2456 (N_2456,N_1607,N_1707);
or U2457 (N_2457,N_1735,N_1793);
nand U2458 (N_2458,N_1047,N_1194);
xor U2459 (N_2459,N_1121,N_1476);
nor U2460 (N_2460,N_1080,N_1443);
or U2461 (N_2461,N_1193,N_1807);
xnor U2462 (N_2462,N_1402,N_1431);
and U2463 (N_2463,N_1647,N_1680);
or U2464 (N_2464,N_1697,N_1150);
nor U2465 (N_2465,N_1497,N_1154);
nand U2466 (N_2466,N_1521,N_1540);
and U2467 (N_2467,N_1702,N_1033);
and U2468 (N_2468,N_1766,N_1621);
or U2469 (N_2469,N_1058,N_1041);
nand U2470 (N_2470,N_1595,N_1327);
xnor U2471 (N_2471,N_1394,N_1344);
or U2472 (N_2472,N_1125,N_1103);
xnor U2473 (N_2473,N_1989,N_1017);
xnor U2474 (N_2474,N_1160,N_1984);
nor U2475 (N_2475,N_1650,N_1490);
nor U2476 (N_2476,N_1060,N_1851);
nor U2477 (N_2477,N_1774,N_1211);
and U2478 (N_2478,N_1429,N_1225);
nand U2479 (N_2479,N_1688,N_1498);
xor U2480 (N_2480,N_1771,N_1353);
xnor U2481 (N_2481,N_1513,N_1823);
nand U2482 (N_2482,N_1113,N_1782);
or U2483 (N_2483,N_1442,N_1780);
and U2484 (N_2484,N_1818,N_1751);
and U2485 (N_2485,N_1207,N_1138);
or U2486 (N_2486,N_1273,N_1890);
and U2487 (N_2487,N_1026,N_1555);
or U2488 (N_2488,N_1004,N_1518);
nor U2489 (N_2489,N_1250,N_1263);
nor U2490 (N_2490,N_1445,N_1899);
or U2491 (N_2491,N_1803,N_1933);
and U2492 (N_2492,N_1285,N_1684);
xnor U2493 (N_2493,N_1878,N_1197);
nand U2494 (N_2494,N_1161,N_1231);
and U2495 (N_2495,N_1996,N_1547);
and U2496 (N_2496,N_1600,N_1214);
nand U2497 (N_2497,N_1894,N_1532);
or U2498 (N_2498,N_1828,N_1190);
nand U2499 (N_2499,N_1687,N_1023);
nor U2500 (N_2500,N_1101,N_1203);
and U2501 (N_2501,N_1142,N_1853);
and U2502 (N_2502,N_1808,N_1502);
xnor U2503 (N_2503,N_1815,N_1089);
nor U2504 (N_2504,N_1878,N_1439);
nand U2505 (N_2505,N_1220,N_1586);
and U2506 (N_2506,N_1324,N_1849);
xnor U2507 (N_2507,N_1937,N_1670);
nand U2508 (N_2508,N_1103,N_1006);
and U2509 (N_2509,N_1257,N_1355);
nand U2510 (N_2510,N_1801,N_1103);
nand U2511 (N_2511,N_1542,N_1403);
or U2512 (N_2512,N_1468,N_1624);
and U2513 (N_2513,N_1635,N_1782);
or U2514 (N_2514,N_1039,N_1354);
or U2515 (N_2515,N_1432,N_1483);
nand U2516 (N_2516,N_1062,N_1299);
and U2517 (N_2517,N_1215,N_1556);
nand U2518 (N_2518,N_1583,N_1800);
or U2519 (N_2519,N_1976,N_1235);
nor U2520 (N_2520,N_1693,N_1153);
nor U2521 (N_2521,N_1421,N_1230);
and U2522 (N_2522,N_1250,N_1350);
nor U2523 (N_2523,N_1602,N_1934);
or U2524 (N_2524,N_1196,N_1983);
or U2525 (N_2525,N_1939,N_1807);
nand U2526 (N_2526,N_1845,N_1012);
xor U2527 (N_2527,N_1253,N_1035);
xor U2528 (N_2528,N_1360,N_1805);
nand U2529 (N_2529,N_1106,N_1020);
nand U2530 (N_2530,N_1831,N_1044);
and U2531 (N_2531,N_1475,N_1438);
xnor U2532 (N_2532,N_1927,N_1796);
nand U2533 (N_2533,N_1299,N_1215);
and U2534 (N_2534,N_1957,N_1406);
or U2535 (N_2535,N_1402,N_1603);
nor U2536 (N_2536,N_1666,N_1299);
and U2537 (N_2537,N_1159,N_1832);
and U2538 (N_2538,N_1042,N_1498);
xor U2539 (N_2539,N_1947,N_1875);
or U2540 (N_2540,N_1521,N_1171);
or U2541 (N_2541,N_1310,N_1662);
xnor U2542 (N_2542,N_1085,N_1768);
or U2543 (N_2543,N_1575,N_1785);
and U2544 (N_2544,N_1880,N_1641);
or U2545 (N_2545,N_1539,N_1472);
or U2546 (N_2546,N_1880,N_1803);
xor U2547 (N_2547,N_1158,N_1205);
xor U2548 (N_2548,N_1528,N_1142);
nor U2549 (N_2549,N_1666,N_1560);
or U2550 (N_2550,N_1589,N_1514);
nor U2551 (N_2551,N_1642,N_1105);
or U2552 (N_2552,N_1118,N_1471);
nor U2553 (N_2553,N_1780,N_1660);
and U2554 (N_2554,N_1086,N_1515);
and U2555 (N_2555,N_1869,N_1487);
nor U2556 (N_2556,N_1336,N_1164);
nand U2557 (N_2557,N_1838,N_1344);
xor U2558 (N_2558,N_1284,N_1070);
xor U2559 (N_2559,N_1706,N_1079);
nor U2560 (N_2560,N_1876,N_1394);
or U2561 (N_2561,N_1667,N_1137);
nand U2562 (N_2562,N_1439,N_1484);
nor U2563 (N_2563,N_1711,N_1664);
nor U2564 (N_2564,N_1346,N_1983);
nand U2565 (N_2565,N_1714,N_1702);
nor U2566 (N_2566,N_1897,N_1815);
nand U2567 (N_2567,N_1268,N_1044);
or U2568 (N_2568,N_1544,N_1510);
xnor U2569 (N_2569,N_1437,N_1246);
nor U2570 (N_2570,N_1602,N_1423);
nor U2571 (N_2571,N_1540,N_1549);
nand U2572 (N_2572,N_1895,N_1090);
nand U2573 (N_2573,N_1545,N_1594);
nand U2574 (N_2574,N_1873,N_1482);
nand U2575 (N_2575,N_1328,N_1568);
or U2576 (N_2576,N_1614,N_1816);
nor U2577 (N_2577,N_1199,N_1541);
xor U2578 (N_2578,N_1118,N_1975);
xnor U2579 (N_2579,N_1841,N_1616);
or U2580 (N_2580,N_1205,N_1884);
xor U2581 (N_2581,N_1301,N_1439);
nor U2582 (N_2582,N_1312,N_1013);
or U2583 (N_2583,N_1252,N_1088);
nand U2584 (N_2584,N_1435,N_1605);
and U2585 (N_2585,N_1326,N_1929);
nand U2586 (N_2586,N_1272,N_1666);
nor U2587 (N_2587,N_1161,N_1651);
nand U2588 (N_2588,N_1449,N_1395);
or U2589 (N_2589,N_1932,N_1363);
or U2590 (N_2590,N_1246,N_1287);
xnor U2591 (N_2591,N_1813,N_1194);
and U2592 (N_2592,N_1007,N_1125);
xor U2593 (N_2593,N_1696,N_1690);
xor U2594 (N_2594,N_1754,N_1868);
or U2595 (N_2595,N_1880,N_1058);
or U2596 (N_2596,N_1815,N_1540);
nand U2597 (N_2597,N_1175,N_1501);
nand U2598 (N_2598,N_1699,N_1573);
and U2599 (N_2599,N_1124,N_1290);
nand U2600 (N_2600,N_1011,N_1328);
xor U2601 (N_2601,N_1842,N_1358);
or U2602 (N_2602,N_1584,N_1855);
xor U2603 (N_2603,N_1479,N_1464);
or U2604 (N_2604,N_1902,N_1275);
nand U2605 (N_2605,N_1672,N_1774);
nor U2606 (N_2606,N_1412,N_1649);
or U2607 (N_2607,N_1265,N_1505);
xor U2608 (N_2608,N_1411,N_1752);
and U2609 (N_2609,N_1375,N_1516);
xor U2610 (N_2610,N_1481,N_1567);
nand U2611 (N_2611,N_1532,N_1072);
nand U2612 (N_2612,N_1595,N_1655);
nor U2613 (N_2613,N_1743,N_1396);
or U2614 (N_2614,N_1506,N_1269);
nor U2615 (N_2615,N_1476,N_1936);
nand U2616 (N_2616,N_1323,N_1804);
or U2617 (N_2617,N_1063,N_1361);
xor U2618 (N_2618,N_1725,N_1356);
xnor U2619 (N_2619,N_1658,N_1721);
nor U2620 (N_2620,N_1527,N_1741);
nand U2621 (N_2621,N_1899,N_1774);
or U2622 (N_2622,N_1890,N_1806);
nor U2623 (N_2623,N_1917,N_1272);
nand U2624 (N_2624,N_1916,N_1366);
nor U2625 (N_2625,N_1325,N_1464);
nor U2626 (N_2626,N_1747,N_1625);
nor U2627 (N_2627,N_1223,N_1310);
and U2628 (N_2628,N_1328,N_1491);
nor U2629 (N_2629,N_1738,N_1580);
nor U2630 (N_2630,N_1160,N_1249);
and U2631 (N_2631,N_1451,N_1706);
nor U2632 (N_2632,N_1542,N_1965);
xnor U2633 (N_2633,N_1906,N_1825);
nand U2634 (N_2634,N_1591,N_1738);
and U2635 (N_2635,N_1325,N_1803);
nand U2636 (N_2636,N_1981,N_1031);
nor U2637 (N_2637,N_1740,N_1185);
nand U2638 (N_2638,N_1965,N_1910);
nand U2639 (N_2639,N_1155,N_1148);
or U2640 (N_2640,N_1117,N_1318);
and U2641 (N_2641,N_1373,N_1632);
and U2642 (N_2642,N_1029,N_1382);
nor U2643 (N_2643,N_1788,N_1464);
or U2644 (N_2644,N_1594,N_1527);
nand U2645 (N_2645,N_1391,N_1197);
and U2646 (N_2646,N_1686,N_1015);
nand U2647 (N_2647,N_1283,N_1438);
xnor U2648 (N_2648,N_1619,N_1883);
or U2649 (N_2649,N_1437,N_1176);
xnor U2650 (N_2650,N_1192,N_1272);
nor U2651 (N_2651,N_1028,N_1653);
and U2652 (N_2652,N_1277,N_1438);
xnor U2653 (N_2653,N_1222,N_1617);
and U2654 (N_2654,N_1410,N_1258);
nand U2655 (N_2655,N_1190,N_1676);
or U2656 (N_2656,N_1629,N_1302);
and U2657 (N_2657,N_1691,N_1032);
and U2658 (N_2658,N_1688,N_1272);
or U2659 (N_2659,N_1122,N_1102);
xor U2660 (N_2660,N_1862,N_1987);
and U2661 (N_2661,N_1727,N_1998);
nand U2662 (N_2662,N_1097,N_1391);
and U2663 (N_2663,N_1135,N_1684);
nor U2664 (N_2664,N_1027,N_1366);
xor U2665 (N_2665,N_1139,N_1252);
or U2666 (N_2666,N_1123,N_1775);
nor U2667 (N_2667,N_1832,N_1331);
and U2668 (N_2668,N_1140,N_1285);
xnor U2669 (N_2669,N_1591,N_1602);
or U2670 (N_2670,N_1490,N_1774);
nor U2671 (N_2671,N_1332,N_1981);
or U2672 (N_2672,N_1945,N_1494);
and U2673 (N_2673,N_1860,N_1012);
xnor U2674 (N_2674,N_1077,N_1363);
nor U2675 (N_2675,N_1629,N_1287);
nor U2676 (N_2676,N_1518,N_1876);
or U2677 (N_2677,N_1425,N_1123);
nor U2678 (N_2678,N_1873,N_1238);
or U2679 (N_2679,N_1852,N_1021);
nor U2680 (N_2680,N_1328,N_1293);
nand U2681 (N_2681,N_1985,N_1983);
xnor U2682 (N_2682,N_1787,N_1732);
xnor U2683 (N_2683,N_1040,N_1971);
and U2684 (N_2684,N_1971,N_1112);
nand U2685 (N_2685,N_1903,N_1661);
nor U2686 (N_2686,N_1371,N_1378);
nor U2687 (N_2687,N_1067,N_1469);
or U2688 (N_2688,N_1314,N_1369);
nor U2689 (N_2689,N_1266,N_1853);
or U2690 (N_2690,N_1853,N_1346);
xnor U2691 (N_2691,N_1993,N_1463);
and U2692 (N_2692,N_1569,N_1782);
or U2693 (N_2693,N_1528,N_1918);
nand U2694 (N_2694,N_1572,N_1891);
nand U2695 (N_2695,N_1205,N_1892);
and U2696 (N_2696,N_1137,N_1538);
and U2697 (N_2697,N_1550,N_1498);
xor U2698 (N_2698,N_1851,N_1461);
nand U2699 (N_2699,N_1467,N_1211);
or U2700 (N_2700,N_1349,N_1508);
nor U2701 (N_2701,N_1766,N_1500);
and U2702 (N_2702,N_1351,N_1213);
xor U2703 (N_2703,N_1107,N_1971);
or U2704 (N_2704,N_1198,N_1605);
nor U2705 (N_2705,N_1108,N_1712);
and U2706 (N_2706,N_1086,N_1893);
nand U2707 (N_2707,N_1941,N_1286);
or U2708 (N_2708,N_1322,N_1120);
nand U2709 (N_2709,N_1694,N_1950);
xor U2710 (N_2710,N_1952,N_1965);
nand U2711 (N_2711,N_1563,N_1582);
or U2712 (N_2712,N_1032,N_1747);
nand U2713 (N_2713,N_1944,N_1665);
or U2714 (N_2714,N_1666,N_1316);
xor U2715 (N_2715,N_1551,N_1753);
or U2716 (N_2716,N_1061,N_1214);
nand U2717 (N_2717,N_1163,N_1656);
and U2718 (N_2718,N_1287,N_1680);
or U2719 (N_2719,N_1600,N_1343);
nor U2720 (N_2720,N_1494,N_1558);
nand U2721 (N_2721,N_1330,N_1217);
nor U2722 (N_2722,N_1123,N_1319);
and U2723 (N_2723,N_1120,N_1050);
nor U2724 (N_2724,N_1768,N_1468);
xnor U2725 (N_2725,N_1155,N_1259);
nand U2726 (N_2726,N_1541,N_1678);
and U2727 (N_2727,N_1470,N_1587);
nor U2728 (N_2728,N_1270,N_1585);
or U2729 (N_2729,N_1875,N_1098);
xnor U2730 (N_2730,N_1708,N_1611);
and U2731 (N_2731,N_1221,N_1601);
or U2732 (N_2732,N_1634,N_1685);
nor U2733 (N_2733,N_1522,N_1540);
nand U2734 (N_2734,N_1026,N_1432);
or U2735 (N_2735,N_1153,N_1326);
xor U2736 (N_2736,N_1093,N_1484);
nor U2737 (N_2737,N_1055,N_1002);
and U2738 (N_2738,N_1374,N_1242);
and U2739 (N_2739,N_1252,N_1126);
xnor U2740 (N_2740,N_1584,N_1205);
nand U2741 (N_2741,N_1042,N_1533);
nor U2742 (N_2742,N_1409,N_1735);
or U2743 (N_2743,N_1249,N_1948);
or U2744 (N_2744,N_1594,N_1941);
and U2745 (N_2745,N_1246,N_1312);
or U2746 (N_2746,N_1964,N_1421);
nor U2747 (N_2747,N_1430,N_1377);
or U2748 (N_2748,N_1757,N_1372);
nand U2749 (N_2749,N_1422,N_1487);
xor U2750 (N_2750,N_1836,N_1464);
and U2751 (N_2751,N_1144,N_1145);
or U2752 (N_2752,N_1615,N_1362);
nand U2753 (N_2753,N_1267,N_1219);
nor U2754 (N_2754,N_1189,N_1417);
nand U2755 (N_2755,N_1310,N_1758);
and U2756 (N_2756,N_1416,N_1941);
or U2757 (N_2757,N_1848,N_1157);
nand U2758 (N_2758,N_1520,N_1198);
or U2759 (N_2759,N_1878,N_1697);
nor U2760 (N_2760,N_1837,N_1698);
xor U2761 (N_2761,N_1343,N_1020);
or U2762 (N_2762,N_1852,N_1831);
nand U2763 (N_2763,N_1640,N_1690);
and U2764 (N_2764,N_1024,N_1154);
nand U2765 (N_2765,N_1390,N_1853);
xor U2766 (N_2766,N_1409,N_1151);
or U2767 (N_2767,N_1066,N_1140);
xor U2768 (N_2768,N_1200,N_1253);
or U2769 (N_2769,N_1786,N_1330);
nor U2770 (N_2770,N_1867,N_1420);
nand U2771 (N_2771,N_1792,N_1795);
and U2772 (N_2772,N_1732,N_1232);
nor U2773 (N_2773,N_1548,N_1117);
or U2774 (N_2774,N_1343,N_1376);
or U2775 (N_2775,N_1283,N_1630);
and U2776 (N_2776,N_1454,N_1675);
nor U2777 (N_2777,N_1641,N_1835);
and U2778 (N_2778,N_1853,N_1802);
and U2779 (N_2779,N_1856,N_1250);
xor U2780 (N_2780,N_1557,N_1164);
nand U2781 (N_2781,N_1399,N_1974);
nand U2782 (N_2782,N_1303,N_1553);
nor U2783 (N_2783,N_1182,N_1433);
nor U2784 (N_2784,N_1217,N_1070);
xor U2785 (N_2785,N_1114,N_1385);
xnor U2786 (N_2786,N_1965,N_1106);
xnor U2787 (N_2787,N_1825,N_1969);
or U2788 (N_2788,N_1461,N_1603);
or U2789 (N_2789,N_1469,N_1943);
xor U2790 (N_2790,N_1463,N_1786);
or U2791 (N_2791,N_1630,N_1439);
nand U2792 (N_2792,N_1792,N_1727);
and U2793 (N_2793,N_1811,N_1493);
and U2794 (N_2794,N_1799,N_1842);
or U2795 (N_2795,N_1957,N_1323);
and U2796 (N_2796,N_1352,N_1136);
or U2797 (N_2797,N_1439,N_1057);
and U2798 (N_2798,N_1176,N_1006);
nand U2799 (N_2799,N_1191,N_1545);
and U2800 (N_2800,N_1175,N_1117);
and U2801 (N_2801,N_1230,N_1663);
nand U2802 (N_2802,N_1893,N_1865);
nor U2803 (N_2803,N_1501,N_1151);
xnor U2804 (N_2804,N_1993,N_1561);
xor U2805 (N_2805,N_1572,N_1090);
or U2806 (N_2806,N_1015,N_1540);
or U2807 (N_2807,N_1976,N_1045);
nand U2808 (N_2808,N_1142,N_1882);
nor U2809 (N_2809,N_1334,N_1341);
xor U2810 (N_2810,N_1906,N_1385);
xnor U2811 (N_2811,N_1901,N_1219);
and U2812 (N_2812,N_1417,N_1629);
nor U2813 (N_2813,N_1886,N_1740);
or U2814 (N_2814,N_1516,N_1621);
xnor U2815 (N_2815,N_1152,N_1038);
or U2816 (N_2816,N_1744,N_1626);
nand U2817 (N_2817,N_1521,N_1269);
or U2818 (N_2818,N_1557,N_1407);
nand U2819 (N_2819,N_1131,N_1598);
nand U2820 (N_2820,N_1475,N_1879);
nor U2821 (N_2821,N_1152,N_1418);
or U2822 (N_2822,N_1956,N_1614);
nand U2823 (N_2823,N_1940,N_1628);
nand U2824 (N_2824,N_1994,N_1865);
or U2825 (N_2825,N_1373,N_1763);
nor U2826 (N_2826,N_1110,N_1504);
nor U2827 (N_2827,N_1669,N_1114);
nand U2828 (N_2828,N_1907,N_1955);
xnor U2829 (N_2829,N_1807,N_1773);
xnor U2830 (N_2830,N_1352,N_1008);
or U2831 (N_2831,N_1435,N_1612);
xor U2832 (N_2832,N_1803,N_1459);
nand U2833 (N_2833,N_1933,N_1343);
and U2834 (N_2834,N_1210,N_1769);
xnor U2835 (N_2835,N_1550,N_1820);
xor U2836 (N_2836,N_1768,N_1993);
xor U2837 (N_2837,N_1156,N_1768);
nor U2838 (N_2838,N_1453,N_1711);
nor U2839 (N_2839,N_1674,N_1155);
xor U2840 (N_2840,N_1245,N_1492);
nand U2841 (N_2841,N_1173,N_1252);
nand U2842 (N_2842,N_1863,N_1324);
nor U2843 (N_2843,N_1032,N_1385);
xor U2844 (N_2844,N_1195,N_1190);
and U2845 (N_2845,N_1292,N_1724);
or U2846 (N_2846,N_1887,N_1498);
nand U2847 (N_2847,N_1005,N_1514);
and U2848 (N_2848,N_1909,N_1727);
and U2849 (N_2849,N_1918,N_1560);
xnor U2850 (N_2850,N_1896,N_1098);
nand U2851 (N_2851,N_1600,N_1509);
and U2852 (N_2852,N_1775,N_1522);
nor U2853 (N_2853,N_1137,N_1439);
nor U2854 (N_2854,N_1677,N_1754);
and U2855 (N_2855,N_1269,N_1548);
xor U2856 (N_2856,N_1841,N_1394);
or U2857 (N_2857,N_1099,N_1187);
or U2858 (N_2858,N_1586,N_1480);
xor U2859 (N_2859,N_1353,N_1798);
nand U2860 (N_2860,N_1478,N_1174);
xnor U2861 (N_2861,N_1355,N_1459);
or U2862 (N_2862,N_1619,N_1529);
or U2863 (N_2863,N_1148,N_1839);
nand U2864 (N_2864,N_1539,N_1054);
nand U2865 (N_2865,N_1548,N_1508);
or U2866 (N_2866,N_1337,N_1118);
and U2867 (N_2867,N_1658,N_1392);
xor U2868 (N_2868,N_1281,N_1518);
or U2869 (N_2869,N_1411,N_1724);
or U2870 (N_2870,N_1688,N_1636);
or U2871 (N_2871,N_1638,N_1734);
and U2872 (N_2872,N_1899,N_1880);
nand U2873 (N_2873,N_1749,N_1895);
xor U2874 (N_2874,N_1958,N_1693);
and U2875 (N_2875,N_1835,N_1270);
nor U2876 (N_2876,N_1866,N_1220);
nand U2877 (N_2877,N_1506,N_1475);
nor U2878 (N_2878,N_1434,N_1247);
xnor U2879 (N_2879,N_1638,N_1303);
and U2880 (N_2880,N_1519,N_1697);
nand U2881 (N_2881,N_1314,N_1380);
nor U2882 (N_2882,N_1664,N_1268);
nand U2883 (N_2883,N_1774,N_1259);
nor U2884 (N_2884,N_1467,N_1961);
nand U2885 (N_2885,N_1809,N_1853);
and U2886 (N_2886,N_1890,N_1239);
and U2887 (N_2887,N_1233,N_1405);
nand U2888 (N_2888,N_1864,N_1030);
or U2889 (N_2889,N_1810,N_1435);
xnor U2890 (N_2890,N_1369,N_1618);
xor U2891 (N_2891,N_1948,N_1686);
or U2892 (N_2892,N_1661,N_1459);
and U2893 (N_2893,N_1386,N_1136);
nor U2894 (N_2894,N_1197,N_1799);
nor U2895 (N_2895,N_1358,N_1610);
nand U2896 (N_2896,N_1897,N_1253);
nand U2897 (N_2897,N_1121,N_1597);
xnor U2898 (N_2898,N_1155,N_1130);
nand U2899 (N_2899,N_1264,N_1533);
nor U2900 (N_2900,N_1135,N_1535);
nor U2901 (N_2901,N_1111,N_1312);
nand U2902 (N_2902,N_1469,N_1701);
xor U2903 (N_2903,N_1979,N_1448);
nor U2904 (N_2904,N_1089,N_1352);
nor U2905 (N_2905,N_1260,N_1566);
and U2906 (N_2906,N_1685,N_1514);
and U2907 (N_2907,N_1072,N_1411);
nand U2908 (N_2908,N_1155,N_1029);
nand U2909 (N_2909,N_1644,N_1384);
nor U2910 (N_2910,N_1975,N_1131);
nand U2911 (N_2911,N_1222,N_1356);
or U2912 (N_2912,N_1899,N_1893);
and U2913 (N_2913,N_1594,N_1062);
or U2914 (N_2914,N_1313,N_1859);
nand U2915 (N_2915,N_1989,N_1598);
xnor U2916 (N_2916,N_1919,N_1334);
or U2917 (N_2917,N_1432,N_1751);
or U2918 (N_2918,N_1540,N_1747);
nand U2919 (N_2919,N_1630,N_1995);
and U2920 (N_2920,N_1593,N_1769);
nor U2921 (N_2921,N_1177,N_1208);
or U2922 (N_2922,N_1865,N_1391);
nand U2923 (N_2923,N_1114,N_1847);
nor U2924 (N_2924,N_1275,N_1770);
xor U2925 (N_2925,N_1027,N_1763);
and U2926 (N_2926,N_1271,N_1132);
xor U2927 (N_2927,N_1335,N_1992);
xor U2928 (N_2928,N_1720,N_1035);
nor U2929 (N_2929,N_1185,N_1591);
xnor U2930 (N_2930,N_1573,N_1172);
nor U2931 (N_2931,N_1400,N_1943);
nor U2932 (N_2932,N_1048,N_1785);
nor U2933 (N_2933,N_1309,N_1153);
nor U2934 (N_2934,N_1350,N_1491);
or U2935 (N_2935,N_1895,N_1424);
nor U2936 (N_2936,N_1875,N_1630);
nand U2937 (N_2937,N_1815,N_1785);
and U2938 (N_2938,N_1344,N_1857);
or U2939 (N_2939,N_1607,N_1510);
and U2940 (N_2940,N_1658,N_1085);
nand U2941 (N_2941,N_1320,N_1088);
and U2942 (N_2942,N_1848,N_1592);
xor U2943 (N_2943,N_1256,N_1174);
or U2944 (N_2944,N_1969,N_1943);
nor U2945 (N_2945,N_1872,N_1090);
nor U2946 (N_2946,N_1987,N_1768);
and U2947 (N_2947,N_1207,N_1089);
nand U2948 (N_2948,N_1594,N_1322);
xnor U2949 (N_2949,N_1209,N_1253);
xor U2950 (N_2950,N_1130,N_1931);
xnor U2951 (N_2951,N_1526,N_1986);
xor U2952 (N_2952,N_1554,N_1907);
and U2953 (N_2953,N_1919,N_1732);
nor U2954 (N_2954,N_1757,N_1564);
or U2955 (N_2955,N_1916,N_1876);
or U2956 (N_2956,N_1931,N_1965);
or U2957 (N_2957,N_1668,N_1371);
nor U2958 (N_2958,N_1856,N_1511);
and U2959 (N_2959,N_1879,N_1710);
and U2960 (N_2960,N_1505,N_1073);
nor U2961 (N_2961,N_1198,N_1111);
xor U2962 (N_2962,N_1810,N_1120);
xor U2963 (N_2963,N_1665,N_1838);
and U2964 (N_2964,N_1429,N_1884);
or U2965 (N_2965,N_1261,N_1079);
nand U2966 (N_2966,N_1342,N_1956);
nand U2967 (N_2967,N_1823,N_1557);
xor U2968 (N_2968,N_1889,N_1887);
nor U2969 (N_2969,N_1975,N_1907);
xnor U2970 (N_2970,N_1100,N_1012);
and U2971 (N_2971,N_1439,N_1799);
xor U2972 (N_2972,N_1816,N_1227);
and U2973 (N_2973,N_1194,N_1230);
nand U2974 (N_2974,N_1749,N_1087);
or U2975 (N_2975,N_1985,N_1555);
nor U2976 (N_2976,N_1359,N_1318);
xnor U2977 (N_2977,N_1278,N_1914);
or U2978 (N_2978,N_1872,N_1516);
or U2979 (N_2979,N_1966,N_1295);
nand U2980 (N_2980,N_1660,N_1517);
xnor U2981 (N_2981,N_1917,N_1950);
and U2982 (N_2982,N_1425,N_1857);
nor U2983 (N_2983,N_1830,N_1627);
nor U2984 (N_2984,N_1925,N_1836);
xnor U2985 (N_2985,N_1985,N_1449);
xor U2986 (N_2986,N_1998,N_1421);
nor U2987 (N_2987,N_1713,N_1687);
xnor U2988 (N_2988,N_1122,N_1745);
and U2989 (N_2989,N_1758,N_1790);
nor U2990 (N_2990,N_1978,N_1143);
xor U2991 (N_2991,N_1684,N_1680);
and U2992 (N_2992,N_1541,N_1596);
nand U2993 (N_2993,N_1204,N_1993);
or U2994 (N_2994,N_1388,N_1924);
nor U2995 (N_2995,N_1800,N_1441);
or U2996 (N_2996,N_1935,N_1733);
nand U2997 (N_2997,N_1970,N_1160);
nor U2998 (N_2998,N_1962,N_1811);
nor U2999 (N_2999,N_1828,N_1722);
xnor U3000 (N_3000,N_2212,N_2600);
or U3001 (N_3001,N_2035,N_2065);
and U3002 (N_3002,N_2272,N_2576);
xnor U3003 (N_3003,N_2870,N_2311);
nor U3004 (N_3004,N_2275,N_2526);
xor U3005 (N_3005,N_2442,N_2683);
nor U3006 (N_3006,N_2350,N_2131);
and U3007 (N_3007,N_2684,N_2935);
and U3008 (N_3008,N_2573,N_2174);
or U3009 (N_3009,N_2293,N_2114);
nor U3010 (N_3010,N_2173,N_2578);
xnor U3011 (N_3011,N_2037,N_2844);
nand U3012 (N_3012,N_2495,N_2728);
xnor U3013 (N_3013,N_2997,N_2286);
nor U3014 (N_3014,N_2787,N_2671);
nor U3015 (N_3015,N_2553,N_2108);
and U3016 (N_3016,N_2920,N_2497);
xor U3017 (N_3017,N_2024,N_2023);
xor U3018 (N_3018,N_2511,N_2030);
or U3019 (N_3019,N_2313,N_2807);
xnor U3020 (N_3020,N_2784,N_2762);
and U3021 (N_3021,N_2727,N_2849);
or U3022 (N_3022,N_2999,N_2195);
nor U3023 (N_3023,N_2458,N_2247);
xor U3024 (N_3024,N_2720,N_2305);
and U3025 (N_3025,N_2322,N_2220);
xor U3026 (N_3026,N_2358,N_2089);
xor U3027 (N_3027,N_2123,N_2067);
nand U3028 (N_3028,N_2763,N_2813);
nand U3029 (N_3029,N_2388,N_2042);
nor U3030 (N_3030,N_2421,N_2517);
nor U3031 (N_3031,N_2982,N_2349);
xor U3032 (N_3032,N_2981,N_2282);
or U3033 (N_3033,N_2060,N_2596);
and U3034 (N_3034,N_2280,N_2484);
and U3035 (N_3035,N_2008,N_2529);
or U3036 (N_3036,N_2003,N_2096);
xor U3037 (N_3037,N_2348,N_2736);
and U3038 (N_3038,N_2558,N_2869);
nor U3039 (N_3039,N_2045,N_2423);
or U3040 (N_3040,N_2678,N_2256);
xor U3041 (N_3041,N_2629,N_2375);
nor U3042 (N_3042,N_2960,N_2907);
or U3043 (N_3043,N_2798,N_2461);
xnor U3044 (N_3044,N_2858,N_2191);
nand U3045 (N_3045,N_2382,N_2536);
or U3046 (N_3046,N_2758,N_2038);
xor U3047 (N_3047,N_2347,N_2779);
nor U3048 (N_3048,N_2092,N_2319);
nor U3049 (N_3049,N_2144,N_2821);
and U3050 (N_3050,N_2519,N_2948);
nand U3051 (N_3051,N_2409,N_2770);
and U3052 (N_3052,N_2002,N_2925);
nor U3053 (N_3053,N_2261,N_2047);
nor U3054 (N_3054,N_2694,N_2102);
and U3055 (N_3055,N_2545,N_2569);
xnor U3056 (N_3056,N_2662,N_2039);
and U3057 (N_3057,N_2974,N_2147);
and U3058 (N_3058,N_2182,N_2524);
and U3059 (N_3059,N_2508,N_2051);
xor U3060 (N_3060,N_2118,N_2747);
nor U3061 (N_3061,N_2165,N_2062);
nor U3062 (N_3062,N_2730,N_2766);
or U3063 (N_3063,N_2289,N_2143);
nand U3064 (N_3064,N_2676,N_2721);
or U3065 (N_3065,N_2091,N_2107);
and U3066 (N_3066,N_2128,N_2203);
xor U3067 (N_3067,N_2263,N_2797);
nand U3068 (N_3068,N_2538,N_2396);
or U3069 (N_3069,N_2176,N_2132);
xnor U3070 (N_3070,N_2453,N_2777);
and U3071 (N_3071,N_2259,N_2656);
and U3072 (N_3072,N_2200,N_2244);
or U3073 (N_3073,N_2947,N_2837);
nor U3074 (N_3074,N_2215,N_2796);
nor U3075 (N_3075,N_2876,N_2959);
nand U3076 (N_3076,N_2056,N_2253);
xor U3077 (N_3077,N_2429,N_2480);
nand U3078 (N_3078,N_2510,N_2991);
and U3079 (N_3079,N_2563,N_2468);
nand U3080 (N_3080,N_2390,N_2125);
or U3081 (N_3081,N_2250,N_2514);
and U3082 (N_3082,N_2740,N_2902);
xor U3083 (N_3083,N_2428,N_2521);
nand U3084 (N_3084,N_2665,N_2823);
nand U3085 (N_3085,N_2994,N_2326);
nand U3086 (N_3086,N_2462,N_2842);
xnor U3087 (N_3087,N_2507,N_2626);
nor U3088 (N_3088,N_2954,N_2376);
nand U3089 (N_3089,N_2893,N_2279);
xor U3090 (N_3090,N_2828,N_2969);
and U3091 (N_3091,N_2093,N_2454);
and U3092 (N_3092,N_2044,N_2196);
xnor U3093 (N_3093,N_2978,N_2599);
nor U3094 (N_3094,N_2713,N_2416);
nand U3095 (N_3095,N_2638,N_2465);
nand U3096 (N_3096,N_2082,N_2815);
and U3097 (N_3097,N_2682,N_2373);
and U3098 (N_3098,N_2417,N_2567);
nand U3099 (N_3099,N_2254,N_2792);
and U3100 (N_3100,N_2587,N_2729);
and U3101 (N_3101,N_2820,N_2891);
nand U3102 (N_3102,N_2722,N_2185);
nand U3103 (N_3103,N_2169,N_2381);
and U3104 (N_3104,N_2258,N_2550);
or U3105 (N_3105,N_2238,N_2219);
nand U3106 (N_3106,N_2257,N_2485);
nor U3107 (N_3107,N_2213,N_2101);
nand U3108 (N_3108,N_2865,N_2325);
nand U3109 (N_3109,N_2631,N_2591);
nor U3110 (N_3110,N_2360,N_2854);
and U3111 (N_3111,N_2308,N_2698);
or U3112 (N_3112,N_2337,N_2150);
xnor U3113 (N_3113,N_2316,N_2644);
xnor U3114 (N_3114,N_2885,N_2509);
and U3115 (N_3115,N_2868,N_2264);
nor U3116 (N_3116,N_2365,N_2085);
or U3117 (N_3117,N_2448,N_2913);
nor U3118 (N_3118,N_2774,N_2690);
nand U3119 (N_3119,N_2470,N_2702);
or U3120 (N_3120,N_2007,N_2934);
xnor U3121 (N_3121,N_2731,N_2776);
xnor U3122 (N_3122,N_2921,N_2696);
or U3123 (N_3123,N_2896,N_2703);
or U3124 (N_3124,N_2335,N_2601);
and U3125 (N_3125,N_2928,N_2034);
xor U3126 (N_3126,N_2245,N_2803);
xnor U3127 (N_3127,N_2119,N_2831);
xor U3128 (N_3128,N_2383,N_2148);
and U3129 (N_3129,N_2834,N_2384);
nand U3130 (N_3130,N_2100,N_2754);
or U3131 (N_3131,N_2363,N_2490);
or U3132 (N_3132,N_2801,N_2782);
nand U3133 (N_3133,N_2989,N_2836);
xnor U3134 (N_3134,N_2752,N_2369);
xor U3135 (N_3135,N_2218,N_2975);
and U3136 (N_3136,N_2287,N_2548);
or U3137 (N_3137,N_2446,N_2415);
and U3138 (N_3138,N_2967,N_2370);
nand U3139 (N_3139,N_2001,N_2641);
nor U3140 (N_3140,N_2945,N_2068);
xor U3141 (N_3141,N_2004,N_2496);
nand U3142 (N_3142,N_2239,N_2126);
or U3143 (N_3143,N_2328,N_2340);
nor U3144 (N_3144,N_2177,N_2192);
xnor U3145 (N_3145,N_2883,N_2564);
or U3146 (N_3146,N_2299,N_2315);
and U3147 (N_3147,N_2594,N_2406);
nand U3148 (N_3148,N_2016,N_2931);
or U3149 (N_3149,N_2367,N_2265);
or U3150 (N_3150,N_2804,N_2281);
and U3151 (N_3151,N_2221,N_2847);
or U3152 (N_3152,N_2582,N_2839);
nand U3153 (N_3153,N_2886,N_2602);
or U3154 (N_3154,N_2664,N_2958);
nand U3155 (N_3155,N_2990,N_2492);
and U3156 (N_3156,N_2320,N_2133);
nor U3157 (N_3157,N_2022,N_2592);
nand U3158 (N_3158,N_2046,N_2426);
or U3159 (N_3159,N_2788,N_2314);
nor U3160 (N_3160,N_2693,N_2867);
nor U3161 (N_3161,N_2850,N_2194);
nor U3162 (N_3162,N_2912,N_2642);
xnor U3163 (N_3163,N_2033,N_2106);
nand U3164 (N_3164,N_2086,N_2742);
nor U3165 (N_3165,N_2162,N_2477);
xnor U3166 (N_3166,N_2819,N_2400);
nor U3167 (N_3167,N_2310,N_2809);
xnor U3168 (N_3168,N_2649,N_2043);
nor U3169 (N_3169,N_2104,N_2539);
nor U3170 (N_3170,N_2775,N_2533);
xor U3171 (N_3171,N_2905,N_2881);
nand U3172 (N_3172,N_2827,N_2057);
or U3173 (N_3173,N_2394,N_2441);
xor U3174 (N_3174,N_2741,N_2466);
and U3175 (N_3175,N_2149,N_2010);
and U3176 (N_3176,N_2674,N_2791);
nor U3177 (N_3177,N_2436,N_2765);
and U3178 (N_3178,N_2204,N_2892);
xor U3179 (N_3179,N_2083,N_2606);
nand U3180 (N_3180,N_2654,N_2237);
xor U3181 (N_3181,N_2963,N_2338);
nand U3182 (N_3182,N_2262,N_2956);
nand U3183 (N_3183,N_2499,N_2120);
xor U3184 (N_3184,N_2832,N_2546);
xnor U3185 (N_3185,N_2880,N_2525);
or U3186 (N_3186,N_2135,N_2352);
nor U3187 (N_3187,N_2542,N_2653);
nor U3188 (N_3188,N_2049,N_2838);
or U3189 (N_3189,N_2528,N_2923);
nand U3190 (N_3190,N_2380,N_2321);
or U3191 (N_3191,N_2235,N_2202);
and U3192 (N_3192,N_2852,N_2603);
and U3193 (N_3193,N_2904,N_2447);
and U3194 (N_3194,N_2781,N_2494);
nand U3195 (N_3195,N_2968,N_2399);
xor U3196 (N_3196,N_2712,N_2686);
and U3197 (N_3197,N_2732,N_2652);
or U3198 (N_3198,N_2541,N_2572);
and U3199 (N_3199,N_2859,N_2789);
xnor U3200 (N_3200,N_2005,N_2493);
nand U3201 (N_3201,N_2650,N_2814);
nor U3202 (N_3202,N_2580,N_2012);
nand U3203 (N_3203,N_2866,N_2233);
and U3204 (N_3204,N_2739,N_2924);
and U3205 (N_3205,N_2605,N_2706);
and U3206 (N_3206,N_2906,N_2655);
nand U3207 (N_3207,N_2748,N_2817);
and U3208 (N_3208,N_2414,N_2473);
and U3209 (N_3209,N_2878,N_2938);
nor U3210 (N_3210,N_2168,N_2872);
xnor U3211 (N_3211,N_2307,N_2330);
or U3212 (N_3212,N_2590,N_2936);
nor U3213 (N_3213,N_2961,N_2113);
nand U3214 (N_3214,N_2616,N_2687);
xnor U3215 (N_3215,N_2216,N_2087);
nor U3216 (N_3216,N_2306,N_2675);
or U3217 (N_3217,N_2794,N_2901);
and U3218 (N_3218,N_2175,N_2139);
or U3219 (N_3219,N_2234,N_2449);
and U3220 (N_3220,N_2780,N_2709);
nor U3221 (N_3221,N_2040,N_2361);
or U3222 (N_3222,N_2768,N_2027);
and U3223 (N_3223,N_2669,N_2184);
nor U3224 (N_3224,N_2598,N_2899);
or U3225 (N_3225,N_2908,N_2648);
and U3226 (N_3226,N_2625,N_2094);
and U3227 (N_3227,N_2769,N_2456);
nand U3228 (N_3228,N_2438,N_2515);
xor U3229 (N_3229,N_2110,N_2750);
or U3230 (N_3230,N_2577,N_2585);
nor U3231 (N_3231,N_2211,N_2952);
xnor U3232 (N_3232,N_2719,N_2705);
or U3233 (N_3233,N_2324,N_2544);
and U3234 (N_3234,N_2372,N_2230);
nand U3235 (N_3235,N_2159,N_2806);
xor U3236 (N_3236,N_2764,N_2620);
nor U3237 (N_3237,N_2304,N_2617);
xnor U3238 (N_3238,N_2993,N_2391);
or U3239 (N_3239,N_2846,N_2597);
xor U3240 (N_3240,N_2922,N_2555);
and U3241 (N_3241,N_2189,N_2312);
and U3242 (N_3242,N_2171,N_2063);
and U3243 (N_3243,N_2953,N_2637);
xnor U3244 (N_3244,N_2080,N_2670);
xor U3245 (N_3245,N_2198,N_2249);
and U3246 (N_3246,N_2055,N_2339);
or U3247 (N_3247,N_2717,N_2518);
nand U3248 (N_3248,N_2986,N_2209);
or U3249 (N_3249,N_2240,N_2164);
and U3250 (N_3250,N_2006,N_2479);
and U3251 (N_3251,N_2889,N_2437);
or U3252 (N_3252,N_2716,N_2504);
or U3253 (N_3253,N_2520,N_2464);
and U3254 (N_3254,N_2505,N_2983);
xor U3255 (N_3255,N_2927,N_2746);
nor U3256 (N_3256,N_2048,N_2988);
nand U3257 (N_3257,N_2972,N_2374);
or U3258 (N_3258,N_2751,N_2588);
xnor U3259 (N_3259,N_2459,N_2207);
nor U3260 (N_3260,N_2193,N_2691);
nor U3261 (N_3261,N_2995,N_2018);
or U3262 (N_3262,N_2405,N_2574);
nor U3263 (N_3263,N_2955,N_2749);
xnor U3264 (N_3264,N_2579,N_2443);
nor U3265 (N_3265,N_2608,N_2724);
and U3266 (N_3266,N_2738,N_2513);
nor U3267 (N_3267,N_2659,N_2822);
or U3268 (N_3268,N_2980,N_2392);
nor U3269 (N_3269,N_2401,N_2829);
or U3270 (N_3270,N_2460,N_2292);
xnor U3271 (N_3271,N_2041,N_2343);
xnor U3272 (N_3272,N_2105,N_2530);
or U3273 (N_3273,N_2267,N_2622);
xor U3274 (N_3274,N_2333,N_2645);
xor U3275 (N_3275,N_2317,N_2556);
or U3276 (N_3276,N_2795,N_2917);
nor U3277 (N_3277,N_2054,N_2695);
nand U3278 (N_3278,N_2962,N_2915);
and U3279 (N_3279,N_2666,N_2640);
nor U3280 (N_3280,N_2420,N_2957);
nand U3281 (N_3281,N_2668,N_2403);
and U3282 (N_3282,N_2759,N_2735);
nor U3283 (N_3283,N_2651,N_2757);
and U3284 (N_3284,N_2069,N_2604);
or U3285 (N_3285,N_2743,N_2121);
nand U3286 (N_3286,N_2680,N_2166);
and U3287 (N_3287,N_2444,N_2761);
and U3288 (N_3288,N_2767,N_2855);
xnor U3289 (N_3289,N_2595,N_2714);
and U3290 (N_3290,N_2697,N_2078);
nor U3291 (N_3291,N_2549,N_2476);
nor U3292 (N_3292,N_2845,N_2187);
and U3293 (N_3293,N_2064,N_2088);
nand U3294 (N_3294,N_2583,N_2707);
or U3295 (N_3295,N_2463,N_2910);
or U3296 (N_3296,N_2701,N_2812);
nor U3297 (N_3297,N_2557,N_2501);
xor U3298 (N_3298,N_2297,N_2607);
and U3299 (N_3299,N_2783,N_2909);
nand U3300 (N_3300,N_2115,N_2074);
or U3301 (N_3301,N_2346,N_2430);
xnor U3302 (N_3302,N_2229,N_2076);
or U3303 (N_3303,N_2887,N_2619);
or U3304 (N_3304,N_2786,N_2565);
xor U3305 (N_3305,N_2685,N_2932);
nand U3306 (N_3306,N_2704,N_2290);
nor U3307 (N_3307,N_2689,N_2295);
nand U3308 (N_3308,N_2816,N_2547);
and U3309 (N_3309,N_2071,N_2527);
nand U3310 (N_3310,N_2097,N_2073);
nor U3311 (N_3311,N_2623,N_2540);
xor U3312 (N_3312,N_2014,N_2482);
nor U3313 (N_3313,N_2543,N_2025);
and U3314 (N_3314,N_2944,N_2793);
or U3315 (N_3315,N_2425,N_2435);
nand U3316 (N_3316,N_2679,N_2481);
xor U3317 (N_3317,N_2966,N_2646);
nand U3318 (N_3318,N_2790,N_2179);
nor U3319 (N_3319,N_2861,N_2560);
xor U3320 (N_3320,N_2532,N_2673);
xnor U3321 (N_3321,N_2283,N_2571);
and U3322 (N_3322,N_2288,N_2422);
nand U3323 (N_3323,N_2660,N_2357);
nand U3324 (N_3324,N_2052,N_2635);
nand U3325 (N_3325,N_2302,N_2241);
nand U3326 (N_3326,N_2418,N_2726);
and U3327 (N_3327,N_2949,N_2411);
nor U3328 (N_3328,N_2612,N_2116);
nor U3329 (N_3329,N_2445,N_2516);
or U3330 (N_3330,N_2627,N_2170);
nor U3331 (N_3331,N_2964,N_2353);
nand U3332 (N_3332,N_2874,N_2404);
xor U3333 (N_3333,N_2756,N_2075);
nand U3334 (N_3334,N_2753,N_2138);
or U3335 (N_3335,N_2483,N_2090);
nand U3336 (N_3336,N_2992,N_2487);
xnor U3337 (N_3337,N_2140,N_2163);
or U3338 (N_3338,N_2489,N_2366);
xor U3339 (N_3339,N_2882,N_2581);
or U3340 (N_3340,N_2395,N_2636);
and U3341 (N_3341,N_2141,N_2851);
xnor U3342 (N_3342,N_2672,N_2061);
xnor U3343 (N_3343,N_2737,N_2835);
nor U3344 (N_3344,N_2354,N_2633);
or U3345 (N_3345,N_2879,N_2408);
and U3346 (N_3346,N_2551,N_2965);
xnor U3347 (N_3347,N_2853,N_2996);
nand U3348 (N_3348,N_2589,N_2875);
or U3349 (N_3349,N_2586,N_2658);
xnor U3350 (N_3350,N_2531,N_2309);
nand U3351 (N_3351,N_2611,N_2561);
xnor U3352 (N_3352,N_2773,N_2273);
and U3353 (N_3353,N_2900,N_2028);
and U3354 (N_3354,N_2232,N_2810);
nand U3355 (N_3355,N_2331,N_2937);
nor U3356 (N_3356,N_2255,N_2142);
xor U3357 (N_3357,N_2700,N_2918);
or U3358 (N_3358,N_2197,N_2841);
nand U3359 (N_3359,N_2095,N_2268);
or U3360 (N_3360,N_2575,N_2486);
xnor U3361 (N_3361,N_2613,N_2032);
nor U3362 (N_3362,N_2228,N_2225);
nor U3363 (N_3363,N_2718,N_2632);
xnor U3364 (N_3364,N_2760,N_2130);
xor U3365 (N_3365,N_2826,N_2248);
nor U3366 (N_3366,N_2387,N_2535);
and U3367 (N_3367,N_2802,N_2020);
nand U3368 (N_3368,N_2205,N_2451);
or U3369 (N_3369,N_2621,N_2491);
nor U3370 (N_3370,N_2036,N_2199);
nand U3371 (N_3371,N_2274,N_2345);
nand U3372 (N_3372,N_2856,N_2457);
or U3373 (N_3373,N_2158,N_2634);
xor U3374 (N_3374,N_2208,N_2186);
and U3375 (N_3375,N_2500,N_2933);
and U3376 (N_3376,N_2231,N_2471);
or U3377 (N_3377,N_2152,N_2318);
nand U3378 (N_3378,N_2364,N_2568);
xnor U3379 (N_3379,N_2725,N_2503);
nand U3380 (N_3380,N_2332,N_2440);
nor U3381 (N_3381,N_2217,N_2843);
or U3382 (N_3382,N_2145,N_2013);
or U3383 (N_3383,N_2183,N_2871);
xnor U3384 (N_3384,N_2647,N_2534);
or U3385 (N_3385,N_2562,N_2498);
xnor U3386 (N_3386,N_2772,N_2294);
nor U3387 (N_3387,N_2895,N_2808);
nand U3388 (N_3388,N_2877,N_2552);
nand U3389 (N_3389,N_2081,N_2252);
xor U3390 (N_3390,N_2973,N_2474);
nand U3391 (N_3391,N_2236,N_2929);
or U3392 (N_3392,N_2688,N_2998);
nor U3393 (N_3393,N_2157,N_2873);
or U3394 (N_3394,N_2432,N_2112);
xnor U3395 (N_3395,N_2223,N_2084);
or U3396 (N_3396,N_2342,N_2070);
xnor U3397 (N_3397,N_2303,N_2941);
nand U3398 (N_3398,N_2711,N_2291);
nor U3399 (N_3399,N_2111,N_2341);
nand U3400 (N_3400,N_2136,N_2916);
or U3401 (N_3401,N_2710,N_2951);
nor U3402 (N_3402,N_2172,N_2566);
xor U3403 (N_3403,N_2864,N_2251);
nand U3404 (N_3404,N_2059,N_2919);
xnor U3405 (N_3405,N_2434,N_2377);
or U3406 (N_3406,N_2890,N_2800);
nand U3407 (N_3407,N_2134,N_2296);
and U3408 (N_3408,N_2077,N_2624);
xnor U3409 (N_3409,N_2593,N_2336);
and U3410 (N_3410,N_2017,N_2942);
xor U3411 (N_3411,N_2433,N_2692);
nor U3412 (N_3412,N_2210,N_2260);
nor U3413 (N_3413,N_2072,N_2026);
nand U3414 (N_3414,N_2630,N_2609);
or U3415 (N_3415,N_2271,N_2833);
and U3416 (N_3416,N_2431,N_2276);
or U3417 (N_3417,N_2888,N_2488);
xnor U3418 (N_3418,N_2351,N_2897);
nand U3419 (N_3419,N_2413,N_2009);
or U3420 (N_3420,N_2155,N_2472);
or U3421 (N_3421,N_2015,N_2570);
nand U3422 (N_3422,N_2584,N_2277);
and U3423 (N_3423,N_2512,N_2848);
nand U3424 (N_3424,N_2153,N_2554);
nor U3425 (N_3425,N_2911,N_2950);
xor U3426 (N_3426,N_2379,N_2805);
and U3427 (N_3427,N_2266,N_2327);
or U3428 (N_3428,N_2242,N_2939);
nand U3429 (N_3429,N_2610,N_2019);
or U3430 (N_3430,N_2031,N_2356);
and U3431 (N_3431,N_2246,N_2270);
or U3432 (N_3432,N_2733,N_2243);
nand U3433 (N_3433,N_2227,N_2412);
xnor U3434 (N_3434,N_2984,N_2278);
nor U3435 (N_3435,N_2661,N_2222);
and U3436 (N_3436,N_2011,N_2469);
nor U3437 (N_3437,N_2681,N_2402);
nor U3438 (N_3438,N_2419,N_2161);
nor U3439 (N_3439,N_2976,N_2639);
xor U3440 (N_3440,N_2439,N_2523);
or U3441 (N_3441,N_2914,N_2190);
nand U3442 (N_3442,N_2894,N_2334);
or U3443 (N_3443,N_2427,N_2502);
xnor U3444 (N_3444,N_2977,N_2066);
and U3445 (N_3445,N_2109,N_2537);
nor U3446 (N_3446,N_2329,N_2344);
and U3447 (N_3447,N_2151,N_2079);
nor U3448 (N_3448,N_2825,N_2559);
or U3449 (N_3449,N_2677,N_2785);
nand U3450 (N_3450,N_2643,N_2284);
xnor U3451 (N_3451,N_2863,N_2424);
or U3452 (N_3452,N_2146,N_2188);
nor U3453 (N_3453,N_2506,N_2201);
nand U3454 (N_3454,N_2214,N_2478);
nand U3455 (N_3455,N_2930,N_2154);
nand U3456 (N_3456,N_2386,N_2522);
nand U3457 (N_3457,N_2389,N_2298);
nor U3458 (N_3458,N_2378,N_2224);
and U3459 (N_3459,N_2467,N_2771);
and U3460 (N_3460,N_2618,N_2397);
and U3461 (N_3461,N_2818,N_2050);
nand U3462 (N_3462,N_2124,N_2778);
nand U3463 (N_3463,N_2407,N_2811);
and U3464 (N_3464,N_2099,N_2987);
xnor U3465 (N_3465,N_2475,N_2300);
or U3466 (N_3466,N_2615,N_2301);
or U3467 (N_3467,N_2744,N_2614);
xnor U3468 (N_3468,N_2667,N_2799);
and U3469 (N_3469,N_2180,N_2450);
or U3470 (N_3470,N_2884,N_2455);
nand U3471 (N_3471,N_2860,N_2943);
or U3472 (N_3472,N_2103,N_2715);
nor U3473 (N_3473,N_2903,N_2355);
nand U3474 (N_3474,N_2167,N_2362);
or U3475 (N_3475,N_2160,N_2452);
nand U3476 (N_3476,N_2385,N_2181);
xnor U3477 (N_3477,N_2940,N_2708);
or U3478 (N_3478,N_2755,N_2156);
nand U3479 (N_3479,N_2946,N_2862);
xor U3480 (N_3480,N_2628,N_2734);
xor U3481 (N_3481,N_2137,N_2699);
nor U3482 (N_3482,N_2723,N_2129);
xnor U3483 (N_3483,N_2371,N_2926);
nor U3484 (N_3484,N_2058,N_2122);
nor U3485 (N_3485,N_2359,N_2657);
and U3486 (N_3486,N_2745,N_2000);
or U3487 (N_3487,N_2206,N_2285);
xor U3488 (N_3488,N_2117,N_2029);
or U3489 (N_3489,N_2410,N_2127);
xor U3490 (N_3490,N_2226,N_2663);
or U3491 (N_3491,N_2398,N_2971);
nor U3492 (N_3492,N_2970,N_2053);
and U3493 (N_3493,N_2857,N_2368);
or U3494 (N_3494,N_2979,N_2840);
or U3495 (N_3495,N_2830,N_2323);
nor U3496 (N_3496,N_2098,N_2021);
xnor U3497 (N_3497,N_2393,N_2824);
or U3498 (N_3498,N_2269,N_2898);
and U3499 (N_3499,N_2985,N_2178);
or U3500 (N_3500,N_2870,N_2282);
and U3501 (N_3501,N_2531,N_2931);
xnor U3502 (N_3502,N_2413,N_2275);
nand U3503 (N_3503,N_2955,N_2624);
xor U3504 (N_3504,N_2504,N_2864);
and U3505 (N_3505,N_2393,N_2980);
xor U3506 (N_3506,N_2381,N_2388);
nor U3507 (N_3507,N_2156,N_2392);
nand U3508 (N_3508,N_2455,N_2371);
and U3509 (N_3509,N_2683,N_2181);
or U3510 (N_3510,N_2469,N_2716);
xor U3511 (N_3511,N_2455,N_2413);
xnor U3512 (N_3512,N_2694,N_2944);
or U3513 (N_3513,N_2871,N_2079);
nor U3514 (N_3514,N_2877,N_2906);
nor U3515 (N_3515,N_2624,N_2127);
and U3516 (N_3516,N_2013,N_2281);
nor U3517 (N_3517,N_2157,N_2421);
and U3518 (N_3518,N_2760,N_2549);
or U3519 (N_3519,N_2020,N_2923);
xnor U3520 (N_3520,N_2818,N_2721);
and U3521 (N_3521,N_2579,N_2269);
nor U3522 (N_3522,N_2497,N_2635);
xnor U3523 (N_3523,N_2828,N_2795);
xnor U3524 (N_3524,N_2675,N_2117);
and U3525 (N_3525,N_2171,N_2574);
xor U3526 (N_3526,N_2746,N_2903);
xor U3527 (N_3527,N_2367,N_2449);
nand U3528 (N_3528,N_2400,N_2048);
nand U3529 (N_3529,N_2728,N_2524);
and U3530 (N_3530,N_2303,N_2615);
or U3531 (N_3531,N_2754,N_2017);
xor U3532 (N_3532,N_2057,N_2888);
nor U3533 (N_3533,N_2266,N_2295);
or U3534 (N_3534,N_2356,N_2201);
nand U3535 (N_3535,N_2488,N_2702);
or U3536 (N_3536,N_2776,N_2595);
and U3537 (N_3537,N_2151,N_2538);
or U3538 (N_3538,N_2067,N_2846);
and U3539 (N_3539,N_2613,N_2310);
or U3540 (N_3540,N_2462,N_2872);
nand U3541 (N_3541,N_2543,N_2076);
or U3542 (N_3542,N_2080,N_2054);
nand U3543 (N_3543,N_2508,N_2230);
xor U3544 (N_3544,N_2941,N_2638);
nand U3545 (N_3545,N_2458,N_2870);
xnor U3546 (N_3546,N_2578,N_2295);
or U3547 (N_3547,N_2485,N_2638);
xor U3548 (N_3548,N_2110,N_2223);
xnor U3549 (N_3549,N_2643,N_2528);
nor U3550 (N_3550,N_2643,N_2572);
nand U3551 (N_3551,N_2764,N_2740);
xnor U3552 (N_3552,N_2771,N_2256);
and U3553 (N_3553,N_2357,N_2572);
or U3554 (N_3554,N_2962,N_2109);
nand U3555 (N_3555,N_2260,N_2602);
nand U3556 (N_3556,N_2215,N_2736);
or U3557 (N_3557,N_2492,N_2959);
nand U3558 (N_3558,N_2703,N_2613);
nand U3559 (N_3559,N_2525,N_2780);
xor U3560 (N_3560,N_2348,N_2819);
xor U3561 (N_3561,N_2478,N_2615);
xor U3562 (N_3562,N_2077,N_2087);
nand U3563 (N_3563,N_2412,N_2828);
xor U3564 (N_3564,N_2904,N_2672);
and U3565 (N_3565,N_2457,N_2123);
nand U3566 (N_3566,N_2116,N_2242);
xnor U3567 (N_3567,N_2590,N_2805);
xnor U3568 (N_3568,N_2979,N_2087);
or U3569 (N_3569,N_2215,N_2083);
or U3570 (N_3570,N_2801,N_2097);
nor U3571 (N_3571,N_2428,N_2814);
nor U3572 (N_3572,N_2180,N_2631);
or U3573 (N_3573,N_2091,N_2716);
and U3574 (N_3574,N_2733,N_2315);
nand U3575 (N_3575,N_2700,N_2806);
xor U3576 (N_3576,N_2997,N_2313);
nand U3577 (N_3577,N_2755,N_2845);
and U3578 (N_3578,N_2268,N_2910);
or U3579 (N_3579,N_2635,N_2122);
xnor U3580 (N_3580,N_2710,N_2248);
or U3581 (N_3581,N_2931,N_2462);
nand U3582 (N_3582,N_2614,N_2681);
nand U3583 (N_3583,N_2914,N_2980);
nor U3584 (N_3584,N_2262,N_2426);
nand U3585 (N_3585,N_2909,N_2256);
nor U3586 (N_3586,N_2758,N_2153);
nand U3587 (N_3587,N_2552,N_2453);
nor U3588 (N_3588,N_2840,N_2724);
and U3589 (N_3589,N_2857,N_2836);
and U3590 (N_3590,N_2400,N_2823);
nor U3591 (N_3591,N_2070,N_2884);
xnor U3592 (N_3592,N_2599,N_2828);
and U3593 (N_3593,N_2300,N_2738);
and U3594 (N_3594,N_2722,N_2604);
and U3595 (N_3595,N_2071,N_2202);
or U3596 (N_3596,N_2305,N_2974);
xnor U3597 (N_3597,N_2030,N_2528);
or U3598 (N_3598,N_2043,N_2501);
or U3599 (N_3599,N_2289,N_2979);
nor U3600 (N_3600,N_2640,N_2974);
nor U3601 (N_3601,N_2163,N_2742);
or U3602 (N_3602,N_2081,N_2334);
and U3603 (N_3603,N_2301,N_2162);
and U3604 (N_3604,N_2454,N_2950);
and U3605 (N_3605,N_2041,N_2360);
nand U3606 (N_3606,N_2693,N_2644);
xnor U3607 (N_3607,N_2199,N_2790);
nor U3608 (N_3608,N_2220,N_2534);
and U3609 (N_3609,N_2961,N_2478);
or U3610 (N_3610,N_2947,N_2509);
xnor U3611 (N_3611,N_2565,N_2774);
nand U3612 (N_3612,N_2366,N_2459);
xnor U3613 (N_3613,N_2848,N_2940);
nand U3614 (N_3614,N_2294,N_2729);
and U3615 (N_3615,N_2907,N_2115);
and U3616 (N_3616,N_2140,N_2039);
or U3617 (N_3617,N_2139,N_2019);
nor U3618 (N_3618,N_2913,N_2603);
nor U3619 (N_3619,N_2842,N_2205);
xnor U3620 (N_3620,N_2629,N_2258);
xor U3621 (N_3621,N_2714,N_2072);
nand U3622 (N_3622,N_2941,N_2702);
xnor U3623 (N_3623,N_2593,N_2869);
nand U3624 (N_3624,N_2440,N_2340);
nand U3625 (N_3625,N_2480,N_2942);
or U3626 (N_3626,N_2164,N_2080);
or U3627 (N_3627,N_2547,N_2616);
and U3628 (N_3628,N_2791,N_2389);
xnor U3629 (N_3629,N_2491,N_2045);
xnor U3630 (N_3630,N_2529,N_2728);
nand U3631 (N_3631,N_2115,N_2460);
or U3632 (N_3632,N_2763,N_2627);
nor U3633 (N_3633,N_2671,N_2512);
or U3634 (N_3634,N_2865,N_2015);
nand U3635 (N_3635,N_2481,N_2967);
nand U3636 (N_3636,N_2660,N_2710);
or U3637 (N_3637,N_2718,N_2741);
nand U3638 (N_3638,N_2048,N_2934);
nand U3639 (N_3639,N_2491,N_2142);
and U3640 (N_3640,N_2237,N_2752);
nand U3641 (N_3641,N_2452,N_2549);
and U3642 (N_3642,N_2621,N_2287);
and U3643 (N_3643,N_2148,N_2289);
and U3644 (N_3644,N_2450,N_2735);
and U3645 (N_3645,N_2239,N_2943);
and U3646 (N_3646,N_2845,N_2939);
xor U3647 (N_3647,N_2985,N_2414);
or U3648 (N_3648,N_2887,N_2768);
xnor U3649 (N_3649,N_2438,N_2682);
or U3650 (N_3650,N_2396,N_2488);
nand U3651 (N_3651,N_2896,N_2073);
nor U3652 (N_3652,N_2044,N_2217);
nor U3653 (N_3653,N_2792,N_2131);
or U3654 (N_3654,N_2761,N_2098);
xnor U3655 (N_3655,N_2823,N_2301);
and U3656 (N_3656,N_2957,N_2674);
and U3657 (N_3657,N_2311,N_2670);
xnor U3658 (N_3658,N_2779,N_2783);
or U3659 (N_3659,N_2773,N_2201);
nor U3660 (N_3660,N_2248,N_2398);
or U3661 (N_3661,N_2586,N_2314);
and U3662 (N_3662,N_2209,N_2885);
nor U3663 (N_3663,N_2922,N_2396);
and U3664 (N_3664,N_2423,N_2563);
nand U3665 (N_3665,N_2631,N_2759);
nand U3666 (N_3666,N_2970,N_2333);
xnor U3667 (N_3667,N_2741,N_2511);
nor U3668 (N_3668,N_2399,N_2824);
xor U3669 (N_3669,N_2579,N_2215);
or U3670 (N_3670,N_2135,N_2137);
and U3671 (N_3671,N_2535,N_2884);
xor U3672 (N_3672,N_2860,N_2390);
or U3673 (N_3673,N_2283,N_2530);
or U3674 (N_3674,N_2513,N_2899);
nor U3675 (N_3675,N_2710,N_2046);
nand U3676 (N_3676,N_2120,N_2538);
nor U3677 (N_3677,N_2816,N_2926);
nor U3678 (N_3678,N_2916,N_2599);
xor U3679 (N_3679,N_2694,N_2930);
nor U3680 (N_3680,N_2775,N_2929);
and U3681 (N_3681,N_2956,N_2237);
nor U3682 (N_3682,N_2517,N_2537);
nand U3683 (N_3683,N_2160,N_2582);
nand U3684 (N_3684,N_2331,N_2414);
and U3685 (N_3685,N_2630,N_2490);
or U3686 (N_3686,N_2979,N_2481);
nor U3687 (N_3687,N_2234,N_2444);
nor U3688 (N_3688,N_2195,N_2625);
nand U3689 (N_3689,N_2168,N_2878);
xnor U3690 (N_3690,N_2698,N_2718);
xor U3691 (N_3691,N_2223,N_2687);
nor U3692 (N_3692,N_2492,N_2803);
xnor U3693 (N_3693,N_2452,N_2886);
xor U3694 (N_3694,N_2623,N_2499);
or U3695 (N_3695,N_2148,N_2422);
nand U3696 (N_3696,N_2228,N_2911);
and U3697 (N_3697,N_2996,N_2994);
or U3698 (N_3698,N_2295,N_2705);
or U3699 (N_3699,N_2705,N_2445);
or U3700 (N_3700,N_2499,N_2062);
and U3701 (N_3701,N_2912,N_2011);
nor U3702 (N_3702,N_2303,N_2945);
or U3703 (N_3703,N_2571,N_2595);
nand U3704 (N_3704,N_2052,N_2278);
or U3705 (N_3705,N_2483,N_2227);
or U3706 (N_3706,N_2024,N_2570);
nand U3707 (N_3707,N_2767,N_2351);
nor U3708 (N_3708,N_2037,N_2346);
nor U3709 (N_3709,N_2631,N_2987);
or U3710 (N_3710,N_2586,N_2968);
or U3711 (N_3711,N_2283,N_2046);
nand U3712 (N_3712,N_2392,N_2125);
and U3713 (N_3713,N_2997,N_2134);
nand U3714 (N_3714,N_2155,N_2314);
nor U3715 (N_3715,N_2453,N_2742);
and U3716 (N_3716,N_2795,N_2298);
nand U3717 (N_3717,N_2535,N_2270);
nor U3718 (N_3718,N_2328,N_2580);
or U3719 (N_3719,N_2561,N_2163);
or U3720 (N_3720,N_2499,N_2522);
and U3721 (N_3721,N_2486,N_2204);
nand U3722 (N_3722,N_2781,N_2904);
or U3723 (N_3723,N_2306,N_2495);
or U3724 (N_3724,N_2737,N_2999);
nand U3725 (N_3725,N_2050,N_2650);
nand U3726 (N_3726,N_2388,N_2919);
xor U3727 (N_3727,N_2501,N_2315);
nor U3728 (N_3728,N_2533,N_2357);
or U3729 (N_3729,N_2791,N_2278);
xor U3730 (N_3730,N_2983,N_2918);
nand U3731 (N_3731,N_2072,N_2471);
nor U3732 (N_3732,N_2870,N_2482);
xor U3733 (N_3733,N_2682,N_2291);
or U3734 (N_3734,N_2388,N_2944);
and U3735 (N_3735,N_2220,N_2118);
xor U3736 (N_3736,N_2220,N_2119);
nand U3737 (N_3737,N_2944,N_2049);
and U3738 (N_3738,N_2958,N_2843);
and U3739 (N_3739,N_2461,N_2074);
xor U3740 (N_3740,N_2984,N_2550);
and U3741 (N_3741,N_2204,N_2299);
or U3742 (N_3742,N_2353,N_2794);
xnor U3743 (N_3743,N_2609,N_2324);
nor U3744 (N_3744,N_2626,N_2740);
nand U3745 (N_3745,N_2352,N_2420);
xor U3746 (N_3746,N_2067,N_2336);
nor U3747 (N_3747,N_2798,N_2547);
nand U3748 (N_3748,N_2036,N_2736);
xnor U3749 (N_3749,N_2120,N_2610);
nand U3750 (N_3750,N_2210,N_2440);
nand U3751 (N_3751,N_2140,N_2077);
nand U3752 (N_3752,N_2815,N_2237);
and U3753 (N_3753,N_2884,N_2345);
or U3754 (N_3754,N_2266,N_2658);
or U3755 (N_3755,N_2852,N_2949);
nand U3756 (N_3756,N_2068,N_2554);
and U3757 (N_3757,N_2607,N_2299);
nor U3758 (N_3758,N_2818,N_2491);
nand U3759 (N_3759,N_2473,N_2440);
xnor U3760 (N_3760,N_2995,N_2912);
and U3761 (N_3761,N_2455,N_2700);
and U3762 (N_3762,N_2652,N_2094);
nand U3763 (N_3763,N_2007,N_2592);
nor U3764 (N_3764,N_2377,N_2421);
and U3765 (N_3765,N_2939,N_2035);
nand U3766 (N_3766,N_2168,N_2296);
nor U3767 (N_3767,N_2337,N_2448);
nand U3768 (N_3768,N_2841,N_2326);
nor U3769 (N_3769,N_2859,N_2529);
and U3770 (N_3770,N_2031,N_2277);
and U3771 (N_3771,N_2196,N_2825);
or U3772 (N_3772,N_2783,N_2110);
nor U3773 (N_3773,N_2092,N_2540);
nor U3774 (N_3774,N_2639,N_2645);
xor U3775 (N_3775,N_2741,N_2682);
and U3776 (N_3776,N_2005,N_2201);
and U3777 (N_3777,N_2856,N_2206);
nor U3778 (N_3778,N_2905,N_2197);
nand U3779 (N_3779,N_2919,N_2247);
nand U3780 (N_3780,N_2883,N_2772);
or U3781 (N_3781,N_2826,N_2456);
or U3782 (N_3782,N_2189,N_2368);
or U3783 (N_3783,N_2934,N_2745);
and U3784 (N_3784,N_2063,N_2704);
and U3785 (N_3785,N_2775,N_2970);
or U3786 (N_3786,N_2799,N_2057);
nand U3787 (N_3787,N_2883,N_2829);
xnor U3788 (N_3788,N_2789,N_2035);
nand U3789 (N_3789,N_2192,N_2289);
xnor U3790 (N_3790,N_2895,N_2742);
nor U3791 (N_3791,N_2239,N_2326);
nor U3792 (N_3792,N_2199,N_2457);
or U3793 (N_3793,N_2763,N_2749);
nor U3794 (N_3794,N_2165,N_2493);
nand U3795 (N_3795,N_2358,N_2735);
and U3796 (N_3796,N_2321,N_2861);
nand U3797 (N_3797,N_2332,N_2708);
nand U3798 (N_3798,N_2662,N_2888);
nor U3799 (N_3799,N_2514,N_2854);
nand U3800 (N_3800,N_2303,N_2758);
and U3801 (N_3801,N_2850,N_2860);
xor U3802 (N_3802,N_2681,N_2236);
or U3803 (N_3803,N_2366,N_2771);
nand U3804 (N_3804,N_2140,N_2744);
nor U3805 (N_3805,N_2529,N_2350);
nor U3806 (N_3806,N_2176,N_2981);
xor U3807 (N_3807,N_2534,N_2401);
nand U3808 (N_3808,N_2908,N_2849);
or U3809 (N_3809,N_2136,N_2069);
nand U3810 (N_3810,N_2197,N_2152);
and U3811 (N_3811,N_2940,N_2790);
nand U3812 (N_3812,N_2133,N_2927);
or U3813 (N_3813,N_2394,N_2565);
nor U3814 (N_3814,N_2977,N_2661);
or U3815 (N_3815,N_2483,N_2415);
or U3816 (N_3816,N_2833,N_2589);
nand U3817 (N_3817,N_2282,N_2571);
and U3818 (N_3818,N_2046,N_2099);
xnor U3819 (N_3819,N_2392,N_2919);
nand U3820 (N_3820,N_2357,N_2226);
and U3821 (N_3821,N_2793,N_2939);
or U3822 (N_3822,N_2479,N_2980);
or U3823 (N_3823,N_2043,N_2611);
and U3824 (N_3824,N_2507,N_2762);
nor U3825 (N_3825,N_2788,N_2987);
xnor U3826 (N_3826,N_2902,N_2977);
nor U3827 (N_3827,N_2684,N_2141);
and U3828 (N_3828,N_2783,N_2725);
nor U3829 (N_3829,N_2609,N_2257);
and U3830 (N_3830,N_2059,N_2142);
or U3831 (N_3831,N_2198,N_2248);
nand U3832 (N_3832,N_2379,N_2958);
nand U3833 (N_3833,N_2821,N_2834);
nand U3834 (N_3834,N_2561,N_2547);
nand U3835 (N_3835,N_2176,N_2734);
xnor U3836 (N_3836,N_2494,N_2714);
nor U3837 (N_3837,N_2952,N_2306);
nor U3838 (N_3838,N_2674,N_2754);
xnor U3839 (N_3839,N_2976,N_2486);
nor U3840 (N_3840,N_2500,N_2350);
xnor U3841 (N_3841,N_2291,N_2273);
nor U3842 (N_3842,N_2376,N_2402);
nor U3843 (N_3843,N_2861,N_2529);
nand U3844 (N_3844,N_2507,N_2676);
or U3845 (N_3845,N_2997,N_2910);
or U3846 (N_3846,N_2672,N_2502);
xor U3847 (N_3847,N_2749,N_2903);
nor U3848 (N_3848,N_2126,N_2154);
or U3849 (N_3849,N_2401,N_2114);
or U3850 (N_3850,N_2268,N_2444);
nand U3851 (N_3851,N_2421,N_2341);
xnor U3852 (N_3852,N_2243,N_2330);
or U3853 (N_3853,N_2367,N_2067);
and U3854 (N_3854,N_2824,N_2068);
nand U3855 (N_3855,N_2947,N_2106);
or U3856 (N_3856,N_2502,N_2750);
nor U3857 (N_3857,N_2535,N_2382);
and U3858 (N_3858,N_2184,N_2842);
nor U3859 (N_3859,N_2033,N_2623);
nand U3860 (N_3860,N_2716,N_2486);
or U3861 (N_3861,N_2317,N_2338);
nor U3862 (N_3862,N_2847,N_2362);
or U3863 (N_3863,N_2765,N_2824);
nand U3864 (N_3864,N_2801,N_2743);
and U3865 (N_3865,N_2325,N_2207);
or U3866 (N_3866,N_2002,N_2990);
and U3867 (N_3867,N_2411,N_2531);
xor U3868 (N_3868,N_2151,N_2899);
nor U3869 (N_3869,N_2544,N_2593);
xnor U3870 (N_3870,N_2281,N_2111);
or U3871 (N_3871,N_2786,N_2107);
nand U3872 (N_3872,N_2765,N_2955);
nand U3873 (N_3873,N_2528,N_2688);
xnor U3874 (N_3874,N_2811,N_2242);
or U3875 (N_3875,N_2968,N_2729);
nor U3876 (N_3876,N_2206,N_2464);
and U3877 (N_3877,N_2976,N_2591);
nor U3878 (N_3878,N_2429,N_2353);
nand U3879 (N_3879,N_2369,N_2029);
xnor U3880 (N_3880,N_2186,N_2300);
xnor U3881 (N_3881,N_2921,N_2344);
nor U3882 (N_3882,N_2198,N_2924);
nand U3883 (N_3883,N_2767,N_2657);
nand U3884 (N_3884,N_2739,N_2663);
and U3885 (N_3885,N_2483,N_2812);
or U3886 (N_3886,N_2262,N_2108);
or U3887 (N_3887,N_2852,N_2216);
nand U3888 (N_3888,N_2875,N_2644);
xor U3889 (N_3889,N_2651,N_2458);
xor U3890 (N_3890,N_2960,N_2447);
nand U3891 (N_3891,N_2411,N_2126);
nor U3892 (N_3892,N_2599,N_2979);
and U3893 (N_3893,N_2258,N_2714);
nand U3894 (N_3894,N_2933,N_2517);
xor U3895 (N_3895,N_2857,N_2694);
xor U3896 (N_3896,N_2337,N_2818);
nor U3897 (N_3897,N_2708,N_2104);
or U3898 (N_3898,N_2259,N_2241);
and U3899 (N_3899,N_2807,N_2699);
and U3900 (N_3900,N_2554,N_2931);
or U3901 (N_3901,N_2014,N_2757);
and U3902 (N_3902,N_2712,N_2655);
or U3903 (N_3903,N_2431,N_2556);
nor U3904 (N_3904,N_2035,N_2667);
xnor U3905 (N_3905,N_2383,N_2178);
xnor U3906 (N_3906,N_2062,N_2802);
and U3907 (N_3907,N_2625,N_2693);
xor U3908 (N_3908,N_2504,N_2082);
xnor U3909 (N_3909,N_2746,N_2865);
and U3910 (N_3910,N_2854,N_2335);
nor U3911 (N_3911,N_2882,N_2197);
xnor U3912 (N_3912,N_2609,N_2245);
or U3913 (N_3913,N_2324,N_2751);
nor U3914 (N_3914,N_2866,N_2183);
nor U3915 (N_3915,N_2080,N_2396);
and U3916 (N_3916,N_2666,N_2350);
nand U3917 (N_3917,N_2635,N_2231);
or U3918 (N_3918,N_2775,N_2154);
or U3919 (N_3919,N_2177,N_2664);
nand U3920 (N_3920,N_2794,N_2141);
or U3921 (N_3921,N_2042,N_2175);
xor U3922 (N_3922,N_2945,N_2326);
nand U3923 (N_3923,N_2314,N_2808);
nor U3924 (N_3924,N_2835,N_2370);
and U3925 (N_3925,N_2728,N_2986);
xnor U3926 (N_3926,N_2440,N_2513);
or U3927 (N_3927,N_2856,N_2325);
or U3928 (N_3928,N_2862,N_2489);
nand U3929 (N_3929,N_2593,N_2061);
nand U3930 (N_3930,N_2258,N_2381);
and U3931 (N_3931,N_2066,N_2548);
or U3932 (N_3932,N_2320,N_2139);
xnor U3933 (N_3933,N_2411,N_2825);
or U3934 (N_3934,N_2802,N_2339);
and U3935 (N_3935,N_2459,N_2349);
and U3936 (N_3936,N_2952,N_2894);
or U3937 (N_3937,N_2544,N_2062);
and U3938 (N_3938,N_2269,N_2222);
and U3939 (N_3939,N_2128,N_2706);
and U3940 (N_3940,N_2394,N_2895);
xnor U3941 (N_3941,N_2575,N_2733);
nand U3942 (N_3942,N_2561,N_2760);
and U3943 (N_3943,N_2198,N_2602);
and U3944 (N_3944,N_2836,N_2775);
nand U3945 (N_3945,N_2031,N_2408);
xnor U3946 (N_3946,N_2804,N_2344);
nor U3947 (N_3947,N_2101,N_2256);
nor U3948 (N_3948,N_2516,N_2263);
and U3949 (N_3949,N_2924,N_2401);
xor U3950 (N_3950,N_2252,N_2984);
or U3951 (N_3951,N_2141,N_2064);
and U3952 (N_3952,N_2682,N_2300);
or U3953 (N_3953,N_2275,N_2175);
and U3954 (N_3954,N_2935,N_2358);
and U3955 (N_3955,N_2829,N_2045);
xor U3956 (N_3956,N_2690,N_2960);
nand U3957 (N_3957,N_2595,N_2116);
nor U3958 (N_3958,N_2820,N_2807);
nor U3959 (N_3959,N_2332,N_2186);
nand U3960 (N_3960,N_2738,N_2021);
nand U3961 (N_3961,N_2720,N_2312);
nand U3962 (N_3962,N_2289,N_2061);
nor U3963 (N_3963,N_2748,N_2068);
or U3964 (N_3964,N_2292,N_2284);
nor U3965 (N_3965,N_2918,N_2039);
nor U3966 (N_3966,N_2719,N_2499);
or U3967 (N_3967,N_2965,N_2665);
nand U3968 (N_3968,N_2291,N_2933);
xnor U3969 (N_3969,N_2840,N_2366);
or U3970 (N_3970,N_2033,N_2900);
nand U3971 (N_3971,N_2596,N_2267);
xnor U3972 (N_3972,N_2469,N_2077);
nor U3973 (N_3973,N_2456,N_2658);
or U3974 (N_3974,N_2174,N_2128);
nor U3975 (N_3975,N_2232,N_2496);
and U3976 (N_3976,N_2896,N_2724);
xor U3977 (N_3977,N_2318,N_2112);
nand U3978 (N_3978,N_2402,N_2584);
nand U3979 (N_3979,N_2901,N_2433);
nand U3980 (N_3980,N_2980,N_2751);
nor U3981 (N_3981,N_2429,N_2599);
nand U3982 (N_3982,N_2216,N_2618);
xnor U3983 (N_3983,N_2096,N_2046);
xnor U3984 (N_3984,N_2952,N_2015);
and U3985 (N_3985,N_2047,N_2322);
nand U3986 (N_3986,N_2047,N_2159);
and U3987 (N_3987,N_2678,N_2193);
nand U3988 (N_3988,N_2669,N_2125);
xor U3989 (N_3989,N_2430,N_2154);
nand U3990 (N_3990,N_2940,N_2716);
nor U3991 (N_3991,N_2309,N_2779);
nand U3992 (N_3992,N_2590,N_2270);
and U3993 (N_3993,N_2956,N_2526);
nand U3994 (N_3994,N_2559,N_2464);
and U3995 (N_3995,N_2908,N_2075);
and U3996 (N_3996,N_2774,N_2215);
nor U3997 (N_3997,N_2655,N_2456);
nand U3998 (N_3998,N_2996,N_2234);
or U3999 (N_3999,N_2790,N_2439);
nand U4000 (N_4000,N_3908,N_3108);
nand U4001 (N_4001,N_3030,N_3243);
or U4002 (N_4002,N_3647,N_3023);
and U4003 (N_4003,N_3858,N_3754);
xor U4004 (N_4004,N_3360,N_3233);
and U4005 (N_4005,N_3819,N_3280);
xnor U4006 (N_4006,N_3800,N_3135);
nand U4007 (N_4007,N_3864,N_3015);
nand U4008 (N_4008,N_3551,N_3724);
nand U4009 (N_4009,N_3425,N_3902);
or U4010 (N_4010,N_3056,N_3466);
nand U4011 (N_4011,N_3500,N_3198);
nand U4012 (N_4012,N_3658,N_3315);
and U4013 (N_4013,N_3675,N_3103);
nor U4014 (N_4014,N_3751,N_3296);
or U4015 (N_4015,N_3561,N_3531);
xor U4016 (N_4016,N_3123,N_3119);
nand U4017 (N_4017,N_3390,N_3041);
or U4018 (N_4018,N_3283,N_3447);
xor U4019 (N_4019,N_3455,N_3672);
and U4020 (N_4020,N_3710,N_3320);
xnor U4021 (N_4021,N_3072,N_3017);
nor U4022 (N_4022,N_3657,N_3225);
nand U4023 (N_4023,N_3837,N_3345);
and U4024 (N_4024,N_3095,N_3289);
xnor U4025 (N_4025,N_3768,N_3856);
xnor U4026 (N_4026,N_3701,N_3730);
xor U4027 (N_4027,N_3610,N_3996);
nor U4028 (N_4028,N_3388,N_3354);
nor U4029 (N_4029,N_3480,N_3204);
or U4030 (N_4030,N_3890,N_3544);
or U4031 (N_4031,N_3887,N_3536);
xnor U4032 (N_4032,N_3293,N_3039);
nor U4033 (N_4033,N_3840,N_3763);
and U4034 (N_4034,N_3779,N_3138);
nand U4035 (N_4035,N_3679,N_3736);
nand U4036 (N_4036,N_3308,N_3980);
nor U4037 (N_4037,N_3275,N_3579);
nor U4038 (N_4038,N_3891,N_3992);
or U4039 (N_4039,N_3967,N_3300);
or U4040 (N_4040,N_3196,N_3405);
and U4041 (N_4041,N_3146,N_3916);
xor U4042 (N_4042,N_3001,N_3033);
or U4043 (N_4043,N_3997,N_3912);
and U4044 (N_4044,N_3968,N_3562);
xor U4045 (N_4045,N_3875,N_3825);
nand U4046 (N_4046,N_3370,N_3978);
xor U4047 (N_4047,N_3230,N_3594);
and U4048 (N_4048,N_3708,N_3118);
or U4049 (N_4049,N_3437,N_3598);
xor U4050 (N_4050,N_3219,N_3650);
xnor U4051 (N_4051,N_3442,N_3934);
nor U4052 (N_4052,N_3584,N_3575);
and U4053 (N_4053,N_3974,N_3136);
nor U4054 (N_4054,N_3646,N_3660);
and U4055 (N_4055,N_3845,N_3306);
nor U4056 (N_4056,N_3347,N_3120);
nor U4057 (N_4057,N_3712,N_3319);
xnor U4058 (N_4058,N_3060,N_3478);
or U4059 (N_4059,N_3578,N_3559);
xor U4060 (N_4060,N_3424,N_3543);
or U4061 (N_4061,N_3915,N_3951);
nor U4062 (N_4062,N_3873,N_3704);
or U4063 (N_4063,N_3782,N_3117);
or U4064 (N_4064,N_3324,N_3178);
nor U4065 (N_4065,N_3924,N_3629);
and U4066 (N_4066,N_3317,N_3218);
and U4067 (N_4067,N_3600,N_3541);
xnor U4068 (N_4068,N_3372,N_3250);
nor U4069 (N_4069,N_3142,N_3385);
and U4070 (N_4070,N_3294,N_3008);
and U4071 (N_4071,N_3130,N_3511);
or U4072 (N_4072,N_3369,N_3412);
nor U4073 (N_4073,N_3674,N_3400);
nor U4074 (N_4074,N_3638,N_3426);
nor U4075 (N_4075,N_3316,N_3731);
and U4076 (N_4076,N_3451,N_3334);
nor U4077 (N_4077,N_3419,N_3247);
xor U4078 (N_4078,N_3262,N_3242);
xnor U4079 (N_4079,N_3038,N_3376);
nand U4080 (N_4080,N_3770,N_3078);
xnor U4081 (N_4081,N_3663,N_3959);
or U4082 (N_4082,N_3277,N_3666);
nor U4083 (N_4083,N_3036,N_3014);
nand U4084 (N_4084,N_3756,N_3645);
and U4085 (N_4085,N_3711,N_3605);
nor U4086 (N_4086,N_3778,N_3127);
nor U4087 (N_4087,N_3668,N_3154);
nor U4088 (N_4088,N_3043,N_3506);
xor U4089 (N_4089,N_3841,N_3947);
nor U4090 (N_4090,N_3504,N_3012);
nor U4091 (N_4091,N_3789,N_3172);
nor U4092 (N_4092,N_3749,N_3299);
or U4093 (N_4093,N_3486,N_3410);
or U4094 (N_4094,N_3199,N_3568);
nor U4095 (N_4095,N_3362,N_3615);
xor U4096 (N_4096,N_3796,N_3395);
nor U4097 (N_4097,N_3368,N_3384);
or U4098 (N_4098,N_3682,N_3279);
nand U4099 (N_4099,N_3878,N_3070);
xnor U4100 (N_4100,N_3281,N_3530);
or U4101 (N_4101,N_3469,N_3398);
xor U4102 (N_4102,N_3539,N_3642);
xor U4103 (N_4103,N_3088,N_3440);
or U4104 (N_4104,N_3152,N_3352);
xnor U4105 (N_4105,N_3031,N_3583);
xor U4106 (N_4106,N_3823,N_3684);
nand U4107 (N_4107,N_3683,N_3367);
and U4108 (N_4108,N_3322,N_3827);
nor U4109 (N_4109,N_3507,N_3760);
xnor U4110 (N_4110,N_3702,N_3637);
and U4111 (N_4111,N_3689,N_3415);
and U4112 (N_4112,N_3581,N_3599);
or U4113 (N_4113,N_3695,N_3465);
nand U4114 (N_4114,N_3098,N_3641);
xor U4115 (N_4115,N_3170,N_3555);
nand U4116 (N_4116,N_3804,N_3874);
nor U4117 (N_4117,N_3591,N_3574);
or U4118 (N_4118,N_3365,N_3810);
or U4119 (N_4119,N_3175,N_3972);
nor U4120 (N_4120,N_3656,N_3991);
nor U4121 (N_4121,N_3066,N_3595);
nand U4122 (N_4122,N_3457,N_3560);
xor U4123 (N_4123,N_3470,N_3240);
xor U4124 (N_4124,N_3255,N_3776);
nor U4125 (N_4125,N_3732,N_3512);
xnor U4126 (N_4126,N_3417,N_3257);
xnor U4127 (N_4127,N_3328,N_3743);
xor U4128 (N_4128,N_3502,N_3490);
and U4129 (N_4129,N_3402,N_3721);
xnor U4130 (N_4130,N_3314,N_3807);
or U4131 (N_4131,N_3636,N_3818);
nand U4132 (N_4132,N_3025,N_3083);
xnor U4133 (N_4133,N_3349,N_3843);
nand U4134 (N_4134,N_3834,N_3895);
or U4135 (N_4135,N_3602,N_3378);
nand U4136 (N_4136,N_3460,N_3366);
xnor U4137 (N_4137,N_3644,N_3898);
nor U4138 (N_4138,N_3508,N_3940);
or U4139 (N_4139,N_3572,N_3518);
nand U4140 (N_4140,N_3665,N_3746);
xnor U4141 (N_4141,N_3163,N_3753);
or U4142 (N_4142,N_3212,N_3726);
and U4143 (N_4143,N_3052,N_3964);
nor U4144 (N_4144,N_3271,N_3527);
xnor U4145 (N_4145,N_3046,N_3116);
nand U4146 (N_4146,N_3958,N_3601);
xor U4147 (N_4147,N_3510,N_3729);
nor U4148 (N_4148,N_3829,N_3587);
or U4149 (N_4149,N_3206,N_3229);
and U4150 (N_4150,N_3209,N_3945);
and U4151 (N_4151,N_3521,N_3464);
and U4152 (N_4152,N_3471,N_3846);
nor U4153 (N_4153,N_3582,N_3093);
and U4154 (N_4154,N_3592,N_3970);
and U4155 (N_4155,N_3948,N_3694);
xnor U4156 (N_4156,N_3462,N_3005);
nand U4157 (N_4157,N_3420,N_3439);
or U4158 (N_4158,N_3074,N_3792);
nor U4159 (N_4159,N_3549,N_3727);
and U4160 (N_4160,N_3662,N_3886);
xor U4161 (N_4161,N_3930,N_3487);
and U4162 (N_4162,N_3748,N_3685);
nand U4163 (N_4163,N_3516,N_3006);
nor U4164 (N_4164,N_3358,N_3932);
nor U4165 (N_4165,N_3573,N_3075);
or U4166 (N_4166,N_3386,N_3801);
nand U4167 (N_4167,N_3361,N_3326);
xnor U4168 (N_4168,N_3422,N_3058);
and U4169 (N_4169,N_3885,N_3654);
xnor U4170 (N_4170,N_3849,N_3520);
xor U4171 (N_4171,N_3459,N_3794);
xnor U4172 (N_4172,N_3099,N_3797);
and U4173 (N_4173,N_3826,N_3923);
and U4174 (N_4174,N_3109,N_3757);
or U4175 (N_4175,N_3483,N_3079);
nand U4176 (N_4176,N_3373,N_3215);
nor U4177 (N_4177,N_3383,N_3403);
or U4178 (N_4178,N_3999,N_3073);
nand U4179 (N_4179,N_3900,N_3697);
nand U4180 (N_4180,N_3336,N_3389);
nor U4181 (N_4181,N_3452,N_3408);
nand U4182 (N_4182,N_3976,N_3505);
or U4183 (N_4183,N_3344,N_3171);
nand U4184 (N_4184,N_3738,N_3145);
and U4185 (N_4185,N_3670,N_3631);
and U4186 (N_4186,N_3037,N_3993);
nor U4187 (N_4187,N_3780,N_3282);
and U4188 (N_4188,N_3833,N_3522);
nand U4189 (N_4189,N_3310,N_3298);
xor U4190 (N_4190,N_3029,N_3189);
and U4191 (N_4191,N_3104,N_3194);
nand U4192 (N_4192,N_3356,N_3421);
nor U4193 (N_4193,N_3621,N_3946);
nand U4194 (N_4194,N_3463,N_3064);
xor U4195 (N_4195,N_3981,N_3741);
nor U4196 (N_4196,N_3153,N_3667);
nor U4197 (N_4197,N_3936,N_3272);
nor U4198 (N_4198,N_3725,N_3355);
nor U4199 (N_4199,N_3238,N_3054);
or U4200 (N_4200,N_3953,N_3589);
nor U4201 (N_4201,N_3774,N_3224);
xor U4202 (N_4202,N_3817,N_3449);
nor U4203 (N_4203,N_3211,N_3329);
xnor U4204 (N_4204,N_3144,N_3766);
and U4205 (N_4205,N_3918,N_3911);
or U4206 (N_4206,N_3382,N_3570);
nand U4207 (N_4207,N_3394,N_3803);
or U4208 (N_4208,N_3020,N_3884);
xnor U4209 (N_4209,N_3205,N_3245);
nand U4210 (N_4210,N_3261,N_3609);
nor U4211 (N_4211,N_3453,N_3990);
nand U4212 (N_4212,N_3822,N_3450);
nor U4213 (N_4213,N_3473,N_3484);
nor U4214 (N_4214,N_3596,N_3643);
xnor U4215 (N_4215,N_3290,N_3167);
or U4216 (N_4216,N_3392,N_3185);
nand U4217 (N_4217,N_3134,N_3556);
nor U4218 (N_4218,N_3671,N_3824);
nor U4219 (N_4219,N_3839,N_3513);
xnor U4220 (N_4220,N_3901,N_3139);
xor U4221 (N_4221,N_3112,N_3847);
or U4222 (N_4222,N_3416,N_3339);
and U4223 (N_4223,N_3423,N_3065);
nand U4224 (N_4224,N_3313,N_3528);
nand U4225 (N_4225,N_3611,N_3264);
xnor U4226 (N_4226,N_3303,N_3853);
nor U4227 (N_4227,N_3396,N_3155);
xnor U4228 (N_4228,N_3047,N_3761);
and U4229 (N_4229,N_3485,N_3069);
and U4230 (N_4230,N_3297,N_3100);
nor U4231 (N_4231,N_3433,N_3016);
nor U4232 (N_4232,N_3003,N_3184);
nand U4233 (N_4233,N_3499,N_3622);
xor U4234 (N_4234,N_3969,N_3111);
nor U4235 (N_4235,N_3497,N_3831);
and U4236 (N_4236,N_3221,N_3795);
and U4237 (N_4237,N_3995,N_3232);
or U4238 (N_4238,N_3742,N_3961);
xnor U4239 (N_4239,N_3799,N_3860);
xnor U4240 (N_4240,N_3124,N_3374);
or U4241 (N_4241,N_3220,N_3141);
and U4242 (N_4242,N_3034,N_3576);
xor U4243 (N_4243,N_3678,N_3254);
nor U4244 (N_4244,N_3381,N_3955);
or U4245 (N_4245,N_3949,N_3191);
nor U4246 (N_4246,N_3021,N_3022);
nor U4247 (N_4247,N_3150,N_3889);
xor U4248 (N_4248,N_3377,N_3379);
or U4249 (N_4249,N_3087,N_3195);
nor U4250 (N_4250,N_3613,N_3019);
nor U4251 (N_4251,N_3399,N_3616);
nor U4252 (N_4252,N_3226,N_3503);
nor U4253 (N_4253,N_3481,N_3208);
nand U4254 (N_4254,N_3181,N_3444);
nor U4255 (N_4255,N_3523,N_3933);
xnor U4256 (N_4256,N_3156,N_3942);
or U4257 (N_4257,N_3567,N_3919);
xor U4258 (N_4258,N_3431,N_3681);
nand U4259 (N_4259,N_3129,N_3716);
nand U4260 (N_4260,N_3438,N_3820);
and U4261 (N_4261,N_3705,N_3180);
or U4262 (N_4262,N_3871,N_3861);
xor U4263 (N_4263,N_3593,N_3532);
nand U4264 (N_4264,N_3494,N_3302);
or U4265 (N_4265,N_3698,N_3435);
xnor U4266 (N_4266,N_3010,N_3051);
and U4267 (N_4267,N_3203,N_3237);
or U4268 (N_4268,N_3265,N_3387);
nand U4269 (N_4269,N_3661,N_3113);
nand U4270 (N_4270,N_3357,N_3013);
xnor U4271 (N_4271,N_3540,N_3735);
nand U4272 (N_4272,N_3558,N_3659);
xor U4273 (N_4273,N_3063,N_3406);
or U4274 (N_4274,N_3956,N_3926);
or U4275 (N_4275,N_3082,N_3632);
xor U4276 (N_4276,N_3904,N_3784);
and U4277 (N_4277,N_3619,N_3569);
or U4278 (N_4278,N_3563,N_3851);
nand U4279 (N_4279,N_3312,N_3193);
or U4280 (N_4280,N_3910,N_3872);
nand U4281 (N_4281,N_3882,N_3688);
or U4282 (N_4282,N_3606,N_3351);
or U4283 (N_4283,N_3246,N_3318);
nor U4284 (N_4284,N_3327,N_3241);
or U4285 (N_4285,N_3723,N_3917);
and U4286 (N_4286,N_3691,N_3603);
xor U4287 (N_4287,N_3838,N_3899);
nand U4288 (N_4288,N_3863,N_3983);
nor U4289 (N_4289,N_3168,N_3216);
xnor U4290 (N_4290,N_3696,N_3836);
xnor U4291 (N_4291,N_3341,N_3121);
nor U4292 (N_4292,N_3448,N_3966);
nor U4293 (N_4293,N_3110,N_3542);
or U4294 (N_4294,N_3210,N_3640);
and U4295 (N_4295,N_3089,N_3335);
nor U4296 (N_4296,N_3786,N_3166);
nand U4297 (N_4297,N_3894,N_3311);
nor U4298 (N_4298,N_3982,N_3548);
and U4299 (N_4299,N_3325,N_3977);
nand U4300 (N_4300,N_3907,N_3519);
xnor U4301 (N_4301,N_3720,N_3222);
or U4302 (N_4302,N_3055,N_3085);
xnor U4303 (N_4303,N_3077,N_3295);
nand U4304 (N_4304,N_3538,N_3533);
nor U4305 (N_4305,N_3931,N_3040);
or U4306 (N_4306,N_3174,N_3635);
nor U4307 (N_4307,N_3639,N_3348);
and U4308 (N_4308,N_3517,N_3653);
xor U4309 (N_4309,N_3292,N_3258);
nand U4310 (N_4310,N_3467,N_3762);
nor U4311 (N_4311,N_3401,N_3190);
and U4312 (N_4312,N_3002,N_3363);
nand U4313 (N_4313,N_3734,N_3699);
nand U4314 (N_4314,N_3868,N_3700);
nor U4315 (N_4315,N_3750,N_3739);
nor U4316 (N_4316,N_3061,N_3769);
xnor U4317 (N_4317,N_3855,N_3765);
xnor U4318 (N_4318,N_3719,N_3159);
or U4319 (N_4319,N_3284,N_3427);
and U4320 (N_4320,N_3346,N_3943);
or U4321 (N_4321,N_3580,N_3301);
xor U4322 (N_4322,N_3565,N_3380);
and U4323 (N_4323,N_3273,N_3101);
nand U4324 (N_4324,N_3649,N_3535);
xnor U4325 (N_4325,N_3514,N_3914);
or U4326 (N_4326,N_3627,N_3090);
nor U4327 (N_4327,N_3989,N_3620);
xor U4328 (N_4328,N_3086,N_3007);
nor U4329 (N_4329,N_3143,N_3617);
nand U4330 (N_4330,N_3717,N_3028);
or U4331 (N_4331,N_3263,N_3122);
xor U4332 (N_4332,N_3935,N_3706);
or U4333 (N_4333,N_3353,N_3909);
or U4334 (N_4334,N_3937,N_3870);
or U4335 (N_4335,N_3728,N_3011);
nor U4336 (N_4336,N_3092,N_3137);
or U4337 (N_4337,N_3553,N_3239);
or U4338 (N_4338,N_3626,N_3928);
or U4339 (N_4339,N_3722,N_3821);
nand U4340 (N_4340,N_3759,N_3883);
nand U4341 (N_4341,N_3084,N_3905);
or U4342 (N_4342,N_3550,N_3067);
nand U4343 (N_4343,N_3498,N_3160);
xnor U4344 (N_4344,N_3375,N_3350);
or U4345 (N_4345,N_3235,N_3474);
nor U4346 (N_4346,N_3256,N_3546);
nor U4347 (N_4347,N_3492,N_3781);
nand U4348 (N_4348,N_3454,N_3252);
and U4349 (N_4349,N_3529,N_3248);
or U4350 (N_4350,N_3251,N_3775);
nor U4351 (N_4351,N_3618,N_3340);
xnor U4352 (N_4352,N_3126,N_3305);
xor U4353 (N_4353,N_3957,N_3411);
or U4354 (N_4354,N_3950,N_3903);
nand U4355 (N_4355,N_3888,N_3461);
nor U4356 (N_4356,N_3938,N_3285);
nand U4357 (N_4357,N_3133,N_3515);
nor U4358 (N_4358,N_3049,N_3552);
and U4359 (N_4359,N_3468,N_3094);
and U4360 (N_4360,N_3475,N_3231);
nand U4361 (N_4361,N_3128,N_3404);
and U4362 (N_4362,N_3059,N_3288);
nand U4363 (N_4363,N_3877,N_3922);
and U4364 (N_4364,N_3182,N_3489);
and U4365 (N_4365,N_3633,N_3534);
and U4366 (N_4366,N_3342,N_3815);
nand U4367 (N_4367,N_3554,N_3169);
nor U4368 (N_4368,N_3577,N_3026);
nor U4369 (N_4369,N_3045,N_3321);
xor U4370 (N_4370,N_3274,N_3161);
or U4371 (N_4371,N_3501,N_3869);
and U4372 (N_4372,N_3755,N_3844);
xor U4373 (N_4373,N_3758,N_3814);
xnor U4374 (N_4374,N_3234,N_3414);
nor U4375 (N_4375,N_3441,N_3050);
or U4376 (N_4376,N_3429,N_3409);
xnor U4377 (N_4377,N_3690,N_3364);
xor U4378 (N_4378,N_3880,N_3566);
and U4379 (N_4379,N_3939,N_3893);
or U4380 (N_4380,N_3162,N_3867);
or U4381 (N_4381,N_3048,N_3608);
and U4382 (N_4382,N_3703,N_3876);
and U4383 (N_4383,N_3269,N_3693);
nand U4384 (N_4384,N_3971,N_3097);
and U4385 (N_4385,N_3973,N_3979);
nor U4386 (N_4386,N_3524,N_3267);
and U4387 (N_4387,N_3625,N_3680);
nor U4388 (N_4388,N_3333,N_3952);
xnor U4389 (N_4389,N_3733,N_3715);
or U4390 (N_4390,N_3805,N_3165);
nand U4391 (N_4391,N_3027,N_3213);
nor U4392 (N_4392,N_3391,N_3044);
nor U4393 (N_4393,N_3173,N_3249);
xnor U4394 (N_4394,N_3482,N_3651);
and U4395 (N_4395,N_3197,N_3148);
nand U4396 (N_4396,N_3597,N_3107);
and U4397 (N_4397,N_3897,N_3188);
nor U4398 (N_4398,N_3881,N_3009);
xor U4399 (N_4399,N_3686,N_3802);
and U4400 (N_4400,N_3812,N_3852);
xnor U4401 (N_4401,N_3132,N_3920);
or U4402 (N_4402,N_3445,N_3998);
or U4403 (N_4403,N_3227,N_3496);
nand U4404 (N_4404,N_3744,N_3176);
nand U4405 (N_4405,N_3630,N_3547);
nor U4406 (N_4406,N_3747,N_3268);
xnor U4407 (N_4407,N_3062,N_3177);
xnor U4408 (N_4408,N_3309,N_3266);
or U4409 (N_4409,N_3183,N_3186);
or U4410 (N_4410,N_3418,N_3987);
nand U4411 (N_4411,N_3509,N_3772);
and U4412 (N_4412,N_3018,N_3842);
nand U4413 (N_4413,N_3371,N_3223);
xnor U4414 (N_4414,N_3397,N_3892);
nor U4415 (N_4415,N_3607,N_3434);
xor U4416 (N_4416,N_3963,N_3745);
nand U4417 (N_4417,N_3771,N_3446);
nand U4418 (N_4418,N_3105,N_3432);
nor U4419 (N_4419,N_3024,N_3585);
xor U4420 (N_4420,N_3790,N_3343);
or U4421 (N_4421,N_3714,N_3588);
and U4422 (N_4422,N_3436,N_3865);
nor U4423 (N_4423,N_3491,N_3332);
and U4424 (N_4424,N_3835,N_3428);
or U4425 (N_4425,N_3071,N_3207);
xor U4426 (N_4426,N_3413,N_3655);
xor U4427 (N_4427,N_3456,N_3236);
nor U4428 (N_4428,N_3323,N_3260);
nand U4429 (N_4429,N_3330,N_3828);
nand U4430 (N_4430,N_3214,N_3811);
nor U4431 (N_4431,N_3004,N_3859);
nand U4432 (N_4432,N_3793,N_3830);
xnor U4433 (N_4433,N_3147,N_3151);
or U4434 (N_4434,N_3164,N_3954);
xnor U4435 (N_4435,N_3525,N_3359);
nor U4436 (N_4436,N_3944,N_3896);
or U4437 (N_4437,N_3783,N_3557);
nor U4438 (N_4438,N_3673,N_3278);
nand U4439 (N_4439,N_3081,N_3798);
nor U4440 (N_4440,N_3458,N_3848);
or U4441 (N_4441,N_3692,N_3407);
and U4442 (N_4442,N_3975,N_3476);
or U4443 (N_4443,N_3125,N_3338);
nand U4444 (N_4444,N_3985,N_3965);
and U4445 (N_4445,N_3179,N_3477);
and U4446 (N_4446,N_3791,N_3816);
or U4447 (N_4447,N_3192,N_3808);
nor U4448 (N_4448,N_3925,N_3545);
nand U4449 (N_4449,N_3590,N_3737);
and U4450 (N_4450,N_3664,N_3276);
nand U4451 (N_4451,N_3057,N_3676);
or U4452 (N_4452,N_3488,N_3986);
xor U4453 (N_4453,N_3076,N_3927);
and U4454 (N_4454,N_3787,N_3624);
or U4455 (N_4455,N_3604,N_3201);
xnor U4456 (N_4456,N_3994,N_3287);
and U4457 (N_4457,N_3053,N_3228);
nor U4458 (N_4458,N_3866,N_3158);
nor U4459 (N_4459,N_3921,N_3850);
xnor U4460 (N_4460,N_3862,N_3628);
nand U4461 (N_4461,N_3687,N_3102);
nor U4462 (N_4462,N_3291,N_3244);
and U4463 (N_4463,N_3187,N_3767);
or U4464 (N_4464,N_3202,N_3479);
or U4465 (N_4465,N_3253,N_3586);
nand U4466 (N_4466,N_3984,N_3495);
and U4467 (N_4467,N_3106,N_3493);
xnor U4468 (N_4468,N_3140,N_3788);
nand U4469 (N_4469,N_3806,N_3809);
nor U4470 (N_4470,N_3707,N_3612);
nor U4471 (N_4471,N_3304,N_3042);
xnor U4472 (N_4472,N_3857,N_3929);
nor U4473 (N_4473,N_3764,N_3115);
nor U4474 (N_4474,N_3752,N_3114);
or U4475 (N_4475,N_3669,N_3854);
nor U4476 (N_4476,N_3740,N_3032);
nand U4477 (N_4477,N_3080,N_3906);
xnor U4478 (N_4478,N_3091,N_3096);
xnor U4479 (N_4479,N_3962,N_3393);
xnor U4480 (N_4480,N_3623,N_3614);
or U4481 (N_4481,N_3785,N_3537);
and U4482 (N_4482,N_3677,N_3157);
nand U4483 (N_4483,N_3709,N_3472);
or U4484 (N_4484,N_3307,N_3286);
and U4485 (N_4485,N_3634,N_3713);
nor U4486 (N_4486,N_3259,N_3000);
nor U4487 (N_4487,N_3960,N_3430);
nand U4488 (N_4488,N_3652,N_3035);
xor U4489 (N_4489,N_3832,N_3718);
xnor U4490 (N_4490,N_3648,N_3217);
xor U4491 (N_4491,N_3813,N_3913);
and U4492 (N_4492,N_3337,N_3571);
nor U4493 (N_4493,N_3068,N_3988);
and U4494 (N_4494,N_3131,N_3200);
nor U4495 (N_4495,N_3777,N_3564);
nand U4496 (N_4496,N_3879,N_3270);
and U4497 (N_4497,N_3526,N_3941);
and U4498 (N_4498,N_3443,N_3149);
or U4499 (N_4499,N_3331,N_3773);
xor U4500 (N_4500,N_3474,N_3013);
and U4501 (N_4501,N_3730,N_3114);
nor U4502 (N_4502,N_3431,N_3552);
or U4503 (N_4503,N_3849,N_3338);
xnor U4504 (N_4504,N_3194,N_3976);
and U4505 (N_4505,N_3251,N_3107);
nor U4506 (N_4506,N_3732,N_3300);
or U4507 (N_4507,N_3682,N_3070);
or U4508 (N_4508,N_3543,N_3437);
xnor U4509 (N_4509,N_3093,N_3473);
xnor U4510 (N_4510,N_3403,N_3479);
xor U4511 (N_4511,N_3883,N_3477);
nand U4512 (N_4512,N_3886,N_3763);
nor U4513 (N_4513,N_3548,N_3923);
or U4514 (N_4514,N_3837,N_3551);
nand U4515 (N_4515,N_3303,N_3015);
nor U4516 (N_4516,N_3834,N_3415);
or U4517 (N_4517,N_3784,N_3489);
xor U4518 (N_4518,N_3948,N_3699);
or U4519 (N_4519,N_3313,N_3453);
or U4520 (N_4520,N_3772,N_3189);
nor U4521 (N_4521,N_3202,N_3828);
or U4522 (N_4522,N_3175,N_3648);
nand U4523 (N_4523,N_3292,N_3639);
xor U4524 (N_4524,N_3102,N_3314);
nand U4525 (N_4525,N_3771,N_3644);
nor U4526 (N_4526,N_3565,N_3451);
nor U4527 (N_4527,N_3098,N_3148);
nand U4528 (N_4528,N_3172,N_3028);
or U4529 (N_4529,N_3777,N_3420);
nand U4530 (N_4530,N_3697,N_3878);
and U4531 (N_4531,N_3941,N_3927);
or U4532 (N_4532,N_3708,N_3385);
nor U4533 (N_4533,N_3309,N_3464);
nor U4534 (N_4534,N_3756,N_3809);
or U4535 (N_4535,N_3633,N_3504);
nand U4536 (N_4536,N_3429,N_3495);
and U4537 (N_4537,N_3325,N_3027);
xor U4538 (N_4538,N_3095,N_3353);
or U4539 (N_4539,N_3820,N_3735);
and U4540 (N_4540,N_3074,N_3648);
nand U4541 (N_4541,N_3708,N_3197);
or U4542 (N_4542,N_3060,N_3089);
or U4543 (N_4543,N_3290,N_3238);
and U4544 (N_4544,N_3057,N_3472);
and U4545 (N_4545,N_3371,N_3075);
and U4546 (N_4546,N_3367,N_3353);
or U4547 (N_4547,N_3216,N_3121);
and U4548 (N_4548,N_3221,N_3032);
nor U4549 (N_4549,N_3304,N_3176);
nand U4550 (N_4550,N_3636,N_3473);
nand U4551 (N_4551,N_3761,N_3576);
nor U4552 (N_4552,N_3716,N_3492);
and U4553 (N_4553,N_3909,N_3243);
xnor U4554 (N_4554,N_3159,N_3018);
or U4555 (N_4555,N_3535,N_3932);
xor U4556 (N_4556,N_3812,N_3741);
nor U4557 (N_4557,N_3213,N_3754);
nand U4558 (N_4558,N_3720,N_3326);
or U4559 (N_4559,N_3568,N_3188);
or U4560 (N_4560,N_3112,N_3489);
xnor U4561 (N_4561,N_3008,N_3762);
or U4562 (N_4562,N_3912,N_3626);
nand U4563 (N_4563,N_3858,N_3850);
xor U4564 (N_4564,N_3724,N_3654);
xor U4565 (N_4565,N_3652,N_3937);
nand U4566 (N_4566,N_3594,N_3995);
nor U4567 (N_4567,N_3295,N_3852);
nand U4568 (N_4568,N_3993,N_3602);
and U4569 (N_4569,N_3063,N_3066);
nand U4570 (N_4570,N_3274,N_3296);
nand U4571 (N_4571,N_3097,N_3223);
and U4572 (N_4572,N_3314,N_3614);
and U4573 (N_4573,N_3846,N_3822);
nor U4574 (N_4574,N_3756,N_3539);
nand U4575 (N_4575,N_3870,N_3217);
nor U4576 (N_4576,N_3639,N_3214);
xor U4577 (N_4577,N_3765,N_3890);
or U4578 (N_4578,N_3797,N_3049);
and U4579 (N_4579,N_3720,N_3147);
xnor U4580 (N_4580,N_3372,N_3735);
nand U4581 (N_4581,N_3362,N_3635);
or U4582 (N_4582,N_3764,N_3816);
nor U4583 (N_4583,N_3450,N_3612);
xor U4584 (N_4584,N_3366,N_3425);
or U4585 (N_4585,N_3679,N_3047);
nand U4586 (N_4586,N_3433,N_3686);
nand U4587 (N_4587,N_3496,N_3446);
and U4588 (N_4588,N_3669,N_3060);
or U4589 (N_4589,N_3659,N_3890);
and U4590 (N_4590,N_3063,N_3658);
nor U4591 (N_4591,N_3425,N_3385);
xnor U4592 (N_4592,N_3376,N_3068);
xnor U4593 (N_4593,N_3615,N_3204);
and U4594 (N_4594,N_3198,N_3601);
nor U4595 (N_4595,N_3485,N_3221);
nand U4596 (N_4596,N_3071,N_3220);
or U4597 (N_4597,N_3092,N_3106);
nand U4598 (N_4598,N_3030,N_3701);
nand U4599 (N_4599,N_3913,N_3410);
or U4600 (N_4600,N_3768,N_3024);
xnor U4601 (N_4601,N_3520,N_3397);
or U4602 (N_4602,N_3373,N_3542);
nand U4603 (N_4603,N_3272,N_3048);
xor U4604 (N_4604,N_3668,N_3355);
xor U4605 (N_4605,N_3217,N_3434);
or U4606 (N_4606,N_3516,N_3175);
or U4607 (N_4607,N_3811,N_3308);
or U4608 (N_4608,N_3722,N_3311);
or U4609 (N_4609,N_3089,N_3512);
nand U4610 (N_4610,N_3846,N_3190);
and U4611 (N_4611,N_3856,N_3359);
nor U4612 (N_4612,N_3797,N_3422);
nor U4613 (N_4613,N_3576,N_3615);
nor U4614 (N_4614,N_3634,N_3424);
and U4615 (N_4615,N_3212,N_3539);
nor U4616 (N_4616,N_3289,N_3036);
xor U4617 (N_4617,N_3520,N_3372);
or U4618 (N_4618,N_3620,N_3977);
xnor U4619 (N_4619,N_3214,N_3470);
nor U4620 (N_4620,N_3773,N_3291);
or U4621 (N_4621,N_3448,N_3980);
or U4622 (N_4622,N_3843,N_3403);
or U4623 (N_4623,N_3257,N_3862);
xnor U4624 (N_4624,N_3257,N_3936);
or U4625 (N_4625,N_3766,N_3735);
or U4626 (N_4626,N_3120,N_3607);
nor U4627 (N_4627,N_3564,N_3799);
or U4628 (N_4628,N_3687,N_3530);
or U4629 (N_4629,N_3506,N_3385);
xor U4630 (N_4630,N_3266,N_3100);
and U4631 (N_4631,N_3850,N_3420);
and U4632 (N_4632,N_3095,N_3418);
or U4633 (N_4633,N_3328,N_3849);
or U4634 (N_4634,N_3544,N_3134);
nand U4635 (N_4635,N_3092,N_3850);
nor U4636 (N_4636,N_3225,N_3339);
and U4637 (N_4637,N_3832,N_3263);
nand U4638 (N_4638,N_3657,N_3697);
and U4639 (N_4639,N_3314,N_3141);
nor U4640 (N_4640,N_3736,N_3447);
nand U4641 (N_4641,N_3419,N_3226);
or U4642 (N_4642,N_3023,N_3097);
nand U4643 (N_4643,N_3134,N_3607);
or U4644 (N_4644,N_3884,N_3462);
or U4645 (N_4645,N_3088,N_3196);
xor U4646 (N_4646,N_3691,N_3162);
or U4647 (N_4647,N_3139,N_3643);
nor U4648 (N_4648,N_3524,N_3850);
or U4649 (N_4649,N_3815,N_3122);
xnor U4650 (N_4650,N_3941,N_3873);
nand U4651 (N_4651,N_3528,N_3797);
nand U4652 (N_4652,N_3102,N_3535);
xnor U4653 (N_4653,N_3221,N_3261);
nor U4654 (N_4654,N_3460,N_3452);
and U4655 (N_4655,N_3160,N_3410);
and U4656 (N_4656,N_3182,N_3284);
xnor U4657 (N_4657,N_3706,N_3763);
and U4658 (N_4658,N_3359,N_3984);
or U4659 (N_4659,N_3710,N_3602);
nand U4660 (N_4660,N_3724,N_3728);
and U4661 (N_4661,N_3724,N_3850);
nor U4662 (N_4662,N_3954,N_3124);
or U4663 (N_4663,N_3854,N_3501);
and U4664 (N_4664,N_3947,N_3300);
nor U4665 (N_4665,N_3569,N_3589);
and U4666 (N_4666,N_3673,N_3392);
nor U4667 (N_4667,N_3484,N_3039);
and U4668 (N_4668,N_3358,N_3016);
nor U4669 (N_4669,N_3078,N_3814);
nand U4670 (N_4670,N_3060,N_3348);
nand U4671 (N_4671,N_3576,N_3697);
nor U4672 (N_4672,N_3607,N_3405);
nor U4673 (N_4673,N_3659,N_3370);
nand U4674 (N_4674,N_3614,N_3617);
xnor U4675 (N_4675,N_3316,N_3946);
nor U4676 (N_4676,N_3176,N_3900);
and U4677 (N_4677,N_3437,N_3084);
xor U4678 (N_4678,N_3180,N_3528);
xor U4679 (N_4679,N_3433,N_3459);
nand U4680 (N_4680,N_3711,N_3204);
nor U4681 (N_4681,N_3236,N_3664);
and U4682 (N_4682,N_3718,N_3140);
xor U4683 (N_4683,N_3068,N_3003);
xnor U4684 (N_4684,N_3606,N_3294);
xor U4685 (N_4685,N_3615,N_3932);
xnor U4686 (N_4686,N_3310,N_3473);
xor U4687 (N_4687,N_3827,N_3873);
xor U4688 (N_4688,N_3647,N_3696);
nand U4689 (N_4689,N_3632,N_3512);
nand U4690 (N_4690,N_3604,N_3012);
nor U4691 (N_4691,N_3214,N_3821);
nor U4692 (N_4692,N_3654,N_3417);
or U4693 (N_4693,N_3783,N_3433);
nor U4694 (N_4694,N_3094,N_3035);
or U4695 (N_4695,N_3321,N_3998);
and U4696 (N_4696,N_3318,N_3269);
nand U4697 (N_4697,N_3629,N_3584);
nand U4698 (N_4698,N_3381,N_3049);
xor U4699 (N_4699,N_3204,N_3274);
nor U4700 (N_4700,N_3173,N_3215);
nand U4701 (N_4701,N_3509,N_3609);
or U4702 (N_4702,N_3481,N_3091);
or U4703 (N_4703,N_3634,N_3083);
nand U4704 (N_4704,N_3519,N_3554);
and U4705 (N_4705,N_3659,N_3774);
or U4706 (N_4706,N_3630,N_3272);
nand U4707 (N_4707,N_3854,N_3271);
or U4708 (N_4708,N_3388,N_3959);
or U4709 (N_4709,N_3578,N_3164);
nor U4710 (N_4710,N_3897,N_3542);
or U4711 (N_4711,N_3596,N_3264);
nor U4712 (N_4712,N_3205,N_3756);
nor U4713 (N_4713,N_3078,N_3064);
nor U4714 (N_4714,N_3189,N_3961);
xor U4715 (N_4715,N_3812,N_3152);
and U4716 (N_4716,N_3557,N_3700);
nand U4717 (N_4717,N_3409,N_3661);
and U4718 (N_4718,N_3779,N_3986);
nand U4719 (N_4719,N_3735,N_3596);
or U4720 (N_4720,N_3998,N_3533);
nor U4721 (N_4721,N_3260,N_3473);
or U4722 (N_4722,N_3553,N_3693);
nand U4723 (N_4723,N_3914,N_3407);
and U4724 (N_4724,N_3967,N_3976);
nand U4725 (N_4725,N_3589,N_3722);
xnor U4726 (N_4726,N_3384,N_3405);
xnor U4727 (N_4727,N_3203,N_3316);
or U4728 (N_4728,N_3589,N_3815);
nand U4729 (N_4729,N_3521,N_3442);
or U4730 (N_4730,N_3310,N_3521);
xor U4731 (N_4731,N_3428,N_3929);
nand U4732 (N_4732,N_3381,N_3303);
and U4733 (N_4733,N_3711,N_3524);
nand U4734 (N_4734,N_3298,N_3394);
or U4735 (N_4735,N_3665,N_3715);
nor U4736 (N_4736,N_3466,N_3773);
nor U4737 (N_4737,N_3760,N_3883);
nand U4738 (N_4738,N_3189,N_3570);
nor U4739 (N_4739,N_3897,N_3629);
xnor U4740 (N_4740,N_3956,N_3227);
or U4741 (N_4741,N_3114,N_3875);
and U4742 (N_4742,N_3225,N_3455);
or U4743 (N_4743,N_3308,N_3283);
xnor U4744 (N_4744,N_3959,N_3174);
xor U4745 (N_4745,N_3125,N_3724);
nor U4746 (N_4746,N_3514,N_3468);
and U4747 (N_4747,N_3188,N_3333);
xor U4748 (N_4748,N_3772,N_3610);
nor U4749 (N_4749,N_3925,N_3566);
nand U4750 (N_4750,N_3640,N_3540);
xnor U4751 (N_4751,N_3228,N_3426);
nand U4752 (N_4752,N_3742,N_3501);
and U4753 (N_4753,N_3531,N_3759);
xnor U4754 (N_4754,N_3577,N_3864);
or U4755 (N_4755,N_3505,N_3660);
xnor U4756 (N_4756,N_3592,N_3270);
or U4757 (N_4757,N_3281,N_3164);
and U4758 (N_4758,N_3371,N_3655);
nor U4759 (N_4759,N_3931,N_3356);
nor U4760 (N_4760,N_3704,N_3970);
nor U4761 (N_4761,N_3582,N_3726);
or U4762 (N_4762,N_3603,N_3747);
nand U4763 (N_4763,N_3502,N_3035);
nand U4764 (N_4764,N_3554,N_3895);
and U4765 (N_4765,N_3578,N_3248);
nand U4766 (N_4766,N_3054,N_3308);
and U4767 (N_4767,N_3036,N_3247);
and U4768 (N_4768,N_3725,N_3689);
and U4769 (N_4769,N_3429,N_3978);
nor U4770 (N_4770,N_3498,N_3766);
xnor U4771 (N_4771,N_3494,N_3047);
xnor U4772 (N_4772,N_3602,N_3786);
and U4773 (N_4773,N_3208,N_3098);
nor U4774 (N_4774,N_3340,N_3963);
or U4775 (N_4775,N_3706,N_3080);
nor U4776 (N_4776,N_3251,N_3160);
xor U4777 (N_4777,N_3581,N_3171);
and U4778 (N_4778,N_3935,N_3454);
nor U4779 (N_4779,N_3216,N_3329);
xnor U4780 (N_4780,N_3982,N_3960);
xor U4781 (N_4781,N_3595,N_3697);
xor U4782 (N_4782,N_3187,N_3255);
nand U4783 (N_4783,N_3571,N_3818);
nand U4784 (N_4784,N_3350,N_3392);
or U4785 (N_4785,N_3646,N_3449);
nor U4786 (N_4786,N_3571,N_3483);
nand U4787 (N_4787,N_3710,N_3637);
nor U4788 (N_4788,N_3866,N_3562);
nor U4789 (N_4789,N_3881,N_3242);
nor U4790 (N_4790,N_3004,N_3513);
or U4791 (N_4791,N_3639,N_3069);
or U4792 (N_4792,N_3420,N_3330);
nor U4793 (N_4793,N_3898,N_3936);
xnor U4794 (N_4794,N_3846,N_3354);
or U4795 (N_4795,N_3454,N_3390);
nand U4796 (N_4796,N_3786,N_3261);
nand U4797 (N_4797,N_3231,N_3055);
and U4798 (N_4798,N_3753,N_3113);
nor U4799 (N_4799,N_3646,N_3485);
xnor U4800 (N_4800,N_3002,N_3966);
nor U4801 (N_4801,N_3102,N_3959);
xor U4802 (N_4802,N_3740,N_3985);
xor U4803 (N_4803,N_3338,N_3304);
and U4804 (N_4804,N_3184,N_3990);
nand U4805 (N_4805,N_3954,N_3190);
nor U4806 (N_4806,N_3445,N_3989);
xnor U4807 (N_4807,N_3100,N_3184);
or U4808 (N_4808,N_3938,N_3228);
or U4809 (N_4809,N_3170,N_3884);
nand U4810 (N_4810,N_3531,N_3737);
nor U4811 (N_4811,N_3002,N_3258);
nor U4812 (N_4812,N_3806,N_3917);
or U4813 (N_4813,N_3819,N_3874);
nor U4814 (N_4814,N_3290,N_3705);
xnor U4815 (N_4815,N_3621,N_3925);
or U4816 (N_4816,N_3080,N_3256);
nand U4817 (N_4817,N_3363,N_3195);
and U4818 (N_4818,N_3975,N_3376);
or U4819 (N_4819,N_3558,N_3206);
nand U4820 (N_4820,N_3507,N_3586);
and U4821 (N_4821,N_3383,N_3926);
nand U4822 (N_4822,N_3209,N_3976);
nand U4823 (N_4823,N_3671,N_3040);
and U4824 (N_4824,N_3427,N_3907);
xor U4825 (N_4825,N_3959,N_3877);
and U4826 (N_4826,N_3009,N_3185);
nand U4827 (N_4827,N_3586,N_3653);
or U4828 (N_4828,N_3424,N_3878);
and U4829 (N_4829,N_3905,N_3634);
nor U4830 (N_4830,N_3880,N_3003);
or U4831 (N_4831,N_3004,N_3926);
and U4832 (N_4832,N_3907,N_3141);
nand U4833 (N_4833,N_3624,N_3454);
nor U4834 (N_4834,N_3817,N_3058);
xor U4835 (N_4835,N_3837,N_3460);
and U4836 (N_4836,N_3704,N_3056);
nand U4837 (N_4837,N_3810,N_3897);
nand U4838 (N_4838,N_3759,N_3673);
or U4839 (N_4839,N_3485,N_3487);
or U4840 (N_4840,N_3302,N_3525);
or U4841 (N_4841,N_3735,N_3737);
nand U4842 (N_4842,N_3719,N_3032);
xor U4843 (N_4843,N_3503,N_3293);
nor U4844 (N_4844,N_3191,N_3567);
nand U4845 (N_4845,N_3187,N_3059);
nor U4846 (N_4846,N_3945,N_3358);
and U4847 (N_4847,N_3200,N_3097);
nand U4848 (N_4848,N_3156,N_3997);
and U4849 (N_4849,N_3350,N_3135);
and U4850 (N_4850,N_3534,N_3138);
nor U4851 (N_4851,N_3202,N_3079);
nand U4852 (N_4852,N_3030,N_3592);
and U4853 (N_4853,N_3980,N_3551);
nor U4854 (N_4854,N_3657,N_3747);
or U4855 (N_4855,N_3317,N_3999);
nor U4856 (N_4856,N_3115,N_3350);
nor U4857 (N_4857,N_3236,N_3800);
nand U4858 (N_4858,N_3166,N_3080);
or U4859 (N_4859,N_3701,N_3075);
nand U4860 (N_4860,N_3333,N_3244);
nor U4861 (N_4861,N_3125,N_3069);
nor U4862 (N_4862,N_3153,N_3683);
nor U4863 (N_4863,N_3737,N_3843);
nand U4864 (N_4864,N_3728,N_3615);
nand U4865 (N_4865,N_3951,N_3646);
nand U4866 (N_4866,N_3522,N_3965);
nand U4867 (N_4867,N_3544,N_3627);
nor U4868 (N_4868,N_3788,N_3488);
xor U4869 (N_4869,N_3433,N_3498);
or U4870 (N_4870,N_3550,N_3408);
or U4871 (N_4871,N_3315,N_3377);
nand U4872 (N_4872,N_3674,N_3020);
nor U4873 (N_4873,N_3741,N_3226);
xnor U4874 (N_4874,N_3535,N_3018);
and U4875 (N_4875,N_3925,N_3175);
nor U4876 (N_4876,N_3265,N_3280);
or U4877 (N_4877,N_3176,N_3460);
xnor U4878 (N_4878,N_3125,N_3486);
nand U4879 (N_4879,N_3569,N_3065);
and U4880 (N_4880,N_3941,N_3100);
or U4881 (N_4881,N_3036,N_3761);
xnor U4882 (N_4882,N_3506,N_3029);
nor U4883 (N_4883,N_3699,N_3968);
or U4884 (N_4884,N_3499,N_3060);
nand U4885 (N_4885,N_3229,N_3666);
xnor U4886 (N_4886,N_3092,N_3410);
nor U4887 (N_4887,N_3611,N_3968);
xor U4888 (N_4888,N_3681,N_3992);
nand U4889 (N_4889,N_3049,N_3252);
nor U4890 (N_4890,N_3178,N_3839);
xnor U4891 (N_4891,N_3433,N_3113);
nor U4892 (N_4892,N_3519,N_3895);
nor U4893 (N_4893,N_3090,N_3833);
xor U4894 (N_4894,N_3786,N_3507);
nand U4895 (N_4895,N_3285,N_3217);
or U4896 (N_4896,N_3848,N_3411);
or U4897 (N_4897,N_3184,N_3787);
xnor U4898 (N_4898,N_3243,N_3170);
nor U4899 (N_4899,N_3268,N_3399);
xor U4900 (N_4900,N_3160,N_3043);
xnor U4901 (N_4901,N_3478,N_3043);
nor U4902 (N_4902,N_3706,N_3425);
nand U4903 (N_4903,N_3193,N_3109);
or U4904 (N_4904,N_3628,N_3708);
and U4905 (N_4905,N_3726,N_3732);
nor U4906 (N_4906,N_3900,N_3781);
and U4907 (N_4907,N_3771,N_3611);
or U4908 (N_4908,N_3388,N_3975);
or U4909 (N_4909,N_3313,N_3251);
nor U4910 (N_4910,N_3111,N_3678);
xnor U4911 (N_4911,N_3732,N_3534);
nor U4912 (N_4912,N_3558,N_3331);
nor U4913 (N_4913,N_3486,N_3153);
nor U4914 (N_4914,N_3014,N_3720);
and U4915 (N_4915,N_3787,N_3366);
xor U4916 (N_4916,N_3325,N_3351);
nor U4917 (N_4917,N_3234,N_3070);
xnor U4918 (N_4918,N_3392,N_3708);
or U4919 (N_4919,N_3297,N_3503);
xor U4920 (N_4920,N_3705,N_3889);
nor U4921 (N_4921,N_3812,N_3209);
xnor U4922 (N_4922,N_3081,N_3777);
nor U4923 (N_4923,N_3399,N_3561);
nor U4924 (N_4924,N_3709,N_3199);
nor U4925 (N_4925,N_3462,N_3092);
xor U4926 (N_4926,N_3849,N_3766);
nor U4927 (N_4927,N_3440,N_3679);
nand U4928 (N_4928,N_3146,N_3407);
nor U4929 (N_4929,N_3798,N_3015);
or U4930 (N_4930,N_3936,N_3414);
and U4931 (N_4931,N_3921,N_3021);
and U4932 (N_4932,N_3811,N_3934);
nand U4933 (N_4933,N_3444,N_3029);
nand U4934 (N_4934,N_3002,N_3105);
xor U4935 (N_4935,N_3286,N_3963);
nor U4936 (N_4936,N_3442,N_3092);
nor U4937 (N_4937,N_3563,N_3313);
nand U4938 (N_4938,N_3325,N_3734);
nor U4939 (N_4939,N_3528,N_3711);
xnor U4940 (N_4940,N_3624,N_3913);
nor U4941 (N_4941,N_3412,N_3218);
nor U4942 (N_4942,N_3668,N_3885);
nor U4943 (N_4943,N_3690,N_3060);
nand U4944 (N_4944,N_3725,N_3041);
xor U4945 (N_4945,N_3344,N_3177);
nor U4946 (N_4946,N_3066,N_3147);
or U4947 (N_4947,N_3628,N_3726);
and U4948 (N_4948,N_3521,N_3549);
nor U4949 (N_4949,N_3639,N_3434);
nand U4950 (N_4950,N_3268,N_3956);
or U4951 (N_4951,N_3599,N_3634);
xor U4952 (N_4952,N_3302,N_3401);
nand U4953 (N_4953,N_3424,N_3382);
nand U4954 (N_4954,N_3402,N_3008);
and U4955 (N_4955,N_3929,N_3800);
or U4956 (N_4956,N_3747,N_3881);
and U4957 (N_4957,N_3834,N_3491);
nand U4958 (N_4958,N_3172,N_3440);
xnor U4959 (N_4959,N_3238,N_3053);
nand U4960 (N_4960,N_3704,N_3938);
nand U4961 (N_4961,N_3073,N_3000);
nor U4962 (N_4962,N_3154,N_3310);
or U4963 (N_4963,N_3940,N_3781);
xnor U4964 (N_4964,N_3711,N_3612);
nand U4965 (N_4965,N_3296,N_3129);
and U4966 (N_4966,N_3800,N_3612);
or U4967 (N_4967,N_3406,N_3433);
or U4968 (N_4968,N_3812,N_3285);
and U4969 (N_4969,N_3484,N_3361);
xnor U4970 (N_4970,N_3871,N_3991);
nor U4971 (N_4971,N_3525,N_3380);
nand U4972 (N_4972,N_3724,N_3273);
xnor U4973 (N_4973,N_3171,N_3087);
or U4974 (N_4974,N_3808,N_3958);
nor U4975 (N_4975,N_3924,N_3916);
xor U4976 (N_4976,N_3677,N_3351);
nand U4977 (N_4977,N_3495,N_3882);
xnor U4978 (N_4978,N_3851,N_3825);
xor U4979 (N_4979,N_3958,N_3821);
and U4980 (N_4980,N_3454,N_3580);
and U4981 (N_4981,N_3338,N_3896);
nor U4982 (N_4982,N_3778,N_3229);
nand U4983 (N_4983,N_3431,N_3466);
xor U4984 (N_4984,N_3830,N_3297);
xnor U4985 (N_4985,N_3693,N_3979);
nand U4986 (N_4986,N_3969,N_3283);
xor U4987 (N_4987,N_3765,N_3638);
xnor U4988 (N_4988,N_3899,N_3577);
xnor U4989 (N_4989,N_3450,N_3909);
or U4990 (N_4990,N_3068,N_3269);
and U4991 (N_4991,N_3833,N_3656);
nand U4992 (N_4992,N_3647,N_3770);
xnor U4993 (N_4993,N_3391,N_3735);
xnor U4994 (N_4994,N_3277,N_3331);
nand U4995 (N_4995,N_3267,N_3106);
or U4996 (N_4996,N_3492,N_3902);
or U4997 (N_4997,N_3968,N_3785);
or U4998 (N_4998,N_3350,N_3209);
and U4999 (N_4999,N_3329,N_3548);
xnor UO_0 (O_0,N_4996,N_4653);
or UO_1 (O_1,N_4117,N_4939);
nor UO_2 (O_2,N_4380,N_4932);
xor UO_3 (O_3,N_4554,N_4128);
nor UO_4 (O_4,N_4130,N_4086);
nor UO_5 (O_5,N_4234,N_4146);
xnor UO_6 (O_6,N_4351,N_4539);
or UO_7 (O_7,N_4375,N_4541);
and UO_8 (O_8,N_4288,N_4749);
and UO_9 (O_9,N_4543,N_4807);
and UO_10 (O_10,N_4024,N_4880);
nand UO_11 (O_11,N_4339,N_4691);
or UO_12 (O_12,N_4497,N_4673);
and UO_13 (O_13,N_4726,N_4233);
nand UO_14 (O_14,N_4356,N_4484);
nand UO_15 (O_15,N_4781,N_4569);
or UO_16 (O_16,N_4040,N_4796);
xnor UO_17 (O_17,N_4737,N_4424);
nand UO_18 (O_18,N_4202,N_4685);
nor UO_19 (O_19,N_4382,N_4631);
xor UO_20 (O_20,N_4455,N_4283);
nor UO_21 (O_21,N_4946,N_4046);
nor UO_22 (O_22,N_4217,N_4099);
nand UO_23 (O_23,N_4537,N_4406);
nand UO_24 (O_24,N_4296,N_4558);
nand UO_25 (O_25,N_4640,N_4094);
xnor UO_26 (O_26,N_4269,N_4582);
xor UO_27 (O_27,N_4889,N_4710);
and UO_28 (O_28,N_4785,N_4010);
nand UO_29 (O_29,N_4170,N_4335);
nor UO_30 (O_30,N_4384,N_4836);
xor UO_31 (O_31,N_4022,N_4858);
and UO_32 (O_32,N_4227,N_4731);
nor UO_33 (O_33,N_4910,N_4120);
nor UO_34 (O_34,N_4614,N_4125);
nor UO_35 (O_35,N_4316,N_4936);
nand UO_36 (O_36,N_4465,N_4913);
or UO_37 (O_37,N_4183,N_4089);
nand UO_38 (O_38,N_4386,N_4722);
or UO_39 (O_39,N_4463,N_4839);
nand UO_40 (O_40,N_4238,N_4468);
or UO_41 (O_41,N_4795,N_4724);
nand UO_42 (O_42,N_4633,N_4563);
or UO_43 (O_43,N_4439,N_4719);
or UO_44 (O_44,N_4123,N_4925);
xor UO_45 (O_45,N_4573,N_4766);
and UO_46 (O_46,N_4167,N_4560);
or UO_47 (O_47,N_4216,N_4490);
nand UO_48 (O_48,N_4866,N_4716);
nor UO_49 (O_49,N_4743,N_4141);
and UO_50 (O_50,N_4136,N_4599);
and UO_51 (O_51,N_4021,N_4548);
nor UO_52 (O_52,N_4254,N_4707);
and UO_53 (O_53,N_4776,N_4505);
nor UO_54 (O_54,N_4262,N_4818);
or UO_55 (O_55,N_4597,N_4054);
nand UO_56 (O_56,N_4688,N_4196);
nand UO_57 (O_57,N_4295,N_4650);
and UO_58 (O_58,N_4039,N_4188);
xor UO_59 (O_59,N_4590,N_4281);
xor UO_60 (O_60,N_4088,N_4938);
or UO_61 (O_61,N_4323,N_4066);
nand UO_62 (O_62,N_4534,N_4634);
or UO_63 (O_63,N_4052,N_4213);
nor UO_64 (O_64,N_4594,N_4903);
or UO_65 (O_65,N_4044,N_4844);
or UO_66 (O_66,N_4638,N_4608);
and UO_67 (O_67,N_4003,N_4008);
and UO_68 (O_68,N_4538,N_4133);
nor UO_69 (O_69,N_4437,N_4280);
and UO_70 (O_70,N_4469,N_4076);
xnor UO_71 (O_71,N_4603,N_4043);
nand UO_72 (O_72,N_4364,N_4636);
and UO_73 (O_73,N_4292,N_4585);
nand UO_74 (O_74,N_4943,N_4026);
and UO_75 (O_75,N_4096,N_4810);
and UO_76 (O_76,N_4751,N_4359);
nand UO_77 (O_77,N_4253,N_4293);
or UO_78 (O_78,N_4207,N_4070);
xor UO_79 (O_79,N_4260,N_4532);
nor UO_80 (O_80,N_4201,N_4881);
or UO_81 (O_81,N_4799,N_4429);
or UO_82 (O_82,N_4273,N_4310);
and UO_83 (O_83,N_4276,N_4075);
or UO_84 (O_84,N_4690,N_4647);
xor UO_85 (O_85,N_4454,N_4362);
xnor UO_86 (O_86,N_4224,N_4471);
nand UO_87 (O_87,N_4615,N_4734);
and UO_88 (O_88,N_4456,N_4015);
and UO_89 (O_89,N_4999,N_4990);
xor UO_90 (O_90,N_4474,N_4873);
xnor UO_91 (O_91,N_4870,N_4042);
xnor UO_92 (O_92,N_4676,N_4431);
nand UO_93 (O_93,N_4047,N_4643);
nor UO_94 (O_94,N_4971,N_4361);
xor UO_95 (O_95,N_4250,N_4980);
nand UO_96 (O_96,N_4624,N_4137);
and UO_97 (O_97,N_4703,N_4579);
nor UO_98 (O_98,N_4111,N_4122);
nor UO_99 (O_99,N_4846,N_4535);
xnor UO_100 (O_100,N_4907,N_4383);
nand UO_101 (O_101,N_4480,N_4800);
and UO_102 (O_102,N_4435,N_4164);
xor UO_103 (O_103,N_4399,N_4682);
xnor UO_104 (O_104,N_4758,N_4906);
nor UO_105 (O_105,N_4859,N_4034);
or UO_106 (O_106,N_4869,N_4901);
xnor UO_107 (O_107,N_4536,N_4268);
and UO_108 (O_108,N_4817,N_4320);
or UO_109 (O_109,N_4526,N_4433);
or UO_110 (O_110,N_4392,N_4552);
and UO_111 (O_111,N_4885,N_4746);
xnor UO_112 (O_112,N_4082,N_4181);
nor UO_113 (O_113,N_4438,N_4065);
nand UO_114 (O_114,N_4923,N_4395);
nand UO_115 (O_115,N_4815,N_4307);
or UO_116 (O_116,N_4491,N_4699);
or UO_117 (O_117,N_4246,N_4951);
nor UO_118 (O_118,N_4408,N_4162);
and UO_119 (O_119,N_4728,N_4374);
or UO_120 (O_120,N_4430,N_4212);
nor UO_121 (O_121,N_4589,N_4805);
nor UO_122 (O_122,N_4460,N_4328);
nor UO_123 (O_123,N_4860,N_4466);
nand UO_124 (O_124,N_4753,N_4847);
or UO_125 (O_125,N_4459,N_4500);
and UO_126 (O_126,N_4530,N_4888);
nand UO_127 (O_127,N_4998,N_4166);
or UO_128 (O_128,N_4477,N_4571);
nor UO_129 (O_129,N_4108,N_4826);
xor UO_130 (O_130,N_4326,N_4440);
and UO_131 (O_131,N_4112,N_4325);
or UO_132 (O_132,N_4527,N_4191);
nor UO_133 (O_133,N_4791,N_4632);
nor UO_134 (O_134,N_4405,N_4182);
or UO_135 (O_135,N_4786,N_4747);
or UO_136 (O_136,N_4899,N_4777);
and UO_137 (O_137,N_4033,N_4169);
nor UO_138 (O_138,N_4531,N_4772);
nor UO_139 (O_139,N_4160,N_4100);
or UO_140 (O_140,N_4489,N_4308);
and UO_141 (O_141,N_4414,N_4451);
or UO_142 (O_142,N_4354,N_4995);
nand UO_143 (O_143,N_4327,N_4171);
nand UO_144 (O_144,N_4921,N_4740);
or UO_145 (O_145,N_4586,N_4522);
nor UO_146 (O_146,N_4069,N_4237);
and UO_147 (O_147,N_4315,N_4656);
nor UO_148 (O_148,N_4891,N_4139);
xor UO_149 (O_149,N_4265,N_4988);
nand UO_150 (O_150,N_4483,N_4997);
and UO_151 (O_151,N_4666,N_4841);
nand UO_152 (O_152,N_4612,N_4765);
nor UO_153 (O_153,N_4116,N_4816);
xor UO_154 (O_154,N_4360,N_4507);
and UO_155 (O_155,N_4173,N_4159);
or UO_156 (O_156,N_4161,N_4398);
nand UO_157 (O_157,N_4769,N_4119);
xor UO_158 (O_158,N_4780,N_4447);
xnor UO_159 (O_159,N_4371,N_4984);
and UO_160 (O_160,N_4723,N_4613);
nand UO_161 (O_161,N_4969,N_4849);
and UO_162 (O_162,N_4397,N_4197);
nor UO_163 (O_163,N_4966,N_4959);
nand UO_164 (O_164,N_4324,N_4245);
and UO_165 (O_165,N_4620,N_4598);
nand UO_166 (O_166,N_4363,N_4550);
or UO_167 (O_167,N_4078,N_4672);
xnor UO_168 (O_168,N_4801,N_4508);
nand UO_169 (O_169,N_4627,N_4485);
nor UO_170 (O_170,N_4622,N_4302);
and UO_171 (O_171,N_4516,N_4900);
or UO_172 (O_172,N_4091,N_4732);
nor UO_173 (O_173,N_4670,N_4001);
and UO_174 (O_174,N_4274,N_4898);
xor UO_175 (O_175,N_4194,N_4220);
and UO_176 (O_176,N_4605,N_4085);
xor UO_177 (O_177,N_4645,N_4566);
xnor UO_178 (O_178,N_4270,N_4714);
or UO_179 (O_179,N_4006,N_4114);
nand UO_180 (O_180,N_4572,N_4868);
and UO_181 (O_181,N_4072,N_4309);
nor UO_182 (O_182,N_4426,N_4228);
nor UO_183 (O_183,N_4317,N_4652);
nand UO_184 (O_184,N_4291,N_4659);
or UO_185 (O_185,N_4894,N_4215);
xnor UO_186 (O_186,N_4129,N_4808);
xor UO_187 (O_187,N_4488,N_4045);
or UO_188 (O_188,N_4333,N_4427);
nand UO_189 (O_189,N_4979,N_4496);
or UO_190 (O_190,N_4559,N_4068);
nand UO_191 (O_191,N_4294,N_4940);
xnor UO_192 (O_192,N_4448,N_4442);
nor UO_193 (O_193,N_4287,N_4994);
nor UO_194 (O_194,N_4093,N_4762);
nand UO_195 (O_195,N_4745,N_4754);
and UO_196 (O_196,N_4919,N_4748);
and UO_197 (O_197,N_4176,N_4140);
nor UO_198 (O_198,N_4711,N_4057);
nand UO_199 (O_199,N_4761,N_4696);
nor UO_200 (O_200,N_4893,N_4546);
or UO_201 (O_201,N_4446,N_4823);
nand UO_202 (O_202,N_4229,N_4417);
or UO_203 (O_203,N_4098,N_4105);
xnor UO_204 (O_204,N_4214,N_4118);
and UO_205 (O_205,N_4882,N_4681);
xnor UO_206 (O_206,N_4461,N_4963);
xnor UO_207 (O_207,N_4148,N_4739);
and UO_208 (O_208,N_4662,N_4501);
xor UO_209 (O_209,N_4368,N_4942);
and UO_210 (O_210,N_4574,N_4520);
and UO_211 (O_211,N_4916,N_4974);
and UO_212 (O_212,N_4038,N_4187);
and UO_213 (O_213,N_4400,N_4486);
and UO_214 (O_214,N_4156,N_4286);
or UO_215 (O_215,N_4350,N_4012);
nor UO_216 (O_216,N_4718,N_4694);
nor UO_217 (O_217,N_4577,N_4390);
xor UO_218 (O_218,N_4947,N_4177);
nor UO_219 (O_219,N_4352,N_4131);
xnor UO_220 (O_220,N_4080,N_4478);
and UO_221 (O_221,N_4056,N_4679);
xnor UO_222 (O_222,N_4510,N_4581);
nand UO_223 (O_223,N_4935,N_4023);
and UO_224 (O_224,N_4492,N_4266);
and UO_225 (O_225,N_4109,N_4025);
nand UO_226 (O_226,N_4272,N_4264);
and UO_227 (O_227,N_4370,N_4886);
xnor UO_228 (O_228,N_4157,N_4124);
or UO_229 (O_229,N_4300,N_4824);
xor UO_230 (O_230,N_4048,N_4693);
nor UO_231 (O_231,N_4991,N_4175);
and UO_232 (O_232,N_4784,N_4110);
xnor UO_233 (O_233,N_4180,N_4837);
nor UO_234 (O_234,N_4879,N_4902);
nor UO_235 (O_235,N_4037,N_4230);
xnor UO_236 (O_236,N_4713,N_4404);
nand UO_237 (O_237,N_4441,N_4609);
nand UO_238 (O_238,N_4499,N_4113);
xor UO_239 (O_239,N_4231,N_4412);
or UO_240 (O_240,N_4578,N_4204);
nand UO_241 (O_241,N_4792,N_4002);
or UO_242 (O_242,N_4704,N_4811);
nor UO_243 (O_243,N_4321,N_4163);
and UO_244 (O_244,N_4625,N_4556);
or UO_245 (O_245,N_4016,N_4472);
xnor UO_246 (O_246,N_4289,N_4700);
nor UO_247 (O_247,N_4411,N_4387);
or UO_248 (O_248,N_4402,N_4329);
xnor UO_249 (O_249,N_4961,N_4768);
or UO_250 (O_250,N_4821,N_4575);
or UO_251 (O_251,N_4298,N_4542);
nor UO_252 (O_252,N_4927,N_4871);
nand UO_253 (O_253,N_4493,N_4420);
nand UO_254 (O_254,N_4349,N_4968);
or UO_255 (O_255,N_4583,N_4611);
xor UO_256 (O_256,N_4106,N_4121);
and UO_257 (O_257,N_4305,N_4004);
nor UO_258 (O_258,N_4528,N_4000);
nor UO_259 (O_259,N_4263,N_4580);
xnor UO_260 (O_260,N_4628,N_4596);
and UO_261 (O_261,N_4330,N_4917);
xnor UO_262 (O_262,N_4861,N_4067);
nor UO_263 (O_263,N_4962,N_4557);
xor UO_264 (O_264,N_4674,N_4487);
and UO_265 (O_265,N_4436,N_4401);
nor UO_266 (O_266,N_4422,N_4789);
nand UO_267 (O_267,N_4804,N_4648);
xor UO_268 (O_268,N_4388,N_4244);
xnor UO_269 (O_269,N_4020,N_4095);
nand UO_270 (O_270,N_4208,N_4771);
xnor UO_271 (O_271,N_4032,N_4081);
or UO_272 (O_272,N_4313,N_4322);
nor UO_273 (O_273,N_4107,N_4820);
nor UO_274 (O_274,N_4144,N_4084);
xor UO_275 (O_275,N_4481,N_4705);
nor UO_276 (O_276,N_4922,N_4147);
nand UO_277 (O_277,N_4240,N_4948);
and UO_278 (O_278,N_4014,N_4783);
nor UO_279 (O_279,N_4418,N_4249);
and UO_280 (O_280,N_4958,N_4186);
and UO_281 (O_281,N_4934,N_4914);
xor UO_282 (O_282,N_4190,N_4825);
or UO_283 (O_283,N_4983,N_4145);
nor UO_284 (O_284,N_4874,N_4941);
or UO_285 (O_285,N_4883,N_4878);
or UO_286 (O_286,N_4256,N_4547);
xnor UO_287 (O_287,N_4926,N_4251);
nor UO_288 (O_288,N_4760,N_4062);
nor UO_289 (O_289,N_4284,N_4555);
nor UO_290 (O_290,N_4945,N_4778);
xor UO_291 (O_291,N_4956,N_4282);
nor UO_292 (O_292,N_4449,N_4138);
xnor UO_293 (O_293,N_4275,N_4153);
nand UO_294 (O_294,N_4982,N_4950);
or UO_295 (O_295,N_4908,N_4890);
and UO_296 (O_296,N_4415,N_4050);
and UO_297 (O_297,N_4104,N_4079);
nor UO_298 (O_298,N_4813,N_4987);
or UO_299 (O_299,N_4909,N_4005);
xnor UO_300 (O_300,N_4267,N_4606);
or UO_301 (O_301,N_4450,N_4053);
nor UO_302 (O_302,N_4425,N_4862);
xnor UO_303 (O_303,N_4524,N_4657);
and UO_304 (O_304,N_4416,N_4318);
nor UO_305 (O_305,N_4521,N_4011);
and UO_306 (O_306,N_4049,N_4239);
or UO_307 (O_307,N_4338,N_4848);
nand UO_308 (O_308,N_4730,N_4346);
xor UO_309 (O_309,N_4976,N_4756);
xor UO_310 (O_310,N_4797,N_4017);
nand UO_311 (O_311,N_4055,N_4061);
xnor UO_312 (O_312,N_4013,N_4028);
xor UO_313 (O_313,N_4561,N_4036);
and UO_314 (O_314,N_4090,N_4219);
and UO_315 (O_315,N_4671,N_4952);
xnor UO_316 (O_316,N_4252,N_4115);
and UO_317 (O_317,N_4604,N_4413);
and UO_318 (O_318,N_4993,N_4464);
xnor UO_319 (O_319,N_4519,N_4132);
and UO_320 (O_320,N_4986,N_4931);
and UO_321 (O_321,N_4509,N_4863);
and UO_322 (O_322,N_4788,N_4225);
and UO_323 (O_323,N_4030,N_4630);
or UO_324 (O_324,N_4185,N_4518);
xor UO_325 (O_325,N_4831,N_4576);
and UO_326 (O_326,N_4829,N_4729);
or UO_327 (O_327,N_4083,N_4835);
nand UO_328 (O_328,N_4767,N_4378);
or UO_329 (O_329,N_4301,N_4782);
nand UO_330 (O_330,N_4646,N_4060);
and UO_331 (O_331,N_4334,N_4851);
nor UO_332 (O_332,N_4553,N_4709);
xnor UO_333 (O_333,N_4635,N_4506);
xor UO_334 (O_334,N_4134,N_4358);
and UO_335 (O_335,N_4258,N_4641);
and UO_336 (O_336,N_4297,N_4348);
and UO_337 (O_337,N_4517,N_4904);
and UO_338 (O_338,N_4852,N_4843);
nor UO_339 (O_339,N_4341,N_4453);
or UO_340 (O_340,N_4494,N_4445);
or UO_341 (O_341,N_4798,N_4515);
xnor UO_342 (O_342,N_4198,N_4353);
xnor UO_343 (O_343,N_4314,N_4680);
xnor UO_344 (O_344,N_4222,N_4706);
xnor UO_345 (O_345,N_4475,N_4975);
nor UO_346 (O_346,N_4376,N_4235);
nand UO_347 (O_347,N_4365,N_4850);
xor UO_348 (O_348,N_4617,N_4944);
xor UO_349 (O_349,N_4311,N_4261);
xor UO_350 (O_350,N_4051,N_4304);
nor UO_351 (O_351,N_4074,N_4814);
and UO_352 (O_352,N_4992,N_4467);
nand UO_353 (O_353,N_4503,N_4396);
and UO_354 (O_354,N_4545,N_4369);
nor UO_355 (O_355,N_4549,N_4741);
xor UO_356 (O_356,N_4059,N_4241);
nor UO_357 (O_357,N_4142,N_4920);
or UO_358 (O_358,N_4179,N_4720);
xnor UO_359 (O_359,N_4856,N_4794);
nor UO_360 (O_360,N_4695,N_4677);
nand UO_361 (O_361,N_4742,N_4892);
nand UO_362 (O_362,N_4833,N_4564);
xnor UO_363 (O_363,N_4512,N_4271);
nor UO_364 (O_364,N_4853,N_4389);
and UO_365 (O_365,N_4336,N_4462);
nand UO_366 (O_366,N_4964,N_4570);
nor UO_367 (O_367,N_4343,N_4877);
nor UO_368 (O_368,N_4689,N_4102);
nand UO_369 (O_369,N_4827,N_4840);
nand UO_370 (O_370,N_4684,N_4629);
nand UO_371 (O_371,N_4277,N_4683);
nor UO_372 (O_372,N_4668,N_4009);
nand UO_373 (O_373,N_4151,N_4193);
and UO_374 (O_374,N_4533,N_4027);
xor UO_375 (O_375,N_4357,N_4502);
and UO_376 (O_376,N_4593,N_4812);
xor UO_377 (O_377,N_4725,N_4344);
nor UO_378 (O_378,N_4347,N_4058);
or UO_379 (O_379,N_4664,N_4618);
xor UO_380 (O_380,N_4774,N_4540);
xnor UO_381 (O_381,N_4733,N_4372);
nand UO_382 (O_382,N_4409,N_4981);
or UO_383 (O_383,N_4621,N_4092);
xor UO_384 (O_384,N_4912,N_4588);
nand UO_385 (O_385,N_4701,N_4007);
or UO_386 (O_386,N_4514,N_4665);
and UO_387 (O_387,N_4591,N_4595);
nand UO_388 (O_388,N_4930,N_4929);
xor UO_389 (O_389,N_4255,N_4031);
xnor UO_390 (O_390,N_4443,N_4355);
xor UO_391 (O_391,N_4150,N_4623);
or UO_392 (O_392,N_4457,N_4525);
or UO_393 (O_393,N_4290,N_4637);
xor UO_394 (O_394,N_4434,N_4381);
or UO_395 (O_395,N_4154,N_4757);
or UO_396 (O_396,N_4895,N_4452);
nor UO_397 (O_397,N_4565,N_4562);
nand UO_398 (O_398,N_4391,N_4949);
nor UO_399 (O_399,N_4421,N_4965);
nand UO_400 (O_400,N_4223,N_4232);
nand UO_401 (O_401,N_4236,N_4143);
nor UO_402 (O_402,N_4736,N_4189);
and UO_403 (O_403,N_4331,N_4832);
nor UO_404 (O_404,N_4248,N_4977);
nand UO_405 (O_405,N_4367,N_4616);
xnor UO_406 (O_406,N_4667,N_4178);
and UO_407 (O_407,N_4955,N_4041);
and UO_408 (O_408,N_4855,N_4864);
or UO_409 (O_409,N_4649,N_4911);
and UO_410 (O_410,N_4924,N_4639);
and UO_411 (O_411,N_4970,N_4199);
xor UO_412 (O_412,N_4385,N_4126);
nand UO_413 (O_413,N_4819,N_4750);
xor UO_414 (O_414,N_4513,N_4644);
and UO_415 (O_415,N_4752,N_4279);
xor UO_416 (O_416,N_4149,N_4174);
nand UO_417 (O_417,N_4345,N_4601);
xnor UO_418 (O_418,N_4407,N_4332);
and UO_419 (O_419,N_4218,N_4830);
nand UO_420 (O_420,N_4366,N_4155);
xor UO_421 (O_421,N_4087,N_4567);
xnor UO_422 (O_422,N_4838,N_4379);
or UO_423 (O_423,N_4568,N_4319);
xor UO_424 (O_424,N_4872,N_4989);
xor UO_425 (O_425,N_4035,N_4790);
nand UO_426 (O_426,N_4960,N_4764);
nand UO_427 (O_427,N_4168,N_4479);
nand UO_428 (O_428,N_4602,N_4205);
or UO_429 (O_429,N_4192,N_4259);
and UO_430 (O_430,N_4299,N_4592);
nor UO_431 (O_431,N_4802,N_4933);
xor UO_432 (O_432,N_4698,N_4773);
nand UO_433 (O_433,N_4822,N_4744);
nand UO_434 (O_434,N_4654,N_4905);
nand UO_435 (O_435,N_4473,N_4377);
nand UO_436 (O_436,N_4470,N_4019);
and UO_437 (O_437,N_4787,N_4097);
nand UO_438 (O_438,N_4206,N_4854);
or UO_439 (O_439,N_4077,N_4721);
nand UO_440 (O_440,N_4763,N_4103);
or UO_441 (O_441,N_4029,N_4972);
and UO_442 (O_442,N_4793,N_4779);
or UO_443 (O_443,N_4073,N_4626);
nand UO_444 (O_444,N_4727,N_4152);
nand UO_445 (O_445,N_4511,N_4865);
nand UO_446 (O_446,N_4809,N_4896);
xor UO_447 (O_447,N_4071,N_4954);
and UO_448 (O_448,N_4211,N_4697);
nor UO_449 (O_449,N_4101,N_4342);
and UO_450 (O_450,N_4444,N_4803);
and UO_451 (O_451,N_4584,N_4708);
nand UO_452 (O_452,N_4410,N_4675);
nand UO_453 (O_453,N_4498,N_4340);
xor UO_454 (O_454,N_4953,N_4337);
and UO_455 (O_455,N_4610,N_4165);
or UO_456 (O_456,N_4619,N_4875);
nand UO_457 (O_457,N_4278,N_4312);
or UO_458 (O_458,N_4018,N_4247);
and UO_459 (O_459,N_4458,N_4985);
nand UO_460 (O_460,N_4957,N_4928);
nand UO_461 (O_461,N_4967,N_4226);
nand UO_462 (O_462,N_4978,N_4755);
or UO_463 (O_463,N_4482,N_4200);
nand UO_464 (O_464,N_4738,N_4686);
nor UO_465 (O_465,N_4828,N_4423);
nand UO_466 (O_466,N_4887,N_4918);
nand UO_467 (O_467,N_4242,N_4687);
nor UO_468 (O_468,N_4775,N_4373);
xnor UO_469 (O_469,N_4063,N_4973);
nor UO_470 (O_470,N_4857,N_4915);
nand UO_471 (O_471,N_4806,N_4257);
or UO_472 (O_472,N_4495,N_4712);
nand UO_473 (O_473,N_4209,N_4158);
and UO_474 (O_474,N_4658,N_4867);
or UO_475 (O_475,N_4770,N_4393);
or UO_476 (O_476,N_4285,N_4834);
and UO_477 (O_477,N_4661,N_4476);
and UO_478 (O_478,N_4127,N_4306);
nand UO_479 (O_479,N_4243,N_4655);
and UO_480 (O_480,N_4715,N_4669);
or UO_481 (O_481,N_4607,N_4184);
and UO_482 (O_482,N_4735,N_4544);
nor UO_483 (O_483,N_4432,N_4660);
nand UO_484 (O_484,N_4195,N_4303);
nand UO_485 (O_485,N_4884,N_4523);
xor UO_486 (O_486,N_4551,N_4210);
nor UO_487 (O_487,N_4419,N_4394);
and UO_488 (O_488,N_4897,N_4876);
or UO_489 (O_489,N_4651,N_4221);
nor UO_490 (O_490,N_4702,N_4692);
nand UO_491 (O_491,N_4678,N_4428);
xor UO_492 (O_492,N_4203,N_4759);
or UO_493 (O_493,N_4504,N_4403);
xnor UO_494 (O_494,N_4600,N_4842);
nand UO_495 (O_495,N_4172,N_4937);
xor UO_496 (O_496,N_4064,N_4717);
xor UO_497 (O_497,N_4135,N_4845);
nand UO_498 (O_498,N_4663,N_4587);
xnor UO_499 (O_499,N_4642,N_4529);
nand UO_500 (O_500,N_4710,N_4606);
nand UO_501 (O_501,N_4936,N_4938);
or UO_502 (O_502,N_4596,N_4126);
nor UO_503 (O_503,N_4001,N_4929);
or UO_504 (O_504,N_4482,N_4607);
and UO_505 (O_505,N_4797,N_4938);
or UO_506 (O_506,N_4176,N_4524);
and UO_507 (O_507,N_4973,N_4081);
or UO_508 (O_508,N_4614,N_4224);
or UO_509 (O_509,N_4941,N_4824);
nor UO_510 (O_510,N_4936,N_4388);
xor UO_511 (O_511,N_4522,N_4244);
xor UO_512 (O_512,N_4679,N_4364);
nand UO_513 (O_513,N_4594,N_4069);
nor UO_514 (O_514,N_4867,N_4365);
or UO_515 (O_515,N_4034,N_4557);
nand UO_516 (O_516,N_4218,N_4202);
nand UO_517 (O_517,N_4989,N_4189);
nor UO_518 (O_518,N_4316,N_4078);
nand UO_519 (O_519,N_4300,N_4855);
or UO_520 (O_520,N_4288,N_4858);
nand UO_521 (O_521,N_4522,N_4261);
nand UO_522 (O_522,N_4124,N_4095);
nand UO_523 (O_523,N_4852,N_4184);
and UO_524 (O_524,N_4758,N_4582);
xnor UO_525 (O_525,N_4191,N_4939);
nor UO_526 (O_526,N_4138,N_4790);
and UO_527 (O_527,N_4722,N_4357);
and UO_528 (O_528,N_4176,N_4752);
nor UO_529 (O_529,N_4489,N_4179);
or UO_530 (O_530,N_4019,N_4650);
xor UO_531 (O_531,N_4881,N_4195);
or UO_532 (O_532,N_4498,N_4877);
xnor UO_533 (O_533,N_4072,N_4975);
xor UO_534 (O_534,N_4868,N_4238);
nand UO_535 (O_535,N_4701,N_4081);
nand UO_536 (O_536,N_4241,N_4123);
xnor UO_537 (O_537,N_4861,N_4730);
xnor UO_538 (O_538,N_4773,N_4418);
xnor UO_539 (O_539,N_4508,N_4598);
nor UO_540 (O_540,N_4480,N_4362);
nor UO_541 (O_541,N_4900,N_4509);
nand UO_542 (O_542,N_4460,N_4785);
xor UO_543 (O_543,N_4574,N_4935);
or UO_544 (O_544,N_4216,N_4550);
xnor UO_545 (O_545,N_4465,N_4914);
xnor UO_546 (O_546,N_4530,N_4149);
nor UO_547 (O_547,N_4610,N_4175);
or UO_548 (O_548,N_4240,N_4349);
nor UO_549 (O_549,N_4330,N_4788);
or UO_550 (O_550,N_4767,N_4528);
xor UO_551 (O_551,N_4342,N_4068);
nor UO_552 (O_552,N_4183,N_4007);
nor UO_553 (O_553,N_4398,N_4178);
nand UO_554 (O_554,N_4094,N_4971);
xnor UO_555 (O_555,N_4447,N_4621);
nor UO_556 (O_556,N_4899,N_4739);
and UO_557 (O_557,N_4268,N_4155);
or UO_558 (O_558,N_4437,N_4861);
nor UO_559 (O_559,N_4140,N_4727);
nor UO_560 (O_560,N_4635,N_4082);
nand UO_561 (O_561,N_4240,N_4678);
or UO_562 (O_562,N_4885,N_4399);
xnor UO_563 (O_563,N_4589,N_4975);
xor UO_564 (O_564,N_4520,N_4366);
or UO_565 (O_565,N_4489,N_4050);
and UO_566 (O_566,N_4752,N_4601);
xor UO_567 (O_567,N_4745,N_4532);
and UO_568 (O_568,N_4225,N_4677);
xor UO_569 (O_569,N_4863,N_4192);
or UO_570 (O_570,N_4201,N_4896);
nand UO_571 (O_571,N_4157,N_4244);
and UO_572 (O_572,N_4716,N_4422);
and UO_573 (O_573,N_4302,N_4160);
and UO_574 (O_574,N_4667,N_4689);
xor UO_575 (O_575,N_4593,N_4415);
nor UO_576 (O_576,N_4814,N_4810);
and UO_577 (O_577,N_4263,N_4175);
xnor UO_578 (O_578,N_4493,N_4741);
nor UO_579 (O_579,N_4910,N_4561);
nand UO_580 (O_580,N_4664,N_4444);
and UO_581 (O_581,N_4461,N_4804);
nand UO_582 (O_582,N_4212,N_4917);
nand UO_583 (O_583,N_4140,N_4417);
nand UO_584 (O_584,N_4326,N_4890);
and UO_585 (O_585,N_4338,N_4206);
or UO_586 (O_586,N_4470,N_4385);
nor UO_587 (O_587,N_4105,N_4394);
and UO_588 (O_588,N_4407,N_4189);
xor UO_589 (O_589,N_4189,N_4714);
nor UO_590 (O_590,N_4907,N_4119);
and UO_591 (O_591,N_4357,N_4422);
xor UO_592 (O_592,N_4347,N_4880);
or UO_593 (O_593,N_4451,N_4557);
xnor UO_594 (O_594,N_4823,N_4918);
nor UO_595 (O_595,N_4069,N_4989);
nand UO_596 (O_596,N_4072,N_4676);
nand UO_597 (O_597,N_4991,N_4859);
nor UO_598 (O_598,N_4135,N_4126);
and UO_599 (O_599,N_4064,N_4025);
nor UO_600 (O_600,N_4107,N_4443);
or UO_601 (O_601,N_4446,N_4026);
nor UO_602 (O_602,N_4864,N_4985);
nor UO_603 (O_603,N_4986,N_4823);
or UO_604 (O_604,N_4899,N_4974);
nand UO_605 (O_605,N_4279,N_4601);
and UO_606 (O_606,N_4792,N_4847);
or UO_607 (O_607,N_4338,N_4967);
xnor UO_608 (O_608,N_4541,N_4135);
xor UO_609 (O_609,N_4193,N_4324);
nand UO_610 (O_610,N_4625,N_4728);
xnor UO_611 (O_611,N_4792,N_4715);
nor UO_612 (O_612,N_4754,N_4836);
nor UO_613 (O_613,N_4757,N_4133);
nand UO_614 (O_614,N_4300,N_4998);
nor UO_615 (O_615,N_4845,N_4625);
and UO_616 (O_616,N_4325,N_4146);
or UO_617 (O_617,N_4281,N_4820);
xor UO_618 (O_618,N_4717,N_4585);
nand UO_619 (O_619,N_4061,N_4284);
or UO_620 (O_620,N_4183,N_4849);
xor UO_621 (O_621,N_4329,N_4420);
or UO_622 (O_622,N_4414,N_4048);
or UO_623 (O_623,N_4565,N_4687);
and UO_624 (O_624,N_4542,N_4883);
and UO_625 (O_625,N_4171,N_4576);
or UO_626 (O_626,N_4124,N_4243);
nor UO_627 (O_627,N_4848,N_4795);
or UO_628 (O_628,N_4390,N_4529);
and UO_629 (O_629,N_4623,N_4983);
and UO_630 (O_630,N_4598,N_4820);
xor UO_631 (O_631,N_4014,N_4151);
or UO_632 (O_632,N_4205,N_4676);
nand UO_633 (O_633,N_4314,N_4533);
or UO_634 (O_634,N_4468,N_4713);
nand UO_635 (O_635,N_4509,N_4749);
xor UO_636 (O_636,N_4677,N_4942);
and UO_637 (O_637,N_4716,N_4272);
and UO_638 (O_638,N_4892,N_4302);
nand UO_639 (O_639,N_4685,N_4727);
nor UO_640 (O_640,N_4411,N_4373);
nor UO_641 (O_641,N_4802,N_4619);
or UO_642 (O_642,N_4395,N_4307);
xor UO_643 (O_643,N_4568,N_4595);
nor UO_644 (O_644,N_4374,N_4698);
or UO_645 (O_645,N_4801,N_4374);
or UO_646 (O_646,N_4610,N_4942);
xnor UO_647 (O_647,N_4048,N_4412);
nor UO_648 (O_648,N_4579,N_4947);
nor UO_649 (O_649,N_4968,N_4889);
and UO_650 (O_650,N_4921,N_4831);
nor UO_651 (O_651,N_4806,N_4542);
xor UO_652 (O_652,N_4861,N_4447);
xor UO_653 (O_653,N_4086,N_4264);
xor UO_654 (O_654,N_4131,N_4948);
nor UO_655 (O_655,N_4307,N_4448);
nor UO_656 (O_656,N_4014,N_4823);
nor UO_657 (O_657,N_4164,N_4961);
or UO_658 (O_658,N_4884,N_4576);
and UO_659 (O_659,N_4117,N_4378);
or UO_660 (O_660,N_4485,N_4228);
nand UO_661 (O_661,N_4313,N_4031);
or UO_662 (O_662,N_4149,N_4685);
and UO_663 (O_663,N_4501,N_4224);
xor UO_664 (O_664,N_4305,N_4171);
xor UO_665 (O_665,N_4380,N_4281);
or UO_666 (O_666,N_4440,N_4837);
and UO_667 (O_667,N_4568,N_4708);
or UO_668 (O_668,N_4603,N_4120);
xnor UO_669 (O_669,N_4935,N_4579);
and UO_670 (O_670,N_4834,N_4659);
nor UO_671 (O_671,N_4371,N_4369);
nor UO_672 (O_672,N_4204,N_4361);
xor UO_673 (O_673,N_4959,N_4277);
and UO_674 (O_674,N_4797,N_4337);
and UO_675 (O_675,N_4244,N_4305);
and UO_676 (O_676,N_4109,N_4411);
and UO_677 (O_677,N_4300,N_4825);
or UO_678 (O_678,N_4200,N_4375);
xnor UO_679 (O_679,N_4966,N_4746);
or UO_680 (O_680,N_4230,N_4331);
nor UO_681 (O_681,N_4540,N_4591);
xor UO_682 (O_682,N_4362,N_4113);
or UO_683 (O_683,N_4830,N_4672);
and UO_684 (O_684,N_4019,N_4816);
nor UO_685 (O_685,N_4575,N_4636);
or UO_686 (O_686,N_4406,N_4514);
nand UO_687 (O_687,N_4603,N_4627);
nor UO_688 (O_688,N_4331,N_4176);
nand UO_689 (O_689,N_4638,N_4936);
nor UO_690 (O_690,N_4207,N_4632);
nor UO_691 (O_691,N_4459,N_4446);
nor UO_692 (O_692,N_4250,N_4955);
nor UO_693 (O_693,N_4602,N_4004);
xnor UO_694 (O_694,N_4069,N_4807);
and UO_695 (O_695,N_4503,N_4208);
or UO_696 (O_696,N_4013,N_4427);
nor UO_697 (O_697,N_4206,N_4389);
nor UO_698 (O_698,N_4657,N_4959);
nor UO_699 (O_699,N_4589,N_4795);
and UO_700 (O_700,N_4489,N_4833);
or UO_701 (O_701,N_4689,N_4924);
or UO_702 (O_702,N_4559,N_4822);
and UO_703 (O_703,N_4778,N_4568);
nand UO_704 (O_704,N_4352,N_4619);
xor UO_705 (O_705,N_4708,N_4363);
or UO_706 (O_706,N_4752,N_4134);
xnor UO_707 (O_707,N_4997,N_4634);
nand UO_708 (O_708,N_4195,N_4842);
nor UO_709 (O_709,N_4988,N_4779);
and UO_710 (O_710,N_4188,N_4743);
xnor UO_711 (O_711,N_4005,N_4377);
xor UO_712 (O_712,N_4695,N_4433);
nor UO_713 (O_713,N_4112,N_4037);
xor UO_714 (O_714,N_4207,N_4675);
nor UO_715 (O_715,N_4750,N_4591);
nand UO_716 (O_716,N_4414,N_4271);
or UO_717 (O_717,N_4451,N_4996);
and UO_718 (O_718,N_4912,N_4668);
nand UO_719 (O_719,N_4717,N_4076);
xnor UO_720 (O_720,N_4219,N_4843);
nor UO_721 (O_721,N_4150,N_4800);
nand UO_722 (O_722,N_4314,N_4276);
xnor UO_723 (O_723,N_4172,N_4092);
xnor UO_724 (O_724,N_4344,N_4783);
or UO_725 (O_725,N_4582,N_4524);
xnor UO_726 (O_726,N_4863,N_4024);
nand UO_727 (O_727,N_4619,N_4562);
and UO_728 (O_728,N_4599,N_4310);
nand UO_729 (O_729,N_4830,N_4077);
or UO_730 (O_730,N_4429,N_4825);
or UO_731 (O_731,N_4418,N_4623);
nor UO_732 (O_732,N_4514,N_4538);
or UO_733 (O_733,N_4163,N_4020);
nor UO_734 (O_734,N_4564,N_4501);
and UO_735 (O_735,N_4702,N_4046);
or UO_736 (O_736,N_4047,N_4058);
or UO_737 (O_737,N_4434,N_4771);
nor UO_738 (O_738,N_4529,N_4498);
nand UO_739 (O_739,N_4516,N_4402);
xor UO_740 (O_740,N_4828,N_4712);
nand UO_741 (O_741,N_4856,N_4089);
nand UO_742 (O_742,N_4395,N_4254);
and UO_743 (O_743,N_4625,N_4944);
nor UO_744 (O_744,N_4116,N_4736);
nor UO_745 (O_745,N_4833,N_4003);
xor UO_746 (O_746,N_4100,N_4233);
xor UO_747 (O_747,N_4451,N_4559);
or UO_748 (O_748,N_4902,N_4413);
nor UO_749 (O_749,N_4767,N_4904);
xor UO_750 (O_750,N_4286,N_4954);
or UO_751 (O_751,N_4621,N_4521);
or UO_752 (O_752,N_4912,N_4124);
xor UO_753 (O_753,N_4234,N_4002);
nand UO_754 (O_754,N_4554,N_4137);
and UO_755 (O_755,N_4942,N_4225);
nor UO_756 (O_756,N_4232,N_4155);
xnor UO_757 (O_757,N_4655,N_4024);
nor UO_758 (O_758,N_4107,N_4878);
and UO_759 (O_759,N_4473,N_4146);
and UO_760 (O_760,N_4743,N_4900);
xor UO_761 (O_761,N_4616,N_4575);
xor UO_762 (O_762,N_4149,N_4138);
or UO_763 (O_763,N_4272,N_4780);
nand UO_764 (O_764,N_4859,N_4717);
and UO_765 (O_765,N_4946,N_4723);
xor UO_766 (O_766,N_4637,N_4034);
or UO_767 (O_767,N_4395,N_4245);
nor UO_768 (O_768,N_4592,N_4864);
nor UO_769 (O_769,N_4045,N_4087);
xor UO_770 (O_770,N_4518,N_4056);
nor UO_771 (O_771,N_4269,N_4257);
and UO_772 (O_772,N_4617,N_4381);
nor UO_773 (O_773,N_4482,N_4333);
nand UO_774 (O_774,N_4016,N_4477);
xnor UO_775 (O_775,N_4711,N_4084);
or UO_776 (O_776,N_4450,N_4536);
xor UO_777 (O_777,N_4805,N_4331);
xnor UO_778 (O_778,N_4844,N_4749);
and UO_779 (O_779,N_4911,N_4536);
and UO_780 (O_780,N_4689,N_4382);
and UO_781 (O_781,N_4786,N_4061);
xnor UO_782 (O_782,N_4647,N_4776);
and UO_783 (O_783,N_4531,N_4941);
or UO_784 (O_784,N_4323,N_4362);
xor UO_785 (O_785,N_4782,N_4290);
nor UO_786 (O_786,N_4037,N_4585);
and UO_787 (O_787,N_4772,N_4080);
nand UO_788 (O_788,N_4685,N_4631);
and UO_789 (O_789,N_4019,N_4725);
nand UO_790 (O_790,N_4565,N_4517);
nor UO_791 (O_791,N_4678,N_4505);
or UO_792 (O_792,N_4565,N_4198);
xor UO_793 (O_793,N_4477,N_4249);
nand UO_794 (O_794,N_4952,N_4785);
nor UO_795 (O_795,N_4526,N_4535);
or UO_796 (O_796,N_4543,N_4062);
nand UO_797 (O_797,N_4943,N_4739);
nand UO_798 (O_798,N_4483,N_4024);
xor UO_799 (O_799,N_4875,N_4297);
nor UO_800 (O_800,N_4595,N_4216);
xnor UO_801 (O_801,N_4160,N_4393);
nand UO_802 (O_802,N_4836,N_4283);
and UO_803 (O_803,N_4427,N_4120);
or UO_804 (O_804,N_4250,N_4631);
xor UO_805 (O_805,N_4649,N_4275);
xor UO_806 (O_806,N_4470,N_4530);
nor UO_807 (O_807,N_4108,N_4127);
and UO_808 (O_808,N_4495,N_4028);
xnor UO_809 (O_809,N_4544,N_4862);
nor UO_810 (O_810,N_4618,N_4156);
or UO_811 (O_811,N_4636,N_4571);
nor UO_812 (O_812,N_4775,N_4563);
nand UO_813 (O_813,N_4219,N_4549);
xnor UO_814 (O_814,N_4779,N_4490);
or UO_815 (O_815,N_4205,N_4514);
and UO_816 (O_816,N_4504,N_4553);
and UO_817 (O_817,N_4774,N_4824);
nand UO_818 (O_818,N_4118,N_4683);
nor UO_819 (O_819,N_4838,N_4384);
and UO_820 (O_820,N_4819,N_4016);
nor UO_821 (O_821,N_4766,N_4845);
and UO_822 (O_822,N_4019,N_4145);
nand UO_823 (O_823,N_4012,N_4683);
nand UO_824 (O_824,N_4778,N_4912);
xnor UO_825 (O_825,N_4204,N_4760);
nand UO_826 (O_826,N_4930,N_4253);
xnor UO_827 (O_827,N_4538,N_4619);
and UO_828 (O_828,N_4216,N_4504);
nor UO_829 (O_829,N_4040,N_4120);
nor UO_830 (O_830,N_4546,N_4377);
xor UO_831 (O_831,N_4360,N_4506);
nand UO_832 (O_832,N_4633,N_4323);
or UO_833 (O_833,N_4635,N_4523);
and UO_834 (O_834,N_4984,N_4601);
xor UO_835 (O_835,N_4446,N_4966);
or UO_836 (O_836,N_4681,N_4304);
or UO_837 (O_837,N_4086,N_4690);
xor UO_838 (O_838,N_4803,N_4673);
nor UO_839 (O_839,N_4916,N_4711);
nand UO_840 (O_840,N_4201,N_4322);
xnor UO_841 (O_841,N_4121,N_4459);
nand UO_842 (O_842,N_4936,N_4333);
xor UO_843 (O_843,N_4160,N_4266);
nand UO_844 (O_844,N_4915,N_4790);
xor UO_845 (O_845,N_4771,N_4885);
or UO_846 (O_846,N_4800,N_4980);
and UO_847 (O_847,N_4260,N_4546);
nand UO_848 (O_848,N_4075,N_4925);
xnor UO_849 (O_849,N_4353,N_4976);
nor UO_850 (O_850,N_4424,N_4764);
xor UO_851 (O_851,N_4098,N_4425);
or UO_852 (O_852,N_4513,N_4551);
xor UO_853 (O_853,N_4069,N_4344);
and UO_854 (O_854,N_4430,N_4052);
or UO_855 (O_855,N_4893,N_4456);
xnor UO_856 (O_856,N_4396,N_4575);
or UO_857 (O_857,N_4902,N_4475);
and UO_858 (O_858,N_4103,N_4112);
and UO_859 (O_859,N_4409,N_4304);
nand UO_860 (O_860,N_4982,N_4344);
or UO_861 (O_861,N_4743,N_4081);
xnor UO_862 (O_862,N_4471,N_4526);
xor UO_863 (O_863,N_4496,N_4463);
nor UO_864 (O_864,N_4756,N_4245);
and UO_865 (O_865,N_4260,N_4672);
and UO_866 (O_866,N_4861,N_4759);
nor UO_867 (O_867,N_4979,N_4526);
nand UO_868 (O_868,N_4518,N_4791);
nor UO_869 (O_869,N_4666,N_4849);
and UO_870 (O_870,N_4562,N_4673);
nand UO_871 (O_871,N_4892,N_4834);
nor UO_872 (O_872,N_4499,N_4741);
xor UO_873 (O_873,N_4921,N_4770);
nor UO_874 (O_874,N_4482,N_4528);
or UO_875 (O_875,N_4003,N_4608);
xnor UO_876 (O_876,N_4268,N_4313);
and UO_877 (O_877,N_4307,N_4777);
xnor UO_878 (O_878,N_4813,N_4271);
nand UO_879 (O_879,N_4067,N_4675);
nor UO_880 (O_880,N_4818,N_4097);
and UO_881 (O_881,N_4807,N_4044);
nand UO_882 (O_882,N_4207,N_4199);
and UO_883 (O_883,N_4643,N_4561);
xnor UO_884 (O_884,N_4951,N_4108);
xor UO_885 (O_885,N_4984,N_4109);
xor UO_886 (O_886,N_4146,N_4249);
nand UO_887 (O_887,N_4160,N_4371);
or UO_888 (O_888,N_4759,N_4553);
or UO_889 (O_889,N_4921,N_4737);
nand UO_890 (O_890,N_4931,N_4343);
nor UO_891 (O_891,N_4385,N_4967);
or UO_892 (O_892,N_4004,N_4427);
nor UO_893 (O_893,N_4224,N_4730);
and UO_894 (O_894,N_4309,N_4911);
or UO_895 (O_895,N_4848,N_4046);
or UO_896 (O_896,N_4171,N_4901);
nor UO_897 (O_897,N_4240,N_4013);
or UO_898 (O_898,N_4411,N_4890);
xnor UO_899 (O_899,N_4432,N_4139);
nand UO_900 (O_900,N_4676,N_4717);
or UO_901 (O_901,N_4072,N_4390);
xor UO_902 (O_902,N_4871,N_4995);
nand UO_903 (O_903,N_4226,N_4249);
nand UO_904 (O_904,N_4873,N_4528);
or UO_905 (O_905,N_4689,N_4753);
or UO_906 (O_906,N_4364,N_4008);
or UO_907 (O_907,N_4051,N_4855);
nor UO_908 (O_908,N_4016,N_4623);
xnor UO_909 (O_909,N_4874,N_4331);
or UO_910 (O_910,N_4522,N_4162);
nor UO_911 (O_911,N_4145,N_4702);
and UO_912 (O_912,N_4464,N_4377);
xnor UO_913 (O_913,N_4887,N_4276);
and UO_914 (O_914,N_4362,N_4007);
and UO_915 (O_915,N_4453,N_4144);
xor UO_916 (O_916,N_4995,N_4454);
and UO_917 (O_917,N_4404,N_4671);
xnor UO_918 (O_918,N_4672,N_4670);
and UO_919 (O_919,N_4249,N_4046);
nand UO_920 (O_920,N_4780,N_4901);
nand UO_921 (O_921,N_4389,N_4364);
xor UO_922 (O_922,N_4039,N_4292);
nand UO_923 (O_923,N_4655,N_4310);
and UO_924 (O_924,N_4903,N_4597);
nor UO_925 (O_925,N_4394,N_4265);
xor UO_926 (O_926,N_4875,N_4206);
or UO_927 (O_927,N_4540,N_4845);
nand UO_928 (O_928,N_4337,N_4652);
and UO_929 (O_929,N_4495,N_4511);
and UO_930 (O_930,N_4784,N_4005);
nand UO_931 (O_931,N_4590,N_4040);
and UO_932 (O_932,N_4030,N_4069);
nand UO_933 (O_933,N_4250,N_4696);
or UO_934 (O_934,N_4233,N_4588);
and UO_935 (O_935,N_4272,N_4054);
and UO_936 (O_936,N_4709,N_4850);
or UO_937 (O_937,N_4268,N_4492);
nand UO_938 (O_938,N_4702,N_4974);
nand UO_939 (O_939,N_4642,N_4293);
nand UO_940 (O_940,N_4387,N_4212);
xor UO_941 (O_941,N_4873,N_4747);
nand UO_942 (O_942,N_4818,N_4755);
nand UO_943 (O_943,N_4407,N_4449);
and UO_944 (O_944,N_4557,N_4468);
nand UO_945 (O_945,N_4245,N_4459);
or UO_946 (O_946,N_4407,N_4428);
nand UO_947 (O_947,N_4517,N_4848);
nand UO_948 (O_948,N_4191,N_4144);
nor UO_949 (O_949,N_4107,N_4608);
and UO_950 (O_950,N_4142,N_4433);
nand UO_951 (O_951,N_4734,N_4788);
xnor UO_952 (O_952,N_4096,N_4856);
or UO_953 (O_953,N_4595,N_4387);
nor UO_954 (O_954,N_4643,N_4040);
or UO_955 (O_955,N_4908,N_4171);
nand UO_956 (O_956,N_4832,N_4468);
nor UO_957 (O_957,N_4334,N_4216);
or UO_958 (O_958,N_4858,N_4548);
xor UO_959 (O_959,N_4585,N_4179);
nand UO_960 (O_960,N_4601,N_4472);
xor UO_961 (O_961,N_4131,N_4912);
and UO_962 (O_962,N_4678,N_4539);
or UO_963 (O_963,N_4617,N_4948);
nor UO_964 (O_964,N_4771,N_4394);
nor UO_965 (O_965,N_4222,N_4244);
and UO_966 (O_966,N_4076,N_4488);
or UO_967 (O_967,N_4479,N_4097);
and UO_968 (O_968,N_4943,N_4769);
and UO_969 (O_969,N_4961,N_4108);
and UO_970 (O_970,N_4860,N_4056);
xor UO_971 (O_971,N_4097,N_4689);
and UO_972 (O_972,N_4535,N_4532);
xor UO_973 (O_973,N_4580,N_4057);
or UO_974 (O_974,N_4548,N_4488);
nor UO_975 (O_975,N_4981,N_4740);
nand UO_976 (O_976,N_4418,N_4324);
or UO_977 (O_977,N_4109,N_4289);
nor UO_978 (O_978,N_4627,N_4551);
and UO_979 (O_979,N_4740,N_4852);
xnor UO_980 (O_980,N_4044,N_4274);
nand UO_981 (O_981,N_4344,N_4382);
or UO_982 (O_982,N_4872,N_4618);
or UO_983 (O_983,N_4421,N_4740);
and UO_984 (O_984,N_4471,N_4380);
and UO_985 (O_985,N_4519,N_4823);
nor UO_986 (O_986,N_4200,N_4003);
or UO_987 (O_987,N_4813,N_4938);
or UO_988 (O_988,N_4326,N_4163);
or UO_989 (O_989,N_4795,N_4587);
nand UO_990 (O_990,N_4638,N_4585);
nand UO_991 (O_991,N_4534,N_4116);
nand UO_992 (O_992,N_4692,N_4938);
nor UO_993 (O_993,N_4692,N_4438);
or UO_994 (O_994,N_4690,N_4042);
or UO_995 (O_995,N_4614,N_4784);
or UO_996 (O_996,N_4589,N_4422);
nor UO_997 (O_997,N_4996,N_4477);
nand UO_998 (O_998,N_4309,N_4062);
xor UO_999 (O_999,N_4929,N_4254);
endmodule