module basic_500_3000_500_15_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_347,In_128);
nor U1 (N_1,In_325,In_248);
xnor U2 (N_2,In_384,In_396);
nor U3 (N_3,In_395,In_392);
nand U4 (N_4,In_198,In_57);
nand U5 (N_5,In_59,In_357);
and U6 (N_6,In_235,In_213);
nand U7 (N_7,In_363,In_473);
nand U8 (N_8,In_63,In_24);
nor U9 (N_9,In_191,In_484);
and U10 (N_10,In_405,In_138);
nand U11 (N_11,In_452,In_38);
nor U12 (N_12,In_418,In_237);
xnor U13 (N_13,In_121,In_48);
nor U14 (N_14,In_348,In_284);
and U15 (N_15,In_375,In_17);
xor U16 (N_16,In_87,In_261);
nor U17 (N_17,In_426,In_136);
nand U18 (N_18,In_303,In_156);
and U19 (N_19,In_196,In_374);
or U20 (N_20,In_293,In_155);
or U21 (N_21,In_360,In_144);
and U22 (N_22,In_41,In_294);
nand U23 (N_23,In_328,In_349);
or U24 (N_24,In_234,In_66);
nand U25 (N_25,In_414,In_182);
nor U26 (N_26,In_68,In_30);
nor U27 (N_27,In_70,In_65);
and U28 (N_28,In_290,In_166);
nand U29 (N_29,In_483,In_232);
and U30 (N_30,In_252,In_139);
and U31 (N_31,In_269,In_117);
xor U32 (N_32,In_11,In_238);
nand U33 (N_33,In_310,In_437);
nand U34 (N_34,In_254,In_211);
and U35 (N_35,In_250,In_297);
nand U36 (N_36,In_226,In_147);
or U37 (N_37,In_258,In_8);
nor U38 (N_38,In_399,In_280);
or U39 (N_39,In_377,In_407);
nand U40 (N_40,In_150,In_390);
nor U41 (N_41,In_169,In_108);
nand U42 (N_42,In_340,In_130);
and U43 (N_43,In_338,In_435);
or U44 (N_44,In_380,In_351);
nor U45 (N_45,In_80,In_105);
nor U46 (N_46,In_436,In_402);
nor U47 (N_47,In_445,In_382);
and U48 (N_48,In_123,In_22);
and U49 (N_49,In_200,In_321);
or U50 (N_50,In_164,In_79);
nor U51 (N_51,In_486,In_223);
nand U52 (N_52,In_316,In_255);
xor U53 (N_53,In_115,In_352);
nor U54 (N_54,In_20,In_85);
and U55 (N_55,In_214,In_141);
xor U56 (N_56,In_387,In_165);
nand U57 (N_57,In_151,In_39);
nor U58 (N_58,In_163,In_314);
nand U59 (N_59,In_247,In_460);
and U60 (N_60,In_461,In_344);
or U61 (N_61,In_192,In_172);
or U62 (N_62,In_64,In_378);
nor U63 (N_63,In_113,In_112);
nand U64 (N_64,In_116,In_89);
and U65 (N_65,In_459,In_127);
nand U66 (N_66,In_187,In_446);
or U67 (N_67,In_370,In_170);
nand U68 (N_68,In_388,In_137);
or U69 (N_69,In_448,In_83);
nor U70 (N_70,In_109,In_225);
and U71 (N_71,In_14,In_286);
nand U72 (N_72,In_84,In_391);
and U73 (N_73,In_21,In_222);
nand U74 (N_74,In_94,In_404);
nand U75 (N_75,In_145,In_309);
and U76 (N_76,In_272,In_288);
and U77 (N_77,In_364,In_133);
or U78 (N_78,In_249,In_494);
nor U79 (N_79,In_32,In_443);
and U80 (N_80,In_28,In_300);
nand U81 (N_81,In_330,In_468);
nand U82 (N_82,In_323,In_474);
nor U83 (N_83,In_311,In_273);
and U84 (N_84,In_126,In_184);
and U85 (N_85,In_171,In_168);
and U86 (N_86,In_206,In_148);
nand U87 (N_87,In_190,In_240);
nor U88 (N_88,In_134,In_203);
or U89 (N_89,In_4,In_422);
or U90 (N_90,In_274,In_244);
nor U91 (N_91,In_317,In_478);
or U92 (N_92,In_413,In_42);
and U93 (N_93,In_119,In_408);
nor U94 (N_94,In_81,In_209);
and U95 (N_95,In_231,In_86);
xnor U96 (N_96,In_427,In_406);
or U97 (N_97,In_415,In_356);
nor U98 (N_98,In_264,In_471);
or U99 (N_99,In_282,In_266);
or U100 (N_100,In_224,In_424);
and U101 (N_101,In_322,In_246);
and U102 (N_102,In_416,In_161);
or U103 (N_103,In_10,In_29);
or U104 (N_104,In_5,In_178);
or U105 (N_105,In_227,In_174);
nand U106 (N_106,In_475,In_101);
nor U107 (N_107,In_37,In_194);
and U108 (N_108,In_393,In_90);
nor U109 (N_109,In_152,In_346);
nor U110 (N_110,In_495,In_104);
nor U111 (N_111,In_215,In_103);
nand U112 (N_112,In_270,In_99);
nand U113 (N_113,In_146,In_98);
nor U114 (N_114,In_132,In_239);
nor U115 (N_115,In_485,In_7);
nand U116 (N_116,In_498,In_299);
nand U117 (N_117,In_308,In_434);
and U118 (N_118,In_36,In_97);
or U119 (N_119,In_464,In_219);
nor U120 (N_120,In_275,In_491);
nor U121 (N_121,In_135,In_467);
nand U122 (N_122,In_447,In_373);
and U123 (N_123,In_401,In_315);
and U124 (N_124,In_173,In_193);
nor U125 (N_125,In_55,In_444);
nor U126 (N_126,In_362,In_440);
nand U127 (N_127,In_449,In_319);
nand U128 (N_128,In_279,In_381);
and U129 (N_129,In_221,In_15);
or U130 (N_130,In_49,In_16);
nor U131 (N_131,In_409,In_490);
xnor U132 (N_132,In_253,In_432);
nor U133 (N_133,In_389,In_285);
and U134 (N_134,In_358,In_180);
nand U135 (N_135,In_27,In_359);
and U136 (N_136,In_78,In_210);
and U137 (N_137,In_431,In_442);
nor U138 (N_138,In_75,In_241);
and U139 (N_139,In_430,In_74);
nor U140 (N_140,In_267,In_218);
nand U141 (N_141,In_296,In_457);
or U142 (N_142,In_106,In_175);
nand U143 (N_143,In_125,In_228);
or U144 (N_144,In_201,In_383);
nor U145 (N_145,In_92,In_167);
or U146 (N_146,In_312,In_34);
nand U147 (N_147,In_394,In_499);
xor U148 (N_148,In_410,In_292);
and U149 (N_149,In_230,In_281);
and U150 (N_150,In_260,In_369);
nand U151 (N_151,In_3,In_428);
nand U152 (N_152,In_276,In_33);
nand U153 (N_153,In_53,In_243);
nand U154 (N_154,In_331,In_496);
or U155 (N_155,In_236,In_111);
nor U156 (N_156,In_333,In_76);
nand U157 (N_157,In_259,In_417);
nor U158 (N_158,In_301,In_477);
and U159 (N_159,In_2,In_385);
or U160 (N_160,In_176,In_283);
nand U161 (N_161,In_412,In_188);
and U162 (N_162,In_454,In_423);
nand U163 (N_163,In_229,In_463);
nand U164 (N_164,In_307,In_455);
or U165 (N_165,In_419,In_93);
or U166 (N_166,In_96,In_204);
nand U167 (N_167,In_54,In_361);
nand U168 (N_168,In_158,In_289);
or U169 (N_169,In_306,In_487);
xor U170 (N_170,In_277,In_304);
nand U171 (N_171,In_372,In_398);
and U172 (N_172,In_52,In_397);
or U173 (N_173,In_199,In_45);
nand U174 (N_174,In_479,In_489);
or U175 (N_175,In_313,In_386);
or U176 (N_176,In_82,In_476);
nor U177 (N_177,In_324,In_140);
or U178 (N_178,In_343,In_162);
and U179 (N_179,In_492,In_149);
nand U180 (N_180,In_451,In_6);
or U181 (N_181,In_107,In_441);
nor U182 (N_182,In_43,In_450);
or U183 (N_183,In_403,In_154);
nand U184 (N_184,In_302,In_497);
or U185 (N_185,In_124,In_298);
or U186 (N_186,In_50,In_71);
and U187 (N_187,In_62,In_212);
nor U188 (N_188,In_9,In_35);
nand U189 (N_189,In_263,In_371);
or U190 (N_190,In_207,In_482);
or U191 (N_191,In_353,In_18);
or U192 (N_192,In_329,In_339);
or U193 (N_193,In_466,In_72);
and U194 (N_194,In_185,In_271);
and U195 (N_195,In_23,In_189);
or U196 (N_196,In_12,In_488);
nand U197 (N_197,In_143,In_77);
or U198 (N_198,In_268,In_100);
and U199 (N_199,In_291,In_425);
nand U200 (N_200,N_73,In_217);
or U201 (N_201,N_60,N_115);
and U202 (N_202,N_102,N_62);
and U203 (N_203,N_160,In_129);
or U204 (N_204,In_157,N_125);
or U205 (N_205,N_113,In_400);
nor U206 (N_206,N_87,N_130);
or U207 (N_207,In_122,N_98);
nor U208 (N_208,N_18,N_153);
nand U209 (N_209,N_33,N_191);
and U210 (N_210,In_368,In_118);
and U211 (N_211,N_68,N_78);
nand U212 (N_212,N_91,N_96);
xnor U213 (N_213,N_37,N_19);
nor U214 (N_214,In_0,In_480);
and U215 (N_215,In_257,In_183);
nand U216 (N_216,N_190,N_136);
or U217 (N_217,N_44,N_5);
and U218 (N_218,N_69,N_141);
nand U219 (N_219,N_181,N_114);
or U220 (N_220,N_71,In_470);
xor U221 (N_221,N_144,In_242);
and U222 (N_222,In_481,N_120);
nor U223 (N_223,N_170,In_334);
or U224 (N_224,N_47,N_151);
nand U225 (N_225,N_199,In_453);
nor U226 (N_226,N_74,N_196);
nor U227 (N_227,N_67,N_110);
nand U228 (N_228,N_122,In_456);
and U229 (N_229,In_114,N_27);
xor U230 (N_230,N_180,N_16);
nand U231 (N_231,N_127,N_58);
nor U232 (N_232,In_95,N_3);
and U233 (N_233,N_81,In_429);
or U234 (N_234,In_278,N_10);
nor U235 (N_235,In_265,N_145);
and U236 (N_236,N_34,N_111);
nor U237 (N_237,N_172,In_411);
and U238 (N_238,N_20,In_195);
xor U239 (N_239,In_131,In_465);
nand U240 (N_240,In_202,In_1);
nor U241 (N_241,N_107,N_198);
or U242 (N_242,In_67,N_30);
nor U243 (N_243,N_168,In_73);
or U244 (N_244,In_341,N_41);
nor U245 (N_245,N_133,N_86);
and U246 (N_246,In_19,In_159);
nor U247 (N_247,N_171,N_162);
nand U248 (N_248,In_26,N_21);
and U249 (N_249,N_12,N_105);
nor U250 (N_250,In_320,N_36);
and U251 (N_251,In_245,N_26);
nor U252 (N_252,In_354,N_97);
or U253 (N_253,N_189,In_69);
or U254 (N_254,In_469,N_85);
nor U255 (N_255,In_433,N_15);
and U256 (N_256,N_152,N_24);
or U257 (N_257,In_181,N_89);
nor U258 (N_258,In_305,N_43);
nor U259 (N_259,In_439,In_177);
and U260 (N_260,In_355,N_59);
and U261 (N_261,N_179,N_75);
xor U262 (N_262,In_56,N_65);
nor U263 (N_263,N_175,In_251);
nand U264 (N_264,In_365,In_366);
and U265 (N_265,N_148,N_147);
or U266 (N_266,In_216,In_256);
or U267 (N_267,N_195,N_157);
or U268 (N_268,In_262,N_51);
or U269 (N_269,N_80,N_95);
and U270 (N_270,N_29,N_174);
or U271 (N_271,N_11,N_119);
xor U272 (N_272,N_139,In_472);
and U273 (N_273,N_117,N_84);
nand U274 (N_274,N_116,In_318);
nor U275 (N_275,In_345,In_142);
xor U276 (N_276,N_132,N_45);
and U277 (N_277,In_153,N_158);
xnor U278 (N_278,N_88,In_295);
and U279 (N_279,In_102,In_350);
or U280 (N_280,N_77,N_137);
nor U281 (N_281,N_94,N_138);
nand U282 (N_282,N_169,In_110);
nand U283 (N_283,In_208,N_14);
and U284 (N_284,In_120,N_23);
and U285 (N_285,In_46,In_438);
or U286 (N_286,N_48,N_129);
nand U287 (N_287,N_104,N_142);
or U288 (N_288,N_123,N_177);
and U289 (N_289,N_9,N_99);
nor U290 (N_290,N_56,N_22);
or U291 (N_291,In_421,N_92);
nor U292 (N_292,N_112,N_118);
and U293 (N_293,N_140,N_156);
and U294 (N_294,N_63,N_83);
nor U295 (N_295,In_205,N_173);
nand U296 (N_296,In_47,In_367);
nand U297 (N_297,N_165,In_60);
nor U298 (N_298,In_326,N_167);
xor U299 (N_299,In_462,N_108);
and U300 (N_300,N_13,N_155);
or U301 (N_301,N_39,N_46);
nand U302 (N_302,N_176,N_194);
or U303 (N_303,N_17,N_70);
and U304 (N_304,N_76,In_342);
and U305 (N_305,In_327,N_7);
nand U306 (N_306,N_55,In_197);
nor U307 (N_307,N_6,N_187);
nor U308 (N_308,N_188,N_28);
nand U309 (N_309,In_88,N_53);
nor U310 (N_310,N_25,N_106);
nor U311 (N_311,N_154,N_103);
xnor U312 (N_312,N_4,In_160);
or U313 (N_313,N_150,N_124);
nor U314 (N_314,N_143,N_93);
xnor U315 (N_315,N_49,N_2);
nand U316 (N_316,N_31,N_146);
xor U317 (N_317,In_25,N_8);
or U318 (N_318,In_337,N_101);
or U319 (N_319,In_233,N_186);
and U320 (N_320,In_420,N_109);
xnor U321 (N_321,N_149,N_1);
or U322 (N_322,In_335,In_287);
nor U323 (N_323,N_35,In_91);
and U324 (N_324,In_336,In_493);
and U325 (N_325,In_332,N_197);
nor U326 (N_326,N_0,In_379);
and U327 (N_327,N_32,N_64);
nand U328 (N_328,In_40,N_184);
nand U329 (N_329,In_376,N_79);
nand U330 (N_330,N_182,N_61);
nand U331 (N_331,N_50,N_82);
or U332 (N_332,In_13,In_51);
and U333 (N_333,N_57,In_458);
xor U334 (N_334,N_161,N_90);
or U335 (N_335,In_179,N_164);
or U336 (N_336,N_131,N_72);
nand U337 (N_337,N_126,N_128);
nand U338 (N_338,N_166,N_193);
or U339 (N_339,In_220,In_44);
nor U340 (N_340,N_66,N_159);
and U341 (N_341,N_183,N_54);
and U342 (N_342,N_163,N_40);
and U343 (N_343,In_186,In_31);
or U344 (N_344,In_58,N_38);
xor U345 (N_345,N_42,N_178);
nand U346 (N_346,N_192,In_61);
nand U347 (N_347,N_134,N_121);
nor U348 (N_348,N_185,N_135);
and U349 (N_349,N_100,N_52);
or U350 (N_350,N_100,In_46);
and U351 (N_351,N_165,In_458);
or U352 (N_352,N_36,In_160);
nand U353 (N_353,N_84,N_143);
and U354 (N_354,N_146,N_67);
or U355 (N_355,N_120,In_480);
or U356 (N_356,N_32,N_175);
nor U357 (N_357,In_472,N_141);
nand U358 (N_358,In_197,In_208);
nand U359 (N_359,N_76,N_116);
xnor U360 (N_360,In_335,N_121);
nor U361 (N_361,N_38,N_61);
and U362 (N_362,N_23,N_85);
nand U363 (N_363,N_34,N_184);
nor U364 (N_364,N_42,In_186);
nor U365 (N_365,N_97,N_45);
nor U366 (N_366,In_19,N_166);
and U367 (N_367,N_152,N_18);
or U368 (N_368,N_15,N_199);
nor U369 (N_369,N_59,N_97);
nand U370 (N_370,In_318,In_295);
nor U371 (N_371,N_99,N_30);
nor U372 (N_372,N_70,N_19);
nor U373 (N_373,N_149,N_155);
and U374 (N_374,N_52,In_183);
nand U375 (N_375,In_181,N_43);
and U376 (N_376,N_25,In_242);
nand U377 (N_377,In_220,In_197);
nor U378 (N_378,N_74,N_178);
or U379 (N_379,In_480,N_21);
and U380 (N_380,N_123,In_245);
or U381 (N_381,In_95,In_420);
nand U382 (N_382,N_121,N_49);
or U383 (N_383,In_186,N_95);
nor U384 (N_384,In_217,N_135);
nand U385 (N_385,N_62,N_28);
nand U386 (N_386,N_8,N_68);
or U387 (N_387,N_70,In_453);
nand U388 (N_388,N_77,N_175);
or U389 (N_389,In_327,N_184);
or U390 (N_390,N_24,In_472);
nand U391 (N_391,N_116,N_139);
nand U392 (N_392,N_53,N_31);
nand U393 (N_393,N_135,N_84);
or U394 (N_394,N_164,In_183);
nor U395 (N_395,N_34,N_53);
nor U396 (N_396,N_70,In_179);
or U397 (N_397,N_74,N_86);
nand U398 (N_398,N_193,N_64);
xor U399 (N_399,In_337,N_11);
nor U400 (N_400,N_392,N_316);
or U401 (N_401,N_232,N_346);
nand U402 (N_402,N_317,N_321);
and U403 (N_403,N_347,N_333);
or U404 (N_404,N_214,N_255);
or U405 (N_405,N_258,N_216);
nand U406 (N_406,N_228,N_261);
or U407 (N_407,N_269,N_301);
or U408 (N_408,N_324,N_229);
and U409 (N_409,N_376,N_221);
nand U410 (N_410,N_274,N_318);
nor U411 (N_411,N_243,N_254);
and U412 (N_412,N_302,N_234);
and U413 (N_413,N_357,N_391);
or U414 (N_414,N_387,N_287);
or U415 (N_415,N_215,N_390);
or U416 (N_416,N_297,N_209);
nand U417 (N_417,N_275,N_311);
nand U418 (N_418,N_354,N_252);
nor U419 (N_419,N_265,N_383);
nor U420 (N_420,N_338,N_398);
and U421 (N_421,N_378,N_325);
nor U422 (N_422,N_217,N_204);
nand U423 (N_423,N_304,N_223);
nand U424 (N_424,N_277,N_386);
nand U425 (N_425,N_271,N_279);
or U426 (N_426,N_245,N_349);
and U427 (N_427,N_353,N_374);
and U428 (N_428,N_247,N_388);
and U429 (N_429,N_328,N_300);
and U430 (N_430,N_267,N_283);
nor U431 (N_431,N_241,N_239);
or U432 (N_432,N_259,N_322);
nor U433 (N_433,N_291,N_264);
nand U434 (N_434,N_394,N_364);
and U435 (N_435,N_395,N_377);
xnor U436 (N_436,N_230,N_385);
nor U437 (N_437,N_224,N_396);
and U438 (N_438,N_220,N_244);
xnor U439 (N_439,N_315,N_352);
or U440 (N_440,N_335,N_235);
nand U441 (N_441,N_358,N_238);
and U442 (N_442,N_226,N_249);
nand U443 (N_443,N_266,N_337);
and U444 (N_444,N_257,N_336);
xnor U445 (N_445,N_272,N_202);
or U446 (N_446,N_281,N_280);
nor U447 (N_447,N_231,N_295);
or U448 (N_448,N_366,N_323);
nor U449 (N_449,N_360,N_330);
nand U450 (N_450,N_299,N_222);
xnor U451 (N_451,N_286,N_240);
or U452 (N_452,N_298,N_310);
nand U453 (N_453,N_368,N_227);
nor U454 (N_454,N_359,N_290);
or U455 (N_455,N_305,N_250);
nor U456 (N_456,N_268,N_344);
nand U457 (N_457,N_362,N_242);
nor U458 (N_458,N_262,N_367);
or U459 (N_459,N_276,N_375);
or U460 (N_460,N_350,N_251);
and U461 (N_461,N_208,N_289);
and U462 (N_462,N_319,N_273);
nor U463 (N_463,N_236,N_293);
nor U464 (N_464,N_203,N_329);
or U465 (N_465,N_294,N_397);
nor U466 (N_466,N_314,N_369);
nand U467 (N_467,N_355,N_356);
nor U468 (N_468,N_211,N_206);
xor U469 (N_469,N_343,N_399);
or U470 (N_470,N_341,N_373);
xnor U471 (N_471,N_308,N_246);
nor U472 (N_472,N_263,N_312);
nor U473 (N_473,N_361,N_292);
and U474 (N_474,N_309,N_389);
nor U475 (N_475,N_288,N_379);
nor U476 (N_476,N_320,N_307);
nand U477 (N_477,N_348,N_225);
nor U478 (N_478,N_331,N_253);
and U479 (N_479,N_339,N_218);
or U480 (N_480,N_363,N_207);
nor U481 (N_481,N_284,N_210);
or U482 (N_482,N_332,N_200);
and U483 (N_483,N_237,N_365);
nor U484 (N_484,N_248,N_256);
nand U485 (N_485,N_282,N_340);
or U486 (N_486,N_372,N_201);
or U487 (N_487,N_303,N_260);
nand U488 (N_488,N_306,N_213);
nor U489 (N_489,N_393,N_380);
and U490 (N_490,N_381,N_326);
or U491 (N_491,N_334,N_345);
and U492 (N_492,N_278,N_327);
nand U493 (N_493,N_342,N_285);
or U494 (N_494,N_270,N_371);
xor U495 (N_495,N_370,N_313);
nand U496 (N_496,N_205,N_351);
xor U497 (N_497,N_212,N_296);
xnor U498 (N_498,N_382,N_219);
nor U499 (N_499,N_384,N_233);
nand U500 (N_500,N_235,N_228);
xnor U501 (N_501,N_286,N_275);
or U502 (N_502,N_231,N_230);
nand U503 (N_503,N_306,N_308);
xor U504 (N_504,N_206,N_224);
or U505 (N_505,N_334,N_206);
or U506 (N_506,N_383,N_335);
and U507 (N_507,N_313,N_220);
nor U508 (N_508,N_397,N_228);
nand U509 (N_509,N_216,N_233);
xor U510 (N_510,N_394,N_233);
and U511 (N_511,N_297,N_353);
and U512 (N_512,N_397,N_280);
nor U513 (N_513,N_244,N_300);
nor U514 (N_514,N_334,N_259);
xor U515 (N_515,N_252,N_283);
xor U516 (N_516,N_344,N_221);
or U517 (N_517,N_346,N_358);
nor U518 (N_518,N_383,N_280);
and U519 (N_519,N_336,N_329);
nor U520 (N_520,N_332,N_389);
nor U521 (N_521,N_303,N_242);
and U522 (N_522,N_331,N_257);
or U523 (N_523,N_370,N_379);
or U524 (N_524,N_286,N_393);
xnor U525 (N_525,N_250,N_301);
nand U526 (N_526,N_357,N_390);
and U527 (N_527,N_212,N_342);
or U528 (N_528,N_216,N_396);
or U529 (N_529,N_216,N_361);
nand U530 (N_530,N_356,N_376);
nand U531 (N_531,N_327,N_218);
or U532 (N_532,N_301,N_288);
and U533 (N_533,N_335,N_202);
nor U534 (N_534,N_231,N_285);
xor U535 (N_535,N_367,N_303);
nand U536 (N_536,N_334,N_366);
nand U537 (N_537,N_256,N_221);
nor U538 (N_538,N_295,N_206);
and U539 (N_539,N_304,N_366);
nor U540 (N_540,N_278,N_293);
and U541 (N_541,N_259,N_317);
and U542 (N_542,N_349,N_279);
or U543 (N_543,N_342,N_203);
xnor U544 (N_544,N_273,N_350);
nand U545 (N_545,N_369,N_289);
nor U546 (N_546,N_389,N_293);
nand U547 (N_547,N_372,N_224);
or U548 (N_548,N_315,N_293);
xor U549 (N_549,N_306,N_283);
or U550 (N_550,N_366,N_226);
nor U551 (N_551,N_277,N_354);
and U552 (N_552,N_280,N_337);
nand U553 (N_553,N_351,N_326);
or U554 (N_554,N_347,N_299);
and U555 (N_555,N_398,N_367);
or U556 (N_556,N_269,N_236);
xnor U557 (N_557,N_340,N_300);
nor U558 (N_558,N_241,N_276);
or U559 (N_559,N_222,N_210);
nand U560 (N_560,N_275,N_289);
or U561 (N_561,N_396,N_291);
and U562 (N_562,N_257,N_386);
nor U563 (N_563,N_335,N_284);
or U564 (N_564,N_321,N_369);
or U565 (N_565,N_310,N_252);
or U566 (N_566,N_229,N_228);
nor U567 (N_567,N_316,N_332);
and U568 (N_568,N_371,N_374);
and U569 (N_569,N_308,N_309);
and U570 (N_570,N_346,N_215);
nand U571 (N_571,N_333,N_382);
nor U572 (N_572,N_337,N_352);
or U573 (N_573,N_384,N_275);
or U574 (N_574,N_332,N_269);
xor U575 (N_575,N_218,N_232);
and U576 (N_576,N_235,N_327);
nand U577 (N_577,N_283,N_222);
xnor U578 (N_578,N_395,N_310);
nor U579 (N_579,N_212,N_233);
nand U580 (N_580,N_225,N_258);
xnor U581 (N_581,N_201,N_309);
nor U582 (N_582,N_359,N_334);
xor U583 (N_583,N_311,N_203);
nor U584 (N_584,N_298,N_233);
nand U585 (N_585,N_385,N_294);
nand U586 (N_586,N_371,N_335);
or U587 (N_587,N_279,N_382);
and U588 (N_588,N_223,N_370);
or U589 (N_589,N_203,N_276);
or U590 (N_590,N_299,N_219);
nand U591 (N_591,N_208,N_384);
and U592 (N_592,N_376,N_399);
or U593 (N_593,N_321,N_287);
nor U594 (N_594,N_272,N_350);
nor U595 (N_595,N_393,N_261);
nor U596 (N_596,N_252,N_309);
nor U597 (N_597,N_328,N_399);
xnor U598 (N_598,N_319,N_341);
and U599 (N_599,N_295,N_245);
xnor U600 (N_600,N_522,N_541);
or U601 (N_601,N_478,N_416);
nand U602 (N_602,N_509,N_427);
or U603 (N_603,N_533,N_549);
or U604 (N_604,N_513,N_546);
nand U605 (N_605,N_531,N_449);
and U606 (N_606,N_443,N_410);
nor U607 (N_607,N_464,N_406);
and U608 (N_608,N_479,N_588);
nor U609 (N_609,N_581,N_493);
and U610 (N_610,N_508,N_448);
nor U611 (N_611,N_466,N_554);
nand U612 (N_612,N_439,N_413);
or U613 (N_613,N_419,N_552);
and U614 (N_614,N_545,N_491);
nand U615 (N_615,N_441,N_593);
and U616 (N_616,N_584,N_572);
or U617 (N_617,N_409,N_577);
and U618 (N_618,N_511,N_418);
and U619 (N_619,N_518,N_526);
xor U620 (N_620,N_598,N_415);
nand U621 (N_621,N_405,N_411);
nand U622 (N_622,N_542,N_543);
xnor U623 (N_623,N_467,N_477);
and U624 (N_624,N_459,N_507);
and U625 (N_625,N_517,N_489);
or U626 (N_626,N_426,N_597);
and U627 (N_627,N_504,N_514);
xnor U628 (N_628,N_521,N_516);
xnor U629 (N_629,N_553,N_428);
and U630 (N_630,N_456,N_472);
nor U631 (N_631,N_569,N_515);
nand U632 (N_632,N_571,N_412);
or U633 (N_633,N_529,N_500);
xnor U634 (N_634,N_583,N_566);
or U635 (N_635,N_403,N_595);
or U636 (N_636,N_570,N_442);
and U637 (N_637,N_528,N_422);
and U638 (N_638,N_447,N_591);
nand U639 (N_639,N_495,N_524);
or U640 (N_640,N_460,N_436);
or U641 (N_641,N_505,N_401);
or U642 (N_642,N_590,N_594);
nand U643 (N_643,N_487,N_499);
nor U644 (N_644,N_455,N_434);
or U645 (N_645,N_475,N_417);
and U646 (N_646,N_537,N_488);
nand U647 (N_647,N_574,N_432);
nor U648 (N_648,N_462,N_471);
nand U649 (N_649,N_536,N_437);
xor U650 (N_650,N_481,N_433);
nor U651 (N_651,N_527,N_497);
nor U652 (N_652,N_438,N_453);
nor U653 (N_653,N_450,N_586);
and U654 (N_654,N_454,N_476);
or U655 (N_655,N_496,N_452);
nand U656 (N_656,N_544,N_540);
nand U657 (N_657,N_430,N_402);
or U658 (N_658,N_482,N_525);
nand U659 (N_659,N_589,N_538);
and U660 (N_660,N_469,N_400);
and U661 (N_661,N_473,N_444);
nor U662 (N_662,N_520,N_480);
xor U663 (N_663,N_492,N_461);
and U664 (N_664,N_532,N_458);
and U665 (N_665,N_568,N_558);
xnor U666 (N_666,N_451,N_424);
and U667 (N_667,N_502,N_494);
nor U668 (N_668,N_567,N_557);
nor U669 (N_669,N_440,N_408);
or U670 (N_670,N_592,N_523);
nand U671 (N_671,N_535,N_548);
or U672 (N_672,N_539,N_551);
xnor U673 (N_673,N_575,N_599);
xnor U674 (N_674,N_431,N_573);
or U675 (N_675,N_423,N_420);
or U676 (N_676,N_582,N_446);
xor U677 (N_677,N_506,N_519);
xnor U678 (N_678,N_404,N_407);
and U679 (N_679,N_486,N_445);
nand U680 (N_680,N_435,N_587);
and U681 (N_681,N_425,N_562);
or U682 (N_682,N_560,N_564);
or U683 (N_683,N_547,N_484);
or U684 (N_684,N_421,N_465);
or U685 (N_685,N_498,N_510);
nand U686 (N_686,N_585,N_474);
and U687 (N_687,N_512,N_565);
or U688 (N_688,N_468,N_463);
and U689 (N_689,N_503,N_563);
or U690 (N_690,N_559,N_470);
or U691 (N_691,N_576,N_483);
nand U692 (N_692,N_457,N_555);
or U693 (N_693,N_579,N_429);
and U694 (N_694,N_530,N_580);
nor U695 (N_695,N_556,N_501);
or U696 (N_696,N_578,N_596);
or U697 (N_697,N_534,N_485);
or U698 (N_698,N_550,N_490);
and U699 (N_699,N_414,N_561);
or U700 (N_700,N_519,N_578);
and U701 (N_701,N_590,N_449);
and U702 (N_702,N_494,N_480);
and U703 (N_703,N_538,N_484);
and U704 (N_704,N_538,N_403);
or U705 (N_705,N_554,N_402);
or U706 (N_706,N_580,N_460);
and U707 (N_707,N_508,N_413);
nor U708 (N_708,N_417,N_496);
and U709 (N_709,N_424,N_597);
and U710 (N_710,N_473,N_461);
nor U711 (N_711,N_433,N_474);
and U712 (N_712,N_477,N_422);
nand U713 (N_713,N_576,N_584);
xor U714 (N_714,N_482,N_454);
and U715 (N_715,N_456,N_478);
and U716 (N_716,N_537,N_405);
and U717 (N_717,N_432,N_578);
and U718 (N_718,N_471,N_433);
or U719 (N_719,N_519,N_437);
nand U720 (N_720,N_466,N_582);
nor U721 (N_721,N_470,N_427);
and U722 (N_722,N_584,N_416);
and U723 (N_723,N_537,N_492);
nor U724 (N_724,N_523,N_565);
nor U725 (N_725,N_568,N_511);
and U726 (N_726,N_568,N_493);
nand U727 (N_727,N_536,N_468);
nor U728 (N_728,N_587,N_483);
or U729 (N_729,N_475,N_568);
nor U730 (N_730,N_477,N_400);
nor U731 (N_731,N_558,N_482);
or U732 (N_732,N_417,N_572);
nor U733 (N_733,N_494,N_560);
or U734 (N_734,N_490,N_450);
or U735 (N_735,N_554,N_421);
xor U736 (N_736,N_524,N_402);
nor U737 (N_737,N_571,N_525);
and U738 (N_738,N_555,N_535);
nand U739 (N_739,N_513,N_403);
nand U740 (N_740,N_414,N_465);
and U741 (N_741,N_540,N_530);
nor U742 (N_742,N_462,N_426);
or U743 (N_743,N_530,N_546);
nor U744 (N_744,N_456,N_448);
or U745 (N_745,N_443,N_551);
or U746 (N_746,N_429,N_545);
or U747 (N_747,N_595,N_511);
nand U748 (N_748,N_571,N_447);
and U749 (N_749,N_456,N_470);
nand U750 (N_750,N_514,N_453);
or U751 (N_751,N_458,N_557);
and U752 (N_752,N_517,N_523);
nor U753 (N_753,N_587,N_416);
and U754 (N_754,N_572,N_548);
and U755 (N_755,N_489,N_433);
nor U756 (N_756,N_540,N_579);
nor U757 (N_757,N_473,N_459);
and U758 (N_758,N_489,N_544);
nand U759 (N_759,N_463,N_577);
nand U760 (N_760,N_576,N_595);
nand U761 (N_761,N_505,N_502);
or U762 (N_762,N_489,N_422);
or U763 (N_763,N_433,N_522);
and U764 (N_764,N_418,N_579);
xnor U765 (N_765,N_481,N_465);
nor U766 (N_766,N_584,N_445);
xnor U767 (N_767,N_594,N_438);
nand U768 (N_768,N_466,N_542);
xor U769 (N_769,N_516,N_478);
nor U770 (N_770,N_414,N_536);
and U771 (N_771,N_510,N_551);
xnor U772 (N_772,N_564,N_519);
or U773 (N_773,N_410,N_574);
and U774 (N_774,N_558,N_446);
or U775 (N_775,N_454,N_427);
and U776 (N_776,N_432,N_547);
or U777 (N_777,N_550,N_589);
nor U778 (N_778,N_587,N_418);
or U779 (N_779,N_573,N_596);
or U780 (N_780,N_558,N_407);
nand U781 (N_781,N_566,N_424);
nor U782 (N_782,N_436,N_413);
nand U783 (N_783,N_499,N_461);
and U784 (N_784,N_428,N_573);
or U785 (N_785,N_412,N_574);
or U786 (N_786,N_489,N_594);
nand U787 (N_787,N_538,N_508);
or U788 (N_788,N_496,N_454);
and U789 (N_789,N_594,N_457);
nor U790 (N_790,N_567,N_464);
nor U791 (N_791,N_447,N_542);
and U792 (N_792,N_400,N_415);
xnor U793 (N_793,N_565,N_415);
nand U794 (N_794,N_463,N_512);
and U795 (N_795,N_416,N_545);
nor U796 (N_796,N_466,N_568);
xor U797 (N_797,N_456,N_461);
and U798 (N_798,N_521,N_483);
nor U799 (N_799,N_426,N_528);
nor U800 (N_800,N_700,N_604);
or U801 (N_801,N_785,N_663);
nor U802 (N_802,N_646,N_668);
nand U803 (N_803,N_774,N_671);
nand U804 (N_804,N_740,N_795);
nor U805 (N_805,N_623,N_702);
and U806 (N_806,N_756,N_788);
and U807 (N_807,N_735,N_699);
nor U808 (N_808,N_741,N_679);
or U809 (N_809,N_636,N_796);
xor U810 (N_810,N_747,N_710);
xnor U811 (N_811,N_658,N_790);
and U812 (N_812,N_654,N_778);
nor U813 (N_813,N_752,N_672);
or U814 (N_814,N_733,N_789);
xor U815 (N_815,N_688,N_734);
nand U816 (N_816,N_727,N_686);
or U817 (N_817,N_715,N_664);
xor U818 (N_818,N_690,N_632);
nand U819 (N_819,N_609,N_704);
xor U820 (N_820,N_651,N_626);
nor U821 (N_821,N_726,N_683);
nor U822 (N_822,N_713,N_798);
nand U823 (N_823,N_607,N_717);
and U824 (N_824,N_770,N_766);
nor U825 (N_825,N_714,N_708);
nor U826 (N_826,N_744,N_682);
nor U827 (N_827,N_701,N_603);
nor U828 (N_828,N_753,N_638);
and U829 (N_829,N_653,N_670);
or U830 (N_830,N_760,N_655);
or U831 (N_831,N_650,N_724);
nand U832 (N_832,N_678,N_755);
nand U833 (N_833,N_685,N_611);
xor U834 (N_834,N_660,N_773);
xor U835 (N_835,N_792,N_705);
nor U836 (N_836,N_703,N_782);
nor U837 (N_837,N_754,N_677);
and U838 (N_838,N_693,N_739);
and U839 (N_839,N_698,N_648);
nor U840 (N_840,N_743,N_649);
nand U841 (N_841,N_721,N_736);
xnor U842 (N_842,N_723,N_681);
and U843 (N_843,N_634,N_657);
nand U844 (N_844,N_745,N_794);
or U845 (N_845,N_777,N_627);
and U846 (N_846,N_628,N_771);
or U847 (N_847,N_605,N_709);
and U848 (N_848,N_775,N_706);
nand U849 (N_849,N_793,N_711);
or U850 (N_850,N_748,N_621);
xor U851 (N_851,N_641,N_761);
nor U852 (N_852,N_791,N_661);
xor U853 (N_853,N_637,N_662);
and U854 (N_854,N_624,N_780);
or U855 (N_855,N_784,N_783);
nand U856 (N_856,N_767,N_676);
nand U857 (N_857,N_787,N_797);
nor U858 (N_858,N_722,N_692);
or U859 (N_859,N_675,N_749);
xnor U860 (N_860,N_613,N_799);
and U861 (N_861,N_635,N_718);
or U862 (N_862,N_725,N_751);
xor U863 (N_863,N_757,N_696);
or U864 (N_864,N_625,N_615);
nand U865 (N_865,N_732,N_776);
nor U866 (N_866,N_630,N_786);
nor U867 (N_867,N_762,N_758);
or U868 (N_868,N_765,N_644);
and U869 (N_869,N_695,N_645);
nor U870 (N_870,N_729,N_608);
or U871 (N_871,N_667,N_694);
nand U872 (N_872,N_666,N_652);
or U873 (N_873,N_669,N_687);
and U874 (N_874,N_622,N_712);
or U875 (N_875,N_716,N_659);
nor U876 (N_876,N_781,N_737);
or U877 (N_877,N_738,N_689);
and U878 (N_878,N_731,N_763);
nor U879 (N_879,N_759,N_633);
or U880 (N_880,N_742,N_750);
or U881 (N_881,N_647,N_720);
or U882 (N_882,N_618,N_779);
or U883 (N_883,N_610,N_772);
nor U884 (N_884,N_606,N_665);
and U885 (N_885,N_697,N_612);
or U886 (N_886,N_768,N_746);
or U887 (N_887,N_601,N_769);
nor U888 (N_888,N_719,N_600);
nor U889 (N_889,N_674,N_640);
xnor U890 (N_890,N_642,N_629);
xor U891 (N_891,N_691,N_643);
nor U892 (N_892,N_764,N_631);
nor U893 (N_893,N_730,N_673);
or U894 (N_894,N_614,N_619);
nand U895 (N_895,N_707,N_620);
nor U896 (N_896,N_639,N_602);
nor U897 (N_897,N_684,N_617);
and U898 (N_898,N_728,N_616);
nand U899 (N_899,N_656,N_680);
nor U900 (N_900,N_699,N_713);
and U901 (N_901,N_709,N_653);
and U902 (N_902,N_640,N_688);
nand U903 (N_903,N_683,N_737);
nand U904 (N_904,N_672,N_667);
nand U905 (N_905,N_742,N_746);
or U906 (N_906,N_757,N_694);
and U907 (N_907,N_668,N_688);
and U908 (N_908,N_652,N_667);
and U909 (N_909,N_756,N_725);
and U910 (N_910,N_639,N_784);
or U911 (N_911,N_774,N_673);
or U912 (N_912,N_764,N_789);
and U913 (N_913,N_780,N_741);
nand U914 (N_914,N_665,N_667);
or U915 (N_915,N_646,N_715);
nand U916 (N_916,N_676,N_759);
nand U917 (N_917,N_736,N_694);
or U918 (N_918,N_605,N_632);
or U919 (N_919,N_670,N_769);
and U920 (N_920,N_628,N_768);
nor U921 (N_921,N_724,N_771);
or U922 (N_922,N_797,N_647);
or U923 (N_923,N_678,N_726);
xor U924 (N_924,N_633,N_783);
and U925 (N_925,N_662,N_744);
nand U926 (N_926,N_697,N_668);
nand U927 (N_927,N_621,N_676);
nor U928 (N_928,N_618,N_605);
nor U929 (N_929,N_674,N_637);
xor U930 (N_930,N_791,N_749);
xor U931 (N_931,N_752,N_772);
and U932 (N_932,N_698,N_758);
nand U933 (N_933,N_741,N_733);
xor U934 (N_934,N_665,N_647);
nand U935 (N_935,N_613,N_647);
nor U936 (N_936,N_717,N_639);
and U937 (N_937,N_642,N_679);
or U938 (N_938,N_609,N_714);
nand U939 (N_939,N_702,N_723);
nor U940 (N_940,N_692,N_749);
and U941 (N_941,N_631,N_630);
or U942 (N_942,N_684,N_764);
and U943 (N_943,N_680,N_658);
xor U944 (N_944,N_670,N_606);
nand U945 (N_945,N_675,N_787);
xnor U946 (N_946,N_733,N_604);
nand U947 (N_947,N_797,N_719);
and U948 (N_948,N_761,N_663);
nor U949 (N_949,N_799,N_740);
and U950 (N_950,N_641,N_798);
nand U951 (N_951,N_745,N_779);
and U952 (N_952,N_798,N_744);
nand U953 (N_953,N_728,N_719);
nand U954 (N_954,N_741,N_621);
nand U955 (N_955,N_796,N_786);
xnor U956 (N_956,N_661,N_781);
and U957 (N_957,N_775,N_602);
nand U958 (N_958,N_760,N_649);
nand U959 (N_959,N_768,N_648);
nor U960 (N_960,N_799,N_712);
nor U961 (N_961,N_791,N_780);
or U962 (N_962,N_729,N_751);
nor U963 (N_963,N_769,N_771);
nor U964 (N_964,N_759,N_621);
nand U965 (N_965,N_683,N_612);
or U966 (N_966,N_764,N_639);
nand U967 (N_967,N_662,N_601);
and U968 (N_968,N_776,N_632);
nand U969 (N_969,N_733,N_715);
nand U970 (N_970,N_765,N_631);
or U971 (N_971,N_705,N_608);
or U972 (N_972,N_716,N_751);
nor U973 (N_973,N_614,N_719);
and U974 (N_974,N_601,N_610);
and U975 (N_975,N_637,N_750);
nand U976 (N_976,N_713,N_706);
or U977 (N_977,N_626,N_722);
nor U978 (N_978,N_676,N_784);
xnor U979 (N_979,N_789,N_799);
xnor U980 (N_980,N_745,N_780);
or U981 (N_981,N_640,N_629);
and U982 (N_982,N_775,N_790);
nand U983 (N_983,N_638,N_657);
nor U984 (N_984,N_641,N_742);
nor U985 (N_985,N_646,N_630);
or U986 (N_986,N_716,N_752);
or U987 (N_987,N_778,N_727);
and U988 (N_988,N_727,N_647);
xnor U989 (N_989,N_697,N_706);
or U990 (N_990,N_744,N_710);
xnor U991 (N_991,N_609,N_710);
nor U992 (N_992,N_641,N_697);
xor U993 (N_993,N_676,N_712);
nand U994 (N_994,N_658,N_647);
nor U995 (N_995,N_743,N_696);
nor U996 (N_996,N_688,N_768);
nand U997 (N_997,N_761,N_783);
nor U998 (N_998,N_636,N_706);
nand U999 (N_999,N_788,N_660);
nor U1000 (N_1000,N_892,N_987);
and U1001 (N_1001,N_848,N_884);
xnor U1002 (N_1002,N_973,N_971);
nor U1003 (N_1003,N_843,N_916);
nand U1004 (N_1004,N_890,N_812);
nand U1005 (N_1005,N_970,N_867);
nor U1006 (N_1006,N_962,N_938);
nand U1007 (N_1007,N_830,N_908);
or U1008 (N_1008,N_968,N_839);
nand U1009 (N_1009,N_826,N_868);
nor U1010 (N_1010,N_978,N_917);
and U1011 (N_1011,N_947,N_915);
xor U1012 (N_1012,N_899,N_929);
nand U1013 (N_1013,N_952,N_911);
or U1014 (N_1014,N_896,N_931);
nor U1015 (N_1015,N_967,N_894);
and U1016 (N_1016,N_838,N_898);
or U1017 (N_1017,N_945,N_999);
and U1018 (N_1018,N_893,N_831);
and U1019 (N_1019,N_974,N_849);
and U1020 (N_1020,N_914,N_981);
nand U1021 (N_1021,N_804,N_948);
xor U1022 (N_1022,N_811,N_821);
and U1023 (N_1023,N_888,N_877);
or U1024 (N_1024,N_958,N_913);
or U1025 (N_1025,N_969,N_886);
nand U1026 (N_1026,N_875,N_858);
nor U1027 (N_1027,N_901,N_840);
nor U1028 (N_1028,N_865,N_955);
nand U1029 (N_1029,N_975,N_926);
nand U1030 (N_1030,N_942,N_961);
xor U1031 (N_1031,N_927,N_869);
xnor U1032 (N_1032,N_957,N_936);
or U1033 (N_1033,N_860,N_944);
nand U1034 (N_1034,N_977,N_979);
nor U1035 (N_1035,N_910,N_963);
and U1036 (N_1036,N_930,N_994);
nor U1037 (N_1037,N_984,N_923);
and U1038 (N_1038,N_976,N_940);
and U1039 (N_1039,N_881,N_924);
nand U1040 (N_1040,N_998,N_837);
nand U1041 (N_1041,N_925,N_906);
nand U1042 (N_1042,N_835,N_847);
nand U1043 (N_1043,N_982,N_902);
and U1044 (N_1044,N_833,N_941);
xor U1045 (N_1045,N_820,N_841);
nor U1046 (N_1046,N_949,N_856);
or U1047 (N_1047,N_922,N_806);
and U1048 (N_1048,N_934,N_828);
or U1049 (N_1049,N_844,N_939);
nand U1050 (N_1050,N_862,N_943);
xnor U1051 (N_1051,N_907,N_817);
nand U1052 (N_1052,N_953,N_960);
nor U1053 (N_1053,N_813,N_964);
or U1054 (N_1054,N_905,N_951);
nand U1055 (N_1055,N_803,N_861);
or U1056 (N_1056,N_823,N_810);
nor U1057 (N_1057,N_864,N_990);
or U1058 (N_1058,N_985,N_956);
xnor U1059 (N_1059,N_850,N_991);
nand U1060 (N_1060,N_874,N_816);
and U1061 (N_1061,N_887,N_895);
and U1062 (N_1062,N_972,N_808);
nand U1063 (N_1063,N_801,N_937);
nor U1064 (N_1064,N_883,N_824);
and U1065 (N_1065,N_919,N_845);
nand U1066 (N_1066,N_891,N_912);
or U1067 (N_1067,N_903,N_854);
and U1068 (N_1068,N_851,N_954);
nand U1069 (N_1069,N_880,N_871);
or U1070 (N_1070,N_989,N_983);
nand U1071 (N_1071,N_863,N_993);
and U1072 (N_1072,N_921,N_873);
and U1073 (N_1073,N_885,N_897);
nor U1074 (N_1074,N_932,N_819);
and U1075 (N_1075,N_827,N_870);
and U1076 (N_1076,N_805,N_855);
nand U1077 (N_1077,N_852,N_857);
xnor U1078 (N_1078,N_900,N_814);
xnor U1079 (N_1079,N_904,N_822);
nor U1080 (N_1080,N_997,N_966);
or U1081 (N_1081,N_882,N_872);
nor U1082 (N_1082,N_818,N_800);
and U1083 (N_1083,N_933,N_866);
and U1084 (N_1084,N_959,N_988);
and U1085 (N_1085,N_825,N_807);
nor U1086 (N_1086,N_878,N_834);
or U1087 (N_1087,N_928,N_829);
xnor U1088 (N_1088,N_859,N_909);
nor U1089 (N_1089,N_889,N_876);
or U1090 (N_1090,N_832,N_815);
nand U1091 (N_1091,N_853,N_965);
xor U1092 (N_1092,N_809,N_986);
and U1093 (N_1093,N_992,N_842);
nor U1094 (N_1094,N_879,N_980);
xor U1095 (N_1095,N_946,N_846);
nor U1096 (N_1096,N_802,N_996);
and U1097 (N_1097,N_995,N_935);
or U1098 (N_1098,N_950,N_836);
and U1099 (N_1099,N_918,N_920);
and U1100 (N_1100,N_943,N_944);
nor U1101 (N_1101,N_812,N_884);
nand U1102 (N_1102,N_954,N_943);
and U1103 (N_1103,N_824,N_865);
nand U1104 (N_1104,N_922,N_997);
and U1105 (N_1105,N_836,N_969);
nor U1106 (N_1106,N_821,N_851);
xnor U1107 (N_1107,N_974,N_956);
and U1108 (N_1108,N_984,N_958);
nor U1109 (N_1109,N_908,N_947);
or U1110 (N_1110,N_899,N_861);
and U1111 (N_1111,N_826,N_971);
nand U1112 (N_1112,N_888,N_955);
nand U1113 (N_1113,N_870,N_820);
or U1114 (N_1114,N_853,N_896);
and U1115 (N_1115,N_802,N_810);
and U1116 (N_1116,N_841,N_967);
nor U1117 (N_1117,N_880,N_838);
or U1118 (N_1118,N_853,N_934);
or U1119 (N_1119,N_816,N_803);
or U1120 (N_1120,N_807,N_853);
nand U1121 (N_1121,N_824,N_826);
xnor U1122 (N_1122,N_932,N_856);
or U1123 (N_1123,N_901,N_905);
nand U1124 (N_1124,N_887,N_988);
or U1125 (N_1125,N_915,N_890);
xnor U1126 (N_1126,N_828,N_938);
nand U1127 (N_1127,N_931,N_825);
nand U1128 (N_1128,N_977,N_830);
nor U1129 (N_1129,N_992,N_868);
xor U1130 (N_1130,N_979,N_988);
xnor U1131 (N_1131,N_932,N_813);
nor U1132 (N_1132,N_973,N_995);
nand U1133 (N_1133,N_923,N_800);
xor U1134 (N_1134,N_996,N_863);
or U1135 (N_1135,N_900,N_887);
or U1136 (N_1136,N_882,N_995);
nand U1137 (N_1137,N_826,N_948);
xor U1138 (N_1138,N_989,N_839);
nor U1139 (N_1139,N_800,N_872);
or U1140 (N_1140,N_933,N_851);
and U1141 (N_1141,N_861,N_864);
and U1142 (N_1142,N_939,N_928);
nand U1143 (N_1143,N_819,N_880);
xnor U1144 (N_1144,N_887,N_944);
and U1145 (N_1145,N_869,N_831);
or U1146 (N_1146,N_938,N_813);
nor U1147 (N_1147,N_822,N_821);
nand U1148 (N_1148,N_976,N_972);
nand U1149 (N_1149,N_907,N_968);
xnor U1150 (N_1150,N_937,N_847);
nor U1151 (N_1151,N_870,N_835);
nand U1152 (N_1152,N_814,N_843);
and U1153 (N_1153,N_987,N_967);
nor U1154 (N_1154,N_804,N_924);
xor U1155 (N_1155,N_995,N_947);
or U1156 (N_1156,N_819,N_806);
or U1157 (N_1157,N_829,N_970);
nand U1158 (N_1158,N_852,N_865);
nand U1159 (N_1159,N_984,N_806);
and U1160 (N_1160,N_959,N_812);
and U1161 (N_1161,N_868,N_870);
nor U1162 (N_1162,N_976,N_865);
or U1163 (N_1163,N_887,N_856);
or U1164 (N_1164,N_895,N_973);
and U1165 (N_1165,N_829,N_938);
nand U1166 (N_1166,N_866,N_915);
nand U1167 (N_1167,N_847,N_979);
nand U1168 (N_1168,N_881,N_936);
nand U1169 (N_1169,N_972,N_912);
or U1170 (N_1170,N_904,N_919);
or U1171 (N_1171,N_814,N_866);
or U1172 (N_1172,N_993,N_882);
or U1173 (N_1173,N_991,N_944);
nand U1174 (N_1174,N_821,N_874);
and U1175 (N_1175,N_887,N_935);
or U1176 (N_1176,N_888,N_952);
xor U1177 (N_1177,N_848,N_935);
nand U1178 (N_1178,N_930,N_985);
or U1179 (N_1179,N_913,N_846);
nor U1180 (N_1180,N_841,N_961);
and U1181 (N_1181,N_957,N_830);
or U1182 (N_1182,N_833,N_906);
and U1183 (N_1183,N_880,N_933);
and U1184 (N_1184,N_976,N_876);
nand U1185 (N_1185,N_849,N_859);
xnor U1186 (N_1186,N_931,N_814);
xnor U1187 (N_1187,N_949,N_887);
xnor U1188 (N_1188,N_993,N_881);
or U1189 (N_1189,N_919,N_962);
and U1190 (N_1190,N_805,N_966);
nor U1191 (N_1191,N_883,N_901);
or U1192 (N_1192,N_874,N_922);
nand U1193 (N_1193,N_883,N_861);
and U1194 (N_1194,N_859,N_985);
or U1195 (N_1195,N_896,N_835);
and U1196 (N_1196,N_987,N_883);
nand U1197 (N_1197,N_974,N_896);
nand U1198 (N_1198,N_970,N_932);
nand U1199 (N_1199,N_922,N_883);
nand U1200 (N_1200,N_1123,N_1084);
and U1201 (N_1201,N_1089,N_1037);
and U1202 (N_1202,N_1019,N_1166);
or U1203 (N_1203,N_1119,N_1046);
nand U1204 (N_1204,N_1014,N_1076);
and U1205 (N_1205,N_1000,N_1135);
nor U1206 (N_1206,N_1103,N_1008);
nand U1207 (N_1207,N_1171,N_1177);
nand U1208 (N_1208,N_1102,N_1018);
and U1209 (N_1209,N_1054,N_1043);
nor U1210 (N_1210,N_1130,N_1004);
and U1211 (N_1211,N_1086,N_1170);
xor U1212 (N_1212,N_1028,N_1193);
nand U1213 (N_1213,N_1082,N_1017);
or U1214 (N_1214,N_1021,N_1097);
xnor U1215 (N_1215,N_1080,N_1175);
or U1216 (N_1216,N_1049,N_1173);
nand U1217 (N_1217,N_1184,N_1114);
or U1218 (N_1218,N_1109,N_1144);
xor U1219 (N_1219,N_1006,N_1002);
nand U1220 (N_1220,N_1143,N_1094);
and U1221 (N_1221,N_1067,N_1005);
nor U1222 (N_1222,N_1011,N_1192);
or U1223 (N_1223,N_1156,N_1125);
and U1224 (N_1224,N_1083,N_1085);
or U1225 (N_1225,N_1105,N_1133);
and U1226 (N_1226,N_1035,N_1093);
xor U1227 (N_1227,N_1120,N_1190);
or U1228 (N_1228,N_1064,N_1142);
or U1229 (N_1229,N_1167,N_1196);
or U1230 (N_1230,N_1013,N_1088);
nor U1231 (N_1231,N_1077,N_1039);
xnor U1232 (N_1232,N_1153,N_1110);
or U1233 (N_1233,N_1157,N_1069);
nand U1234 (N_1234,N_1051,N_1195);
xor U1235 (N_1235,N_1141,N_1023);
or U1236 (N_1236,N_1198,N_1068);
or U1237 (N_1237,N_1052,N_1048);
and U1238 (N_1238,N_1118,N_1148);
xnor U1239 (N_1239,N_1010,N_1078);
nor U1240 (N_1240,N_1191,N_1117);
or U1241 (N_1241,N_1159,N_1158);
or U1242 (N_1242,N_1095,N_1022);
nand U1243 (N_1243,N_1180,N_1079);
and U1244 (N_1244,N_1147,N_1182);
nand U1245 (N_1245,N_1003,N_1134);
and U1246 (N_1246,N_1063,N_1070);
nor U1247 (N_1247,N_1194,N_1055);
nand U1248 (N_1248,N_1127,N_1185);
xor U1249 (N_1249,N_1197,N_1174);
nand U1250 (N_1250,N_1031,N_1057);
nand U1251 (N_1251,N_1062,N_1074);
nor U1252 (N_1252,N_1030,N_1199);
xor U1253 (N_1253,N_1045,N_1179);
xnor U1254 (N_1254,N_1016,N_1189);
nand U1255 (N_1255,N_1115,N_1188);
nand U1256 (N_1256,N_1108,N_1100);
nor U1257 (N_1257,N_1160,N_1096);
and U1258 (N_1258,N_1163,N_1146);
nor U1259 (N_1259,N_1101,N_1140);
xor U1260 (N_1260,N_1099,N_1149);
nand U1261 (N_1261,N_1073,N_1027);
or U1262 (N_1262,N_1107,N_1165);
nor U1263 (N_1263,N_1050,N_1026);
nor U1264 (N_1264,N_1169,N_1007);
or U1265 (N_1265,N_1025,N_1187);
nand U1266 (N_1266,N_1111,N_1139);
xnor U1267 (N_1267,N_1042,N_1081);
or U1268 (N_1268,N_1181,N_1058);
and U1269 (N_1269,N_1124,N_1178);
or U1270 (N_1270,N_1155,N_1113);
nor U1271 (N_1271,N_1024,N_1075);
nand U1272 (N_1272,N_1121,N_1092);
nor U1273 (N_1273,N_1009,N_1168);
and U1274 (N_1274,N_1029,N_1065);
nor U1275 (N_1275,N_1090,N_1056);
nor U1276 (N_1276,N_1132,N_1106);
and U1277 (N_1277,N_1128,N_1152);
nand U1278 (N_1278,N_1071,N_1150);
or U1279 (N_1279,N_1034,N_1176);
nor U1280 (N_1280,N_1164,N_1116);
nor U1281 (N_1281,N_1047,N_1126);
nor U1282 (N_1282,N_1066,N_1151);
or U1283 (N_1283,N_1138,N_1131);
or U1284 (N_1284,N_1104,N_1145);
nor U1285 (N_1285,N_1036,N_1015);
nor U1286 (N_1286,N_1183,N_1112);
nand U1287 (N_1287,N_1053,N_1137);
nor U1288 (N_1288,N_1012,N_1162);
or U1289 (N_1289,N_1161,N_1098);
and U1290 (N_1290,N_1038,N_1060);
nand U1291 (N_1291,N_1059,N_1061);
nor U1292 (N_1292,N_1154,N_1136);
and U1293 (N_1293,N_1072,N_1033);
nand U1294 (N_1294,N_1129,N_1172);
and U1295 (N_1295,N_1041,N_1122);
nand U1296 (N_1296,N_1087,N_1032);
and U1297 (N_1297,N_1044,N_1040);
and U1298 (N_1298,N_1091,N_1020);
xnor U1299 (N_1299,N_1186,N_1001);
nand U1300 (N_1300,N_1152,N_1118);
nand U1301 (N_1301,N_1118,N_1056);
nand U1302 (N_1302,N_1010,N_1012);
or U1303 (N_1303,N_1019,N_1060);
nor U1304 (N_1304,N_1183,N_1061);
or U1305 (N_1305,N_1141,N_1031);
nor U1306 (N_1306,N_1052,N_1146);
or U1307 (N_1307,N_1123,N_1090);
nand U1308 (N_1308,N_1031,N_1054);
nand U1309 (N_1309,N_1084,N_1139);
or U1310 (N_1310,N_1070,N_1000);
xor U1311 (N_1311,N_1031,N_1019);
or U1312 (N_1312,N_1102,N_1154);
xnor U1313 (N_1313,N_1115,N_1189);
nor U1314 (N_1314,N_1063,N_1048);
nor U1315 (N_1315,N_1054,N_1182);
nand U1316 (N_1316,N_1009,N_1151);
or U1317 (N_1317,N_1008,N_1182);
nor U1318 (N_1318,N_1003,N_1026);
nor U1319 (N_1319,N_1135,N_1114);
nor U1320 (N_1320,N_1008,N_1164);
and U1321 (N_1321,N_1106,N_1014);
and U1322 (N_1322,N_1126,N_1067);
nand U1323 (N_1323,N_1022,N_1065);
nand U1324 (N_1324,N_1186,N_1072);
xor U1325 (N_1325,N_1166,N_1065);
nor U1326 (N_1326,N_1111,N_1090);
or U1327 (N_1327,N_1079,N_1063);
nand U1328 (N_1328,N_1053,N_1087);
or U1329 (N_1329,N_1040,N_1144);
nor U1330 (N_1330,N_1143,N_1078);
nor U1331 (N_1331,N_1008,N_1067);
and U1332 (N_1332,N_1164,N_1151);
or U1333 (N_1333,N_1048,N_1080);
or U1334 (N_1334,N_1005,N_1004);
xnor U1335 (N_1335,N_1008,N_1135);
nand U1336 (N_1336,N_1071,N_1012);
and U1337 (N_1337,N_1146,N_1033);
nand U1338 (N_1338,N_1189,N_1165);
and U1339 (N_1339,N_1097,N_1056);
and U1340 (N_1340,N_1087,N_1150);
or U1341 (N_1341,N_1193,N_1019);
or U1342 (N_1342,N_1106,N_1031);
or U1343 (N_1343,N_1002,N_1141);
nand U1344 (N_1344,N_1018,N_1183);
nand U1345 (N_1345,N_1178,N_1183);
or U1346 (N_1346,N_1007,N_1140);
or U1347 (N_1347,N_1155,N_1045);
and U1348 (N_1348,N_1123,N_1162);
or U1349 (N_1349,N_1046,N_1135);
nand U1350 (N_1350,N_1188,N_1179);
and U1351 (N_1351,N_1119,N_1091);
nand U1352 (N_1352,N_1144,N_1149);
and U1353 (N_1353,N_1145,N_1117);
xor U1354 (N_1354,N_1062,N_1067);
nand U1355 (N_1355,N_1039,N_1183);
nor U1356 (N_1356,N_1046,N_1036);
or U1357 (N_1357,N_1023,N_1119);
nand U1358 (N_1358,N_1120,N_1077);
xor U1359 (N_1359,N_1108,N_1153);
and U1360 (N_1360,N_1117,N_1171);
or U1361 (N_1361,N_1045,N_1184);
or U1362 (N_1362,N_1092,N_1073);
nor U1363 (N_1363,N_1138,N_1174);
and U1364 (N_1364,N_1077,N_1156);
nand U1365 (N_1365,N_1152,N_1184);
nor U1366 (N_1366,N_1141,N_1119);
and U1367 (N_1367,N_1195,N_1115);
nand U1368 (N_1368,N_1030,N_1071);
nand U1369 (N_1369,N_1057,N_1176);
nand U1370 (N_1370,N_1143,N_1052);
and U1371 (N_1371,N_1033,N_1047);
and U1372 (N_1372,N_1031,N_1104);
and U1373 (N_1373,N_1117,N_1065);
nor U1374 (N_1374,N_1049,N_1194);
or U1375 (N_1375,N_1084,N_1114);
and U1376 (N_1376,N_1067,N_1083);
and U1377 (N_1377,N_1184,N_1053);
or U1378 (N_1378,N_1157,N_1120);
xnor U1379 (N_1379,N_1126,N_1094);
and U1380 (N_1380,N_1184,N_1157);
nand U1381 (N_1381,N_1129,N_1166);
nand U1382 (N_1382,N_1136,N_1179);
xnor U1383 (N_1383,N_1040,N_1096);
nor U1384 (N_1384,N_1109,N_1118);
or U1385 (N_1385,N_1149,N_1148);
nor U1386 (N_1386,N_1137,N_1100);
nand U1387 (N_1387,N_1164,N_1049);
nand U1388 (N_1388,N_1118,N_1025);
nor U1389 (N_1389,N_1186,N_1050);
xor U1390 (N_1390,N_1182,N_1022);
and U1391 (N_1391,N_1105,N_1037);
nor U1392 (N_1392,N_1011,N_1037);
nor U1393 (N_1393,N_1165,N_1028);
nor U1394 (N_1394,N_1017,N_1162);
nand U1395 (N_1395,N_1123,N_1045);
nand U1396 (N_1396,N_1009,N_1048);
nand U1397 (N_1397,N_1165,N_1044);
xor U1398 (N_1398,N_1104,N_1096);
nand U1399 (N_1399,N_1154,N_1021);
nand U1400 (N_1400,N_1249,N_1224);
or U1401 (N_1401,N_1388,N_1328);
nand U1402 (N_1402,N_1392,N_1274);
nor U1403 (N_1403,N_1341,N_1348);
xnor U1404 (N_1404,N_1276,N_1396);
and U1405 (N_1405,N_1266,N_1288);
nor U1406 (N_1406,N_1383,N_1327);
nand U1407 (N_1407,N_1267,N_1311);
and U1408 (N_1408,N_1221,N_1277);
xnor U1409 (N_1409,N_1344,N_1256);
nand U1410 (N_1410,N_1250,N_1360);
nor U1411 (N_1411,N_1232,N_1300);
nand U1412 (N_1412,N_1317,N_1316);
nand U1413 (N_1413,N_1282,N_1320);
nor U1414 (N_1414,N_1314,N_1245);
xnor U1415 (N_1415,N_1270,N_1229);
nor U1416 (N_1416,N_1322,N_1399);
and U1417 (N_1417,N_1375,N_1200);
or U1418 (N_1418,N_1337,N_1319);
xor U1419 (N_1419,N_1389,N_1204);
or U1420 (N_1420,N_1332,N_1269);
nor U1421 (N_1421,N_1377,N_1285);
or U1422 (N_1422,N_1325,N_1299);
nor U1423 (N_1423,N_1238,N_1236);
and U1424 (N_1424,N_1211,N_1247);
and U1425 (N_1425,N_1227,N_1290);
nor U1426 (N_1426,N_1234,N_1380);
and U1427 (N_1427,N_1203,N_1286);
or U1428 (N_1428,N_1202,N_1304);
nand U1429 (N_1429,N_1361,N_1363);
or U1430 (N_1430,N_1350,N_1384);
and U1431 (N_1431,N_1382,N_1297);
nand U1432 (N_1432,N_1346,N_1235);
nand U1433 (N_1433,N_1351,N_1289);
nand U1434 (N_1434,N_1205,N_1394);
and U1435 (N_1435,N_1226,N_1324);
and U1436 (N_1436,N_1349,N_1230);
or U1437 (N_1437,N_1353,N_1217);
nor U1438 (N_1438,N_1241,N_1386);
and U1439 (N_1439,N_1261,N_1268);
nand U1440 (N_1440,N_1362,N_1292);
and U1441 (N_1441,N_1284,N_1264);
nor U1442 (N_1442,N_1242,N_1218);
or U1443 (N_1443,N_1315,N_1215);
nor U1444 (N_1444,N_1368,N_1279);
xnor U1445 (N_1445,N_1259,N_1296);
and U1446 (N_1446,N_1251,N_1335);
or U1447 (N_1447,N_1240,N_1312);
nor U1448 (N_1448,N_1365,N_1381);
xor U1449 (N_1449,N_1228,N_1372);
nor U1450 (N_1450,N_1207,N_1310);
nor U1451 (N_1451,N_1246,N_1379);
and U1452 (N_1452,N_1303,N_1356);
nor U1453 (N_1453,N_1343,N_1201);
or U1454 (N_1454,N_1273,N_1254);
or U1455 (N_1455,N_1301,N_1263);
and U1456 (N_1456,N_1366,N_1244);
or U1457 (N_1457,N_1378,N_1354);
and U1458 (N_1458,N_1252,N_1305);
or U1459 (N_1459,N_1209,N_1222);
nor U1460 (N_1460,N_1339,N_1223);
and U1461 (N_1461,N_1371,N_1345);
nand U1462 (N_1462,N_1253,N_1306);
nand U1463 (N_1463,N_1321,N_1326);
nor U1464 (N_1464,N_1347,N_1287);
xnor U1465 (N_1465,N_1271,N_1364);
and U1466 (N_1466,N_1260,N_1237);
nand U1467 (N_1467,N_1367,N_1342);
and U1468 (N_1468,N_1374,N_1295);
or U1469 (N_1469,N_1313,N_1278);
or U1470 (N_1470,N_1220,N_1291);
and U1471 (N_1471,N_1309,N_1283);
xnor U1472 (N_1472,N_1393,N_1280);
nor U1473 (N_1473,N_1208,N_1231);
or U1474 (N_1474,N_1272,N_1355);
and U1475 (N_1475,N_1357,N_1395);
xor U1476 (N_1476,N_1333,N_1216);
or U1477 (N_1477,N_1262,N_1212);
or U1478 (N_1478,N_1323,N_1206);
nor U1479 (N_1479,N_1308,N_1336);
nand U1480 (N_1480,N_1390,N_1376);
or U1481 (N_1481,N_1298,N_1275);
nand U1482 (N_1482,N_1329,N_1391);
nand U1483 (N_1483,N_1213,N_1330);
nand U1484 (N_1484,N_1331,N_1398);
or U1485 (N_1485,N_1293,N_1239);
or U1486 (N_1486,N_1233,N_1359);
or U1487 (N_1487,N_1302,N_1258);
or U1488 (N_1488,N_1318,N_1294);
and U1489 (N_1489,N_1352,N_1257);
nor U1490 (N_1490,N_1255,N_1334);
nor U1491 (N_1491,N_1210,N_1281);
or U1492 (N_1492,N_1265,N_1338);
nor U1493 (N_1493,N_1358,N_1370);
or U1494 (N_1494,N_1243,N_1397);
nand U1495 (N_1495,N_1385,N_1248);
or U1496 (N_1496,N_1214,N_1307);
and U1497 (N_1497,N_1225,N_1369);
nand U1498 (N_1498,N_1387,N_1340);
or U1499 (N_1499,N_1219,N_1373);
xnor U1500 (N_1500,N_1260,N_1369);
xnor U1501 (N_1501,N_1361,N_1398);
nor U1502 (N_1502,N_1318,N_1295);
xor U1503 (N_1503,N_1204,N_1305);
or U1504 (N_1504,N_1269,N_1352);
nand U1505 (N_1505,N_1242,N_1385);
or U1506 (N_1506,N_1205,N_1354);
or U1507 (N_1507,N_1262,N_1359);
xor U1508 (N_1508,N_1286,N_1280);
or U1509 (N_1509,N_1365,N_1208);
and U1510 (N_1510,N_1300,N_1207);
or U1511 (N_1511,N_1218,N_1270);
and U1512 (N_1512,N_1364,N_1377);
and U1513 (N_1513,N_1365,N_1247);
xnor U1514 (N_1514,N_1257,N_1262);
nor U1515 (N_1515,N_1388,N_1335);
or U1516 (N_1516,N_1293,N_1220);
or U1517 (N_1517,N_1399,N_1299);
nand U1518 (N_1518,N_1301,N_1381);
and U1519 (N_1519,N_1303,N_1204);
and U1520 (N_1520,N_1380,N_1369);
nor U1521 (N_1521,N_1230,N_1220);
nor U1522 (N_1522,N_1304,N_1332);
nor U1523 (N_1523,N_1300,N_1268);
or U1524 (N_1524,N_1219,N_1377);
nor U1525 (N_1525,N_1378,N_1298);
and U1526 (N_1526,N_1302,N_1225);
nor U1527 (N_1527,N_1393,N_1230);
xnor U1528 (N_1528,N_1218,N_1385);
and U1529 (N_1529,N_1290,N_1357);
nand U1530 (N_1530,N_1356,N_1278);
and U1531 (N_1531,N_1290,N_1296);
and U1532 (N_1532,N_1284,N_1218);
nor U1533 (N_1533,N_1310,N_1247);
and U1534 (N_1534,N_1364,N_1320);
nor U1535 (N_1535,N_1367,N_1270);
nand U1536 (N_1536,N_1252,N_1374);
and U1537 (N_1537,N_1255,N_1376);
or U1538 (N_1538,N_1212,N_1244);
nor U1539 (N_1539,N_1384,N_1369);
and U1540 (N_1540,N_1213,N_1231);
and U1541 (N_1541,N_1231,N_1330);
and U1542 (N_1542,N_1320,N_1271);
nor U1543 (N_1543,N_1349,N_1263);
or U1544 (N_1544,N_1394,N_1298);
and U1545 (N_1545,N_1266,N_1386);
xor U1546 (N_1546,N_1265,N_1299);
nor U1547 (N_1547,N_1240,N_1217);
and U1548 (N_1548,N_1334,N_1362);
and U1549 (N_1549,N_1296,N_1306);
or U1550 (N_1550,N_1241,N_1302);
and U1551 (N_1551,N_1215,N_1213);
and U1552 (N_1552,N_1263,N_1363);
or U1553 (N_1553,N_1307,N_1326);
xor U1554 (N_1554,N_1356,N_1248);
nor U1555 (N_1555,N_1234,N_1385);
nor U1556 (N_1556,N_1249,N_1231);
nand U1557 (N_1557,N_1360,N_1254);
nand U1558 (N_1558,N_1374,N_1352);
nor U1559 (N_1559,N_1245,N_1320);
or U1560 (N_1560,N_1395,N_1240);
nand U1561 (N_1561,N_1373,N_1257);
nor U1562 (N_1562,N_1207,N_1315);
nand U1563 (N_1563,N_1204,N_1254);
nor U1564 (N_1564,N_1211,N_1387);
and U1565 (N_1565,N_1226,N_1389);
and U1566 (N_1566,N_1236,N_1364);
nand U1567 (N_1567,N_1250,N_1265);
and U1568 (N_1568,N_1397,N_1302);
xnor U1569 (N_1569,N_1266,N_1360);
and U1570 (N_1570,N_1280,N_1215);
and U1571 (N_1571,N_1368,N_1283);
nor U1572 (N_1572,N_1230,N_1279);
or U1573 (N_1573,N_1290,N_1253);
nand U1574 (N_1574,N_1360,N_1329);
nand U1575 (N_1575,N_1316,N_1328);
nor U1576 (N_1576,N_1377,N_1248);
xnor U1577 (N_1577,N_1251,N_1348);
or U1578 (N_1578,N_1236,N_1233);
nand U1579 (N_1579,N_1307,N_1345);
nand U1580 (N_1580,N_1371,N_1387);
nor U1581 (N_1581,N_1295,N_1285);
and U1582 (N_1582,N_1278,N_1307);
and U1583 (N_1583,N_1337,N_1397);
and U1584 (N_1584,N_1363,N_1209);
xor U1585 (N_1585,N_1326,N_1375);
nor U1586 (N_1586,N_1347,N_1326);
nor U1587 (N_1587,N_1263,N_1300);
nor U1588 (N_1588,N_1278,N_1390);
nor U1589 (N_1589,N_1235,N_1383);
nor U1590 (N_1590,N_1346,N_1297);
nor U1591 (N_1591,N_1340,N_1335);
or U1592 (N_1592,N_1393,N_1294);
nand U1593 (N_1593,N_1382,N_1301);
and U1594 (N_1594,N_1334,N_1344);
or U1595 (N_1595,N_1316,N_1394);
or U1596 (N_1596,N_1324,N_1317);
nand U1597 (N_1597,N_1274,N_1275);
nor U1598 (N_1598,N_1353,N_1234);
nor U1599 (N_1599,N_1371,N_1327);
or U1600 (N_1600,N_1418,N_1424);
and U1601 (N_1601,N_1595,N_1425);
and U1602 (N_1602,N_1591,N_1528);
nand U1603 (N_1603,N_1489,N_1509);
or U1604 (N_1604,N_1477,N_1561);
and U1605 (N_1605,N_1423,N_1476);
and U1606 (N_1606,N_1408,N_1438);
xor U1607 (N_1607,N_1463,N_1593);
xor U1608 (N_1608,N_1565,N_1519);
nand U1609 (N_1609,N_1479,N_1483);
nor U1610 (N_1610,N_1566,N_1574);
nor U1611 (N_1611,N_1536,N_1441);
nor U1612 (N_1612,N_1572,N_1410);
nand U1613 (N_1613,N_1541,N_1471);
and U1614 (N_1614,N_1472,N_1559);
nand U1615 (N_1615,N_1415,N_1568);
and U1616 (N_1616,N_1551,N_1419);
and U1617 (N_1617,N_1475,N_1432);
nor U1618 (N_1618,N_1417,N_1445);
and U1619 (N_1619,N_1433,N_1443);
nor U1620 (N_1620,N_1465,N_1490);
or U1621 (N_1621,N_1436,N_1546);
and U1622 (N_1622,N_1567,N_1409);
nand U1623 (N_1623,N_1526,N_1442);
or U1624 (N_1624,N_1531,N_1404);
xor U1625 (N_1625,N_1511,N_1462);
nand U1626 (N_1626,N_1598,N_1557);
and U1627 (N_1627,N_1422,N_1599);
or U1628 (N_1628,N_1553,N_1579);
xor U1629 (N_1629,N_1468,N_1429);
or U1630 (N_1630,N_1555,N_1493);
xor U1631 (N_1631,N_1495,N_1427);
nor U1632 (N_1632,N_1570,N_1460);
and U1633 (N_1633,N_1401,N_1510);
nand U1634 (N_1634,N_1416,N_1560);
and U1635 (N_1635,N_1485,N_1459);
and U1636 (N_1636,N_1525,N_1597);
xor U1637 (N_1637,N_1512,N_1558);
and U1638 (N_1638,N_1480,N_1543);
nand U1639 (N_1639,N_1503,N_1529);
and U1640 (N_1640,N_1521,N_1542);
xnor U1641 (N_1641,N_1478,N_1486);
or U1642 (N_1642,N_1469,N_1513);
nand U1643 (N_1643,N_1467,N_1447);
nand U1644 (N_1644,N_1548,N_1446);
and U1645 (N_1645,N_1589,N_1538);
xor U1646 (N_1646,N_1573,N_1596);
nor U1647 (N_1647,N_1474,N_1584);
nand U1648 (N_1648,N_1544,N_1554);
nor U1649 (N_1649,N_1564,N_1498);
nor U1650 (N_1650,N_1547,N_1497);
nor U1651 (N_1651,N_1535,N_1583);
or U1652 (N_1652,N_1403,N_1481);
xor U1653 (N_1653,N_1507,N_1407);
and U1654 (N_1654,N_1435,N_1414);
and U1655 (N_1655,N_1545,N_1585);
nor U1656 (N_1656,N_1426,N_1552);
or U1657 (N_1657,N_1492,N_1444);
nand U1658 (N_1658,N_1540,N_1452);
nor U1659 (N_1659,N_1451,N_1496);
nand U1660 (N_1660,N_1488,N_1508);
or U1661 (N_1661,N_1412,N_1580);
xor U1662 (N_1662,N_1400,N_1502);
nand U1663 (N_1663,N_1491,N_1581);
nor U1664 (N_1664,N_1549,N_1517);
or U1665 (N_1665,N_1537,N_1448);
and U1666 (N_1666,N_1437,N_1505);
nand U1667 (N_1667,N_1587,N_1501);
nor U1668 (N_1668,N_1430,N_1516);
and U1669 (N_1669,N_1473,N_1482);
nor U1670 (N_1670,N_1523,N_1420);
nand U1671 (N_1671,N_1450,N_1457);
or U1672 (N_1672,N_1456,N_1569);
xor U1673 (N_1673,N_1504,N_1461);
and U1674 (N_1674,N_1402,N_1454);
nand U1675 (N_1675,N_1588,N_1571);
or U1676 (N_1676,N_1434,N_1440);
xnor U1677 (N_1677,N_1453,N_1464);
nor U1678 (N_1678,N_1562,N_1577);
and U1679 (N_1679,N_1431,N_1594);
or U1680 (N_1680,N_1439,N_1406);
nand U1681 (N_1681,N_1532,N_1518);
and U1682 (N_1682,N_1522,N_1458);
or U1683 (N_1683,N_1582,N_1586);
nand U1684 (N_1684,N_1411,N_1455);
and U1685 (N_1685,N_1592,N_1494);
nand U1686 (N_1686,N_1506,N_1515);
nor U1687 (N_1687,N_1524,N_1484);
and U1688 (N_1688,N_1533,N_1428);
nand U1689 (N_1689,N_1421,N_1534);
or U1690 (N_1690,N_1530,N_1520);
nor U1691 (N_1691,N_1563,N_1550);
nor U1692 (N_1692,N_1487,N_1514);
nor U1693 (N_1693,N_1413,N_1578);
xor U1694 (N_1694,N_1405,N_1466);
nor U1695 (N_1695,N_1470,N_1556);
and U1696 (N_1696,N_1500,N_1449);
or U1697 (N_1697,N_1590,N_1527);
or U1698 (N_1698,N_1576,N_1539);
and U1699 (N_1699,N_1575,N_1499);
nor U1700 (N_1700,N_1587,N_1505);
nor U1701 (N_1701,N_1569,N_1464);
and U1702 (N_1702,N_1525,N_1519);
and U1703 (N_1703,N_1552,N_1425);
or U1704 (N_1704,N_1479,N_1499);
nand U1705 (N_1705,N_1562,N_1599);
or U1706 (N_1706,N_1545,N_1503);
and U1707 (N_1707,N_1481,N_1594);
nor U1708 (N_1708,N_1586,N_1510);
and U1709 (N_1709,N_1421,N_1419);
nor U1710 (N_1710,N_1522,N_1417);
nand U1711 (N_1711,N_1485,N_1419);
nand U1712 (N_1712,N_1421,N_1592);
or U1713 (N_1713,N_1575,N_1467);
or U1714 (N_1714,N_1478,N_1523);
nand U1715 (N_1715,N_1429,N_1505);
nor U1716 (N_1716,N_1510,N_1430);
nand U1717 (N_1717,N_1436,N_1533);
nor U1718 (N_1718,N_1501,N_1440);
or U1719 (N_1719,N_1503,N_1455);
nand U1720 (N_1720,N_1424,N_1501);
nand U1721 (N_1721,N_1533,N_1515);
nand U1722 (N_1722,N_1466,N_1421);
or U1723 (N_1723,N_1550,N_1425);
and U1724 (N_1724,N_1528,N_1552);
or U1725 (N_1725,N_1431,N_1461);
nand U1726 (N_1726,N_1555,N_1590);
nand U1727 (N_1727,N_1439,N_1417);
or U1728 (N_1728,N_1434,N_1422);
xnor U1729 (N_1729,N_1565,N_1488);
nor U1730 (N_1730,N_1424,N_1542);
or U1731 (N_1731,N_1473,N_1407);
and U1732 (N_1732,N_1507,N_1433);
nand U1733 (N_1733,N_1486,N_1477);
nor U1734 (N_1734,N_1545,N_1516);
nor U1735 (N_1735,N_1411,N_1593);
and U1736 (N_1736,N_1541,N_1543);
nor U1737 (N_1737,N_1431,N_1508);
or U1738 (N_1738,N_1464,N_1496);
nand U1739 (N_1739,N_1424,N_1551);
or U1740 (N_1740,N_1524,N_1544);
xnor U1741 (N_1741,N_1555,N_1565);
or U1742 (N_1742,N_1431,N_1526);
or U1743 (N_1743,N_1593,N_1586);
and U1744 (N_1744,N_1536,N_1517);
nand U1745 (N_1745,N_1540,N_1554);
nand U1746 (N_1746,N_1402,N_1419);
xnor U1747 (N_1747,N_1559,N_1435);
nor U1748 (N_1748,N_1567,N_1556);
nand U1749 (N_1749,N_1521,N_1547);
nand U1750 (N_1750,N_1532,N_1566);
nand U1751 (N_1751,N_1548,N_1428);
and U1752 (N_1752,N_1493,N_1537);
xor U1753 (N_1753,N_1470,N_1498);
or U1754 (N_1754,N_1493,N_1577);
or U1755 (N_1755,N_1420,N_1442);
or U1756 (N_1756,N_1505,N_1545);
nor U1757 (N_1757,N_1405,N_1410);
nand U1758 (N_1758,N_1549,N_1587);
nor U1759 (N_1759,N_1444,N_1525);
or U1760 (N_1760,N_1555,N_1575);
nor U1761 (N_1761,N_1483,N_1508);
nand U1762 (N_1762,N_1566,N_1520);
nand U1763 (N_1763,N_1506,N_1493);
and U1764 (N_1764,N_1516,N_1526);
or U1765 (N_1765,N_1469,N_1431);
and U1766 (N_1766,N_1549,N_1443);
nand U1767 (N_1767,N_1584,N_1536);
nand U1768 (N_1768,N_1450,N_1508);
and U1769 (N_1769,N_1518,N_1494);
and U1770 (N_1770,N_1594,N_1464);
or U1771 (N_1771,N_1401,N_1426);
or U1772 (N_1772,N_1510,N_1420);
nand U1773 (N_1773,N_1417,N_1458);
or U1774 (N_1774,N_1434,N_1458);
nor U1775 (N_1775,N_1475,N_1531);
nand U1776 (N_1776,N_1549,N_1558);
or U1777 (N_1777,N_1522,N_1574);
or U1778 (N_1778,N_1435,N_1491);
or U1779 (N_1779,N_1547,N_1525);
or U1780 (N_1780,N_1514,N_1570);
nor U1781 (N_1781,N_1506,N_1571);
nor U1782 (N_1782,N_1546,N_1422);
or U1783 (N_1783,N_1574,N_1599);
or U1784 (N_1784,N_1505,N_1503);
and U1785 (N_1785,N_1445,N_1459);
nand U1786 (N_1786,N_1424,N_1466);
and U1787 (N_1787,N_1501,N_1443);
nor U1788 (N_1788,N_1406,N_1493);
nor U1789 (N_1789,N_1438,N_1458);
xor U1790 (N_1790,N_1458,N_1520);
nor U1791 (N_1791,N_1435,N_1581);
and U1792 (N_1792,N_1598,N_1483);
xor U1793 (N_1793,N_1503,N_1520);
or U1794 (N_1794,N_1586,N_1592);
or U1795 (N_1795,N_1465,N_1545);
or U1796 (N_1796,N_1597,N_1523);
xor U1797 (N_1797,N_1403,N_1411);
nor U1798 (N_1798,N_1547,N_1448);
nor U1799 (N_1799,N_1582,N_1420);
nand U1800 (N_1800,N_1648,N_1623);
nor U1801 (N_1801,N_1655,N_1699);
xor U1802 (N_1802,N_1702,N_1660);
nor U1803 (N_1803,N_1711,N_1675);
and U1804 (N_1804,N_1767,N_1677);
or U1805 (N_1805,N_1792,N_1734);
or U1806 (N_1806,N_1770,N_1785);
or U1807 (N_1807,N_1708,N_1682);
nor U1808 (N_1808,N_1728,N_1688);
or U1809 (N_1809,N_1704,N_1741);
nand U1810 (N_1810,N_1672,N_1755);
nor U1811 (N_1811,N_1766,N_1636);
xor U1812 (N_1812,N_1680,N_1723);
and U1813 (N_1813,N_1600,N_1798);
and U1814 (N_1814,N_1662,N_1773);
nor U1815 (N_1815,N_1628,N_1753);
or U1816 (N_1816,N_1709,N_1697);
nand U1817 (N_1817,N_1657,N_1629);
or U1818 (N_1818,N_1713,N_1687);
nor U1819 (N_1819,N_1787,N_1790);
nand U1820 (N_1820,N_1645,N_1668);
and U1821 (N_1821,N_1640,N_1779);
or U1822 (N_1822,N_1769,N_1611);
nand U1823 (N_1823,N_1671,N_1650);
and U1824 (N_1824,N_1693,N_1703);
or U1825 (N_1825,N_1617,N_1701);
nand U1826 (N_1826,N_1724,N_1742);
nor U1827 (N_1827,N_1663,N_1794);
and U1828 (N_1828,N_1762,N_1620);
nor U1829 (N_1829,N_1758,N_1780);
or U1830 (N_1830,N_1615,N_1729);
nand U1831 (N_1831,N_1642,N_1759);
or U1832 (N_1832,N_1637,N_1696);
and U1833 (N_1833,N_1646,N_1659);
nor U1834 (N_1834,N_1788,N_1643);
nor U1835 (N_1835,N_1684,N_1797);
nor U1836 (N_1836,N_1695,N_1707);
nor U1837 (N_1837,N_1745,N_1653);
and U1838 (N_1838,N_1781,N_1722);
or U1839 (N_1839,N_1782,N_1743);
or U1840 (N_1840,N_1606,N_1602);
nand U1841 (N_1841,N_1764,N_1661);
nand U1842 (N_1842,N_1667,N_1656);
or U1843 (N_1843,N_1618,N_1717);
xnor U1844 (N_1844,N_1778,N_1774);
nand U1845 (N_1845,N_1720,N_1624);
nor U1846 (N_1846,N_1613,N_1754);
nand U1847 (N_1847,N_1666,N_1705);
nand U1848 (N_1848,N_1799,N_1768);
nand U1849 (N_1849,N_1749,N_1691);
and U1850 (N_1850,N_1689,N_1761);
nor U1851 (N_1851,N_1683,N_1725);
nand U1852 (N_1852,N_1679,N_1738);
nand U1853 (N_1853,N_1706,N_1612);
nor U1854 (N_1854,N_1789,N_1748);
nor U1855 (N_1855,N_1669,N_1710);
nand U1856 (N_1856,N_1760,N_1601);
xnor U1857 (N_1857,N_1721,N_1783);
nand U1858 (N_1858,N_1639,N_1673);
xnor U1859 (N_1859,N_1791,N_1647);
or U1860 (N_1860,N_1775,N_1736);
nor U1861 (N_1861,N_1652,N_1700);
and U1862 (N_1862,N_1670,N_1616);
and U1863 (N_1863,N_1746,N_1777);
and U1864 (N_1864,N_1651,N_1609);
and U1865 (N_1865,N_1737,N_1765);
xnor U1866 (N_1866,N_1772,N_1719);
or U1867 (N_1867,N_1603,N_1622);
xor U1868 (N_1868,N_1727,N_1739);
and U1869 (N_1869,N_1756,N_1751);
nand U1870 (N_1870,N_1690,N_1625);
xor U1871 (N_1871,N_1744,N_1604);
and U1872 (N_1872,N_1776,N_1757);
nor U1873 (N_1873,N_1784,N_1674);
or U1874 (N_1874,N_1658,N_1750);
or U1875 (N_1875,N_1610,N_1712);
or U1876 (N_1876,N_1641,N_1681);
or U1877 (N_1877,N_1678,N_1793);
or U1878 (N_1878,N_1771,N_1664);
and U1879 (N_1879,N_1698,N_1715);
nand U1880 (N_1880,N_1731,N_1726);
nand U1881 (N_1881,N_1635,N_1665);
and U1882 (N_1882,N_1714,N_1644);
nand U1883 (N_1883,N_1608,N_1732);
and U1884 (N_1884,N_1735,N_1716);
or U1885 (N_1885,N_1638,N_1676);
nand U1886 (N_1886,N_1786,N_1796);
xnor U1887 (N_1887,N_1631,N_1718);
nor U1888 (N_1888,N_1747,N_1633);
nor U1889 (N_1889,N_1634,N_1733);
nand U1890 (N_1890,N_1685,N_1632);
or U1891 (N_1891,N_1694,N_1607);
nor U1892 (N_1892,N_1649,N_1730);
nor U1893 (N_1893,N_1752,N_1627);
and U1894 (N_1894,N_1692,N_1740);
or U1895 (N_1895,N_1763,N_1605);
nand U1896 (N_1896,N_1621,N_1795);
nor U1897 (N_1897,N_1654,N_1614);
or U1898 (N_1898,N_1630,N_1626);
nand U1899 (N_1899,N_1686,N_1619);
or U1900 (N_1900,N_1775,N_1674);
or U1901 (N_1901,N_1667,N_1739);
nor U1902 (N_1902,N_1790,N_1604);
xor U1903 (N_1903,N_1690,N_1688);
nor U1904 (N_1904,N_1618,N_1710);
nor U1905 (N_1905,N_1693,N_1635);
xnor U1906 (N_1906,N_1741,N_1600);
and U1907 (N_1907,N_1770,N_1679);
or U1908 (N_1908,N_1603,N_1789);
nand U1909 (N_1909,N_1610,N_1710);
nor U1910 (N_1910,N_1779,N_1759);
nor U1911 (N_1911,N_1639,N_1607);
nor U1912 (N_1912,N_1743,N_1615);
nor U1913 (N_1913,N_1723,N_1726);
nor U1914 (N_1914,N_1685,N_1604);
nand U1915 (N_1915,N_1737,N_1725);
nand U1916 (N_1916,N_1682,N_1649);
nand U1917 (N_1917,N_1679,N_1642);
nand U1918 (N_1918,N_1615,N_1759);
and U1919 (N_1919,N_1727,N_1635);
and U1920 (N_1920,N_1621,N_1752);
or U1921 (N_1921,N_1773,N_1607);
and U1922 (N_1922,N_1777,N_1776);
nand U1923 (N_1923,N_1742,N_1792);
and U1924 (N_1924,N_1702,N_1741);
and U1925 (N_1925,N_1740,N_1691);
nor U1926 (N_1926,N_1687,N_1769);
or U1927 (N_1927,N_1698,N_1664);
xor U1928 (N_1928,N_1750,N_1775);
nand U1929 (N_1929,N_1675,N_1603);
and U1930 (N_1930,N_1776,N_1758);
or U1931 (N_1931,N_1629,N_1656);
nor U1932 (N_1932,N_1721,N_1774);
nand U1933 (N_1933,N_1707,N_1756);
and U1934 (N_1934,N_1633,N_1799);
or U1935 (N_1935,N_1614,N_1681);
and U1936 (N_1936,N_1742,N_1638);
nor U1937 (N_1937,N_1618,N_1795);
and U1938 (N_1938,N_1640,N_1657);
and U1939 (N_1939,N_1734,N_1770);
or U1940 (N_1940,N_1606,N_1766);
and U1941 (N_1941,N_1752,N_1784);
or U1942 (N_1942,N_1669,N_1600);
nor U1943 (N_1943,N_1712,N_1611);
nand U1944 (N_1944,N_1624,N_1724);
or U1945 (N_1945,N_1770,N_1784);
and U1946 (N_1946,N_1654,N_1655);
or U1947 (N_1947,N_1670,N_1736);
or U1948 (N_1948,N_1763,N_1619);
and U1949 (N_1949,N_1733,N_1618);
xnor U1950 (N_1950,N_1763,N_1706);
or U1951 (N_1951,N_1729,N_1708);
or U1952 (N_1952,N_1663,N_1735);
or U1953 (N_1953,N_1649,N_1651);
xor U1954 (N_1954,N_1796,N_1652);
or U1955 (N_1955,N_1611,N_1645);
or U1956 (N_1956,N_1736,N_1725);
or U1957 (N_1957,N_1685,N_1663);
or U1958 (N_1958,N_1606,N_1640);
nand U1959 (N_1959,N_1626,N_1793);
nand U1960 (N_1960,N_1797,N_1618);
nor U1961 (N_1961,N_1793,N_1714);
nor U1962 (N_1962,N_1617,N_1793);
and U1963 (N_1963,N_1798,N_1601);
nand U1964 (N_1964,N_1709,N_1797);
nand U1965 (N_1965,N_1604,N_1631);
and U1966 (N_1966,N_1663,N_1782);
xor U1967 (N_1967,N_1745,N_1704);
or U1968 (N_1968,N_1722,N_1717);
nor U1969 (N_1969,N_1683,N_1632);
or U1970 (N_1970,N_1779,N_1774);
and U1971 (N_1971,N_1744,N_1777);
or U1972 (N_1972,N_1710,N_1663);
xnor U1973 (N_1973,N_1730,N_1617);
and U1974 (N_1974,N_1780,N_1680);
or U1975 (N_1975,N_1748,N_1744);
nor U1976 (N_1976,N_1744,N_1646);
and U1977 (N_1977,N_1738,N_1639);
nor U1978 (N_1978,N_1654,N_1747);
xor U1979 (N_1979,N_1710,N_1608);
nor U1980 (N_1980,N_1685,N_1728);
and U1981 (N_1981,N_1725,N_1716);
and U1982 (N_1982,N_1701,N_1678);
and U1983 (N_1983,N_1743,N_1682);
nand U1984 (N_1984,N_1728,N_1726);
nor U1985 (N_1985,N_1727,N_1662);
xor U1986 (N_1986,N_1729,N_1786);
or U1987 (N_1987,N_1751,N_1785);
and U1988 (N_1988,N_1712,N_1718);
or U1989 (N_1989,N_1737,N_1646);
nand U1990 (N_1990,N_1682,N_1795);
or U1991 (N_1991,N_1633,N_1753);
or U1992 (N_1992,N_1744,N_1608);
or U1993 (N_1993,N_1623,N_1607);
or U1994 (N_1994,N_1601,N_1781);
or U1995 (N_1995,N_1784,N_1631);
and U1996 (N_1996,N_1764,N_1702);
nor U1997 (N_1997,N_1676,N_1700);
and U1998 (N_1998,N_1776,N_1678);
and U1999 (N_1999,N_1749,N_1753);
nand U2000 (N_2000,N_1942,N_1949);
or U2001 (N_2001,N_1866,N_1848);
xnor U2002 (N_2002,N_1981,N_1882);
xor U2003 (N_2003,N_1997,N_1965);
and U2004 (N_2004,N_1864,N_1881);
nor U2005 (N_2005,N_1956,N_1998);
or U2006 (N_2006,N_1903,N_1976);
xnor U2007 (N_2007,N_1802,N_1800);
nand U2008 (N_2008,N_1854,N_1911);
and U2009 (N_2009,N_1839,N_1850);
nand U2010 (N_2010,N_1885,N_1992);
xor U2011 (N_2011,N_1963,N_1807);
nand U2012 (N_2012,N_1991,N_1805);
nor U2013 (N_2013,N_1899,N_1862);
nand U2014 (N_2014,N_1833,N_1817);
and U2015 (N_2015,N_1892,N_1818);
nor U2016 (N_2016,N_1896,N_1948);
and U2017 (N_2017,N_1910,N_1970);
or U2018 (N_2018,N_1951,N_1927);
or U2019 (N_2019,N_1883,N_1984);
or U2020 (N_2020,N_1943,N_1977);
and U2021 (N_2021,N_1897,N_1995);
and U2022 (N_2022,N_1929,N_1823);
and U2023 (N_2023,N_1863,N_1962);
or U2024 (N_2024,N_1928,N_1810);
nor U2025 (N_2025,N_1867,N_1968);
or U2026 (N_2026,N_1923,N_1989);
nand U2027 (N_2027,N_1934,N_1925);
nor U2028 (N_2028,N_1905,N_1974);
nor U2029 (N_2029,N_1874,N_1808);
and U2030 (N_2030,N_1842,N_1827);
or U2031 (N_2031,N_1861,N_1830);
or U2032 (N_2032,N_1868,N_1947);
or U2033 (N_2033,N_1857,N_1824);
and U2034 (N_2034,N_1975,N_1819);
or U2035 (N_2035,N_1811,N_1846);
or U2036 (N_2036,N_1834,N_1994);
or U2037 (N_2037,N_1804,N_1865);
or U2038 (N_2038,N_1849,N_1987);
or U2039 (N_2039,N_1941,N_1843);
xor U2040 (N_2040,N_1806,N_1930);
or U2041 (N_2041,N_1856,N_1946);
and U2042 (N_2042,N_1958,N_1888);
nand U2043 (N_2043,N_1999,N_1954);
xor U2044 (N_2044,N_1877,N_1822);
nand U2045 (N_2045,N_1921,N_1935);
xnor U2046 (N_2046,N_1851,N_1973);
and U2047 (N_2047,N_1858,N_1893);
nor U2048 (N_2048,N_1985,N_1960);
and U2049 (N_2049,N_1845,N_1915);
nand U2050 (N_2050,N_1964,N_1966);
or U2051 (N_2051,N_1828,N_1918);
nor U2052 (N_2052,N_1979,N_1957);
nand U2053 (N_2053,N_1990,N_1853);
or U2054 (N_2054,N_1878,N_1838);
and U2055 (N_2055,N_1876,N_1955);
nor U2056 (N_2056,N_1801,N_1870);
or U2057 (N_2057,N_1939,N_1847);
or U2058 (N_2058,N_1887,N_1836);
nor U2059 (N_2059,N_1931,N_1936);
or U2060 (N_2060,N_1944,N_1873);
nand U2061 (N_2061,N_1815,N_1829);
or U2062 (N_2062,N_1803,N_1891);
and U2063 (N_2063,N_1837,N_1913);
and U2064 (N_2064,N_1986,N_1926);
and U2065 (N_2065,N_1826,N_1831);
nand U2066 (N_2066,N_1821,N_1832);
nand U2067 (N_2067,N_1961,N_1982);
nand U2068 (N_2068,N_1809,N_1914);
xnor U2069 (N_2069,N_1884,N_1814);
and U2070 (N_2070,N_1904,N_1901);
nand U2071 (N_2071,N_1967,N_1938);
nor U2072 (N_2072,N_1855,N_1906);
or U2073 (N_2073,N_1875,N_1889);
and U2074 (N_2074,N_1907,N_1971);
xnor U2075 (N_2075,N_1859,N_1912);
nand U2076 (N_2076,N_1860,N_1812);
nor U2077 (N_2077,N_1813,N_1872);
nor U2078 (N_2078,N_1886,N_1890);
and U2079 (N_2079,N_1945,N_1895);
nand U2080 (N_2080,N_1880,N_1983);
nor U2081 (N_2081,N_1993,N_1898);
xnor U2082 (N_2082,N_1953,N_1869);
or U2083 (N_2083,N_1852,N_1950);
or U2084 (N_2084,N_1969,N_1916);
or U2085 (N_2085,N_1920,N_1825);
xnor U2086 (N_2086,N_1902,N_1933);
nand U2087 (N_2087,N_1940,N_1919);
nand U2088 (N_2088,N_1988,N_1937);
nand U2089 (N_2089,N_1922,N_1900);
nand U2090 (N_2090,N_1980,N_1996);
nor U2091 (N_2091,N_1820,N_1841);
nand U2092 (N_2092,N_1879,N_1871);
or U2093 (N_2093,N_1932,N_1952);
or U2094 (N_2094,N_1894,N_1917);
nor U2095 (N_2095,N_1978,N_1908);
nand U2096 (N_2096,N_1924,N_1909);
nor U2097 (N_2097,N_1844,N_1816);
nand U2098 (N_2098,N_1959,N_1835);
nor U2099 (N_2099,N_1840,N_1972);
and U2100 (N_2100,N_1827,N_1947);
nor U2101 (N_2101,N_1848,N_1898);
nand U2102 (N_2102,N_1930,N_1862);
nor U2103 (N_2103,N_1997,N_1887);
and U2104 (N_2104,N_1919,N_1822);
or U2105 (N_2105,N_1839,N_1956);
or U2106 (N_2106,N_1833,N_1892);
nand U2107 (N_2107,N_1950,N_1879);
and U2108 (N_2108,N_1893,N_1849);
or U2109 (N_2109,N_1992,N_1896);
xor U2110 (N_2110,N_1841,N_1836);
nand U2111 (N_2111,N_1966,N_1962);
and U2112 (N_2112,N_1864,N_1811);
or U2113 (N_2113,N_1933,N_1847);
and U2114 (N_2114,N_1981,N_1832);
nand U2115 (N_2115,N_1948,N_1965);
or U2116 (N_2116,N_1852,N_1942);
nand U2117 (N_2117,N_1943,N_1970);
nand U2118 (N_2118,N_1864,N_1806);
and U2119 (N_2119,N_1985,N_1993);
and U2120 (N_2120,N_1840,N_1872);
or U2121 (N_2121,N_1835,N_1916);
nand U2122 (N_2122,N_1816,N_1925);
or U2123 (N_2123,N_1922,N_1889);
xor U2124 (N_2124,N_1818,N_1905);
or U2125 (N_2125,N_1981,N_1809);
nand U2126 (N_2126,N_1806,N_1872);
or U2127 (N_2127,N_1800,N_1810);
nor U2128 (N_2128,N_1842,N_1828);
nand U2129 (N_2129,N_1834,N_1889);
nor U2130 (N_2130,N_1936,N_1955);
nor U2131 (N_2131,N_1805,N_1863);
nor U2132 (N_2132,N_1981,N_1875);
nor U2133 (N_2133,N_1914,N_1976);
nor U2134 (N_2134,N_1992,N_1952);
nor U2135 (N_2135,N_1993,N_1828);
and U2136 (N_2136,N_1992,N_1965);
nand U2137 (N_2137,N_1891,N_1927);
or U2138 (N_2138,N_1800,N_1917);
and U2139 (N_2139,N_1862,N_1956);
and U2140 (N_2140,N_1993,N_1885);
xor U2141 (N_2141,N_1874,N_1816);
nor U2142 (N_2142,N_1949,N_1937);
nor U2143 (N_2143,N_1808,N_1915);
nor U2144 (N_2144,N_1861,N_1901);
nor U2145 (N_2145,N_1860,N_1937);
xnor U2146 (N_2146,N_1875,N_1879);
and U2147 (N_2147,N_1872,N_1942);
and U2148 (N_2148,N_1820,N_1882);
nor U2149 (N_2149,N_1989,N_1829);
nor U2150 (N_2150,N_1836,N_1821);
or U2151 (N_2151,N_1809,N_1936);
or U2152 (N_2152,N_1993,N_1987);
and U2153 (N_2153,N_1849,N_1965);
or U2154 (N_2154,N_1991,N_1838);
and U2155 (N_2155,N_1808,N_1905);
nand U2156 (N_2156,N_1861,N_1970);
or U2157 (N_2157,N_1803,N_1935);
or U2158 (N_2158,N_1977,N_1817);
nand U2159 (N_2159,N_1975,N_1955);
nand U2160 (N_2160,N_1880,N_1871);
nor U2161 (N_2161,N_1909,N_1894);
and U2162 (N_2162,N_1821,N_1841);
and U2163 (N_2163,N_1834,N_1807);
nor U2164 (N_2164,N_1996,N_1961);
or U2165 (N_2165,N_1969,N_1998);
or U2166 (N_2166,N_1976,N_1990);
or U2167 (N_2167,N_1908,N_1913);
and U2168 (N_2168,N_1821,N_1861);
nor U2169 (N_2169,N_1944,N_1874);
or U2170 (N_2170,N_1899,N_1965);
nor U2171 (N_2171,N_1840,N_1888);
and U2172 (N_2172,N_1858,N_1887);
nor U2173 (N_2173,N_1959,N_1924);
or U2174 (N_2174,N_1858,N_1865);
or U2175 (N_2175,N_1850,N_1829);
or U2176 (N_2176,N_1812,N_1869);
and U2177 (N_2177,N_1973,N_1913);
nor U2178 (N_2178,N_1862,N_1953);
and U2179 (N_2179,N_1936,N_1864);
nand U2180 (N_2180,N_1886,N_1993);
nand U2181 (N_2181,N_1921,N_1809);
or U2182 (N_2182,N_1867,N_1987);
or U2183 (N_2183,N_1953,N_1893);
nand U2184 (N_2184,N_1869,N_1811);
or U2185 (N_2185,N_1963,N_1873);
nand U2186 (N_2186,N_1902,N_1957);
and U2187 (N_2187,N_1979,N_1823);
and U2188 (N_2188,N_1845,N_1969);
and U2189 (N_2189,N_1814,N_1872);
nand U2190 (N_2190,N_1977,N_1933);
xnor U2191 (N_2191,N_1933,N_1822);
and U2192 (N_2192,N_1973,N_1904);
or U2193 (N_2193,N_1942,N_1963);
or U2194 (N_2194,N_1833,N_1965);
nand U2195 (N_2195,N_1936,N_1998);
nand U2196 (N_2196,N_1979,N_1811);
nor U2197 (N_2197,N_1972,N_1809);
nand U2198 (N_2198,N_1940,N_1851);
nand U2199 (N_2199,N_1954,N_1993);
or U2200 (N_2200,N_2039,N_2059);
or U2201 (N_2201,N_2035,N_2187);
nor U2202 (N_2202,N_2163,N_2164);
nor U2203 (N_2203,N_2085,N_2152);
nor U2204 (N_2204,N_2132,N_2155);
nand U2205 (N_2205,N_2173,N_2034);
nand U2206 (N_2206,N_2150,N_2065);
nor U2207 (N_2207,N_2148,N_2041);
nand U2208 (N_2208,N_2190,N_2158);
nand U2209 (N_2209,N_2104,N_2133);
nor U2210 (N_2210,N_2197,N_2151);
nor U2211 (N_2211,N_2018,N_2087);
xnor U2212 (N_2212,N_2052,N_2171);
nor U2213 (N_2213,N_2166,N_2169);
and U2214 (N_2214,N_2023,N_2075);
nor U2215 (N_2215,N_2057,N_2128);
or U2216 (N_2216,N_2020,N_2061);
or U2217 (N_2217,N_2101,N_2116);
or U2218 (N_2218,N_2091,N_2015);
or U2219 (N_2219,N_2198,N_2115);
xor U2220 (N_2220,N_2014,N_2185);
or U2221 (N_2221,N_2043,N_2009);
nor U2222 (N_2222,N_2086,N_2064);
and U2223 (N_2223,N_2017,N_2131);
and U2224 (N_2224,N_2141,N_2097);
or U2225 (N_2225,N_2093,N_2145);
nor U2226 (N_2226,N_2025,N_2120);
nand U2227 (N_2227,N_2144,N_2160);
nand U2228 (N_2228,N_2050,N_2099);
or U2229 (N_2229,N_2032,N_2137);
nor U2230 (N_2230,N_2107,N_2047);
or U2231 (N_2231,N_2054,N_2003);
nand U2232 (N_2232,N_2080,N_2095);
or U2233 (N_2233,N_2109,N_2146);
nor U2234 (N_2234,N_2139,N_2130);
and U2235 (N_2235,N_2196,N_2177);
nand U2236 (N_2236,N_2103,N_2188);
nand U2237 (N_2237,N_2172,N_2077);
nand U2238 (N_2238,N_2011,N_2090);
and U2239 (N_2239,N_2111,N_2005);
or U2240 (N_2240,N_2036,N_2094);
xor U2241 (N_2241,N_2167,N_2089);
nand U2242 (N_2242,N_2176,N_2175);
nor U2243 (N_2243,N_2021,N_2063);
or U2244 (N_2244,N_2027,N_2037);
xnor U2245 (N_2245,N_2049,N_2121);
nand U2246 (N_2246,N_2078,N_2118);
or U2247 (N_2247,N_2016,N_2181);
or U2248 (N_2248,N_2042,N_2186);
or U2249 (N_2249,N_2001,N_2066);
xnor U2250 (N_2250,N_2199,N_2100);
and U2251 (N_2251,N_2125,N_2098);
nor U2252 (N_2252,N_2082,N_2123);
or U2253 (N_2253,N_2142,N_2083);
nor U2254 (N_2254,N_2008,N_2012);
nand U2255 (N_2255,N_2108,N_2070);
or U2256 (N_2256,N_2074,N_2106);
and U2257 (N_2257,N_2182,N_2113);
and U2258 (N_2258,N_2067,N_2045);
or U2259 (N_2259,N_2192,N_2129);
nor U2260 (N_2260,N_2117,N_2040);
nand U2261 (N_2261,N_2048,N_2072);
xnor U2262 (N_2262,N_2162,N_2161);
nor U2263 (N_2263,N_2028,N_2156);
nor U2264 (N_2264,N_2159,N_2051);
nor U2265 (N_2265,N_2127,N_2168);
nor U2266 (N_2266,N_2053,N_2126);
and U2267 (N_2267,N_2134,N_2007);
and U2268 (N_2268,N_2143,N_2096);
nor U2269 (N_2269,N_2149,N_2124);
or U2270 (N_2270,N_2030,N_2105);
and U2271 (N_2271,N_2004,N_2102);
nand U2272 (N_2272,N_2062,N_2033);
xor U2273 (N_2273,N_2140,N_2079);
or U2274 (N_2274,N_2058,N_2193);
nor U2275 (N_2275,N_2071,N_2179);
nand U2276 (N_2276,N_2092,N_2138);
or U2277 (N_2277,N_2189,N_2060);
xor U2278 (N_2278,N_2114,N_2147);
and U2279 (N_2279,N_2019,N_2112);
or U2280 (N_2280,N_2044,N_2076);
nand U2281 (N_2281,N_2024,N_2006);
and U2282 (N_2282,N_2136,N_2174);
nor U2283 (N_2283,N_2084,N_2157);
nand U2284 (N_2284,N_2081,N_2013);
nor U2285 (N_2285,N_2031,N_2153);
and U2286 (N_2286,N_2056,N_2010);
nor U2287 (N_2287,N_2002,N_2122);
nand U2288 (N_2288,N_2184,N_2000);
and U2289 (N_2289,N_2195,N_2068);
or U2290 (N_2290,N_2055,N_2170);
nand U2291 (N_2291,N_2191,N_2178);
and U2292 (N_2292,N_2180,N_2029);
nand U2293 (N_2293,N_2110,N_2073);
nor U2294 (N_2294,N_2183,N_2135);
and U2295 (N_2295,N_2069,N_2154);
and U2296 (N_2296,N_2119,N_2194);
nor U2297 (N_2297,N_2026,N_2022);
nand U2298 (N_2298,N_2165,N_2038);
or U2299 (N_2299,N_2046,N_2088);
and U2300 (N_2300,N_2041,N_2123);
nor U2301 (N_2301,N_2075,N_2053);
and U2302 (N_2302,N_2031,N_2174);
nand U2303 (N_2303,N_2055,N_2131);
nand U2304 (N_2304,N_2143,N_2196);
nor U2305 (N_2305,N_2128,N_2069);
or U2306 (N_2306,N_2018,N_2026);
xnor U2307 (N_2307,N_2029,N_2116);
xnor U2308 (N_2308,N_2111,N_2127);
xor U2309 (N_2309,N_2087,N_2058);
nor U2310 (N_2310,N_2088,N_2084);
nand U2311 (N_2311,N_2104,N_2112);
and U2312 (N_2312,N_2047,N_2087);
or U2313 (N_2313,N_2126,N_2166);
or U2314 (N_2314,N_2019,N_2080);
and U2315 (N_2315,N_2193,N_2192);
xor U2316 (N_2316,N_2109,N_2183);
or U2317 (N_2317,N_2198,N_2195);
or U2318 (N_2318,N_2058,N_2180);
xor U2319 (N_2319,N_2121,N_2048);
nor U2320 (N_2320,N_2092,N_2122);
nor U2321 (N_2321,N_2149,N_2091);
nand U2322 (N_2322,N_2051,N_2017);
nand U2323 (N_2323,N_2021,N_2008);
nor U2324 (N_2324,N_2108,N_2028);
and U2325 (N_2325,N_2041,N_2133);
xnor U2326 (N_2326,N_2016,N_2003);
nor U2327 (N_2327,N_2154,N_2075);
and U2328 (N_2328,N_2076,N_2190);
xor U2329 (N_2329,N_2088,N_2147);
and U2330 (N_2330,N_2190,N_2096);
nor U2331 (N_2331,N_2136,N_2168);
nor U2332 (N_2332,N_2038,N_2046);
and U2333 (N_2333,N_2118,N_2194);
or U2334 (N_2334,N_2133,N_2055);
and U2335 (N_2335,N_2134,N_2025);
and U2336 (N_2336,N_2174,N_2111);
or U2337 (N_2337,N_2052,N_2046);
nand U2338 (N_2338,N_2173,N_2015);
and U2339 (N_2339,N_2099,N_2046);
and U2340 (N_2340,N_2055,N_2091);
nor U2341 (N_2341,N_2059,N_2001);
and U2342 (N_2342,N_2192,N_2161);
and U2343 (N_2343,N_2096,N_2066);
nor U2344 (N_2344,N_2124,N_2066);
or U2345 (N_2345,N_2189,N_2172);
or U2346 (N_2346,N_2089,N_2005);
xor U2347 (N_2347,N_2005,N_2159);
or U2348 (N_2348,N_2155,N_2044);
nor U2349 (N_2349,N_2173,N_2080);
nor U2350 (N_2350,N_2058,N_2132);
nor U2351 (N_2351,N_2198,N_2095);
and U2352 (N_2352,N_2178,N_2148);
and U2353 (N_2353,N_2014,N_2094);
and U2354 (N_2354,N_2168,N_2124);
nand U2355 (N_2355,N_2149,N_2077);
xnor U2356 (N_2356,N_2013,N_2082);
and U2357 (N_2357,N_2076,N_2103);
and U2358 (N_2358,N_2145,N_2156);
nor U2359 (N_2359,N_2005,N_2172);
or U2360 (N_2360,N_2076,N_2146);
or U2361 (N_2361,N_2098,N_2103);
nand U2362 (N_2362,N_2027,N_2167);
and U2363 (N_2363,N_2011,N_2072);
nand U2364 (N_2364,N_2149,N_2001);
nor U2365 (N_2365,N_2179,N_2096);
xnor U2366 (N_2366,N_2067,N_2033);
and U2367 (N_2367,N_2187,N_2130);
xnor U2368 (N_2368,N_2021,N_2062);
nand U2369 (N_2369,N_2142,N_2067);
and U2370 (N_2370,N_2071,N_2061);
nand U2371 (N_2371,N_2054,N_2012);
and U2372 (N_2372,N_2074,N_2060);
nand U2373 (N_2373,N_2120,N_2183);
or U2374 (N_2374,N_2089,N_2079);
and U2375 (N_2375,N_2078,N_2004);
and U2376 (N_2376,N_2015,N_2165);
and U2377 (N_2377,N_2039,N_2190);
or U2378 (N_2378,N_2052,N_2069);
xnor U2379 (N_2379,N_2017,N_2130);
or U2380 (N_2380,N_2074,N_2103);
and U2381 (N_2381,N_2023,N_2127);
nor U2382 (N_2382,N_2164,N_2182);
and U2383 (N_2383,N_2174,N_2130);
nand U2384 (N_2384,N_2007,N_2035);
or U2385 (N_2385,N_2144,N_2017);
nor U2386 (N_2386,N_2002,N_2142);
xor U2387 (N_2387,N_2174,N_2116);
and U2388 (N_2388,N_2199,N_2158);
nor U2389 (N_2389,N_2134,N_2084);
and U2390 (N_2390,N_2122,N_2044);
nor U2391 (N_2391,N_2169,N_2185);
and U2392 (N_2392,N_2156,N_2023);
or U2393 (N_2393,N_2046,N_2044);
and U2394 (N_2394,N_2195,N_2132);
or U2395 (N_2395,N_2055,N_2038);
nand U2396 (N_2396,N_2090,N_2164);
or U2397 (N_2397,N_2098,N_2150);
nand U2398 (N_2398,N_2001,N_2159);
and U2399 (N_2399,N_2135,N_2125);
nand U2400 (N_2400,N_2328,N_2360);
nor U2401 (N_2401,N_2279,N_2305);
and U2402 (N_2402,N_2315,N_2340);
nor U2403 (N_2403,N_2200,N_2311);
and U2404 (N_2404,N_2239,N_2260);
nand U2405 (N_2405,N_2399,N_2325);
and U2406 (N_2406,N_2378,N_2346);
nor U2407 (N_2407,N_2262,N_2398);
nor U2408 (N_2408,N_2268,N_2206);
xnor U2409 (N_2409,N_2396,N_2240);
or U2410 (N_2410,N_2233,N_2236);
nor U2411 (N_2411,N_2245,N_2283);
nand U2412 (N_2412,N_2292,N_2261);
or U2413 (N_2413,N_2372,N_2229);
nor U2414 (N_2414,N_2308,N_2388);
or U2415 (N_2415,N_2324,N_2291);
or U2416 (N_2416,N_2278,N_2251);
nor U2417 (N_2417,N_2384,N_2216);
nor U2418 (N_2418,N_2242,N_2212);
xnor U2419 (N_2419,N_2366,N_2263);
nor U2420 (N_2420,N_2376,N_2287);
and U2421 (N_2421,N_2395,N_2286);
nand U2422 (N_2422,N_2375,N_2220);
nand U2423 (N_2423,N_2297,N_2390);
or U2424 (N_2424,N_2252,N_2290);
nand U2425 (N_2425,N_2322,N_2243);
or U2426 (N_2426,N_2364,N_2392);
nor U2427 (N_2427,N_2339,N_2202);
and U2428 (N_2428,N_2285,N_2337);
or U2429 (N_2429,N_2205,N_2365);
nand U2430 (N_2430,N_2389,N_2320);
nand U2431 (N_2431,N_2344,N_2303);
nor U2432 (N_2432,N_2317,N_2271);
nand U2433 (N_2433,N_2246,N_2379);
or U2434 (N_2434,N_2218,N_2314);
or U2435 (N_2435,N_2210,N_2357);
nand U2436 (N_2436,N_2345,N_2255);
nor U2437 (N_2437,N_2310,N_2241);
or U2438 (N_2438,N_2333,N_2358);
or U2439 (N_2439,N_2335,N_2288);
or U2440 (N_2440,N_2321,N_2351);
or U2441 (N_2441,N_2282,N_2341);
or U2442 (N_2442,N_2259,N_2383);
nand U2443 (N_2443,N_2382,N_2294);
nand U2444 (N_2444,N_2237,N_2387);
nor U2445 (N_2445,N_2264,N_2250);
or U2446 (N_2446,N_2352,N_2391);
or U2447 (N_2447,N_2369,N_2397);
nand U2448 (N_2448,N_2217,N_2276);
and U2449 (N_2449,N_2232,N_2373);
nand U2450 (N_2450,N_2371,N_2281);
or U2451 (N_2451,N_2309,N_2270);
nand U2452 (N_2452,N_2209,N_2329);
nor U2453 (N_2453,N_2211,N_2207);
xnor U2454 (N_2454,N_2223,N_2221);
or U2455 (N_2455,N_2277,N_2256);
nand U2456 (N_2456,N_2316,N_2258);
or U2457 (N_2457,N_2273,N_2306);
nand U2458 (N_2458,N_2332,N_2295);
nand U2459 (N_2459,N_2253,N_2235);
nor U2460 (N_2460,N_2298,N_2374);
and U2461 (N_2461,N_2368,N_2267);
nor U2462 (N_2462,N_2386,N_2224);
and U2463 (N_2463,N_2234,N_2296);
or U2464 (N_2464,N_2302,N_2204);
nand U2465 (N_2465,N_2331,N_2367);
and U2466 (N_2466,N_2319,N_2214);
nand U2467 (N_2467,N_2330,N_2394);
nand U2468 (N_2468,N_2353,N_2363);
or U2469 (N_2469,N_2327,N_2201);
or U2470 (N_2470,N_2393,N_2342);
or U2471 (N_2471,N_2272,N_2284);
and U2472 (N_2472,N_2257,N_2334);
and U2473 (N_2473,N_2265,N_2348);
nor U2474 (N_2474,N_2381,N_2343);
nor U2475 (N_2475,N_2304,N_2350);
xor U2476 (N_2476,N_2230,N_2222);
and U2477 (N_2477,N_2248,N_2370);
nand U2478 (N_2478,N_2269,N_2238);
nor U2479 (N_2479,N_2359,N_2213);
or U2480 (N_2480,N_2249,N_2231);
nand U2481 (N_2481,N_2203,N_2307);
nor U2482 (N_2482,N_2227,N_2356);
nand U2483 (N_2483,N_2380,N_2361);
nand U2484 (N_2484,N_2354,N_2318);
and U2485 (N_2485,N_2338,N_2347);
or U2486 (N_2486,N_2299,N_2362);
nand U2487 (N_2487,N_2247,N_2323);
xor U2488 (N_2488,N_2301,N_2226);
nand U2489 (N_2489,N_2349,N_2289);
and U2490 (N_2490,N_2275,N_2215);
nand U2491 (N_2491,N_2219,N_2377);
and U2492 (N_2492,N_2280,N_2208);
or U2493 (N_2493,N_2312,N_2336);
or U2494 (N_2494,N_2244,N_2326);
or U2495 (N_2495,N_2274,N_2266);
and U2496 (N_2496,N_2293,N_2254);
or U2497 (N_2497,N_2385,N_2225);
nand U2498 (N_2498,N_2300,N_2355);
xor U2499 (N_2499,N_2228,N_2313);
and U2500 (N_2500,N_2268,N_2360);
xnor U2501 (N_2501,N_2265,N_2366);
and U2502 (N_2502,N_2220,N_2255);
and U2503 (N_2503,N_2216,N_2388);
nor U2504 (N_2504,N_2272,N_2378);
nand U2505 (N_2505,N_2230,N_2394);
and U2506 (N_2506,N_2296,N_2277);
or U2507 (N_2507,N_2376,N_2279);
and U2508 (N_2508,N_2223,N_2382);
or U2509 (N_2509,N_2270,N_2312);
and U2510 (N_2510,N_2262,N_2238);
or U2511 (N_2511,N_2291,N_2394);
xnor U2512 (N_2512,N_2318,N_2369);
or U2513 (N_2513,N_2284,N_2223);
or U2514 (N_2514,N_2226,N_2308);
and U2515 (N_2515,N_2248,N_2349);
xor U2516 (N_2516,N_2238,N_2348);
xnor U2517 (N_2517,N_2287,N_2342);
nor U2518 (N_2518,N_2395,N_2267);
nor U2519 (N_2519,N_2294,N_2362);
nand U2520 (N_2520,N_2249,N_2243);
xor U2521 (N_2521,N_2328,N_2222);
or U2522 (N_2522,N_2330,N_2325);
xor U2523 (N_2523,N_2344,N_2259);
xor U2524 (N_2524,N_2344,N_2364);
or U2525 (N_2525,N_2302,N_2245);
nand U2526 (N_2526,N_2256,N_2212);
xor U2527 (N_2527,N_2222,N_2327);
and U2528 (N_2528,N_2244,N_2258);
nor U2529 (N_2529,N_2263,N_2231);
or U2530 (N_2530,N_2286,N_2331);
and U2531 (N_2531,N_2340,N_2277);
or U2532 (N_2532,N_2308,N_2337);
nor U2533 (N_2533,N_2355,N_2245);
and U2534 (N_2534,N_2330,N_2337);
and U2535 (N_2535,N_2284,N_2325);
nand U2536 (N_2536,N_2365,N_2382);
or U2537 (N_2537,N_2251,N_2372);
or U2538 (N_2538,N_2307,N_2311);
nor U2539 (N_2539,N_2245,N_2378);
and U2540 (N_2540,N_2280,N_2228);
xor U2541 (N_2541,N_2378,N_2286);
or U2542 (N_2542,N_2350,N_2374);
or U2543 (N_2543,N_2202,N_2318);
and U2544 (N_2544,N_2290,N_2357);
nor U2545 (N_2545,N_2355,N_2364);
or U2546 (N_2546,N_2283,N_2371);
nor U2547 (N_2547,N_2329,N_2202);
xnor U2548 (N_2548,N_2230,N_2211);
xnor U2549 (N_2549,N_2221,N_2348);
and U2550 (N_2550,N_2325,N_2306);
or U2551 (N_2551,N_2269,N_2290);
nor U2552 (N_2552,N_2285,N_2215);
xnor U2553 (N_2553,N_2232,N_2399);
or U2554 (N_2554,N_2202,N_2211);
and U2555 (N_2555,N_2310,N_2213);
and U2556 (N_2556,N_2208,N_2217);
nor U2557 (N_2557,N_2303,N_2302);
xnor U2558 (N_2558,N_2383,N_2287);
nor U2559 (N_2559,N_2216,N_2311);
and U2560 (N_2560,N_2368,N_2297);
or U2561 (N_2561,N_2255,N_2347);
or U2562 (N_2562,N_2396,N_2208);
nor U2563 (N_2563,N_2215,N_2277);
or U2564 (N_2564,N_2393,N_2385);
nor U2565 (N_2565,N_2384,N_2388);
nor U2566 (N_2566,N_2323,N_2391);
xnor U2567 (N_2567,N_2353,N_2392);
nor U2568 (N_2568,N_2299,N_2331);
xor U2569 (N_2569,N_2371,N_2315);
nand U2570 (N_2570,N_2323,N_2399);
nand U2571 (N_2571,N_2329,N_2397);
xnor U2572 (N_2572,N_2379,N_2329);
nand U2573 (N_2573,N_2354,N_2293);
or U2574 (N_2574,N_2213,N_2383);
or U2575 (N_2575,N_2367,N_2268);
and U2576 (N_2576,N_2368,N_2340);
and U2577 (N_2577,N_2395,N_2324);
nor U2578 (N_2578,N_2207,N_2270);
or U2579 (N_2579,N_2232,N_2242);
and U2580 (N_2580,N_2397,N_2215);
or U2581 (N_2581,N_2255,N_2321);
xnor U2582 (N_2582,N_2372,N_2262);
nand U2583 (N_2583,N_2291,N_2240);
or U2584 (N_2584,N_2260,N_2341);
and U2585 (N_2585,N_2357,N_2207);
and U2586 (N_2586,N_2338,N_2276);
and U2587 (N_2587,N_2298,N_2232);
nand U2588 (N_2588,N_2391,N_2309);
or U2589 (N_2589,N_2250,N_2301);
nand U2590 (N_2590,N_2346,N_2297);
and U2591 (N_2591,N_2345,N_2236);
and U2592 (N_2592,N_2258,N_2326);
or U2593 (N_2593,N_2337,N_2227);
xnor U2594 (N_2594,N_2345,N_2357);
nor U2595 (N_2595,N_2203,N_2375);
nor U2596 (N_2596,N_2261,N_2392);
and U2597 (N_2597,N_2395,N_2234);
or U2598 (N_2598,N_2333,N_2238);
nand U2599 (N_2599,N_2335,N_2298);
nor U2600 (N_2600,N_2429,N_2463);
nand U2601 (N_2601,N_2476,N_2549);
nand U2602 (N_2602,N_2492,N_2455);
nand U2603 (N_2603,N_2590,N_2504);
or U2604 (N_2604,N_2449,N_2412);
and U2605 (N_2605,N_2406,N_2519);
nor U2606 (N_2606,N_2525,N_2490);
nand U2607 (N_2607,N_2523,N_2530);
or U2608 (N_2608,N_2408,N_2532);
and U2609 (N_2609,N_2464,N_2582);
nor U2610 (N_2610,N_2460,N_2401);
nand U2611 (N_2611,N_2511,N_2407);
nor U2612 (N_2612,N_2415,N_2566);
and U2613 (N_2613,N_2559,N_2453);
xnor U2614 (N_2614,N_2447,N_2423);
and U2615 (N_2615,N_2482,N_2572);
nor U2616 (N_2616,N_2534,N_2461);
and U2617 (N_2617,N_2467,N_2466);
and U2618 (N_2618,N_2574,N_2470);
xnor U2619 (N_2619,N_2521,N_2578);
xnor U2620 (N_2620,N_2434,N_2477);
nor U2621 (N_2621,N_2419,N_2430);
or U2622 (N_2622,N_2550,N_2531);
nor U2623 (N_2623,N_2465,N_2595);
or U2624 (N_2624,N_2493,N_2551);
xor U2625 (N_2625,N_2579,N_2506);
or U2626 (N_2626,N_2581,N_2480);
and U2627 (N_2627,N_2468,N_2562);
nand U2628 (N_2628,N_2588,N_2418);
or U2629 (N_2629,N_2565,N_2560);
nor U2630 (N_2630,N_2503,N_2599);
or U2631 (N_2631,N_2478,N_2402);
xnor U2632 (N_2632,N_2433,N_2427);
and U2633 (N_2633,N_2440,N_2567);
xor U2634 (N_2634,N_2598,N_2553);
nor U2635 (N_2635,N_2454,N_2444);
or U2636 (N_2636,N_2414,N_2556);
xor U2637 (N_2637,N_2594,N_2403);
and U2638 (N_2638,N_2577,N_2555);
nor U2639 (N_2639,N_2538,N_2452);
or U2640 (N_2640,N_2536,N_2587);
and U2641 (N_2641,N_2526,N_2518);
nand U2642 (N_2642,N_2507,N_2462);
or U2643 (N_2643,N_2416,N_2410);
or U2644 (N_2644,N_2573,N_2400);
nor U2645 (N_2645,N_2580,N_2435);
or U2646 (N_2646,N_2443,N_2500);
or U2647 (N_2647,N_2576,N_2437);
nand U2648 (N_2648,N_2527,N_2589);
nor U2649 (N_2649,N_2485,N_2596);
nand U2650 (N_2650,N_2510,N_2546);
xor U2651 (N_2651,N_2489,N_2529);
nand U2652 (N_2652,N_2422,N_2585);
or U2653 (N_2653,N_2513,N_2543);
nand U2654 (N_2654,N_2545,N_2475);
nor U2655 (N_2655,N_2591,N_2471);
and U2656 (N_2656,N_2458,N_2450);
and U2657 (N_2657,N_2584,N_2438);
nand U2658 (N_2658,N_2428,N_2508);
nor U2659 (N_2659,N_2514,N_2439);
nand U2660 (N_2660,N_2424,N_2457);
and U2661 (N_2661,N_2451,N_2495);
nand U2662 (N_2662,N_2487,N_2570);
nor U2663 (N_2663,N_2533,N_2547);
nor U2664 (N_2664,N_2569,N_2420);
and U2665 (N_2665,N_2484,N_2586);
nand U2666 (N_2666,N_2528,N_2575);
nor U2667 (N_2667,N_2524,N_2431);
and U2668 (N_2668,N_2554,N_2542);
nor U2669 (N_2669,N_2516,N_2405);
nor U2670 (N_2670,N_2488,N_2501);
nor U2671 (N_2671,N_2563,N_2446);
or U2672 (N_2672,N_2502,N_2491);
nor U2673 (N_2673,N_2441,N_2459);
and U2674 (N_2674,N_2535,N_2411);
nand U2675 (N_2675,N_2515,N_2522);
nor U2676 (N_2676,N_2512,N_2558);
nor U2677 (N_2677,N_2421,N_2472);
nand U2678 (N_2678,N_2483,N_2442);
nor U2679 (N_2679,N_2593,N_2561);
nor U2680 (N_2680,N_2517,N_2592);
and U2681 (N_2681,N_2456,N_2544);
nor U2682 (N_2682,N_2436,N_2499);
and U2683 (N_2683,N_2520,N_2426);
nor U2684 (N_2684,N_2552,N_2432);
nand U2685 (N_2685,N_2497,N_2496);
nand U2686 (N_2686,N_2539,N_2486);
or U2687 (N_2687,N_2597,N_2425);
xnor U2688 (N_2688,N_2557,N_2404);
and U2689 (N_2689,N_2537,N_2417);
nor U2690 (N_2690,N_2548,N_2564);
and U2691 (N_2691,N_2474,N_2571);
or U2692 (N_2692,N_2540,N_2413);
nand U2693 (N_2693,N_2469,N_2479);
xor U2694 (N_2694,N_2541,N_2448);
xnor U2695 (N_2695,N_2505,N_2494);
and U2696 (N_2696,N_2409,N_2481);
nand U2697 (N_2697,N_2509,N_2445);
nand U2698 (N_2698,N_2473,N_2498);
nor U2699 (N_2699,N_2583,N_2568);
or U2700 (N_2700,N_2503,N_2519);
or U2701 (N_2701,N_2418,N_2566);
and U2702 (N_2702,N_2547,N_2492);
or U2703 (N_2703,N_2464,N_2547);
xnor U2704 (N_2704,N_2426,N_2524);
nor U2705 (N_2705,N_2491,N_2473);
or U2706 (N_2706,N_2440,N_2507);
and U2707 (N_2707,N_2513,N_2575);
or U2708 (N_2708,N_2519,N_2570);
nor U2709 (N_2709,N_2571,N_2553);
nor U2710 (N_2710,N_2507,N_2477);
or U2711 (N_2711,N_2538,N_2512);
and U2712 (N_2712,N_2571,N_2533);
and U2713 (N_2713,N_2454,N_2598);
or U2714 (N_2714,N_2413,N_2406);
and U2715 (N_2715,N_2490,N_2516);
or U2716 (N_2716,N_2570,N_2577);
xor U2717 (N_2717,N_2412,N_2401);
nand U2718 (N_2718,N_2503,N_2552);
or U2719 (N_2719,N_2400,N_2419);
or U2720 (N_2720,N_2444,N_2520);
and U2721 (N_2721,N_2519,N_2571);
and U2722 (N_2722,N_2580,N_2429);
nor U2723 (N_2723,N_2408,N_2445);
nand U2724 (N_2724,N_2463,N_2502);
and U2725 (N_2725,N_2496,N_2500);
nand U2726 (N_2726,N_2494,N_2484);
nor U2727 (N_2727,N_2405,N_2492);
nor U2728 (N_2728,N_2472,N_2467);
or U2729 (N_2729,N_2441,N_2403);
xnor U2730 (N_2730,N_2521,N_2593);
nand U2731 (N_2731,N_2537,N_2581);
or U2732 (N_2732,N_2576,N_2532);
nand U2733 (N_2733,N_2552,N_2494);
or U2734 (N_2734,N_2408,N_2583);
nor U2735 (N_2735,N_2542,N_2446);
and U2736 (N_2736,N_2481,N_2552);
and U2737 (N_2737,N_2588,N_2422);
and U2738 (N_2738,N_2554,N_2524);
nand U2739 (N_2739,N_2562,N_2523);
nand U2740 (N_2740,N_2563,N_2570);
nand U2741 (N_2741,N_2476,N_2579);
nand U2742 (N_2742,N_2572,N_2492);
nand U2743 (N_2743,N_2487,N_2427);
nor U2744 (N_2744,N_2574,N_2425);
or U2745 (N_2745,N_2542,N_2462);
and U2746 (N_2746,N_2470,N_2541);
and U2747 (N_2747,N_2456,N_2576);
or U2748 (N_2748,N_2531,N_2422);
or U2749 (N_2749,N_2545,N_2492);
and U2750 (N_2750,N_2450,N_2577);
nor U2751 (N_2751,N_2437,N_2442);
nand U2752 (N_2752,N_2529,N_2516);
nor U2753 (N_2753,N_2544,N_2580);
nor U2754 (N_2754,N_2451,N_2588);
xor U2755 (N_2755,N_2596,N_2599);
and U2756 (N_2756,N_2508,N_2578);
nor U2757 (N_2757,N_2413,N_2492);
and U2758 (N_2758,N_2436,N_2477);
xnor U2759 (N_2759,N_2474,N_2585);
or U2760 (N_2760,N_2439,N_2471);
or U2761 (N_2761,N_2447,N_2464);
or U2762 (N_2762,N_2469,N_2585);
xor U2763 (N_2763,N_2586,N_2492);
or U2764 (N_2764,N_2422,N_2425);
or U2765 (N_2765,N_2543,N_2532);
nor U2766 (N_2766,N_2595,N_2460);
or U2767 (N_2767,N_2410,N_2475);
nor U2768 (N_2768,N_2472,N_2404);
nor U2769 (N_2769,N_2568,N_2410);
nor U2770 (N_2770,N_2410,N_2412);
and U2771 (N_2771,N_2430,N_2449);
nand U2772 (N_2772,N_2525,N_2583);
and U2773 (N_2773,N_2554,N_2471);
and U2774 (N_2774,N_2568,N_2519);
or U2775 (N_2775,N_2574,N_2401);
and U2776 (N_2776,N_2475,N_2570);
or U2777 (N_2777,N_2479,N_2418);
nand U2778 (N_2778,N_2451,N_2490);
and U2779 (N_2779,N_2468,N_2573);
and U2780 (N_2780,N_2473,N_2567);
and U2781 (N_2781,N_2425,N_2598);
and U2782 (N_2782,N_2571,N_2425);
nand U2783 (N_2783,N_2563,N_2517);
and U2784 (N_2784,N_2431,N_2486);
nand U2785 (N_2785,N_2489,N_2436);
nor U2786 (N_2786,N_2514,N_2512);
nor U2787 (N_2787,N_2583,N_2406);
nand U2788 (N_2788,N_2438,N_2591);
nand U2789 (N_2789,N_2426,N_2457);
xnor U2790 (N_2790,N_2413,N_2484);
and U2791 (N_2791,N_2427,N_2470);
and U2792 (N_2792,N_2489,N_2443);
or U2793 (N_2793,N_2462,N_2504);
nor U2794 (N_2794,N_2548,N_2452);
and U2795 (N_2795,N_2461,N_2533);
or U2796 (N_2796,N_2557,N_2516);
nand U2797 (N_2797,N_2578,N_2448);
and U2798 (N_2798,N_2402,N_2535);
and U2799 (N_2799,N_2588,N_2517);
and U2800 (N_2800,N_2611,N_2672);
or U2801 (N_2801,N_2647,N_2777);
xnor U2802 (N_2802,N_2735,N_2604);
or U2803 (N_2803,N_2600,N_2711);
nand U2804 (N_2804,N_2772,N_2615);
xnor U2805 (N_2805,N_2757,N_2646);
or U2806 (N_2806,N_2743,N_2715);
xor U2807 (N_2807,N_2667,N_2731);
or U2808 (N_2808,N_2751,N_2704);
and U2809 (N_2809,N_2679,N_2783);
or U2810 (N_2810,N_2789,N_2763);
and U2811 (N_2811,N_2775,N_2795);
or U2812 (N_2812,N_2706,N_2678);
or U2813 (N_2813,N_2657,N_2787);
or U2814 (N_2814,N_2788,N_2725);
or U2815 (N_2815,N_2652,N_2702);
nand U2816 (N_2816,N_2753,N_2796);
or U2817 (N_2817,N_2637,N_2768);
nor U2818 (N_2818,N_2693,N_2792);
and U2819 (N_2819,N_2690,N_2684);
nor U2820 (N_2820,N_2614,N_2724);
nand U2821 (N_2821,N_2670,N_2707);
and U2822 (N_2822,N_2630,N_2764);
and U2823 (N_2823,N_2688,N_2761);
nand U2824 (N_2824,N_2713,N_2746);
nor U2825 (N_2825,N_2698,N_2744);
xor U2826 (N_2826,N_2628,N_2649);
xor U2827 (N_2827,N_2709,N_2755);
and U2828 (N_2828,N_2603,N_2616);
and U2829 (N_2829,N_2639,N_2606);
and U2830 (N_2830,N_2786,N_2634);
nand U2831 (N_2831,N_2691,N_2656);
and U2832 (N_2832,N_2723,N_2700);
and U2833 (N_2833,N_2726,N_2754);
nor U2834 (N_2834,N_2780,N_2608);
or U2835 (N_2835,N_2699,N_2607);
or U2836 (N_2836,N_2750,N_2633);
and U2837 (N_2837,N_2640,N_2625);
and U2838 (N_2838,N_2676,N_2624);
nor U2839 (N_2839,N_2722,N_2716);
nor U2840 (N_2840,N_2650,N_2636);
xnor U2841 (N_2841,N_2797,N_2645);
nand U2842 (N_2842,N_2794,N_2718);
xnor U2843 (N_2843,N_2766,N_2728);
or U2844 (N_2844,N_2791,N_2685);
nor U2845 (N_2845,N_2692,N_2623);
nand U2846 (N_2846,N_2681,N_2785);
or U2847 (N_2847,N_2714,N_2626);
nand U2848 (N_2848,N_2641,N_2612);
or U2849 (N_2849,N_2708,N_2793);
or U2850 (N_2850,N_2621,N_2737);
nor U2851 (N_2851,N_2659,N_2701);
nor U2852 (N_2852,N_2631,N_2651);
or U2853 (N_2853,N_2605,N_2696);
or U2854 (N_2854,N_2770,N_2643);
or U2855 (N_2855,N_2655,N_2799);
nor U2856 (N_2856,N_2627,N_2662);
or U2857 (N_2857,N_2776,N_2779);
nand U2858 (N_2858,N_2663,N_2682);
xor U2859 (N_2859,N_2674,N_2760);
nand U2860 (N_2860,N_2617,N_2664);
or U2861 (N_2861,N_2654,N_2620);
and U2862 (N_2862,N_2703,N_2727);
or U2863 (N_2863,N_2671,N_2665);
nor U2864 (N_2864,N_2730,N_2677);
xor U2865 (N_2865,N_2683,N_2778);
nand U2866 (N_2866,N_2781,N_2712);
nand U2867 (N_2867,N_2610,N_2784);
or U2868 (N_2868,N_2748,N_2613);
nand U2869 (N_2869,N_2686,N_2756);
or U2870 (N_2870,N_2762,N_2773);
and U2871 (N_2871,N_2609,N_2644);
nor U2872 (N_2872,N_2798,N_2790);
nand U2873 (N_2873,N_2721,N_2673);
nor U2874 (N_2874,N_2738,N_2745);
nand U2875 (N_2875,N_2759,N_2668);
and U2876 (N_2876,N_2710,N_2648);
or U2877 (N_2877,N_2782,N_2752);
nand U2878 (N_2878,N_2734,N_2632);
nand U2879 (N_2879,N_2622,N_2739);
nor U2880 (N_2880,N_2732,N_2741);
or U2881 (N_2881,N_2618,N_2705);
and U2882 (N_2882,N_2689,N_2602);
and U2883 (N_2883,N_2767,N_2747);
or U2884 (N_2884,N_2695,N_2680);
and U2885 (N_2885,N_2720,N_2660);
nand U2886 (N_2886,N_2697,N_2638);
nor U2887 (N_2887,N_2666,N_2687);
and U2888 (N_2888,N_2642,N_2758);
or U2889 (N_2889,N_2733,N_2601);
or U2890 (N_2890,N_2653,N_2729);
and U2891 (N_2891,N_2774,N_2736);
nor U2892 (N_2892,N_2771,N_2740);
and U2893 (N_2893,N_2694,N_2765);
or U2894 (N_2894,N_2661,N_2658);
xor U2895 (N_2895,N_2619,N_2719);
xor U2896 (N_2896,N_2629,N_2635);
xnor U2897 (N_2897,N_2669,N_2749);
nor U2898 (N_2898,N_2769,N_2717);
and U2899 (N_2899,N_2742,N_2675);
and U2900 (N_2900,N_2770,N_2753);
xor U2901 (N_2901,N_2616,N_2680);
xor U2902 (N_2902,N_2685,N_2768);
nand U2903 (N_2903,N_2778,N_2797);
xnor U2904 (N_2904,N_2633,N_2658);
and U2905 (N_2905,N_2605,N_2785);
xor U2906 (N_2906,N_2751,N_2630);
xnor U2907 (N_2907,N_2769,N_2700);
nor U2908 (N_2908,N_2703,N_2646);
xnor U2909 (N_2909,N_2728,N_2638);
nor U2910 (N_2910,N_2670,N_2765);
nor U2911 (N_2911,N_2725,N_2700);
or U2912 (N_2912,N_2614,N_2653);
nand U2913 (N_2913,N_2691,N_2717);
and U2914 (N_2914,N_2718,N_2671);
and U2915 (N_2915,N_2754,N_2762);
or U2916 (N_2916,N_2752,N_2749);
nand U2917 (N_2917,N_2762,N_2682);
nand U2918 (N_2918,N_2791,N_2763);
nor U2919 (N_2919,N_2641,N_2756);
and U2920 (N_2920,N_2717,N_2777);
nor U2921 (N_2921,N_2624,N_2601);
or U2922 (N_2922,N_2691,N_2644);
or U2923 (N_2923,N_2673,N_2738);
nand U2924 (N_2924,N_2667,N_2705);
nor U2925 (N_2925,N_2672,N_2724);
nor U2926 (N_2926,N_2754,N_2605);
nand U2927 (N_2927,N_2771,N_2624);
or U2928 (N_2928,N_2761,N_2737);
nor U2929 (N_2929,N_2647,N_2685);
xnor U2930 (N_2930,N_2623,N_2669);
nand U2931 (N_2931,N_2761,N_2700);
or U2932 (N_2932,N_2622,N_2791);
nand U2933 (N_2933,N_2713,N_2724);
xnor U2934 (N_2934,N_2723,N_2780);
nor U2935 (N_2935,N_2711,N_2609);
and U2936 (N_2936,N_2795,N_2607);
or U2937 (N_2937,N_2676,N_2763);
and U2938 (N_2938,N_2746,N_2605);
and U2939 (N_2939,N_2760,N_2768);
and U2940 (N_2940,N_2703,N_2677);
nor U2941 (N_2941,N_2706,N_2624);
and U2942 (N_2942,N_2696,N_2781);
or U2943 (N_2943,N_2683,N_2651);
xnor U2944 (N_2944,N_2604,N_2738);
nand U2945 (N_2945,N_2641,N_2781);
or U2946 (N_2946,N_2632,N_2661);
nor U2947 (N_2947,N_2789,N_2648);
nand U2948 (N_2948,N_2641,N_2706);
or U2949 (N_2949,N_2768,N_2680);
or U2950 (N_2950,N_2747,N_2624);
or U2951 (N_2951,N_2601,N_2783);
nor U2952 (N_2952,N_2631,N_2704);
and U2953 (N_2953,N_2762,N_2721);
or U2954 (N_2954,N_2739,N_2650);
nand U2955 (N_2955,N_2605,N_2649);
or U2956 (N_2956,N_2710,N_2749);
xnor U2957 (N_2957,N_2793,N_2700);
xor U2958 (N_2958,N_2633,N_2714);
or U2959 (N_2959,N_2637,N_2739);
xnor U2960 (N_2960,N_2684,N_2642);
or U2961 (N_2961,N_2757,N_2767);
or U2962 (N_2962,N_2703,N_2794);
or U2963 (N_2963,N_2732,N_2769);
xor U2964 (N_2964,N_2641,N_2663);
nand U2965 (N_2965,N_2761,N_2657);
and U2966 (N_2966,N_2653,N_2737);
nand U2967 (N_2967,N_2687,N_2775);
and U2968 (N_2968,N_2685,N_2718);
nand U2969 (N_2969,N_2761,N_2791);
and U2970 (N_2970,N_2726,N_2627);
and U2971 (N_2971,N_2672,N_2697);
and U2972 (N_2972,N_2768,N_2754);
and U2973 (N_2973,N_2710,N_2727);
nand U2974 (N_2974,N_2665,N_2638);
and U2975 (N_2975,N_2614,N_2643);
nand U2976 (N_2976,N_2728,N_2655);
nand U2977 (N_2977,N_2749,N_2608);
nor U2978 (N_2978,N_2754,N_2727);
and U2979 (N_2979,N_2703,N_2603);
and U2980 (N_2980,N_2644,N_2711);
or U2981 (N_2981,N_2780,N_2777);
nor U2982 (N_2982,N_2617,N_2703);
nand U2983 (N_2983,N_2626,N_2745);
nor U2984 (N_2984,N_2649,N_2777);
and U2985 (N_2985,N_2709,N_2619);
xor U2986 (N_2986,N_2759,N_2775);
and U2987 (N_2987,N_2673,N_2621);
nand U2988 (N_2988,N_2664,N_2654);
and U2989 (N_2989,N_2640,N_2693);
and U2990 (N_2990,N_2621,N_2686);
nor U2991 (N_2991,N_2763,N_2772);
nor U2992 (N_2992,N_2766,N_2665);
xnor U2993 (N_2993,N_2736,N_2761);
and U2994 (N_2994,N_2753,N_2736);
nand U2995 (N_2995,N_2792,N_2683);
nor U2996 (N_2996,N_2605,N_2681);
nand U2997 (N_2997,N_2728,N_2690);
xnor U2998 (N_2998,N_2604,N_2600);
nor U2999 (N_2999,N_2673,N_2761);
nand UO_0 (O_0,N_2949,N_2998);
nand UO_1 (O_1,N_2941,N_2931);
nor UO_2 (O_2,N_2828,N_2809);
or UO_3 (O_3,N_2878,N_2895);
or UO_4 (O_4,N_2824,N_2842);
or UO_5 (O_5,N_2983,N_2839);
and UO_6 (O_6,N_2989,N_2913);
nand UO_7 (O_7,N_2830,N_2880);
or UO_8 (O_8,N_2819,N_2951);
and UO_9 (O_9,N_2822,N_2816);
nor UO_10 (O_10,N_2806,N_2827);
xor UO_11 (O_11,N_2897,N_2835);
and UO_12 (O_12,N_2975,N_2922);
and UO_13 (O_13,N_2920,N_2866);
nor UO_14 (O_14,N_2899,N_2890);
nand UO_15 (O_15,N_2982,N_2805);
nand UO_16 (O_16,N_2834,N_2848);
nor UO_17 (O_17,N_2843,N_2995);
or UO_18 (O_18,N_2971,N_2981);
and UO_19 (O_19,N_2801,N_2831);
and UO_20 (O_20,N_2921,N_2847);
nand UO_21 (O_21,N_2851,N_2962);
nor UO_22 (O_22,N_2905,N_2912);
or UO_23 (O_23,N_2810,N_2877);
or UO_24 (O_24,N_2940,N_2859);
and UO_25 (O_25,N_2825,N_2944);
nand UO_26 (O_26,N_2889,N_2803);
and UO_27 (O_27,N_2832,N_2891);
xnor UO_28 (O_28,N_2939,N_2856);
nor UO_29 (O_29,N_2833,N_2829);
xnor UO_30 (O_30,N_2928,N_2954);
and UO_31 (O_31,N_2838,N_2820);
and UO_32 (O_32,N_2894,N_2868);
nand UO_33 (O_33,N_2821,N_2896);
or UO_34 (O_34,N_2948,N_2858);
nand UO_35 (O_35,N_2898,N_2872);
xor UO_36 (O_36,N_2996,N_2903);
nand UO_37 (O_37,N_2811,N_2930);
nand UO_38 (O_38,N_2970,N_2867);
nor UO_39 (O_39,N_2815,N_2945);
nor UO_40 (O_40,N_2870,N_2906);
nor UO_41 (O_41,N_2955,N_2804);
and UO_42 (O_42,N_2862,N_2854);
and UO_43 (O_43,N_2884,N_2875);
or UO_44 (O_44,N_2850,N_2966);
and UO_45 (O_45,N_2909,N_2886);
nor UO_46 (O_46,N_2857,N_2873);
nor UO_47 (O_47,N_2882,N_2855);
nor UO_48 (O_48,N_2800,N_2911);
nor UO_49 (O_49,N_2865,N_2919);
nor UO_50 (O_50,N_2893,N_2938);
xnor UO_51 (O_51,N_2943,N_2910);
and UO_52 (O_52,N_2860,N_2874);
nor UO_53 (O_53,N_2991,N_2881);
or UO_54 (O_54,N_2925,N_2963);
xnor UO_55 (O_55,N_2826,N_2876);
or UO_56 (O_56,N_2802,N_2902);
nand UO_57 (O_57,N_2869,N_2888);
nor UO_58 (O_58,N_2953,N_2836);
and UO_59 (O_59,N_2993,N_2861);
or UO_60 (O_60,N_2946,N_2837);
and UO_61 (O_61,N_2932,N_2988);
xor UO_62 (O_62,N_2915,N_2957);
nor UO_63 (O_63,N_2845,N_2997);
nor UO_64 (O_64,N_2968,N_2918);
nand UO_65 (O_65,N_2960,N_2977);
xnor UO_66 (O_66,N_2952,N_2935);
nor UO_67 (O_67,N_2979,N_2947);
and UO_68 (O_68,N_2950,N_2958);
nand UO_69 (O_69,N_2907,N_2934);
and UO_70 (O_70,N_2841,N_2987);
and UO_71 (O_71,N_2901,N_2813);
nand UO_72 (O_72,N_2942,N_2863);
nor UO_73 (O_73,N_2818,N_2852);
or UO_74 (O_74,N_2900,N_2959);
nor UO_75 (O_75,N_2864,N_2929);
xnor UO_76 (O_76,N_2840,N_2853);
nand UO_77 (O_77,N_2926,N_2978);
and UO_78 (O_78,N_2904,N_2817);
or UO_79 (O_79,N_2917,N_2986);
xnor UO_80 (O_80,N_2933,N_2883);
nor UO_81 (O_81,N_2976,N_2980);
and UO_82 (O_82,N_2956,N_2936);
or UO_83 (O_83,N_2923,N_2846);
or UO_84 (O_84,N_2823,N_2892);
nand UO_85 (O_85,N_2812,N_2984);
nand UO_86 (O_86,N_2961,N_2908);
nor UO_87 (O_87,N_2814,N_2990);
or UO_88 (O_88,N_2973,N_2807);
nand UO_89 (O_89,N_2964,N_2844);
nand UO_90 (O_90,N_2924,N_2871);
nand UO_91 (O_91,N_2914,N_2879);
nand UO_92 (O_92,N_2937,N_2916);
nand UO_93 (O_93,N_2972,N_2885);
nor UO_94 (O_94,N_2985,N_2974);
and UO_95 (O_95,N_2927,N_2965);
nand UO_96 (O_96,N_2887,N_2994);
or UO_97 (O_97,N_2999,N_2808);
and UO_98 (O_98,N_2849,N_2992);
nand UO_99 (O_99,N_2969,N_2967);
nand UO_100 (O_100,N_2862,N_2975);
nand UO_101 (O_101,N_2967,N_2935);
and UO_102 (O_102,N_2950,N_2801);
nand UO_103 (O_103,N_2916,N_2864);
and UO_104 (O_104,N_2993,N_2804);
xnor UO_105 (O_105,N_2952,N_2987);
nand UO_106 (O_106,N_2921,N_2851);
nor UO_107 (O_107,N_2954,N_2867);
nor UO_108 (O_108,N_2988,N_2801);
or UO_109 (O_109,N_2884,N_2852);
nor UO_110 (O_110,N_2921,N_2936);
nor UO_111 (O_111,N_2897,N_2970);
or UO_112 (O_112,N_2824,N_2920);
nand UO_113 (O_113,N_2859,N_2872);
nor UO_114 (O_114,N_2866,N_2864);
nand UO_115 (O_115,N_2903,N_2989);
nor UO_116 (O_116,N_2955,N_2842);
nor UO_117 (O_117,N_2937,N_2867);
or UO_118 (O_118,N_2999,N_2850);
nand UO_119 (O_119,N_2997,N_2909);
or UO_120 (O_120,N_2803,N_2848);
nor UO_121 (O_121,N_2984,N_2896);
or UO_122 (O_122,N_2999,N_2826);
nor UO_123 (O_123,N_2882,N_2980);
and UO_124 (O_124,N_2911,N_2851);
or UO_125 (O_125,N_2905,N_2831);
nor UO_126 (O_126,N_2919,N_2967);
nor UO_127 (O_127,N_2823,N_2952);
nor UO_128 (O_128,N_2938,N_2984);
or UO_129 (O_129,N_2813,N_2909);
nor UO_130 (O_130,N_2989,N_2896);
or UO_131 (O_131,N_2858,N_2856);
or UO_132 (O_132,N_2986,N_2933);
nor UO_133 (O_133,N_2927,N_2848);
or UO_134 (O_134,N_2972,N_2998);
and UO_135 (O_135,N_2815,N_2996);
nor UO_136 (O_136,N_2853,N_2935);
or UO_137 (O_137,N_2901,N_2974);
xnor UO_138 (O_138,N_2848,N_2919);
xor UO_139 (O_139,N_2917,N_2935);
nor UO_140 (O_140,N_2985,N_2992);
nand UO_141 (O_141,N_2964,N_2999);
and UO_142 (O_142,N_2987,N_2810);
and UO_143 (O_143,N_2925,N_2873);
nor UO_144 (O_144,N_2983,N_2831);
and UO_145 (O_145,N_2901,N_2899);
and UO_146 (O_146,N_2842,N_2876);
or UO_147 (O_147,N_2958,N_2981);
nor UO_148 (O_148,N_2883,N_2981);
or UO_149 (O_149,N_2809,N_2865);
nor UO_150 (O_150,N_2993,N_2930);
nor UO_151 (O_151,N_2810,N_2949);
and UO_152 (O_152,N_2837,N_2820);
nor UO_153 (O_153,N_2905,N_2925);
and UO_154 (O_154,N_2870,N_2810);
and UO_155 (O_155,N_2988,N_2900);
and UO_156 (O_156,N_2865,N_2889);
or UO_157 (O_157,N_2887,N_2868);
nand UO_158 (O_158,N_2881,N_2948);
and UO_159 (O_159,N_2846,N_2905);
nand UO_160 (O_160,N_2853,N_2912);
nor UO_161 (O_161,N_2801,N_2892);
nand UO_162 (O_162,N_2923,N_2803);
xnor UO_163 (O_163,N_2850,N_2841);
and UO_164 (O_164,N_2935,N_2828);
xnor UO_165 (O_165,N_2984,N_2976);
or UO_166 (O_166,N_2800,N_2845);
and UO_167 (O_167,N_2962,N_2852);
and UO_168 (O_168,N_2848,N_2821);
xnor UO_169 (O_169,N_2858,N_2853);
nand UO_170 (O_170,N_2854,N_2898);
or UO_171 (O_171,N_2939,N_2983);
nor UO_172 (O_172,N_2995,N_2872);
xor UO_173 (O_173,N_2997,N_2889);
xor UO_174 (O_174,N_2965,N_2987);
or UO_175 (O_175,N_2823,N_2927);
nor UO_176 (O_176,N_2998,N_2928);
nand UO_177 (O_177,N_2845,N_2967);
nand UO_178 (O_178,N_2982,N_2868);
nor UO_179 (O_179,N_2896,N_2961);
or UO_180 (O_180,N_2904,N_2830);
nand UO_181 (O_181,N_2988,N_2852);
and UO_182 (O_182,N_2910,N_2800);
nand UO_183 (O_183,N_2864,N_2881);
nand UO_184 (O_184,N_2919,N_2820);
nand UO_185 (O_185,N_2884,N_2919);
nand UO_186 (O_186,N_2998,N_2863);
nor UO_187 (O_187,N_2846,N_2810);
and UO_188 (O_188,N_2893,N_2846);
or UO_189 (O_189,N_2980,N_2948);
or UO_190 (O_190,N_2918,N_2875);
nand UO_191 (O_191,N_2905,N_2948);
or UO_192 (O_192,N_2839,N_2979);
and UO_193 (O_193,N_2818,N_2967);
nor UO_194 (O_194,N_2901,N_2806);
nor UO_195 (O_195,N_2976,N_2943);
nand UO_196 (O_196,N_2889,N_2939);
or UO_197 (O_197,N_2938,N_2878);
nand UO_198 (O_198,N_2905,N_2909);
nor UO_199 (O_199,N_2925,N_2918);
or UO_200 (O_200,N_2869,N_2958);
nand UO_201 (O_201,N_2806,N_2911);
nor UO_202 (O_202,N_2958,N_2911);
nor UO_203 (O_203,N_2849,N_2805);
or UO_204 (O_204,N_2868,N_2803);
xnor UO_205 (O_205,N_2949,N_2957);
nand UO_206 (O_206,N_2988,N_2807);
nor UO_207 (O_207,N_2988,N_2830);
or UO_208 (O_208,N_2824,N_2865);
and UO_209 (O_209,N_2859,N_2809);
and UO_210 (O_210,N_2880,N_2956);
nor UO_211 (O_211,N_2827,N_2982);
nor UO_212 (O_212,N_2974,N_2892);
nand UO_213 (O_213,N_2858,N_2876);
nor UO_214 (O_214,N_2951,N_2886);
or UO_215 (O_215,N_2920,N_2881);
or UO_216 (O_216,N_2979,N_2939);
and UO_217 (O_217,N_2805,N_2947);
and UO_218 (O_218,N_2981,N_2908);
nand UO_219 (O_219,N_2841,N_2823);
nand UO_220 (O_220,N_2923,N_2834);
or UO_221 (O_221,N_2922,N_2878);
xor UO_222 (O_222,N_2986,N_2811);
nor UO_223 (O_223,N_2999,N_2864);
nand UO_224 (O_224,N_2825,N_2856);
nor UO_225 (O_225,N_2959,N_2989);
or UO_226 (O_226,N_2831,N_2968);
nor UO_227 (O_227,N_2898,N_2900);
nor UO_228 (O_228,N_2961,N_2903);
and UO_229 (O_229,N_2849,N_2821);
nor UO_230 (O_230,N_2813,N_2973);
xor UO_231 (O_231,N_2823,N_2935);
nor UO_232 (O_232,N_2860,N_2935);
or UO_233 (O_233,N_2890,N_2953);
or UO_234 (O_234,N_2876,N_2889);
nor UO_235 (O_235,N_2874,N_2836);
or UO_236 (O_236,N_2887,N_2965);
nor UO_237 (O_237,N_2935,N_2986);
nand UO_238 (O_238,N_2943,N_2984);
nor UO_239 (O_239,N_2801,N_2841);
or UO_240 (O_240,N_2835,N_2898);
nand UO_241 (O_241,N_2927,N_2973);
and UO_242 (O_242,N_2861,N_2822);
and UO_243 (O_243,N_2876,N_2979);
nand UO_244 (O_244,N_2925,N_2863);
nor UO_245 (O_245,N_2893,N_2981);
and UO_246 (O_246,N_2972,N_2895);
and UO_247 (O_247,N_2907,N_2935);
or UO_248 (O_248,N_2855,N_2897);
nand UO_249 (O_249,N_2866,N_2865);
or UO_250 (O_250,N_2839,N_2997);
or UO_251 (O_251,N_2922,N_2946);
nor UO_252 (O_252,N_2877,N_2889);
nand UO_253 (O_253,N_2907,N_2909);
or UO_254 (O_254,N_2846,N_2980);
nor UO_255 (O_255,N_2863,N_2888);
and UO_256 (O_256,N_2881,N_2834);
nand UO_257 (O_257,N_2803,N_2827);
or UO_258 (O_258,N_2866,N_2931);
or UO_259 (O_259,N_2843,N_2862);
and UO_260 (O_260,N_2880,N_2847);
nor UO_261 (O_261,N_2952,N_2945);
and UO_262 (O_262,N_2893,N_2877);
nand UO_263 (O_263,N_2882,N_2853);
or UO_264 (O_264,N_2994,N_2967);
and UO_265 (O_265,N_2937,N_2956);
and UO_266 (O_266,N_2953,N_2929);
nor UO_267 (O_267,N_2877,N_2834);
or UO_268 (O_268,N_2999,N_2848);
and UO_269 (O_269,N_2990,N_2957);
nor UO_270 (O_270,N_2884,N_2849);
or UO_271 (O_271,N_2993,N_2869);
and UO_272 (O_272,N_2885,N_2915);
xor UO_273 (O_273,N_2881,N_2923);
or UO_274 (O_274,N_2891,N_2993);
or UO_275 (O_275,N_2925,N_2992);
or UO_276 (O_276,N_2820,N_2804);
and UO_277 (O_277,N_2890,N_2837);
xnor UO_278 (O_278,N_2983,N_2878);
and UO_279 (O_279,N_2825,N_2948);
and UO_280 (O_280,N_2930,N_2857);
xnor UO_281 (O_281,N_2814,N_2878);
xnor UO_282 (O_282,N_2971,N_2859);
nor UO_283 (O_283,N_2909,N_2887);
nor UO_284 (O_284,N_2845,N_2915);
and UO_285 (O_285,N_2903,N_2950);
nor UO_286 (O_286,N_2943,N_2884);
or UO_287 (O_287,N_2964,N_2850);
nor UO_288 (O_288,N_2875,N_2996);
nand UO_289 (O_289,N_2978,N_2880);
nor UO_290 (O_290,N_2914,N_2834);
nand UO_291 (O_291,N_2858,N_2976);
nor UO_292 (O_292,N_2968,N_2868);
and UO_293 (O_293,N_2900,N_2935);
xor UO_294 (O_294,N_2895,N_2874);
nand UO_295 (O_295,N_2925,N_2881);
nor UO_296 (O_296,N_2883,N_2869);
nand UO_297 (O_297,N_2907,N_2916);
and UO_298 (O_298,N_2937,N_2823);
or UO_299 (O_299,N_2946,N_2881);
or UO_300 (O_300,N_2885,N_2963);
xnor UO_301 (O_301,N_2872,N_2874);
nand UO_302 (O_302,N_2854,N_2975);
or UO_303 (O_303,N_2894,N_2982);
nor UO_304 (O_304,N_2932,N_2862);
or UO_305 (O_305,N_2847,N_2825);
and UO_306 (O_306,N_2899,N_2817);
or UO_307 (O_307,N_2882,N_2927);
and UO_308 (O_308,N_2807,N_2997);
nand UO_309 (O_309,N_2874,N_2946);
nor UO_310 (O_310,N_2930,N_2870);
and UO_311 (O_311,N_2914,N_2955);
or UO_312 (O_312,N_2966,N_2881);
or UO_313 (O_313,N_2955,N_2891);
nand UO_314 (O_314,N_2850,N_2837);
nand UO_315 (O_315,N_2927,N_2936);
and UO_316 (O_316,N_2837,N_2914);
nor UO_317 (O_317,N_2807,N_2965);
and UO_318 (O_318,N_2912,N_2805);
nor UO_319 (O_319,N_2873,N_2949);
and UO_320 (O_320,N_2832,N_2977);
and UO_321 (O_321,N_2905,N_2893);
nand UO_322 (O_322,N_2963,N_2989);
and UO_323 (O_323,N_2972,N_2835);
or UO_324 (O_324,N_2806,N_2839);
nor UO_325 (O_325,N_2879,N_2962);
nor UO_326 (O_326,N_2828,N_2991);
xor UO_327 (O_327,N_2967,N_2983);
nand UO_328 (O_328,N_2868,N_2921);
xnor UO_329 (O_329,N_2892,N_2886);
nor UO_330 (O_330,N_2822,N_2874);
or UO_331 (O_331,N_2880,N_2865);
or UO_332 (O_332,N_2848,N_2853);
and UO_333 (O_333,N_2873,N_2814);
nand UO_334 (O_334,N_2901,N_2884);
or UO_335 (O_335,N_2939,N_2960);
nor UO_336 (O_336,N_2939,N_2825);
xnor UO_337 (O_337,N_2894,N_2888);
nand UO_338 (O_338,N_2947,N_2843);
nand UO_339 (O_339,N_2989,N_2916);
nand UO_340 (O_340,N_2985,N_2965);
xnor UO_341 (O_341,N_2865,N_2932);
nor UO_342 (O_342,N_2914,N_2818);
or UO_343 (O_343,N_2915,N_2807);
or UO_344 (O_344,N_2979,N_2855);
or UO_345 (O_345,N_2932,N_2986);
and UO_346 (O_346,N_2932,N_2992);
nand UO_347 (O_347,N_2830,N_2959);
xnor UO_348 (O_348,N_2882,N_2992);
nor UO_349 (O_349,N_2964,N_2823);
nor UO_350 (O_350,N_2998,N_2885);
xnor UO_351 (O_351,N_2966,N_2960);
nand UO_352 (O_352,N_2984,N_2989);
nand UO_353 (O_353,N_2915,N_2976);
nor UO_354 (O_354,N_2991,N_2846);
or UO_355 (O_355,N_2970,N_2918);
xnor UO_356 (O_356,N_2940,N_2849);
nor UO_357 (O_357,N_2881,N_2866);
and UO_358 (O_358,N_2920,N_2825);
nor UO_359 (O_359,N_2940,N_2910);
nor UO_360 (O_360,N_2893,N_2815);
nor UO_361 (O_361,N_2812,N_2928);
xnor UO_362 (O_362,N_2988,N_2946);
nor UO_363 (O_363,N_2986,N_2959);
or UO_364 (O_364,N_2860,N_2825);
or UO_365 (O_365,N_2993,N_2885);
or UO_366 (O_366,N_2922,N_2988);
xnor UO_367 (O_367,N_2934,N_2882);
nor UO_368 (O_368,N_2824,N_2843);
nand UO_369 (O_369,N_2972,N_2884);
nor UO_370 (O_370,N_2800,N_2924);
nand UO_371 (O_371,N_2992,N_2891);
xnor UO_372 (O_372,N_2892,N_2901);
nor UO_373 (O_373,N_2960,N_2982);
or UO_374 (O_374,N_2852,N_2810);
or UO_375 (O_375,N_2998,N_2800);
and UO_376 (O_376,N_2991,N_2955);
nor UO_377 (O_377,N_2845,N_2850);
nand UO_378 (O_378,N_2966,N_2945);
nor UO_379 (O_379,N_2858,N_2889);
nand UO_380 (O_380,N_2852,N_2849);
or UO_381 (O_381,N_2956,N_2879);
or UO_382 (O_382,N_2997,N_2987);
nor UO_383 (O_383,N_2868,N_2989);
xor UO_384 (O_384,N_2905,N_2873);
or UO_385 (O_385,N_2879,N_2822);
or UO_386 (O_386,N_2847,N_2889);
nor UO_387 (O_387,N_2860,N_2977);
or UO_388 (O_388,N_2832,N_2865);
xnor UO_389 (O_389,N_2971,N_2816);
xnor UO_390 (O_390,N_2984,N_2988);
nor UO_391 (O_391,N_2946,N_2987);
and UO_392 (O_392,N_2905,N_2961);
nand UO_393 (O_393,N_2887,N_2877);
xor UO_394 (O_394,N_2890,N_2932);
nand UO_395 (O_395,N_2995,N_2846);
nor UO_396 (O_396,N_2914,N_2929);
xor UO_397 (O_397,N_2926,N_2948);
or UO_398 (O_398,N_2938,N_2822);
nand UO_399 (O_399,N_2936,N_2812);
or UO_400 (O_400,N_2900,N_2953);
nand UO_401 (O_401,N_2929,N_2947);
nand UO_402 (O_402,N_2982,N_2845);
or UO_403 (O_403,N_2955,N_2852);
or UO_404 (O_404,N_2986,N_2877);
nand UO_405 (O_405,N_2835,N_2905);
or UO_406 (O_406,N_2978,N_2805);
nand UO_407 (O_407,N_2865,N_2939);
nor UO_408 (O_408,N_2924,N_2977);
or UO_409 (O_409,N_2942,N_2986);
nand UO_410 (O_410,N_2894,N_2934);
nand UO_411 (O_411,N_2805,N_2814);
and UO_412 (O_412,N_2882,N_2942);
or UO_413 (O_413,N_2897,N_2946);
or UO_414 (O_414,N_2939,N_2897);
and UO_415 (O_415,N_2820,N_2900);
or UO_416 (O_416,N_2914,N_2938);
nor UO_417 (O_417,N_2996,N_2952);
or UO_418 (O_418,N_2964,N_2994);
nor UO_419 (O_419,N_2989,N_2815);
and UO_420 (O_420,N_2897,N_2981);
nand UO_421 (O_421,N_2865,N_2984);
or UO_422 (O_422,N_2835,N_2971);
and UO_423 (O_423,N_2982,N_2811);
xor UO_424 (O_424,N_2882,N_2848);
nand UO_425 (O_425,N_2817,N_2869);
nor UO_426 (O_426,N_2847,N_2967);
and UO_427 (O_427,N_2850,N_2813);
nand UO_428 (O_428,N_2817,N_2872);
or UO_429 (O_429,N_2995,N_2817);
or UO_430 (O_430,N_2882,N_2973);
or UO_431 (O_431,N_2917,N_2882);
nor UO_432 (O_432,N_2935,N_2852);
nand UO_433 (O_433,N_2952,N_2965);
and UO_434 (O_434,N_2910,N_2915);
or UO_435 (O_435,N_2955,N_2826);
nor UO_436 (O_436,N_2875,N_2828);
or UO_437 (O_437,N_2925,N_2948);
and UO_438 (O_438,N_2988,N_2889);
and UO_439 (O_439,N_2969,N_2971);
or UO_440 (O_440,N_2854,N_2834);
nor UO_441 (O_441,N_2837,N_2996);
nand UO_442 (O_442,N_2828,N_2934);
nor UO_443 (O_443,N_2833,N_2922);
and UO_444 (O_444,N_2989,N_2828);
or UO_445 (O_445,N_2801,N_2922);
nor UO_446 (O_446,N_2840,N_2808);
or UO_447 (O_447,N_2814,N_2920);
or UO_448 (O_448,N_2984,N_2947);
nand UO_449 (O_449,N_2878,N_2931);
nand UO_450 (O_450,N_2868,N_2976);
xor UO_451 (O_451,N_2843,N_2900);
and UO_452 (O_452,N_2873,N_2803);
nand UO_453 (O_453,N_2807,N_2916);
nand UO_454 (O_454,N_2971,N_2953);
nor UO_455 (O_455,N_2940,N_2929);
nor UO_456 (O_456,N_2922,N_2890);
and UO_457 (O_457,N_2933,N_2975);
or UO_458 (O_458,N_2941,N_2942);
and UO_459 (O_459,N_2829,N_2923);
nor UO_460 (O_460,N_2894,N_2874);
or UO_461 (O_461,N_2895,N_2993);
or UO_462 (O_462,N_2908,N_2895);
nor UO_463 (O_463,N_2880,N_2813);
nand UO_464 (O_464,N_2927,N_2854);
nand UO_465 (O_465,N_2831,N_2981);
and UO_466 (O_466,N_2816,N_2979);
xor UO_467 (O_467,N_2843,N_2958);
nor UO_468 (O_468,N_2863,N_2948);
xor UO_469 (O_469,N_2948,N_2933);
or UO_470 (O_470,N_2990,N_2922);
and UO_471 (O_471,N_2819,N_2912);
and UO_472 (O_472,N_2930,N_2914);
nor UO_473 (O_473,N_2933,N_2832);
nor UO_474 (O_474,N_2887,N_2808);
nand UO_475 (O_475,N_2818,N_2896);
nor UO_476 (O_476,N_2835,N_2872);
or UO_477 (O_477,N_2845,N_2918);
and UO_478 (O_478,N_2887,N_2938);
nor UO_479 (O_479,N_2927,N_2833);
or UO_480 (O_480,N_2856,N_2966);
or UO_481 (O_481,N_2834,N_2853);
nor UO_482 (O_482,N_2939,N_2812);
nor UO_483 (O_483,N_2858,N_2994);
and UO_484 (O_484,N_2844,N_2915);
nor UO_485 (O_485,N_2831,N_2834);
nand UO_486 (O_486,N_2880,N_2846);
nand UO_487 (O_487,N_2994,N_2853);
or UO_488 (O_488,N_2943,N_2817);
and UO_489 (O_489,N_2849,N_2801);
xnor UO_490 (O_490,N_2847,N_2958);
nor UO_491 (O_491,N_2853,N_2851);
or UO_492 (O_492,N_2993,N_2876);
xnor UO_493 (O_493,N_2976,N_2842);
or UO_494 (O_494,N_2851,N_2825);
nor UO_495 (O_495,N_2830,N_2907);
xnor UO_496 (O_496,N_2913,N_2962);
and UO_497 (O_497,N_2969,N_2825);
or UO_498 (O_498,N_2921,N_2858);
or UO_499 (O_499,N_2947,N_2868);
endmodule