module basic_500_3000_500_30_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_413,In_120);
or U1 (N_1,In_16,In_71);
or U2 (N_2,In_7,In_282);
or U3 (N_3,In_254,In_290);
nand U4 (N_4,In_193,In_409);
or U5 (N_5,In_471,In_299);
nor U6 (N_6,In_434,In_258);
and U7 (N_7,In_363,In_489);
nand U8 (N_8,In_239,In_224);
xnor U9 (N_9,In_26,In_345);
or U10 (N_10,In_68,In_190);
nor U11 (N_11,In_12,In_165);
or U12 (N_12,In_463,In_72);
xnor U13 (N_13,In_469,In_244);
xnor U14 (N_14,In_129,In_40);
xnor U15 (N_15,In_309,In_252);
xnor U16 (N_16,In_86,In_454);
nor U17 (N_17,In_470,In_215);
xor U18 (N_18,In_20,In_283);
xnor U19 (N_19,In_286,In_81);
xor U20 (N_20,In_130,In_269);
nor U21 (N_21,In_343,In_268);
and U22 (N_22,In_274,In_55);
or U23 (N_23,In_101,In_160);
xor U24 (N_24,In_364,In_385);
xnor U25 (N_25,In_1,In_420);
nand U26 (N_26,In_14,In_361);
or U27 (N_27,In_419,In_310);
nor U28 (N_28,In_432,In_30);
nor U29 (N_29,In_125,In_455);
nand U30 (N_30,In_292,In_227);
or U31 (N_31,In_243,In_330);
or U32 (N_32,In_328,In_300);
or U33 (N_33,In_382,In_303);
nand U34 (N_34,In_146,In_387);
nand U35 (N_35,In_51,In_38);
nor U36 (N_36,In_184,In_76);
xor U37 (N_37,In_168,In_152);
xor U38 (N_38,In_459,In_34);
nor U39 (N_39,In_314,In_205);
or U40 (N_40,In_82,In_477);
nand U41 (N_41,In_226,In_186);
nand U42 (N_42,In_183,In_42);
xnor U43 (N_43,In_355,In_416);
xor U44 (N_44,In_480,In_497);
xnor U45 (N_45,In_85,In_230);
nand U46 (N_46,In_9,In_223);
and U47 (N_47,In_366,In_149);
nand U48 (N_48,In_144,In_36);
or U49 (N_49,In_496,In_5);
xor U50 (N_50,In_108,In_196);
nor U51 (N_51,In_93,In_114);
xnor U52 (N_52,In_62,In_450);
xnor U53 (N_53,In_327,In_429);
nor U54 (N_54,In_19,In_356);
nand U55 (N_55,In_468,In_380);
or U56 (N_56,In_123,In_231);
and U57 (N_57,In_358,In_192);
nand U58 (N_58,In_92,In_119);
or U59 (N_59,In_201,In_242);
nor U60 (N_60,In_465,In_462);
nand U61 (N_61,In_444,In_383);
nor U62 (N_62,In_272,In_482);
or U63 (N_63,In_381,In_112);
or U64 (N_64,In_460,In_445);
xor U65 (N_65,In_237,In_296);
nand U66 (N_66,In_372,In_298);
and U67 (N_67,In_393,In_411);
or U68 (N_68,In_344,In_334);
xor U69 (N_69,In_256,In_234);
xnor U70 (N_70,In_475,In_317);
nand U71 (N_71,In_287,In_261);
and U72 (N_72,In_294,In_247);
nand U73 (N_73,In_404,In_248);
and U74 (N_74,In_199,In_483);
nor U75 (N_75,In_246,In_403);
nor U76 (N_76,In_285,In_228);
nand U77 (N_77,In_349,In_306);
and U78 (N_78,In_388,In_464);
nand U79 (N_79,In_249,In_56);
and U80 (N_80,In_24,In_219);
nor U81 (N_81,In_21,In_316);
and U82 (N_82,In_453,In_80);
nand U83 (N_83,In_77,In_166);
nand U84 (N_84,In_105,In_426);
xor U85 (N_85,In_182,In_367);
or U86 (N_86,In_195,In_335);
nand U87 (N_87,In_422,In_238);
or U88 (N_88,In_473,In_425);
or U89 (N_89,In_25,In_360);
xor U90 (N_90,In_315,In_29);
or U91 (N_91,In_107,In_132);
nor U92 (N_92,In_63,In_297);
and U93 (N_93,In_479,In_438);
xnor U94 (N_94,In_69,In_275);
nand U95 (N_95,In_379,In_163);
nor U96 (N_96,In_188,In_67);
nor U97 (N_97,In_407,In_308);
nor U98 (N_98,In_245,In_441);
or U99 (N_99,In_378,In_135);
nor U100 (N_100,N_16,In_435);
or U101 (N_101,In_94,In_41);
xnor U102 (N_102,In_106,N_4);
or U103 (N_103,In_498,In_45);
and U104 (N_104,In_213,N_83);
and U105 (N_105,In_194,In_96);
nand U106 (N_106,In_395,In_78);
xnor U107 (N_107,In_347,In_39);
xnor U108 (N_108,In_37,N_92);
nor U109 (N_109,In_284,In_3);
nand U110 (N_110,In_52,In_126);
nor U111 (N_111,In_342,In_493);
or U112 (N_112,N_21,In_302);
or U113 (N_113,In_266,In_392);
nor U114 (N_114,In_97,In_439);
xnor U115 (N_115,N_66,In_4);
nor U116 (N_116,N_0,N_29);
or U117 (N_117,N_44,In_103);
and U118 (N_118,In_412,In_140);
nor U119 (N_119,In_336,N_1);
nor U120 (N_120,In_305,In_415);
xnor U121 (N_121,In_43,In_177);
xor U122 (N_122,In_447,In_353);
nand U123 (N_123,In_264,N_95);
and U124 (N_124,In_88,N_76);
nand U125 (N_125,In_136,In_484);
and U126 (N_126,In_157,In_117);
xor U127 (N_127,In_396,N_62);
and U128 (N_128,In_145,In_458);
and U129 (N_129,In_348,N_5);
xor U130 (N_130,In_331,In_49);
nand U131 (N_131,In_389,N_3);
nand U132 (N_132,N_89,In_318);
nor U133 (N_133,In_427,In_276);
nand U134 (N_134,In_250,In_321);
xor U135 (N_135,In_15,In_492);
xor U136 (N_136,In_398,In_390);
nor U137 (N_137,N_37,In_164);
nor U138 (N_138,In_373,In_148);
nor U139 (N_139,N_26,In_11);
nor U140 (N_140,N_35,N_7);
nand U141 (N_141,N_57,In_170);
nand U142 (N_142,In_28,In_394);
nor U143 (N_143,In_359,In_337);
nor U144 (N_144,In_323,N_71);
xnor U145 (N_145,In_70,N_24);
or U146 (N_146,In_210,In_255);
nand U147 (N_147,In_122,In_48);
nor U148 (N_148,In_433,In_259);
nor U149 (N_149,N_68,N_15);
nor U150 (N_150,N_53,In_84);
or U151 (N_151,In_240,In_257);
nand U152 (N_152,In_178,N_74);
xnor U153 (N_153,In_265,In_35);
and U154 (N_154,In_60,N_79);
or U155 (N_155,In_155,In_339);
xor U156 (N_156,In_325,In_467);
or U157 (N_157,In_279,In_357);
nand U158 (N_158,N_81,In_174);
nor U159 (N_159,In_446,N_22);
and U160 (N_160,In_365,N_49);
nand U161 (N_161,In_391,In_362);
and U162 (N_162,In_311,In_233);
and U163 (N_163,N_31,In_262);
xnor U164 (N_164,N_10,In_486);
xnor U165 (N_165,In_151,In_437);
or U166 (N_166,In_288,In_137);
or U167 (N_167,In_191,In_376);
and U168 (N_168,In_211,In_127);
nand U169 (N_169,In_291,In_495);
nand U170 (N_170,In_18,N_45);
xnor U171 (N_171,In_212,In_214);
xnor U172 (N_172,In_216,N_84);
nand U173 (N_173,N_19,In_6);
and U174 (N_174,In_64,In_457);
nor U175 (N_175,N_75,In_278);
and U176 (N_176,In_488,In_225);
xor U177 (N_177,In_222,N_36);
nor U178 (N_178,N_47,In_198);
xnor U179 (N_179,In_147,In_485);
or U180 (N_180,In_59,In_352);
nand U181 (N_181,In_273,In_100);
or U182 (N_182,N_42,In_65);
and U183 (N_183,N_51,In_430);
and U184 (N_184,N_97,In_370);
xnor U185 (N_185,N_88,In_143);
and U186 (N_186,In_478,In_124);
nand U187 (N_187,N_63,In_340);
nand U188 (N_188,In_270,N_70);
and U189 (N_189,N_56,In_402);
nand U190 (N_190,In_377,In_121);
nor U191 (N_191,In_424,In_253);
nor U192 (N_192,In_46,In_118);
nor U193 (N_193,In_281,N_86);
xor U194 (N_194,N_40,N_94);
nand U195 (N_195,In_161,In_456);
and U196 (N_196,In_171,In_58);
or U197 (N_197,In_418,N_77);
xor U198 (N_198,In_481,In_139);
nor U199 (N_199,In_267,In_154);
or U200 (N_200,N_99,In_301);
nor U201 (N_201,N_150,N_46);
or U202 (N_202,N_170,N_154);
and U203 (N_203,In_156,N_13);
nand U204 (N_204,In_312,N_91);
nor U205 (N_205,In_181,In_280);
and U206 (N_206,N_164,N_191);
nor U207 (N_207,N_136,N_184);
and U208 (N_208,N_162,N_102);
xor U209 (N_209,In_371,In_61);
xor U210 (N_210,In_490,In_134);
xnor U211 (N_211,In_260,N_157);
and U212 (N_212,N_106,In_241);
or U213 (N_213,In_289,N_145);
nor U214 (N_214,N_23,In_74);
nor U215 (N_215,In_406,In_87);
or U216 (N_216,N_65,In_142);
and U217 (N_217,N_137,In_113);
and U218 (N_218,In_319,N_188);
nand U219 (N_219,N_126,N_161);
nand U220 (N_220,In_197,In_13);
nor U221 (N_221,In_232,In_102);
or U222 (N_222,In_410,In_384);
and U223 (N_223,N_166,N_190);
xor U224 (N_224,In_448,In_354);
nand U225 (N_225,N_48,N_73);
nor U226 (N_226,In_22,N_138);
and U227 (N_227,N_110,In_436);
xor U228 (N_228,N_152,N_197);
or U229 (N_229,In_218,In_73);
and U230 (N_230,In_54,N_30);
and U231 (N_231,In_322,N_174);
xnor U232 (N_232,In_110,In_172);
and U233 (N_233,In_115,In_326);
xor U234 (N_234,In_79,N_39);
xnor U235 (N_235,N_171,N_167);
or U236 (N_236,N_125,In_99);
nand U237 (N_237,N_149,In_185);
and U238 (N_238,In_57,N_69);
and U239 (N_239,N_41,N_72);
or U240 (N_240,N_153,In_452);
nor U241 (N_241,N_59,N_130);
nor U242 (N_242,N_112,In_346);
nor U243 (N_243,In_324,N_193);
nand U244 (N_244,N_159,In_428);
nor U245 (N_245,N_176,N_93);
nor U246 (N_246,In_138,In_374);
or U247 (N_247,N_148,In_167);
nand U248 (N_248,N_105,In_31);
and U249 (N_249,In_451,N_121);
or U250 (N_250,In_350,N_158);
and U251 (N_251,In_83,In_200);
or U252 (N_252,In_189,N_101);
nand U253 (N_253,In_162,In_133);
xnor U254 (N_254,N_52,In_221);
or U255 (N_255,In_461,N_108);
xor U256 (N_256,In_408,In_338);
or U257 (N_257,In_442,N_128);
and U258 (N_258,N_18,N_151);
and U259 (N_259,N_109,N_169);
nor U260 (N_260,In_414,N_115);
nand U261 (N_261,N_165,N_180);
or U262 (N_262,N_198,In_229);
nand U263 (N_263,In_89,N_182);
xor U264 (N_264,In_369,N_133);
nand U265 (N_265,In_179,In_401);
and U266 (N_266,N_186,N_78);
xnor U267 (N_267,N_54,N_173);
or U268 (N_268,N_140,In_313);
nor U269 (N_269,N_9,In_368);
and U270 (N_270,In_175,In_440);
nand U271 (N_271,In_33,In_332);
nor U272 (N_272,N_196,N_17);
nor U273 (N_273,N_127,N_134);
and U274 (N_274,N_192,In_397);
or U275 (N_275,In_431,N_111);
or U276 (N_276,N_25,In_75);
nor U277 (N_277,N_124,In_0);
xor U278 (N_278,In_329,In_220);
nor U279 (N_279,In_47,N_55);
xnor U280 (N_280,In_405,In_251);
xor U281 (N_281,In_386,N_27);
nor U282 (N_282,In_8,N_123);
or U283 (N_283,In_443,N_147);
nor U284 (N_284,In_141,In_27);
and U285 (N_285,In_399,N_8);
xnor U286 (N_286,In_466,In_66);
nor U287 (N_287,In_499,In_217);
nor U288 (N_288,N_58,In_2);
xor U289 (N_289,In_304,N_143);
xnor U290 (N_290,N_172,N_61);
and U291 (N_291,In_491,In_202);
xor U292 (N_292,In_95,In_494);
xor U293 (N_293,N_122,In_487);
nor U294 (N_294,In_10,In_307);
and U295 (N_295,In_236,N_113);
and U296 (N_296,N_177,N_100);
or U297 (N_297,N_135,N_82);
xor U298 (N_298,In_104,N_6);
nor U299 (N_299,In_277,N_187);
xnor U300 (N_300,N_245,In_417);
or U301 (N_301,In_150,In_17);
nand U302 (N_302,N_265,In_90);
xor U303 (N_303,N_287,N_38);
xnor U304 (N_304,In_159,In_295);
nor U305 (N_305,N_264,In_449);
nor U306 (N_306,N_279,In_208);
and U307 (N_307,N_28,N_299);
nor U308 (N_308,N_199,N_118);
xor U309 (N_309,N_239,N_240);
or U310 (N_310,N_274,N_212);
or U311 (N_311,N_217,N_87);
and U312 (N_312,N_218,In_23);
nand U313 (N_313,In_204,In_169);
and U314 (N_314,N_211,In_421);
nor U315 (N_315,N_258,N_67);
nor U316 (N_316,N_243,N_98);
nor U317 (N_317,In_207,N_160);
nand U318 (N_318,N_60,N_263);
and U319 (N_319,N_248,N_298);
nand U320 (N_320,N_291,N_215);
nor U321 (N_321,In_320,N_293);
nor U322 (N_322,N_266,N_114);
nand U323 (N_323,In_109,In_271);
and U324 (N_324,N_288,N_11);
and U325 (N_325,N_33,N_282);
nor U326 (N_326,N_194,N_219);
or U327 (N_327,N_276,N_119);
and U328 (N_328,In_50,N_233);
nand U329 (N_329,N_281,N_270);
or U330 (N_330,N_247,N_117);
nor U331 (N_331,N_183,In_158);
or U332 (N_332,N_32,N_43);
xor U333 (N_333,N_246,N_203);
nor U334 (N_334,N_252,N_286);
nor U335 (N_335,N_210,N_256);
and U336 (N_336,N_257,N_242);
and U337 (N_337,N_12,In_351);
and U338 (N_338,In_235,N_216);
nand U339 (N_339,N_201,N_185);
or U340 (N_340,N_220,N_131);
and U341 (N_341,N_221,N_107);
or U342 (N_342,N_146,N_168);
nor U343 (N_343,N_280,N_120);
nand U344 (N_344,N_273,In_203);
or U345 (N_345,N_14,N_284);
nand U346 (N_346,N_64,N_231);
nand U347 (N_347,N_234,N_223);
xnor U348 (N_348,N_225,In_375);
nor U349 (N_349,N_235,In_187);
and U350 (N_350,N_260,N_238);
xor U351 (N_351,N_229,N_209);
and U352 (N_352,N_179,N_255);
xor U353 (N_353,N_278,N_296);
or U354 (N_354,In_474,N_132);
and U355 (N_355,N_129,N_141);
xnor U356 (N_356,N_163,N_272);
xor U357 (N_357,N_228,In_180);
nand U358 (N_358,In_153,N_207);
nor U359 (N_359,In_91,N_85);
nor U360 (N_360,N_295,N_214);
or U361 (N_361,In_293,N_253);
nor U362 (N_362,N_104,N_289);
nand U363 (N_363,N_181,N_222);
or U364 (N_364,In_341,N_230);
and U365 (N_365,N_269,In_423);
nor U366 (N_366,N_144,In_116);
xor U367 (N_367,N_202,In_400);
xnor U368 (N_368,N_50,N_80);
nor U369 (N_369,In_476,In_173);
nand U370 (N_370,N_156,N_290);
or U371 (N_371,N_277,N_189);
nor U372 (N_372,N_268,N_139);
nand U373 (N_373,In_176,N_116);
and U374 (N_374,N_208,N_2);
or U375 (N_375,N_250,N_226);
xor U376 (N_376,In_472,In_111);
and U377 (N_377,In_206,N_283);
or U378 (N_378,N_195,N_142);
nor U379 (N_379,In_32,N_178);
nor U380 (N_380,In_209,N_262);
nor U381 (N_381,In_53,N_254);
or U382 (N_382,N_213,In_128);
or U383 (N_383,N_204,N_241);
nor U384 (N_384,N_294,N_206);
xor U385 (N_385,N_224,N_251);
and U386 (N_386,N_200,In_131);
nor U387 (N_387,In_333,In_263);
and U388 (N_388,N_155,N_275);
xnor U389 (N_389,N_244,N_96);
nand U390 (N_390,N_232,In_98);
nand U391 (N_391,N_292,N_249);
nand U392 (N_392,N_237,N_285);
or U393 (N_393,N_90,N_236);
or U394 (N_394,N_175,N_205);
or U395 (N_395,N_34,N_20);
nor U396 (N_396,N_259,N_297);
nor U397 (N_397,N_261,N_271);
and U398 (N_398,N_103,N_267);
and U399 (N_399,In_44,N_227);
nand U400 (N_400,N_331,N_373);
nand U401 (N_401,N_388,N_310);
and U402 (N_402,N_366,N_303);
xor U403 (N_403,N_367,N_370);
xor U404 (N_404,N_372,N_332);
xor U405 (N_405,N_344,N_336);
or U406 (N_406,N_318,N_365);
nor U407 (N_407,N_325,N_322);
nor U408 (N_408,N_377,N_347);
and U409 (N_409,N_333,N_398);
nor U410 (N_410,N_345,N_371);
and U411 (N_411,N_330,N_312);
and U412 (N_412,N_384,N_328);
or U413 (N_413,N_306,N_391);
nor U414 (N_414,N_350,N_383);
nor U415 (N_415,N_315,N_349);
and U416 (N_416,N_357,N_339);
xor U417 (N_417,N_378,N_399);
nor U418 (N_418,N_319,N_343);
nand U419 (N_419,N_364,N_369);
nor U420 (N_420,N_393,N_341);
xnor U421 (N_421,N_316,N_351);
and U422 (N_422,N_385,N_368);
or U423 (N_423,N_394,N_327);
nor U424 (N_424,N_324,N_314);
nor U425 (N_425,N_362,N_342);
nand U426 (N_426,N_337,N_356);
xnor U427 (N_427,N_305,N_361);
and U428 (N_428,N_389,N_363);
nor U429 (N_429,N_334,N_374);
nor U430 (N_430,N_340,N_317);
nor U431 (N_431,N_321,N_307);
and U432 (N_432,N_375,N_386);
xor U433 (N_433,N_308,N_392);
and U434 (N_434,N_354,N_348);
and U435 (N_435,N_376,N_326);
xor U436 (N_436,N_358,N_320);
nand U437 (N_437,N_352,N_335);
nand U438 (N_438,N_311,N_380);
xnor U439 (N_439,N_397,N_379);
nor U440 (N_440,N_359,N_301);
xnor U441 (N_441,N_355,N_309);
or U442 (N_442,N_329,N_387);
nand U443 (N_443,N_353,N_302);
and U444 (N_444,N_346,N_395);
xnor U445 (N_445,N_390,N_381);
nor U446 (N_446,N_360,N_323);
xnor U447 (N_447,N_300,N_382);
nor U448 (N_448,N_338,N_304);
and U449 (N_449,N_313,N_396);
xor U450 (N_450,N_321,N_306);
xor U451 (N_451,N_324,N_395);
nor U452 (N_452,N_301,N_321);
nor U453 (N_453,N_387,N_372);
nand U454 (N_454,N_373,N_374);
or U455 (N_455,N_385,N_312);
xnor U456 (N_456,N_375,N_377);
and U457 (N_457,N_311,N_379);
xnor U458 (N_458,N_304,N_345);
nor U459 (N_459,N_388,N_326);
xnor U460 (N_460,N_386,N_352);
or U461 (N_461,N_369,N_314);
nand U462 (N_462,N_322,N_361);
or U463 (N_463,N_387,N_317);
nor U464 (N_464,N_321,N_325);
xnor U465 (N_465,N_305,N_339);
xor U466 (N_466,N_311,N_309);
nand U467 (N_467,N_331,N_302);
nand U468 (N_468,N_330,N_394);
or U469 (N_469,N_320,N_376);
xnor U470 (N_470,N_376,N_340);
nor U471 (N_471,N_390,N_329);
or U472 (N_472,N_314,N_379);
and U473 (N_473,N_363,N_307);
and U474 (N_474,N_390,N_313);
or U475 (N_475,N_322,N_365);
nor U476 (N_476,N_357,N_346);
nand U477 (N_477,N_315,N_301);
nor U478 (N_478,N_392,N_390);
or U479 (N_479,N_355,N_336);
and U480 (N_480,N_357,N_386);
xnor U481 (N_481,N_330,N_396);
nor U482 (N_482,N_320,N_328);
nor U483 (N_483,N_376,N_351);
and U484 (N_484,N_331,N_311);
nand U485 (N_485,N_374,N_340);
nand U486 (N_486,N_337,N_363);
nor U487 (N_487,N_307,N_324);
and U488 (N_488,N_347,N_363);
and U489 (N_489,N_389,N_375);
or U490 (N_490,N_321,N_320);
and U491 (N_491,N_350,N_339);
nor U492 (N_492,N_305,N_360);
and U493 (N_493,N_301,N_318);
or U494 (N_494,N_356,N_378);
and U495 (N_495,N_312,N_374);
and U496 (N_496,N_386,N_315);
and U497 (N_497,N_380,N_316);
or U498 (N_498,N_380,N_379);
nor U499 (N_499,N_396,N_382);
xor U500 (N_500,N_433,N_418);
or U501 (N_501,N_458,N_416);
xor U502 (N_502,N_457,N_404);
xor U503 (N_503,N_431,N_469);
nor U504 (N_504,N_405,N_437);
and U505 (N_505,N_406,N_407);
nand U506 (N_506,N_443,N_441);
nand U507 (N_507,N_483,N_460);
or U508 (N_508,N_446,N_475);
xor U509 (N_509,N_488,N_421);
nor U510 (N_510,N_449,N_444);
nand U511 (N_511,N_493,N_450);
or U512 (N_512,N_445,N_452);
xor U513 (N_513,N_456,N_497);
xor U514 (N_514,N_439,N_453);
xnor U515 (N_515,N_464,N_447);
and U516 (N_516,N_420,N_403);
and U517 (N_517,N_415,N_409);
xor U518 (N_518,N_468,N_473);
and U519 (N_519,N_498,N_417);
and U520 (N_520,N_489,N_459);
nand U521 (N_521,N_430,N_425);
and U522 (N_522,N_451,N_479);
and U523 (N_523,N_478,N_429);
xnor U524 (N_524,N_462,N_481);
and U525 (N_525,N_414,N_465);
nor U526 (N_526,N_484,N_486);
xor U527 (N_527,N_492,N_419);
xor U528 (N_528,N_472,N_435);
or U529 (N_529,N_455,N_423);
nor U530 (N_530,N_410,N_466);
and U531 (N_531,N_436,N_476);
or U532 (N_532,N_411,N_474);
or U533 (N_533,N_408,N_448);
xnor U534 (N_534,N_434,N_426);
xor U535 (N_535,N_495,N_470);
or U536 (N_536,N_482,N_477);
and U537 (N_537,N_487,N_412);
nand U538 (N_538,N_424,N_494);
nand U539 (N_539,N_402,N_499);
or U540 (N_540,N_467,N_471);
and U541 (N_541,N_496,N_440);
or U542 (N_542,N_400,N_428);
and U543 (N_543,N_485,N_442);
nor U544 (N_544,N_454,N_432);
or U545 (N_545,N_427,N_438);
nor U546 (N_546,N_422,N_463);
nand U547 (N_547,N_491,N_490);
nand U548 (N_548,N_461,N_413);
and U549 (N_549,N_401,N_480);
or U550 (N_550,N_467,N_416);
or U551 (N_551,N_477,N_408);
xnor U552 (N_552,N_466,N_405);
or U553 (N_553,N_445,N_433);
nor U554 (N_554,N_471,N_413);
and U555 (N_555,N_478,N_497);
or U556 (N_556,N_465,N_475);
xnor U557 (N_557,N_430,N_477);
nand U558 (N_558,N_489,N_485);
nor U559 (N_559,N_449,N_485);
and U560 (N_560,N_484,N_429);
xnor U561 (N_561,N_480,N_438);
nand U562 (N_562,N_476,N_457);
and U563 (N_563,N_420,N_485);
nand U564 (N_564,N_446,N_420);
nand U565 (N_565,N_433,N_425);
nand U566 (N_566,N_429,N_425);
nor U567 (N_567,N_444,N_470);
xnor U568 (N_568,N_426,N_414);
xor U569 (N_569,N_400,N_423);
nor U570 (N_570,N_441,N_476);
or U571 (N_571,N_413,N_497);
nor U572 (N_572,N_472,N_468);
or U573 (N_573,N_489,N_469);
or U574 (N_574,N_400,N_472);
xor U575 (N_575,N_437,N_431);
nor U576 (N_576,N_482,N_468);
or U577 (N_577,N_446,N_404);
nand U578 (N_578,N_434,N_473);
nor U579 (N_579,N_466,N_486);
nand U580 (N_580,N_482,N_409);
or U581 (N_581,N_400,N_486);
and U582 (N_582,N_451,N_449);
and U583 (N_583,N_428,N_457);
and U584 (N_584,N_400,N_415);
xnor U585 (N_585,N_458,N_480);
and U586 (N_586,N_489,N_411);
nor U587 (N_587,N_425,N_437);
nor U588 (N_588,N_400,N_439);
or U589 (N_589,N_466,N_433);
and U590 (N_590,N_491,N_409);
and U591 (N_591,N_433,N_408);
xnor U592 (N_592,N_438,N_451);
xor U593 (N_593,N_478,N_491);
nor U594 (N_594,N_443,N_425);
xnor U595 (N_595,N_464,N_402);
or U596 (N_596,N_440,N_457);
nor U597 (N_597,N_469,N_487);
xor U598 (N_598,N_481,N_410);
and U599 (N_599,N_462,N_468);
and U600 (N_600,N_581,N_532);
or U601 (N_601,N_548,N_531);
and U602 (N_602,N_511,N_563);
xor U603 (N_603,N_572,N_550);
nand U604 (N_604,N_533,N_544);
and U605 (N_605,N_569,N_504);
xnor U606 (N_606,N_552,N_509);
xnor U607 (N_607,N_502,N_521);
nor U608 (N_608,N_591,N_564);
nor U609 (N_609,N_534,N_561);
nand U610 (N_610,N_545,N_595);
nand U611 (N_611,N_556,N_589);
or U612 (N_612,N_524,N_537);
nand U613 (N_613,N_508,N_555);
nor U614 (N_614,N_528,N_599);
nand U615 (N_615,N_574,N_571);
or U616 (N_616,N_566,N_505);
or U617 (N_617,N_547,N_515);
or U618 (N_618,N_551,N_584);
or U619 (N_619,N_516,N_542);
or U620 (N_620,N_559,N_568);
xnor U621 (N_621,N_580,N_510);
xnor U622 (N_622,N_573,N_519);
nor U623 (N_623,N_562,N_553);
and U624 (N_624,N_575,N_565);
nand U625 (N_625,N_535,N_594);
nand U626 (N_626,N_525,N_549);
or U627 (N_627,N_507,N_530);
xnor U628 (N_628,N_520,N_543);
and U629 (N_629,N_592,N_597);
xnor U630 (N_630,N_598,N_513);
or U631 (N_631,N_588,N_567);
nand U632 (N_632,N_546,N_576);
nand U633 (N_633,N_512,N_503);
or U634 (N_634,N_585,N_529);
or U635 (N_635,N_514,N_560);
or U636 (N_636,N_554,N_570);
nor U637 (N_637,N_577,N_527);
nor U638 (N_638,N_583,N_500);
or U639 (N_639,N_501,N_523);
and U640 (N_640,N_558,N_540);
xor U641 (N_641,N_582,N_587);
nor U642 (N_642,N_593,N_538);
or U643 (N_643,N_596,N_586);
and U644 (N_644,N_536,N_539);
and U645 (N_645,N_518,N_506);
or U646 (N_646,N_578,N_541);
nor U647 (N_647,N_522,N_590);
nor U648 (N_648,N_557,N_579);
nor U649 (N_649,N_526,N_517);
or U650 (N_650,N_590,N_596);
xnor U651 (N_651,N_558,N_593);
nor U652 (N_652,N_564,N_506);
or U653 (N_653,N_525,N_541);
and U654 (N_654,N_580,N_511);
nand U655 (N_655,N_523,N_506);
nor U656 (N_656,N_551,N_562);
nand U657 (N_657,N_559,N_545);
xnor U658 (N_658,N_561,N_514);
xor U659 (N_659,N_555,N_551);
or U660 (N_660,N_524,N_585);
nand U661 (N_661,N_556,N_549);
nand U662 (N_662,N_537,N_528);
nand U663 (N_663,N_572,N_583);
nand U664 (N_664,N_584,N_577);
or U665 (N_665,N_534,N_543);
and U666 (N_666,N_555,N_587);
and U667 (N_667,N_585,N_586);
nor U668 (N_668,N_523,N_502);
or U669 (N_669,N_586,N_568);
or U670 (N_670,N_511,N_537);
and U671 (N_671,N_582,N_589);
and U672 (N_672,N_548,N_501);
nor U673 (N_673,N_507,N_567);
nor U674 (N_674,N_598,N_592);
or U675 (N_675,N_509,N_538);
or U676 (N_676,N_535,N_597);
nand U677 (N_677,N_506,N_560);
nand U678 (N_678,N_547,N_554);
nor U679 (N_679,N_585,N_582);
nor U680 (N_680,N_500,N_547);
and U681 (N_681,N_539,N_548);
xnor U682 (N_682,N_522,N_551);
xnor U683 (N_683,N_573,N_501);
nor U684 (N_684,N_594,N_516);
and U685 (N_685,N_503,N_597);
nand U686 (N_686,N_515,N_557);
or U687 (N_687,N_504,N_529);
and U688 (N_688,N_527,N_587);
or U689 (N_689,N_589,N_500);
xor U690 (N_690,N_598,N_523);
nand U691 (N_691,N_545,N_553);
xor U692 (N_692,N_525,N_598);
or U693 (N_693,N_509,N_562);
xor U694 (N_694,N_590,N_595);
nor U695 (N_695,N_515,N_541);
or U696 (N_696,N_524,N_559);
and U697 (N_697,N_583,N_589);
nor U698 (N_698,N_500,N_522);
nand U699 (N_699,N_599,N_534);
or U700 (N_700,N_675,N_660);
nand U701 (N_701,N_679,N_621);
xor U702 (N_702,N_619,N_611);
or U703 (N_703,N_656,N_642);
nor U704 (N_704,N_681,N_652);
or U705 (N_705,N_622,N_643);
and U706 (N_706,N_641,N_682);
nor U707 (N_707,N_620,N_699);
and U708 (N_708,N_655,N_683);
xnor U709 (N_709,N_697,N_646);
nor U710 (N_710,N_669,N_657);
and U711 (N_711,N_670,N_626);
nand U712 (N_712,N_639,N_605);
or U713 (N_713,N_618,N_674);
or U714 (N_714,N_654,N_609);
and U715 (N_715,N_623,N_671);
and U716 (N_716,N_695,N_616);
or U717 (N_717,N_661,N_608);
or U718 (N_718,N_628,N_696);
nand U719 (N_719,N_668,N_647);
or U720 (N_720,N_630,N_662);
and U721 (N_721,N_612,N_613);
nand U722 (N_722,N_676,N_680);
nand U723 (N_723,N_601,N_645);
nor U724 (N_724,N_610,N_667);
xnor U725 (N_725,N_625,N_694);
nor U726 (N_726,N_693,N_690);
nand U727 (N_727,N_658,N_666);
xor U728 (N_728,N_673,N_637);
or U729 (N_729,N_692,N_603);
nand U730 (N_730,N_672,N_677);
or U731 (N_731,N_698,N_653);
and U732 (N_732,N_615,N_633);
and U733 (N_733,N_691,N_665);
and U734 (N_734,N_624,N_600);
and U735 (N_735,N_664,N_689);
or U736 (N_736,N_685,N_686);
xnor U737 (N_737,N_687,N_604);
nand U738 (N_738,N_632,N_678);
xor U739 (N_739,N_617,N_684);
nand U740 (N_740,N_631,N_659);
nand U741 (N_741,N_634,N_638);
xnor U742 (N_742,N_636,N_651);
xnor U743 (N_743,N_649,N_644);
nor U744 (N_744,N_640,N_602);
and U745 (N_745,N_607,N_606);
nor U746 (N_746,N_650,N_614);
or U747 (N_747,N_627,N_688);
and U748 (N_748,N_629,N_663);
nor U749 (N_749,N_648,N_635);
xor U750 (N_750,N_602,N_685);
xor U751 (N_751,N_644,N_602);
nor U752 (N_752,N_639,N_667);
xor U753 (N_753,N_676,N_695);
nand U754 (N_754,N_680,N_645);
xnor U755 (N_755,N_612,N_637);
or U756 (N_756,N_623,N_694);
xnor U757 (N_757,N_610,N_682);
or U758 (N_758,N_629,N_690);
xor U759 (N_759,N_633,N_653);
xnor U760 (N_760,N_609,N_680);
or U761 (N_761,N_685,N_676);
nor U762 (N_762,N_636,N_654);
and U763 (N_763,N_613,N_693);
and U764 (N_764,N_646,N_616);
or U765 (N_765,N_618,N_621);
and U766 (N_766,N_633,N_691);
nor U767 (N_767,N_632,N_616);
or U768 (N_768,N_644,N_673);
or U769 (N_769,N_602,N_652);
xor U770 (N_770,N_636,N_606);
or U771 (N_771,N_663,N_672);
nand U772 (N_772,N_675,N_690);
and U773 (N_773,N_644,N_636);
nand U774 (N_774,N_622,N_657);
nor U775 (N_775,N_656,N_611);
nand U776 (N_776,N_614,N_676);
xnor U777 (N_777,N_649,N_647);
nor U778 (N_778,N_614,N_669);
and U779 (N_779,N_627,N_672);
nor U780 (N_780,N_672,N_675);
nor U781 (N_781,N_697,N_612);
or U782 (N_782,N_695,N_625);
xor U783 (N_783,N_654,N_601);
nor U784 (N_784,N_681,N_672);
nor U785 (N_785,N_637,N_663);
and U786 (N_786,N_698,N_662);
nor U787 (N_787,N_641,N_652);
nand U788 (N_788,N_633,N_686);
nand U789 (N_789,N_656,N_622);
xnor U790 (N_790,N_657,N_659);
nand U791 (N_791,N_670,N_622);
or U792 (N_792,N_698,N_630);
or U793 (N_793,N_647,N_678);
or U794 (N_794,N_639,N_673);
nand U795 (N_795,N_664,N_609);
nand U796 (N_796,N_637,N_651);
and U797 (N_797,N_663,N_623);
xor U798 (N_798,N_649,N_688);
or U799 (N_799,N_643,N_665);
and U800 (N_800,N_776,N_761);
nor U801 (N_801,N_740,N_748);
and U802 (N_802,N_736,N_779);
and U803 (N_803,N_770,N_771);
xor U804 (N_804,N_723,N_726);
xor U805 (N_805,N_714,N_793);
xor U806 (N_806,N_700,N_715);
nand U807 (N_807,N_737,N_719);
nor U808 (N_808,N_759,N_769);
and U809 (N_809,N_787,N_735);
nand U810 (N_810,N_727,N_754);
xor U811 (N_811,N_745,N_774);
nor U812 (N_812,N_794,N_712);
nor U813 (N_813,N_733,N_799);
xnor U814 (N_814,N_717,N_706);
xnor U815 (N_815,N_742,N_705);
nor U816 (N_816,N_708,N_729);
and U817 (N_817,N_757,N_724);
xnor U818 (N_818,N_707,N_743);
or U819 (N_819,N_789,N_752);
nor U820 (N_820,N_788,N_734);
and U821 (N_821,N_790,N_775);
nor U822 (N_822,N_744,N_751);
nor U823 (N_823,N_750,N_728);
nand U824 (N_824,N_763,N_746);
nand U825 (N_825,N_755,N_782);
nor U826 (N_826,N_773,N_731);
nand U827 (N_827,N_718,N_749);
and U828 (N_828,N_783,N_768);
nand U829 (N_829,N_756,N_765);
xnor U830 (N_830,N_777,N_795);
and U831 (N_831,N_732,N_710);
nor U832 (N_832,N_781,N_797);
or U833 (N_833,N_762,N_720);
nand U834 (N_834,N_709,N_753);
nor U835 (N_835,N_716,N_703);
nand U836 (N_836,N_791,N_796);
and U837 (N_837,N_798,N_760);
nand U838 (N_838,N_741,N_713);
and U839 (N_839,N_778,N_764);
or U840 (N_840,N_767,N_738);
nand U841 (N_841,N_725,N_784);
or U842 (N_842,N_747,N_780);
or U843 (N_843,N_772,N_711);
or U844 (N_844,N_721,N_792);
and U845 (N_845,N_730,N_766);
xnor U846 (N_846,N_702,N_758);
or U847 (N_847,N_704,N_786);
and U848 (N_848,N_701,N_739);
nor U849 (N_849,N_722,N_785);
nor U850 (N_850,N_793,N_733);
xor U851 (N_851,N_770,N_755);
nor U852 (N_852,N_738,N_779);
xnor U853 (N_853,N_790,N_784);
nor U854 (N_854,N_788,N_735);
xnor U855 (N_855,N_711,N_770);
or U856 (N_856,N_760,N_755);
nand U857 (N_857,N_772,N_740);
nand U858 (N_858,N_749,N_717);
xor U859 (N_859,N_766,N_740);
nor U860 (N_860,N_777,N_701);
nor U861 (N_861,N_707,N_776);
nand U862 (N_862,N_796,N_716);
and U863 (N_863,N_717,N_712);
and U864 (N_864,N_732,N_761);
nand U865 (N_865,N_738,N_791);
nand U866 (N_866,N_742,N_737);
nor U867 (N_867,N_731,N_794);
and U868 (N_868,N_741,N_770);
or U869 (N_869,N_715,N_714);
or U870 (N_870,N_739,N_768);
or U871 (N_871,N_749,N_774);
xnor U872 (N_872,N_753,N_742);
and U873 (N_873,N_759,N_753);
or U874 (N_874,N_734,N_765);
nand U875 (N_875,N_737,N_749);
nand U876 (N_876,N_782,N_767);
xnor U877 (N_877,N_786,N_708);
nor U878 (N_878,N_724,N_765);
nor U879 (N_879,N_796,N_778);
nand U880 (N_880,N_743,N_728);
nor U881 (N_881,N_798,N_705);
and U882 (N_882,N_793,N_722);
xor U883 (N_883,N_722,N_712);
or U884 (N_884,N_704,N_700);
nor U885 (N_885,N_709,N_769);
nand U886 (N_886,N_775,N_703);
or U887 (N_887,N_795,N_711);
nor U888 (N_888,N_761,N_703);
or U889 (N_889,N_722,N_748);
nor U890 (N_890,N_706,N_738);
xor U891 (N_891,N_796,N_792);
or U892 (N_892,N_789,N_775);
nor U893 (N_893,N_760,N_767);
xnor U894 (N_894,N_733,N_769);
nand U895 (N_895,N_721,N_742);
and U896 (N_896,N_750,N_709);
and U897 (N_897,N_730,N_700);
or U898 (N_898,N_710,N_778);
xor U899 (N_899,N_708,N_776);
nand U900 (N_900,N_856,N_868);
or U901 (N_901,N_851,N_878);
or U902 (N_902,N_838,N_847);
nor U903 (N_903,N_881,N_870);
or U904 (N_904,N_840,N_846);
and U905 (N_905,N_895,N_875);
nand U906 (N_906,N_811,N_828);
or U907 (N_907,N_869,N_820);
or U908 (N_908,N_844,N_810);
and U909 (N_909,N_864,N_843);
and U910 (N_910,N_830,N_888);
nor U911 (N_911,N_836,N_824);
and U912 (N_912,N_800,N_803);
nor U913 (N_913,N_812,N_892);
xnor U914 (N_914,N_802,N_852);
nor U915 (N_915,N_872,N_866);
nand U916 (N_916,N_849,N_808);
and U917 (N_917,N_816,N_841);
nor U918 (N_918,N_890,N_822);
nand U919 (N_919,N_814,N_805);
nor U920 (N_920,N_880,N_845);
xnor U921 (N_921,N_882,N_877);
and U922 (N_922,N_813,N_891);
xnor U923 (N_923,N_853,N_848);
or U924 (N_924,N_819,N_809);
or U925 (N_925,N_860,N_807);
and U926 (N_926,N_818,N_885);
or U927 (N_927,N_894,N_835);
and U928 (N_928,N_893,N_873);
and U929 (N_929,N_861,N_874);
xor U930 (N_930,N_834,N_823);
nor U931 (N_931,N_829,N_883);
xor U932 (N_932,N_837,N_821);
nand U933 (N_933,N_876,N_865);
xor U934 (N_934,N_867,N_871);
nand U935 (N_935,N_879,N_826);
or U936 (N_936,N_898,N_896);
and U937 (N_937,N_850,N_858);
and U938 (N_938,N_839,N_833);
nand U939 (N_939,N_827,N_815);
nor U940 (N_940,N_831,N_859);
and U941 (N_941,N_801,N_854);
nand U942 (N_942,N_884,N_825);
xor U943 (N_943,N_817,N_842);
nand U944 (N_944,N_855,N_804);
nor U945 (N_945,N_899,N_832);
and U946 (N_946,N_897,N_806);
nor U947 (N_947,N_886,N_863);
nor U948 (N_948,N_887,N_889);
nand U949 (N_949,N_862,N_857);
nor U950 (N_950,N_874,N_801);
xnor U951 (N_951,N_819,N_815);
or U952 (N_952,N_852,N_820);
nor U953 (N_953,N_823,N_872);
xnor U954 (N_954,N_896,N_837);
or U955 (N_955,N_882,N_856);
nor U956 (N_956,N_823,N_840);
xnor U957 (N_957,N_873,N_867);
nand U958 (N_958,N_876,N_843);
xor U959 (N_959,N_808,N_837);
nand U960 (N_960,N_897,N_869);
nand U961 (N_961,N_849,N_837);
nor U962 (N_962,N_879,N_863);
nand U963 (N_963,N_895,N_864);
or U964 (N_964,N_850,N_811);
and U965 (N_965,N_875,N_801);
or U966 (N_966,N_816,N_891);
xnor U967 (N_967,N_848,N_846);
and U968 (N_968,N_800,N_809);
and U969 (N_969,N_863,N_865);
nor U970 (N_970,N_810,N_881);
nor U971 (N_971,N_827,N_845);
and U972 (N_972,N_833,N_803);
nor U973 (N_973,N_894,N_895);
nor U974 (N_974,N_894,N_870);
nor U975 (N_975,N_894,N_829);
nand U976 (N_976,N_854,N_893);
xor U977 (N_977,N_841,N_882);
xnor U978 (N_978,N_824,N_862);
or U979 (N_979,N_866,N_809);
nand U980 (N_980,N_807,N_867);
nand U981 (N_981,N_831,N_852);
and U982 (N_982,N_815,N_841);
and U983 (N_983,N_831,N_819);
and U984 (N_984,N_894,N_890);
xnor U985 (N_985,N_812,N_849);
and U986 (N_986,N_823,N_882);
nand U987 (N_987,N_824,N_820);
and U988 (N_988,N_897,N_868);
or U989 (N_989,N_878,N_865);
xnor U990 (N_990,N_824,N_801);
xnor U991 (N_991,N_837,N_856);
or U992 (N_992,N_887,N_843);
or U993 (N_993,N_824,N_800);
and U994 (N_994,N_843,N_899);
nor U995 (N_995,N_887,N_855);
nand U996 (N_996,N_828,N_853);
nor U997 (N_997,N_805,N_830);
nand U998 (N_998,N_868,N_857);
or U999 (N_999,N_841,N_806);
and U1000 (N_1000,N_909,N_900);
nor U1001 (N_1001,N_910,N_916);
xor U1002 (N_1002,N_968,N_906);
nand U1003 (N_1003,N_964,N_912);
or U1004 (N_1004,N_911,N_932);
xor U1005 (N_1005,N_908,N_933);
and U1006 (N_1006,N_904,N_928);
nor U1007 (N_1007,N_953,N_944);
and U1008 (N_1008,N_957,N_979);
or U1009 (N_1009,N_925,N_959);
and U1010 (N_1010,N_978,N_951);
and U1011 (N_1011,N_982,N_935);
and U1012 (N_1012,N_965,N_969);
and U1013 (N_1013,N_994,N_989);
xor U1014 (N_1014,N_983,N_998);
or U1015 (N_1015,N_960,N_922);
and U1016 (N_1016,N_946,N_981);
xnor U1017 (N_1017,N_921,N_923);
nand U1018 (N_1018,N_966,N_941);
nand U1019 (N_1019,N_976,N_992);
and U1020 (N_1020,N_929,N_926);
nand U1021 (N_1021,N_985,N_917);
or U1022 (N_1022,N_984,N_938);
nor U1023 (N_1023,N_963,N_987);
or U1024 (N_1024,N_939,N_940);
nor U1025 (N_1025,N_972,N_996);
xor U1026 (N_1026,N_991,N_943);
nand U1027 (N_1027,N_924,N_902);
or U1028 (N_1028,N_915,N_927);
and U1029 (N_1029,N_970,N_950);
or U1030 (N_1030,N_988,N_967);
xnor U1031 (N_1031,N_920,N_945);
nand U1032 (N_1032,N_997,N_993);
nor U1033 (N_1033,N_971,N_942);
xor U1034 (N_1034,N_974,N_936);
nor U1035 (N_1035,N_973,N_977);
and U1036 (N_1036,N_952,N_956);
or U1037 (N_1037,N_961,N_930);
and U1038 (N_1038,N_901,N_958);
and U1039 (N_1039,N_919,N_995);
nor U1040 (N_1040,N_949,N_948);
nor U1041 (N_1041,N_955,N_937);
or U1042 (N_1042,N_990,N_931);
and U1043 (N_1043,N_913,N_962);
nor U1044 (N_1044,N_954,N_914);
and U1045 (N_1045,N_934,N_947);
or U1046 (N_1046,N_986,N_903);
nor U1047 (N_1047,N_999,N_918);
xnor U1048 (N_1048,N_975,N_905);
nand U1049 (N_1049,N_907,N_980);
nand U1050 (N_1050,N_956,N_927);
and U1051 (N_1051,N_912,N_956);
xnor U1052 (N_1052,N_932,N_976);
or U1053 (N_1053,N_995,N_999);
nor U1054 (N_1054,N_986,N_908);
and U1055 (N_1055,N_945,N_978);
xor U1056 (N_1056,N_944,N_975);
and U1057 (N_1057,N_991,N_915);
or U1058 (N_1058,N_985,N_920);
nor U1059 (N_1059,N_971,N_986);
nand U1060 (N_1060,N_928,N_980);
and U1061 (N_1061,N_927,N_953);
nand U1062 (N_1062,N_950,N_909);
and U1063 (N_1063,N_982,N_998);
or U1064 (N_1064,N_981,N_977);
or U1065 (N_1065,N_983,N_996);
or U1066 (N_1066,N_911,N_971);
xor U1067 (N_1067,N_967,N_912);
nand U1068 (N_1068,N_999,N_974);
or U1069 (N_1069,N_933,N_930);
nor U1070 (N_1070,N_983,N_902);
or U1071 (N_1071,N_946,N_907);
nand U1072 (N_1072,N_983,N_917);
and U1073 (N_1073,N_999,N_925);
xnor U1074 (N_1074,N_903,N_981);
or U1075 (N_1075,N_945,N_981);
xor U1076 (N_1076,N_952,N_980);
and U1077 (N_1077,N_913,N_935);
nand U1078 (N_1078,N_941,N_985);
nor U1079 (N_1079,N_998,N_928);
and U1080 (N_1080,N_935,N_926);
and U1081 (N_1081,N_922,N_972);
or U1082 (N_1082,N_931,N_995);
nand U1083 (N_1083,N_967,N_940);
or U1084 (N_1084,N_928,N_939);
nor U1085 (N_1085,N_966,N_931);
nand U1086 (N_1086,N_920,N_926);
nor U1087 (N_1087,N_977,N_947);
or U1088 (N_1088,N_981,N_987);
or U1089 (N_1089,N_986,N_989);
xor U1090 (N_1090,N_918,N_962);
nor U1091 (N_1091,N_984,N_961);
nor U1092 (N_1092,N_909,N_970);
nand U1093 (N_1093,N_987,N_933);
nand U1094 (N_1094,N_913,N_989);
nor U1095 (N_1095,N_939,N_925);
xnor U1096 (N_1096,N_958,N_917);
xnor U1097 (N_1097,N_975,N_991);
and U1098 (N_1098,N_983,N_997);
nand U1099 (N_1099,N_989,N_976);
nor U1100 (N_1100,N_1086,N_1088);
nand U1101 (N_1101,N_1091,N_1053);
xnor U1102 (N_1102,N_1098,N_1030);
nor U1103 (N_1103,N_1023,N_1095);
nor U1104 (N_1104,N_1071,N_1032);
nor U1105 (N_1105,N_1037,N_1009);
or U1106 (N_1106,N_1072,N_1094);
nor U1107 (N_1107,N_1007,N_1042);
xor U1108 (N_1108,N_1001,N_1074);
nand U1109 (N_1109,N_1063,N_1038);
or U1110 (N_1110,N_1041,N_1051);
nor U1111 (N_1111,N_1093,N_1054);
nand U1112 (N_1112,N_1097,N_1073);
xor U1113 (N_1113,N_1021,N_1022);
nand U1114 (N_1114,N_1067,N_1016);
nor U1115 (N_1115,N_1092,N_1004);
or U1116 (N_1116,N_1084,N_1031);
nand U1117 (N_1117,N_1026,N_1078);
xnor U1118 (N_1118,N_1024,N_1096);
nor U1119 (N_1119,N_1005,N_1058);
and U1120 (N_1120,N_1008,N_1057);
xor U1121 (N_1121,N_1002,N_1028);
nand U1122 (N_1122,N_1066,N_1013);
nand U1123 (N_1123,N_1003,N_1059);
xnor U1124 (N_1124,N_1044,N_1046);
and U1125 (N_1125,N_1012,N_1089);
or U1126 (N_1126,N_1061,N_1048);
xor U1127 (N_1127,N_1077,N_1060);
xor U1128 (N_1128,N_1018,N_1019);
nand U1129 (N_1129,N_1040,N_1015);
and U1130 (N_1130,N_1085,N_1027);
nor U1131 (N_1131,N_1025,N_1070);
nand U1132 (N_1132,N_1000,N_1056);
xor U1133 (N_1133,N_1049,N_1082);
nor U1134 (N_1134,N_1052,N_1029);
nor U1135 (N_1135,N_1075,N_1010);
or U1136 (N_1136,N_1087,N_1068);
and U1137 (N_1137,N_1081,N_1069);
xor U1138 (N_1138,N_1065,N_1090);
nor U1139 (N_1139,N_1099,N_1006);
or U1140 (N_1140,N_1045,N_1020);
xnor U1141 (N_1141,N_1014,N_1033);
and U1142 (N_1142,N_1039,N_1050);
nor U1143 (N_1143,N_1062,N_1079);
nor U1144 (N_1144,N_1076,N_1080);
or U1145 (N_1145,N_1036,N_1055);
xor U1146 (N_1146,N_1064,N_1047);
xor U1147 (N_1147,N_1043,N_1035);
and U1148 (N_1148,N_1017,N_1083);
xnor U1149 (N_1149,N_1034,N_1011);
xor U1150 (N_1150,N_1037,N_1069);
xnor U1151 (N_1151,N_1075,N_1098);
and U1152 (N_1152,N_1044,N_1065);
and U1153 (N_1153,N_1054,N_1099);
and U1154 (N_1154,N_1056,N_1043);
nand U1155 (N_1155,N_1014,N_1030);
nor U1156 (N_1156,N_1035,N_1092);
and U1157 (N_1157,N_1004,N_1036);
nor U1158 (N_1158,N_1060,N_1005);
or U1159 (N_1159,N_1037,N_1084);
nor U1160 (N_1160,N_1096,N_1038);
nor U1161 (N_1161,N_1005,N_1006);
or U1162 (N_1162,N_1057,N_1088);
or U1163 (N_1163,N_1088,N_1071);
and U1164 (N_1164,N_1007,N_1036);
or U1165 (N_1165,N_1032,N_1013);
or U1166 (N_1166,N_1087,N_1018);
nand U1167 (N_1167,N_1007,N_1086);
nor U1168 (N_1168,N_1002,N_1072);
nor U1169 (N_1169,N_1094,N_1075);
and U1170 (N_1170,N_1099,N_1080);
or U1171 (N_1171,N_1074,N_1031);
and U1172 (N_1172,N_1097,N_1065);
nand U1173 (N_1173,N_1044,N_1054);
nor U1174 (N_1174,N_1069,N_1043);
and U1175 (N_1175,N_1002,N_1054);
nor U1176 (N_1176,N_1033,N_1052);
xnor U1177 (N_1177,N_1091,N_1015);
nand U1178 (N_1178,N_1041,N_1006);
nand U1179 (N_1179,N_1039,N_1057);
and U1180 (N_1180,N_1009,N_1033);
xnor U1181 (N_1181,N_1078,N_1074);
and U1182 (N_1182,N_1088,N_1099);
xor U1183 (N_1183,N_1029,N_1031);
and U1184 (N_1184,N_1026,N_1039);
or U1185 (N_1185,N_1098,N_1032);
or U1186 (N_1186,N_1014,N_1062);
or U1187 (N_1187,N_1014,N_1069);
nor U1188 (N_1188,N_1088,N_1007);
nand U1189 (N_1189,N_1046,N_1090);
nor U1190 (N_1190,N_1050,N_1056);
nand U1191 (N_1191,N_1066,N_1058);
xnor U1192 (N_1192,N_1083,N_1075);
and U1193 (N_1193,N_1099,N_1036);
or U1194 (N_1194,N_1072,N_1019);
nor U1195 (N_1195,N_1058,N_1035);
xor U1196 (N_1196,N_1045,N_1040);
or U1197 (N_1197,N_1021,N_1058);
xnor U1198 (N_1198,N_1025,N_1051);
nand U1199 (N_1199,N_1083,N_1093);
and U1200 (N_1200,N_1161,N_1159);
nor U1201 (N_1201,N_1180,N_1116);
nand U1202 (N_1202,N_1164,N_1196);
or U1203 (N_1203,N_1167,N_1154);
nand U1204 (N_1204,N_1193,N_1128);
nand U1205 (N_1205,N_1145,N_1134);
xnor U1206 (N_1206,N_1187,N_1178);
xor U1207 (N_1207,N_1166,N_1138);
nor U1208 (N_1208,N_1107,N_1182);
and U1209 (N_1209,N_1109,N_1165);
nand U1210 (N_1210,N_1197,N_1174);
nand U1211 (N_1211,N_1133,N_1170);
xnor U1212 (N_1212,N_1160,N_1151);
xor U1213 (N_1213,N_1155,N_1100);
xnor U1214 (N_1214,N_1137,N_1142);
nand U1215 (N_1215,N_1139,N_1156);
nor U1216 (N_1216,N_1189,N_1188);
nor U1217 (N_1217,N_1104,N_1121);
xnor U1218 (N_1218,N_1130,N_1126);
nor U1219 (N_1219,N_1129,N_1198);
nor U1220 (N_1220,N_1191,N_1173);
and U1221 (N_1221,N_1163,N_1108);
xor U1222 (N_1222,N_1131,N_1162);
xor U1223 (N_1223,N_1105,N_1127);
xor U1224 (N_1224,N_1195,N_1184);
nand U1225 (N_1225,N_1111,N_1106);
nor U1226 (N_1226,N_1113,N_1147);
and U1227 (N_1227,N_1192,N_1144);
nand U1228 (N_1228,N_1115,N_1181);
nor U1229 (N_1229,N_1149,N_1148);
and U1230 (N_1230,N_1194,N_1136);
xnor U1231 (N_1231,N_1177,N_1146);
xor U1232 (N_1232,N_1176,N_1114);
nor U1233 (N_1233,N_1101,N_1119);
xnor U1234 (N_1234,N_1117,N_1112);
nand U1235 (N_1235,N_1102,N_1152);
and U1236 (N_1236,N_1150,N_1143);
nand U1237 (N_1237,N_1172,N_1169);
nor U1238 (N_1238,N_1123,N_1118);
nand U1239 (N_1239,N_1110,N_1103);
nor U1240 (N_1240,N_1175,N_1132);
nand U1241 (N_1241,N_1199,N_1157);
nor U1242 (N_1242,N_1171,N_1190);
or U1243 (N_1243,N_1185,N_1168);
and U1244 (N_1244,N_1120,N_1124);
or U1245 (N_1245,N_1125,N_1135);
nor U1246 (N_1246,N_1179,N_1183);
or U1247 (N_1247,N_1153,N_1141);
and U1248 (N_1248,N_1186,N_1158);
or U1249 (N_1249,N_1122,N_1140);
xnor U1250 (N_1250,N_1185,N_1151);
or U1251 (N_1251,N_1148,N_1167);
xor U1252 (N_1252,N_1122,N_1138);
nor U1253 (N_1253,N_1160,N_1136);
nor U1254 (N_1254,N_1102,N_1122);
nand U1255 (N_1255,N_1114,N_1182);
nand U1256 (N_1256,N_1119,N_1174);
nand U1257 (N_1257,N_1115,N_1196);
nor U1258 (N_1258,N_1108,N_1121);
or U1259 (N_1259,N_1115,N_1194);
xnor U1260 (N_1260,N_1183,N_1102);
nor U1261 (N_1261,N_1163,N_1109);
xor U1262 (N_1262,N_1184,N_1179);
nand U1263 (N_1263,N_1199,N_1178);
or U1264 (N_1264,N_1131,N_1135);
nand U1265 (N_1265,N_1194,N_1108);
nand U1266 (N_1266,N_1191,N_1110);
and U1267 (N_1267,N_1160,N_1179);
nor U1268 (N_1268,N_1171,N_1117);
xnor U1269 (N_1269,N_1197,N_1115);
xor U1270 (N_1270,N_1121,N_1116);
xor U1271 (N_1271,N_1181,N_1113);
nor U1272 (N_1272,N_1107,N_1106);
and U1273 (N_1273,N_1102,N_1184);
nand U1274 (N_1274,N_1187,N_1192);
nand U1275 (N_1275,N_1163,N_1190);
nand U1276 (N_1276,N_1119,N_1138);
nand U1277 (N_1277,N_1116,N_1140);
xnor U1278 (N_1278,N_1131,N_1122);
nor U1279 (N_1279,N_1180,N_1195);
nand U1280 (N_1280,N_1137,N_1165);
nand U1281 (N_1281,N_1120,N_1189);
xor U1282 (N_1282,N_1159,N_1181);
xor U1283 (N_1283,N_1106,N_1173);
xor U1284 (N_1284,N_1110,N_1101);
nand U1285 (N_1285,N_1180,N_1147);
xnor U1286 (N_1286,N_1195,N_1142);
xnor U1287 (N_1287,N_1158,N_1117);
nor U1288 (N_1288,N_1156,N_1157);
xnor U1289 (N_1289,N_1165,N_1183);
and U1290 (N_1290,N_1181,N_1175);
nor U1291 (N_1291,N_1162,N_1103);
nand U1292 (N_1292,N_1119,N_1113);
nand U1293 (N_1293,N_1191,N_1189);
or U1294 (N_1294,N_1133,N_1110);
xnor U1295 (N_1295,N_1167,N_1115);
nand U1296 (N_1296,N_1197,N_1159);
or U1297 (N_1297,N_1183,N_1103);
xor U1298 (N_1298,N_1133,N_1140);
and U1299 (N_1299,N_1129,N_1171);
xor U1300 (N_1300,N_1202,N_1232);
nor U1301 (N_1301,N_1229,N_1220);
or U1302 (N_1302,N_1216,N_1294);
or U1303 (N_1303,N_1224,N_1276);
xnor U1304 (N_1304,N_1272,N_1239);
nor U1305 (N_1305,N_1251,N_1255);
nand U1306 (N_1306,N_1291,N_1277);
nand U1307 (N_1307,N_1295,N_1211);
and U1308 (N_1308,N_1227,N_1269);
xor U1309 (N_1309,N_1209,N_1242);
and U1310 (N_1310,N_1244,N_1204);
nor U1311 (N_1311,N_1285,N_1250);
nand U1312 (N_1312,N_1258,N_1252);
and U1313 (N_1313,N_1282,N_1207);
or U1314 (N_1314,N_1208,N_1225);
xnor U1315 (N_1315,N_1230,N_1206);
and U1316 (N_1316,N_1212,N_1288);
or U1317 (N_1317,N_1274,N_1289);
and U1318 (N_1318,N_1284,N_1218);
nor U1319 (N_1319,N_1270,N_1201);
nand U1320 (N_1320,N_1249,N_1219);
nor U1321 (N_1321,N_1233,N_1205);
nor U1322 (N_1322,N_1240,N_1245);
nand U1323 (N_1323,N_1271,N_1223);
and U1324 (N_1324,N_1298,N_1247);
nor U1325 (N_1325,N_1283,N_1237);
nor U1326 (N_1326,N_1200,N_1238);
nor U1327 (N_1327,N_1254,N_1273);
nand U1328 (N_1328,N_1263,N_1241);
and U1329 (N_1329,N_1275,N_1226);
nor U1330 (N_1330,N_1278,N_1296);
or U1331 (N_1331,N_1246,N_1256);
or U1332 (N_1332,N_1217,N_1297);
nand U1333 (N_1333,N_1293,N_1261);
or U1334 (N_1334,N_1210,N_1268);
nand U1335 (N_1335,N_1290,N_1248);
or U1336 (N_1336,N_1222,N_1257);
xor U1337 (N_1337,N_1221,N_1292);
and U1338 (N_1338,N_1266,N_1236);
xor U1339 (N_1339,N_1281,N_1253);
xnor U1340 (N_1340,N_1286,N_1228);
nor U1341 (N_1341,N_1262,N_1279);
or U1342 (N_1342,N_1265,N_1267);
or U1343 (N_1343,N_1260,N_1214);
nand U1344 (N_1344,N_1280,N_1243);
nor U1345 (N_1345,N_1213,N_1231);
and U1346 (N_1346,N_1234,N_1299);
xor U1347 (N_1347,N_1235,N_1215);
nor U1348 (N_1348,N_1259,N_1264);
nand U1349 (N_1349,N_1287,N_1203);
xor U1350 (N_1350,N_1289,N_1227);
nor U1351 (N_1351,N_1214,N_1233);
nand U1352 (N_1352,N_1252,N_1212);
nor U1353 (N_1353,N_1237,N_1201);
and U1354 (N_1354,N_1288,N_1289);
nand U1355 (N_1355,N_1254,N_1274);
or U1356 (N_1356,N_1284,N_1220);
or U1357 (N_1357,N_1236,N_1222);
xor U1358 (N_1358,N_1222,N_1215);
xor U1359 (N_1359,N_1202,N_1239);
and U1360 (N_1360,N_1202,N_1294);
xor U1361 (N_1361,N_1274,N_1257);
or U1362 (N_1362,N_1230,N_1242);
and U1363 (N_1363,N_1213,N_1278);
nor U1364 (N_1364,N_1289,N_1251);
or U1365 (N_1365,N_1280,N_1251);
and U1366 (N_1366,N_1224,N_1286);
or U1367 (N_1367,N_1274,N_1250);
nand U1368 (N_1368,N_1252,N_1266);
or U1369 (N_1369,N_1216,N_1215);
or U1370 (N_1370,N_1272,N_1231);
xor U1371 (N_1371,N_1269,N_1218);
nand U1372 (N_1372,N_1276,N_1204);
or U1373 (N_1373,N_1209,N_1293);
xnor U1374 (N_1374,N_1220,N_1261);
xor U1375 (N_1375,N_1251,N_1224);
nand U1376 (N_1376,N_1205,N_1271);
or U1377 (N_1377,N_1243,N_1216);
or U1378 (N_1378,N_1227,N_1291);
nor U1379 (N_1379,N_1235,N_1238);
or U1380 (N_1380,N_1287,N_1297);
xnor U1381 (N_1381,N_1256,N_1274);
nand U1382 (N_1382,N_1228,N_1278);
xnor U1383 (N_1383,N_1221,N_1296);
and U1384 (N_1384,N_1297,N_1214);
nand U1385 (N_1385,N_1206,N_1284);
and U1386 (N_1386,N_1261,N_1246);
or U1387 (N_1387,N_1201,N_1233);
nand U1388 (N_1388,N_1235,N_1252);
nand U1389 (N_1389,N_1212,N_1257);
and U1390 (N_1390,N_1258,N_1256);
xor U1391 (N_1391,N_1295,N_1251);
nand U1392 (N_1392,N_1288,N_1295);
xnor U1393 (N_1393,N_1220,N_1234);
or U1394 (N_1394,N_1283,N_1203);
xor U1395 (N_1395,N_1238,N_1250);
xnor U1396 (N_1396,N_1202,N_1236);
nor U1397 (N_1397,N_1273,N_1265);
or U1398 (N_1398,N_1288,N_1293);
xnor U1399 (N_1399,N_1255,N_1260);
and U1400 (N_1400,N_1345,N_1349);
nand U1401 (N_1401,N_1361,N_1335);
nand U1402 (N_1402,N_1359,N_1311);
xnor U1403 (N_1403,N_1332,N_1352);
nor U1404 (N_1404,N_1360,N_1379);
and U1405 (N_1405,N_1363,N_1397);
and U1406 (N_1406,N_1340,N_1372);
nand U1407 (N_1407,N_1326,N_1386);
nor U1408 (N_1408,N_1317,N_1394);
xnor U1409 (N_1409,N_1371,N_1342);
xor U1410 (N_1410,N_1374,N_1313);
and U1411 (N_1411,N_1316,N_1355);
and U1412 (N_1412,N_1344,N_1350);
nand U1413 (N_1413,N_1329,N_1353);
nor U1414 (N_1414,N_1376,N_1306);
nand U1415 (N_1415,N_1341,N_1347);
and U1416 (N_1416,N_1330,N_1339);
nor U1417 (N_1417,N_1358,N_1310);
and U1418 (N_1418,N_1377,N_1322);
nor U1419 (N_1419,N_1343,N_1334);
or U1420 (N_1420,N_1388,N_1328);
nor U1421 (N_1421,N_1314,N_1324);
nor U1422 (N_1422,N_1336,N_1318);
xnor U1423 (N_1423,N_1348,N_1373);
xnor U1424 (N_1424,N_1384,N_1395);
nand U1425 (N_1425,N_1365,N_1375);
or U1426 (N_1426,N_1382,N_1368);
xor U1427 (N_1427,N_1387,N_1305);
nand U1428 (N_1428,N_1303,N_1319);
and U1429 (N_1429,N_1308,N_1370);
xor U1430 (N_1430,N_1301,N_1315);
xnor U1431 (N_1431,N_1389,N_1369);
xnor U1432 (N_1432,N_1385,N_1337);
or U1433 (N_1433,N_1323,N_1367);
xnor U1434 (N_1434,N_1300,N_1390);
xor U1435 (N_1435,N_1351,N_1383);
nor U1436 (N_1436,N_1307,N_1338);
xnor U1437 (N_1437,N_1396,N_1302);
and U1438 (N_1438,N_1380,N_1392);
xnor U1439 (N_1439,N_1331,N_1393);
and U1440 (N_1440,N_1391,N_1378);
and U1441 (N_1441,N_1398,N_1362);
or U1442 (N_1442,N_1304,N_1333);
and U1443 (N_1443,N_1366,N_1321);
nand U1444 (N_1444,N_1312,N_1354);
nand U1445 (N_1445,N_1320,N_1309);
xor U1446 (N_1446,N_1346,N_1327);
nand U1447 (N_1447,N_1325,N_1357);
nand U1448 (N_1448,N_1356,N_1364);
nor U1449 (N_1449,N_1399,N_1381);
xnor U1450 (N_1450,N_1396,N_1306);
nand U1451 (N_1451,N_1304,N_1369);
xnor U1452 (N_1452,N_1354,N_1378);
and U1453 (N_1453,N_1361,N_1357);
and U1454 (N_1454,N_1364,N_1300);
and U1455 (N_1455,N_1395,N_1331);
nand U1456 (N_1456,N_1346,N_1324);
xnor U1457 (N_1457,N_1387,N_1336);
xor U1458 (N_1458,N_1320,N_1381);
and U1459 (N_1459,N_1312,N_1329);
nor U1460 (N_1460,N_1352,N_1376);
xnor U1461 (N_1461,N_1337,N_1378);
or U1462 (N_1462,N_1379,N_1326);
nor U1463 (N_1463,N_1338,N_1339);
nand U1464 (N_1464,N_1332,N_1365);
xnor U1465 (N_1465,N_1358,N_1362);
and U1466 (N_1466,N_1398,N_1349);
and U1467 (N_1467,N_1309,N_1385);
and U1468 (N_1468,N_1315,N_1344);
nand U1469 (N_1469,N_1376,N_1383);
nand U1470 (N_1470,N_1352,N_1373);
and U1471 (N_1471,N_1347,N_1326);
and U1472 (N_1472,N_1398,N_1371);
nand U1473 (N_1473,N_1347,N_1327);
and U1474 (N_1474,N_1339,N_1325);
nand U1475 (N_1475,N_1312,N_1383);
xor U1476 (N_1476,N_1325,N_1311);
or U1477 (N_1477,N_1323,N_1311);
and U1478 (N_1478,N_1346,N_1319);
nor U1479 (N_1479,N_1364,N_1313);
and U1480 (N_1480,N_1343,N_1353);
or U1481 (N_1481,N_1324,N_1344);
or U1482 (N_1482,N_1332,N_1339);
and U1483 (N_1483,N_1318,N_1382);
nor U1484 (N_1484,N_1358,N_1394);
and U1485 (N_1485,N_1374,N_1341);
xnor U1486 (N_1486,N_1391,N_1392);
nor U1487 (N_1487,N_1329,N_1315);
nand U1488 (N_1488,N_1364,N_1344);
and U1489 (N_1489,N_1332,N_1363);
nand U1490 (N_1490,N_1335,N_1350);
or U1491 (N_1491,N_1380,N_1369);
xnor U1492 (N_1492,N_1381,N_1303);
xor U1493 (N_1493,N_1303,N_1350);
nor U1494 (N_1494,N_1349,N_1330);
xor U1495 (N_1495,N_1344,N_1333);
and U1496 (N_1496,N_1371,N_1384);
xor U1497 (N_1497,N_1302,N_1352);
nor U1498 (N_1498,N_1329,N_1335);
xnor U1499 (N_1499,N_1346,N_1397);
nand U1500 (N_1500,N_1461,N_1470);
or U1501 (N_1501,N_1434,N_1422);
or U1502 (N_1502,N_1442,N_1469);
nor U1503 (N_1503,N_1454,N_1490);
nand U1504 (N_1504,N_1426,N_1456);
nor U1505 (N_1505,N_1416,N_1493);
nand U1506 (N_1506,N_1427,N_1455);
nand U1507 (N_1507,N_1462,N_1492);
and U1508 (N_1508,N_1480,N_1430);
and U1509 (N_1509,N_1438,N_1499);
xor U1510 (N_1510,N_1436,N_1495);
nor U1511 (N_1511,N_1453,N_1423);
nor U1512 (N_1512,N_1404,N_1451);
nand U1513 (N_1513,N_1484,N_1467);
xor U1514 (N_1514,N_1415,N_1431);
xor U1515 (N_1515,N_1466,N_1450);
nor U1516 (N_1516,N_1474,N_1457);
xor U1517 (N_1517,N_1472,N_1494);
and U1518 (N_1518,N_1409,N_1446);
xnor U1519 (N_1519,N_1440,N_1489);
nand U1520 (N_1520,N_1443,N_1401);
xnor U1521 (N_1521,N_1497,N_1411);
and U1522 (N_1522,N_1447,N_1441);
nand U1523 (N_1523,N_1475,N_1465);
and U1524 (N_1524,N_1452,N_1464);
xor U1525 (N_1525,N_1437,N_1471);
xnor U1526 (N_1526,N_1458,N_1413);
nor U1527 (N_1527,N_1425,N_1410);
and U1528 (N_1528,N_1476,N_1478);
xor U1529 (N_1529,N_1496,N_1463);
nand U1530 (N_1530,N_1412,N_1479);
or U1531 (N_1531,N_1485,N_1473);
and U1532 (N_1532,N_1486,N_1417);
nor U1533 (N_1533,N_1477,N_1406);
nand U1534 (N_1534,N_1419,N_1444);
and U1535 (N_1535,N_1403,N_1498);
and U1536 (N_1536,N_1435,N_1428);
or U1537 (N_1537,N_1400,N_1482);
nor U1538 (N_1538,N_1491,N_1433);
and U1539 (N_1539,N_1468,N_1488);
xor U1540 (N_1540,N_1429,N_1481);
nand U1541 (N_1541,N_1424,N_1487);
or U1542 (N_1542,N_1449,N_1408);
xnor U1543 (N_1543,N_1460,N_1448);
nor U1544 (N_1544,N_1439,N_1402);
xor U1545 (N_1545,N_1432,N_1483);
nor U1546 (N_1546,N_1445,N_1459);
nor U1547 (N_1547,N_1407,N_1421);
xnor U1548 (N_1548,N_1420,N_1414);
and U1549 (N_1549,N_1418,N_1405);
or U1550 (N_1550,N_1493,N_1492);
or U1551 (N_1551,N_1447,N_1435);
nor U1552 (N_1552,N_1484,N_1450);
or U1553 (N_1553,N_1467,N_1470);
xor U1554 (N_1554,N_1439,N_1463);
xor U1555 (N_1555,N_1462,N_1451);
or U1556 (N_1556,N_1419,N_1463);
and U1557 (N_1557,N_1453,N_1400);
xor U1558 (N_1558,N_1431,N_1405);
xor U1559 (N_1559,N_1407,N_1416);
xor U1560 (N_1560,N_1454,N_1402);
nand U1561 (N_1561,N_1460,N_1440);
and U1562 (N_1562,N_1466,N_1464);
nand U1563 (N_1563,N_1485,N_1483);
nor U1564 (N_1564,N_1446,N_1443);
xor U1565 (N_1565,N_1466,N_1414);
or U1566 (N_1566,N_1466,N_1458);
xor U1567 (N_1567,N_1461,N_1478);
xor U1568 (N_1568,N_1403,N_1468);
nor U1569 (N_1569,N_1498,N_1494);
and U1570 (N_1570,N_1455,N_1475);
nand U1571 (N_1571,N_1435,N_1441);
or U1572 (N_1572,N_1494,N_1448);
nor U1573 (N_1573,N_1448,N_1421);
nor U1574 (N_1574,N_1415,N_1424);
nor U1575 (N_1575,N_1442,N_1452);
xnor U1576 (N_1576,N_1464,N_1430);
and U1577 (N_1577,N_1469,N_1495);
and U1578 (N_1578,N_1444,N_1457);
and U1579 (N_1579,N_1430,N_1492);
and U1580 (N_1580,N_1456,N_1493);
and U1581 (N_1581,N_1470,N_1435);
or U1582 (N_1582,N_1438,N_1488);
and U1583 (N_1583,N_1437,N_1457);
nor U1584 (N_1584,N_1456,N_1437);
or U1585 (N_1585,N_1441,N_1434);
nand U1586 (N_1586,N_1484,N_1427);
or U1587 (N_1587,N_1443,N_1452);
and U1588 (N_1588,N_1413,N_1474);
nand U1589 (N_1589,N_1497,N_1432);
nand U1590 (N_1590,N_1494,N_1470);
and U1591 (N_1591,N_1496,N_1477);
or U1592 (N_1592,N_1444,N_1456);
nand U1593 (N_1593,N_1479,N_1413);
or U1594 (N_1594,N_1452,N_1406);
nor U1595 (N_1595,N_1492,N_1456);
and U1596 (N_1596,N_1416,N_1400);
nor U1597 (N_1597,N_1407,N_1446);
xnor U1598 (N_1598,N_1427,N_1458);
and U1599 (N_1599,N_1401,N_1430);
xor U1600 (N_1600,N_1502,N_1580);
nor U1601 (N_1601,N_1564,N_1528);
nand U1602 (N_1602,N_1592,N_1534);
xnor U1603 (N_1603,N_1518,N_1544);
xor U1604 (N_1604,N_1586,N_1530);
nor U1605 (N_1605,N_1574,N_1531);
and U1606 (N_1606,N_1510,N_1538);
or U1607 (N_1607,N_1526,N_1519);
nor U1608 (N_1608,N_1514,N_1557);
xor U1609 (N_1609,N_1571,N_1539);
and U1610 (N_1610,N_1578,N_1550);
and U1611 (N_1611,N_1535,N_1547);
nor U1612 (N_1612,N_1554,N_1591);
or U1613 (N_1613,N_1559,N_1575);
or U1614 (N_1614,N_1569,N_1537);
nand U1615 (N_1615,N_1542,N_1572);
xor U1616 (N_1616,N_1561,N_1565);
xnor U1617 (N_1617,N_1509,N_1541);
nand U1618 (N_1618,N_1582,N_1545);
and U1619 (N_1619,N_1562,N_1525);
xor U1620 (N_1620,N_1506,N_1556);
xor U1621 (N_1621,N_1508,N_1517);
or U1622 (N_1622,N_1524,N_1560);
or U1623 (N_1623,N_1563,N_1555);
nand U1624 (N_1624,N_1595,N_1553);
and U1625 (N_1625,N_1579,N_1511);
and U1626 (N_1626,N_1599,N_1540);
and U1627 (N_1627,N_1570,N_1503);
and U1628 (N_1628,N_1529,N_1513);
xnor U1629 (N_1629,N_1521,N_1551);
and U1630 (N_1630,N_1549,N_1512);
nor U1631 (N_1631,N_1507,N_1533);
xnor U1632 (N_1632,N_1577,N_1596);
nor U1633 (N_1633,N_1594,N_1500);
and U1634 (N_1634,N_1588,N_1505);
and U1635 (N_1635,N_1590,N_1584);
and U1636 (N_1636,N_1598,N_1548);
nand U1637 (N_1637,N_1527,N_1593);
nand U1638 (N_1638,N_1585,N_1552);
and U1639 (N_1639,N_1573,N_1566);
and U1640 (N_1640,N_1581,N_1589);
and U1641 (N_1641,N_1597,N_1558);
or U1642 (N_1642,N_1536,N_1587);
and U1643 (N_1643,N_1523,N_1532);
nand U1644 (N_1644,N_1543,N_1567);
nand U1645 (N_1645,N_1576,N_1568);
nor U1646 (N_1646,N_1504,N_1583);
and U1647 (N_1647,N_1522,N_1516);
nor U1648 (N_1648,N_1515,N_1520);
and U1649 (N_1649,N_1546,N_1501);
or U1650 (N_1650,N_1514,N_1594);
nand U1651 (N_1651,N_1532,N_1585);
or U1652 (N_1652,N_1588,N_1569);
and U1653 (N_1653,N_1564,N_1546);
and U1654 (N_1654,N_1578,N_1594);
xor U1655 (N_1655,N_1519,N_1535);
nand U1656 (N_1656,N_1507,N_1571);
or U1657 (N_1657,N_1591,N_1573);
and U1658 (N_1658,N_1536,N_1589);
and U1659 (N_1659,N_1537,N_1524);
nor U1660 (N_1660,N_1549,N_1544);
or U1661 (N_1661,N_1564,N_1580);
or U1662 (N_1662,N_1590,N_1503);
xnor U1663 (N_1663,N_1580,N_1565);
nand U1664 (N_1664,N_1566,N_1516);
and U1665 (N_1665,N_1556,N_1572);
xnor U1666 (N_1666,N_1500,N_1537);
xnor U1667 (N_1667,N_1585,N_1586);
nor U1668 (N_1668,N_1540,N_1523);
nand U1669 (N_1669,N_1536,N_1580);
xnor U1670 (N_1670,N_1547,N_1578);
nor U1671 (N_1671,N_1547,N_1524);
nand U1672 (N_1672,N_1558,N_1556);
xnor U1673 (N_1673,N_1513,N_1506);
or U1674 (N_1674,N_1534,N_1548);
or U1675 (N_1675,N_1532,N_1533);
nor U1676 (N_1676,N_1575,N_1512);
or U1677 (N_1677,N_1522,N_1541);
or U1678 (N_1678,N_1584,N_1525);
nand U1679 (N_1679,N_1531,N_1552);
or U1680 (N_1680,N_1529,N_1587);
xor U1681 (N_1681,N_1567,N_1556);
or U1682 (N_1682,N_1586,N_1535);
nand U1683 (N_1683,N_1527,N_1507);
xnor U1684 (N_1684,N_1500,N_1562);
and U1685 (N_1685,N_1592,N_1571);
nand U1686 (N_1686,N_1529,N_1595);
nand U1687 (N_1687,N_1501,N_1533);
nor U1688 (N_1688,N_1573,N_1593);
or U1689 (N_1689,N_1518,N_1563);
and U1690 (N_1690,N_1543,N_1516);
or U1691 (N_1691,N_1571,N_1538);
xor U1692 (N_1692,N_1594,N_1575);
xnor U1693 (N_1693,N_1540,N_1552);
nor U1694 (N_1694,N_1544,N_1571);
and U1695 (N_1695,N_1582,N_1566);
or U1696 (N_1696,N_1522,N_1521);
nand U1697 (N_1697,N_1569,N_1517);
nor U1698 (N_1698,N_1568,N_1503);
or U1699 (N_1699,N_1550,N_1584);
xor U1700 (N_1700,N_1618,N_1690);
nor U1701 (N_1701,N_1678,N_1687);
nor U1702 (N_1702,N_1634,N_1676);
or U1703 (N_1703,N_1670,N_1612);
and U1704 (N_1704,N_1631,N_1623);
xor U1705 (N_1705,N_1692,N_1607);
nand U1706 (N_1706,N_1668,N_1602);
nor U1707 (N_1707,N_1673,N_1650);
nor U1708 (N_1708,N_1667,N_1620);
nor U1709 (N_1709,N_1686,N_1640);
xnor U1710 (N_1710,N_1675,N_1601);
nor U1711 (N_1711,N_1688,N_1666);
nand U1712 (N_1712,N_1665,N_1639);
nand U1713 (N_1713,N_1630,N_1699);
or U1714 (N_1714,N_1658,N_1677);
nand U1715 (N_1715,N_1651,N_1672);
nor U1716 (N_1716,N_1619,N_1679);
nor U1717 (N_1717,N_1641,N_1671);
nor U1718 (N_1718,N_1695,N_1661);
nand U1719 (N_1719,N_1697,N_1604);
nand U1720 (N_1720,N_1683,N_1660);
xor U1721 (N_1721,N_1608,N_1696);
and U1722 (N_1722,N_1689,N_1637);
or U1723 (N_1723,N_1609,N_1647);
nor U1724 (N_1724,N_1664,N_1603);
nand U1725 (N_1725,N_1614,N_1627);
and U1726 (N_1726,N_1662,N_1633);
nand U1727 (N_1727,N_1621,N_1652);
or U1728 (N_1728,N_1653,N_1636);
xor U1729 (N_1729,N_1628,N_1610);
xnor U1730 (N_1730,N_1682,N_1654);
or U1731 (N_1731,N_1625,N_1656);
and U1732 (N_1732,N_1645,N_1698);
or U1733 (N_1733,N_1606,N_1624);
nor U1734 (N_1734,N_1642,N_1600);
and U1735 (N_1735,N_1644,N_1629);
and U1736 (N_1736,N_1657,N_1674);
nand U1737 (N_1737,N_1691,N_1643);
nand U1738 (N_1738,N_1685,N_1635);
nand U1739 (N_1739,N_1655,N_1669);
nor U1740 (N_1740,N_1622,N_1638);
nand U1741 (N_1741,N_1693,N_1681);
and U1742 (N_1742,N_1684,N_1648);
nor U1743 (N_1743,N_1663,N_1611);
nor U1744 (N_1744,N_1694,N_1646);
nor U1745 (N_1745,N_1613,N_1615);
or U1746 (N_1746,N_1632,N_1626);
or U1747 (N_1747,N_1617,N_1649);
nor U1748 (N_1748,N_1659,N_1616);
nor U1749 (N_1749,N_1680,N_1605);
nand U1750 (N_1750,N_1676,N_1645);
or U1751 (N_1751,N_1667,N_1636);
and U1752 (N_1752,N_1656,N_1605);
or U1753 (N_1753,N_1628,N_1688);
nor U1754 (N_1754,N_1666,N_1609);
nand U1755 (N_1755,N_1694,N_1658);
xnor U1756 (N_1756,N_1610,N_1670);
xnor U1757 (N_1757,N_1691,N_1626);
and U1758 (N_1758,N_1675,N_1642);
xnor U1759 (N_1759,N_1695,N_1613);
xnor U1760 (N_1760,N_1612,N_1694);
xnor U1761 (N_1761,N_1607,N_1620);
xnor U1762 (N_1762,N_1648,N_1642);
nand U1763 (N_1763,N_1622,N_1647);
nand U1764 (N_1764,N_1674,N_1668);
or U1765 (N_1765,N_1617,N_1656);
nor U1766 (N_1766,N_1620,N_1668);
or U1767 (N_1767,N_1637,N_1666);
and U1768 (N_1768,N_1687,N_1609);
nand U1769 (N_1769,N_1640,N_1684);
xnor U1770 (N_1770,N_1672,N_1679);
or U1771 (N_1771,N_1636,N_1643);
and U1772 (N_1772,N_1606,N_1663);
nand U1773 (N_1773,N_1672,N_1682);
or U1774 (N_1774,N_1620,N_1621);
nand U1775 (N_1775,N_1674,N_1669);
or U1776 (N_1776,N_1626,N_1628);
or U1777 (N_1777,N_1692,N_1638);
nor U1778 (N_1778,N_1605,N_1684);
xor U1779 (N_1779,N_1658,N_1657);
nor U1780 (N_1780,N_1687,N_1642);
and U1781 (N_1781,N_1630,N_1697);
or U1782 (N_1782,N_1696,N_1631);
nor U1783 (N_1783,N_1636,N_1621);
nand U1784 (N_1784,N_1698,N_1655);
nand U1785 (N_1785,N_1660,N_1666);
nor U1786 (N_1786,N_1606,N_1657);
xor U1787 (N_1787,N_1613,N_1686);
nand U1788 (N_1788,N_1634,N_1636);
and U1789 (N_1789,N_1692,N_1654);
nand U1790 (N_1790,N_1632,N_1624);
nand U1791 (N_1791,N_1644,N_1615);
and U1792 (N_1792,N_1632,N_1628);
nor U1793 (N_1793,N_1600,N_1654);
and U1794 (N_1794,N_1677,N_1669);
xnor U1795 (N_1795,N_1663,N_1680);
and U1796 (N_1796,N_1602,N_1665);
xnor U1797 (N_1797,N_1652,N_1620);
nor U1798 (N_1798,N_1629,N_1601);
or U1799 (N_1799,N_1656,N_1612);
xnor U1800 (N_1800,N_1777,N_1736);
nor U1801 (N_1801,N_1796,N_1757);
nor U1802 (N_1802,N_1778,N_1782);
nand U1803 (N_1803,N_1791,N_1719);
or U1804 (N_1804,N_1784,N_1787);
nand U1805 (N_1805,N_1767,N_1763);
xor U1806 (N_1806,N_1722,N_1738);
nor U1807 (N_1807,N_1771,N_1724);
and U1808 (N_1808,N_1776,N_1740);
and U1809 (N_1809,N_1758,N_1788);
nand U1810 (N_1810,N_1704,N_1733);
nand U1811 (N_1811,N_1750,N_1799);
and U1812 (N_1812,N_1793,N_1751);
or U1813 (N_1813,N_1747,N_1701);
or U1814 (N_1814,N_1730,N_1785);
or U1815 (N_1815,N_1781,N_1735);
nand U1816 (N_1816,N_1727,N_1737);
nor U1817 (N_1817,N_1762,N_1749);
and U1818 (N_1818,N_1710,N_1798);
and U1819 (N_1819,N_1706,N_1744);
or U1820 (N_1820,N_1734,N_1726);
and U1821 (N_1821,N_1790,N_1728);
nand U1822 (N_1822,N_1780,N_1765);
xor U1823 (N_1823,N_1729,N_1752);
nor U1824 (N_1824,N_1774,N_1794);
or U1825 (N_1825,N_1797,N_1715);
nand U1826 (N_1826,N_1741,N_1714);
or U1827 (N_1827,N_1756,N_1773);
nor U1828 (N_1828,N_1713,N_1712);
or U1829 (N_1829,N_1742,N_1775);
nand U1830 (N_1830,N_1789,N_1703);
or U1831 (N_1831,N_1766,N_1720);
or U1832 (N_1832,N_1721,N_1770);
or U1833 (N_1833,N_1755,N_1753);
or U1834 (N_1834,N_1718,N_1760);
xor U1835 (N_1835,N_1709,N_1702);
and U1836 (N_1836,N_1754,N_1743);
xnor U1837 (N_1837,N_1700,N_1764);
xnor U1838 (N_1838,N_1716,N_1792);
and U1839 (N_1839,N_1768,N_1731);
or U1840 (N_1840,N_1705,N_1748);
or U1841 (N_1841,N_1779,N_1786);
or U1842 (N_1842,N_1717,N_1739);
and U1843 (N_1843,N_1725,N_1769);
xnor U1844 (N_1844,N_1783,N_1761);
xor U1845 (N_1845,N_1795,N_1759);
or U1846 (N_1846,N_1711,N_1772);
or U1847 (N_1847,N_1745,N_1707);
or U1848 (N_1848,N_1732,N_1746);
or U1849 (N_1849,N_1708,N_1723);
or U1850 (N_1850,N_1716,N_1754);
and U1851 (N_1851,N_1775,N_1740);
nor U1852 (N_1852,N_1724,N_1789);
xnor U1853 (N_1853,N_1775,N_1724);
or U1854 (N_1854,N_1780,N_1703);
xnor U1855 (N_1855,N_1778,N_1744);
and U1856 (N_1856,N_1783,N_1759);
or U1857 (N_1857,N_1733,N_1701);
nand U1858 (N_1858,N_1755,N_1703);
or U1859 (N_1859,N_1792,N_1790);
nor U1860 (N_1860,N_1739,N_1715);
and U1861 (N_1861,N_1752,N_1731);
or U1862 (N_1862,N_1733,N_1754);
and U1863 (N_1863,N_1704,N_1795);
and U1864 (N_1864,N_1712,N_1782);
or U1865 (N_1865,N_1719,N_1787);
nand U1866 (N_1866,N_1798,N_1752);
and U1867 (N_1867,N_1758,N_1745);
and U1868 (N_1868,N_1723,N_1758);
xnor U1869 (N_1869,N_1720,N_1754);
or U1870 (N_1870,N_1756,N_1722);
and U1871 (N_1871,N_1783,N_1764);
and U1872 (N_1872,N_1755,N_1795);
or U1873 (N_1873,N_1739,N_1772);
xnor U1874 (N_1874,N_1735,N_1764);
or U1875 (N_1875,N_1741,N_1790);
or U1876 (N_1876,N_1741,N_1756);
or U1877 (N_1877,N_1748,N_1710);
nor U1878 (N_1878,N_1780,N_1737);
nor U1879 (N_1879,N_1744,N_1798);
and U1880 (N_1880,N_1789,N_1706);
and U1881 (N_1881,N_1774,N_1732);
and U1882 (N_1882,N_1779,N_1771);
or U1883 (N_1883,N_1720,N_1757);
and U1884 (N_1884,N_1729,N_1741);
xor U1885 (N_1885,N_1738,N_1724);
xnor U1886 (N_1886,N_1759,N_1771);
nor U1887 (N_1887,N_1718,N_1757);
nand U1888 (N_1888,N_1715,N_1789);
xnor U1889 (N_1889,N_1749,N_1787);
nand U1890 (N_1890,N_1776,N_1738);
or U1891 (N_1891,N_1740,N_1785);
and U1892 (N_1892,N_1702,N_1712);
and U1893 (N_1893,N_1750,N_1709);
nand U1894 (N_1894,N_1767,N_1771);
and U1895 (N_1895,N_1719,N_1765);
nand U1896 (N_1896,N_1722,N_1747);
nand U1897 (N_1897,N_1712,N_1768);
xor U1898 (N_1898,N_1733,N_1721);
or U1899 (N_1899,N_1704,N_1742);
nor U1900 (N_1900,N_1859,N_1895);
xor U1901 (N_1901,N_1826,N_1862);
xor U1902 (N_1902,N_1844,N_1817);
xnor U1903 (N_1903,N_1877,N_1875);
nor U1904 (N_1904,N_1812,N_1821);
nand U1905 (N_1905,N_1848,N_1855);
nor U1906 (N_1906,N_1898,N_1813);
nor U1907 (N_1907,N_1883,N_1889);
nor U1908 (N_1908,N_1894,N_1831);
and U1909 (N_1909,N_1884,N_1888);
and U1910 (N_1910,N_1864,N_1845);
and U1911 (N_1911,N_1835,N_1870);
xor U1912 (N_1912,N_1827,N_1882);
or U1913 (N_1913,N_1881,N_1869);
nor U1914 (N_1914,N_1833,N_1816);
and U1915 (N_1915,N_1861,N_1856);
or U1916 (N_1916,N_1846,N_1868);
nand U1917 (N_1917,N_1892,N_1838);
xnor U1918 (N_1918,N_1890,N_1893);
or U1919 (N_1919,N_1829,N_1841);
nor U1920 (N_1920,N_1886,N_1876);
nor U1921 (N_1921,N_1822,N_1824);
xor U1922 (N_1922,N_1880,N_1878);
or U1923 (N_1923,N_1887,N_1857);
or U1924 (N_1924,N_1820,N_1805);
nor U1925 (N_1925,N_1872,N_1891);
nor U1926 (N_1926,N_1804,N_1832);
nand U1927 (N_1927,N_1871,N_1834);
nand U1928 (N_1928,N_1825,N_1819);
xor U1929 (N_1929,N_1849,N_1806);
xnor U1930 (N_1930,N_1863,N_1896);
xor U1931 (N_1931,N_1818,N_1807);
xnor U1932 (N_1932,N_1874,N_1866);
nand U1933 (N_1933,N_1837,N_1853);
nand U1934 (N_1934,N_1865,N_1801);
nand U1935 (N_1935,N_1808,N_1854);
xor U1936 (N_1936,N_1899,N_1852);
or U1937 (N_1937,N_1850,N_1860);
or U1938 (N_1938,N_1867,N_1802);
xnor U1939 (N_1939,N_1836,N_1815);
nand U1940 (N_1940,N_1858,N_1873);
xnor U1941 (N_1941,N_1810,N_1879);
xor U1942 (N_1942,N_1830,N_1843);
and U1943 (N_1943,N_1803,N_1809);
nor U1944 (N_1944,N_1811,N_1839);
nor U1945 (N_1945,N_1828,N_1814);
nand U1946 (N_1946,N_1842,N_1851);
or U1947 (N_1947,N_1840,N_1897);
and U1948 (N_1948,N_1885,N_1847);
or U1949 (N_1949,N_1823,N_1800);
xnor U1950 (N_1950,N_1809,N_1808);
xor U1951 (N_1951,N_1818,N_1880);
nor U1952 (N_1952,N_1861,N_1895);
xor U1953 (N_1953,N_1883,N_1836);
or U1954 (N_1954,N_1845,N_1802);
nor U1955 (N_1955,N_1874,N_1855);
xor U1956 (N_1956,N_1890,N_1846);
and U1957 (N_1957,N_1814,N_1800);
nand U1958 (N_1958,N_1876,N_1842);
nor U1959 (N_1959,N_1810,N_1837);
nor U1960 (N_1960,N_1884,N_1806);
and U1961 (N_1961,N_1856,N_1875);
xor U1962 (N_1962,N_1878,N_1860);
xor U1963 (N_1963,N_1802,N_1817);
nor U1964 (N_1964,N_1884,N_1837);
or U1965 (N_1965,N_1824,N_1803);
nor U1966 (N_1966,N_1840,N_1835);
or U1967 (N_1967,N_1816,N_1887);
nor U1968 (N_1968,N_1884,N_1851);
and U1969 (N_1969,N_1830,N_1807);
nand U1970 (N_1970,N_1870,N_1884);
nand U1971 (N_1971,N_1801,N_1877);
and U1972 (N_1972,N_1850,N_1863);
nor U1973 (N_1973,N_1865,N_1887);
xor U1974 (N_1974,N_1822,N_1841);
nor U1975 (N_1975,N_1849,N_1813);
xor U1976 (N_1976,N_1829,N_1814);
and U1977 (N_1977,N_1896,N_1829);
xnor U1978 (N_1978,N_1882,N_1801);
xor U1979 (N_1979,N_1874,N_1895);
nor U1980 (N_1980,N_1855,N_1868);
or U1981 (N_1981,N_1863,N_1815);
or U1982 (N_1982,N_1804,N_1834);
nor U1983 (N_1983,N_1826,N_1805);
nand U1984 (N_1984,N_1860,N_1893);
nand U1985 (N_1985,N_1877,N_1881);
xor U1986 (N_1986,N_1838,N_1860);
nor U1987 (N_1987,N_1808,N_1881);
or U1988 (N_1988,N_1801,N_1822);
or U1989 (N_1989,N_1876,N_1877);
and U1990 (N_1990,N_1814,N_1827);
or U1991 (N_1991,N_1839,N_1865);
nor U1992 (N_1992,N_1801,N_1888);
nor U1993 (N_1993,N_1870,N_1856);
xor U1994 (N_1994,N_1861,N_1887);
and U1995 (N_1995,N_1883,N_1811);
and U1996 (N_1996,N_1886,N_1864);
or U1997 (N_1997,N_1821,N_1808);
xnor U1998 (N_1998,N_1843,N_1874);
or U1999 (N_1999,N_1817,N_1804);
and U2000 (N_2000,N_1966,N_1928);
nand U2001 (N_2001,N_1967,N_1993);
or U2002 (N_2002,N_1912,N_1918);
and U2003 (N_2003,N_1929,N_1963);
nand U2004 (N_2004,N_1933,N_1985);
nand U2005 (N_2005,N_1907,N_1909);
nand U2006 (N_2006,N_1986,N_1936);
and U2007 (N_2007,N_1943,N_1983);
or U2008 (N_2008,N_1922,N_1908);
nand U2009 (N_2009,N_1952,N_1919);
nand U2010 (N_2010,N_1931,N_1914);
or U2011 (N_2011,N_1942,N_1934);
or U2012 (N_2012,N_1956,N_1930);
and U2013 (N_2013,N_1945,N_1997);
nor U2014 (N_2014,N_1944,N_1958);
nor U2015 (N_2015,N_1935,N_1987);
or U2016 (N_2016,N_1906,N_1996);
xnor U2017 (N_2017,N_1948,N_1968);
nand U2018 (N_2018,N_1980,N_1969);
nor U2019 (N_2019,N_1917,N_1981);
nor U2020 (N_2020,N_1960,N_1911);
nand U2021 (N_2021,N_1939,N_1998);
and U2022 (N_2022,N_1999,N_1905);
nand U2023 (N_2023,N_1989,N_1940);
or U2024 (N_2024,N_1916,N_1923);
nor U2025 (N_2025,N_1988,N_1913);
and U2026 (N_2026,N_1946,N_1965);
nor U2027 (N_2027,N_1957,N_1927);
xnor U2028 (N_2028,N_1950,N_1924);
xnor U2029 (N_2029,N_1925,N_1949);
and U2030 (N_2030,N_1941,N_1955);
nor U2031 (N_2031,N_1990,N_1953);
and U2032 (N_2032,N_1959,N_1974);
nor U2033 (N_2033,N_1995,N_1951);
or U2034 (N_2034,N_1982,N_1991);
or U2035 (N_2035,N_1938,N_1978);
and U2036 (N_2036,N_1984,N_1962);
nand U2037 (N_2037,N_1902,N_1977);
or U2038 (N_2038,N_1979,N_1915);
nand U2039 (N_2039,N_1901,N_1926);
nor U2040 (N_2040,N_1900,N_1975);
nand U2041 (N_2041,N_1937,N_1932);
or U2042 (N_2042,N_1964,N_1992);
nor U2043 (N_2043,N_1971,N_1970);
nand U2044 (N_2044,N_1973,N_1976);
or U2045 (N_2045,N_1961,N_1954);
or U2046 (N_2046,N_1994,N_1903);
and U2047 (N_2047,N_1904,N_1921);
or U2048 (N_2048,N_1910,N_1920);
or U2049 (N_2049,N_1947,N_1972);
nand U2050 (N_2050,N_1903,N_1970);
nor U2051 (N_2051,N_1998,N_1960);
nor U2052 (N_2052,N_1908,N_1923);
and U2053 (N_2053,N_1922,N_1992);
xor U2054 (N_2054,N_1961,N_1960);
and U2055 (N_2055,N_1910,N_1900);
or U2056 (N_2056,N_1912,N_1969);
nand U2057 (N_2057,N_1904,N_1924);
nor U2058 (N_2058,N_1933,N_1964);
or U2059 (N_2059,N_1945,N_1967);
xnor U2060 (N_2060,N_1929,N_1983);
xnor U2061 (N_2061,N_1939,N_1969);
nand U2062 (N_2062,N_1978,N_1906);
nand U2063 (N_2063,N_1948,N_1964);
xnor U2064 (N_2064,N_1900,N_1996);
xnor U2065 (N_2065,N_1942,N_1973);
and U2066 (N_2066,N_1946,N_1908);
nand U2067 (N_2067,N_1994,N_1954);
nand U2068 (N_2068,N_1949,N_1960);
xnor U2069 (N_2069,N_1949,N_1947);
and U2070 (N_2070,N_1902,N_1985);
xor U2071 (N_2071,N_1901,N_1910);
and U2072 (N_2072,N_1939,N_1973);
nor U2073 (N_2073,N_1955,N_1916);
nand U2074 (N_2074,N_1912,N_1987);
nor U2075 (N_2075,N_1938,N_1903);
or U2076 (N_2076,N_1981,N_1962);
xnor U2077 (N_2077,N_1937,N_1904);
nand U2078 (N_2078,N_1991,N_1934);
or U2079 (N_2079,N_1994,N_1970);
and U2080 (N_2080,N_1918,N_1904);
nor U2081 (N_2081,N_1952,N_1993);
and U2082 (N_2082,N_1941,N_1988);
nand U2083 (N_2083,N_1991,N_1968);
nor U2084 (N_2084,N_1920,N_1975);
nand U2085 (N_2085,N_1971,N_1967);
and U2086 (N_2086,N_1936,N_1931);
or U2087 (N_2087,N_1950,N_1973);
or U2088 (N_2088,N_1983,N_1925);
and U2089 (N_2089,N_1938,N_1910);
nor U2090 (N_2090,N_1905,N_1979);
xnor U2091 (N_2091,N_1943,N_1935);
nand U2092 (N_2092,N_1953,N_1994);
and U2093 (N_2093,N_1909,N_1908);
or U2094 (N_2094,N_1907,N_1980);
or U2095 (N_2095,N_1974,N_1978);
and U2096 (N_2096,N_1936,N_1915);
nor U2097 (N_2097,N_1983,N_1978);
nor U2098 (N_2098,N_1918,N_1925);
or U2099 (N_2099,N_1930,N_1946);
or U2100 (N_2100,N_2076,N_2070);
and U2101 (N_2101,N_2044,N_2085);
xnor U2102 (N_2102,N_2030,N_2074);
xnor U2103 (N_2103,N_2035,N_2036);
xnor U2104 (N_2104,N_2053,N_2081);
xor U2105 (N_2105,N_2090,N_2047);
and U2106 (N_2106,N_2057,N_2040);
xor U2107 (N_2107,N_2094,N_2046);
and U2108 (N_2108,N_2002,N_2003);
and U2109 (N_2109,N_2055,N_2089);
or U2110 (N_2110,N_2012,N_2061);
nand U2111 (N_2111,N_2075,N_2005);
nand U2112 (N_2112,N_2095,N_2058);
or U2113 (N_2113,N_2087,N_2099);
or U2114 (N_2114,N_2026,N_2028);
nor U2115 (N_2115,N_2034,N_2060);
and U2116 (N_2116,N_2049,N_2006);
or U2117 (N_2117,N_2007,N_2022);
nor U2118 (N_2118,N_2069,N_2008);
nor U2119 (N_2119,N_2013,N_2097);
nand U2120 (N_2120,N_2079,N_2033);
nand U2121 (N_2121,N_2045,N_2000);
xnor U2122 (N_2122,N_2011,N_2025);
and U2123 (N_2123,N_2086,N_2015);
or U2124 (N_2124,N_2042,N_2043);
xnor U2125 (N_2125,N_2051,N_2029);
xnor U2126 (N_2126,N_2056,N_2004);
nand U2127 (N_2127,N_2072,N_2093);
and U2128 (N_2128,N_2010,N_2024);
nor U2129 (N_2129,N_2050,N_2017);
and U2130 (N_2130,N_2031,N_2071);
xnor U2131 (N_2131,N_2014,N_2059);
nand U2132 (N_2132,N_2048,N_2001);
and U2133 (N_2133,N_2068,N_2066);
nand U2134 (N_2134,N_2027,N_2009);
or U2135 (N_2135,N_2038,N_2091);
xor U2136 (N_2136,N_2067,N_2078);
xnor U2137 (N_2137,N_2019,N_2023);
nand U2138 (N_2138,N_2084,N_2018);
and U2139 (N_2139,N_2021,N_2092);
xor U2140 (N_2140,N_2064,N_2077);
nor U2141 (N_2141,N_2098,N_2041);
and U2142 (N_2142,N_2052,N_2037);
nand U2143 (N_2143,N_2063,N_2062);
or U2144 (N_2144,N_2073,N_2039);
nor U2145 (N_2145,N_2016,N_2020);
xnor U2146 (N_2146,N_2088,N_2054);
or U2147 (N_2147,N_2080,N_2032);
or U2148 (N_2148,N_2083,N_2082);
nand U2149 (N_2149,N_2096,N_2065);
xnor U2150 (N_2150,N_2097,N_2057);
or U2151 (N_2151,N_2051,N_2018);
and U2152 (N_2152,N_2091,N_2036);
or U2153 (N_2153,N_2092,N_2050);
or U2154 (N_2154,N_2048,N_2092);
nand U2155 (N_2155,N_2030,N_2051);
nor U2156 (N_2156,N_2034,N_2049);
xor U2157 (N_2157,N_2014,N_2017);
nor U2158 (N_2158,N_2051,N_2000);
nor U2159 (N_2159,N_2046,N_2059);
nand U2160 (N_2160,N_2032,N_2036);
nor U2161 (N_2161,N_2041,N_2089);
xor U2162 (N_2162,N_2044,N_2094);
xor U2163 (N_2163,N_2090,N_2000);
nor U2164 (N_2164,N_2033,N_2043);
or U2165 (N_2165,N_2055,N_2025);
xnor U2166 (N_2166,N_2024,N_2099);
and U2167 (N_2167,N_2078,N_2025);
xnor U2168 (N_2168,N_2072,N_2078);
or U2169 (N_2169,N_2099,N_2030);
or U2170 (N_2170,N_2007,N_2037);
xnor U2171 (N_2171,N_2078,N_2092);
nor U2172 (N_2172,N_2003,N_2062);
or U2173 (N_2173,N_2046,N_2093);
nor U2174 (N_2174,N_2084,N_2021);
or U2175 (N_2175,N_2059,N_2062);
or U2176 (N_2176,N_2014,N_2078);
nand U2177 (N_2177,N_2055,N_2007);
or U2178 (N_2178,N_2082,N_2017);
and U2179 (N_2179,N_2074,N_2004);
nor U2180 (N_2180,N_2055,N_2057);
xnor U2181 (N_2181,N_2034,N_2096);
and U2182 (N_2182,N_2085,N_2048);
or U2183 (N_2183,N_2017,N_2080);
nand U2184 (N_2184,N_2060,N_2049);
or U2185 (N_2185,N_2039,N_2021);
and U2186 (N_2186,N_2026,N_2098);
xnor U2187 (N_2187,N_2067,N_2025);
xor U2188 (N_2188,N_2066,N_2082);
and U2189 (N_2189,N_2075,N_2081);
and U2190 (N_2190,N_2046,N_2010);
nor U2191 (N_2191,N_2063,N_2001);
nand U2192 (N_2192,N_2079,N_2098);
nor U2193 (N_2193,N_2067,N_2076);
and U2194 (N_2194,N_2070,N_2049);
and U2195 (N_2195,N_2078,N_2084);
nand U2196 (N_2196,N_2019,N_2076);
xor U2197 (N_2197,N_2060,N_2057);
and U2198 (N_2198,N_2074,N_2052);
nand U2199 (N_2199,N_2028,N_2034);
xnor U2200 (N_2200,N_2159,N_2176);
or U2201 (N_2201,N_2126,N_2181);
and U2202 (N_2202,N_2170,N_2192);
nand U2203 (N_2203,N_2153,N_2136);
nor U2204 (N_2204,N_2116,N_2141);
and U2205 (N_2205,N_2133,N_2182);
nor U2206 (N_2206,N_2190,N_2184);
or U2207 (N_2207,N_2169,N_2188);
and U2208 (N_2208,N_2171,N_2131);
or U2209 (N_2209,N_2179,N_2193);
and U2210 (N_2210,N_2160,N_2105);
nand U2211 (N_2211,N_2122,N_2155);
nor U2212 (N_2212,N_2174,N_2137);
or U2213 (N_2213,N_2127,N_2165);
nand U2214 (N_2214,N_2157,N_2120);
xor U2215 (N_2215,N_2140,N_2199);
nand U2216 (N_2216,N_2119,N_2135);
nor U2217 (N_2217,N_2109,N_2146);
or U2218 (N_2218,N_2194,N_2108);
and U2219 (N_2219,N_2134,N_2191);
xnor U2220 (N_2220,N_2123,N_2197);
nor U2221 (N_2221,N_2173,N_2168);
or U2222 (N_2222,N_2145,N_2147);
nor U2223 (N_2223,N_2150,N_2115);
nor U2224 (N_2224,N_2129,N_2189);
and U2225 (N_2225,N_2196,N_2100);
nand U2226 (N_2226,N_2124,N_2198);
or U2227 (N_2227,N_2172,N_2112);
nand U2228 (N_2228,N_2128,N_2164);
and U2229 (N_2229,N_2156,N_2121);
xnor U2230 (N_2230,N_2142,N_2162);
or U2231 (N_2231,N_2186,N_2166);
or U2232 (N_2232,N_2161,N_2178);
and U2233 (N_2233,N_2167,N_2104);
xnor U2234 (N_2234,N_2148,N_2144);
or U2235 (N_2235,N_2101,N_2125);
or U2236 (N_2236,N_2130,N_2103);
nand U2237 (N_2237,N_2158,N_2187);
and U2238 (N_2238,N_2152,N_2114);
xor U2239 (N_2239,N_2177,N_2110);
nand U2240 (N_2240,N_2195,N_2138);
nor U2241 (N_2241,N_2149,N_2107);
and U2242 (N_2242,N_2183,N_2180);
nand U2243 (N_2243,N_2118,N_2151);
xor U2244 (N_2244,N_2154,N_2175);
nand U2245 (N_2245,N_2132,N_2163);
and U2246 (N_2246,N_2106,N_2102);
xnor U2247 (N_2247,N_2113,N_2143);
xnor U2248 (N_2248,N_2185,N_2139);
and U2249 (N_2249,N_2111,N_2117);
nor U2250 (N_2250,N_2132,N_2136);
nor U2251 (N_2251,N_2160,N_2133);
nor U2252 (N_2252,N_2124,N_2186);
or U2253 (N_2253,N_2116,N_2130);
and U2254 (N_2254,N_2138,N_2146);
nand U2255 (N_2255,N_2173,N_2107);
or U2256 (N_2256,N_2176,N_2118);
nand U2257 (N_2257,N_2102,N_2103);
or U2258 (N_2258,N_2184,N_2107);
or U2259 (N_2259,N_2199,N_2114);
or U2260 (N_2260,N_2115,N_2166);
and U2261 (N_2261,N_2159,N_2141);
xnor U2262 (N_2262,N_2190,N_2180);
and U2263 (N_2263,N_2168,N_2187);
xnor U2264 (N_2264,N_2195,N_2123);
nand U2265 (N_2265,N_2159,N_2112);
or U2266 (N_2266,N_2124,N_2177);
nand U2267 (N_2267,N_2178,N_2148);
and U2268 (N_2268,N_2177,N_2111);
or U2269 (N_2269,N_2186,N_2197);
xor U2270 (N_2270,N_2119,N_2183);
and U2271 (N_2271,N_2169,N_2115);
or U2272 (N_2272,N_2155,N_2165);
nand U2273 (N_2273,N_2172,N_2129);
or U2274 (N_2274,N_2159,N_2124);
nor U2275 (N_2275,N_2160,N_2126);
or U2276 (N_2276,N_2193,N_2161);
or U2277 (N_2277,N_2196,N_2173);
and U2278 (N_2278,N_2141,N_2173);
and U2279 (N_2279,N_2145,N_2149);
or U2280 (N_2280,N_2164,N_2172);
and U2281 (N_2281,N_2170,N_2153);
nor U2282 (N_2282,N_2152,N_2115);
nor U2283 (N_2283,N_2151,N_2144);
xor U2284 (N_2284,N_2190,N_2116);
and U2285 (N_2285,N_2101,N_2107);
and U2286 (N_2286,N_2148,N_2131);
nor U2287 (N_2287,N_2191,N_2104);
or U2288 (N_2288,N_2181,N_2106);
nand U2289 (N_2289,N_2143,N_2123);
xor U2290 (N_2290,N_2189,N_2145);
and U2291 (N_2291,N_2166,N_2144);
nor U2292 (N_2292,N_2113,N_2191);
xor U2293 (N_2293,N_2196,N_2197);
nand U2294 (N_2294,N_2163,N_2179);
and U2295 (N_2295,N_2151,N_2104);
nand U2296 (N_2296,N_2115,N_2144);
nand U2297 (N_2297,N_2195,N_2147);
and U2298 (N_2298,N_2108,N_2191);
or U2299 (N_2299,N_2170,N_2133);
nor U2300 (N_2300,N_2227,N_2215);
and U2301 (N_2301,N_2274,N_2263);
or U2302 (N_2302,N_2270,N_2290);
xnor U2303 (N_2303,N_2241,N_2226);
nor U2304 (N_2304,N_2209,N_2228);
and U2305 (N_2305,N_2295,N_2206);
xor U2306 (N_2306,N_2278,N_2255);
and U2307 (N_2307,N_2266,N_2254);
nor U2308 (N_2308,N_2207,N_2285);
xnor U2309 (N_2309,N_2281,N_2225);
nor U2310 (N_2310,N_2297,N_2247);
nor U2311 (N_2311,N_2298,N_2265);
nor U2312 (N_2312,N_2224,N_2286);
and U2313 (N_2313,N_2212,N_2240);
nor U2314 (N_2314,N_2214,N_2268);
or U2315 (N_2315,N_2252,N_2279);
or U2316 (N_2316,N_2259,N_2291);
xor U2317 (N_2317,N_2216,N_2229);
nand U2318 (N_2318,N_2210,N_2299);
nor U2319 (N_2319,N_2211,N_2235);
nand U2320 (N_2320,N_2269,N_2288);
and U2321 (N_2321,N_2208,N_2292);
nand U2322 (N_2322,N_2251,N_2223);
xnor U2323 (N_2323,N_2239,N_2230);
or U2324 (N_2324,N_2205,N_2284);
nand U2325 (N_2325,N_2253,N_2250);
nand U2326 (N_2326,N_2232,N_2233);
xor U2327 (N_2327,N_2280,N_2258);
and U2328 (N_2328,N_2293,N_2237);
and U2329 (N_2329,N_2244,N_2242);
and U2330 (N_2330,N_2248,N_2236);
or U2331 (N_2331,N_2217,N_2200);
nand U2332 (N_2332,N_2203,N_2282);
xor U2333 (N_2333,N_2246,N_2218);
and U2334 (N_2334,N_2243,N_2272);
xnor U2335 (N_2335,N_2275,N_2245);
or U2336 (N_2336,N_2289,N_2201);
and U2337 (N_2337,N_2267,N_2231);
nand U2338 (N_2338,N_2249,N_2238);
and U2339 (N_2339,N_2287,N_2221);
xor U2340 (N_2340,N_2262,N_2277);
nand U2341 (N_2341,N_2222,N_2219);
nor U2342 (N_2342,N_2204,N_2260);
xnor U2343 (N_2343,N_2296,N_2264);
nor U2344 (N_2344,N_2256,N_2213);
xnor U2345 (N_2345,N_2234,N_2271);
xor U2346 (N_2346,N_2257,N_2294);
nor U2347 (N_2347,N_2220,N_2283);
and U2348 (N_2348,N_2276,N_2261);
and U2349 (N_2349,N_2273,N_2202);
and U2350 (N_2350,N_2207,N_2238);
and U2351 (N_2351,N_2241,N_2286);
nand U2352 (N_2352,N_2258,N_2202);
xnor U2353 (N_2353,N_2281,N_2284);
or U2354 (N_2354,N_2244,N_2258);
nor U2355 (N_2355,N_2203,N_2287);
xor U2356 (N_2356,N_2211,N_2284);
nand U2357 (N_2357,N_2232,N_2222);
nand U2358 (N_2358,N_2262,N_2233);
nand U2359 (N_2359,N_2230,N_2273);
nand U2360 (N_2360,N_2233,N_2207);
nor U2361 (N_2361,N_2256,N_2265);
xor U2362 (N_2362,N_2212,N_2295);
or U2363 (N_2363,N_2282,N_2269);
xnor U2364 (N_2364,N_2261,N_2215);
xor U2365 (N_2365,N_2279,N_2227);
xor U2366 (N_2366,N_2200,N_2263);
nor U2367 (N_2367,N_2206,N_2248);
or U2368 (N_2368,N_2260,N_2230);
or U2369 (N_2369,N_2227,N_2290);
and U2370 (N_2370,N_2236,N_2208);
nor U2371 (N_2371,N_2247,N_2218);
xnor U2372 (N_2372,N_2223,N_2281);
nor U2373 (N_2373,N_2212,N_2266);
and U2374 (N_2374,N_2234,N_2259);
nor U2375 (N_2375,N_2268,N_2210);
xor U2376 (N_2376,N_2290,N_2250);
nand U2377 (N_2377,N_2203,N_2292);
nor U2378 (N_2378,N_2227,N_2277);
nand U2379 (N_2379,N_2296,N_2274);
xnor U2380 (N_2380,N_2266,N_2282);
xnor U2381 (N_2381,N_2246,N_2259);
xor U2382 (N_2382,N_2231,N_2251);
and U2383 (N_2383,N_2279,N_2248);
nor U2384 (N_2384,N_2236,N_2223);
xor U2385 (N_2385,N_2279,N_2265);
and U2386 (N_2386,N_2263,N_2244);
and U2387 (N_2387,N_2282,N_2273);
or U2388 (N_2388,N_2293,N_2282);
xnor U2389 (N_2389,N_2209,N_2240);
and U2390 (N_2390,N_2265,N_2225);
nor U2391 (N_2391,N_2248,N_2283);
nor U2392 (N_2392,N_2295,N_2222);
nand U2393 (N_2393,N_2283,N_2240);
xnor U2394 (N_2394,N_2268,N_2225);
or U2395 (N_2395,N_2283,N_2291);
xnor U2396 (N_2396,N_2240,N_2232);
nand U2397 (N_2397,N_2216,N_2293);
or U2398 (N_2398,N_2233,N_2203);
xor U2399 (N_2399,N_2220,N_2233);
nor U2400 (N_2400,N_2354,N_2340);
nand U2401 (N_2401,N_2380,N_2373);
nor U2402 (N_2402,N_2343,N_2391);
nor U2403 (N_2403,N_2345,N_2344);
nor U2404 (N_2404,N_2311,N_2365);
and U2405 (N_2405,N_2385,N_2336);
nand U2406 (N_2406,N_2337,N_2399);
or U2407 (N_2407,N_2359,N_2371);
nor U2408 (N_2408,N_2375,N_2316);
nand U2409 (N_2409,N_2321,N_2326);
and U2410 (N_2410,N_2388,N_2308);
xor U2411 (N_2411,N_2363,N_2305);
nand U2412 (N_2412,N_2324,N_2333);
nor U2413 (N_2413,N_2335,N_2322);
and U2414 (N_2414,N_2367,N_2353);
nand U2415 (N_2415,N_2355,N_2352);
nand U2416 (N_2416,N_2309,N_2329);
nor U2417 (N_2417,N_2376,N_2350);
and U2418 (N_2418,N_2398,N_2395);
or U2419 (N_2419,N_2392,N_2341);
and U2420 (N_2420,N_2379,N_2307);
or U2421 (N_2421,N_2319,N_2384);
xor U2422 (N_2422,N_2387,N_2342);
nand U2423 (N_2423,N_2323,N_2347);
and U2424 (N_2424,N_2369,N_2349);
nor U2425 (N_2425,N_2358,N_2368);
xor U2426 (N_2426,N_2317,N_2377);
nand U2427 (N_2427,N_2312,N_2300);
nand U2428 (N_2428,N_2310,N_2390);
xor U2429 (N_2429,N_2383,N_2304);
nand U2430 (N_2430,N_2346,N_2378);
nor U2431 (N_2431,N_2364,N_2382);
or U2432 (N_2432,N_2348,N_2331);
and U2433 (N_2433,N_2394,N_2332);
and U2434 (N_2434,N_2318,N_2361);
xnor U2435 (N_2435,N_2374,N_2351);
xor U2436 (N_2436,N_2302,N_2397);
and U2437 (N_2437,N_2328,N_2320);
nor U2438 (N_2438,N_2315,N_2372);
xnor U2439 (N_2439,N_2370,N_2356);
and U2440 (N_2440,N_2330,N_2301);
and U2441 (N_2441,N_2396,N_2334);
and U2442 (N_2442,N_2360,N_2306);
or U2443 (N_2443,N_2327,N_2389);
nor U2444 (N_2444,N_2313,N_2381);
or U2445 (N_2445,N_2386,N_2314);
or U2446 (N_2446,N_2338,N_2362);
nand U2447 (N_2447,N_2366,N_2325);
nand U2448 (N_2448,N_2339,N_2357);
nand U2449 (N_2449,N_2303,N_2393);
nand U2450 (N_2450,N_2337,N_2376);
or U2451 (N_2451,N_2300,N_2357);
or U2452 (N_2452,N_2357,N_2327);
or U2453 (N_2453,N_2312,N_2308);
and U2454 (N_2454,N_2319,N_2325);
nand U2455 (N_2455,N_2319,N_2361);
and U2456 (N_2456,N_2338,N_2360);
or U2457 (N_2457,N_2314,N_2394);
xnor U2458 (N_2458,N_2337,N_2387);
xor U2459 (N_2459,N_2358,N_2317);
nor U2460 (N_2460,N_2378,N_2332);
xnor U2461 (N_2461,N_2332,N_2302);
nor U2462 (N_2462,N_2396,N_2351);
nand U2463 (N_2463,N_2369,N_2321);
nand U2464 (N_2464,N_2366,N_2349);
or U2465 (N_2465,N_2310,N_2365);
xor U2466 (N_2466,N_2396,N_2322);
or U2467 (N_2467,N_2347,N_2364);
xor U2468 (N_2468,N_2365,N_2330);
xor U2469 (N_2469,N_2369,N_2362);
xnor U2470 (N_2470,N_2336,N_2356);
nand U2471 (N_2471,N_2361,N_2312);
and U2472 (N_2472,N_2376,N_2353);
nor U2473 (N_2473,N_2325,N_2362);
or U2474 (N_2474,N_2383,N_2399);
or U2475 (N_2475,N_2363,N_2375);
and U2476 (N_2476,N_2361,N_2351);
or U2477 (N_2477,N_2395,N_2339);
nor U2478 (N_2478,N_2394,N_2320);
xnor U2479 (N_2479,N_2360,N_2352);
xor U2480 (N_2480,N_2342,N_2337);
xor U2481 (N_2481,N_2365,N_2360);
nand U2482 (N_2482,N_2390,N_2307);
xor U2483 (N_2483,N_2354,N_2386);
and U2484 (N_2484,N_2321,N_2362);
nor U2485 (N_2485,N_2306,N_2356);
nor U2486 (N_2486,N_2355,N_2321);
and U2487 (N_2487,N_2363,N_2393);
and U2488 (N_2488,N_2327,N_2391);
nand U2489 (N_2489,N_2319,N_2349);
or U2490 (N_2490,N_2351,N_2312);
xor U2491 (N_2491,N_2358,N_2338);
nor U2492 (N_2492,N_2300,N_2319);
and U2493 (N_2493,N_2305,N_2315);
and U2494 (N_2494,N_2377,N_2331);
xnor U2495 (N_2495,N_2348,N_2329);
or U2496 (N_2496,N_2311,N_2351);
xor U2497 (N_2497,N_2320,N_2325);
nor U2498 (N_2498,N_2302,N_2314);
nand U2499 (N_2499,N_2332,N_2371);
nor U2500 (N_2500,N_2400,N_2428);
nand U2501 (N_2501,N_2461,N_2485);
nand U2502 (N_2502,N_2487,N_2440);
nor U2503 (N_2503,N_2430,N_2481);
xor U2504 (N_2504,N_2410,N_2490);
xor U2505 (N_2505,N_2497,N_2429);
nor U2506 (N_2506,N_2488,N_2418);
nor U2507 (N_2507,N_2435,N_2427);
nor U2508 (N_2508,N_2434,N_2482);
nor U2509 (N_2509,N_2407,N_2443);
or U2510 (N_2510,N_2456,N_2498);
xnor U2511 (N_2511,N_2408,N_2425);
nor U2512 (N_2512,N_2494,N_2477);
or U2513 (N_2513,N_2475,N_2449);
or U2514 (N_2514,N_2484,N_2458);
or U2515 (N_2515,N_2471,N_2433);
and U2516 (N_2516,N_2416,N_2448);
and U2517 (N_2517,N_2415,N_2401);
nand U2518 (N_2518,N_2439,N_2441);
nor U2519 (N_2519,N_2414,N_2432);
nand U2520 (N_2520,N_2499,N_2413);
nand U2521 (N_2521,N_2451,N_2466);
and U2522 (N_2522,N_2454,N_2495);
nor U2523 (N_2523,N_2460,N_2480);
nand U2524 (N_2524,N_2459,N_2476);
nand U2525 (N_2525,N_2404,N_2403);
and U2526 (N_2526,N_2492,N_2457);
nand U2527 (N_2527,N_2470,N_2455);
nor U2528 (N_2528,N_2442,N_2496);
nand U2529 (N_2529,N_2437,N_2468);
or U2530 (N_2530,N_2447,N_2462);
or U2531 (N_2531,N_2467,N_2411);
nor U2532 (N_2532,N_2465,N_2417);
and U2533 (N_2533,N_2446,N_2420);
and U2534 (N_2534,N_2444,N_2486);
nand U2535 (N_2535,N_2450,N_2419);
nand U2536 (N_2536,N_2422,N_2483);
nand U2537 (N_2537,N_2453,N_2426);
xnor U2538 (N_2538,N_2473,N_2445);
nand U2539 (N_2539,N_2452,N_2421);
xnor U2540 (N_2540,N_2405,N_2478);
nand U2541 (N_2541,N_2474,N_2469);
nand U2542 (N_2542,N_2412,N_2431);
and U2543 (N_2543,N_2479,N_2423);
or U2544 (N_2544,N_2491,N_2436);
xor U2545 (N_2545,N_2424,N_2472);
or U2546 (N_2546,N_2463,N_2409);
xor U2547 (N_2547,N_2489,N_2464);
and U2548 (N_2548,N_2402,N_2406);
nand U2549 (N_2549,N_2493,N_2438);
and U2550 (N_2550,N_2433,N_2480);
and U2551 (N_2551,N_2481,N_2495);
or U2552 (N_2552,N_2466,N_2411);
nor U2553 (N_2553,N_2426,N_2465);
nand U2554 (N_2554,N_2450,N_2481);
or U2555 (N_2555,N_2424,N_2490);
nor U2556 (N_2556,N_2420,N_2400);
nand U2557 (N_2557,N_2404,N_2405);
nor U2558 (N_2558,N_2468,N_2435);
or U2559 (N_2559,N_2489,N_2493);
or U2560 (N_2560,N_2401,N_2408);
and U2561 (N_2561,N_2437,N_2424);
and U2562 (N_2562,N_2452,N_2418);
and U2563 (N_2563,N_2499,N_2410);
nand U2564 (N_2564,N_2472,N_2439);
and U2565 (N_2565,N_2442,N_2439);
nand U2566 (N_2566,N_2498,N_2478);
nor U2567 (N_2567,N_2476,N_2488);
nor U2568 (N_2568,N_2425,N_2432);
or U2569 (N_2569,N_2462,N_2467);
or U2570 (N_2570,N_2467,N_2463);
nand U2571 (N_2571,N_2467,N_2401);
and U2572 (N_2572,N_2487,N_2498);
or U2573 (N_2573,N_2401,N_2461);
xor U2574 (N_2574,N_2481,N_2483);
or U2575 (N_2575,N_2400,N_2425);
or U2576 (N_2576,N_2457,N_2445);
and U2577 (N_2577,N_2482,N_2485);
or U2578 (N_2578,N_2468,N_2400);
and U2579 (N_2579,N_2416,N_2459);
xnor U2580 (N_2580,N_2427,N_2464);
nand U2581 (N_2581,N_2403,N_2443);
nand U2582 (N_2582,N_2480,N_2475);
and U2583 (N_2583,N_2409,N_2400);
nand U2584 (N_2584,N_2468,N_2408);
and U2585 (N_2585,N_2466,N_2490);
and U2586 (N_2586,N_2439,N_2490);
xor U2587 (N_2587,N_2420,N_2414);
nor U2588 (N_2588,N_2436,N_2469);
nor U2589 (N_2589,N_2465,N_2415);
xor U2590 (N_2590,N_2403,N_2482);
nand U2591 (N_2591,N_2401,N_2487);
and U2592 (N_2592,N_2447,N_2423);
and U2593 (N_2593,N_2478,N_2438);
nor U2594 (N_2594,N_2428,N_2493);
xor U2595 (N_2595,N_2468,N_2444);
nor U2596 (N_2596,N_2412,N_2480);
or U2597 (N_2597,N_2477,N_2487);
nor U2598 (N_2598,N_2419,N_2451);
or U2599 (N_2599,N_2488,N_2498);
nor U2600 (N_2600,N_2592,N_2571);
nor U2601 (N_2601,N_2520,N_2540);
and U2602 (N_2602,N_2538,N_2503);
or U2603 (N_2603,N_2553,N_2563);
nor U2604 (N_2604,N_2545,N_2599);
nor U2605 (N_2605,N_2574,N_2586);
and U2606 (N_2606,N_2550,N_2513);
or U2607 (N_2607,N_2532,N_2502);
or U2608 (N_2608,N_2544,N_2557);
and U2609 (N_2609,N_2508,N_2556);
nand U2610 (N_2610,N_2512,N_2579);
nand U2611 (N_2611,N_2506,N_2547);
nand U2612 (N_2612,N_2551,N_2581);
nand U2613 (N_2613,N_2504,N_2577);
nor U2614 (N_2614,N_2535,N_2568);
nand U2615 (N_2615,N_2584,N_2505);
nand U2616 (N_2616,N_2522,N_2548);
nand U2617 (N_2617,N_2530,N_2541);
nand U2618 (N_2618,N_2555,N_2539);
and U2619 (N_2619,N_2596,N_2561);
and U2620 (N_2620,N_2582,N_2560);
and U2621 (N_2621,N_2500,N_2529);
nand U2622 (N_2622,N_2507,N_2572);
nand U2623 (N_2623,N_2583,N_2589);
or U2624 (N_2624,N_2569,N_2598);
or U2625 (N_2625,N_2591,N_2587);
and U2626 (N_2626,N_2570,N_2597);
nor U2627 (N_2627,N_2515,N_2527);
or U2628 (N_2628,N_2509,N_2558);
xnor U2629 (N_2629,N_2595,N_2590);
nand U2630 (N_2630,N_2524,N_2542);
nand U2631 (N_2631,N_2501,N_2531);
nor U2632 (N_2632,N_2537,N_2528);
or U2633 (N_2633,N_2593,N_2576);
nor U2634 (N_2634,N_2546,N_2575);
and U2635 (N_2635,N_2518,N_2578);
xnor U2636 (N_2636,N_2559,N_2534);
or U2637 (N_2637,N_2562,N_2565);
or U2638 (N_2638,N_2516,N_2585);
and U2639 (N_2639,N_2549,N_2543);
or U2640 (N_2640,N_2523,N_2521);
and U2641 (N_2641,N_2552,N_2580);
and U2642 (N_2642,N_2511,N_2510);
nor U2643 (N_2643,N_2566,N_2517);
and U2644 (N_2644,N_2567,N_2525);
and U2645 (N_2645,N_2573,N_2519);
nor U2646 (N_2646,N_2564,N_2536);
nor U2647 (N_2647,N_2514,N_2594);
and U2648 (N_2648,N_2588,N_2554);
and U2649 (N_2649,N_2533,N_2526);
nand U2650 (N_2650,N_2574,N_2506);
and U2651 (N_2651,N_2585,N_2590);
or U2652 (N_2652,N_2531,N_2594);
or U2653 (N_2653,N_2502,N_2528);
nor U2654 (N_2654,N_2521,N_2543);
nand U2655 (N_2655,N_2568,N_2547);
and U2656 (N_2656,N_2589,N_2504);
and U2657 (N_2657,N_2526,N_2578);
or U2658 (N_2658,N_2542,N_2540);
or U2659 (N_2659,N_2528,N_2507);
nand U2660 (N_2660,N_2506,N_2565);
xnor U2661 (N_2661,N_2599,N_2526);
or U2662 (N_2662,N_2543,N_2503);
nand U2663 (N_2663,N_2520,N_2599);
nor U2664 (N_2664,N_2516,N_2548);
nand U2665 (N_2665,N_2525,N_2518);
or U2666 (N_2666,N_2557,N_2515);
xor U2667 (N_2667,N_2522,N_2564);
and U2668 (N_2668,N_2540,N_2544);
xor U2669 (N_2669,N_2506,N_2501);
nor U2670 (N_2670,N_2549,N_2590);
and U2671 (N_2671,N_2513,N_2549);
nand U2672 (N_2672,N_2586,N_2522);
nor U2673 (N_2673,N_2537,N_2584);
nand U2674 (N_2674,N_2506,N_2548);
and U2675 (N_2675,N_2596,N_2591);
and U2676 (N_2676,N_2566,N_2575);
and U2677 (N_2677,N_2563,N_2508);
or U2678 (N_2678,N_2510,N_2588);
nor U2679 (N_2679,N_2557,N_2549);
and U2680 (N_2680,N_2574,N_2593);
nor U2681 (N_2681,N_2545,N_2575);
nand U2682 (N_2682,N_2556,N_2576);
or U2683 (N_2683,N_2515,N_2552);
nand U2684 (N_2684,N_2594,N_2524);
or U2685 (N_2685,N_2592,N_2532);
nor U2686 (N_2686,N_2584,N_2525);
nand U2687 (N_2687,N_2573,N_2557);
or U2688 (N_2688,N_2559,N_2539);
xor U2689 (N_2689,N_2519,N_2569);
nor U2690 (N_2690,N_2597,N_2510);
and U2691 (N_2691,N_2596,N_2534);
nor U2692 (N_2692,N_2539,N_2567);
or U2693 (N_2693,N_2526,N_2548);
and U2694 (N_2694,N_2560,N_2500);
xnor U2695 (N_2695,N_2544,N_2508);
nand U2696 (N_2696,N_2590,N_2577);
and U2697 (N_2697,N_2557,N_2529);
or U2698 (N_2698,N_2539,N_2525);
nor U2699 (N_2699,N_2555,N_2595);
or U2700 (N_2700,N_2622,N_2663);
and U2701 (N_2701,N_2685,N_2618);
and U2702 (N_2702,N_2621,N_2698);
nand U2703 (N_2703,N_2649,N_2694);
or U2704 (N_2704,N_2651,N_2690);
xor U2705 (N_2705,N_2607,N_2605);
or U2706 (N_2706,N_2627,N_2639);
xnor U2707 (N_2707,N_2643,N_2667);
or U2708 (N_2708,N_2680,N_2620);
or U2709 (N_2709,N_2682,N_2606);
nand U2710 (N_2710,N_2648,N_2633);
nor U2711 (N_2711,N_2616,N_2637);
and U2712 (N_2712,N_2688,N_2626);
nand U2713 (N_2713,N_2640,N_2679);
and U2714 (N_2714,N_2624,N_2611);
nor U2715 (N_2715,N_2614,N_2656);
xor U2716 (N_2716,N_2675,N_2666);
nand U2717 (N_2717,N_2604,N_2686);
or U2718 (N_2718,N_2670,N_2600);
and U2719 (N_2719,N_2625,N_2684);
and U2720 (N_2720,N_2662,N_2691);
xnor U2721 (N_2721,N_2631,N_2602);
and U2722 (N_2722,N_2623,N_2659);
or U2723 (N_2723,N_2635,N_2664);
and U2724 (N_2724,N_2653,N_2661);
nand U2725 (N_2725,N_2668,N_2617);
and U2726 (N_2726,N_2687,N_2636);
and U2727 (N_2727,N_2655,N_2693);
xnor U2728 (N_2728,N_2645,N_2677);
or U2729 (N_2729,N_2619,N_2658);
and U2730 (N_2730,N_2613,N_2609);
xnor U2731 (N_2731,N_2695,N_2657);
xor U2732 (N_2732,N_2612,N_2654);
nand U2733 (N_2733,N_2672,N_2660);
nor U2734 (N_2734,N_2696,N_2674);
or U2735 (N_2735,N_2683,N_2634);
xnor U2736 (N_2736,N_2652,N_2608);
xnor U2737 (N_2737,N_2699,N_2676);
and U2738 (N_2738,N_2610,N_2650);
or U2739 (N_2739,N_2615,N_2646);
xor U2740 (N_2740,N_2630,N_2628);
and U2741 (N_2741,N_2642,N_2665);
nand U2742 (N_2742,N_2641,N_2692);
and U2743 (N_2743,N_2638,N_2671);
or U2744 (N_2744,N_2673,N_2681);
nor U2745 (N_2745,N_2689,N_2697);
nand U2746 (N_2746,N_2644,N_2678);
xor U2747 (N_2747,N_2603,N_2669);
nor U2748 (N_2748,N_2601,N_2647);
nor U2749 (N_2749,N_2629,N_2632);
nand U2750 (N_2750,N_2612,N_2695);
nand U2751 (N_2751,N_2697,N_2645);
nor U2752 (N_2752,N_2667,N_2679);
nor U2753 (N_2753,N_2685,N_2600);
xnor U2754 (N_2754,N_2624,N_2625);
nand U2755 (N_2755,N_2690,N_2696);
xnor U2756 (N_2756,N_2674,N_2693);
and U2757 (N_2757,N_2609,N_2654);
xor U2758 (N_2758,N_2659,N_2669);
or U2759 (N_2759,N_2692,N_2652);
nor U2760 (N_2760,N_2666,N_2601);
and U2761 (N_2761,N_2639,N_2695);
nor U2762 (N_2762,N_2652,N_2630);
or U2763 (N_2763,N_2645,N_2680);
nand U2764 (N_2764,N_2641,N_2659);
or U2765 (N_2765,N_2605,N_2638);
or U2766 (N_2766,N_2651,N_2620);
and U2767 (N_2767,N_2646,N_2688);
and U2768 (N_2768,N_2601,N_2661);
nor U2769 (N_2769,N_2600,N_2638);
xnor U2770 (N_2770,N_2606,N_2675);
and U2771 (N_2771,N_2676,N_2687);
nor U2772 (N_2772,N_2645,N_2619);
xor U2773 (N_2773,N_2620,N_2656);
and U2774 (N_2774,N_2648,N_2695);
and U2775 (N_2775,N_2684,N_2621);
xnor U2776 (N_2776,N_2622,N_2623);
nand U2777 (N_2777,N_2630,N_2649);
nand U2778 (N_2778,N_2657,N_2607);
nand U2779 (N_2779,N_2647,N_2648);
xnor U2780 (N_2780,N_2675,N_2677);
nor U2781 (N_2781,N_2656,N_2616);
nor U2782 (N_2782,N_2649,N_2677);
and U2783 (N_2783,N_2632,N_2641);
nor U2784 (N_2784,N_2638,N_2641);
nand U2785 (N_2785,N_2652,N_2635);
or U2786 (N_2786,N_2607,N_2678);
and U2787 (N_2787,N_2675,N_2603);
nand U2788 (N_2788,N_2643,N_2682);
or U2789 (N_2789,N_2642,N_2657);
nor U2790 (N_2790,N_2603,N_2646);
xnor U2791 (N_2791,N_2686,N_2638);
and U2792 (N_2792,N_2607,N_2637);
or U2793 (N_2793,N_2621,N_2685);
or U2794 (N_2794,N_2674,N_2639);
and U2795 (N_2795,N_2695,N_2608);
or U2796 (N_2796,N_2641,N_2649);
or U2797 (N_2797,N_2683,N_2633);
nor U2798 (N_2798,N_2668,N_2654);
and U2799 (N_2799,N_2632,N_2671);
or U2800 (N_2800,N_2771,N_2735);
nand U2801 (N_2801,N_2719,N_2728);
and U2802 (N_2802,N_2713,N_2737);
nand U2803 (N_2803,N_2712,N_2784);
and U2804 (N_2804,N_2791,N_2703);
nor U2805 (N_2805,N_2774,N_2776);
nor U2806 (N_2806,N_2792,N_2757);
nand U2807 (N_2807,N_2781,N_2724);
xor U2808 (N_2808,N_2708,N_2755);
nand U2809 (N_2809,N_2782,N_2716);
xnor U2810 (N_2810,N_2778,N_2769);
nor U2811 (N_2811,N_2785,N_2794);
or U2812 (N_2812,N_2715,N_2718);
and U2813 (N_2813,N_2752,N_2783);
nand U2814 (N_2814,N_2761,N_2707);
or U2815 (N_2815,N_2738,N_2779);
and U2816 (N_2816,N_2705,N_2709);
and U2817 (N_2817,N_2795,N_2740);
or U2818 (N_2818,N_2727,N_2797);
and U2819 (N_2819,N_2704,N_2788);
and U2820 (N_2820,N_2762,N_2750);
or U2821 (N_2821,N_2736,N_2786);
nor U2822 (N_2822,N_2729,N_2717);
nand U2823 (N_2823,N_2700,N_2766);
or U2824 (N_2824,N_2739,N_2722);
or U2825 (N_2825,N_2725,N_2731);
or U2826 (N_2826,N_2772,N_2799);
nand U2827 (N_2827,N_2730,N_2726);
xnor U2828 (N_2828,N_2777,N_2796);
or U2829 (N_2829,N_2734,N_2758);
nor U2830 (N_2830,N_2751,N_2741);
and U2831 (N_2831,N_2787,N_2790);
and U2832 (N_2832,N_2793,N_2773);
xnor U2833 (N_2833,N_2720,N_2780);
nor U2834 (N_2834,N_2742,N_2768);
xor U2835 (N_2835,N_2754,N_2711);
nand U2836 (N_2836,N_2759,N_2764);
or U2837 (N_2837,N_2714,N_2753);
nor U2838 (N_2838,N_2733,N_2763);
or U2839 (N_2839,N_2721,N_2747);
nand U2840 (N_2840,N_2748,N_2749);
and U2841 (N_2841,N_2756,N_2798);
and U2842 (N_2842,N_2745,N_2710);
and U2843 (N_2843,N_2744,N_2723);
and U2844 (N_2844,N_2789,N_2746);
and U2845 (N_2845,N_2701,N_2760);
and U2846 (N_2846,N_2765,N_2767);
or U2847 (N_2847,N_2702,N_2743);
nand U2848 (N_2848,N_2770,N_2706);
and U2849 (N_2849,N_2732,N_2775);
or U2850 (N_2850,N_2744,N_2790);
and U2851 (N_2851,N_2712,N_2750);
and U2852 (N_2852,N_2731,N_2784);
xnor U2853 (N_2853,N_2777,N_2700);
or U2854 (N_2854,N_2751,N_2791);
xnor U2855 (N_2855,N_2761,N_2788);
and U2856 (N_2856,N_2739,N_2784);
and U2857 (N_2857,N_2758,N_2737);
xor U2858 (N_2858,N_2714,N_2739);
or U2859 (N_2859,N_2713,N_2789);
nor U2860 (N_2860,N_2733,N_2747);
or U2861 (N_2861,N_2735,N_2750);
xnor U2862 (N_2862,N_2741,N_2711);
nand U2863 (N_2863,N_2713,N_2757);
and U2864 (N_2864,N_2717,N_2723);
nand U2865 (N_2865,N_2785,N_2730);
nor U2866 (N_2866,N_2787,N_2765);
nand U2867 (N_2867,N_2793,N_2718);
and U2868 (N_2868,N_2701,N_2758);
and U2869 (N_2869,N_2773,N_2708);
xor U2870 (N_2870,N_2770,N_2725);
and U2871 (N_2871,N_2791,N_2733);
nand U2872 (N_2872,N_2716,N_2742);
nor U2873 (N_2873,N_2764,N_2704);
or U2874 (N_2874,N_2785,N_2728);
or U2875 (N_2875,N_2700,N_2733);
xnor U2876 (N_2876,N_2783,N_2781);
nor U2877 (N_2877,N_2712,N_2721);
or U2878 (N_2878,N_2754,N_2753);
or U2879 (N_2879,N_2733,N_2796);
nand U2880 (N_2880,N_2787,N_2785);
nand U2881 (N_2881,N_2725,N_2716);
xnor U2882 (N_2882,N_2791,N_2767);
nor U2883 (N_2883,N_2774,N_2789);
nand U2884 (N_2884,N_2706,N_2776);
or U2885 (N_2885,N_2753,N_2774);
xor U2886 (N_2886,N_2783,N_2753);
or U2887 (N_2887,N_2792,N_2797);
or U2888 (N_2888,N_2776,N_2724);
xnor U2889 (N_2889,N_2735,N_2729);
and U2890 (N_2890,N_2705,N_2746);
nand U2891 (N_2891,N_2775,N_2761);
or U2892 (N_2892,N_2720,N_2789);
nand U2893 (N_2893,N_2700,N_2763);
and U2894 (N_2894,N_2754,N_2755);
and U2895 (N_2895,N_2762,N_2788);
or U2896 (N_2896,N_2737,N_2771);
xor U2897 (N_2897,N_2799,N_2713);
nor U2898 (N_2898,N_2733,N_2776);
nor U2899 (N_2899,N_2766,N_2781);
and U2900 (N_2900,N_2803,N_2893);
nand U2901 (N_2901,N_2843,N_2811);
xnor U2902 (N_2902,N_2875,N_2819);
or U2903 (N_2903,N_2810,N_2822);
and U2904 (N_2904,N_2885,N_2823);
and U2905 (N_2905,N_2820,N_2897);
nand U2906 (N_2906,N_2880,N_2829);
nand U2907 (N_2907,N_2848,N_2881);
xor U2908 (N_2908,N_2864,N_2835);
or U2909 (N_2909,N_2806,N_2802);
and U2910 (N_2910,N_2895,N_2812);
xor U2911 (N_2911,N_2873,N_2852);
nand U2912 (N_2912,N_2827,N_2872);
or U2913 (N_2913,N_2834,N_2836);
xor U2914 (N_2914,N_2861,N_2825);
or U2915 (N_2915,N_2866,N_2874);
xor U2916 (N_2916,N_2883,N_2869);
nor U2917 (N_2917,N_2804,N_2830);
nor U2918 (N_2918,N_2847,N_2809);
and U2919 (N_2919,N_2807,N_2894);
and U2920 (N_2920,N_2832,N_2800);
nand U2921 (N_2921,N_2886,N_2887);
and U2922 (N_2922,N_2817,N_2840);
xnor U2923 (N_2923,N_2862,N_2871);
nor U2924 (N_2924,N_2853,N_2870);
xnor U2925 (N_2925,N_2876,N_2860);
xnor U2926 (N_2926,N_2867,N_2898);
and U2927 (N_2927,N_2816,N_2808);
nand U2928 (N_2928,N_2859,N_2828);
or U2929 (N_2929,N_2814,N_2839);
nand U2930 (N_2930,N_2824,N_2899);
or U2931 (N_2931,N_2856,N_2882);
or U2932 (N_2932,N_2879,N_2858);
and U2933 (N_2933,N_2838,N_2877);
and U2934 (N_2934,N_2850,N_2896);
or U2935 (N_2935,N_2855,N_2818);
and U2936 (N_2936,N_2846,N_2842);
nor U2937 (N_2937,N_2865,N_2849);
nor U2938 (N_2938,N_2813,N_2837);
xor U2939 (N_2939,N_2851,N_2857);
nor U2940 (N_2940,N_2854,N_2844);
and U2941 (N_2941,N_2831,N_2801);
xnor U2942 (N_2942,N_2878,N_2821);
nand U2943 (N_2943,N_2892,N_2841);
nor U2944 (N_2944,N_2833,N_2891);
or U2945 (N_2945,N_2845,N_2890);
nor U2946 (N_2946,N_2826,N_2863);
xor U2947 (N_2947,N_2868,N_2815);
nand U2948 (N_2948,N_2889,N_2884);
or U2949 (N_2949,N_2805,N_2888);
or U2950 (N_2950,N_2892,N_2826);
or U2951 (N_2951,N_2853,N_2886);
or U2952 (N_2952,N_2897,N_2819);
xor U2953 (N_2953,N_2863,N_2839);
nand U2954 (N_2954,N_2895,N_2897);
xnor U2955 (N_2955,N_2833,N_2846);
nand U2956 (N_2956,N_2890,N_2885);
and U2957 (N_2957,N_2841,N_2884);
and U2958 (N_2958,N_2829,N_2843);
nor U2959 (N_2959,N_2835,N_2873);
nand U2960 (N_2960,N_2818,N_2878);
nand U2961 (N_2961,N_2874,N_2807);
and U2962 (N_2962,N_2818,N_2808);
xnor U2963 (N_2963,N_2865,N_2883);
nor U2964 (N_2964,N_2851,N_2802);
and U2965 (N_2965,N_2899,N_2875);
and U2966 (N_2966,N_2817,N_2811);
nor U2967 (N_2967,N_2848,N_2863);
nor U2968 (N_2968,N_2847,N_2829);
nor U2969 (N_2969,N_2892,N_2851);
nand U2970 (N_2970,N_2841,N_2853);
and U2971 (N_2971,N_2823,N_2826);
nor U2972 (N_2972,N_2867,N_2852);
nand U2973 (N_2973,N_2846,N_2882);
and U2974 (N_2974,N_2895,N_2892);
nand U2975 (N_2975,N_2875,N_2845);
xor U2976 (N_2976,N_2884,N_2877);
or U2977 (N_2977,N_2844,N_2811);
or U2978 (N_2978,N_2870,N_2868);
and U2979 (N_2979,N_2816,N_2880);
or U2980 (N_2980,N_2818,N_2892);
xnor U2981 (N_2981,N_2853,N_2896);
and U2982 (N_2982,N_2870,N_2859);
nand U2983 (N_2983,N_2864,N_2885);
xnor U2984 (N_2984,N_2868,N_2885);
nand U2985 (N_2985,N_2862,N_2831);
nor U2986 (N_2986,N_2836,N_2843);
and U2987 (N_2987,N_2860,N_2811);
nor U2988 (N_2988,N_2814,N_2838);
and U2989 (N_2989,N_2806,N_2864);
xnor U2990 (N_2990,N_2870,N_2825);
and U2991 (N_2991,N_2866,N_2892);
xnor U2992 (N_2992,N_2854,N_2895);
nor U2993 (N_2993,N_2813,N_2860);
or U2994 (N_2994,N_2880,N_2847);
xor U2995 (N_2995,N_2882,N_2859);
or U2996 (N_2996,N_2863,N_2818);
or U2997 (N_2997,N_2847,N_2835);
nor U2998 (N_2998,N_2806,N_2824);
xor U2999 (N_2999,N_2842,N_2820);
nand UO_0 (O_0,N_2928,N_2906);
xor UO_1 (O_1,N_2997,N_2983);
nor UO_2 (O_2,N_2965,N_2923);
or UO_3 (O_3,N_2957,N_2987);
and UO_4 (O_4,N_2932,N_2918);
or UO_5 (O_5,N_2976,N_2930);
or UO_6 (O_6,N_2980,N_2922);
xor UO_7 (O_7,N_2908,N_2971);
xnor UO_8 (O_8,N_2989,N_2933);
and UO_9 (O_9,N_2979,N_2953);
nor UO_10 (O_10,N_2938,N_2984);
or UO_11 (O_11,N_2963,N_2916);
and UO_12 (O_12,N_2982,N_2919);
xor UO_13 (O_13,N_2939,N_2956);
nand UO_14 (O_14,N_2934,N_2941);
and UO_15 (O_15,N_2986,N_2921);
and UO_16 (O_16,N_2936,N_2926);
and UO_17 (O_17,N_2943,N_2972);
and UO_18 (O_18,N_2970,N_2998);
nor UO_19 (O_19,N_2977,N_2929);
and UO_20 (O_20,N_2966,N_2912);
and UO_21 (O_21,N_2905,N_2935);
or UO_22 (O_22,N_2924,N_2914);
nand UO_23 (O_23,N_2973,N_2990);
or UO_24 (O_24,N_2937,N_2958);
nand UO_25 (O_25,N_2964,N_2969);
nand UO_26 (O_26,N_2968,N_2951);
nand UO_27 (O_27,N_2945,N_2903);
nor UO_28 (O_28,N_2975,N_2901);
or UO_29 (O_29,N_2988,N_2995);
and UO_30 (O_30,N_2967,N_2978);
or UO_31 (O_31,N_2925,N_2915);
nand UO_32 (O_32,N_2999,N_2993);
nor UO_33 (O_33,N_2981,N_2952);
nor UO_34 (O_34,N_2902,N_2920);
or UO_35 (O_35,N_2927,N_2955);
and UO_36 (O_36,N_2910,N_2904);
or UO_37 (O_37,N_2909,N_2961);
xnor UO_38 (O_38,N_2948,N_2940);
and UO_39 (O_39,N_2911,N_2942);
nor UO_40 (O_40,N_2913,N_2931);
or UO_41 (O_41,N_2959,N_2917);
or UO_42 (O_42,N_2954,N_2949);
or UO_43 (O_43,N_2991,N_2992);
and UO_44 (O_44,N_2907,N_2946);
and UO_45 (O_45,N_2996,N_2960);
xnor UO_46 (O_46,N_2985,N_2947);
xnor UO_47 (O_47,N_2950,N_2994);
nor UO_48 (O_48,N_2974,N_2944);
nor UO_49 (O_49,N_2900,N_2962);
xor UO_50 (O_50,N_2996,N_2988);
nand UO_51 (O_51,N_2963,N_2950);
nor UO_52 (O_52,N_2936,N_2975);
nor UO_53 (O_53,N_2985,N_2952);
nor UO_54 (O_54,N_2969,N_2980);
nor UO_55 (O_55,N_2907,N_2959);
and UO_56 (O_56,N_2938,N_2961);
or UO_57 (O_57,N_2934,N_2931);
nor UO_58 (O_58,N_2970,N_2974);
nor UO_59 (O_59,N_2953,N_2909);
xor UO_60 (O_60,N_2971,N_2909);
or UO_61 (O_61,N_2917,N_2913);
or UO_62 (O_62,N_2939,N_2923);
and UO_63 (O_63,N_2924,N_2940);
xnor UO_64 (O_64,N_2916,N_2941);
nor UO_65 (O_65,N_2922,N_2962);
nor UO_66 (O_66,N_2945,N_2926);
nand UO_67 (O_67,N_2998,N_2969);
or UO_68 (O_68,N_2903,N_2932);
nand UO_69 (O_69,N_2987,N_2983);
and UO_70 (O_70,N_2900,N_2983);
nand UO_71 (O_71,N_2923,N_2992);
or UO_72 (O_72,N_2949,N_2929);
or UO_73 (O_73,N_2994,N_2982);
nor UO_74 (O_74,N_2933,N_2917);
and UO_75 (O_75,N_2961,N_2900);
nand UO_76 (O_76,N_2989,N_2942);
nor UO_77 (O_77,N_2972,N_2975);
nand UO_78 (O_78,N_2953,N_2958);
xnor UO_79 (O_79,N_2998,N_2989);
xor UO_80 (O_80,N_2932,N_2925);
and UO_81 (O_81,N_2956,N_2908);
or UO_82 (O_82,N_2979,N_2966);
nor UO_83 (O_83,N_2975,N_2957);
or UO_84 (O_84,N_2938,N_2902);
nand UO_85 (O_85,N_2953,N_2932);
or UO_86 (O_86,N_2901,N_2969);
and UO_87 (O_87,N_2994,N_2976);
or UO_88 (O_88,N_2928,N_2957);
and UO_89 (O_89,N_2916,N_2902);
xor UO_90 (O_90,N_2978,N_2988);
nand UO_91 (O_91,N_2986,N_2925);
nand UO_92 (O_92,N_2934,N_2965);
and UO_93 (O_93,N_2989,N_2977);
nor UO_94 (O_94,N_2902,N_2926);
xor UO_95 (O_95,N_2937,N_2910);
and UO_96 (O_96,N_2966,N_2961);
or UO_97 (O_97,N_2904,N_2968);
nor UO_98 (O_98,N_2912,N_2970);
and UO_99 (O_99,N_2937,N_2900);
nor UO_100 (O_100,N_2915,N_2983);
nand UO_101 (O_101,N_2942,N_2984);
and UO_102 (O_102,N_2986,N_2991);
nor UO_103 (O_103,N_2961,N_2955);
or UO_104 (O_104,N_2908,N_2929);
and UO_105 (O_105,N_2907,N_2999);
and UO_106 (O_106,N_2901,N_2974);
nor UO_107 (O_107,N_2922,N_2967);
or UO_108 (O_108,N_2976,N_2949);
nand UO_109 (O_109,N_2990,N_2938);
or UO_110 (O_110,N_2904,N_2981);
xor UO_111 (O_111,N_2942,N_2949);
nand UO_112 (O_112,N_2970,N_2937);
and UO_113 (O_113,N_2912,N_2913);
xnor UO_114 (O_114,N_2926,N_2958);
xnor UO_115 (O_115,N_2970,N_2972);
and UO_116 (O_116,N_2929,N_2913);
and UO_117 (O_117,N_2914,N_2941);
and UO_118 (O_118,N_2990,N_2915);
nor UO_119 (O_119,N_2940,N_2985);
xnor UO_120 (O_120,N_2988,N_2941);
and UO_121 (O_121,N_2938,N_2933);
xnor UO_122 (O_122,N_2902,N_2974);
nor UO_123 (O_123,N_2986,N_2984);
and UO_124 (O_124,N_2953,N_2936);
nor UO_125 (O_125,N_2910,N_2993);
nand UO_126 (O_126,N_2965,N_2993);
or UO_127 (O_127,N_2900,N_2973);
and UO_128 (O_128,N_2950,N_2969);
nor UO_129 (O_129,N_2908,N_2919);
nor UO_130 (O_130,N_2925,N_2916);
nand UO_131 (O_131,N_2977,N_2955);
xnor UO_132 (O_132,N_2951,N_2981);
nand UO_133 (O_133,N_2951,N_2996);
or UO_134 (O_134,N_2958,N_2991);
xor UO_135 (O_135,N_2970,N_2949);
xnor UO_136 (O_136,N_2959,N_2964);
or UO_137 (O_137,N_2905,N_2995);
nor UO_138 (O_138,N_2922,N_2954);
or UO_139 (O_139,N_2903,N_2960);
and UO_140 (O_140,N_2910,N_2992);
nand UO_141 (O_141,N_2993,N_2997);
nand UO_142 (O_142,N_2989,N_2904);
and UO_143 (O_143,N_2950,N_2919);
or UO_144 (O_144,N_2919,N_2926);
nor UO_145 (O_145,N_2940,N_2910);
nand UO_146 (O_146,N_2965,N_2937);
or UO_147 (O_147,N_2916,N_2906);
and UO_148 (O_148,N_2900,N_2950);
xor UO_149 (O_149,N_2910,N_2999);
and UO_150 (O_150,N_2902,N_2990);
or UO_151 (O_151,N_2927,N_2942);
or UO_152 (O_152,N_2950,N_2997);
or UO_153 (O_153,N_2989,N_2915);
xor UO_154 (O_154,N_2934,N_2936);
and UO_155 (O_155,N_2941,N_2949);
xor UO_156 (O_156,N_2969,N_2970);
and UO_157 (O_157,N_2904,N_2934);
nand UO_158 (O_158,N_2921,N_2984);
or UO_159 (O_159,N_2995,N_2909);
nor UO_160 (O_160,N_2906,N_2945);
or UO_161 (O_161,N_2918,N_2984);
nand UO_162 (O_162,N_2903,N_2938);
and UO_163 (O_163,N_2913,N_2926);
or UO_164 (O_164,N_2902,N_2951);
and UO_165 (O_165,N_2990,N_2925);
xnor UO_166 (O_166,N_2900,N_2928);
and UO_167 (O_167,N_2977,N_2992);
nand UO_168 (O_168,N_2994,N_2964);
nand UO_169 (O_169,N_2985,N_2968);
xor UO_170 (O_170,N_2989,N_2932);
nand UO_171 (O_171,N_2978,N_2952);
xor UO_172 (O_172,N_2940,N_2938);
or UO_173 (O_173,N_2913,N_2910);
nand UO_174 (O_174,N_2988,N_2900);
nor UO_175 (O_175,N_2935,N_2921);
xor UO_176 (O_176,N_2932,N_2958);
and UO_177 (O_177,N_2917,N_2927);
nand UO_178 (O_178,N_2947,N_2973);
nor UO_179 (O_179,N_2947,N_2968);
and UO_180 (O_180,N_2915,N_2972);
nor UO_181 (O_181,N_2919,N_2976);
xnor UO_182 (O_182,N_2901,N_2934);
and UO_183 (O_183,N_2943,N_2944);
nand UO_184 (O_184,N_2990,N_2911);
and UO_185 (O_185,N_2911,N_2985);
or UO_186 (O_186,N_2930,N_2998);
or UO_187 (O_187,N_2977,N_2901);
nand UO_188 (O_188,N_2961,N_2957);
xor UO_189 (O_189,N_2932,N_2999);
nand UO_190 (O_190,N_2935,N_2999);
and UO_191 (O_191,N_2935,N_2994);
nor UO_192 (O_192,N_2967,N_2912);
xor UO_193 (O_193,N_2917,N_2944);
xnor UO_194 (O_194,N_2985,N_2980);
or UO_195 (O_195,N_2966,N_2973);
or UO_196 (O_196,N_2930,N_2980);
nand UO_197 (O_197,N_2990,N_2986);
nand UO_198 (O_198,N_2924,N_2983);
or UO_199 (O_199,N_2960,N_2953);
nand UO_200 (O_200,N_2957,N_2930);
nand UO_201 (O_201,N_2995,N_2947);
and UO_202 (O_202,N_2977,N_2922);
xnor UO_203 (O_203,N_2951,N_2952);
nand UO_204 (O_204,N_2903,N_2955);
nand UO_205 (O_205,N_2998,N_2967);
and UO_206 (O_206,N_2960,N_2949);
nand UO_207 (O_207,N_2970,N_2906);
and UO_208 (O_208,N_2956,N_2918);
nand UO_209 (O_209,N_2985,N_2993);
nor UO_210 (O_210,N_2961,N_2981);
and UO_211 (O_211,N_2975,N_2909);
nor UO_212 (O_212,N_2984,N_2991);
and UO_213 (O_213,N_2952,N_2942);
and UO_214 (O_214,N_2923,N_2947);
nand UO_215 (O_215,N_2902,N_2936);
nor UO_216 (O_216,N_2903,N_2984);
xnor UO_217 (O_217,N_2968,N_2913);
nand UO_218 (O_218,N_2990,N_2952);
nand UO_219 (O_219,N_2983,N_2904);
nor UO_220 (O_220,N_2906,N_2905);
or UO_221 (O_221,N_2997,N_2973);
nor UO_222 (O_222,N_2923,N_2977);
xnor UO_223 (O_223,N_2976,N_2900);
xor UO_224 (O_224,N_2935,N_2983);
nor UO_225 (O_225,N_2928,N_2956);
nand UO_226 (O_226,N_2977,N_2967);
and UO_227 (O_227,N_2961,N_2945);
nor UO_228 (O_228,N_2998,N_2925);
xnor UO_229 (O_229,N_2937,N_2901);
xor UO_230 (O_230,N_2947,N_2903);
nand UO_231 (O_231,N_2932,N_2997);
xnor UO_232 (O_232,N_2995,N_2972);
or UO_233 (O_233,N_2963,N_2989);
and UO_234 (O_234,N_2995,N_2991);
nor UO_235 (O_235,N_2969,N_2999);
nor UO_236 (O_236,N_2903,N_2998);
xnor UO_237 (O_237,N_2984,N_2951);
xnor UO_238 (O_238,N_2900,N_2929);
nand UO_239 (O_239,N_2924,N_2956);
xnor UO_240 (O_240,N_2987,N_2976);
xnor UO_241 (O_241,N_2998,N_2932);
nor UO_242 (O_242,N_2922,N_2976);
nand UO_243 (O_243,N_2949,N_2922);
and UO_244 (O_244,N_2981,N_2960);
nor UO_245 (O_245,N_2914,N_2986);
xor UO_246 (O_246,N_2934,N_2970);
and UO_247 (O_247,N_2913,N_2906);
nand UO_248 (O_248,N_2960,N_2928);
or UO_249 (O_249,N_2906,N_2949);
or UO_250 (O_250,N_2958,N_2979);
and UO_251 (O_251,N_2987,N_2991);
and UO_252 (O_252,N_2916,N_2961);
and UO_253 (O_253,N_2932,N_2985);
or UO_254 (O_254,N_2996,N_2989);
or UO_255 (O_255,N_2946,N_2986);
or UO_256 (O_256,N_2939,N_2949);
xnor UO_257 (O_257,N_2919,N_2910);
xnor UO_258 (O_258,N_2987,N_2980);
nor UO_259 (O_259,N_2958,N_2957);
or UO_260 (O_260,N_2931,N_2922);
nand UO_261 (O_261,N_2965,N_2974);
or UO_262 (O_262,N_2916,N_2940);
xor UO_263 (O_263,N_2942,N_2937);
nand UO_264 (O_264,N_2969,N_2954);
nor UO_265 (O_265,N_2905,N_2959);
nor UO_266 (O_266,N_2968,N_2920);
xor UO_267 (O_267,N_2979,N_2903);
xor UO_268 (O_268,N_2905,N_2976);
and UO_269 (O_269,N_2939,N_2950);
xor UO_270 (O_270,N_2951,N_2959);
nor UO_271 (O_271,N_2941,N_2907);
and UO_272 (O_272,N_2911,N_2969);
nor UO_273 (O_273,N_2909,N_2960);
xor UO_274 (O_274,N_2909,N_2983);
or UO_275 (O_275,N_2933,N_2982);
nand UO_276 (O_276,N_2953,N_2910);
nand UO_277 (O_277,N_2967,N_2973);
nand UO_278 (O_278,N_2917,N_2963);
nor UO_279 (O_279,N_2904,N_2995);
nor UO_280 (O_280,N_2901,N_2962);
nor UO_281 (O_281,N_2944,N_2937);
or UO_282 (O_282,N_2931,N_2954);
nor UO_283 (O_283,N_2983,N_2907);
nor UO_284 (O_284,N_2939,N_2999);
nor UO_285 (O_285,N_2902,N_2967);
xor UO_286 (O_286,N_2901,N_2902);
or UO_287 (O_287,N_2978,N_2979);
xor UO_288 (O_288,N_2994,N_2958);
xnor UO_289 (O_289,N_2950,N_2915);
nand UO_290 (O_290,N_2935,N_2977);
xnor UO_291 (O_291,N_2913,N_2963);
and UO_292 (O_292,N_2919,N_2989);
and UO_293 (O_293,N_2936,N_2994);
xnor UO_294 (O_294,N_2943,N_2954);
nand UO_295 (O_295,N_2998,N_2927);
and UO_296 (O_296,N_2949,N_2908);
nor UO_297 (O_297,N_2929,N_2999);
or UO_298 (O_298,N_2977,N_2933);
and UO_299 (O_299,N_2975,N_2934);
nor UO_300 (O_300,N_2904,N_2947);
and UO_301 (O_301,N_2943,N_2970);
xor UO_302 (O_302,N_2935,N_2934);
xor UO_303 (O_303,N_2909,N_2901);
or UO_304 (O_304,N_2990,N_2917);
and UO_305 (O_305,N_2931,N_2964);
nor UO_306 (O_306,N_2936,N_2965);
and UO_307 (O_307,N_2956,N_2969);
and UO_308 (O_308,N_2997,N_2922);
or UO_309 (O_309,N_2949,N_2930);
nor UO_310 (O_310,N_2981,N_2956);
or UO_311 (O_311,N_2907,N_2989);
nand UO_312 (O_312,N_2914,N_2933);
and UO_313 (O_313,N_2964,N_2903);
nor UO_314 (O_314,N_2954,N_2952);
nor UO_315 (O_315,N_2974,N_2913);
and UO_316 (O_316,N_2907,N_2948);
xor UO_317 (O_317,N_2993,N_2944);
nand UO_318 (O_318,N_2958,N_2934);
xor UO_319 (O_319,N_2983,N_2921);
xor UO_320 (O_320,N_2907,N_2908);
nor UO_321 (O_321,N_2906,N_2998);
or UO_322 (O_322,N_2996,N_2965);
nand UO_323 (O_323,N_2938,N_2954);
and UO_324 (O_324,N_2949,N_2958);
and UO_325 (O_325,N_2919,N_2954);
and UO_326 (O_326,N_2924,N_2988);
xor UO_327 (O_327,N_2949,N_2927);
xnor UO_328 (O_328,N_2943,N_2923);
xor UO_329 (O_329,N_2904,N_2972);
or UO_330 (O_330,N_2994,N_2925);
or UO_331 (O_331,N_2989,N_2918);
or UO_332 (O_332,N_2976,N_2907);
or UO_333 (O_333,N_2998,N_2972);
nand UO_334 (O_334,N_2924,N_2975);
nor UO_335 (O_335,N_2918,N_2952);
xor UO_336 (O_336,N_2940,N_2956);
nor UO_337 (O_337,N_2992,N_2960);
nor UO_338 (O_338,N_2961,N_2985);
nand UO_339 (O_339,N_2971,N_2973);
xnor UO_340 (O_340,N_2979,N_2977);
or UO_341 (O_341,N_2961,N_2910);
xor UO_342 (O_342,N_2986,N_2902);
or UO_343 (O_343,N_2947,N_2943);
nand UO_344 (O_344,N_2976,N_2901);
nand UO_345 (O_345,N_2926,N_2973);
xnor UO_346 (O_346,N_2926,N_2994);
xor UO_347 (O_347,N_2918,N_2991);
nand UO_348 (O_348,N_2976,N_2913);
and UO_349 (O_349,N_2988,N_2904);
xnor UO_350 (O_350,N_2927,N_2984);
nor UO_351 (O_351,N_2907,N_2936);
or UO_352 (O_352,N_2929,N_2958);
or UO_353 (O_353,N_2994,N_2913);
and UO_354 (O_354,N_2984,N_2902);
xor UO_355 (O_355,N_2949,N_2963);
nor UO_356 (O_356,N_2981,N_2908);
nand UO_357 (O_357,N_2985,N_2962);
or UO_358 (O_358,N_2985,N_2939);
and UO_359 (O_359,N_2924,N_2923);
xor UO_360 (O_360,N_2944,N_2992);
nor UO_361 (O_361,N_2966,N_2964);
nand UO_362 (O_362,N_2966,N_2929);
nor UO_363 (O_363,N_2974,N_2973);
nand UO_364 (O_364,N_2944,N_2933);
nand UO_365 (O_365,N_2913,N_2993);
or UO_366 (O_366,N_2922,N_2939);
and UO_367 (O_367,N_2928,N_2929);
or UO_368 (O_368,N_2972,N_2950);
nor UO_369 (O_369,N_2928,N_2905);
nor UO_370 (O_370,N_2940,N_2926);
xor UO_371 (O_371,N_2915,N_2949);
and UO_372 (O_372,N_2934,N_2940);
nand UO_373 (O_373,N_2919,N_2968);
nor UO_374 (O_374,N_2912,N_2962);
and UO_375 (O_375,N_2924,N_2907);
or UO_376 (O_376,N_2970,N_2913);
nor UO_377 (O_377,N_2970,N_2923);
nor UO_378 (O_378,N_2929,N_2985);
and UO_379 (O_379,N_2937,N_2904);
xor UO_380 (O_380,N_2933,N_2946);
xnor UO_381 (O_381,N_2997,N_2924);
nand UO_382 (O_382,N_2954,N_2964);
and UO_383 (O_383,N_2941,N_2982);
nor UO_384 (O_384,N_2968,N_2989);
nand UO_385 (O_385,N_2964,N_2943);
or UO_386 (O_386,N_2995,N_2989);
and UO_387 (O_387,N_2920,N_2912);
nand UO_388 (O_388,N_2936,N_2931);
xnor UO_389 (O_389,N_2952,N_2925);
or UO_390 (O_390,N_2942,N_2943);
or UO_391 (O_391,N_2934,N_2933);
and UO_392 (O_392,N_2984,N_2900);
nand UO_393 (O_393,N_2936,N_2972);
and UO_394 (O_394,N_2937,N_2960);
nor UO_395 (O_395,N_2986,N_2907);
xnor UO_396 (O_396,N_2962,N_2967);
or UO_397 (O_397,N_2964,N_2948);
or UO_398 (O_398,N_2992,N_2997);
or UO_399 (O_399,N_2946,N_2989);
nor UO_400 (O_400,N_2919,N_2963);
nor UO_401 (O_401,N_2942,N_2996);
or UO_402 (O_402,N_2923,N_2925);
and UO_403 (O_403,N_2998,N_2949);
nand UO_404 (O_404,N_2971,N_2914);
or UO_405 (O_405,N_2934,N_2980);
or UO_406 (O_406,N_2943,N_2936);
xnor UO_407 (O_407,N_2910,N_2972);
and UO_408 (O_408,N_2965,N_2911);
xnor UO_409 (O_409,N_2938,N_2962);
xnor UO_410 (O_410,N_2942,N_2981);
xnor UO_411 (O_411,N_2942,N_2978);
nand UO_412 (O_412,N_2969,N_2960);
and UO_413 (O_413,N_2915,N_2923);
or UO_414 (O_414,N_2933,N_2954);
nor UO_415 (O_415,N_2974,N_2952);
xor UO_416 (O_416,N_2975,N_2945);
nand UO_417 (O_417,N_2937,N_2936);
or UO_418 (O_418,N_2953,N_2952);
nand UO_419 (O_419,N_2963,N_2981);
and UO_420 (O_420,N_2933,N_2976);
nand UO_421 (O_421,N_2974,N_2908);
or UO_422 (O_422,N_2927,N_2946);
or UO_423 (O_423,N_2907,N_2915);
xor UO_424 (O_424,N_2946,N_2929);
nand UO_425 (O_425,N_2936,N_2991);
and UO_426 (O_426,N_2952,N_2914);
and UO_427 (O_427,N_2908,N_2937);
nor UO_428 (O_428,N_2941,N_2997);
nand UO_429 (O_429,N_2953,N_2988);
and UO_430 (O_430,N_2952,N_2902);
xnor UO_431 (O_431,N_2910,N_2976);
and UO_432 (O_432,N_2986,N_2973);
or UO_433 (O_433,N_2926,N_2993);
or UO_434 (O_434,N_2970,N_2959);
or UO_435 (O_435,N_2957,N_2919);
and UO_436 (O_436,N_2984,N_2944);
nand UO_437 (O_437,N_2948,N_2922);
or UO_438 (O_438,N_2994,N_2966);
nand UO_439 (O_439,N_2980,N_2991);
or UO_440 (O_440,N_2976,N_2906);
and UO_441 (O_441,N_2949,N_2905);
nand UO_442 (O_442,N_2998,N_2933);
or UO_443 (O_443,N_2912,N_2911);
and UO_444 (O_444,N_2940,N_2997);
nor UO_445 (O_445,N_2974,N_2916);
nor UO_446 (O_446,N_2912,N_2934);
nand UO_447 (O_447,N_2905,N_2923);
nor UO_448 (O_448,N_2960,N_2930);
nand UO_449 (O_449,N_2967,N_2959);
nand UO_450 (O_450,N_2967,N_2939);
and UO_451 (O_451,N_2955,N_2967);
nand UO_452 (O_452,N_2950,N_2968);
or UO_453 (O_453,N_2910,N_2951);
nor UO_454 (O_454,N_2933,N_2903);
and UO_455 (O_455,N_2913,N_2916);
nor UO_456 (O_456,N_2942,N_2972);
or UO_457 (O_457,N_2905,N_2903);
and UO_458 (O_458,N_2909,N_2926);
and UO_459 (O_459,N_2915,N_2940);
or UO_460 (O_460,N_2942,N_2906);
xnor UO_461 (O_461,N_2999,N_2918);
nor UO_462 (O_462,N_2916,N_2955);
or UO_463 (O_463,N_2972,N_2903);
xor UO_464 (O_464,N_2974,N_2958);
nand UO_465 (O_465,N_2917,N_2979);
xor UO_466 (O_466,N_2968,N_2990);
nor UO_467 (O_467,N_2998,N_2986);
nor UO_468 (O_468,N_2933,N_2937);
nor UO_469 (O_469,N_2941,N_2985);
nor UO_470 (O_470,N_2952,N_2923);
or UO_471 (O_471,N_2988,N_2928);
or UO_472 (O_472,N_2945,N_2947);
and UO_473 (O_473,N_2908,N_2906);
and UO_474 (O_474,N_2903,N_2925);
or UO_475 (O_475,N_2956,N_2959);
and UO_476 (O_476,N_2939,N_2977);
nand UO_477 (O_477,N_2992,N_2951);
xnor UO_478 (O_478,N_2939,N_2918);
nor UO_479 (O_479,N_2939,N_2969);
and UO_480 (O_480,N_2957,N_2934);
nor UO_481 (O_481,N_2922,N_2990);
and UO_482 (O_482,N_2914,N_2991);
nor UO_483 (O_483,N_2945,N_2916);
or UO_484 (O_484,N_2905,N_2900);
and UO_485 (O_485,N_2909,N_2987);
xor UO_486 (O_486,N_2930,N_2909);
xnor UO_487 (O_487,N_2925,N_2933);
and UO_488 (O_488,N_2959,N_2975);
and UO_489 (O_489,N_2923,N_2919);
xor UO_490 (O_490,N_2934,N_2902);
xnor UO_491 (O_491,N_2958,N_2970);
and UO_492 (O_492,N_2961,N_2942);
xnor UO_493 (O_493,N_2945,N_2954);
or UO_494 (O_494,N_2963,N_2903);
or UO_495 (O_495,N_2987,N_2973);
nand UO_496 (O_496,N_2962,N_2928);
nand UO_497 (O_497,N_2996,N_2912);
nor UO_498 (O_498,N_2942,N_2997);
xnor UO_499 (O_499,N_2972,N_2902);
endmodule