module basic_3000_30000_3500_60_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_2789,In_895);
and U1 (N_1,In_2209,In_73);
or U2 (N_2,In_2131,In_934);
or U3 (N_3,In_1572,In_56);
xor U4 (N_4,In_1749,In_373);
or U5 (N_5,In_118,In_1427);
or U6 (N_6,In_1971,In_211);
and U7 (N_7,In_628,In_2323);
xor U8 (N_8,In_748,In_497);
and U9 (N_9,In_1881,In_1762);
nand U10 (N_10,In_653,In_1428);
xor U11 (N_11,In_2260,In_760);
or U12 (N_12,In_2073,In_2654);
nor U13 (N_13,In_161,In_1928);
or U14 (N_14,In_1310,In_1676);
nand U15 (N_15,In_1872,In_2103);
xnor U16 (N_16,In_1908,In_1142);
nand U17 (N_17,In_1441,In_1827);
xnor U18 (N_18,In_2432,In_1770);
nand U19 (N_19,In_2025,In_1537);
xor U20 (N_20,In_1470,In_474);
or U21 (N_21,In_657,In_1498);
nor U22 (N_22,In_709,In_806);
or U23 (N_23,In_517,In_326);
and U24 (N_24,In_1471,In_213);
or U25 (N_25,In_402,In_2520);
nand U26 (N_26,In_2058,In_2094);
nor U27 (N_27,In_2879,In_2697);
and U28 (N_28,In_1829,In_1461);
or U29 (N_29,In_1303,In_2017);
and U30 (N_30,In_2881,In_2882);
nand U31 (N_31,In_1245,In_1631);
nor U32 (N_32,In_1816,In_2134);
nand U33 (N_33,In_570,In_1033);
nor U34 (N_34,In_1091,In_611);
or U35 (N_35,In_1269,In_691);
or U36 (N_36,In_218,In_2326);
xor U37 (N_37,In_410,In_2913);
nor U38 (N_38,In_1440,In_1768);
or U39 (N_39,In_2829,In_114);
and U40 (N_40,In_879,In_2346);
and U41 (N_41,In_2428,In_1579);
xnor U42 (N_42,In_222,In_65);
nand U43 (N_43,In_2948,In_1696);
nor U44 (N_44,In_2767,In_324);
nor U45 (N_45,In_2386,In_661);
and U46 (N_46,In_1165,In_1358);
xnor U47 (N_47,In_273,In_1279);
and U48 (N_48,In_1840,In_2825);
or U49 (N_49,In_589,In_2987);
nand U50 (N_50,In_1945,In_2537);
xor U51 (N_51,In_2007,In_972);
or U52 (N_52,In_2979,In_2037);
nand U53 (N_53,In_292,In_2999);
xnor U54 (N_54,In_2641,In_966);
xor U55 (N_55,In_1502,In_365);
nor U56 (N_56,In_244,In_254);
and U57 (N_57,In_988,In_2120);
or U58 (N_58,In_2500,In_742);
nor U59 (N_59,In_1174,In_1511);
nor U60 (N_60,In_1521,In_2168);
nor U61 (N_61,In_1843,In_2454);
nor U62 (N_62,In_142,In_307);
and U63 (N_63,In_2099,In_2587);
and U64 (N_64,In_2779,In_2297);
nand U65 (N_65,In_1841,In_1071);
xor U66 (N_66,In_2033,In_524);
or U67 (N_67,In_2307,In_1981);
xnor U68 (N_68,In_1281,In_2807);
nor U69 (N_69,In_2281,In_235);
and U70 (N_70,In_1691,In_917);
or U71 (N_71,In_1481,In_430);
nor U72 (N_72,In_996,In_2092);
xnor U73 (N_73,In_1853,In_2889);
nor U74 (N_74,In_1718,In_2242);
nand U75 (N_75,In_2304,In_915);
xor U76 (N_76,In_2378,In_2546);
xnor U77 (N_77,In_868,In_2236);
nand U78 (N_78,In_801,In_2111);
nand U79 (N_79,In_1237,In_2851);
xnor U80 (N_80,In_1658,In_1675);
and U81 (N_81,In_2202,In_2868);
xnor U82 (N_82,In_1261,In_2536);
xor U83 (N_83,In_2241,In_156);
and U84 (N_84,In_420,In_382);
or U85 (N_85,In_2726,In_1622);
nand U86 (N_86,In_2569,In_287);
xnor U87 (N_87,In_2350,In_2270);
and U88 (N_88,In_1247,In_1611);
or U89 (N_89,In_484,In_1367);
xnor U90 (N_90,In_592,In_2353);
xor U91 (N_91,In_1680,In_1545);
or U92 (N_92,In_622,In_2718);
or U93 (N_93,In_1251,In_660);
nand U94 (N_94,In_2351,In_2405);
nor U95 (N_95,In_1201,In_638);
nand U96 (N_96,In_2959,In_2574);
nand U97 (N_97,In_1751,In_1713);
and U98 (N_98,In_1534,In_1554);
and U99 (N_99,In_625,In_1487);
nor U100 (N_100,In_931,In_648);
nand U101 (N_101,In_2674,In_2395);
and U102 (N_102,In_1295,In_250);
nor U103 (N_103,In_1815,In_2700);
nor U104 (N_104,In_2832,In_1746);
or U105 (N_105,In_2330,In_62);
nor U106 (N_106,In_2356,In_473);
xor U107 (N_107,In_520,In_659);
nor U108 (N_108,In_198,In_332);
xor U109 (N_109,In_500,In_199);
nor U110 (N_110,In_1342,In_1535);
xor U111 (N_111,In_761,In_2671);
xnor U112 (N_112,In_94,In_1507);
xor U113 (N_113,In_1596,In_792);
xnor U114 (N_114,In_275,In_2963);
xnor U115 (N_115,In_2176,In_2684);
and U116 (N_116,In_2827,In_1);
or U117 (N_117,In_2429,In_1810);
and U118 (N_118,In_391,In_2178);
nand U119 (N_119,In_1469,In_1108);
nand U120 (N_120,In_2720,In_2298);
or U121 (N_121,In_428,In_1285);
or U122 (N_122,In_1066,In_745);
and U123 (N_123,In_1255,In_131);
or U124 (N_124,In_2918,In_906);
nand U125 (N_125,In_2699,In_579);
xnor U126 (N_126,In_1500,In_1377);
xnor U127 (N_127,In_945,In_1651);
and U128 (N_128,In_2044,In_2690);
and U129 (N_129,In_2483,In_1681);
nor U130 (N_130,In_2045,In_2565);
xnor U131 (N_131,In_833,In_1114);
xnor U132 (N_132,In_2371,In_1378);
and U133 (N_133,In_1542,In_2524);
nand U134 (N_134,In_357,In_680);
xor U135 (N_135,In_1664,In_1182);
nand U136 (N_136,In_81,In_1733);
nor U137 (N_137,In_2530,In_303);
and U138 (N_138,In_195,In_468);
or U139 (N_139,In_781,In_900);
or U140 (N_140,In_259,In_165);
or U141 (N_141,In_1570,In_1308);
nor U142 (N_142,In_1380,In_604);
nand U143 (N_143,In_2581,In_1972);
and U144 (N_144,In_2138,In_2757);
xnor U145 (N_145,In_1786,In_2054);
xnor U146 (N_146,In_2375,In_70);
nor U147 (N_147,In_2600,In_567);
nor U148 (N_148,In_2908,In_2820);
nor U149 (N_149,In_898,In_358);
nor U150 (N_150,In_92,In_1757);
and U151 (N_151,In_2397,In_2137);
xor U152 (N_152,In_1646,In_1501);
or U153 (N_153,In_1429,In_2919);
nand U154 (N_154,In_1687,In_2655);
or U155 (N_155,In_172,In_706);
xor U156 (N_156,In_713,In_2156);
nand U157 (N_157,In_393,In_2701);
and U158 (N_158,In_378,In_1458);
nor U159 (N_159,In_2442,In_2257);
nand U160 (N_160,In_2437,In_1519);
nor U161 (N_161,In_1421,In_2883);
nand U162 (N_162,In_1300,In_1288);
nor U163 (N_163,In_1929,In_1027);
or U164 (N_164,In_1386,In_459);
xnor U165 (N_165,In_2512,In_1573);
nand U166 (N_166,In_557,In_1640);
and U167 (N_167,In_107,In_89);
nor U168 (N_168,In_1890,In_2614);
or U169 (N_169,In_1650,In_846);
xnor U170 (N_170,In_400,In_2036);
and U171 (N_171,In_2592,In_2104);
and U172 (N_172,In_1065,In_636);
xnor U173 (N_173,In_2848,In_1606);
xor U174 (N_174,In_369,In_1709);
nor U175 (N_175,In_2423,In_479);
nand U176 (N_176,In_1963,In_509);
xor U177 (N_177,In_2184,In_2552);
nor U178 (N_178,In_729,In_1638);
nor U179 (N_179,In_2462,In_1067);
nor U180 (N_180,In_1807,In_362);
xor U181 (N_181,In_2471,In_187);
nand U182 (N_182,In_605,In_2164);
nor U183 (N_183,In_2172,In_901);
or U184 (N_184,In_1144,In_2840);
or U185 (N_185,In_80,In_2802);
xnor U186 (N_186,In_1394,In_734);
xor U187 (N_187,In_2446,In_2831);
xnor U188 (N_188,In_2694,In_1665);
nand U189 (N_189,In_201,In_1097);
or U190 (N_190,In_2933,In_776);
nor U191 (N_191,In_2905,In_1878);
nand U192 (N_192,In_1912,In_285);
and U193 (N_193,In_1524,In_1900);
and U194 (N_194,In_1785,In_586);
nand U195 (N_195,In_2285,In_1047);
nand U196 (N_196,In_2998,In_54);
nand U197 (N_197,In_746,In_805);
nor U198 (N_198,In_682,In_85);
nor U199 (N_199,In_2775,In_1924);
nor U200 (N_200,In_2736,In_2125);
or U201 (N_201,In_2810,In_2459);
and U202 (N_202,In_329,In_328);
nor U203 (N_203,In_2336,In_1381);
nand U204 (N_204,In_2452,In_1660);
xor U205 (N_205,In_2362,In_2381);
nand U206 (N_206,In_2162,In_2254);
nor U207 (N_207,In_1761,In_225);
xor U208 (N_208,In_2766,In_2838);
or U209 (N_209,In_1043,In_1857);
nor U210 (N_210,In_907,In_1617);
nand U211 (N_211,In_2890,In_2739);
or U212 (N_212,In_535,In_614);
nor U213 (N_213,In_878,In_488);
nor U214 (N_214,In_1172,In_1045);
and U215 (N_215,In_2174,In_1203);
and U216 (N_216,In_1565,In_920);
or U217 (N_217,In_2447,In_2481);
or U218 (N_218,In_866,In_2426);
xor U219 (N_219,In_1880,In_1339);
nor U220 (N_220,In_79,In_2361);
and U221 (N_221,In_2862,In_1276);
nor U222 (N_222,In_1003,In_2598);
xor U223 (N_223,In_1164,In_1867);
nor U224 (N_224,In_2294,In_1149);
nand U225 (N_225,In_652,In_404);
xor U226 (N_226,In_1546,In_597);
nand U227 (N_227,In_2216,In_2567);
and U228 (N_228,In_756,In_1992);
nor U229 (N_229,In_1959,In_1375);
xor U230 (N_230,In_301,In_1384);
nand U231 (N_231,In_2124,In_457);
and U232 (N_232,In_1459,In_825);
or U233 (N_233,In_82,In_1183);
or U234 (N_234,In_1609,In_2163);
or U235 (N_235,In_1050,In_316);
nor U236 (N_236,In_2101,In_1153);
nor U237 (N_237,In_1395,In_1913);
nand U238 (N_238,In_2510,In_1802);
xor U239 (N_239,In_747,In_645);
and U240 (N_240,In_2155,In_1350);
nand U241 (N_241,In_72,In_1316);
xor U242 (N_242,In_2728,In_1781);
nor U243 (N_243,In_2219,In_574);
and U244 (N_244,In_1443,In_1671);
and U245 (N_245,In_1086,In_874);
nand U246 (N_246,In_1294,In_101);
and U247 (N_247,In_1776,In_753);
xnor U248 (N_248,In_1520,In_505);
or U249 (N_249,In_1348,In_2899);
xor U250 (N_250,In_811,In_1355);
nand U251 (N_251,In_647,In_774);
and U252 (N_252,In_2066,In_1766);
and U253 (N_253,In_2801,In_1845);
nand U254 (N_254,In_1042,In_455);
and U255 (N_255,In_556,In_1111);
xnor U256 (N_256,In_1764,In_280);
or U257 (N_257,In_2649,In_704);
and U258 (N_258,In_317,In_1817);
and U259 (N_259,In_2860,In_1644);
nand U260 (N_260,In_2836,In_1057);
and U261 (N_261,In_2263,In_1922);
xor U262 (N_262,In_2553,In_1119);
nand U263 (N_263,In_1264,In_1448);
nor U264 (N_264,In_1527,In_764);
and U265 (N_265,In_193,In_1997);
or U266 (N_266,In_736,In_1844);
and U267 (N_267,In_651,In_1645);
nand U268 (N_268,In_2746,In_260);
nor U269 (N_269,In_1287,In_434);
nand U270 (N_270,In_2144,In_529);
and U271 (N_271,In_2608,In_2891);
nor U272 (N_272,In_309,In_339);
nand U273 (N_273,In_1087,In_2482);
or U274 (N_274,In_421,In_1438);
xor U275 (N_275,In_1224,In_1915);
nor U276 (N_276,In_2605,In_2011);
nand U277 (N_277,In_1726,In_663);
or U278 (N_278,In_1455,In_914);
xnor U279 (N_279,In_2075,In_471);
xor U280 (N_280,In_1508,In_2215);
and U281 (N_281,In_1998,In_705);
or U282 (N_282,In_2169,In_646);
nor U283 (N_283,In_1836,In_1098);
xor U284 (N_284,In_2522,In_150);
or U285 (N_285,In_88,In_1124);
nor U286 (N_286,In_284,In_2339);
and U287 (N_287,In_1413,In_2849);
xnor U288 (N_288,In_1560,In_2855);
xor U289 (N_289,In_134,In_1662);
nand U290 (N_290,In_2213,In_445);
nor U291 (N_291,In_2142,In_1422);
xnor U292 (N_292,In_1110,In_281);
nor U293 (N_293,In_1636,In_1385);
nor U294 (N_294,In_2610,In_2010);
and U295 (N_295,In_780,In_2874);
or U296 (N_296,In_1714,In_684);
nor U297 (N_297,In_2976,In_1150);
nor U298 (N_298,In_1873,In_2093);
nand U299 (N_299,In_2404,In_2100);
or U300 (N_300,In_1383,In_1474);
xor U301 (N_301,In_2352,In_192);
and U302 (N_302,In_23,In_2941);
nor U303 (N_303,In_2764,In_1062);
and U304 (N_304,In_2239,In_2795);
xor U305 (N_305,In_2514,In_1029);
nand U306 (N_306,In_2528,In_2455);
nand U307 (N_307,In_962,In_2539);
and U308 (N_308,In_245,In_135);
nor U309 (N_309,In_2477,In_2803);
nand U310 (N_310,In_2666,In_2053);
nor U311 (N_311,In_274,In_2515);
or U312 (N_312,In_1876,In_28);
nand U313 (N_313,In_644,In_288);
nand U314 (N_314,In_208,In_2493);
or U315 (N_315,In_2559,In_930);
nand U316 (N_316,In_1208,In_237);
nand U317 (N_317,In_2098,In_2661);
nor U318 (N_318,In_880,In_951);
nand U319 (N_319,In_456,In_2875);
nand U320 (N_320,In_2813,In_561);
nor U321 (N_321,In_1954,In_512);
nor U322 (N_322,In_1813,In_1051);
nand U323 (N_323,In_738,In_2083);
nor U324 (N_324,In_1258,In_15);
or U325 (N_325,In_998,In_1143);
nand U326 (N_326,In_1263,In_2095);
nor U327 (N_327,In_669,In_385);
or U328 (N_328,In_1784,In_2668);
xnor U329 (N_329,In_315,In_2897);
nand U330 (N_330,In_629,In_1748);
and U331 (N_331,In_2824,In_995);
xor U332 (N_332,In_1801,In_163);
xnor U333 (N_333,In_1171,In_1979);
xor U334 (N_334,In_2118,In_2016);
nand U335 (N_335,In_2814,In_1397);
nor U336 (N_336,In_1591,In_1738);
or U337 (N_337,In_2609,In_767);
xor U338 (N_338,In_1629,In_789);
nand U339 (N_339,In_105,In_2845);
nor U340 (N_340,In_1734,In_876);
xnor U341 (N_341,In_340,In_1444);
or U342 (N_342,In_1884,In_1132);
nor U343 (N_343,In_342,In_1755);
nand U344 (N_344,In_203,In_947);
nor U345 (N_345,In_1669,In_849);
and U346 (N_346,In_2320,In_1811);
nand U347 (N_347,In_2618,In_1456);
or U348 (N_348,In_2904,In_2582);
nand U349 (N_349,In_550,In_2505);
or U350 (N_350,In_2809,In_982);
nand U351 (N_351,In_2002,In_853);
and U352 (N_352,In_1575,In_848);
xor U353 (N_353,In_726,In_2906);
and U354 (N_354,In_1637,In_1219);
xnor U355 (N_355,In_306,In_953);
xor U356 (N_356,In_1152,In_2096);
xnor U357 (N_357,In_214,In_212);
nand U358 (N_358,In_2047,In_2222);
and U359 (N_359,In_443,In_1404);
xnor U360 (N_360,In_14,In_2744);
nor U361 (N_361,In_2921,In_2617);
nand U362 (N_362,In_991,In_802);
xnor U363 (N_363,In_599,In_1541);
nor U364 (N_364,In_609,In_236);
and U365 (N_365,In_302,In_718);
xnor U366 (N_366,In_1126,In_2151);
xor U367 (N_367,In_266,In_110);
or U368 (N_368,In_1018,In_1403);
or U369 (N_369,In_1994,In_2364);
and U370 (N_370,In_2498,In_2244);
nor U371 (N_371,In_202,In_397);
and U372 (N_372,In_1101,In_2737);
xor U373 (N_373,In_847,In_2237);
or U374 (N_374,In_986,In_1191);
nor U375 (N_375,In_1475,In_2197);
nor U376 (N_376,In_416,In_2639);
xor U377 (N_377,In_1788,In_440);
nand U378 (N_378,In_1293,In_102);
xnor U379 (N_379,In_1023,In_1777);
nor U380 (N_380,In_1655,In_2986);
and U381 (N_381,In_1396,In_739);
xor U382 (N_382,In_2063,In_1100);
and U383 (N_383,In_2338,In_2458);
xor U384 (N_384,In_1272,In_1222);
xnor U385 (N_385,In_1105,In_1286);
nor U386 (N_386,In_837,In_634);
xor U387 (N_387,In_1490,In_2431);
nand U388 (N_388,In_2055,In_2488);
nand U389 (N_389,In_1720,In_419);
nand U390 (N_390,In_1539,In_1235);
and U391 (N_391,In_2210,In_1808);
or U392 (N_392,In_1948,In_2698);
and U393 (N_393,In_668,In_2086);
xor U394 (N_394,In_9,In_1564);
or U395 (N_395,In_44,In_1343);
and U396 (N_396,In_1154,In_2416);
xor U397 (N_397,In_415,In_1055);
xor U398 (N_398,In_1918,In_1892);
nor U399 (N_399,In_2040,In_1012);
and U400 (N_400,In_2422,In_681);
nor U401 (N_401,In_1592,In_2758);
or U402 (N_402,In_2563,In_1790);
and U403 (N_403,In_575,In_1567);
nor U404 (N_404,In_2032,In_241);
or U405 (N_405,In_1837,In_2686);
or U406 (N_406,In_2975,In_2024);
xnor U407 (N_407,In_690,In_1059);
nand U408 (N_408,In_560,In_537);
xnor U409 (N_409,In_2776,In_2384);
nand U410 (N_410,In_1075,In_396);
nor U411 (N_411,In_1512,In_1988);
xor U412 (N_412,In_1906,In_671);
xor U413 (N_413,In_637,In_478);
and U414 (N_414,In_1002,In_779);
xnor U415 (N_415,In_2826,In_1717);
and U416 (N_416,In_836,In_1980);
or U417 (N_417,In_2105,In_294);
xor U418 (N_418,In_749,In_832);
nand U419 (N_419,In_279,In_2745);
xnor U420 (N_420,In_148,In_48);
nand U421 (N_421,In_1550,In_2635);
and U422 (N_422,In_769,In_298);
or U423 (N_423,In_1227,In_1522);
xnor U424 (N_424,In_2453,In_45);
xnor U425 (N_425,In_1001,In_2227);
nor U426 (N_426,In_1698,In_788);
or U427 (N_427,In_2557,In_2132);
or U428 (N_428,In_2368,In_2410);
or U429 (N_429,In_731,In_2859);
and U430 (N_430,In_2780,In_2950);
or U431 (N_431,In_1327,In_1076);
xnor U432 (N_432,In_1453,In_850);
or U433 (N_433,In_2189,In_1724);
nor U434 (N_434,In_2566,In_501);
and U435 (N_435,In_2880,In_1695);
xor U436 (N_436,In_167,In_460);
or U437 (N_437,In_508,In_728);
nand U438 (N_438,In_424,In_2268);
or U439 (N_439,In_1728,In_1036);
and U440 (N_440,In_1814,In_2276);
xnor U441 (N_441,In_470,In_57);
xor U442 (N_442,In_1238,In_444);
xor U443 (N_443,In_1409,In_95);
or U444 (N_444,In_1582,In_2473);
or U445 (N_445,In_1292,In_374);
or U446 (N_446,In_2958,In_2910);
and U447 (N_447,In_1771,In_770);
nor U448 (N_448,In_448,In_626);
and U449 (N_449,In_124,In_883);
or U450 (N_450,In_308,In_1209);
nor U451 (N_451,In_2708,In_1946);
nor U452 (N_452,In_2220,In_2759);
or U453 (N_453,In_68,In_399);
nand U454 (N_454,In_1186,In_997);
nand U455 (N_455,In_2529,In_139);
xor U456 (N_456,In_2980,In_2903);
nor U457 (N_457,In_2997,In_818);
nor U458 (N_458,In_1792,In_1398);
and U459 (N_459,In_2932,In_861);
or U460 (N_460,In_2318,In_2008);
or U461 (N_461,In_1479,In_145);
xor U462 (N_462,In_2262,In_1334);
and U463 (N_463,In_2577,In_2894);
xnor U464 (N_464,In_1241,In_844);
and U465 (N_465,In_2012,In_2374);
or U466 (N_466,In_314,In_2433);
xnor U467 (N_467,In_674,In_1095);
or U468 (N_468,In_491,In_784);
nand U469 (N_469,In_2141,In_2266);
or U470 (N_470,In_2517,In_2203);
nor U471 (N_471,In_240,In_2601);
or U472 (N_472,In_1859,In_1585);
nor U473 (N_473,In_768,In_1052);
and U474 (N_474,In_954,In_2108);
nor U475 (N_475,In_2143,In_2409);
or U476 (N_476,In_290,In_1060);
or U477 (N_477,In_76,In_2013);
xnor U478 (N_478,In_856,In_231);
or U479 (N_479,In_1216,In_125);
and U480 (N_480,In_194,In_1901);
xnor U481 (N_481,In_1712,In_2427);
xnor U482 (N_482,In_2344,In_149);
and U483 (N_483,In_1962,In_2106);
nor U484 (N_484,In_527,In_969);
nand U485 (N_485,In_2248,In_1608);
and U486 (N_486,In_2370,In_2243);
and U487 (N_487,In_1943,In_741);
xor U488 (N_488,In_2456,In_2171);
nor U489 (N_489,In_1547,In_1435);
and U490 (N_490,In_2333,In_2751);
and U491 (N_491,In_1434,In_1252);
nand U492 (N_492,In_2199,In_1666);
or U493 (N_493,In_312,In_2665);
and U494 (N_494,In_467,In_1909);
or U495 (N_495,In_2296,In_364);
xor U496 (N_496,In_2067,In_354);
and U497 (N_497,In_2360,In_255);
nand U498 (N_498,In_1407,In_1898);
or U499 (N_499,In_2696,In_50);
xor U500 (N_500,In_249,In_2878);
and U501 (N_501,N_497,N_238);
or U502 (N_502,In_2161,In_2018);
nor U503 (N_503,N_56,N_16);
or U504 (N_504,In_2562,In_318);
and U505 (N_505,In_2818,In_1330);
and U506 (N_506,In_49,In_1365);
and U507 (N_507,In_1847,In_1484);
nor U508 (N_508,In_2369,In_504);
xnor U509 (N_509,N_312,In_723);
nand U510 (N_510,N_479,In_2660);
or U511 (N_511,In_2200,In_69);
xor U512 (N_512,In_1702,In_1745);
nand U513 (N_513,In_2387,In_2974);
or U514 (N_514,N_52,In_1820);
and U515 (N_515,In_1947,N_426);
and U516 (N_516,In_1151,N_428);
xnor U517 (N_517,N_379,N_129);
nor U518 (N_518,N_7,In_624);
xor U519 (N_519,In_572,N_119);
and U520 (N_520,In_1588,In_346);
and U521 (N_521,In_2490,In_270);
or U522 (N_522,In_2123,N_217);
or U523 (N_523,In_1604,N_42);
and U524 (N_524,In_799,In_2561);
and U525 (N_525,In_2359,In_1780);
or U526 (N_526,N_464,In_2122);
and U527 (N_527,In_961,In_2463);
xor U528 (N_528,In_1184,In_1041);
and U529 (N_529,In_1268,In_2928);
or U530 (N_530,In_2977,In_842);
xor U531 (N_531,In_1233,In_2183);
or U532 (N_532,In_1274,In_1016);
nor U533 (N_533,In_785,N_272);
or U534 (N_534,In_401,N_283);
xor U535 (N_535,In_499,In_2211);
and U536 (N_536,In_2277,N_323);
nor U537 (N_537,In_2863,In_1584);
and U538 (N_538,In_687,In_1831);
nor U539 (N_539,N_386,In_1797);
xnor U540 (N_540,In_819,In_137);
or U541 (N_541,In_2636,In_2450);
or U542 (N_542,In_476,N_437);
and U543 (N_543,In_515,In_1064);
xor U544 (N_544,In_493,In_1360);
nand U545 (N_545,In_1914,In_719);
nor U546 (N_546,In_822,N_355);
and U547 (N_547,In_2425,In_971);
xor U548 (N_548,In_772,In_1194);
nand U549 (N_549,In_1791,In_860);
xnor U550 (N_550,In_205,In_363);
nor U551 (N_551,In_1180,In_2020);
nand U552 (N_552,In_1849,In_2877);
nand U553 (N_553,In_126,In_2738);
xor U554 (N_554,In_2533,In_896);
nor U555 (N_555,N_225,In_322);
nor U556 (N_556,In_699,In_2673);
nand U557 (N_557,In_1862,N_76);
xor U558 (N_558,In_937,In_1445);
nor U559 (N_559,In_2006,In_2460);
nor U560 (N_560,In_569,In_1491);
nor U561 (N_561,In_2247,N_168);
nand U562 (N_562,N_324,In_441);
nand U563 (N_563,In_1044,In_403);
xor U564 (N_564,In_620,In_1145);
nand U565 (N_565,In_5,In_2624);
or U566 (N_566,In_2850,In_2403);
xnor U567 (N_567,In_2710,In_513);
nand U568 (N_568,In_2642,In_1178);
nand U569 (N_569,N_218,In_2499);
nor U570 (N_570,In_2724,In_2470);
and U571 (N_571,In_2564,In_1169);
nor U572 (N_572,N_423,In_2451);
nand U573 (N_573,In_591,In_1812);
or U574 (N_574,N_381,In_217);
or U575 (N_575,In_170,In_1307);
or U576 (N_576,In_610,N_484);
xnor U577 (N_577,In_83,In_935);
nor U578 (N_578,In_1505,In_2508);
nand U579 (N_579,In_2588,N_35);
xor U580 (N_580,In_831,In_1767);
nor U581 (N_581,In_175,N_3);
nand U582 (N_582,In_2074,In_925);
nor U583 (N_583,N_214,In_2149);
xor U584 (N_584,In_1433,In_119);
and U585 (N_585,In_183,In_2773);
and U586 (N_586,In_1454,In_2382);
nand U587 (N_587,In_965,In_2283);
nand U588 (N_588,N_399,In_744);
nand U589 (N_589,In_1830,In_1538);
and U590 (N_590,In_1008,In_2261);
xnor U591 (N_591,N_370,In_1193);
nor U592 (N_592,In_960,In_1961);
xnor U593 (N_593,In_1942,In_2584);
xor U594 (N_594,In_1414,In_1690);
nand U595 (N_595,In_1599,N_50);
nor U596 (N_596,In_2116,In_1319);
xor U597 (N_597,In_350,In_447);
xor U598 (N_598,In_2743,In_580);
and U599 (N_599,N_253,In_2117);
nor U600 (N_600,N_84,N_442);
xnor U601 (N_601,In_2599,In_1084);
xnor U602 (N_602,N_452,In_1860);
nor U603 (N_603,In_224,In_2424);
nor U604 (N_604,In_2633,In_2954);
or U605 (N_605,N_384,In_168);
nand U606 (N_606,In_1405,In_1402);
nand U607 (N_607,In_596,In_2873);
nor U608 (N_608,In_1530,In_2026);
or U609 (N_609,In_2441,In_35);
or U610 (N_610,In_100,In_2658);
and U611 (N_611,N_316,In_2571);
and U612 (N_612,N_154,In_595);
nor U613 (N_613,In_775,In_530);
xnor U614 (N_614,In_1305,In_1262);
or U615 (N_615,In_238,In_1423);
xor U616 (N_616,In_2677,N_106);
or U617 (N_617,In_2621,N_162);
xor U618 (N_618,In_2867,In_1982);
nor U619 (N_619,In_492,In_2769);
xnor U620 (N_620,In_2231,In_2735);
nor U621 (N_621,In_2644,In_616);
and U622 (N_622,N_333,In_2019);
nor U623 (N_623,In_1225,In_1206);
nor U624 (N_624,In_407,N_315);
nor U625 (N_625,In_1993,In_2082);
and U626 (N_626,In_1703,In_356);
and U627 (N_627,In_1950,In_111);
and U628 (N_628,In_2469,N_346);
nor U629 (N_629,N_203,N_161);
and U630 (N_630,In_438,In_523);
nor U631 (N_631,In_1432,In_1026);
nor U632 (N_632,N_302,In_826);
or U633 (N_633,In_2255,In_353);
or U634 (N_634,In_2579,N_494);
xnor U635 (N_635,N_107,In_1868);
xor U636 (N_636,In_1607,In_594);
nand U637 (N_637,In_475,N_98);
xor U638 (N_638,In_2693,In_411);
nand U639 (N_639,In_1480,N_258);
or U640 (N_640,In_1509,In_1969);
and U641 (N_641,In_1796,In_927);
xor U642 (N_642,N_115,In_1389);
xor U643 (N_643,In_1118,In_2722);
nand U644 (N_644,In_2729,N_69);
and U645 (N_645,In_388,In_1408);
or U646 (N_646,N_164,N_151);
nand U647 (N_647,In_2043,In_708);
nor U648 (N_648,In_234,N_138);
nor U649 (N_649,In_272,N_15);
and U650 (N_650,In_2388,In_394);
and U651 (N_651,In_1278,N_184);
or U652 (N_652,In_1516,In_166);
nand U653 (N_653,N_44,In_1325);
or U654 (N_654,In_1063,In_2606);
or U655 (N_655,N_347,In_1559);
nor U656 (N_656,In_221,In_2730);
or U657 (N_657,N_461,In_940);
or U658 (N_658,N_257,N_210);
nand U659 (N_659,In_251,In_2663);
or U660 (N_660,In_2823,In_1937);
nor U661 (N_661,N_10,In_1320);
nand U662 (N_662,In_2989,In_795);
and U663 (N_663,In_2264,In_1120);
or U664 (N_664,N_486,In_1089);
and U665 (N_665,In_656,In_2365);
and U666 (N_666,N_185,N_392);
xnor U667 (N_667,In_178,In_2492);
xor U668 (N_668,N_20,In_2349);
xnor U669 (N_669,In_2833,In_1804);
nor U670 (N_670,In_1205,In_1744);
xnor U671 (N_671,In_1934,In_1202);
and U672 (N_672,N_265,In_1010);
nor U673 (N_673,In_2472,In_20);
nand U674 (N_674,In_1321,In_2185);
xnor U675 (N_675,In_1763,In_19);
xnor U676 (N_676,In_2130,N_466);
xor U677 (N_677,In_2152,In_602);
xnor U678 (N_678,N_13,In_2967);
nand U679 (N_679,In_2519,In_2888);
or U680 (N_680,In_355,In_1447);
and U681 (N_681,N_47,In_2944);
and U682 (N_682,In_613,In_2476);
and U683 (N_683,In_1437,In_138);
nor U684 (N_684,N_160,In_899);
and U685 (N_685,In_538,In_159);
nand U686 (N_686,N_19,In_1213);
nand U687 (N_687,In_1392,In_2235);
xor U688 (N_688,In_2170,In_1187);
and U689 (N_689,N_144,In_1472);
nand U690 (N_690,In_2080,In_598);
xor U691 (N_691,In_2790,In_173);
and U692 (N_692,In_295,In_2021);
nand U693 (N_693,In_1215,In_1936);
xnor U694 (N_694,In_1944,In_413);
xnor U695 (N_695,N_36,In_151);
nand U696 (N_696,In_2650,In_1821);
nor U697 (N_697,N_314,In_841);
nor U698 (N_698,In_1173,In_1123);
nand U699 (N_699,In_2627,In_1577);
nand U700 (N_700,In_1250,In_2952);
nor U701 (N_701,In_859,In_141);
and U702 (N_702,In_2805,N_59);
or U703 (N_703,In_2417,In_2691);
xor U704 (N_704,In_140,In_964);
nor U705 (N_705,In_1902,In_1185);
nor U706 (N_706,In_2865,In_1113);
or U707 (N_707,In_360,In_2558);
nor U708 (N_708,In_271,In_1376);
and U709 (N_709,In_693,In_1104);
and U710 (N_710,In_903,In_2792);
nor U711 (N_711,N_30,In_2190);
and U712 (N_712,In_1705,In_2061);
or U713 (N_713,N_235,In_2314);
nor U714 (N_714,N_388,In_1439);
xor U715 (N_715,N_17,In_117);
and U716 (N_716,In_1157,In_2319);
or U717 (N_717,In_1338,In_41);
or U718 (N_718,In_325,In_1426);
nor U719 (N_719,In_1431,In_794);
nand U720 (N_720,In_2844,In_477);
nand U721 (N_721,In_1078,In_2872);
or U722 (N_722,N_43,In_2794);
nand U723 (N_723,In_398,N_402);
or U724 (N_724,In_967,N_369);
nand U725 (N_725,In_2586,In_980);
nand U726 (N_726,In_2821,N_443);
and U727 (N_727,In_1058,N_433);
xnor U728 (N_728,In_2180,In_29);
and U729 (N_729,In_450,In_2616);
or U730 (N_730,In_1514,In_1312);
and U731 (N_731,In_160,In_2206);
nand U732 (N_732,In_345,In_2363);
xor U733 (N_733,In_1927,In_919);
or U734 (N_734,N_425,N_222);
or U735 (N_735,In_2175,In_551);
nand U736 (N_736,In_2069,N_291);
nor U737 (N_737,In_1563,In_1372);
nand U738 (N_738,In_701,In_1499);
nor U739 (N_739,In_536,In_2484);
xnor U740 (N_740,N_249,In_619);
nand U741 (N_741,In_632,N_361);
xor U742 (N_742,In_2925,N_348);
or U743 (N_743,In_1891,In_2526);
nor U744 (N_744,N_389,In_2835);
nand U745 (N_745,In_654,In_372);
nand U746 (N_746,N_67,N_290);
and U747 (N_747,In_689,In_2418);
or U748 (N_748,In_2090,In_968);
or U749 (N_749,In_754,In_387);
nand U750 (N_750,In_526,N_147);
or U751 (N_751,In_2870,N_487);
nor U752 (N_752,N_244,In_1015);
and U753 (N_753,N_396,In_34);
or U754 (N_754,In_2896,In_1290);
or U755 (N_755,In_2996,In_1275);
xor U756 (N_756,In_1885,In_932);
xor U757 (N_757,In_2953,In_1601);
or U758 (N_758,In_2556,In_1468);
or U759 (N_759,In_2158,In_1694);
xor U760 (N_760,In_521,In_2380);
or U761 (N_761,In_423,In_2278);
nor U762 (N_762,In_46,In_32);
or U763 (N_763,N_137,In_539);
nor U764 (N_764,N_71,In_2039);
nand U765 (N_765,In_2188,N_321);
nand U766 (N_766,In_1742,In_1879);
xor U767 (N_767,In_1673,In_615);
nand U768 (N_768,In_1926,In_291);
and U769 (N_769,In_2186,In_1832);
xnor U770 (N_770,In_2031,In_1659);
or U771 (N_771,In_531,In_712);
or U772 (N_772,In_999,In_2572);
nor U773 (N_773,In_608,In_643);
nor U774 (N_774,In_1566,In_1463);
nand U775 (N_775,In_750,In_1800);
nand U776 (N_776,In_540,In_451);
nor U777 (N_777,In_1858,In_720);
and U778 (N_778,In_2408,N_387);
and U779 (N_779,In_2274,N_170);
xor U780 (N_780,N_174,N_248);
nand U781 (N_781,In_1077,In_2316);
or U782 (N_782,In_809,In_278);
nor U783 (N_783,In_1839,In_265);
nand U784 (N_784,In_43,In_559);
or U785 (N_785,In_1109,In_1332);
xnor U786 (N_786,N_134,In_1888);
xnor U787 (N_787,In_546,In_1406);
xor U788 (N_788,N_362,In_1240);
or U789 (N_789,In_16,N_459);
xnor U790 (N_790,N_401,In_1568);
or U791 (N_791,N_318,In_2267);
and U792 (N_792,In_2280,N_376);
xor U793 (N_793,In_1919,In_2513);
or U794 (N_794,N_234,In_1496);
or U795 (N_795,In_563,In_2940);
xor U796 (N_796,In_38,In_2549);
nor U797 (N_797,In_1628,In_1368);
nor U798 (N_798,In_2626,N_213);
nand U799 (N_799,In_2819,N_237);
xor U800 (N_800,In_232,N_308);
nor U801 (N_801,N_462,In_1618);
nor U802 (N_802,In_1798,In_2652);
xor U803 (N_803,In_2334,N_394);
or U804 (N_804,In_1092,In_1482);
nor U805 (N_805,In_2496,In_106);
and U806 (N_806,In_2902,N_406);
nand U807 (N_807,N_419,In_297);
nand U808 (N_808,In_1682,N_187);
nor U809 (N_809,In_182,In_1930);
or U810 (N_810,N_31,N_463);
nor U811 (N_811,In_334,In_2303);
and U812 (N_812,In_2784,N_27);
and U813 (N_813,In_1977,N_492);
nor U814 (N_814,N_349,In_1163);
xor U815 (N_815,N_311,In_2343);
nand U816 (N_816,In_2828,In_2911);
or U817 (N_817,In_2643,In_239);
xor U818 (N_818,In_1034,In_717);
and U819 (N_819,In_1903,In_2014);
nand U820 (N_820,In_1506,In_2962);
or U821 (N_821,N_471,In_348);
nor U822 (N_822,In_1181,In_2651);
nor U823 (N_823,In_122,N_57);
and U824 (N_824,In_558,In_757);
nor U825 (N_825,In_2858,In_2407);
nor U826 (N_826,N_171,In_581);
or U827 (N_827,In_1989,N_310);
or U828 (N_828,In_2341,In_2540);
nand U829 (N_829,N_284,In_2224);
xnor U830 (N_830,In_152,In_2154);
nand U831 (N_831,In_11,In_2659);
or U832 (N_832,In_1418,In_2541);
xnor U833 (N_833,N_322,In_47);
or U834 (N_834,In_894,N_227);
nor U835 (N_835,In_2548,In_2982);
or U836 (N_836,In_331,In_1917);
nand U837 (N_837,In_707,In_2246);
and U838 (N_838,In_2449,In_1907);
nor U839 (N_839,In_1576,In_506);
nor U840 (N_840,In_1218,In_2181);
nand U841 (N_841,In_1970,In_2233);
nor U842 (N_842,N_116,In_1156);
xnor U843 (N_843,In_1641,In_1580);
nand U844 (N_844,In_683,In_511);
or U845 (N_845,In_1686,N_8);
nor U846 (N_846,In_1616,In_1155);
nor U847 (N_847,In_2507,N_211);
nand U848 (N_848,In_973,In_2709);
or U849 (N_849,In_1886,In_2984);
xor U850 (N_850,N_232,N_498);
nor U851 (N_851,In_1625,In_262);
and U852 (N_852,In_630,N_55);
and U853 (N_853,In_2419,In_2402);
xor U854 (N_854,In_2783,In_820);
xnor U855 (N_855,N_202,In_1590);
or U856 (N_856,In_2379,N_303);
nor U857 (N_857,N_328,In_1846);
or U858 (N_858,In_1976,In_75);
or U859 (N_859,In_1996,In_2992);
nor U860 (N_860,In_918,N_282);
nor U861 (N_861,N_289,In_33);
nor U862 (N_862,In_910,In_64);
nor U863 (N_863,In_2377,In_1707);
xor U864 (N_864,In_1103,In_2847);
and U865 (N_865,In_823,In_607);
xor U866 (N_866,N_141,In_2619);
and U867 (N_867,N_157,N_72);
or U868 (N_868,In_184,In_777);
or U869 (N_869,In_1864,In_1136);
nand U870 (N_870,In_839,In_1693);
or U871 (N_871,N_473,In_1692);
xnor U872 (N_872,In_542,In_665);
or U873 (N_873,In_2160,N_382);
or U874 (N_874,In_1774,In_2781);
nor U875 (N_875,N_354,In_1363);
or U876 (N_876,In_490,In_2893);
and U877 (N_877,In_386,N_37);
or U878 (N_878,In_1605,In_1663);
nor U879 (N_879,In_2107,In_1649);
xnor U880 (N_880,In_1805,In_1464);
xor U881 (N_881,In_722,In_1701);
and U882 (N_882,In_1053,In_2555);
nor U883 (N_883,In_2509,N_489);
xnor U884 (N_884,In_532,In_790);
or U885 (N_885,In_2527,In_1446);
nand U886 (N_886,In_2494,In_2392);
and U887 (N_887,In_1093,In_827);
and U888 (N_888,N_169,In_2272);
nand U889 (N_889,N_435,In_58);
and U890 (N_890,In_144,In_2165);
or U891 (N_891,In_1037,N_383);
or U892 (N_892,In_2637,N_407);
nand U893 (N_893,In_816,N_124);
and U894 (N_894,In_1558,In_1166);
or U895 (N_895,In_93,In_1985);
and U896 (N_896,In_1204,N_374);
nor U897 (N_897,In_1267,In_1731);
xnor U898 (N_898,In_13,In_1722);
nor U899 (N_899,In_1834,In_1895);
or U900 (N_900,In_1230,In_180);
nor U901 (N_901,In_418,In_1176);
or U902 (N_902,N_496,N_465);
nand U903 (N_903,In_1555,In_2534);
xnor U904 (N_904,N_178,In_2886);
nand U905 (N_905,N_475,In_227);
nand U906 (N_906,In_2596,In_1006);
or U907 (N_907,N_292,In_1586);
and U908 (N_908,N_408,N_231);
and U909 (N_909,In_1773,In_2438);
or U910 (N_910,In_190,In_3);
nor U911 (N_911,N_417,In_1387);
xnor U912 (N_912,N_280,In_2657);
nor U913 (N_913,N_48,In_588);
nand U914 (N_914,In_2389,In_223);
nor U915 (N_915,In_2302,In_2909);
nand U916 (N_916,In_2015,In_1708);
and U917 (N_917,In_1932,In_2576);
nand U918 (N_918,In_2603,In_1024);
xor U919 (N_919,In_2861,In_808);
or U920 (N_920,In_1175,N_422);
xnor U921 (N_921,In_871,N_424);
xor U922 (N_922,In_828,In_2312);
xor U923 (N_923,In_1243,In_1207);
and U924 (N_924,N_350,N_183);
or U925 (N_925,In_2315,In_1964);
nor U926 (N_926,In_71,In_1322);
xnor U927 (N_927,In_1270,In_2753);
or U928 (N_928,In_128,In_464);
or U929 (N_929,N_45,In_2786);
nor U930 (N_930,N_270,In_1983);
nand U931 (N_931,In_1280,In_230);
xor U932 (N_932,In_248,In_1968);
nand U933 (N_933,In_1356,In_2279);
xor U934 (N_934,In_1079,In_1345);
nand U935 (N_935,In_435,In_1613);
and U936 (N_936,In_282,In_564);
and U937 (N_937,In_327,In_2256);
nand U938 (N_938,In_1190,In_916);
and U939 (N_939,In_2308,In_1760);
or U940 (N_940,In_522,In_677);
xnor U941 (N_941,N_28,In_2695);
nand U942 (N_942,In_485,In_676);
nand U943 (N_943,In_1975,In_2938);
or U944 (N_944,N_53,In_2892);
xnor U945 (N_945,In_53,In_2914);
xor U946 (N_946,N_21,In_453);
and U947 (N_947,In_943,In_2129);
xor U948 (N_948,N_51,N_409);
nand U949 (N_949,N_208,In_1357);
nor U950 (N_950,N_216,In_2620);
nor U951 (N_951,N_454,In_330);
and U952 (N_952,In_1382,In_2342);
or U953 (N_953,In_2669,In_2275);
and U954 (N_954,N_341,In_2749);
and U955 (N_955,In_2771,In_1344);
nand U956 (N_956,In_1436,N_483);
and U957 (N_957,In_893,In_793);
nor U958 (N_958,N_123,N_130);
nor U959 (N_959,In_2085,In_2194);
or U960 (N_960,N_447,In_1740);
or U961 (N_961,In_1009,In_2615);
and U962 (N_962,N_367,In_1161);
nand U963 (N_963,In_2923,In_612);
nor U964 (N_964,In_2683,In_1851);
and U965 (N_965,In_1921,In_18);
nand U966 (N_966,In_176,N_63);
nor U967 (N_967,In_370,N_421);
xnor U968 (N_968,In_2166,In_796);
nand U969 (N_969,In_2808,In_2201);
nor U970 (N_970,In_442,In_1562);
nor U971 (N_971,In_510,N_221);
nor U972 (N_972,In_486,N_4);
xnor U973 (N_973,In_1657,In_1667);
and U974 (N_974,In_289,In_2538);
and U975 (N_975,In_2725,In_939);
and U976 (N_976,N_9,N_191);
nor U977 (N_977,In_247,N_109);
nor U978 (N_978,In_2223,In_204);
and U979 (N_979,N_274,N_165);
nand U980 (N_980,N_485,N_58);
xnor U981 (N_981,In_2390,In_2293);
nand U982 (N_982,N_180,In_2030);
nand U983 (N_983,In_1769,In_863);
nor U984 (N_984,N_295,In_732);
and U985 (N_985,N_418,In_518);
xnor U986 (N_986,N_136,In_2475);
xor U987 (N_987,In_2084,In_269);
and U988 (N_988,In_2685,In_1674);
nor U989 (N_989,In_2208,In_2837);
nor U990 (N_990,In_200,In_2817);
or U991 (N_991,In_1865,In_1923);
nor U992 (N_992,N_336,In_952);
nor U993 (N_993,In_543,In_1254);
and U994 (N_994,N_177,N_335);
xor U995 (N_995,In_1986,In_2078);
or U996 (N_996,In_2238,In_2945);
or U997 (N_997,In_277,In_1861);
xor U998 (N_998,In_2310,In_1759);
or U999 (N_999,In_1416,In_714);
and U1000 (N_1000,In_1147,N_783);
nand U1001 (N_1001,In_1999,In_2511);
nand U1002 (N_1002,N_537,In_2727);
xor U1003 (N_1003,In_2942,In_549);
nor U1004 (N_1004,N_194,In_2187);
nand U1005 (N_1005,N_104,N_701);
xnor U1006 (N_1006,N_444,N_131);
and U1007 (N_1007,In_762,N_812);
and U1008 (N_1008,N_476,N_166);
or U1009 (N_1009,In_2503,In_2936);
or U1010 (N_1010,In_2554,N_884);
and U1011 (N_1011,In_120,In_1442);
or U1012 (N_1012,In_395,N_250);
or U1013 (N_1013,In_2676,In_1139);
nor U1014 (N_1014,In_1341,N_205);
nand U1015 (N_1015,In_1492,In_215);
xnor U1016 (N_1016,In_1415,N_514);
nor U1017 (N_1017,N_919,N_904);
nand U1018 (N_1018,In_528,N_100);
and U1019 (N_1019,N_995,In_1260);
or U1020 (N_1020,In_2785,In_2580);
nor U1021 (N_1021,In_2301,In_1457);
and U1022 (N_1022,In_25,In_2812);
nor U1023 (N_1023,In_2924,N_879);
nand U1024 (N_1024,N_29,In_703);
or U1025 (N_1025,N_404,In_1284);
nor U1026 (N_1026,N_25,In_1273);
or U1027 (N_1027,In_1072,N_472);
nand U1028 (N_1028,In_1984,In_773);
and U1029 (N_1029,In_1214,In_2731);
or U1030 (N_1030,In_1782,N_307);
nand U1031 (N_1031,N_240,N_189);
nor U1032 (N_1032,In_2114,In_2358);
xor U1033 (N_1033,N_18,In_1140);
and U1034 (N_1034,In_2946,In_662);
nor U1035 (N_1035,N_246,In_1688);
and U1036 (N_1036,In_1729,In_990);
or U1037 (N_1037,In_2922,In_1634);
nand U1038 (N_1038,In_2772,N_737);
and U1039 (N_1039,N_913,In_377);
nor U1040 (N_1040,In_2207,In_2971);
nor U1041 (N_1041,N_618,In_2347);
nand U1042 (N_1042,N_656,In_905);
nand U1043 (N_1043,N_949,In_688);
and U1044 (N_1044,In_2196,In_1299);
xnor U1045 (N_1045,In_1642,N_903);
or U1046 (N_1046,In_1877,N_560);
nor U1047 (N_1047,In_1127,N_204);
xor U1048 (N_1048,N_532,In_1789);
xor U1049 (N_1049,In_2741,N_294);
xor U1050 (N_1050,N_747,In_2796);
and U1051 (N_1051,N_630,In_305);
xor U1052 (N_1052,In_2704,N_915);
nor U1053 (N_1053,In_1393,In_2332);
nor U1054 (N_1054,N_860,In_2250);
and U1055 (N_1055,N_689,In_104);
or U1056 (N_1056,In_2607,In_1595);
nor U1057 (N_1057,N_90,In_2628);
xor U1058 (N_1058,In_758,N_599);
xnor U1059 (N_1059,In_1925,In_1672);
nand U1060 (N_1060,In_855,In_2702);
nand U1061 (N_1061,N_105,In_1198);
nand U1062 (N_1062,In_1329,N_414);
or U1063 (N_1063,N_142,In_1347);
and U1064 (N_1064,In_1417,In_2327);
or U1065 (N_1065,N_300,In_838);
or U1066 (N_1066,N_754,In_1794);
or U1067 (N_1067,In_735,N_163);
nor U1068 (N_1068,In_525,N_750);
or U1069 (N_1069,N_681,N_12);
or U1070 (N_1070,N_611,N_121);
nand U1071 (N_1071,N_512,N_420);
or U1072 (N_1072,In_349,N_763);
nand U1073 (N_1073,In_1146,N_702);
and U1074 (N_1074,In_115,In_2990);
xor U1075 (N_1075,N_840,In_977);
nor U1076 (N_1076,In_1289,In_933);
xor U1077 (N_1077,N_501,In_2797);
nand U1078 (N_1078,N_930,In_1824);
nand U1079 (N_1079,In_1603,In_1028);
and U1080 (N_1080,In_2173,In_2937);
nor U1081 (N_1081,N_984,In_2916);
and U1082 (N_1082,In_889,In_1000);
xnor U1083 (N_1083,In_465,In_902);
xor U1084 (N_1084,In_191,In_2712);
or U1085 (N_1085,N_395,In_1856);
nand U1086 (N_1086,N_872,N_515);
xnor U1087 (N_1087,In_347,In_458);
nor U1088 (N_1088,In_639,In_496);
nand U1089 (N_1089,In_1210,N_523);
and U1090 (N_1090,N_547,In_189);
nor U1091 (N_1091,In_1793,In_854);
and U1092 (N_1092,In_2148,N_60);
or U1093 (N_1093,In_1882,N_644);
or U1094 (N_1094,In_2804,In_1401);
and U1095 (N_1095,In_371,In_2497);
nor U1096 (N_1096,N_922,N_659);
nor U1097 (N_1097,N_994,In_1314);
and U1098 (N_1098,In_601,N_309);
or U1099 (N_1099,In_2415,In_730);
nor U1100 (N_1100,N_590,In_2000);
nor U1101 (N_1101,N_658,In_1624);
or U1102 (N_1102,In_627,N_677);
nand U1103 (N_1103,In_1727,N_843);
xnor U1104 (N_1104,N_327,In_1291);
nor U1105 (N_1105,In_311,In_1633);
nand U1106 (N_1106,In_1974,In_1129);
and U1107 (N_1107,N_793,In_1529);
xnor U1108 (N_1108,In_1517,In_1875);
and U1109 (N_1109,In_2119,N_591);
or U1110 (N_1110,In_1735,In_1819);
nor U1111 (N_1111,In_2357,In_368);
nand U1112 (N_1112,N_690,In_1099);
xor U1113 (N_1113,In_179,N_197);
or U1114 (N_1114,N_828,In_2943);
nor U1115 (N_1115,In_264,In_1298);
nand U1116 (N_1116,In_2853,In_783);
xor U1117 (N_1117,In_2443,N_759);
xnor U1118 (N_1118,In_220,N_831);
or U1119 (N_1119,In_787,N_971);
and U1120 (N_1120,In_1309,N_206);
or U1121 (N_1121,In_829,In_1532);
and U1122 (N_1122,In_1420,In_702);
nand U1123 (N_1123,In_1141,N_732);
xor U1124 (N_1124,N_964,In_258);
and U1125 (N_1125,In_2252,N_713);
and U1126 (N_1126,In_976,In_2761);
xnor U1127 (N_1127,In_1513,In_2939);
nand U1128 (N_1128,N_623,N_377);
xor U1129 (N_1129,N_942,In_8);
or U1130 (N_1130,In_2305,In_2711);
and U1131 (N_1131,In_1085,N_236);
and U1132 (N_1132,In_171,In_98);
xnor U1133 (N_1133,In_2042,N_805);
nand U1134 (N_1134,N_874,N_145);
or U1135 (N_1135,In_2640,In_2815);
nor U1136 (N_1136,In_2523,N_807);
or U1137 (N_1137,N_802,In_1117);
xnor U1138 (N_1138,N_627,In_810);
and U1139 (N_1139,In_1795,N_990);
xor U1140 (N_1140,In_1351,In_1549);
nor U1141 (N_1141,N_636,N_542);
nand U1142 (N_1142,N_522,N_856);
xor U1143 (N_1143,N_541,In_2097);
or U1144 (N_1144,N_548,In_1889);
nor U1145 (N_1145,In_1571,N_719);
nor U1146 (N_1146,N_992,N_155);
xnor U1147 (N_1147,In_323,In_667);
nand U1148 (N_1148,In_1122,In_417);
and U1149 (N_1149,In_1485,In_571);
or U1150 (N_1150,In_1896,In_2072);
xnor U1151 (N_1151,N_778,In_2839);
and U1152 (N_1152,In_1236,In_786);
nor U1153 (N_1153,In_1887,N_101);
nand U1154 (N_1154,N_746,In_1504);
and U1155 (N_1155,N_474,In_2192);
xnor U1156 (N_1156,N_5,In_904);
xor U1157 (N_1157,N_671,In_2435);
or U1158 (N_1158,In_2931,In_2373);
nand U1159 (N_1159,N_956,In_2495);
and U1160 (N_1160,N_526,N_789);
and U1161 (N_1161,In_2740,N_688);
xor U1162 (N_1162,N_175,In_1069);
nor U1163 (N_1163,In_2478,In_1723);
and U1164 (N_1164,N_242,In_989);
xor U1165 (N_1165,N_781,N_808);
and U1166 (N_1166,N_816,In_1670);
nand U1167 (N_1167,N_676,N_207);
or U1168 (N_1168,In_181,N_567);
nand U1169 (N_1169,N_538,In_1685);
nor U1170 (N_1170,In_1476,In_425);
nor U1171 (N_1171,N_449,N_929);
and U1172 (N_1172,In_970,In_909);
or U1173 (N_1173,In_1096,N_862);
xnor U1174 (N_1174,N_456,N_761);
nor U1175 (N_1175,N_525,In_1938);
and U1176 (N_1176,In_884,N_756);
xor U1177 (N_1177,In_436,N_693);
nand U1178 (N_1178,In_162,N_803);
nand U1179 (N_1179,In_1019,In_1991);
xnor U1180 (N_1180,In_2664,N_524);
or U1181 (N_1181,In_1551,N_412);
nand U1182 (N_1182,N_871,N_865);
xor U1183 (N_1183,N_62,In_1753);
xor U1184 (N_1184,In_2273,In_1167);
nand U1185 (N_1185,N_65,N_585);
and U1186 (N_1186,N_298,N_439);
xnor U1187 (N_1187,N_952,In_782);
or U1188 (N_1188,In_2841,N_24);
and U1189 (N_1189,N_580,In_99);
nand U1190 (N_1190,N_950,In_67);
xnor U1191 (N_1191,In_2394,In_2791);
or U1192 (N_1192,N_400,N_112);
and U1193 (N_1193,In_2752,In_1536);
or U1194 (N_1194,N_641,N_985);
nand U1195 (N_1195,N_345,In_1040);
nand U1196 (N_1196,N_881,N_200);
nand U1197 (N_1197,In_1503,N_583);
or U1198 (N_1198,N_586,N_518);
nand U1199 (N_1199,N_563,In_618);
nand U1200 (N_1200,In_2714,N_707);
xnor U1201 (N_1201,In_872,N_743);
or U1202 (N_1202,N_642,In_2479);
and U1203 (N_1203,N_469,N_852);
xor U1204 (N_1204,In_2214,In_2376);
xnor U1205 (N_1205,In_2754,In_10);
or U1206 (N_1206,N_261,In_1452);
nand U1207 (N_1207,In_840,N_830);
and U1208 (N_1208,In_1627,N_695);
nand U1209 (N_1209,N_705,N_912);
xnor U1210 (N_1210,N_286,In_507);
and U1211 (N_1211,N_616,N_770);
xor U1212 (N_1212,N_75,In_293);
nand U1213 (N_1213,In_2887,In_1602);
nand U1214 (N_1214,In_617,In_2340);
or U1215 (N_1215,N_600,N_633);
xnor U1216 (N_1216,In_2028,In_2466);
nor U1217 (N_1217,N_159,In_1011);
or U1218 (N_1218,N_448,N_330);
nand U1219 (N_1219,N_193,N_715);
xor U1220 (N_1220,N_674,In_941);
and U1221 (N_1221,In_2457,N_457);
or U1222 (N_1222,In_2468,In_710);
or U1223 (N_1223,In_814,In_2440);
and U1224 (N_1224,In_1716,In_2793);
xnor U1225 (N_1225,In_1597,In_642);
or U1226 (N_1226,In_1112,N_536);
nor U1227 (N_1227,In_727,In_1318);
nand U1228 (N_1228,N_923,In_1587);
xnor U1229 (N_1229,In_922,In_1234);
or U1230 (N_1230,In_1257,In_2550);
or U1231 (N_1231,N_405,In_2822);
nand U1232 (N_1232,N_6,N_895);
nor U1233 (N_1233,N_212,In_936);
nand U1234 (N_1234,In_446,In_1683);
xnor U1235 (N_1235,N_415,In_1931);
and U1236 (N_1236,In_36,In_715);
xor U1237 (N_1237,In_2843,In_2198);
or U1238 (N_1238,In_1960,In_1916);
nand U1239 (N_1239,In_1495,N_143);
nand U1240 (N_1240,In_2504,In_1460);
nor U1241 (N_1241,N_331,In_695);
nor U1242 (N_1242,In_655,In_2502);
and U1243 (N_1243,In_2679,In_1410);
and U1244 (N_1244,In_1589,In_1741);
nor U1245 (N_1245,In_2050,In_697);
and U1246 (N_1246,In_452,In_759);
nor U1247 (N_1247,In_1199,In_1850);
xor U1248 (N_1248,In_1752,In_519);
nor U1249 (N_1249,In_1825,In_299);
and U1250 (N_1250,In_815,N_570);
xor U1251 (N_1251,In_1540,In_2480);
xor U1252 (N_1252,In_685,N_79);
or U1253 (N_1253,N_960,In_263);
and U1254 (N_1254,In_2348,In_2995);
or U1255 (N_1255,N_593,In_2901);
and U1256 (N_1256,In_376,In_1388);
nor U1257 (N_1257,N_795,In_1179);
nand U1258 (N_1258,N_883,N_342);
or U1259 (N_1259,N_598,In_1828);
or U1260 (N_1260,In_752,In_843);
nor U1261 (N_1261,In_2430,In_950);
xnor U1262 (N_1262,N_561,N_906);
xor U1263 (N_1263,N_122,In_1494);
nor U1264 (N_1264,In_2145,N_550);
nand U1265 (N_1265,In_1353,In_2768);
nor U1266 (N_1266,N_430,In_2842);
xor U1267 (N_1267,In_2983,N_458);
or U1268 (N_1268,N_390,In_544);
xor U1269 (N_1269,N_907,In_979);
and U1270 (N_1270,In_1277,In_2631);
or U1271 (N_1271,In_206,In_555);
xnor U1272 (N_1272,In_1025,N_179);
nor U1273 (N_1273,In_2212,In_1304);
or U1274 (N_1274,N_790,N_722);
nand U1275 (N_1275,In_2816,N_329);
or U1276 (N_1276,In_1806,In_392);
nand U1277 (N_1277,In_582,In_2287);
nand U1278 (N_1278,In_1678,In_2003);
and U1279 (N_1279,In_803,In_924);
nor U1280 (N_1280,In_2383,In_143);
xor U1281 (N_1281,In_1897,In_1953);
or U1282 (N_1282,N_753,N_724);
nor U1283 (N_1283,In_2613,N_751);
and U1284 (N_1284,In_1130,N_698);
or U1285 (N_1285,In_2081,N_545);
nand U1286 (N_1286,In_2733,In_1523);
or U1287 (N_1287,In_1121,In_621);
nor U1288 (N_1288,In_2317,N_827);
and U1289 (N_1289,N_986,N_398);
nand U1290 (N_1290,In_1328,In_1074);
or U1291 (N_1291,In_1049,In_1652);
and U1292 (N_1292,In_882,In_2885);
or U1293 (N_1293,In_1904,N_247);
nor U1294 (N_1294,In_1005,In_1905);
nor U1295 (N_1295,N_352,In_1826);
or U1296 (N_1296,In_1893,In_2981);
nand U1297 (N_1297,In_1778,N_173);
nor U1298 (N_1298,In_1162,N_578);
and U1299 (N_1299,In_2191,N_982);
nor U1300 (N_1300,In_1623,N_650);
nor U1301 (N_1301,In_1958,In_2289);
xnor U1302 (N_1302,N_635,N_140);
nand U1303 (N_1303,In_2895,In_481);
nor U1304 (N_1304,N_1,In_121);
nand U1305 (N_1305,N_468,In_1750);
or U1306 (N_1306,N_978,In_864);
xor U1307 (N_1307,N_645,In_1259);
nand U1308 (N_1308,In_2800,In_1283);
and U1309 (N_1309,In_2027,In_422);
nor U1310 (N_1310,In_1323,N_89);
nor U1311 (N_1311,N_796,N_577);
or U1312 (N_1312,In_1400,N_957);
nor U1313 (N_1313,In_2798,In_268);
nand U1314 (N_1314,N_64,In_2328);
nor U1315 (N_1315,In_577,In_1610);
nor U1316 (N_1316,In_2401,In_2300);
xor U1317 (N_1317,In_1654,N_385);
nor U1318 (N_1318,N_612,In_2623);
nand U1319 (N_1319,In_1583,In_565);
and U1320 (N_1320,N_317,N_135);
xnor U1321 (N_1321,In_2292,In_2670);
xnor U1322 (N_1322,N_799,In_480);
nand U1323 (N_1323,In_1115,In_1107);
nand U1324 (N_1324,N_182,In_1965);
xor U1325 (N_1325,N_279,N_275);
nand U1326 (N_1326,In_454,In_585);
xnor U1327 (N_1327,In_2632,In_157);
xnor U1328 (N_1328,N_103,N_38);
nor U1329 (N_1329,In_1620,In_196);
and U1330 (N_1330,In_2022,N_620);
or U1331 (N_1331,N_397,In_885);
or U1332 (N_1332,In_1626,In_2112);
nor U1333 (N_1333,In_2445,In_336);
and U1334 (N_1334,In_603,In_74);
xor U1335 (N_1335,In_877,In_2420);
xnor U1336 (N_1336,In_1978,N_631);
and U1337 (N_1337,In_2265,N_780);
nand U1338 (N_1338,In_283,In_548);
nand U1339 (N_1339,In_2929,N_337);
and U1340 (N_1340,In_59,In_817);
nand U1341 (N_1341,In_1335,In_2474);
xor U1342 (N_1342,N_2,N_167);
and U1343 (N_1343,N_933,N_555);
or U1344 (N_1344,N_708,N_82);
xor U1345 (N_1345,In_1489,N_565);
or U1346 (N_1346,N_926,In_1533);
nor U1347 (N_1347,In_1391,N_873);
and U1348 (N_1348,In_487,In_2385);
nand U1349 (N_1349,In_469,In_692);
nand U1350 (N_1350,N_804,In_1803);
or U1351 (N_1351,In_1990,In_2719);
or U1352 (N_1352,In_1863,In_2678);
nand U1353 (N_1353,In_1544,N_581);
nor U1354 (N_1354,In_24,N_969);
or U1355 (N_1355,N_495,N_326);
and U1356 (N_1356,In_886,N_558);
nand U1357 (N_1357,N_95,N_720);
xnor U1358 (N_1358,In_1569,In_2345);
and U1359 (N_1359,N_738,N_637);
or U1360 (N_1360,N_87,N_725);
xnor U1361 (N_1361,In_1955,N_975);
xnor U1362 (N_1362,N_277,N_557);
nand U1363 (N_1363,In_1758,In_1557);
or U1364 (N_1364,In_2518,N_520);
nand U1365 (N_1365,N_918,In_1048);
or U1366 (N_1366,N_605,In_1615);
nor U1367 (N_1367,In_1046,In_2917);
or U1368 (N_1368,In_1337,In_1848);
and U1369 (N_1369,In_432,In_1137);
xnor U1370 (N_1370,In_1370,In_1594);
and U1371 (N_1371,N_905,In_2765);
nand U1372 (N_1372,In_2680,N_325);
nor U1373 (N_1373,In_2985,In_158);
xor U1374 (N_1374,In_2068,N_584);
nor U1375 (N_1375,N_911,In_78);
and U1376 (N_1376,In_1061,In_2715);
and U1377 (N_1377,N_219,N_847);
xnor U1378 (N_1378,In_1957,In_584);
or U1379 (N_1379,In_587,N_268);
or U1380 (N_1380,In_2393,N_543);
nor U1381 (N_1381,In_1870,In_813);
and U1382 (N_1382,N_981,In_381);
xor U1383 (N_1383,In_2672,N_769);
xnor U1384 (N_1384,N_41,In_711);
and U1385 (N_1385,In_881,In_154);
and U1386 (N_1386,In_2056,In_2324);
nand U1387 (N_1387,N_776,N_609);
nor U1388 (N_1388,N_841,In_2414);
or U1389 (N_1389,N_506,N_684);
or U1390 (N_1390,In_7,N_987);
or U1391 (N_1391,N_40,In_606);
and U1392 (N_1392,N_158,In_640);
or U1393 (N_1393,In_409,In_1425);
and U1394 (N_1394,In_2788,In_1852);
nand U1395 (N_1395,In_219,N_646);
xnor U1396 (N_1396,In_439,In_1324);
xor U1397 (N_1397,N_953,N_838);
xnor U1398 (N_1398,In_39,N_810);
nor U1399 (N_1399,N_854,N_683);
nor U1400 (N_1400,In_2547,In_2133);
and U1401 (N_1401,In_2688,In_351);
or U1402 (N_1402,In_1271,In_1035);
or U1403 (N_1403,In_1192,In_1369);
nor U1404 (N_1404,In_2593,In_1467);
nor U1405 (N_1405,N_467,In_412);
xnor U1406 (N_1406,In_1424,In_1940);
and U1407 (N_1407,In_2064,N_220);
or U1408 (N_1408,N_771,N_516);
nor U1409 (N_1409,In_1013,In_1787);
nand U1410 (N_1410,In_226,N_993);
nor U1411 (N_1411,N_245,In_2560);
nand U1412 (N_1412,N_488,In_1614);
nor U1413 (N_1413,In_366,N_356);
or U1414 (N_1414,In_957,In_2583);
or U1415 (N_1415,In_673,In_1483);
and U1416 (N_1416,In_1966,In_858);
nand U1417 (N_1417,N_527,N_823);
xnor U1418 (N_1418,N_875,N_539);
and U1419 (N_1419,In_1004,In_686);
and U1420 (N_1420,In_2313,N_814);
nand U1421 (N_1421,In_1326,N_579);
and U1422 (N_1422,In_911,N_652);
and U1423 (N_1423,N_199,In_631);
nand U1424 (N_1424,In_1371,In_2400);
nor U1425 (N_1425,N_614,N_429);
and U1426 (N_1426,In_2035,N_726);
nor U1427 (N_1427,N_481,N_574);
and U1428 (N_1428,N_358,In_2195);
or U1429 (N_1429,In_132,In_887);
xnor U1430 (N_1430,In_1556,N_113);
nor U1431 (N_1431,In_155,In_243);
nand U1432 (N_1432,N_0,N_477);
nand U1433 (N_1433,In_2076,In_2110);
nor U1434 (N_1434,In_1488,N_962);
xnor U1435 (N_1435,In_1719,In_2146);
nand U1436 (N_1436,In_2590,In_2734);
xnor U1437 (N_1437,N_604,N_788);
nor U1438 (N_1438,N_264,N_954);
or U1439 (N_1439,N_917,In_1619);
and U1440 (N_1440,N_787,N_876);
and U1441 (N_1441,N_26,In_800);
xnor U1442 (N_1442,N_667,N_615);
nor U1443 (N_1443,In_2799,In_845);
or U1444 (N_1444,In_2412,N_687);
or U1445 (N_1445,In_2777,In_2689);
xnor U1446 (N_1446,N_943,In_716);
xnor U1447 (N_1447,N_983,N_716);
xor U1448 (N_1448,In_1809,In_1939);
nor U1449 (N_1449,N_634,In_1600);
nand U1450 (N_1450,N_181,In_2721);
xnor U1451 (N_1451,N_869,In_2486);
and U1452 (N_1452,In_2038,In_379);
nor U1453 (N_1453,In_133,In_553);
xnor U1454 (N_1454,N_126,N_861);
nor U1455 (N_1455,N_156,In_834);
and U1456 (N_1456,N_371,In_2732);
nor U1457 (N_1457,N_967,N_427);
xor U1458 (N_1458,In_2489,In_1779);
or U1459 (N_1459,N_740,N_148);
and U1460 (N_1460,N_640,N_85);
or U1461 (N_1461,In_2087,In_2034);
nand U1462 (N_1462,In_109,In_1581);
xor U1463 (N_1463,In_146,In_2140);
or U1464 (N_1464,In_1772,In_489);
nor U1465 (N_1465,N_925,In_462);
or U1466 (N_1466,In_1451,In_2687);
and U1467 (N_1467,In_466,In_2630);
nor U1468 (N_1468,In_890,In_778);
xnor U1469 (N_1469,N_602,In_1518);
and U1470 (N_1470,In_1699,In_91);
and U1471 (N_1471,In_2774,In_1478);
xnor U1472 (N_1472,In_1229,In_1070);
nor U1473 (N_1473,In_408,In_1765);
and U1474 (N_1474,N_503,In_2230);
nand U1475 (N_1475,N_794,In_2284);
and U1476 (N_1476,In_2703,In_2920);
nor U1477 (N_1477,In_2436,In_1297);
or U1478 (N_1478,In_2337,In_1188);
nor U1479 (N_1479,In_913,N_647);
nor U1480 (N_1480,In_1148,N_660);
nand U1481 (N_1481,In_494,N_410);
and U1482 (N_1482,N_285,N_149);
and U1483 (N_1483,N_305,N_882);
and U1484 (N_1484,N_436,N_111);
nor U1485 (N_1485,In_333,N_78);
and U1486 (N_1486,In_1106,N_772);
xor U1487 (N_1487,N_102,In_2057);
and U1488 (N_1488,In_1725,In_2048);
or U1489 (N_1489,N_490,In_1228);
nor U1490 (N_1490,In_2041,In_1933);
nor U1491 (N_1491,N_49,N_998);
nor U1492 (N_1492,In_1661,In_1102);
and U1493 (N_1493,In_2004,N_934);
xnor U1494 (N_1494,N_46,In_1265);
or U1495 (N_1495,N_896,N_287);
or U1496 (N_1496,In_2965,N_977);
nand U1497 (N_1497,In_541,In_2367);
or U1498 (N_1498,N_262,N_742);
nand U1499 (N_1499,N_108,In_449);
nand U1500 (N_1500,N_1345,N_1451);
nor U1501 (N_1501,In_2335,N_989);
xnor U1502 (N_1502,N_944,N_717);
xnor U1503 (N_1503,In_2755,N_569);
xor U1504 (N_1504,In_2421,N_1182);
nor U1505 (N_1505,N_1226,In_63);
nor U1506 (N_1506,In_2960,In_177);
nand U1507 (N_1507,N_1485,N_832);
xnor U1508 (N_1508,N_80,In_1217);
xor U1509 (N_1509,N_664,N_1018);
nor U1510 (N_1510,N_1391,N_529);
or U1511 (N_1511,N_958,In_1007);
nand U1512 (N_1512,In_568,In_2864);
xnor U1513 (N_1513,N_594,In_1855);
nor U1514 (N_1514,In_1030,N_1279);
nor U1515 (N_1515,In_2439,In_2568);
and U1516 (N_1516,N_588,N_1350);
nand U1517 (N_1517,N_1029,In_2288);
nand U1518 (N_1518,N_1372,N_1435);
or U1519 (N_1519,In_1630,N_850);
xnor U1520 (N_1520,In_1223,N_228);
nor U1521 (N_1521,N_1317,In_743);
or U1522 (N_1522,In_384,In_427);
nor U1523 (N_1523,N_817,N_784);
nand U1524 (N_1524,N_745,In_242);
or U1525 (N_1525,N_939,N_1390);
xnor U1526 (N_1526,N_94,N_1036);
xor U1527 (N_1527,In_2531,In_22);
nand U1528 (N_1528,In_737,In_666);
nand U1529 (N_1529,N_899,In_1842);
or U1530 (N_1530,N_800,In_130);
and U1531 (N_1531,In_678,N_1463);
nand U1532 (N_1532,In_2532,In_1088);
and U1533 (N_1533,N_898,N_597);
nor U1534 (N_1534,N_1076,In_593);
or U1535 (N_1535,N_965,N_306);
or U1536 (N_1536,In_2898,In_383);
or U1537 (N_1537,In_2915,In_1056);
and U1538 (N_1538,N_1312,In_2229);
nand U1539 (N_1539,N_1496,N_1493);
and U1540 (N_1540,In_169,N_1297);
or U1541 (N_1541,N_1311,N_1497);
and U1542 (N_1542,N_186,N_278);
nor U1543 (N_1543,In_672,N_1088);
nand U1544 (N_1544,N_1276,N_891);
nor U1545 (N_1545,In_97,N_1346);
or U1546 (N_1546,N_1404,N_1491);
or U1547 (N_1547,In_2742,N_1498);
and U1548 (N_1548,In_1835,In_2834);
nand U1549 (N_1549,N_1443,In_367);
or U1550 (N_1550,N_1064,N_820);
xor U1551 (N_1551,In_1306,N_1338);
nand U1552 (N_1552,N_1039,In_2869);
and U1553 (N_1553,N_1185,In_2286);
nor U1554 (N_1554,N_777,N_509);
xor U1555 (N_1555,In_2760,N_1189);
and U1556 (N_1556,In_873,In_186);
nand U1557 (N_1557,N_607,N_1045);
nand U1558 (N_1558,N_1173,N_1061);
nand U1559 (N_1559,In_857,In_2329);
nand U1560 (N_1560,N_1403,N_77);
nand U1561 (N_1561,In_862,N_1389);
or U1562 (N_1562,In_2218,N_1465);
nor U1563 (N_1563,In_1668,N_86);
nand U1564 (N_1564,N_1203,N_1104);
nand U1565 (N_1565,In_209,In_344);
nand U1566 (N_1566,In_1359,N_961);
nor U1567 (N_1567,In_252,N_608);
xnor U1568 (N_1568,N_727,N_482);
nand U1569 (N_1569,N_1096,In_1553);
nor U1570 (N_1570,N_1233,N_1117);
nor U1571 (N_1571,N_1100,In_1775);
nor U1572 (N_1572,N_1330,In_1313);
xnor U1573 (N_1573,N_792,In_938);
or U1574 (N_1574,N_1003,N_1377);
or U1575 (N_1575,N_572,N_1097);
or U1576 (N_1576,N_948,In_1138);
nor U1577 (N_1577,N_1375,In_658);
or U1578 (N_1578,N_1286,N_68);
nor U1579 (N_1579,In_650,N_1220);
nand U1580 (N_1580,In_2182,N_23);
xnor U1581 (N_1581,In_633,N_1081);
and U1582 (N_1582,In_4,N_1112);
nor U1583 (N_1583,N_1320,In_2253);
and U1584 (N_1584,N_1211,N_256);
xor U1585 (N_1585,In_2625,In_1935);
xnor U1586 (N_1586,In_590,N_1030);
and U1587 (N_1587,In_2290,In_2434);
and U1588 (N_1588,N_1120,N_1352);
xor U1589 (N_1589,N_1208,In_766);
or U1590 (N_1590,N_1167,In_1973);
nand U1591 (N_1591,N_1401,N_849);
nand U1592 (N_1592,N_198,N_1243);
nand U1593 (N_1593,In_1094,In_1754);
nand U1594 (N_1594,N_1075,In_352);
xor U1595 (N_1595,N_1310,N_1103);
xnor U1596 (N_1596,In_164,N_440);
xnor U1597 (N_1597,N_1424,N_880);
nand U1598 (N_1598,N_764,N_1229);
nand U1599 (N_1599,N_1107,N_744);
xnor U1600 (N_1600,N_1057,N_1138);
nand U1601 (N_1601,N_1209,N_587);
and U1602 (N_1602,In_2051,N_625);
xor U1603 (N_1603,N_431,N_132);
nor U1604 (N_1604,N_1074,N_33);
xnor U1605 (N_1605,In_229,In_2852);
and U1606 (N_1606,In_2,N_1011);
or U1607 (N_1607,N_1188,N_1416);
or U1608 (N_1608,N_1444,In_2716);
xor U1609 (N_1609,N_654,N_887);
and U1610 (N_1610,N_319,N_1034);
nand U1611 (N_1611,N_1300,N_1027);
or U1612 (N_1612,N_712,In_2046);
nand U1613 (N_1613,N_768,N_932);
nand U1614 (N_1614,N_1004,N_190);
nor U1615 (N_1615,N_1197,In_2653);
or U1616 (N_1616,N_1328,N_1281);
or U1617 (N_1617,N_478,In_1730);
or U1618 (N_1618,N_209,N_1452);
nand U1619 (N_1619,N_360,N_1380);
xnor U1620 (N_1620,In_1374,N_114);
nand U1621 (N_1621,In_2115,N_1221);
xnor U1622 (N_1622,N_1130,In_1736);
nand U1623 (N_1623,In_2949,In_483);
or U1624 (N_1624,N_1431,N_1418);
nand U1625 (N_1625,N_239,In_1131);
and U1626 (N_1626,N_534,In_649);
nor U1627 (N_1627,N_902,In_1168);
or U1628 (N_1628,In_2126,N_391);
nor U1629 (N_1629,N_1178,In_2662);
or U1630 (N_1630,In_1354,In_534);
or U1631 (N_1631,N_441,N_1482);
nor U1632 (N_1632,In_1679,In_153);
xor U1633 (N_1633,In_1799,N_1216);
and U1634 (N_1634,In_1231,In_1054);
or U1635 (N_1635,N_508,N_1183);
and U1636 (N_1636,In_313,N_556);
nor U1637 (N_1637,N_1355,N_297);
xnor U1638 (N_1638,N_502,N_1262);
or U1639 (N_1639,N_1318,In_2521);
and U1640 (N_1640,In_1510,N_411);
or U1641 (N_1641,In_2271,In_929);
xnor U1642 (N_1642,N_1324,N_901);
xor U1643 (N_1643,N_626,In_1449);
nand U1644 (N_1644,N_1139,N_1478);
nor U1645 (N_1645,N_1228,N_531);
nand U1646 (N_1646,In_547,In_869);
or U1647 (N_1647,In_1526,N_1070);
and U1648 (N_1648,N_1454,N_91);
nand U1649 (N_1649,In_1732,N_1369);
or U1650 (N_1650,N_535,In_959);
nor U1651 (N_1651,N_334,In_2900);
nor U1652 (N_1652,In_502,N_1149);
and U1653 (N_1653,N_665,In_2113);
nand U1654 (N_1654,In_852,N_1357);
nand U1655 (N_1655,N_1239,N_1231);
nand U1656 (N_1656,In_797,In_2372);
nand U1657 (N_1657,N_945,N_937);
or U1658 (N_1658,N_1164,In_1710);
nor U1659 (N_1659,N_226,N_1381);
xor U1660 (N_1660,N_755,N_1438);
or U1661 (N_1661,N_562,In_2249);
or U1662 (N_1662,In_623,N_893);
or U1663 (N_1663,In_1739,In_978);
xor U1664 (N_1664,N_192,N_139);
xor U1665 (N_1665,N_1062,N_1299);
and U1666 (N_1666,N_649,N_619);
nand U1667 (N_1667,In_2089,N_530);
or U1668 (N_1668,In_2234,In_1073);
nor U1669 (N_1669,N_1193,In_740);
nor U1670 (N_1670,In_2259,N_1123);
or U1671 (N_1671,N_1241,N_1268);
and U1672 (N_1672,N_273,N_914);
and U1673 (N_1673,In_2399,N_1334);
and U1674 (N_1674,N_663,N_1019);
nor U1675 (N_1675,N_1225,In_261);
xor U1676 (N_1676,N_752,In_1333);
or U1677 (N_1677,N_438,N_779);
nand U1678 (N_1678,In_1128,N_1155);
nor U1679 (N_1679,In_123,In_2516);
and U1680 (N_1680,In_482,N_88);
nor U1681 (N_1681,N_1373,In_1941);
or U1682 (N_1682,In_2150,N_699);
or U1683 (N_1683,N_1414,N_1005);
nor U1684 (N_1684,N_451,In_1899);
and U1685 (N_1685,In_1612,In_2240);
and U1686 (N_1686,N_1056,N_706);
or U1687 (N_1687,N_1186,N_818);
nand U1688 (N_1688,In_2612,N_224);
nor U1689 (N_1689,In_1528,N_1336);
xor U1690 (N_1690,In_2448,N_809);
and U1691 (N_1691,In_84,In_635);
nand U1692 (N_1692,N_1473,In_955);
xor U1693 (N_1693,In_516,N_1204);
xnor U1694 (N_1694,In_341,N_568);
nor U1695 (N_1695,N_670,N_267);
nand U1696 (N_1696,N_1432,N_1354);
or U1697 (N_1697,In_1486,In_1366);
and U1698 (N_1698,N_908,N_1235);
xnor U1699 (N_1699,N_1249,In_405);
or U1700 (N_1700,In_406,N_196);
and U1701 (N_1701,In_2366,In_1256);
or U1702 (N_1702,N_1412,N_1456);
or U1703 (N_1703,N_1022,In_888);
or U1704 (N_1704,N_920,In_1621);
nor U1705 (N_1705,In_136,In_2444);
xor U1706 (N_1706,In_1246,N_551);
and U1707 (N_1707,N_263,N_1359);
nor U1708 (N_1708,N_34,N_1240);
and U1709 (N_1709,N_353,N_1158);
nor U1710 (N_1710,In_2973,N_1339);
and U1711 (N_1711,In_1689,In_2857);
and U1712 (N_1712,N_638,N_1032);
nand U1713 (N_1713,N_1447,In_1032);
nor U1714 (N_1714,N_1245,In_1082);
xnor U1715 (N_1715,In_830,N_924);
xor U1716 (N_1716,N_1161,N_1212);
nand U1717 (N_1717,In_2102,In_246);
or U1718 (N_1718,In_751,In_1715);
xor U1719 (N_1719,In_2052,N_1044);
nor U1720 (N_1720,N_446,In_1364);
xnor U1721 (N_1721,N_366,N_878);
nor U1722 (N_1722,In_1399,N_1471);
nor U1723 (N_1723,In_253,N_1398);
xnor U1724 (N_1724,N_947,In_2088);
xor U1725 (N_1725,In_2232,N_748);
xnor U1726 (N_1726,N_1215,N_782);
nand U1727 (N_1727,N_972,N_127);
nor U1728 (N_1728,In_562,N_1199);
xnor U1729 (N_1729,In_2993,In_2295);
xor U1730 (N_1730,N_1295,In_431);
and U1731 (N_1731,N_1335,N_1446);
xnor U1732 (N_1732,N_1265,N_1160);
and U1733 (N_1733,In_103,In_721);
nor U1734 (N_1734,In_2136,N_1433);
and U1735 (N_1735,In_2717,N_824);
and U1736 (N_1736,N_592,In_296);
nand U1737 (N_1737,N_1083,N_1437);
and U1738 (N_1738,In_2464,N_83);
or U1739 (N_1739,In_1531,N_1441);
and U1740 (N_1740,In_185,N_675);
nor U1741 (N_1741,N_513,N_1476);
xnor U1742 (N_1742,N_241,In_26);
and U1743 (N_1743,N_892,N_1127);
xor U1744 (N_1744,N_729,In_2411);
xnor U1745 (N_1745,N_897,N_1344);
or U1746 (N_1746,In_1639,In_335);
xor U1747 (N_1747,In_31,N_1102);
nand U1748 (N_1748,N_1316,N_255);
and U1749 (N_1749,In_2926,In_2062);
xor U1750 (N_1750,N_1309,In_1411);
nor U1751 (N_1751,N_900,In_2543);
nand U1752 (N_1752,N_1059,In_2461);
and U1753 (N_1753,In_2204,In_2542);
xnor U1754 (N_1754,In_1450,N_655);
or U1755 (N_1755,In_1266,N_1133);
nand U1756 (N_1756,N_909,In_51);
xor U1757 (N_1757,N_1322,N_505);
nand U1758 (N_1758,N_375,N_1408);
xor U1759 (N_1759,In_1833,N_1121);
or U1760 (N_1760,N_1230,N_511);
nand U1761 (N_1761,N_1449,In_942);
nor U1762 (N_1762,N_128,N_955);
nand U1763 (N_1763,N_1291,N_1023);
nand U1764 (N_1764,In_2811,N_1095);
and U1765 (N_1765,In_1021,N_1043);
or U1766 (N_1766,In_2070,In_2646);
nand U1767 (N_1767,N_927,N_928);
nor U1768 (N_1768,In_2589,N_54);
or U1769 (N_1769,In_1022,N_709);
nor U1770 (N_1770,N_1210,In_228);
xor U1771 (N_1771,N_866,N_365);
xor U1772 (N_1772,N_1371,In_2787);
nand U1773 (N_1773,N_1079,N_403);
or U1774 (N_1774,N_1293,N_351);
nand U1775 (N_1775,In_2978,In_2228);
xnor U1776 (N_1776,N_1046,N_1082);
and U1777 (N_1777,N_851,N_1395);
nor U1778 (N_1778,N_1470,N_1037);
nand U1779 (N_1779,N_1153,N_1007);
nor U1780 (N_1780,In_600,In_576);
and U1781 (N_1781,In_1987,In_2487);
nand U1782 (N_1782,In_1133,In_1083);
nor U1783 (N_1783,N_500,In_1317);
and U1784 (N_1784,N_833,N_1308);
or U1785 (N_1785,N_233,In_343);
or U1786 (N_1786,In_1014,N_1384);
xor U1787 (N_1787,In_60,In_304);
or U1788 (N_1788,N_215,In_2907);
nand U1789 (N_1789,In_1653,N_363);
nor U1790 (N_1790,In_2994,In_2947);
and U1791 (N_1791,N_1187,N_845);
and U1792 (N_1792,In_2291,In_2634);
nand U1793 (N_1793,N_980,In_2545);
nand U1794 (N_1794,N_894,In_2968);
nand U1795 (N_1795,In_1743,In_573);
nand U1796 (N_1796,N_1387,N_172);
nand U1797 (N_1797,N_1172,N_858);
nor U1798 (N_1798,N_1434,N_736);
xor U1799 (N_1799,In_2398,In_698);
and U1800 (N_1800,N_344,N_1129);
nand U1801 (N_1801,In_2467,N_672);
xnor U1802 (N_1802,N_1148,N_710);
and U1803 (N_1803,N_1442,N_848);
nor U1804 (N_1804,N_357,N_566);
and U1805 (N_1805,N_1154,N_1207);
nand U1806 (N_1806,N_552,In_2023);
nand U1807 (N_1807,N_1090,N_1492);
xnor U1808 (N_1808,N_1157,In_108);
nand U1809 (N_1809,N_1073,N_1382);
xor U1810 (N_1810,In_2648,N_1165);
or U1811 (N_1811,In_2585,N_1420);
nand U1812 (N_1812,In_1197,N_1001);
nand U1813 (N_1813,N_1460,N_700);
or U1814 (N_1814,N_434,N_519);
nand U1815 (N_1815,N_1191,N_1329);
xnor U1816 (N_1816,In_958,In_694);
nand U1817 (N_1817,In_1232,In_1116);
nand U1818 (N_1818,N_765,N_1054);
nand U1819 (N_1819,In_77,N_271);
and U1820 (N_1820,N_1307,N_276);
nor U1821 (N_1821,In_1525,In_1823);
and U1822 (N_1822,N_1026,N_1255);
and U1823 (N_1823,N_201,In_2934);
nand U1824 (N_1824,In_2147,N_1325);
and U1825 (N_1825,In_1340,N_1489);
nand U1826 (N_1826,N_1248,N_1232);
nor U1827 (N_1827,N_528,In_870);
nand U1828 (N_1828,N_378,N_1440);
nor U1829 (N_1829,In_2935,In_207);
nor U1830 (N_1830,In_1866,N_1010);
or U1831 (N_1831,N_1136,N_1425);
xor U1832 (N_1832,In_791,N_1163);
and U1833 (N_1833,In_2681,In_375);
xnor U1834 (N_1834,In_984,N_889);
xnor U1835 (N_1835,In_2525,In_2049);
nand U1836 (N_1836,N_1124,In_851);
nor U1837 (N_1837,N_493,N_766);
nor U1838 (N_1838,N_886,N_1128);
or U1839 (N_1839,In_1704,N_470);
and U1840 (N_1840,N_1388,N_1315);
nand U1841 (N_1841,N_976,In_2638);
xor U1842 (N_1842,In_52,N_97);
nor U1843 (N_1843,In_1956,N_133);
nand U1844 (N_1844,N_855,N_372);
and U1845 (N_1845,In_944,N_1490);
xor U1846 (N_1846,N_1303,N_1461);
nor U1847 (N_1847,In_1349,In_2866);
nor U1848 (N_1848,N_455,In_1894);
nand U1849 (N_1849,In_300,In_1226);
or U1850 (N_1850,N_1246,In_426);
xor U1851 (N_1851,N_230,N_741);
nand U1852 (N_1852,In_1822,In_2622);
xnor U1853 (N_1853,N_1277,In_2970);
or U1854 (N_1854,N_1450,In_2391);
and U1855 (N_1855,In_2706,In_2355);
nor U1856 (N_1856,N_96,N_1439);
or U1857 (N_1857,N_575,In_2071);
or U1858 (N_1858,N_1298,N_1296);
nor U1859 (N_1859,N_1427,In_1643);
nand U1860 (N_1860,In_1949,In_310);
or U1861 (N_1861,N_666,N_195);
and U1862 (N_1862,In_495,In_2221);
nand U1863 (N_1863,In_2491,N_846);
nor U1864 (N_1864,N_32,In_216);
and U1865 (N_1865,In_319,N_1110);
and U1866 (N_1866,N_251,In_2128);
or U1867 (N_1867,N_931,In_875);
or U1868 (N_1868,N_1122,N_806);
nand U1869 (N_1869,In_2396,N_1411);
and U1870 (N_1870,N_842,N_1134);
or U1871 (N_1871,N_368,N_1253);
or U1872 (N_1872,In_1031,N_1234);
and U1873 (N_1873,N_1143,N_1237);
nand U1874 (N_1874,In_1135,N_1258);
or U1875 (N_1875,In_2029,N_1275);
or U1876 (N_1876,N_697,N_1114);
nor U1877 (N_1877,N_110,In_926);
nor U1878 (N_1878,In_2544,N_1015);
or U1879 (N_1879,In_804,In_2884);
nand U1880 (N_1880,In_993,In_2413);
or U1881 (N_1881,N_1284,N_606);
xnor U1882 (N_1882,N_1101,In_96);
and U1883 (N_1883,N_1343,N_150);
nand U1884 (N_1884,N_774,N_288);
xor U1885 (N_1885,N_730,N_997);
and U1886 (N_1886,N_313,In_1578);
and U1887 (N_1887,In_1462,N_1337);
xor U1888 (N_1888,N_1483,N_1455);
nor U1889 (N_1889,In_763,N_546);
or U1890 (N_1890,In_1632,In_21);
and U1891 (N_1891,In_2465,N_867);
nand U1892 (N_1892,N_460,N_1351);
and U1893 (N_1893,N_1135,N_480);
xnor U1894 (N_1894,N_252,In_1170);
or U1895 (N_1895,N_1406,N_1145);
nor U1896 (N_1896,N_916,N_1067);
nor U1897 (N_1897,N_1333,N_1190);
and U1898 (N_1898,N_844,N_1181);
xnor U1899 (N_1899,N_1205,In_891);
nand U1900 (N_1900,In_2578,N_704);
or U1901 (N_1901,In_946,In_2406);
nand U1902 (N_1902,In_1177,In_2535);
nor U1903 (N_1903,N_668,N_1374);
and U1904 (N_1904,In_923,In_2854);
nand U1905 (N_1905,In_429,N_510);
xor U1906 (N_1906,In_66,In_2955);
xnor U1907 (N_1907,N_1040,N_66);
xnor U1908 (N_1908,N_1282,N_1111);
or U1909 (N_1909,In_2245,In_1706);
xnor U1910 (N_1910,N_1144,N_1242);
nand U1911 (N_1911,In_2139,In_437);
and U1912 (N_1912,N_692,N_1131);
nor U1913 (N_1913,N_1472,In_1212);
or U1914 (N_1914,N_694,N_1094);
xor U1915 (N_1915,In_2647,N_1146);
xor U1916 (N_1916,In_127,In_921);
xnor U1917 (N_1917,In_257,In_12);
and U1918 (N_1918,In_1189,N_1014);
nor U1919 (N_1919,In_985,In_992);
xnor U1920 (N_1920,N_974,N_1370);
nor U1921 (N_1921,In_361,N_571);
nand U1922 (N_1922,In_1373,In_359);
nor U1923 (N_1923,In_1362,In_2595);
nor U1924 (N_1924,N_1272,In_463);
nor U1925 (N_1925,In_2957,In_1818);
xnor U1926 (N_1926,In_2951,In_1920);
nor U1927 (N_1927,N_1244,N_1459);
nand U1928 (N_1928,N_1341,N_1016);
nor U1929 (N_1929,In_2575,N_450);
nand U1930 (N_1930,N_1421,In_2077);
nand U1931 (N_1931,N_1376,N_1407);
nor U1932 (N_1932,N_653,N_821);
nor U1933 (N_1933,N_1273,N_1031);
nor U1934 (N_1934,N_281,N_1012);
nor U1935 (N_1935,N_1367,N_938);
nor U1936 (N_1936,N_1072,In_1412);
nand U1937 (N_1937,In_321,In_2682);
or U1938 (N_1938,N_1323,In_2153);
xnor U1939 (N_1939,In_908,N_1361);
and U1940 (N_1940,N_453,In_2713);
nor U1941 (N_1941,N_1468,N_81);
nand U1942 (N_1942,In_2157,In_948);
nor U1943 (N_1943,N_662,N_696);
xor U1944 (N_1944,N_1084,In_1838);
or U1945 (N_1945,N_576,In_2707);
nor U1946 (N_1946,In_2135,In_286);
or U1947 (N_1947,N_1171,In_1220);
nor U1948 (N_1948,In_2604,N_1176);
xnor U1949 (N_1949,N_1466,N_786);
or U1950 (N_1950,N_815,N_757);
and U1951 (N_1951,N_1383,N_1214);
nor U1952 (N_1952,N_910,N_549);
and U1953 (N_1953,N_678,N_1348);
nor U1954 (N_1954,In_2179,N_632);
xor U1955 (N_1955,In_1561,In_2723);
nor U1956 (N_1956,In_1911,In_2597);
xnor U1957 (N_1957,N_731,N_1417);
or U1958 (N_1958,N_834,In_1020);
xnor U1959 (N_1959,N_39,N_822);
nor U1960 (N_1960,In_2675,N_1227);
xor U1961 (N_1961,N_1340,N_941);
nand U1962 (N_1962,N_117,N_1342);
nor U1963 (N_1963,In_1656,N_1274);
nand U1964 (N_1964,In_2778,N_22);
nand U1965 (N_1965,N_999,N_1025);
nand U1966 (N_1966,N_269,In_2217);
or U1967 (N_1967,In_2966,N_1224);
nand U1968 (N_1968,N_680,N_1270);
or U1969 (N_1969,N_728,In_974);
or U1970 (N_1970,N_1050,N_1166);
and U1971 (N_1971,N_1195,N_1147);
and U1972 (N_1972,N_836,N_760);
nor U1973 (N_1973,In_1090,In_1346);
and U1974 (N_1974,N_1252,N_864);
and U1975 (N_1975,N_544,In_2309);
xor U1976 (N_1976,N_254,N_1419);
or U1977 (N_1977,In_27,N_1013);
and U1978 (N_1978,In_2109,In_1081);
nand U1979 (N_1979,N_499,N_1379);
and U1980 (N_1980,N_819,N_1151);
and U1981 (N_1981,N_1364,N_734);
xnor U1982 (N_1982,In_2127,N_1487);
nand U1983 (N_1983,N_888,N_629);
xnor U1984 (N_1984,N_1126,In_2331);
xnor U1985 (N_1985,N_1319,In_912);
and U1986 (N_1986,N_1287,In_994);
and U1987 (N_1987,N_1202,N_1467);
xor U1988 (N_1988,N_1099,N_259);
and U1989 (N_1989,N_416,N_223);
nand U1990 (N_1990,In_765,N_343);
xor U1991 (N_1991,In_1747,In_2501);
nand U1992 (N_1992,N_1453,N_517);
nand U1993 (N_1993,N_1238,In_928);
nor U1994 (N_1994,In_2748,N_643);
xnor U1995 (N_1995,N_364,In_1869);
and U1996 (N_1996,N_1141,In_1017);
xor U1997 (N_1997,N_1077,In_86);
or U1998 (N_1998,In_664,In_725);
nor U1999 (N_1999,In_2225,N_1150);
or U2000 (N_2000,N_1567,N_1428);
xnor U2001 (N_2001,In_679,N_801);
nand U2002 (N_2002,N_837,N_1709);
xnor U2003 (N_2003,N_1142,In_1159);
and U2004 (N_2004,In_6,N_1469);
and U2005 (N_2005,N_1041,In_2956);
nor U2006 (N_2006,N_1569,N_1501);
and U2007 (N_2007,N_1448,N_1711);
nand U2008 (N_2008,N_1169,N_1621);
nand U2009 (N_2009,N_1581,In_2321);
nor U2010 (N_2010,In_2159,N_1716);
or U2011 (N_2011,N_1793,N_877);
xor U2012 (N_2012,N_1500,N_1905);
xor U2013 (N_2013,In_2001,N_1691);
xnor U2014 (N_2014,N_1681,N_1289);
nor U2015 (N_2015,N_610,In_1249);
nor U2016 (N_2016,N_1257,N_299);
nor U2017 (N_2017,N_1584,N_1565);
xnor U2018 (N_2018,N_1516,N_1570);
and U2019 (N_2019,N_1977,N_1002);
nand U2020 (N_2020,N_1881,In_1200);
xor U2021 (N_2021,In_37,N_1116);
and U2022 (N_2022,N_93,N_1800);
nand U2023 (N_2023,In_865,In_1552);
xnor U2024 (N_2024,N_1159,In_2009);
or U2025 (N_2025,In_2830,N_1708);
or U2026 (N_2026,N_1599,N_1888);
xnor U2027 (N_2027,In_233,N_1869);
nand U2028 (N_2028,N_839,N_92);
nor U2029 (N_2029,In_1253,N_1766);
xnor U2030 (N_2030,N_1087,N_1937);
xnor U2031 (N_2031,N_936,N_1738);
and U2032 (N_2032,N_1995,N_1086);
nor U2033 (N_2033,N_1368,N_1600);
nand U2034 (N_2034,N_1543,N_1280);
nand U2035 (N_2035,N_1925,N_373);
and U2036 (N_2036,In_1311,N_1589);
xor U2037 (N_2037,N_1770,N_1582);
xor U2038 (N_2038,N_1620,N_1528);
nand U2039 (N_2039,N_176,N_1609);
nor U2040 (N_2040,N_1967,N_1579);
or U2041 (N_2041,N_1829,N_1093);
nor U2042 (N_2042,In_2667,N_188);
or U2043 (N_2043,N_813,N_863);
xnor U2044 (N_2044,N_711,N_1744);
nor U2045 (N_2045,N_293,N_1758);
xor U2046 (N_2046,N_1962,N_1887);
and U2047 (N_2047,N_1657,N_1540);
nor U2048 (N_2048,N_1771,N_1849);
xor U2049 (N_2049,N_1729,N_1658);
or U2050 (N_2050,N_857,In_2856);
and U2051 (N_2051,N_1784,N_1611);
xor U2052 (N_2052,N_1921,N_1961);
xnor U2053 (N_2053,In_1684,N_1590);
xor U2054 (N_2054,N_1913,N_648);
nor U2055 (N_2055,N_1689,N_1653);
or U2056 (N_2056,N_1606,N_951);
nor U2057 (N_2057,N_1200,N_1877);
or U2058 (N_2058,N_1959,N_1973);
xor U2059 (N_2059,N_1347,In_256);
or U2060 (N_2060,In_514,N_1436);
or U2061 (N_2061,N_797,N_1402);
nor U2062 (N_2062,N_1867,N_1017);
or U2063 (N_2063,N_1818,N_1256);
nor U2064 (N_2064,N_1480,N_1477);
nor U2065 (N_2065,N_1494,N_1566);
or U2066 (N_2066,N_829,N_491);
xnor U2067 (N_2067,N_1727,N_1267);
and U2068 (N_2068,In_2763,In_112);
xnor U2069 (N_2069,N_1878,N_1719);
nand U2070 (N_2070,N_1587,N_1445);
or U2071 (N_2071,N_1794,In_1248);
nand U2072 (N_2072,N_1551,In_1301);
or U2073 (N_2073,In_1080,N_1759);
and U2074 (N_2074,N_1971,In_113);
xnor U2075 (N_2075,N_1356,N_739);
xnor U2076 (N_2076,N_1263,N_1720);
or U2077 (N_2077,N_1944,N_1986);
or U2078 (N_2078,N_152,N_1692);
and U2079 (N_2079,N_1386,N_1332);
or U2080 (N_2080,N_1882,N_1515);
and U2081 (N_2081,N_1213,In_55);
xor U2082 (N_2082,N_504,N_1614);
xor U2083 (N_2083,N_1108,N_1697);
xor U2084 (N_2084,N_1085,N_1980);
xor U2085 (N_2085,N_445,N_1671);
and U2086 (N_2086,In_1466,In_1361);
nor U2087 (N_2087,N_1290,N_1885);
or U2088 (N_2088,In_1473,N_1841);
nand U2089 (N_2089,N_1000,N_1791);
nand U2090 (N_2090,N_1278,N_1777);
or U2091 (N_2091,N_1764,N_963);
and U2092 (N_2092,N_1628,N_229);
nor U2093 (N_2093,N_1895,N_1633);
and U2094 (N_2094,N_1942,In_2306);
xor U2095 (N_2095,N_1575,N_1647);
nor U2096 (N_2096,N_1321,In_1195);
or U2097 (N_2097,N_935,N_1904);
and U2098 (N_2098,N_1604,N_380);
and U2099 (N_2099,N_1908,N_1071);
or U2100 (N_2100,N_762,In_2846);
nor U2101 (N_2101,N_1047,N_1999);
nand U2102 (N_2102,N_1285,N_1137);
and U2103 (N_2103,N_1920,N_99);
xnor U2104 (N_2104,N_1786,In_2354);
or U2105 (N_2105,N_1781,N_1871);
nor U2106 (N_2106,N_118,N_1850);
nor U2107 (N_2107,N_1399,N_1513);
nand U2108 (N_2108,In_1039,In_2121);
nand U2109 (N_2109,N_1636,In_2871);
and U2110 (N_2110,N_868,N_1838);
and U2111 (N_2111,N_691,N_596);
and U2112 (N_2112,N_413,N_1748);
nand U2113 (N_2113,N_785,N_1648);
xnor U2114 (N_2114,N_1851,N_1876);
and U2115 (N_2115,N_679,In_1515);
and U2116 (N_2116,N_1559,N_1360);
nand U2117 (N_2117,N_1741,N_1900);
nor U2118 (N_2118,N_1933,N_1723);
nor U2119 (N_2119,In_552,In_1737);
and U2120 (N_2120,N_1747,N_1909);
nand U2121 (N_2121,In_197,In_2762);
xnor U2122 (N_2122,N_1302,N_1832);
or U2123 (N_2123,N_1132,N_432);
nand U2124 (N_2124,N_1612,N_1966);
nand U2125 (N_2125,N_332,N_1254);
or U2126 (N_2126,N_1065,N_1778);
xnor U2127 (N_2127,N_1993,N_1946);
xor U2128 (N_2128,In_1239,N_1283);
nor U2129 (N_2129,N_1522,In_1134);
and U2130 (N_2130,N_521,In_1352);
or U2131 (N_2131,N_1737,In_129);
and U2132 (N_2132,In_2258,N_1140);
or U2133 (N_2133,N_1823,N_1066);
and U2134 (N_2134,N_1969,N_1842);
xnor U2135 (N_2135,N_1665,In_1574);
nor U2136 (N_2136,N_1929,N_1819);
nand U2137 (N_2137,N_767,N_1988);
nor U2138 (N_2138,In_42,N_1734);
xor U2139 (N_2139,N_1886,In_1430);
nor U2140 (N_2140,N_669,N_835);
or U2141 (N_2141,N_1544,N_1830);
nor U2142 (N_2142,N_1479,N_1826);
or U2143 (N_2143,N_1860,N_1409);
and U2144 (N_2144,N_1813,N_1632);
nand U2145 (N_2145,N_1713,N_1413);
nor U2146 (N_2146,N_651,N_1694);
xnor U2147 (N_2147,In_983,N_825);
or U2148 (N_2148,N_1836,N_1080);
nor U2149 (N_2149,N_1520,N_1827);
or U2150 (N_2150,N_1911,In_1995);
and U2151 (N_2151,N_1736,N_1564);
nand U2152 (N_2152,N_1898,In_675);
or U2153 (N_2153,N_1392,In_1244);
nor U2154 (N_2154,In_1697,N_1703);
nor U2155 (N_2155,N_1058,N_1264);
nand U2156 (N_2156,In_2091,N_1809);
nor U2157 (N_2157,N_1288,N_1902);
and U2158 (N_2158,N_1853,N_1617);
xnor U2159 (N_2159,N_1684,N_1638);
and U2160 (N_2160,N_1679,N_1530);
nor U2161 (N_2161,N_1677,N_1523);
nand U2162 (N_2162,In_1756,N_120);
nand U2163 (N_2163,N_1817,In_188);
and U2164 (N_2164,In_1477,N_775);
nor U2165 (N_2165,N_1812,N_1998);
nor U2166 (N_2166,N_266,N_1052);
xnor U2167 (N_2167,N_1981,In_1871);
and U2168 (N_2168,In_2322,N_1847);
nand U2169 (N_2169,N_1735,N_859);
nand U2170 (N_2170,In_1315,In_2506);
xor U2171 (N_2171,N_1746,N_1349);
or U2172 (N_2172,N_1558,N_1538);
and U2173 (N_2173,N_1603,N_1915);
nand U2174 (N_2174,N_1894,N_1542);
nand U2175 (N_2175,N_1688,N_1765);
and U2176 (N_2176,N_1624,In_2969);
xor U2177 (N_2177,N_1313,N_758);
nand U2178 (N_2178,N_1979,N_1639);
xnor U2179 (N_2179,N_1118,N_1685);
nand U2180 (N_2180,N_1327,N_1640);
xnor U2181 (N_2181,N_1822,In_812);
or U2182 (N_2182,N_1511,In_1783);
xnor U2183 (N_2183,In_2629,N_559);
and U2184 (N_2184,N_1752,N_1659);
or U2185 (N_2185,N_1662,N_1702);
nand U2186 (N_2186,In_1951,N_921);
xnor U2187 (N_2187,In_0,In_2573);
nor U2188 (N_2188,N_540,N_1660);
xor U2189 (N_2189,N_1548,N_1301);
and U2190 (N_2190,N_11,N_1634);
nor U2191 (N_2191,In_835,N_1803);
and U2192 (N_2192,In_2551,N_1755);
and U2193 (N_2193,N_1619,N_1839);
xnor U2194 (N_2194,N_1588,N_1583);
nand U2195 (N_2195,N_1970,N_1577);
xor U2196 (N_2196,N_1423,N_1524);
and U2197 (N_2197,N_996,N_1512);
xor U2198 (N_2198,N_1562,N_1947);
xnor U2199 (N_2199,N_1712,N_1721);
and U2200 (N_2200,N_1571,N_940);
xor U2201 (N_2201,N_1831,In_2282);
or U2202 (N_2202,In_116,N_1932);
or U2203 (N_2203,In_2205,N_1563);
or U2204 (N_2204,In_503,N_1535);
and U2205 (N_2205,N_1761,N_1623);
and U2206 (N_2206,N_1678,N_1378);
xnor U2207 (N_2207,In_2912,N_1954);
or U2208 (N_2208,N_1919,In_1497);
nor U2209 (N_2209,In_987,In_2193);
nand U2210 (N_2210,N_1928,N_973);
xnor U2211 (N_2211,N_1177,In_174);
nor U2212 (N_2212,In_276,In_1677);
and U2213 (N_2213,N_1218,N_1890);
nor U2214 (N_2214,In_2079,N_1506);
nor U2215 (N_2215,In_897,N_1796);
or U2216 (N_2216,In_2269,N_1795);
and U2217 (N_2217,In_798,N_1613);
and U2218 (N_2218,N_1618,N_1314);
nor U2219 (N_2219,N_1458,In_2226);
nor U2220 (N_2220,In_1874,In_670);
xnor U2221 (N_2221,N_1602,N_1762);
nor U2222 (N_2222,N_1598,N_1695);
xor U2223 (N_2223,N_507,N_1907);
xnor U2224 (N_2224,N_1811,N_1106);
xor U2225 (N_2225,N_1666,In_2059);
nor U2226 (N_2226,N_661,N_1474);
or U2227 (N_2227,In_755,N_1724);
nand U2228 (N_2228,N_1410,N_1955);
nor U2229 (N_2229,N_1607,N_1576);
and U2230 (N_2230,N_1763,N_1769);
nand U2231 (N_2231,N_1514,N_1682);
xnor U2232 (N_2232,N_890,In_1282);
or U2233 (N_2233,N_1782,N_628);
nand U2234 (N_2234,N_686,In_696);
xor U2235 (N_2235,In_1952,N_1430);
xor U2236 (N_2236,N_1834,N_791);
and U2237 (N_2237,N_304,N_339);
xor U2238 (N_2238,N_1787,N_1910);
nand U2239 (N_2239,N_1663,N_296);
or U2240 (N_2240,N_1864,N_1845);
nand U2241 (N_2241,N_1305,In_90);
nand U2242 (N_2242,N_1875,N_1858);
nand U2243 (N_2243,N_1294,N_1554);
xor U2244 (N_2244,N_1749,N_1024);
or U2245 (N_2245,N_1917,N_1457);
nand U2246 (N_2246,N_1536,N_1630);
nand U2247 (N_2247,N_1790,N_1785);
nand U2248 (N_2248,N_703,N_1651);
xor U2249 (N_2249,N_1884,N_1978);
nor U2250 (N_2250,N_1247,N_1363);
and U2251 (N_2251,In_2060,N_1856);
xor U2252 (N_2252,In_433,N_1510);
xor U2253 (N_2253,N_970,N_1557);
nand U2254 (N_2254,N_1989,N_1518);
nand U2255 (N_2255,N_1595,In_733);
xor U2256 (N_2256,In_1242,N_1306);
nand U2257 (N_2257,N_1008,N_1396);
and U2258 (N_2258,N_1555,N_1053);
xnor U2259 (N_2259,N_1531,N_1868);
xor U2260 (N_2260,In_2251,N_1006);
xnor U2261 (N_2261,In_2972,N_1292);
nor U2262 (N_2262,N_1550,N_1901);
and U2263 (N_2263,N_1503,N_1714);
nor U2264 (N_2264,N_1109,In_771);
or U2265 (N_2265,N_1174,N_826);
xnor U2266 (N_2266,N_1394,In_337);
nand U2267 (N_2267,N_1808,N_125);
nand U2268 (N_2268,N_1400,N_1028);
xor U2269 (N_2269,N_721,N_1561);
nor U2270 (N_2270,N_1960,In_545);
nand U2271 (N_2271,N_946,N_1951);
nor U2272 (N_2272,N_1990,In_61);
nor U2273 (N_2273,N_1366,N_1192);
xor U2274 (N_2274,N_1726,N_1956);
and U2275 (N_2275,N_1170,N_613);
xnor U2276 (N_2276,N_1553,N_1991);
nor U2277 (N_2277,In_2770,In_2611);
xor U2278 (N_2278,In_1068,N_966);
xor U2279 (N_2279,N_1585,N_1475);
nor U2280 (N_2280,N_533,N_1821);
and U2281 (N_2281,In_956,N_1063);
nand U2282 (N_2282,N_1038,N_1405);
or U2283 (N_2283,N_1362,N_1502);
xnor U2284 (N_2284,N_1964,N_1162);
nor U2285 (N_2285,In_1419,N_1304);
or U2286 (N_2286,N_1656,N_1673);
and U2287 (N_2287,In_2991,N_1916);
or U2288 (N_2288,N_1655,N_1680);
nor U2289 (N_2289,In_267,N_1779);
nor U2290 (N_2290,In_1379,N_1353);
and U2291 (N_2291,In_2485,N_1975);
xnor U2292 (N_2292,N_1635,N_1223);
xnor U2293 (N_2293,N_1649,N_1260);
and U2294 (N_2294,N_1021,N_1669);
and U2295 (N_2295,N_1499,N_1848);
nand U2296 (N_2296,N_1664,N_1397);
nor U2297 (N_2297,N_1717,N_1814);
or U2298 (N_2298,N_1594,N_1873);
nand U2299 (N_2299,N_1650,N_1180);
or U2300 (N_2300,N_1840,N_153);
or U2301 (N_2301,N_1945,N_1976);
or U2302 (N_2302,N_1125,N_1707);
xor U2303 (N_2303,N_1844,N_1773);
or U2304 (N_2304,N_1984,In_461);
nand U2305 (N_2305,N_1519,N_1206);
nand U2306 (N_2306,N_959,N_749);
xnor U2307 (N_2307,N_1393,N_1760);
nand U2308 (N_2308,N_1698,N_1622);
or U2309 (N_2309,In_2961,N_340);
nor U2310 (N_2310,In_2988,N_723);
or U2311 (N_2311,N_1119,N_1201);
xor U2312 (N_2312,N_1722,N_1105);
or U2313 (N_2313,N_1532,N_1488);
nand U2314 (N_2314,In_1302,N_1539);
and U2315 (N_2315,N_1217,N_1415);
nand U2316 (N_2316,In_1125,N_1941);
xnor U2317 (N_2317,In_2594,N_1326);
and U2318 (N_2318,N_1892,N_1667);
nor U2319 (N_2319,N_1175,In_892);
nor U2320 (N_2320,N_1939,N_1710);
nand U2321 (N_2321,N_1802,N_1641);
xnor U2322 (N_2322,N_1965,In_807);
nor U2323 (N_2323,N_1742,N_1997);
nand U2324 (N_2324,In_498,N_1776);
nor U2325 (N_2325,N_1699,N_1753);
and U2326 (N_2326,N_1820,N_1940);
or U2327 (N_2327,In_975,N_553);
nand U2328 (N_2328,N_1597,N_1730);
or U2329 (N_2329,N_1807,N_622);
and U2330 (N_2330,In_2656,In_1910);
nor U2331 (N_2331,N_1385,In_30);
nand U2332 (N_2332,N_595,N_1568);
or U2333 (N_2333,N_1271,In_2602);
nand U2334 (N_2334,In_963,N_1768);
nor U2335 (N_2335,N_624,In_1647);
or U2336 (N_2336,N_1504,N_1985);
nor U2337 (N_2337,N_1092,In_2591);
or U2338 (N_2338,N_1705,In_2876);
nor U2339 (N_2339,In_1635,N_1893);
or U2340 (N_2340,N_1732,In_2311);
or U2341 (N_2341,N_243,N_1912);
xnor U2342 (N_2342,N_1852,N_1687);
nand U2343 (N_2343,N_1987,N_1556);
nor U2344 (N_2344,N_1870,In_1390);
nand U2345 (N_2345,In_320,N_988);
nand U2346 (N_2346,N_1676,N_554);
and U2347 (N_2347,N_1331,N_260);
xnor U2348 (N_2348,N_991,N_1484);
xnor U2349 (N_2349,N_601,N_1690);
nor U2350 (N_2350,N_1509,In_1196);
and U2351 (N_2351,N_714,N_1931);
or U2352 (N_2352,N_1042,N_1464);
nand U2353 (N_2353,In_2325,N_1992);
and U2354 (N_2354,In_1336,N_870);
and U2355 (N_2355,In_700,In_1593);
nor U2356 (N_2356,N_1806,N_639);
nand U2357 (N_2357,In_210,In_1221);
xor U2358 (N_2358,N_617,N_564);
nand U2359 (N_2359,In_338,N_359);
nand U2360 (N_2360,N_1646,N_1683);
xnor U2361 (N_2361,N_853,In_2747);
or U2362 (N_2362,In_2705,N_1792);
nand U2363 (N_2363,N_1843,N_1728);
and U2364 (N_2364,N_1596,In_87);
and U2365 (N_2365,N_1069,N_1872);
and U2366 (N_2366,N_1857,In_1211);
nand U2367 (N_2367,N_1549,In_949);
or U2368 (N_2368,N_1194,N_589);
nor U2369 (N_2369,N_1529,N_1974);
or U2370 (N_2370,N_1783,In_414);
xnor U2371 (N_2371,In_1158,In_1711);
nor U2372 (N_2372,N_1943,In_583);
xnor U2373 (N_2373,N_1810,N_1654);
nor U2374 (N_2374,In_1883,N_1527);
nand U2375 (N_2375,N_1772,N_1743);
or U2376 (N_2376,N_1963,N_1804);
and U2377 (N_2377,N_1780,N_1615);
and U2378 (N_2378,N_1828,In_1721);
or U2379 (N_2379,N_1914,N_1824);
nand U2380 (N_2380,N_1700,N_773);
xnor U2381 (N_2381,N_1219,N_1222);
and U2382 (N_2382,N_685,N_1846);
nand U2383 (N_2383,N_1547,In_2756);
or U2384 (N_2384,N_798,N_1899);
xor U2385 (N_2385,N_1938,N_1574);
or U2386 (N_2386,N_1580,N_1068);
nor U2387 (N_2387,In_389,N_1865);
and U2388 (N_2388,N_1521,N_1156);
nor U2389 (N_2389,N_1629,N_1115);
nand U2390 (N_2390,N_1896,N_338);
or U2391 (N_2391,N_657,In_2005);
or U2392 (N_2392,N_1091,N_61);
or U2393 (N_2393,N_1601,N_1674);
xor U2394 (N_2394,N_1983,N_1798);
nand U2395 (N_2395,N_1541,N_1879);
xnor U2396 (N_2396,N_1505,N_1113);
and U2397 (N_2397,N_1948,N_979);
or U2398 (N_2398,N_1701,N_1009);
and U2399 (N_2399,N_1429,In_724);
nor U2400 (N_2400,N_1934,N_1586);
nand U2401 (N_2401,N_1731,N_682);
nor U2402 (N_2402,N_1740,N_1179);
or U2403 (N_2403,N_1365,N_1048);
xnor U2404 (N_2404,N_1251,In_380);
and U2405 (N_2405,N_1837,N_1266);
and U2406 (N_2406,N_718,N_1950);
and U2407 (N_2407,In_566,N_1526);
nand U2408 (N_2408,N_1924,N_1686);
or U2409 (N_2409,N_1261,N_1751);
nor U2410 (N_2410,N_1693,N_1644);
xor U2411 (N_2411,N_1426,In_1465);
and U2412 (N_2412,N_1051,In_2927);
or U2413 (N_2413,N_393,In_1493);
nand U2414 (N_2414,In_40,N_1754);
and U2415 (N_2415,N_1035,N_1815);
nor U2416 (N_2416,In_1548,N_146);
or U2417 (N_2417,N_1996,N_1060);
or U2418 (N_2418,In_2964,N_1715);
and U2419 (N_2419,N_1767,N_1952);
nor U2420 (N_2420,In_1543,N_1098);
or U2421 (N_2421,N_811,N_1578);
and U2422 (N_2422,N_1198,N_573);
nor U2423 (N_2423,N_1855,N_1706);
nor U2424 (N_2424,N_1704,In_1598);
nand U2425 (N_2425,N_1805,N_1049);
xor U2426 (N_2426,In_17,N_1507);
or U2427 (N_2427,In_2299,N_673);
or U2428 (N_2428,N_1801,N_1835);
or U2429 (N_2429,In_2692,N_1797);
nor U2430 (N_2430,N_1642,N_1422);
xor U2431 (N_2431,N_1923,In_2782);
nor U2432 (N_2432,N_1668,N_1670);
xnor U2433 (N_2433,N_621,N_1196);
and U2434 (N_2434,N_1866,N_1953);
nor U2435 (N_2435,N_1625,N_1982);
or U2436 (N_2436,In_390,N_1926);
or U2437 (N_2437,N_1891,N_1750);
and U2438 (N_2438,N_1572,N_1525);
and U2439 (N_2439,N_733,N_1994);
nor U2440 (N_2440,N_1168,N_1799);
nand U2441 (N_2441,N_1922,In_1648);
and U2442 (N_2442,N_1462,N_1152);
nand U2443 (N_2443,N_1906,N_1560);
and U2444 (N_2444,N_582,N_1631);
nand U2445 (N_2445,N_1927,N_74);
nor U2446 (N_2446,N_1184,In_981);
and U2447 (N_2447,N_1774,In_824);
xor U2448 (N_2448,In_867,N_1889);
nor U2449 (N_2449,N_1935,N_1626);
and U2450 (N_2450,N_1481,N_1903);
or U2451 (N_2451,N_1739,N_1972);
xnor U2452 (N_2452,N_1645,N_1637);
nor U2453 (N_2453,N_1958,N_73);
or U2454 (N_2454,N_1591,N_1546);
nand U2455 (N_2455,N_1537,N_1863);
or U2456 (N_2456,In_533,N_1816);
xnor U2457 (N_2457,N_1517,N_1957);
nor U2458 (N_2458,N_1592,N_1675);
and U2459 (N_2459,N_1775,N_1236);
and U2460 (N_2460,N_968,N_1718);
or U2461 (N_2461,N_1269,In_1296);
nor U2462 (N_2462,N_1696,N_1949);
and U2463 (N_2463,N_1627,In_554);
and U2464 (N_2464,In_2806,N_1862);
nand U2465 (N_2465,N_1250,N_1573);
nand U2466 (N_2466,N_1608,N_1883);
nand U2467 (N_2467,N_1508,In_1700);
xnor U2468 (N_2468,N_1918,In_641);
nor U2469 (N_2469,In_578,In_1967);
or U2470 (N_2470,N_1930,In_2645);
nor U2471 (N_2471,N_1880,In_147);
nor U2472 (N_2472,N_1874,N_1661);
or U2473 (N_2473,N_1020,In_2930);
or U2474 (N_2474,In_2750,N_1610);
nor U2475 (N_2475,N_1757,N_1725);
and U2476 (N_2476,N_1358,N_1593);
and U2477 (N_2477,In_1331,In_821);
and U2478 (N_2478,N_320,N_1533);
or U2479 (N_2479,N_735,N_1495);
nor U2480 (N_2480,N_301,N_603);
nand U2481 (N_2481,In_472,N_1652);
nand U2482 (N_2482,In_1854,N_1854);
xor U2483 (N_2483,N_1534,N_70);
nor U2484 (N_2484,N_1033,N_1788);
nor U2485 (N_2485,N_1643,N_1968);
xnor U2486 (N_2486,N_1825,N_1733);
or U2487 (N_2487,N_1756,N_1859);
nand U2488 (N_2488,N_1078,In_1160);
xor U2489 (N_2489,N_1616,N_1745);
xor U2490 (N_2490,N_1936,N_1833);
or U2491 (N_2491,In_1038,N_1486);
or U2492 (N_2492,N_1789,N_1605);
or U2493 (N_2493,N_1259,In_2167);
nand U2494 (N_2494,N_1089,N_1897);
xnor U2495 (N_2495,In_2570,N_1861);
or U2496 (N_2496,In_2177,In_2065);
or U2497 (N_2497,N_1552,N_885);
nand U2498 (N_2498,N_1672,N_1545);
or U2499 (N_2499,N_1055,N_14);
xor U2500 (N_2500,N_2239,N_2344);
nand U2501 (N_2501,N_2298,N_2156);
xnor U2502 (N_2502,N_2022,N_2209);
nand U2503 (N_2503,N_2073,N_2068);
nor U2504 (N_2504,N_2196,N_2017);
nor U2505 (N_2505,N_2304,N_2272);
nor U2506 (N_2506,N_2461,N_2244);
xnor U2507 (N_2507,N_2011,N_2417);
or U2508 (N_2508,N_2320,N_2149);
nor U2509 (N_2509,N_2111,N_2498);
nand U2510 (N_2510,N_2299,N_2015);
and U2511 (N_2511,N_2053,N_2201);
and U2512 (N_2512,N_2186,N_2338);
nand U2513 (N_2513,N_2402,N_2337);
nand U2514 (N_2514,N_2333,N_2019);
or U2515 (N_2515,N_2419,N_2357);
and U2516 (N_2516,N_2311,N_2375);
and U2517 (N_2517,N_2109,N_2356);
nor U2518 (N_2518,N_2308,N_2236);
nor U2519 (N_2519,N_2099,N_2121);
nor U2520 (N_2520,N_2076,N_2067);
and U2521 (N_2521,N_2421,N_2412);
nand U2522 (N_2522,N_2179,N_2314);
xor U2523 (N_2523,N_2413,N_2240);
or U2524 (N_2524,N_2460,N_2012);
and U2525 (N_2525,N_2322,N_2029);
nand U2526 (N_2526,N_2008,N_2214);
and U2527 (N_2527,N_2494,N_2164);
or U2528 (N_2528,N_2098,N_2300);
and U2529 (N_2529,N_2425,N_2075);
nand U2530 (N_2530,N_2282,N_2229);
nor U2531 (N_2531,N_2267,N_2296);
xnor U2532 (N_2532,N_2255,N_2443);
and U2533 (N_2533,N_2444,N_2104);
nand U2534 (N_2534,N_2043,N_2459);
or U2535 (N_2535,N_2090,N_2238);
nand U2536 (N_2536,N_2010,N_2166);
nand U2537 (N_2537,N_2061,N_2409);
or U2538 (N_2538,N_2364,N_2147);
or U2539 (N_2539,N_2354,N_2185);
nor U2540 (N_2540,N_2342,N_2458);
or U2541 (N_2541,N_2235,N_2477);
and U2542 (N_2542,N_2120,N_2007);
nand U2543 (N_2543,N_2231,N_2493);
and U2544 (N_2544,N_2031,N_2188);
nor U2545 (N_2545,N_2431,N_2155);
and U2546 (N_2546,N_2446,N_2327);
xnor U2547 (N_2547,N_2400,N_2290);
nor U2548 (N_2548,N_2315,N_2396);
and U2549 (N_2549,N_2004,N_2297);
nand U2550 (N_2550,N_2097,N_2347);
and U2551 (N_2551,N_2112,N_2197);
nand U2552 (N_2552,N_2441,N_2385);
nand U2553 (N_2553,N_2183,N_2034);
nand U2554 (N_2554,N_2005,N_2167);
xnor U2555 (N_2555,N_2135,N_2318);
nor U2556 (N_2556,N_2093,N_2384);
or U2557 (N_2557,N_2159,N_2449);
or U2558 (N_2558,N_2365,N_2251);
xor U2559 (N_2559,N_2323,N_2452);
nor U2560 (N_2560,N_2095,N_2100);
or U2561 (N_2561,N_2202,N_2285);
and U2562 (N_2562,N_2199,N_2144);
and U2563 (N_2563,N_2113,N_2165);
and U2564 (N_2564,N_2391,N_2062);
or U2565 (N_2565,N_2469,N_2148);
xnor U2566 (N_2566,N_2390,N_2230);
nand U2567 (N_2567,N_2271,N_2268);
and U2568 (N_2568,N_2335,N_2046);
or U2569 (N_2569,N_2142,N_2134);
and U2570 (N_2570,N_2281,N_2085);
or U2571 (N_2571,N_2439,N_2399);
or U2572 (N_2572,N_2146,N_2168);
xor U2573 (N_2573,N_2423,N_2169);
nor U2574 (N_2574,N_2374,N_2457);
and U2575 (N_2575,N_2137,N_2127);
or U2576 (N_2576,N_2198,N_2471);
and U2577 (N_2577,N_2380,N_2432);
or U2578 (N_2578,N_2274,N_2291);
and U2579 (N_2579,N_2130,N_2057);
and U2580 (N_2580,N_2252,N_2484);
nand U2581 (N_2581,N_2232,N_2077);
nor U2582 (N_2582,N_2411,N_2071);
nor U2583 (N_2583,N_2133,N_2486);
nand U2584 (N_2584,N_2348,N_2059);
nor U2585 (N_2585,N_2414,N_2237);
nand U2586 (N_2586,N_2042,N_2079);
nor U2587 (N_2587,N_2386,N_2036);
nor U2588 (N_2588,N_2225,N_2026);
nand U2589 (N_2589,N_2193,N_2138);
and U2590 (N_2590,N_2065,N_2490);
and U2591 (N_2591,N_2456,N_2301);
nor U2592 (N_2592,N_2243,N_2226);
nand U2593 (N_2593,N_2210,N_2270);
xnor U2594 (N_2594,N_2427,N_2454);
nand U2595 (N_2595,N_2448,N_2018);
or U2596 (N_2596,N_2241,N_2035);
nand U2597 (N_2597,N_2455,N_2253);
nor U2598 (N_2598,N_2242,N_2006);
nand U2599 (N_2599,N_2174,N_2211);
nand U2600 (N_2600,N_2420,N_2024);
or U2601 (N_2601,N_2033,N_2309);
nand U2602 (N_2602,N_2064,N_2050);
nor U2603 (N_2603,N_2372,N_2306);
xor U2604 (N_2604,N_2488,N_2125);
or U2605 (N_2605,N_2256,N_2378);
xor U2606 (N_2606,N_2078,N_2480);
xnor U2607 (N_2607,N_2436,N_2037);
and U2608 (N_2608,N_2447,N_2377);
or U2609 (N_2609,N_2361,N_2086);
nand U2610 (N_2610,N_2262,N_2213);
nor U2611 (N_2611,N_2048,N_2161);
nor U2612 (N_2612,N_2353,N_2223);
xor U2613 (N_2613,N_2258,N_2394);
nor U2614 (N_2614,N_2247,N_2286);
or U2615 (N_2615,N_2279,N_2330);
or U2616 (N_2616,N_2143,N_2195);
nand U2617 (N_2617,N_2221,N_2092);
nand U2618 (N_2618,N_2351,N_2101);
or U2619 (N_2619,N_2215,N_2094);
xor U2620 (N_2620,N_2462,N_2157);
nor U2621 (N_2621,N_2191,N_2319);
xnor U2622 (N_2622,N_2212,N_2217);
or U2623 (N_2623,N_2476,N_2328);
or U2624 (N_2624,N_2467,N_2352);
nand U2625 (N_2625,N_2389,N_2021);
nand U2626 (N_2626,N_2136,N_2485);
nand U2627 (N_2627,N_2478,N_2013);
and U2628 (N_2628,N_2336,N_2422);
nand U2629 (N_2629,N_2108,N_2023);
xnor U2630 (N_2630,N_2404,N_2069);
xor U2631 (N_2631,N_2481,N_2295);
or U2632 (N_2632,N_2317,N_2184);
or U2633 (N_2633,N_2141,N_2219);
and U2634 (N_2634,N_2056,N_2140);
nand U2635 (N_2635,N_2126,N_2429);
or U2636 (N_2636,N_2468,N_2265);
xnor U2637 (N_2637,N_2194,N_2181);
nor U2638 (N_2638,N_2233,N_2283);
nand U2639 (N_2639,N_2345,N_2341);
or U2640 (N_2640,N_2359,N_2039);
nand U2641 (N_2641,N_2128,N_2160);
nor U2642 (N_2642,N_2395,N_2131);
nand U2643 (N_2643,N_2055,N_2190);
nand U2644 (N_2644,N_2275,N_2234);
nor U2645 (N_2645,N_2246,N_2139);
or U2646 (N_2646,N_2278,N_2114);
or U2647 (N_2647,N_2316,N_2415);
or U2648 (N_2648,N_2122,N_2313);
or U2649 (N_2649,N_2170,N_2263);
or U2650 (N_2650,N_2366,N_2349);
nand U2651 (N_2651,N_2491,N_2000);
nor U2652 (N_2652,N_2277,N_2387);
nor U2653 (N_2653,N_2074,N_2398);
or U2654 (N_2654,N_2321,N_2116);
or U2655 (N_2655,N_2442,N_2003);
nand U2656 (N_2656,N_2350,N_2371);
or U2657 (N_2657,N_2206,N_2472);
nand U2658 (N_2658,N_2451,N_2189);
and U2659 (N_2659,N_2284,N_2045);
and U2660 (N_2660,N_2379,N_2192);
xnor U2661 (N_2661,N_2401,N_2424);
or U2662 (N_2662,N_2154,N_2176);
and U2663 (N_2663,N_2466,N_2107);
nand U2664 (N_2664,N_2257,N_2473);
and U2665 (N_2665,N_2463,N_2403);
nand U2666 (N_2666,N_2428,N_2080);
or U2667 (N_2667,N_2082,N_2020);
nor U2668 (N_2668,N_2204,N_2066);
nand U2669 (N_2669,N_2025,N_2117);
nor U2670 (N_2670,N_2002,N_2162);
or U2671 (N_2671,N_2177,N_2489);
or U2672 (N_2672,N_2228,N_2200);
nand U2673 (N_2673,N_2091,N_2203);
xnor U2674 (N_2674,N_2096,N_2450);
xnor U2675 (N_2675,N_2216,N_2307);
or U2676 (N_2676,N_2248,N_2180);
xor U2677 (N_2677,N_2260,N_2070);
and U2678 (N_2678,N_2362,N_2329);
nor U2679 (N_2679,N_2483,N_2393);
xnor U2680 (N_2680,N_2051,N_2261);
nor U2681 (N_2681,N_2178,N_2499);
nand U2682 (N_2682,N_2382,N_2266);
xnor U2683 (N_2683,N_2115,N_2249);
and U2684 (N_2684,N_2363,N_2305);
and U2685 (N_2685,N_2102,N_2383);
xnor U2686 (N_2686,N_2292,N_2287);
nand U2687 (N_2687,N_2171,N_2332);
nand U2688 (N_2688,N_2150,N_2250);
or U2689 (N_2689,N_2222,N_2433);
and U2690 (N_2690,N_2310,N_2381);
nor U2691 (N_2691,N_2016,N_2087);
xnor U2692 (N_2692,N_2355,N_2369);
and U2693 (N_2693,N_2325,N_2445);
xor U2694 (N_2694,N_2440,N_2058);
nor U2695 (N_2695,N_2106,N_2208);
nand U2696 (N_2696,N_2482,N_2269);
nor U2697 (N_2697,N_2172,N_2132);
or U2698 (N_2698,N_2118,N_2406);
or U2699 (N_2699,N_2453,N_2001);
and U2700 (N_2700,N_2264,N_2392);
nand U2701 (N_2701,N_2028,N_2302);
xnor U2702 (N_2702,N_2339,N_2294);
or U2703 (N_2703,N_2175,N_2492);
nand U2704 (N_2704,N_2370,N_2105);
xnor U2705 (N_2705,N_2205,N_2324);
or U2706 (N_2706,N_2273,N_2388);
nand U2707 (N_2707,N_2464,N_2129);
and U2708 (N_2708,N_2430,N_2410);
nand U2709 (N_2709,N_2331,N_2303);
and U2710 (N_2710,N_2312,N_2276);
nand U2711 (N_2711,N_2474,N_2081);
nor U2712 (N_2712,N_2437,N_2495);
and U2713 (N_2713,N_2334,N_2416);
nand U2714 (N_2714,N_2435,N_2368);
nand U2715 (N_2715,N_2434,N_2340);
nor U2716 (N_2716,N_2124,N_2052);
or U2717 (N_2717,N_2254,N_2418);
or U2718 (N_2718,N_2373,N_2153);
or U2719 (N_2719,N_2224,N_2426);
and U2720 (N_2720,N_2245,N_2376);
and U2721 (N_2721,N_2479,N_2346);
or U2722 (N_2722,N_2293,N_2009);
nand U2723 (N_2723,N_2083,N_2218);
nor U2724 (N_2724,N_2182,N_2088);
nor U2725 (N_2725,N_2497,N_2358);
nand U2726 (N_2726,N_2049,N_2060);
and U2727 (N_2727,N_2367,N_2465);
and U2728 (N_2728,N_2470,N_2288);
nor U2729 (N_2729,N_2405,N_2173);
and U2730 (N_2730,N_2041,N_2397);
nor U2731 (N_2731,N_2063,N_2084);
nand U2732 (N_2732,N_2259,N_2038);
nor U2733 (N_2733,N_2027,N_2326);
nor U2734 (N_2734,N_2072,N_2207);
nor U2735 (N_2735,N_2496,N_2110);
nand U2736 (N_2736,N_2343,N_2220);
or U2737 (N_2737,N_2030,N_2014);
xnor U2738 (N_2738,N_2151,N_2289);
and U2739 (N_2739,N_2119,N_2152);
nor U2740 (N_2740,N_2044,N_2227);
nor U2741 (N_2741,N_2475,N_2032);
xor U2742 (N_2742,N_2360,N_2054);
nor U2743 (N_2743,N_2158,N_2438);
and U2744 (N_2744,N_2047,N_2280);
and U2745 (N_2745,N_2487,N_2407);
nand U2746 (N_2746,N_2040,N_2103);
and U2747 (N_2747,N_2089,N_2145);
nor U2748 (N_2748,N_2408,N_2163);
and U2749 (N_2749,N_2187,N_2123);
or U2750 (N_2750,N_2309,N_2001);
nor U2751 (N_2751,N_2026,N_2283);
xor U2752 (N_2752,N_2251,N_2493);
nor U2753 (N_2753,N_2325,N_2477);
nor U2754 (N_2754,N_2261,N_2000);
nand U2755 (N_2755,N_2321,N_2280);
and U2756 (N_2756,N_2124,N_2264);
xnor U2757 (N_2757,N_2382,N_2101);
nor U2758 (N_2758,N_2226,N_2438);
nand U2759 (N_2759,N_2166,N_2072);
xnor U2760 (N_2760,N_2446,N_2244);
xor U2761 (N_2761,N_2409,N_2218);
nor U2762 (N_2762,N_2231,N_2355);
and U2763 (N_2763,N_2242,N_2379);
nor U2764 (N_2764,N_2037,N_2215);
nand U2765 (N_2765,N_2179,N_2437);
or U2766 (N_2766,N_2139,N_2304);
nand U2767 (N_2767,N_2239,N_2056);
or U2768 (N_2768,N_2113,N_2042);
nand U2769 (N_2769,N_2124,N_2185);
xor U2770 (N_2770,N_2458,N_2102);
xnor U2771 (N_2771,N_2158,N_2465);
and U2772 (N_2772,N_2275,N_2185);
nor U2773 (N_2773,N_2246,N_2015);
or U2774 (N_2774,N_2479,N_2448);
and U2775 (N_2775,N_2438,N_2201);
or U2776 (N_2776,N_2120,N_2201);
and U2777 (N_2777,N_2296,N_2304);
nor U2778 (N_2778,N_2449,N_2039);
and U2779 (N_2779,N_2474,N_2045);
nand U2780 (N_2780,N_2253,N_2088);
or U2781 (N_2781,N_2387,N_2475);
nor U2782 (N_2782,N_2280,N_2344);
and U2783 (N_2783,N_2310,N_2061);
xnor U2784 (N_2784,N_2317,N_2361);
and U2785 (N_2785,N_2073,N_2262);
nand U2786 (N_2786,N_2149,N_2232);
nor U2787 (N_2787,N_2223,N_2176);
or U2788 (N_2788,N_2059,N_2360);
nand U2789 (N_2789,N_2282,N_2217);
xor U2790 (N_2790,N_2418,N_2274);
or U2791 (N_2791,N_2378,N_2393);
nor U2792 (N_2792,N_2466,N_2058);
xnor U2793 (N_2793,N_2033,N_2101);
and U2794 (N_2794,N_2303,N_2218);
or U2795 (N_2795,N_2003,N_2063);
nor U2796 (N_2796,N_2047,N_2240);
or U2797 (N_2797,N_2417,N_2449);
nand U2798 (N_2798,N_2259,N_2386);
or U2799 (N_2799,N_2073,N_2385);
and U2800 (N_2800,N_2431,N_2051);
nor U2801 (N_2801,N_2096,N_2036);
xor U2802 (N_2802,N_2264,N_2275);
and U2803 (N_2803,N_2393,N_2181);
xor U2804 (N_2804,N_2354,N_2482);
or U2805 (N_2805,N_2435,N_2047);
nor U2806 (N_2806,N_2277,N_2045);
and U2807 (N_2807,N_2025,N_2013);
and U2808 (N_2808,N_2023,N_2268);
nor U2809 (N_2809,N_2497,N_2172);
and U2810 (N_2810,N_2401,N_2438);
nand U2811 (N_2811,N_2052,N_2313);
and U2812 (N_2812,N_2074,N_2080);
nor U2813 (N_2813,N_2136,N_2466);
nor U2814 (N_2814,N_2041,N_2178);
or U2815 (N_2815,N_2315,N_2065);
nand U2816 (N_2816,N_2364,N_2184);
or U2817 (N_2817,N_2066,N_2288);
nor U2818 (N_2818,N_2108,N_2320);
xnor U2819 (N_2819,N_2218,N_2229);
nor U2820 (N_2820,N_2014,N_2436);
nand U2821 (N_2821,N_2002,N_2435);
or U2822 (N_2822,N_2307,N_2122);
and U2823 (N_2823,N_2440,N_2443);
and U2824 (N_2824,N_2038,N_2103);
nor U2825 (N_2825,N_2371,N_2394);
and U2826 (N_2826,N_2247,N_2244);
nor U2827 (N_2827,N_2469,N_2228);
and U2828 (N_2828,N_2418,N_2022);
nand U2829 (N_2829,N_2225,N_2046);
nor U2830 (N_2830,N_2433,N_2343);
or U2831 (N_2831,N_2335,N_2288);
nand U2832 (N_2832,N_2055,N_2057);
nand U2833 (N_2833,N_2472,N_2156);
or U2834 (N_2834,N_2337,N_2060);
nand U2835 (N_2835,N_2365,N_2039);
nand U2836 (N_2836,N_2276,N_2391);
and U2837 (N_2837,N_2043,N_2144);
nand U2838 (N_2838,N_2353,N_2240);
nor U2839 (N_2839,N_2243,N_2179);
nor U2840 (N_2840,N_2180,N_2317);
and U2841 (N_2841,N_2034,N_2016);
xor U2842 (N_2842,N_2318,N_2331);
or U2843 (N_2843,N_2288,N_2456);
or U2844 (N_2844,N_2235,N_2009);
xnor U2845 (N_2845,N_2496,N_2347);
nand U2846 (N_2846,N_2091,N_2060);
nand U2847 (N_2847,N_2019,N_2143);
or U2848 (N_2848,N_2480,N_2115);
and U2849 (N_2849,N_2434,N_2378);
nor U2850 (N_2850,N_2062,N_2274);
and U2851 (N_2851,N_2199,N_2045);
xor U2852 (N_2852,N_2318,N_2420);
nand U2853 (N_2853,N_2211,N_2118);
and U2854 (N_2854,N_2339,N_2412);
nor U2855 (N_2855,N_2342,N_2455);
or U2856 (N_2856,N_2421,N_2448);
nand U2857 (N_2857,N_2213,N_2168);
xor U2858 (N_2858,N_2387,N_2110);
nor U2859 (N_2859,N_2374,N_2009);
or U2860 (N_2860,N_2054,N_2087);
nand U2861 (N_2861,N_2486,N_2487);
and U2862 (N_2862,N_2435,N_2369);
nand U2863 (N_2863,N_2094,N_2180);
xnor U2864 (N_2864,N_2450,N_2142);
xnor U2865 (N_2865,N_2484,N_2441);
xnor U2866 (N_2866,N_2136,N_2016);
xor U2867 (N_2867,N_2255,N_2130);
xor U2868 (N_2868,N_2050,N_2259);
nor U2869 (N_2869,N_2395,N_2489);
nor U2870 (N_2870,N_2122,N_2444);
and U2871 (N_2871,N_2219,N_2491);
nand U2872 (N_2872,N_2499,N_2458);
xnor U2873 (N_2873,N_2338,N_2050);
xor U2874 (N_2874,N_2315,N_2302);
nand U2875 (N_2875,N_2291,N_2017);
and U2876 (N_2876,N_2101,N_2482);
nand U2877 (N_2877,N_2488,N_2353);
and U2878 (N_2878,N_2180,N_2413);
and U2879 (N_2879,N_2458,N_2011);
xor U2880 (N_2880,N_2196,N_2424);
or U2881 (N_2881,N_2243,N_2102);
nor U2882 (N_2882,N_2340,N_2128);
or U2883 (N_2883,N_2348,N_2297);
and U2884 (N_2884,N_2196,N_2486);
nand U2885 (N_2885,N_2459,N_2102);
or U2886 (N_2886,N_2165,N_2486);
or U2887 (N_2887,N_2309,N_2323);
xnor U2888 (N_2888,N_2351,N_2427);
nand U2889 (N_2889,N_2175,N_2385);
nand U2890 (N_2890,N_2289,N_2355);
nor U2891 (N_2891,N_2452,N_2268);
nand U2892 (N_2892,N_2228,N_2437);
xnor U2893 (N_2893,N_2312,N_2130);
xnor U2894 (N_2894,N_2497,N_2198);
xnor U2895 (N_2895,N_2257,N_2099);
nor U2896 (N_2896,N_2272,N_2245);
nand U2897 (N_2897,N_2172,N_2096);
xnor U2898 (N_2898,N_2142,N_2276);
or U2899 (N_2899,N_2006,N_2286);
xor U2900 (N_2900,N_2249,N_2219);
and U2901 (N_2901,N_2322,N_2153);
and U2902 (N_2902,N_2485,N_2274);
nand U2903 (N_2903,N_2311,N_2187);
nand U2904 (N_2904,N_2187,N_2095);
and U2905 (N_2905,N_2111,N_2090);
and U2906 (N_2906,N_2251,N_2096);
xnor U2907 (N_2907,N_2106,N_2158);
nand U2908 (N_2908,N_2060,N_2377);
and U2909 (N_2909,N_2244,N_2365);
nor U2910 (N_2910,N_2007,N_2345);
and U2911 (N_2911,N_2013,N_2196);
or U2912 (N_2912,N_2188,N_2254);
nand U2913 (N_2913,N_2050,N_2071);
nand U2914 (N_2914,N_2076,N_2180);
nand U2915 (N_2915,N_2077,N_2477);
and U2916 (N_2916,N_2414,N_2107);
nor U2917 (N_2917,N_2240,N_2474);
xnor U2918 (N_2918,N_2190,N_2145);
nor U2919 (N_2919,N_2345,N_2027);
nor U2920 (N_2920,N_2360,N_2124);
xor U2921 (N_2921,N_2154,N_2315);
xnor U2922 (N_2922,N_2000,N_2465);
or U2923 (N_2923,N_2152,N_2408);
nor U2924 (N_2924,N_2160,N_2090);
and U2925 (N_2925,N_2159,N_2015);
and U2926 (N_2926,N_2016,N_2058);
or U2927 (N_2927,N_2334,N_2078);
xor U2928 (N_2928,N_2029,N_2439);
xnor U2929 (N_2929,N_2234,N_2173);
nor U2930 (N_2930,N_2009,N_2004);
xnor U2931 (N_2931,N_2221,N_2013);
nand U2932 (N_2932,N_2404,N_2021);
and U2933 (N_2933,N_2441,N_2341);
xnor U2934 (N_2934,N_2320,N_2387);
xnor U2935 (N_2935,N_2431,N_2205);
and U2936 (N_2936,N_2082,N_2078);
and U2937 (N_2937,N_2393,N_2230);
nand U2938 (N_2938,N_2343,N_2138);
nand U2939 (N_2939,N_2085,N_2118);
nor U2940 (N_2940,N_2140,N_2083);
and U2941 (N_2941,N_2071,N_2014);
or U2942 (N_2942,N_2194,N_2204);
or U2943 (N_2943,N_2453,N_2407);
nand U2944 (N_2944,N_2193,N_2293);
xor U2945 (N_2945,N_2351,N_2221);
xor U2946 (N_2946,N_2222,N_2261);
or U2947 (N_2947,N_2394,N_2231);
nor U2948 (N_2948,N_2325,N_2191);
xor U2949 (N_2949,N_2033,N_2053);
and U2950 (N_2950,N_2105,N_2308);
and U2951 (N_2951,N_2197,N_2345);
xor U2952 (N_2952,N_2037,N_2406);
and U2953 (N_2953,N_2349,N_2144);
and U2954 (N_2954,N_2003,N_2001);
xor U2955 (N_2955,N_2480,N_2417);
and U2956 (N_2956,N_2331,N_2139);
nand U2957 (N_2957,N_2188,N_2130);
nor U2958 (N_2958,N_2097,N_2192);
nand U2959 (N_2959,N_2137,N_2426);
xor U2960 (N_2960,N_2435,N_2139);
and U2961 (N_2961,N_2156,N_2023);
and U2962 (N_2962,N_2336,N_2201);
nor U2963 (N_2963,N_2248,N_2186);
or U2964 (N_2964,N_2210,N_2081);
xnor U2965 (N_2965,N_2437,N_2306);
nor U2966 (N_2966,N_2124,N_2170);
and U2967 (N_2967,N_2083,N_2245);
nand U2968 (N_2968,N_2136,N_2150);
nor U2969 (N_2969,N_2379,N_2445);
nand U2970 (N_2970,N_2198,N_2328);
xnor U2971 (N_2971,N_2214,N_2210);
or U2972 (N_2972,N_2370,N_2150);
or U2973 (N_2973,N_2263,N_2438);
or U2974 (N_2974,N_2431,N_2380);
and U2975 (N_2975,N_2154,N_2020);
nor U2976 (N_2976,N_2304,N_2385);
nor U2977 (N_2977,N_2436,N_2480);
nand U2978 (N_2978,N_2264,N_2024);
nand U2979 (N_2979,N_2020,N_2102);
or U2980 (N_2980,N_2280,N_2031);
nand U2981 (N_2981,N_2363,N_2111);
and U2982 (N_2982,N_2392,N_2381);
xor U2983 (N_2983,N_2053,N_2213);
and U2984 (N_2984,N_2212,N_2384);
and U2985 (N_2985,N_2402,N_2495);
or U2986 (N_2986,N_2231,N_2157);
or U2987 (N_2987,N_2209,N_2494);
or U2988 (N_2988,N_2247,N_2175);
nand U2989 (N_2989,N_2099,N_2196);
xor U2990 (N_2990,N_2164,N_2273);
nor U2991 (N_2991,N_2009,N_2396);
nand U2992 (N_2992,N_2482,N_2263);
and U2993 (N_2993,N_2241,N_2021);
nand U2994 (N_2994,N_2434,N_2088);
or U2995 (N_2995,N_2365,N_2487);
nand U2996 (N_2996,N_2401,N_2307);
nand U2997 (N_2997,N_2302,N_2006);
nor U2998 (N_2998,N_2078,N_2362);
xnor U2999 (N_2999,N_2388,N_2413);
nor U3000 (N_3000,N_2854,N_2600);
nor U3001 (N_3001,N_2861,N_2834);
xor U3002 (N_3002,N_2845,N_2869);
xnor U3003 (N_3003,N_2805,N_2786);
nor U3004 (N_3004,N_2978,N_2703);
and U3005 (N_3005,N_2525,N_2524);
xor U3006 (N_3006,N_2716,N_2668);
xnor U3007 (N_3007,N_2530,N_2729);
or U3008 (N_3008,N_2622,N_2577);
nand U3009 (N_3009,N_2724,N_2635);
xnor U3010 (N_3010,N_2645,N_2938);
nor U3011 (N_3011,N_2793,N_2826);
nand U3012 (N_3012,N_2986,N_2999);
or U3013 (N_3013,N_2552,N_2578);
and U3014 (N_3014,N_2897,N_2798);
nand U3015 (N_3015,N_2753,N_2662);
xor U3016 (N_3016,N_2891,N_2658);
nor U3017 (N_3017,N_2732,N_2795);
and U3018 (N_3018,N_2933,N_2997);
and U3019 (N_3019,N_2500,N_2941);
nor U3020 (N_3020,N_2783,N_2603);
and U3021 (N_3021,N_2556,N_2972);
and U3022 (N_3022,N_2537,N_2632);
xor U3023 (N_3023,N_2914,N_2850);
nor U3024 (N_3024,N_2708,N_2613);
xor U3025 (N_3025,N_2792,N_2769);
nand U3026 (N_3026,N_2693,N_2928);
nor U3027 (N_3027,N_2902,N_2947);
nor U3028 (N_3028,N_2871,N_2961);
nor U3029 (N_3029,N_2772,N_2888);
nor U3030 (N_3030,N_2699,N_2735);
and U3031 (N_3031,N_2936,N_2592);
or U3032 (N_3032,N_2679,N_2591);
nor U3033 (N_3033,N_2759,N_2881);
nor U3034 (N_3034,N_2754,N_2589);
nor U3035 (N_3035,N_2559,N_2810);
nor U3036 (N_3036,N_2538,N_2782);
xnor U3037 (N_3037,N_2915,N_2824);
xnor U3038 (N_3038,N_2619,N_2837);
nor U3039 (N_3039,N_2949,N_2706);
or U3040 (N_3040,N_2852,N_2534);
and U3041 (N_3041,N_2670,N_2627);
nand U3042 (N_3042,N_2833,N_2704);
or U3043 (N_3043,N_2916,N_2554);
nor U3044 (N_3044,N_2730,N_2581);
nand U3045 (N_3045,N_2715,N_2757);
xnor U3046 (N_3046,N_2697,N_2975);
xor U3047 (N_3047,N_2889,N_2643);
xnor U3048 (N_3048,N_2701,N_2971);
or U3049 (N_3049,N_2895,N_2504);
and U3050 (N_3050,N_2996,N_2566);
xnor U3051 (N_3051,N_2896,N_2934);
or U3052 (N_3052,N_2940,N_2501);
nor U3053 (N_3053,N_2840,N_2744);
and U3054 (N_3054,N_2980,N_2683);
nand U3055 (N_3055,N_2765,N_2666);
and U3056 (N_3056,N_2580,N_2541);
and U3057 (N_3057,N_2582,N_2721);
or U3058 (N_3058,N_2644,N_2751);
and U3059 (N_3059,N_2848,N_2790);
or U3060 (N_3060,N_2809,N_2521);
nor U3061 (N_3061,N_2954,N_2626);
and U3062 (N_3062,N_2617,N_2512);
xor U3063 (N_3063,N_2791,N_2696);
nand U3064 (N_3064,N_2540,N_2630);
nand U3065 (N_3065,N_2987,N_2728);
and U3066 (N_3066,N_2787,N_2799);
nand U3067 (N_3067,N_2758,N_2962);
xor U3068 (N_3068,N_2719,N_2515);
nor U3069 (N_3069,N_2640,N_2514);
or U3070 (N_3070,N_2857,N_2907);
and U3071 (N_3071,N_2605,N_2688);
nor U3072 (N_3072,N_2988,N_2746);
and U3073 (N_3073,N_2620,N_2846);
and U3074 (N_3074,N_2633,N_2979);
nor U3075 (N_3075,N_2764,N_2808);
nand U3076 (N_3076,N_2939,N_2502);
and U3077 (N_3077,N_2612,N_2748);
or U3078 (N_3078,N_2653,N_2648);
nand U3079 (N_3079,N_2522,N_2647);
nor U3080 (N_3080,N_2796,N_2776);
nand U3081 (N_3081,N_2536,N_2803);
or U3082 (N_3082,N_2761,N_2775);
xnor U3083 (N_3083,N_2637,N_2771);
and U3084 (N_3084,N_2737,N_2678);
and U3085 (N_3085,N_2596,N_2731);
or U3086 (N_3086,N_2767,N_2667);
nand U3087 (N_3087,N_2567,N_2866);
nor U3088 (N_3088,N_2953,N_2563);
nand U3089 (N_3089,N_2905,N_2685);
and U3090 (N_3090,N_2970,N_2562);
nand U3091 (N_3091,N_2608,N_2654);
nand U3092 (N_3092,N_2739,N_2867);
or U3093 (N_3093,N_2526,N_2817);
or U3094 (N_3094,N_2955,N_2991);
nand U3095 (N_3095,N_2836,N_2831);
nand U3096 (N_3096,N_2990,N_2781);
xor U3097 (N_3097,N_2827,N_2646);
or U3098 (N_3098,N_2985,N_2920);
and U3099 (N_3099,N_2887,N_2686);
nor U3100 (N_3100,N_2777,N_2665);
nor U3101 (N_3101,N_2804,N_2872);
nor U3102 (N_3102,N_2569,N_2992);
xor U3103 (N_3103,N_2516,N_2814);
or U3104 (N_3104,N_2820,N_2993);
and U3105 (N_3105,N_2585,N_2952);
nor U3106 (N_3106,N_2838,N_2707);
nor U3107 (N_3107,N_2599,N_2691);
or U3108 (N_3108,N_2963,N_2573);
nor U3109 (N_3109,N_2885,N_2723);
nand U3110 (N_3110,N_2564,N_2998);
nor U3111 (N_3111,N_2863,N_2921);
nand U3112 (N_3112,N_2811,N_2948);
and U3113 (N_3113,N_2511,N_2806);
xor U3114 (N_3114,N_2532,N_2752);
nor U3115 (N_3115,N_2788,N_2880);
or U3116 (N_3116,N_2631,N_2742);
nor U3117 (N_3117,N_2802,N_2832);
nand U3118 (N_3118,N_2908,N_2588);
nand U3119 (N_3119,N_2579,N_2917);
nor U3120 (N_3120,N_2784,N_2960);
xor U3121 (N_3121,N_2584,N_2576);
xnor U3122 (N_3122,N_2506,N_2779);
or U3123 (N_3123,N_2574,N_2884);
xnor U3124 (N_3124,N_2571,N_2904);
nand U3125 (N_3125,N_2642,N_2894);
and U3126 (N_3126,N_2957,N_2956);
nand U3127 (N_3127,N_2713,N_2702);
nor U3128 (N_3128,N_2828,N_2813);
or U3129 (N_3129,N_2763,N_2520);
nand U3130 (N_3130,N_2812,N_2656);
and U3131 (N_3131,N_2964,N_2539);
or U3132 (N_3132,N_2733,N_2821);
xnor U3133 (N_3133,N_2676,N_2565);
nand U3134 (N_3134,N_2590,N_2594);
nand U3135 (N_3135,N_2523,N_2892);
nand U3136 (N_3136,N_2641,N_2692);
nor U3137 (N_3137,N_2655,N_2937);
or U3138 (N_3138,N_2684,N_2950);
nor U3139 (N_3139,N_2965,N_2705);
nand U3140 (N_3140,N_2507,N_2882);
xnor U3141 (N_3141,N_2572,N_2621);
and U3142 (N_3142,N_2968,N_2910);
xor U3143 (N_3143,N_2844,N_2913);
or U3144 (N_3144,N_2551,N_2879);
nand U3145 (N_3145,N_2661,N_2690);
or U3146 (N_3146,N_2529,N_2741);
nor U3147 (N_3147,N_2710,N_2973);
and U3148 (N_3148,N_2624,N_2816);
and U3149 (N_3149,N_2994,N_2636);
xnor U3150 (N_3150,N_2736,N_2597);
nor U3151 (N_3151,N_2595,N_2543);
nand U3152 (N_3152,N_2877,N_2926);
and U3153 (N_3153,N_2918,N_2602);
or U3154 (N_3154,N_2923,N_2760);
nor U3155 (N_3155,N_2510,N_2815);
and U3156 (N_3156,N_2958,N_2568);
nand U3157 (N_3157,N_2652,N_2931);
or U3158 (N_3158,N_2601,N_2528);
and U3159 (N_3159,N_2743,N_2542);
or U3160 (N_3160,N_2976,N_2680);
and U3161 (N_3161,N_2853,N_2943);
xnor U3162 (N_3162,N_2616,N_2677);
or U3163 (N_3163,N_2720,N_2818);
nor U3164 (N_3164,N_2570,N_2995);
and U3165 (N_3165,N_2660,N_2924);
nor U3166 (N_3166,N_2583,N_2780);
nor U3167 (N_3167,N_2835,N_2945);
nor U3168 (N_3168,N_2984,N_2819);
nand U3169 (N_3169,N_2927,N_2778);
nand U3170 (N_3170,N_2919,N_2989);
and U3171 (N_3171,N_2638,N_2909);
nand U3172 (N_3172,N_2575,N_2825);
and U3173 (N_3173,N_2935,N_2858);
xor U3174 (N_3174,N_2823,N_2557);
nor U3175 (N_3175,N_2615,N_2587);
nand U3176 (N_3176,N_2883,N_2714);
xor U3177 (N_3177,N_2614,N_2893);
and U3178 (N_3178,N_2898,N_2906);
xor U3179 (N_3179,N_2982,N_2847);
nand U3180 (N_3180,N_2930,N_2762);
nand U3181 (N_3181,N_2509,N_2586);
xnor U3182 (N_3182,N_2870,N_2681);
nand U3183 (N_3183,N_2698,N_2830);
xor U3184 (N_3184,N_2669,N_2531);
or U3185 (N_3185,N_2868,N_2800);
xnor U3186 (N_3186,N_2773,N_2768);
nand U3187 (N_3187,N_2709,N_2651);
or U3188 (N_3188,N_2722,N_2864);
and U3189 (N_3189,N_2747,N_2750);
nor U3190 (N_3190,N_2983,N_2607);
xor U3191 (N_3191,N_2561,N_2829);
nand U3192 (N_3192,N_2929,N_2900);
or U3193 (N_3193,N_2518,N_2598);
and U3194 (N_3194,N_2673,N_2593);
nand U3195 (N_3195,N_2689,N_2508);
nand U3196 (N_3196,N_2807,N_2755);
nor U3197 (N_3197,N_2674,N_2860);
xor U3198 (N_3198,N_2553,N_2560);
or U3199 (N_3199,N_2547,N_2756);
nor U3200 (N_3200,N_2944,N_2544);
or U3201 (N_3201,N_2634,N_2801);
or U3202 (N_3202,N_2903,N_2946);
nor U3203 (N_3203,N_2650,N_2695);
nor U3204 (N_3204,N_2745,N_2770);
and U3205 (N_3205,N_2628,N_2664);
or U3206 (N_3206,N_2841,N_2873);
or U3207 (N_3207,N_2517,N_2558);
xnor U3208 (N_3208,N_2513,N_2546);
xnor U3209 (N_3209,N_2951,N_2878);
or U3210 (N_3210,N_2505,N_2749);
and U3211 (N_3211,N_2843,N_2639);
and U3212 (N_3212,N_2610,N_2865);
xnor U3213 (N_3213,N_2682,N_2967);
and U3214 (N_3214,N_2727,N_2711);
and U3215 (N_3215,N_2981,N_2663);
nand U3216 (N_3216,N_2527,N_2875);
xnor U3217 (N_3217,N_2901,N_2671);
or U3218 (N_3218,N_2874,N_2842);
xor U3219 (N_3219,N_2851,N_2548);
nand U3220 (N_3220,N_2932,N_2922);
nand U3221 (N_3221,N_2899,N_2659);
nor U3222 (N_3222,N_2550,N_2609);
and U3223 (N_3223,N_2797,N_2738);
xor U3224 (N_3224,N_2625,N_2977);
or U3225 (N_3225,N_2687,N_2911);
or U3226 (N_3226,N_2734,N_2549);
or U3227 (N_3227,N_2611,N_2606);
nor U3228 (N_3228,N_2503,N_2649);
nand U3229 (N_3229,N_2694,N_2672);
or U3230 (N_3230,N_2712,N_2789);
and U3231 (N_3231,N_2912,N_2766);
and U3232 (N_3232,N_2629,N_2700);
or U3233 (N_3233,N_2855,N_2726);
and U3234 (N_3234,N_2839,N_2675);
and U3235 (N_3235,N_2822,N_2849);
and U3236 (N_3236,N_2545,N_2657);
or U3237 (N_3237,N_2886,N_2862);
nor U3238 (N_3238,N_2856,N_2618);
or U3239 (N_3239,N_2925,N_2794);
nand U3240 (N_3240,N_2966,N_2959);
or U3241 (N_3241,N_2725,N_2533);
nor U3242 (N_3242,N_2555,N_2969);
nand U3243 (N_3243,N_2604,N_2535);
and U3244 (N_3244,N_2859,N_2623);
and U3245 (N_3245,N_2774,N_2718);
nor U3246 (N_3246,N_2890,N_2942);
nor U3247 (N_3247,N_2519,N_2876);
nand U3248 (N_3248,N_2740,N_2717);
and U3249 (N_3249,N_2974,N_2785);
and U3250 (N_3250,N_2780,N_2959);
nor U3251 (N_3251,N_2932,N_2830);
xnor U3252 (N_3252,N_2911,N_2921);
xor U3253 (N_3253,N_2520,N_2536);
nor U3254 (N_3254,N_2935,N_2955);
xor U3255 (N_3255,N_2839,N_2520);
xnor U3256 (N_3256,N_2921,N_2638);
and U3257 (N_3257,N_2744,N_2692);
or U3258 (N_3258,N_2621,N_2702);
or U3259 (N_3259,N_2593,N_2741);
or U3260 (N_3260,N_2793,N_2709);
nor U3261 (N_3261,N_2848,N_2839);
nand U3262 (N_3262,N_2751,N_2670);
and U3263 (N_3263,N_2564,N_2982);
nor U3264 (N_3264,N_2918,N_2692);
nor U3265 (N_3265,N_2552,N_2764);
nor U3266 (N_3266,N_2612,N_2894);
and U3267 (N_3267,N_2765,N_2599);
nand U3268 (N_3268,N_2819,N_2719);
or U3269 (N_3269,N_2947,N_2555);
xor U3270 (N_3270,N_2788,N_2618);
nor U3271 (N_3271,N_2716,N_2676);
nor U3272 (N_3272,N_2582,N_2831);
and U3273 (N_3273,N_2861,N_2756);
nand U3274 (N_3274,N_2901,N_2964);
xor U3275 (N_3275,N_2822,N_2553);
nand U3276 (N_3276,N_2953,N_2959);
xnor U3277 (N_3277,N_2984,N_2692);
nand U3278 (N_3278,N_2850,N_2588);
nor U3279 (N_3279,N_2518,N_2613);
nand U3280 (N_3280,N_2986,N_2912);
and U3281 (N_3281,N_2885,N_2796);
xor U3282 (N_3282,N_2966,N_2699);
nand U3283 (N_3283,N_2883,N_2884);
or U3284 (N_3284,N_2917,N_2993);
xnor U3285 (N_3285,N_2655,N_2640);
or U3286 (N_3286,N_2540,N_2845);
nor U3287 (N_3287,N_2758,N_2656);
or U3288 (N_3288,N_2846,N_2501);
or U3289 (N_3289,N_2505,N_2864);
nor U3290 (N_3290,N_2935,N_2828);
xnor U3291 (N_3291,N_2762,N_2885);
xor U3292 (N_3292,N_2659,N_2651);
nor U3293 (N_3293,N_2513,N_2651);
nor U3294 (N_3294,N_2586,N_2669);
nor U3295 (N_3295,N_2956,N_2717);
or U3296 (N_3296,N_2618,N_2621);
xor U3297 (N_3297,N_2689,N_2740);
nor U3298 (N_3298,N_2632,N_2666);
nor U3299 (N_3299,N_2569,N_2651);
xnor U3300 (N_3300,N_2867,N_2632);
and U3301 (N_3301,N_2536,N_2719);
nand U3302 (N_3302,N_2946,N_2931);
xnor U3303 (N_3303,N_2835,N_2599);
xnor U3304 (N_3304,N_2837,N_2979);
nand U3305 (N_3305,N_2733,N_2945);
nand U3306 (N_3306,N_2620,N_2546);
or U3307 (N_3307,N_2639,N_2864);
or U3308 (N_3308,N_2647,N_2712);
nor U3309 (N_3309,N_2532,N_2593);
nor U3310 (N_3310,N_2679,N_2575);
nor U3311 (N_3311,N_2692,N_2891);
or U3312 (N_3312,N_2573,N_2720);
or U3313 (N_3313,N_2530,N_2741);
and U3314 (N_3314,N_2702,N_2717);
nand U3315 (N_3315,N_2556,N_2746);
nor U3316 (N_3316,N_2724,N_2859);
nand U3317 (N_3317,N_2787,N_2623);
and U3318 (N_3318,N_2547,N_2876);
nor U3319 (N_3319,N_2973,N_2965);
nor U3320 (N_3320,N_2615,N_2901);
and U3321 (N_3321,N_2538,N_2981);
xor U3322 (N_3322,N_2691,N_2680);
xnor U3323 (N_3323,N_2967,N_2962);
nor U3324 (N_3324,N_2695,N_2717);
or U3325 (N_3325,N_2781,N_2731);
or U3326 (N_3326,N_2970,N_2533);
nand U3327 (N_3327,N_2803,N_2523);
xor U3328 (N_3328,N_2593,N_2972);
nand U3329 (N_3329,N_2636,N_2877);
nor U3330 (N_3330,N_2611,N_2604);
nand U3331 (N_3331,N_2761,N_2961);
xnor U3332 (N_3332,N_2518,N_2712);
nor U3333 (N_3333,N_2686,N_2873);
and U3334 (N_3334,N_2627,N_2950);
and U3335 (N_3335,N_2958,N_2747);
and U3336 (N_3336,N_2679,N_2594);
nor U3337 (N_3337,N_2797,N_2718);
nor U3338 (N_3338,N_2635,N_2973);
xnor U3339 (N_3339,N_2595,N_2817);
nand U3340 (N_3340,N_2752,N_2878);
xnor U3341 (N_3341,N_2890,N_2508);
nor U3342 (N_3342,N_2742,N_2878);
and U3343 (N_3343,N_2574,N_2747);
nor U3344 (N_3344,N_2928,N_2534);
or U3345 (N_3345,N_2685,N_2759);
nand U3346 (N_3346,N_2875,N_2584);
and U3347 (N_3347,N_2557,N_2551);
or U3348 (N_3348,N_2862,N_2754);
nand U3349 (N_3349,N_2633,N_2725);
xnor U3350 (N_3350,N_2959,N_2848);
or U3351 (N_3351,N_2807,N_2995);
xnor U3352 (N_3352,N_2832,N_2680);
nor U3353 (N_3353,N_2500,N_2601);
nor U3354 (N_3354,N_2900,N_2573);
or U3355 (N_3355,N_2516,N_2560);
xor U3356 (N_3356,N_2782,N_2893);
and U3357 (N_3357,N_2624,N_2920);
nor U3358 (N_3358,N_2709,N_2835);
or U3359 (N_3359,N_2690,N_2827);
and U3360 (N_3360,N_2770,N_2952);
and U3361 (N_3361,N_2796,N_2772);
or U3362 (N_3362,N_2928,N_2583);
and U3363 (N_3363,N_2856,N_2687);
nand U3364 (N_3364,N_2805,N_2710);
and U3365 (N_3365,N_2833,N_2564);
and U3366 (N_3366,N_2530,N_2610);
nor U3367 (N_3367,N_2702,N_2932);
nor U3368 (N_3368,N_2717,N_2954);
or U3369 (N_3369,N_2536,N_2903);
nand U3370 (N_3370,N_2822,N_2607);
nor U3371 (N_3371,N_2686,N_2913);
nand U3372 (N_3372,N_2523,N_2859);
xnor U3373 (N_3373,N_2742,N_2696);
and U3374 (N_3374,N_2710,N_2580);
nor U3375 (N_3375,N_2615,N_2980);
nand U3376 (N_3376,N_2800,N_2813);
xnor U3377 (N_3377,N_2667,N_2827);
nor U3378 (N_3378,N_2516,N_2584);
nor U3379 (N_3379,N_2883,N_2717);
or U3380 (N_3380,N_2569,N_2874);
xor U3381 (N_3381,N_2562,N_2577);
nor U3382 (N_3382,N_2810,N_2744);
nor U3383 (N_3383,N_2801,N_2600);
nor U3384 (N_3384,N_2947,N_2994);
nor U3385 (N_3385,N_2684,N_2838);
or U3386 (N_3386,N_2743,N_2858);
nand U3387 (N_3387,N_2548,N_2568);
nand U3388 (N_3388,N_2655,N_2900);
nand U3389 (N_3389,N_2980,N_2691);
nor U3390 (N_3390,N_2965,N_2785);
nor U3391 (N_3391,N_2824,N_2616);
or U3392 (N_3392,N_2583,N_2975);
and U3393 (N_3393,N_2527,N_2904);
nor U3394 (N_3394,N_2971,N_2993);
nor U3395 (N_3395,N_2650,N_2611);
nand U3396 (N_3396,N_2898,N_2944);
and U3397 (N_3397,N_2635,N_2543);
or U3398 (N_3398,N_2595,N_2745);
nor U3399 (N_3399,N_2875,N_2554);
nor U3400 (N_3400,N_2862,N_2869);
nor U3401 (N_3401,N_2854,N_2924);
and U3402 (N_3402,N_2706,N_2906);
and U3403 (N_3403,N_2849,N_2735);
and U3404 (N_3404,N_2539,N_2884);
nor U3405 (N_3405,N_2725,N_2596);
nand U3406 (N_3406,N_2987,N_2751);
nand U3407 (N_3407,N_2849,N_2700);
nor U3408 (N_3408,N_2640,N_2989);
nand U3409 (N_3409,N_2706,N_2784);
or U3410 (N_3410,N_2691,N_2587);
or U3411 (N_3411,N_2505,N_2941);
xnor U3412 (N_3412,N_2602,N_2522);
nand U3413 (N_3413,N_2651,N_2907);
and U3414 (N_3414,N_2633,N_2834);
nor U3415 (N_3415,N_2663,N_2636);
or U3416 (N_3416,N_2550,N_2714);
nor U3417 (N_3417,N_2896,N_2852);
nor U3418 (N_3418,N_2807,N_2965);
xnor U3419 (N_3419,N_2765,N_2638);
nor U3420 (N_3420,N_2883,N_2626);
xnor U3421 (N_3421,N_2559,N_2524);
xnor U3422 (N_3422,N_2762,N_2744);
nand U3423 (N_3423,N_2750,N_2716);
xor U3424 (N_3424,N_2608,N_2553);
and U3425 (N_3425,N_2511,N_2767);
or U3426 (N_3426,N_2558,N_2749);
nor U3427 (N_3427,N_2509,N_2928);
nor U3428 (N_3428,N_2573,N_2587);
xor U3429 (N_3429,N_2614,N_2574);
or U3430 (N_3430,N_2687,N_2776);
and U3431 (N_3431,N_2920,N_2507);
nand U3432 (N_3432,N_2847,N_2552);
nand U3433 (N_3433,N_2893,N_2844);
xor U3434 (N_3434,N_2515,N_2932);
xnor U3435 (N_3435,N_2601,N_2636);
nor U3436 (N_3436,N_2875,N_2876);
nand U3437 (N_3437,N_2805,N_2718);
or U3438 (N_3438,N_2628,N_2593);
nand U3439 (N_3439,N_2890,N_2898);
nand U3440 (N_3440,N_2738,N_2827);
nor U3441 (N_3441,N_2863,N_2970);
nand U3442 (N_3442,N_2919,N_2780);
xor U3443 (N_3443,N_2580,N_2509);
or U3444 (N_3444,N_2711,N_2972);
xor U3445 (N_3445,N_2863,N_2781);
nand U3446 (N_3446,N_2646,N_2881);
and U3447 (N_3447,N_2729,N_2754);
nor U3448 (N_3448,N_2908,N_2555);
and U3449 (N_3449,N_2544,N_2577);
xnor U3450 (N_3450,N_2658,N_2801);
nor U3451 (N_3451,N_2943,N_2773);
nor U3452 (N_3452,N_2955,N_2607);
xnor U3453 (N_3453,N_2507,N_2565);
nand U3454 (N_3454,N_2910,N_2971);
xor U3455 (N_3455,N_2869,N_2724);
xor U3456 (N_3456,N_2541,N_2827);
or U3457 (N_3457,N_2879,N_2878);
nor U3458 (N_3458,N_2591,N_2983);
xnor U3459 (N_3459,N_2757,N_2776);
nor U3460 (N_3460,N_2591,N_2964);
nand U3461 (N_3461,N_2945,N_2775);
xnor U3462 (N_3462,N_2907,N_2668);
or U3463 (N_3463,N_2625,N_2856);
nor U3464 (N_3464,N_2555,N_2882);
or U3465 (N_3465,N_2900,N_2878);
nor U3466 (N_3466,N_2788,N_2896);
nor U3467 (N_3467,N_2996,N_2513);
or U3468 (N_3468,N_2932,N_2975);
xor U3469 (N_3469,N_2838,N_2681);
nand U3470 (N_3470,N_2662,N_2688);
nand U3471 (N_3471,N_2603,N_2902);
nand U3472 (N_3472,N_2602,N_2867);
xor U3473 (N_3473,N_2758,N_2866);
nor U3474 (N_3474,N_2792,N_2506);
nand U3475 (N_3475,N_2800,N_2831);
or U3476 (N_3476,N_2687,N_2652);
or U3477 (N_3477,N_2586,N_2630);
or U3478 (N_3478,N_2711,N_2511);
xnor U3479 (N_3479,N_2713,N_2667);
xnor U3480 (N_3480,N_2989,N_2635);
nand U3481 (N_3481,N_2913,N_2610);
and U3482 (N_3482,N_2531,N_2989);
nand U3483 (N_3483,N_2508,N_2897);
and U3484 (N_3484,N_2771,N_2604);
and U3485 (N_3485,N_2969,N_2710);
or U3486 (N_3486,N_2524,N_2884);
xnor U3487 (N_3487,N_2822,N_2659);
nand U3488 (N_3488,N_2911,N_2522);
nor U3489 (N_3489,N_2880,N_2570);
or U3490 (N_3490,N_2525,N_2508);
xor U3491 (N_3491,N_2701,N_2881);
and U3492 (N_3492,N_2980,N_2745);
or U3493 (N_3493,N_2783,N_2650);
nor U3494 (N_3494,N_2730,N_2882);
nand U3495 (N_3495,N_2780,N_2553);
and U3496 (N_3496,N_2763,N_2927);
nor U3497 (N_3497,N_2901,N_2884);
nor U3498 (N_3498,N_2965,N_2532);
or U3499 (N_3499,N_2856,N_2788);
nand U3500 (N_3500,N_3482,N_3347);
xnor U3501 (N_3501,N_3226,N_3216);
nand U3502 (N_3502,N_3139,N_3210);
and U3503 (N_3503,N_3477,N_3228);
or U3504 (N_3504,N_3293,N_3271);
nand U3505 (N_3505,N_3042,N_3007);
nand U3506 (N_3506,N_3140,N_3300);
and U3507 (N_3507,N_3261,N_3028);
xor U3508 (N_3508,N_3481,N_3315);
nor U3509 (N_3509,N_3108,N_3051);
xor U3510 (N_3510,N_3471,N_3033);
or U3511 (N_3511,N_3229,N_3157);
xnor U3512 (N_3512,N_3298,N_3381);
nand U3513 (N_3513,N_3379,N_3038);
or U3514 (N_3514,N_3434,N_3318);
xor U3515 (N_3515,N_3333,N_3013);
and U3516 (N_3516,N_3212,N_3225);
nand U3517 (N_3517,N_3485,N_3101);
nand U3518 (N_3518,N_3187,N_3198);
or U3519 (N_3519,N_3325,N_3359);
and U3520 (N_3520,N_3159,N_3001);
xor U3521 (N_3521,N_3447,N_3369);
xnor U3522 (N_3522,N_3155,N_3282);
and U3523 (N_3523,N_3441,N_3009);
nand U3524 (N_3524,N_3150,N_3256);
xor U3525 (N_3525,N_3121,N_3064);
xor U3526 (N_3526,N_3113,N_3094);
or U3527 (N_3527,N_3415,N_3400);
nor U3528 (N_3528,N_3248,N_3492);
or U3529 (N_3529,N_3107,N_3370);
nor U3530 (N_3530,N_3397,N_3403);
xnor U3531 (N_3531,N_3326,N_3346);
nor U3532 (N_3532,N_3382,N_3204);
xnor U3533 (N_3533,N_3221,N_3392);
and U3534 (N_3534,N_3025,N_3335);
nand U3535 (N_3535,N_3254,N_3024);
nand U3536 (N_3536,N_3371,N_3448);
nor U3537 (N_3537,N_3132,N_3004);
nor U3538 (N_3538,N_3037,N_3092);
xor U3539 (N_3539,N_3294,N_3044);
xor U3540 (N_3540,N_3016,N_3205);
or U3541 (N_3541,N_3106,N_3241);
nor U3542 (N_3542,N_3428,N_3242);
and U3543 (N_3543,N_3366,N_3461);
nand U3544 (N_3544,N_3322,N_3022);
xnor U3545 (N_3545,N_3329,N_3170);
xor U3546 (N_3546,N_3003,N_3267);
xnor U3547 (N_3547,N_3088,N_3115);
and U3548 (N_3548,N_3249,N_3017);
xor U3549 (N_3549,N_3144,N_3006);
or U3550 (N_3550,N_3130,N_3474);
nand U3551 (N_3551,N_3288,N_3046);
nand U3552 (N_3552,N_3137,N_3260);
xnor U3553 (N_3553,N_3060,N_3099);
and U3554 (N_3554,N_3194,N_3465);
or U3555 (N_3555,N_3436,N_3026);
xnor U3556 (N_3556,N_3074,N_3036);
nand U3557 (N_3557,N_3151,N_3272);
and U3558 (N_3558,N_3311,N_3011);
or U3559 (N_3559,N_3426,N_3207);
nand U3560 (N_3560,N_3405,N_3131);
xnor U3561 (N_3561,N_3160,N_3197);
xnor U3562 (N_3562,N_3384,N_3427);
nor U3563 (N_3563,N_3123,N_3062);
xnor U3564 (N_3564,N_3320,N_3336);
nand U3565 (N_3565,N_3182,N_3255);
or U3566 (N_3566,N_3104,N_3148);
xnor U3567 (N_3567,N_3245,N_3443);
nor U3568 (N_3568,N_3488,N_3065);
or U3569 (N_3569,N_3296,N_3068);
nor U3570 (N_3570,N_3253,N_3040);
xnor U3571 (N_3571,N_3277,N_3142);
nand U3572 (N_3572,N_3352,N_3124);
nand U3573 (N_3573,N_3444,N_3240);
nand U3574 (N_3574,N_3478,N_3475);
and U3575 (N_3575,N_3164,N_3334);
nor U3576 (N_3576,N_3184,N_3079);
or U3577 (N_3577,N_3105,N_3045);
or U3578 (N_3578,N_3072,N_3401);
or U3579 (N_3579,N_3189,N_3224);
or U3580 (N_3580,N_3243,N_3283);
or U3581 (N_3581,N_3353,N_3377);
xnor U3582 (N_3582,N_3383,N_3070);
or U3583 (N_3583,N_3156,N_3457);
and U3584 (N_3584,N_3404,N_3454);
and U3585 (N_3585,N_3010,N_3368);
and U3586 (N_3586,N_3112,N_3432);
xnor U3587 (N_3587,N_3201,N_3423);
or U3588 (N_3588,N_3129,N_3056);
nor U3589 (N_3589,N_3470,N_3348);
nand U3590 (N_3590,N_3494,N_3340);
or U3591 (N_3591,N_3174,N_3133);
or U3592 (N_3592,N_3186,N_3458);
xor U3593 (N_3593,N_3324,N_3331);
xor U3594 (N_3594,N_3417,N_3493);
and U3595 (N_3595,N_3191,N_3274);
nor U3596 (N_3596,N_3053,N_3034);
and U3597 (N_3597,N_3161,N_3192);
nor U3598 (N_3598,N_3175,N_3143);
or U3599 (N_3599,N_3455,N_3118);
xnor U3600 (N_3600,N_3128,N_3418);
xor U3601 (N_3601,N_3306,N_3414);
xor U3602 (N_3602,N_3343,N_3220);
nor U3603 (N_3603,N_3301,N_3453);
nor U3604 (N_3604,N_3213,N_3179);
and U3605 (N_3605,N_3378,N_3399);
nand U3606 (N_3606,N_3289,N_3354);
nand U3607 (N_3607,N_3167,N_3409);
nand U3608 (N_3608,N_3251,N_3049);
or U3609 (N_3609,N_3077,N_3181);
and U3610 (N_3610,N_3290,N_3349);
nand U3611 (N_3611,N_3116,N_3019);
and U3612 (N_3612,N_3279,N_3075);
nand U3613 (N_3613,N_3345,N_3421);
nor U3614 (N_3614,N_3171,N_3223);
xor U3615 (N_3615,N_3364,N_3412);
or U3616 (N_3616,N_3374,N_3232);
or U3617 (N_3617,N_3424,N_3015);
or U3618 (N_3618,N_3193,N_3269);
or U3619 (N_3619,N_3027,N_3310);
nor U3620 (N_3620,N_3206,N_3375);
nor U3621 (N_3621,N_3141,N_3163);
or U3622 (N_3622,N_3136,N_3168);
nand U3623 (N_3623,N_3446,N_3158);
or U3624 (N_3624,N_3257,N_3278);
nand U3625 (N_3625,N_3052,N_3273);
nand U3626 (N_3626,N_3263,N_3199);
nor U3627 (N_3627,N_3433,N_3351);
xor U3628 (N_3628,N_3445,N_3307);
or U3629 (N_3629,N_3183,N_3344);
nor U3630 (N_3630,N_3236,N_3238);
nand U3631 (N_3631,N_3073,N_3196);
or U3632 (N_3632,N_3319,N_3373);
and U3633 (N_3633,N_3235,N_3147);
nand U3634 (N_3634,N_3048,N_3096);
or U3635 (N_3635,N_3110,N_3005);
and U3636 (N_3636,N_3219,N_3266);
xnor U3637 (N_3637,N_3416,N_3063);
nand U3638 (N_3638,N_3087,N_3463);
xor U3639 (N_3639,N_3165,N_3419);
nand U3640 (N_3640,N_3258,N_3252);
or U3641 (N_3641,N_3084,N_3203);
nor U3642 (N_3642,N_3327,N_3050);
xor U3643 (N_3643,N_3332,N_3102);
xnor U3644 (N_3644,N_3173,N_3291);
nor U3645 (N_3645,N_3080,N_3385);
or U3646 (N_3646,N_3398,N_3341);
and U3647 (N_3647,N_3372,N_3451);
or U3648 (N_3648,N_3227,N_3422);
and U3649 (N_3649,N_3083,N_3029);
and U3650 (N_3650,N_3314,N_3406);
or U3651 (N_3651,N_3305,N_3286);
nor U3652 (N_3652,N_3281,N_3246);
nor U3653 (N_3653,N_3280,N_3337);
and U3654 (N_3654,N_3365,N_3211);
or U3655 (N_3655,N_3247,N_3276);
or U3656 (N_3656,N_3127,N_3302);
or U3657 (N_3657,N_3218,N_3450);
and U3658 (N_3658,N_3390,N_3407);
and U3659 (N_3659,N_3466,N_3497);
xor U3660 (N_3660,N_3032,N_3097);
or U3661 (N_3661,N_3389,N_3002);
nor U3662 (N_3662,N_3393,N_3035);
xnor U3663 (N_3663,N_3120,N_3103);
or U3664 (N_3664,N_3330,N_3442);
xor U3665 (N_3665,N_3185,N_3057);
or U3666 (N_3666,N_3178,N_3491);
or U3667 (N_3667,N_3264,N_3012);
xor U3668 (N_3668,N_3386,N_3230);
or U3669 (N_3669,N_3388,N_3486);
or U3670 (N_3670,N_3100,N_3259);
and U3671 (N_3671,N_3313,N_3287);
xor U3672 (N_3672,N_3410,N_3039);
and U3673 (N_3673,N_3489,N_3483);
xor U3674 (N_3674,N_3089,N_3146);
nor U3675 (N_3675,N_3217,N_3047);
xnor U3676 (N_3676,N_3316,N_3295);
xor U3677 (N_3677,N_3166,N_3473);
and U3678 (N_3678,N_3109,N_3358);
and U3679 (N_3679,N_3233,N_3119);
and U3680 (N_3680,N_3149,N_3195);
nor U3681 (N_3681,N_3342,N_3317);
nand U3682 (N_3682,N_3081,N_3209);
and U3683 (N_3683,N_3043,N_3402);
or U3684 (N_3684,N_3408,N_3425);
nor U3685 (N_3685,N_3055,N_3299);
or U3686 (N_3686,N_3117,N_3188);
and U3687 (N_3687,N_3304,N_3438);
nand U3688 (N_3688,N_3200,N_3265);
and U3689 (N_3689,N_3479,N_3239);
nor U3690 (N_3690,N_3145,N_3495);
and U3691 (N_3691,N_3098,N_3361);
or U3692 (N_3692,N_3122,N_3135);
nor U3693 (N_3693,N_3476,N_3071);
nand U3694 (N_3694,N_3284,N_3484);
or U3695 (N_3695,N_3067,N_3312);
and U3696 (N_3696,N_3008,N_3153);
nor U3697 (N_3697,N_3054,N_3222);
nand U3698 (N_3698,N_3376,N_3059);
xnor U3699 (N_3699,N_3360,N_3462);
and U3700 (N_3700,N_3321,N_3095);
or U3701 (N_3701,N_3268,N_3134);
and U3702 (N_3702,N_3125,N_3328);
xor U3703 (N_3703,N_3262,N_3000);
nand U3704 (N_3704,N_3297,N_3270);
nor U3705 (N_3705,N_3190,N_3114);
and U3706 (N_3706,N_3357,N_3021);
xnor U3707 (N_3707,N_3435,N_3339);
and U3708 (N_3708,N_3411,N_3176);
or U3709 (N_3709,N_3367,N_3472);
and U3710 (N_3710,N_3468,N_3177);
and U3711 (N_3711,N_3093,N_3152);
and U3712 (N_3712,N_3380,N_3387);
xnor U3713 (N_3713,N_3061,N_3469);
and U3714 (N_3714,N_3449,N_3126);
nor U3715 (N_3715,N_3066,N_3413);
nor U3716 (N_3716,N_3430,N_3308);
and U3717 (N_3717,N_3496,N_3459);
or U3718 (N_3718,N_3091,N_3020);
xnor U3719 (N_3719,N_3420,N_3498);
or U3720 (N_3720,N_3292,N_3480);
nand U3721 (N_3721,N_3309,N_3464);
xor U3722 (N_3722,N_3082,N_3323);
nand U3723 (N_3723,N_3439,N_3041);
nand U3724 (N_3724,N_3078,N_3391);
or U3725 (N_3725,N_3394,N_3172);
nand U3726 (N_3726,N_3499,N_3303);
nor U3727 (N_3727,N_3154,N_3076);
or U3728 (N_3728,N_3356,N_3069);
xor U3729 (N_3729,N_3169,N_3030);
nand U3730 (N_3730,N_3237,N_3431);
nor U3731 (N_3731,N_3214,N_3396);
nand U3732 (N_3732,N_3014,N_3215);
nand U3733 (N_3733,N_3437,N_3338);
or U3734 (N_3734,N_3085,N_3162);
nor U3735 (N_3735,N_3362,N_3285);
xor U3736 (N_3736,N_3429,N_3031);
and U3737 (N_3737,N_3058,N_3180);
xnor U3738 (N_3738,N_3440,N_3467);
or U3739 (N_3739,N_3460,N_3452);
xnor U3740 (N_3740,N_3086,N_3456);
and U3741 (N_3741,N_3490,N_3018);
or U3742 (N_3742,N_3355,N_3363);
nand U3743 (N_3743,N_3275,N_3090);
nor U3744 (N_3744,N_3111,N_3023);
and U3745 (N_3745,N_3244,N_3202);
xor U3746 (N_3746,N_3234,N_3208);
xor U3747 (N_3747,N_3138,N_3250);
nand U3748 (N_3748,N_3395,N_3231);
nor U3749 (N_3749,N_3487,N_3350);
nor U3750 (N_3750,N_3462,N_3188);
xor U3751 (N_3751,N_3008,N_3461);
xnor U3752 (N_3752,N_3202,N_3100);
and U3753 (N_3753,N_3083,N_3412);
and U3754 (N_3754,N_3182,N_3028);
nand U3755 (N_3755,N_3002,N_3480);
nand U3756 (N_3756,N_3296,N_3094);
nand U3757 (N_3757,N_3023,N_3402);
and U3758 (N_3758,N_3235,N_3372);
or U3759 (N_3759,N_3279,N_3358);
and U3760 (N_3760,N_3028,N_3475);
nand U3761 (N_3761,N_3049,N_3425);
and U3762 (N_3762,N_3135,N_3325);
and U3763 (N_3763,N_3133,N_3113);
nor U3764 (N_3764,N_3183,N_3464);
xor U3765 (N_3765,N_3465,N_3411);
nand U3766 (N_3766,N_3362,N_3486);
or U3767 (N_3767,N_3416,N_3101);
and U3768 (N_3768,N_3262,N_3084);
xnor U3769 (N_3769,N_3437,N_3260);
and U3770 (N_3770,N_3062,N_3385);
xor U3771 (N_3771,N_3046,N_3128);
xor U3772 (N_3772,N_3142,N_3174);
xnor U3773 (N_3773,N_3072,N_3000);
and U3774 (N_3774,N_3249,N_3149);
nand U3775 (N_3775,N_3347,N_3185);
xor U3776 (N_3776,N_3102,N_3453);
xor U3777 (N_3777,N_3289,N_3399);
xor U3778 (N_3778,N_3038,N_3497);
and U3779 (N_3779,N_3049,N_3074);
or U3780 (N_3780,N_3166,N_3259);
and U3781 (N_3781,N_3384,N_3012);
nand U3782 (N_3782,N_3159,N_3346);
nand U3783 (N_3783,N_3299,N_3406);
and U3784 (N_3784,N_3127,N_3263);
nand U3785 (N_3785,N_3324,N_3036);
nor U3786 (N_3786,N_3228,N_3162);
nor U3787 (N_3787,N_3254,N_3489);
xnor U3788 (N_3788,N_3062,N_3368);
or U3789 (N_3789,N_3428,N_3088);
and U3790 (N_3790,N_3394,N_3212);
nand U3791 (N_3791,N_3064,N_3273);
nand U3792 (N_3792,N_3422,N_3243);
nor U3793 (N_3793,N_3469,N_3256);
or U3794 (N_3794,N_3038,N_3285);
xor U3795 (N_3795,N_3493,N_3356);
nand U3796 (N_3796,N_3271,N_3331);
and U3797 (N_3797,N_3377,N_3350);
nor U3798 (N_3798,N_3106,N_3254);
and U3799 (N_3799,N_3001,N_3077);
nand U3800 (N_3800,N_3372,N_3461);
or U3801 (N_3801,N_3038,N_3330);
nor U3802 (N_3802,N_3390,N_3136);
xnor U3803 (N_3803,N_3129,N_3283);
xor U3804 (N_3804,N_3475,N_3065);
xnor U3805 (N_3805,N_3158,N_3382);
xor U3806 (N_3806,N_3212,N_3399);
nand U3807 (N_3807,N_3328,N_3049);
or U3808 (N_3808,N_3059,N_3064);
nor U3809 (N_3809,N_3493,N_3152);
nand U3810 (N_3810,N_3366,N_3415);
or U3811 (N_3811,N_3026,N_3167);
and U3812 (N_3812,N_3324,N_3364);
xor U3813 (N_3813,N_3279,N_3306);
nand U3814 (N_3814,N_3126,N_3162);
xnor U3815 (N_3815,N_3023,N_3266);
xnor U3816 (N_3816,N_3346,N_3381);
nor U3817 (N_3817,N_3462,N_3029);
xor U3818 (N_3818,N_3203,N_3029);
xor U3819 (N_3819,N_3158,N_3181);
nor U3820 (N_3820,N_3376,N_3329);
xnor U3821 (N_3821,N_3061,N_3185);
nand U3822 (N_3822,N_3023,N_3069);
and U3823 (N_3823,N_3483,N_3335);
nand U3824 (N_3824,N_3239,N_3415);
nor U3825 (N_3825,N_3464,N_3256);
or U3826 (N_3826,N_3346,N_3130);
nor U3827 (N_3827,N_3218,N_3004);
and U3828 (N_3828,N_3107,N_3146);
and U3829 (N_3829,N_3217,N_3174);
nor U3830 (N_3830,N_3107,N_3065);
nor U3831 (N_3831,N_3487,N_3432);
xnor U3832 (N_3832,N_3492,N_3491);
nand U3833 (N_3833,N_3059,N_3057);
and U3834 (N_3834,N_3435,N_3277);
or U3835 (N_3835,N_3170,N_3102);
xnor U3836 (N_3836,N_3476,N_3379);
nand U3837 (N_3837,N_3466,N_3331);
nor U3838 (N_3838,N_3241,N_3378);
and U3839 (N_3839,N_3239,N_3190);
xor U3840 (N_3840,N_3397,N_3123);
xor U3841 (N_3841,N_3131,N_3439);
and U3842 (N_3842,N_3489,N_3488);
or U3843 (N_3843,N_3139,N_3354);
nand U3844 (N_3844,N_3100,N_3362);
xnor U3845 (N_3845,N_3343,N_3150);
or U3846 (N_3846,N_3380,N_3098);
nand U3847 (N_3847,N_3133,N_3381);
nor U3848 (N_3848,N_3041,N_3372);
or U3849 (N_3849,N_3007,N_3206);
nor U3850 (N_3850,N_3043,N_3124);
nor U3851 (N_3851,N_3475,N_3231);
nor U3852 (N_3852,N_3234,N_3323);
nand U3853 (N_3853,N_3484,N_3039);
or U3854 (N_3854,N_3282,N_3321);
nand U3855 (N_3855,N_3001,N_3370);
nor U3856 (N_3856,N_3135,N_3499);
xnor U3857 (N_3857,N_3168,N_3096);
or U3858 (N_3858,N_3459,N_3234);
nor U3859 (N_3859,N_3479,N_3426);
nand U3860 (N_3860,N_3466,N_3324);
and U3861 (N_3861,N_3085,N_3486);
and U3862 (N_3862,N_3152,N_3102);
or U3863 (N_3863,N_3464,N_3476);
or U3864 (N_3864,N_3037,N_3224);
or U3865 (N_3865,N_3210,N_3478);
xnor U3866 (N_3866,N_3463,N_3138);
nand U3867 (N_3867,N_3450,N_3375);
nand U3868 (N_3868,N_3292,N_3417);
or U3869 (N_3869,N_3102,N_3083);
nor U3870 (N_3870,N_3176,N_3329);
or U3871 (N_3871,N_3378,N_3452);
and U3872 (N_3872,N_3223,N_3101);
nand U3873 (N_3873,N_3148,N_3156);
and U3874 (N_3874,N_3178,N_3055);
nand U3875 (N_3875,N_3452,N_3070);
nand U3876 (N_3876,N_3306,N_3427);
or U3877 (N_3877,N_3194,N_3432);
nand U3878 (N_3878,N_3001,N_3097);
or U3879 (N_3879,N_3178,N_3329);
or U3880 (N_3880,N_3200,N_3208);
and U3881 (N_3881,N_3314,N_3070);
or U3882 (N_3882,N_3421,N_3079);
or U3883 (N_3883,N_3254,N_3039);
nand U3884 (N_3884,N_3240,N_3057);
xnor U3885 (N_3885,N_3009,N_3477);
and U3886 (N_3886,N_3019,N_3077);
nor U3887 (N_3887,N_3344,N_3295);
and U3888 (N_3888,N_3426,N_3113);
nand U3889 (N_3889,N_3239,N_3278);
and U3890 (N_3890,N_3326,N_3297);
nand U3891 (N_3891,N_3344,N_3134);
nor U3892 (N_3892,N_3167,N_3407);
nor U3893 (N_3893,N_3083,N_3322);
nand U3894 (N_3894,N_3402,N_3005);
nand U3895 (N_3895,N_3213,N_3192);
nor U3896 (N_3896,N_3135,N_3408);
nor U3897 (N_3897,N_3185,N_3116);
or U3898 (N_3898,N_3286,N_3311);
or U3899 (N_3899,N_3151,N_3295);
nand U3900 (N_3900,N_3015,N_3308);
or U3901 (N_3901,N_3009,N_3450);
xnor U3902 (N_3902,N_3106,N_3393);
xor U3903 (N_3903,N_3446,N_3322);
or U3904 (N_3904,N_3050,N_3011);
nand U3905 (N_3905,N_3245,N_3135);
or U3906 (N_3906,N_3394,N_3303);
and U3907 (N_3907,N_3345,N_3174);
xnor U3908 (N_3908,N_3036,N_3418);
and U3909 (N_3909,N_3271,N_3269);
and U3910 (N_3910,N_3434,N_3479);
xor U3911 (N_3911,N_3378,N_3385);
nand U3912 (N_3912,N_3043,N_3206);
and U3913 (N_3913,N_3220,N_3203);
nand U3914 (N_3914,N_3104,N_3467);
nor U3915 (N_3915,N_3002,N_3341);
and U3916 (N_3916,N_3040,N_3098);
and U3917 (N_3917,N_3058,N_3177);
nand U3918 (N_3918,N_3330,N_3248);
xor U3919 (N_3919,N_3031,N_3064);
nor U3920 (N_3920,N_3286,N_3149);
or U3921 (N_3921,N_3415,N_3422);
nor U3922 (N_3922,N_3307,N_3259);
or U3923 (N_3923,N_3308,N_3371);
and U3924 (N_3924,N_3475,N_3175);
and U3925 (N_3925,N_3351,N_3297);
or U3926 (N_3926,N_3154,N_3339);
or U3927 (N_3927,N_3372,N_3355);
nor U3928 (N_3928,N_3180,N_3234);
nand U3929 (N_3929,N_3301,N_3305);
and U3930 (N_3930,N_3193,N_3383);
xor U3931 (N_3931,N_3008,N_3444);
or U3932 (N_3932,N_3048,N_3487);
xor U3933 (N_3933,N_3056,N_3447);
xnor U3934 (N_3934,N_3128,N_3290);
or U3935 (N_3935,N_3457,N_3351);
nor U3936 (N_3936,N_3269,N_3320);
and U3937 (N_3937,N_3125,N_3205);
nand U3938 (N_3938,N_3231,N_3038);
or U3939 (N_3939,N_3305,N_3410);
nand U3940 (N_3940,N_3265,N_3308);
and U3941 (N_3941,N_3300,N_3397);
and U3942 (N_3942,N_3158,N_3140);
or U3943 (N_3943,N_3298,N_3146);
nor U3944 (N_3944,N_3183,N_3272);
nand U3945 (N_3945,N_3090,N_3228);
and U3946 (N_3946,N_3435,N_3216);
or U3947 (N_3947,N_3450,N_3257);
or U3948 (N_3948,N_3480,N_3288);
nor U3949 (N_3949,N_3422,N_3066);
and U3950 (N_3950,N_3488,N_3002);
nand U3951 (N_3951,N_3268,N_3409);
or U3952 (N_3952,N_3367,N_3233);
xnor U3953 (N_3953,N_3014,N_3221);
nor U3954 (N_3954,N_3423,N_3114);
or U3955 (N_3955,N_3295,N_3300);
or U3956 (N_3956,N_3250,N_3113);
and U3957 (N_3957,N_3092,N_3061);
and U3958 (N_3958,N_3048,N_3118);
nand U3959 (N_3959,N_3340,N_3280);
xnor U3960 (N_3960,N_3445,N_3278);
xor U3961 (N_3961,N_3101,N_3392);
or U3962 (N_3962,N_3486,N_3466);
or U3963 (N_3963,N_3083,N_3461);
nor U3964 (N_3964,N_3130,N_3222);
and U3965 (N_3965,N_3203,N_3139);
nand U3966 (N_3966,N_3351,N_3273);
or U3967 (N_3967,N_3296,N_3166);
or U3968 (N_3968,N_3457,N_3170);
nor U3969 (N_3969,N_3356,N_3245);
or U3970 (N_3970,N_3004,N_3488);
xnor U3971 (N_3971,N_3381,N_3460);
nor U3972 (N_3972,N_3419,N_3075);
and U3973 (N_3973,N_3090,N_3305);
xnor U3974 (N_3974,N_3363,N_3155);
nand U3975 (N_3975,N_3030,N_3111);
nor U3976 (N_3976,N_3247,N_3477);
or U3977 (N_3977,N_3127,N_3499);
and U3978 (N_3978,N_3320,N_3412);
nor U3979 (N_3979,N_3222,N_3126);
or U3980 (N_3980,N_3238,N_3454);
xor U3981 (N_3981,N_3167,N_3344);
and U3982 (N_3982,N_3309,N_3072);
and U3983 (N_3983,N_3106,N_3407);
xor U3984 (N_3984,N_3434,N_3250);
nand U3985 (N_3985,N_3006,N_3343);
or U3986 (N_3986,N_3181,N_3459);
xor U3987 (N_3987,N_3434,N_3212);
or U3988 (N_3988,N_3220,N_3001);
nor U3989 (N_3989,N_3148,N_3375);
nand U3990 (N_3990,N_3101,N_3206);
xor U3991 (N_3991,N_3428,N_3269);
xnor U3992 (N_3992,N_3234,N_3193);
nor U3993 (N_3993,N_3300,N_3469);
xor U3994 (N_3994,N_3214,N_3088);
xnor U3995 (N_3995,N_3164,N_3111);
or U3996 (N_3996,N_3086,N_3471);
or U3997 (N_3997,N_3392,N_3351);
nand U3998 (N_3998,N_3274,N_3346);
nor U3999 (N_3999,N_3478,N_3135);
or U4000 (N_4000,N_3927,N_3545);
xor U4001 (N_4001,N_3577,N_3540);
nor U4002 (N_4002,N_3961,N_3669);
nor U4003 (N_4003,N_3804,N_3680);
and U4004 (N_4004,N_3969,N_3675);
or U4005 (N_4005,N_3596,N_3589);
nand U4006 (N_4006,N_3661,N_3611);
nand U4007 (N_4007,N_3859,N_3614);
nand U4008 (N_4008,N_3549,N_3560);
nand U4009 (N_4009,N_3619,N_3563);
and U4010 (N_4010,N_3728,N_3706);
nand U4011 (N_4011,N_3871,N_3908);
nand U4012 (N_4012,N_3801,N_3509);
and U4013 (N_4013,N_3515,N_3630);
nor U4014 (N_4014,N_3530,N_3655);
nor U4015 (N_4015,N_3808,N_3943);
and U4016 (N_4016,N_3602,N_3899);
or U4017 (N_4017,N_3867,N_3699);
and U4018 (N_4018,N_3725,N_3701);
or U4019 (N_4019,N_3552,N_3894);
and U4020 (N_4020,N_3994,N_3723);
and U4021 (N_4021,N_3637,N_3623);
nand U4022 (N_4022,N_3930,N_3650);
nand U4023 (N_4023,N_3853,N_3874);
nor U4024 (N_4024,N_3793,N_3795);
nor U4025 (N_4025,N_3638,N_3968);
and U4026 (N_4026,N_3852,N_3666);
or U4027 (N_4027,N_3733,N_3771);
xnor U4028 (N_4028,N_3644,N_3950);
and U4029 (N_4029,N_3615,N_3812);
nor U4030 (N_4030,N_3883,N_3700);
xor U4031 (N_4031,N_3869,N_3902);
and U4032 (N_4032,N_3624,N_3963);
nand U4033 (N_4033,N_3708,N_3579);
xnor U4034 (N_4034,N_3752,N_3717);
xnor U4035 (N_4035,N_3756,N_3572);
nor U4036 (N_4036,N_3870,N_3649);
or U4037 (N_4037,N_3999,N_3794);
and U4038 (N_4038,N_3960,N_3763);
and U4039 (N_4039,N_3778,N_3993);
or U4040 (N_4040,N_3974,N_3764);
and U4041 (N_4041,N_3553,N_3651);
nand U4042 (N_4042,N_3737,N_3951);
or U4043 (N_4043,N_3762,N_3842);
nand U4044 (N_4044,N_3525,N_3674);
or U4045 (N_4045,N_3513,N_3645);
nand U4046 (N_4046,N_3508,N_3582);
nand U4047 (N_4047,N_3814,N_3510);
nand U4048 (N_4048,N_3886,N_3914);
nand U4049 (N_4049,N_3940,N_3526);
or U4050 (N_4050,N_3964,N_3824);
or U4051 (N_4051,N_3879,N_3512);
or U4052 (N_4052,N_3988,N_3556);
nor U4053 (N_4053,N_3939,N_3562);
nor U4054 (N_4054,N_3523,N_3640);
and U4055 (N_4055,N_3505,N_3709);
nand U4056 (N_4056,N_3858,N_3621);
xnor U4057 (N_4057,N_3738,N_3838);
or U4058 (N_4058,N_3566,N_3903);
xor U4059 (N_4059,N_3888,N_3834);
nand U4060 (N_4060,N_3885,N_3765);
xnor U4061 (N_4061,N_3920,N_3750);
nand U4062 (N_4062,N_3807,N_3607);
nor U4063 (N_4063,N_3696,N_3681);
nand U4064 (N_4064,N_3689,N_3997);
nor U4065 (N_4065,N_3802,N_3833);
nor U4066 (N_4066,N_3783,N_3517);
and U4067 (N_4067,N_3925,N_3601);
or U4068 (N_4068,N_3845,N_3891);
xnor U4069 (N_4069,N_3503,N_3975);
or U4070 (N_4070,N_3539,N_3736);
and U4071 (N_4071,N_3500,N_3551);
nor U4072 (N_4072,N_3797,N_3606);
xor U4073 (N_4073,N_3986,N_3718);
nand U4074 (N_4074,N_3815,N_3881);
or U4075 (N_4075,N_3840,N_3904);
and U4076 (N_4076,N_3643,N_3864);
xnor U4077 (N_4077,N_3720,N_3844);
nand U4078 (N_4078,N_3861,N_3622);
nor U4079 (N_4079,N_3537,N_3766);
or U4080 (N_4080,N_3590,N_3803);
nand U4081 (N_4081,N_3768,N_3895);
nand U4082 (N_4082,N_3954,N_3825);
nand U4083 (N_4083,N_3584,N_3985);
nor U4084 (N_4084,N_3729,N_3998);
nand U4085 (N_4085,N_3683,N_3702);
or U4086 (N_4086,N_3912,N_3679);
xor U4087 (N_4087,N_3828,N_3713);
xnor U4088 (N_4088,N_3850,N_3820);
or U4089 (N_4089,N_3610,N_3647);
nand U4090 (N_4090,N_3773,N_3529);
nor U4091 (N_4091,N_3664,N_3976);
xor U4092 (N_4092,N_3555,N_3955);
or U4093 (N_4093,N_3693,N_3944);
and U4094 (N_4094,N_3910,N_3884);
xor U4095 (N_4095,N_3520,N_3984);
nand U4096 (N_4096,N_3848,N_3660);
nand U4097 (N_4097,N_3755,N_3548);
nand U4098 (N_4098,N_3957,N_3897);
nor U4099 (N_4099,N_3535,N_3913);
or U4100 (N_4100,N_3550,N_3782);
and U4101 (N_4101,N_3703,N_3949);
or U4102 (N_4102,N_3712,N_3599);
xor U4103 (N_4103,N_3758,N_3924);
nor U4104 (N_4104,N_3597,N_3594);
nand U4105 (N_4105,N_3633,N_3978);
and U4106 (N_4106,N_3936,N_3627);
and U4107 (N_4107,N_3831,N_3952);
and U4108 (N_4108,N_3860,N_3889);
xor U4109 (N_4109,N_3996,N_3629);
or U4110 (N_4110,N_3800,N_3668);
or U4111 (N_4111,N_3928,N_3559);
and U4112 (N_4112,N_3715,N_3934);
nor U4113 (N_4113,N_3571,N_3697);
xor U4114 (N_4114,N_3543,N_3835);
and U4115 (N_4115,N_3598,N_3608);
xnor U4116 (N_4116,N_3719,N_3777);
and U4117 (N_4117,N_3603,N_3652);
or U4118 (N_4118,N_3785,N_3742);
nand U4119 (N_4119,N_3781,N_3747);
and U4120 (N_4120,N_3536,N_3810);
nor U4121 (N_4121,N_3727,N_3648);
or U4122 (N_4122,N_3625,N_3847);
or U4123 (N_4123,N_3732,N_3816);
nand U4124 (N_4124,N_3977,N_3938);
nand U4125 (N_4125,N_3740,N_3919);
or U4126 (N_4126,N_3635,N_3780);
nand U4127 (N_4127,N_3929,N_3704);
or U4128 (N_4128,N_3521,N_3923);
nand U4129 (N_4129,N_3767,N_3887);
and U4130 (N_4130,N_3665,N_3827);
nand U4131 (N_4131,N_3741,N_3863);
and U4132 (N_4132,N_3933,N_3915);
or U4133 (N_4133,N_3872,N_3779);
or U4134 (N_4134,N_3528,N_3605);
nand U4135 (N_4135,N_3504,N_3796);
and U4136 (N_4136,N_3724,N_3965);
xnor U4137 (N_4137,N_3714,N_3642);
nand U4138 (N_4138,N_3770,N_3743);
or U4139 (N_4139,N_3730,N_3685);
and U4140 (N_4140,N_3544,N_3855);
and U4141 (N_4141,N_3739,N_3811);
and U4142 (N_4142,N_3854,N_3684);
or U4143 (N_4143,N_3832,N_3942);
xor U4144 (N_4144,N_3878,N_3524);
and U4145 (N_4145,N_3673,N_3971);
xor U4146 (N_4146,N_3917,N_3532);
nor U4147 (N_4147,N_3641,N_3757);
xor U4148 (N_4148,N_3569,N_3798);
xnor U4149 (N_4149,N_3538,N_3926);
and U4150 (N_4150,N_3901,N_3722);
or U4151 (N_4151,N_3754,N_3829);
or U4152 (N_4152,N_3973,N_3995);
or U4153 (N_4153,N_3721,N_3574);
nor U4154 (N_4154,N_3836,N_3561);
nor U4155 (N_4155,N_3578,N_3972);
and U4156 (N_4156,N_3992,N_3937);
nand U4157 (N_4157,N_3711,N_3705);
nand U4158 (N_4158,N_3516,N_3843);
xor U4159 (N_4159,N_3911,N_3690);
or U4160 (N_4160,N_3533,N_3791);
nor U4161 (N_4161,N_3565,N_3900);
xor U4162 (N_4162,N_3753,N_3688);
and U4163 (N_4163,N_3716,N_3837);
xnor U4164 (N_4164,N_3958,N_3892);
nand U4165 (N_4165,N_3857,N_3979);
nor U4166 (N_4166,N_3658,N_3823);
xor U4167 (N_4167,N_3982,N_3822);
or U4168 (N_4168,N_3731,N_3593);
xor U4169 (N_4169,N_3656,N_3662);
nand U4170 (N_4170,N_3698,N_3769);
nand U4171 (N_4171,N_3695,N_3980);
xor U4172 (N_4172,N_3588,N_3626);
and U4173 (N_4173,N_3546,N_3792);
xnor U4174 (N_4174,N_3581,N_3507);
or U4175 (N_4175,N_3941,N_3789);
and U4176 (N_4176,N_3564,N_3896);
nor U4177 (N_4177,N_3672,N_3609);
xor U4178 (N_4178,N_3600,N_3639);
and U4179 (N_4179,N_3511,N_3947);
nor U4180 (N_4180,N_3726,N_3898);
nor U4181 (N_4181,N_3809,N_3568);
xnor U4182 (N_4182,N_3868,N_3787);
nand U4183 (N_4183,N_3873,N_3813);
or U4184 (N_4184,N_3692,N_3922);
and U4185 (N_4185,N_3604,N_3819);
nor U4186 (N_4186,N_3676,N_3667);
and U4187 (N_4187,N_3557,N_3990);
xnor U4188 (N_4188,N_3531,N_3587);
and U4189 (N_4189,N_3636,N_3612);
xnor U4190 (N_4190,N_3786,N_3983);
or U4191 (N_4191,N_3707,N_3772);
nand U4192 (N_4192,N_3585,N_3541);
and U4193 (N_4193,N_3558,N_3547);
nand U4194 (N_4194,N_3966,N_3514);
and U4195 (N_4195,N_3905,N_3646);
or U4196 (N_4196,N_3970,N_3677);
xnor U4197 (N_4197,N_3893,N_3890);
xor U4198 (N_4198,N_3632,N_3776);
and U4199 (N_4199,N_3631,N_3506);
and U4200 (N_4200,N_3788,N_3967);
xnor U4201 (N_4201,N_3959,N_3962);
nor U4202 (N_4202,N_3710,N_3866);
nor U4203 (N_4203,N_3575,N_3554);
nor U4204 (N_4204,N_3775,N_3907);
or U4205 (N_4205,N_3784,N_3989);
xnor U4206 (N_4206,N_3849,N_3906);
nor U4207 (N_4207,N_3931,N_3580);
xor U4208 (N_4208,N_3634,N_3932);
nand U4209 (N_4209,N_3567,N_3851);
nand U4210 (N_4210,N_3527,N_3981);
or U4211 (N_4211,N_3671,N_3501);
xor U4212 (N_4212,N_3876,N_3805);
nor U4213 (N_4213,N_3613,N_3670);
nor U4214 (N_4214,N_3518,N_3691);
and U4215 (N_4215,N_3856,N_3687);
nor U4216 (N_4216,N_3956,N_3790);
or U4217 (N_4217,N_3522,N_3946);
and U4218 (N_4218,N_3534,N_3846);
and U4219 (N_4219,N_3617,N_3774);
nand U4220 (N_4220,N_3502,N_3841);
nor U4221 (N_4221,N_3595,N_3663);
nor U4222 (N_4222,N_3916,N_3576);
or U4223 (N_4223,N_3760,N_3909);
xnor U4224 (N_4224,N_3657,N_3746);
xnor U4225 (N_4225,N_3953,N_3880);
and U4226 (N_4226,N_3694,N_3748);
and U4227 (N_4227,N_3573,N_3751);
nor U4228 (N_4228,N_3653,N_3749);
and U4229 (N_4229,N_3826,N_3877);
nand U4230 (N_4230,N_3945,N_3839);
xor U4231 (N_4231,N_3618,N_3830);
nand U4232 (N_4232,N_3659,N_3682);
nor U4233 (N_4233,N_3821,N_3806);
nor U4234 (N_4234,N_3628,N_3735);
xnor U4235 (N_4235,N_3948,N_3686);
nor U4236 (N_4236,N_3678,N_3654);
or U4237 (N_4237,N_3620,N_3921);
xnor U4238 (N_4238,N_3865,N_3759);
xor U4239 (N_4239,N_3882,N_3570);
xnor U4240 (N_4240,N_3935,N_3817);
xor U4241 (N_4241,N_3862,N_3761);
xor U4242 (N_4242,N_3744,N_3987);
xor U4243 (N_4243,N_3745,N_3519);
xnor U4244 (N_4244,N_3586,N_3818);
and U4245 (N_4245,N_3591,N_3592);
nor U4246 (N_4246,N_3799,N_3918);
nor U4247 (N_4247,N_3583,N_3542);
nand U4248 (N_4248,N_3991,N_3616);
or U4249 (N_4249,N_3734,N_3875);
nor U4250 (N_4250,N_3638,N_3675);
xor U4251 (N_4251,N_3771,N_3721);
and U4252 (N_4252,N_3939,N_3918);
nand U4253 (N_4253,N_3500,N_3680);
nand U4254 (N_4254,N_3640,N_3860);
xnor U4255 (N_4255,N_3627,N_3736);
xor U4256 (N_4256,N_3595,N_3700);
or U4257 (N_4257,N_3989,N_3751);
or U4258 (N_4258,N_3912,N_3954);
nand U4259 (N_4259,N_3541,N_3623);
or U4260 (N_4260,N_3591,N_3772);
nor U4261 (N_4261,N_3870,N_3953);
or U4262 (N_4262,N_3540,N_3845);
xnor U4263 (N_4263,N_3521,N_3889);
xor U4264 (N_4264,N_3575,N_3876);
and U4265 (N_4265,N_3717,N_3631);
xor U4266 (N_4266,N_3550,N_3985);
nor U4267 (N_4267,N_3899,N_3515);
xnor U4268 (N_4268,N_3900,N_3991);
xor U4269 (N_4269,N_3670,N_3969);
nor U4270 (N_4270,N_3985,N_3872);
xnor U4271 (N_4271,N_3745,N_3888);
and U4272 (N_4272,N_3770,N_3986);
and U4273 (N_4273,N_3993,N_3541);
and U4274 (N_4274,N_3886,N_3702);
or U4275 (N_4275,N_3645,N_3921);
nor U4276 (N_4276,N_3715,N_3983);
nor U4277 (N_4277,N_3789,N_3681);
nor U4278 (N_4278,N_3630,N_3781);
nor U4279 (N_4279,N_3517,N_3963);
or U4280 (N_4280,N_3960,N_3989);
xnor U4281 (N_4281,N_3689,N_3513);
nand U4282 (N_4282,N_3937,N_3890);
nand U4283 (N_4283,N_3907,N_3812);
nand U4284 (N_4284,N_3654,N_3659);
nor U4285 (N_4285,N_3625,N_3636);
nor U4286 (N_4286,N_3598,N_3770);
and U4287 (N_4287,N_3993,N_3642);
or U4288 (N_4288,N_3875,N_3941);
nor U4289 (N_4289,N_3537,N_3560);
nor U4290 (N_4290,N_3934,N_3740);
nand U4291 (N_4291,N_3651,N_3558);
xor U4292 (N_4292,N_3740,N_3949);
nor U4293 (N_4293,N_3896,N_3518);
and U4294 (N_4294,N_3921,N_3748);
and U4295 (N_4295,N_3523,N_3953);
and U4296 (N_4296,N_3553,N_3861);
or U4297 (N_4297,N_3941,N_3567);
xnor U4298 (N_4298,N_3559,N_3949);
nand U4299 (N_4299,N_3811,N_3873);
xnor U4300 (N_4300,N_3788,N_3742);
and U4301 (N_4301,N_3597,N_3715);
or U4302 (N_4302,N_3896,N_3740);
and U4303 (N_4303,N_3828,N_3944);
or U4304 (N_4304,N_3923,N_3525);
nand U4305 (N_4305,N_3560,N_3825);
or U4306 (N_4306,N_3701,N_3615);
xnor U4307 (N_4307,N_3764,N_3677);
xnor U4308 (N_4308,N_3777,N_3563);
nor U4309 (N_4309,N_3635,N_3758);
nand U4310 (N_4310,N_3760,N_3786);
xor U4311 (N_4311,N_3950,N_3984);
and U4312 (N_4312,N_3916,N_3705);
and U4313 (N_4313,N_3952,N_3601);
nand U4314 (N_4314,N_3735,N_3953);
and U4315 (N_4315,N_3690,N_3514);
and U4316 (N_4316,N_3889,N_3877);
nor U4317 (N_4317,N_3646,N_3861);
xor U4318 (N_4318,N_3850,N_3539);
nor U4319 (N_4319,N_3897,N_3713);
nor U4320 (N_4320,N_3920,N_3985);
and U4321 (N_4321,N_3577,N_3775);
nand U4322 (N_4322,N_3950,N_3723);
xnor U4323 (N_4323,N_3667,N_3852);
and U4324 (N_4324,N_3962,N_3852);
xnor U4325 (N_4325,N_3837,N_3986);
xor U4326 (N_4326,N_3598,N_3986);
nand U4327 (N_4327,N_3645,N_3769);
nor U4328 (N_4328,N_3548,N_3684);
and U4329 (N_4329,N_3786,N_3719);
nor U4330 (N_4330,N_3914,N_3641);
and U4331 (N_4331,N_3578,N_3657);
or U4332 (N_4332,N_3599,N_3523);
or U4333 (N_4333,N_3922,N_3763);
nand U4334 (N_4334,N_3863,N_3999);
nand U4335 (N_4335,N_3866,N_3561);
xnor U4336 (N_4336,N_3619,N_3617);
nand U4337 (N_4337,N_3688,N_3966);
xnor U4338 (N_4338,N_3503,N_3818);
nor U4339 (N_4339,N_3867,N_3637);
or U4340 (N_4340,N_3754,N_3594);
xor U4341 (N_4341,N_3705,N_3954);
nand U4342 (N_4342,N_3642,N_3971);
nor U4343 (N_4343,N_3525,N_3513);
or U4344 (N_4344,N_3628,N_3829);
nand U4345 (N_4345,N_3974,N_3816);
xnor U4346 (N_4346,N_3509,N_3741);
nor U4347 (N_4347,N_3865,N_3856);
nor U4348 (N_4348,N_3969,N_3607);
xor U4349 (N_4349,N_3715,N_3560);
or U4350 (N_4350,N_3827,N_3761);
and U4351 (N_4351,N_3666,N_3855);
or U4352 (N_4352,N_3981,N_3895);
nor U4353 (N_4353,N_3793,N_3691);
xnor U4354 (N_4354,N_3946,N_3643);
xor U4355 (N_4355,N_3691,N_3962);
and U4356 (N_4356,N_3836,N_3584);
xnor U4357 (N_4357,N_3786,N_3816);
xor U4358 (N_4358,N_3830,N_3990);
and U4359 (N_4359,N_3652,N_3738);
xor U4360 (N_4360,N_3806,N_3944);
nand U4361 (N_4361,N_3870,N_3941);
nand U4362 (N_4362,N_3982,N_3776);
xor U4363 (N_4363,N_3661,N_3932);
nor U4364 (N_4364,N_3746,N_3546);
and U4365 (N_4365,N_3690,N_3887);
xor U4366 (N_4366,N_3714,N_3665);
nor U4367 (N_4367,N_3787,N_3806);
and U4368 (N_4368,N_3749,N_3923);
or U4369 (N_4369,N_3536,N_3520);
nand U4370 (N_4370,N_3779,N_3788);
nor U4371 (N_4371,N_3941,N_3879);
and U4372 (N_4372,N_3638,N_3996);
or U4373 (N_4373,N_3903,N_3561);
or U4374 (N_4374,N_3679,N_3603);
nor U4375 (N_4375,N_3992,N_3851);
nand U4376 (N_4376,N_3524,N_3612);
nand U4377 (N_4377,N_3962,N_3615);
nand U4378 (N_4378,N_3941,N_3715);
xor U4379 (N_4379,N_3973,N_3987);
nor U4380 (N_4380,N_3978,N_3744);
xnor U4381 (N_4381,N_3992,N_3601);
xor U4382 (N_4382,N_3595,N_3813);
and U4383 (N_4383,N_3928,N_3878);
or U4384 (N_4384,N_3862,N_3740);
nor U4385 (N_4385,N_3946,N_3719);
nand U4386 (N_4386,N_3655,N_3775);
and U4387 (N_4387,N_3919,N_3940);
and U4388 (N_4388,N_3615,N_3534);
and U4389 (N_4389,N_3583,N_3769);
nand U4390 (N_4390,N_3991,N_3838);
or U4391 (N_4391,N_3795,N_3593);
and U4392 (N_4392,N_3748,N_3657);
xnor U4393 (N_4393,N_3614,N_3909);
and U4394 (N_4394,N_3507,N_3987);
xor U4395 (N_4395,N_3691,N_3674);
nor U4396 (N_4396,N_3574,N_3682);
xnor U4397 (N_4397,N_3559,N_3626);
nor U4398 (N_4398,N_3724,N_3676);
nand U4399 (N_4399,N_3616,N_3972);
and U4400 (N_4400,N_3665,N_3721);
xor U4401 (N_4401,N_3931,N_3505);
nor U4402 (N_4402,N_3773,N_3647);
or U4403 (N_4403,N_3660,N_3537);
nor U4404 (N_4404,N_3574,N_3724);
or U4405 (N_4405,N_3867,N_3505);
and U4406 (N_4406,N_3826,N_3711);
nand U4407 (N_4407,N_3996,N_3947);
and U4408 (N_4408,N_3857,N_3720);
xnor U4409 (N_4409,N_3679,N_3872);
and U4410 (N_4410,N_3819,N_3640);
nor U4411 (N_4411,N_3906,N_3801);
nor U4412 (N_4412,N_3707,N_3584);
nor U4413 (N_4413,N_3849,N_3720);
or U4414 (N_4414,N_3903,N_3862);
or U4415 (N_4415,N_3985,N_3974);
and U4416 (N_4416,N_3759,N_3677);
and U4417 (N_4417,N_3745,N_3592);
xnor U4418 (N_4418,N_3877,N_3586);
nor U4419 (N_4419,N_3621,N_3706);
nand U4420 (N_4420,N_3599,N_3851);
xor U4421 (N_4421,N_3573,N_3773);
xor U4422 (N_4422,N_3602,N_3799);
and U4423 (N_4423,N_3948,N_3631);
nand U4424 (N_4424,N_3795,N_3968);
or U4425 (N_4425,N_3920,N_3581);
nor U4426 (N_4426,N_3515,N_3671);
nand U4427 (N_4427,N_3801,N_3633);
nand U4428 (N_4428,N_3802,N_3513);
nor U4429 (N_4429,N_3698,N_3924);
nand U4430 (N_4430,N_3945,N_3728);
or U4431 (N_4431,N_3955,N_3576);
and U4432 (N_4432,N_3808,N_3580);
xnor U4433 (N_4433,N_3595,N_3625);
nor U4434 (N_4434,N_3519,N_3657);
nand U4435 (N_4435,N_3898,N_3684);
nand U4436 (N_4436,N_3957,N_3527);
xnor U4437 (N_4437,N_3650,N_3721);
and U4438 (N_4438,N_3614,N_3815);
and U4439 (N_4439,N_3502,N_3681);
nand U4440 (N_4440,N_3565,N_3641);
and U4441 (N_4441,N_3619,N_3518);
and U4442 (N_4442,N_3735,N_3555);
xor U4443 (N_4443,N_3822,N_3856);
nor U4444 (N_4444,N_3613,N_3945);
xor U4445 (N_4445,N_3972,N_3829);
nor U4446 (N_4446,N_3728,N_3529);
and U4447 (N_4447,N_3578,N_3541);
nand U4448 (N_4448,N_3793,N_3655);
nand U4449 (N_4449,N_3536,N_3945);
nor U4450 (N_4450,N_3863,N_3751);
and U4451 (N_4451,N_3769,N_3768);
and U4452 (N_4452,N_3888,N_3990);
xor U4453 (N_4453,N_3748,N_3824);
or U4454 (N_4454,N_3832,N_3720);
nor U4455 (N_4455,N_3823,N_3649);
and U4456 (N_4456,N_3794,N_3755);
xnor U4457 (N_4457,N_3794,N_3506);
and U4458 (N_4458,N_3564,N_3815);
nor U4459 (N_4459,N_3985,N_3934);
nand U4460 (N_4460,N_3500,N_3860);
nand U4461 (N_4461,N_3927,N_3945);
and U4462 (N_4462,N_3604,N_3613);
nand U4463 (N_4463,N_3852,N_3590);
nand U4464 (N_4464,N_3946,N_3886);
or U4465 (N_4465,N_3803,N_3790);
and U4466 (N_4466,N_3967,N_3541);
xor U4467 (N_4467,N_3568,N_3603);
and U4468 (N_4468,N_3568,N_3864);
or U4469 (N_4469,N_3771,N_3869);
nor U4470 (N_4470,N_3803,N_3501);
nor U4471 (N_4471,N_3911,N_3702);
nor U4472 (N_4472,N_3893,N_3657);
nand U4473 (N_4473,N_3573,N_3630);
nand U4474 (N_4474,N_3844,N_3943);
and U4475 (N_4475,N_3692,N_3576);
nor U4476 (N_4476,N_3605,N_3636);
and U4477 (N_4477,N_3638,N_3631);
nor U4478 (N_4478,N_3651,N_3748);
xnor U4479 (N_4479,N_3984,N_3578);
and U4480 (N_4480,N_3614,N_3979);
nor U4481 (N_4481,N_3578,N_3851);
and U4482 (N_4482,N_3987,N_3784);
and U4483 (N_4483,N_3779,N_3950);
xor U4484 (N_4484,N_3982,N_3718);
nand U4485 (N_4485,N_3852,N_3650);
and U4486 (N_4486,N_3778,N_3516);
nor U4487 (N_4487,N_3925,N_3878);
xnor U4488 (N_4488,N_3664,N_3633);
or U4489 (N_4489,N_3960,N_3602);
xnor U4490 (N_4490,N_3983,N_3621);
and U4491 (N_4491,N_3688,N_3946);
nand U4492 (N_4492,N_3816,N_3645);
xnor U4493 (N_4493,N_3883,N_3775);
and U4494 (N_4494,N_3995,N_3965);
or U4495 (N_4495,N_3930,N_3583);
nor U4496 (N_4496,N_3912,N_3927);
or U4497 (N_4497,N_3938,N_3727);
or U4498 (N_4498,N_3735,N_3996);
nor U4499 (N_4499,N_3614,N_3542);
nor U4500 (N_4500,N_4479,N_4093);
nor U4501 (N_4501,N_4300,N_4239);
xor U4502 (N_4502,N_4148,N_4301);
nor U4503 (N_4503,N_4433,N_4138);
or U4504 (N_4504,N_4183,N_4222);
nand U4505 (N_4505,N_4000,N_4079);
nor U4506 (N_4506,N_4360,N_4071);
nand U4507 (N_4507,N_4388,N_4243);
and U4508 (N_4508,N_4296,N_4132);
nand U4509 (N_4509,N_4114,N_4212);
nand U4510 (N_4510,N_4258,N_4369);
and U4511 (N_4511,N_4175,N_4249);
and U4512 (N_4512,N_4142,N_4282);
xnor U4513 (N_4513,N_4499,N_4234);
nand U4514 (N_4514,N_4029,N_4184);
nor U4515 (N_4515,N_4005,N_4167);
nor U4516 (N_4516,N_4270,N_4072);
and U4517 (N_4517,N_4205,N_4032);
and U4518 (N_4518,N_4008,N_4326);
xnor U4519 (N_4519,N_4204,N_4231);
and U4520 (N_4520,N_4421,N_4195);
or U4521 (N_4521,N_4238,N_4325);
nor U4522 (N_4522,N_4436,N_4059);
or U4523 (N_4523,N_4377,N_4244);
or U4524 (N_4524,N_4080,N_4268);
and U4525 (N_4525,N_4327,N_4474);
xor U4526 (N_4526,N_4434,N_4161);
or U4527 (N_4527,N_4216,N_4030);
or U4528 (N_4528,N_4026,N_4464);
xnor U4529 (N_4529,N_4150,N_4315);
and U4530 (N_4530,N_4082,N_4439);
nor U4531 (N_4531,N_4340,N_4387);
or U4532 (N_4532,N_4101,N_4115);
nor U4533 (N_4533,N_4170,N_4309);
xor U4534 (N_4534,N_4208,N_4061);
nand U4535 (N_4535,N_4437,N_4224);
and U4536 (N_4536,N_4261,N_4135);
xor U4537 (N_4537,N_4203,N_4346);
and U4538 (N_4538,N_4178,N_4223);
nand U4539 (N_4539,N_4073,N_4366);
xor U4540 (N_4540,N_4202,N_4154);
xnor U4541 (N_4541,N_4328,N_4062);
nand U4542 (N_4542,N_4305,N_4453);
and U4543 (N_4543,N_4156,N_4329);
or U4544 (N_4544,N_4050,N_4028);
xor U4545 (N_4545,N_4367,N_4016);
xor U4546 (N_4546,N_4339,N_4102);
xnor U4547 (N_4547,N_4476,N_4343);
nand U4548 (N_4548,N_4198,N_4381);
and U4549 (N_4549,N_4316,N_4482);
xor U4550 (N_4550,N_4283,N_4347);
nor U4551 (N_4551,N_4157,N_4291);
and U4552 (N_4552,N_4496,N_4133);
or U4553 (N_4553,N_4497,N_4067);
or U4554 (N_4554,N_4290,N_4025);
xnor U4555 (N_4555,N_4237,N_4475);
xor U4556 (N_4556,N_4352,N_4292);
or U4557 (N_4557,N_4463,N_4066);
nor U4558 (N_4558,N_4415,N_4351);
xnor U4559 (N_4559,N_4158,N_4117);
nor U4560 (N_4560,N_4179,N_4456);
xor U4561 (N_4561,N_4060,N_4333);
xnor U4562 (N_4562,N_4051,N_4215);
nor U4563 (N_4563,N_4130,N_4100);
nand U4564 (N_4564,N_4484,N_4152);
nand U4565 (N_4565,N_4252,N_4068);
xor U4566 (N_4566,N_4069,N_4012);
or U4567 (N_4567,N_4053,N_4171);
and U4568 (N_4568,N_4103,N_4047);
nand U4569 (N_4569,N_4221,N_4368);
and U4570 (N_4570,N_4407,N_4236);
nand U4571 (N_4571,N_4284,N_4281);
nor U4572 (N_4572,N_4039,N_4162);
and U4573 (N_4573,N_4087,N_4119);
nand U4574 (N_4574,N_4011,N_4332);
xnor U4575 (N_4575,N_4097,N_4277);
or U4576 (N_4576,N_4374,N_4031);
nor U4577 (N_4577,N_4054,N_4017);
or U4578 (N_4578,N_4324,N_4286);
and U4579 (N_4579,N_4376,N_4398);
or U4580 (N_4580,N_4293,N_4489);
and U4581 (N_4581,N_4124,N_4276);
and U4582 (N_4582,N_4354,N_4402);
and U4583 (N_4583,N_4401,N_4413);
nor U4584 (N_4584,N_4058,N_4105);
xnor U4585 (N_4585,N_4396,N_4323);
nor U4586 (N_4586,N_4335,N_4043);
nand U4587 (N_4587,N_4416,N_4266);
nor U4588 (N_4588,N_4227,N_4120);
and U4589 (N_4589,N_4055,N_4126);
xor U4590 (N_4590,N_4228,N_4384);
or U4591 (N_4591,N_4123,N_4090);
nand U4592 (N_4592,N_4450,N_4400);
nor U4593 (N_4593,N_4477,N_4498);
nand U4594 (N_4594,N_4487,N_4107);
nand U4595 (N_4595,N_4108,N_4033);
xor U4596 (N_4596,N_4085,N_4359);
xnor U4597 (N_4597,N_4454,N_4235);
or U4598 (N_4598,N_4313,N_4007);
or U4599 (N_4599,N_4230,N_4040);
xor U4600 (N_4600,N_4151,N_4446);
nor U4601 (N_4601,N_4317,N_4201);
or U4602 (N_4602,N_4096,N_4302);
nor U4603 (N_4603,N_4404,N_4395);
nor U4604 (N_4604,N_4455,N_4425);
and U4605 (N_4605,N_4191,N_4038);
xor U4606 (N_4606,N_4278,N_4188);
or U4607 (N_4607,N_4287,N_4448);
xor U4608 (N_4608,N_4465,N_4263);
nand U4609 (N_4609,N_4155,N_4297);
nor U4610 (N_4610,N_4190,N_4020);
xor U4611 (N_4611,N_4274,N_4273);
xnor U4612 (N_4612,N_4288,N_4037);
nor U4613 (N_4613,N_4417,N_4480);
and U4614 (N_4614,N_4137,N_4163);
nor U4615 (N_4615,N_4219,N_4397);
and U4616 (N_4616,N_4458,N_4122);
and U4617 (N_4617,N_4094,N_4147);
nand U4618 (N_4618,N_4310,N_4298);
nor U4619 (N_4619,N_4414,N_4084);
xnor U4620 (N_4620,N_4176,N_4412);
nor U4621 (N_4621,N_4070,N_4265);
nor U4622 (N_4622,N_4035,N_4468);
and U4623 (N_4623,N_4389,N_4267);
xor U4624 (N_4624,N_4023,N_4419);
nand U4625 (N_4625,N_4182,N_4226);
or U4626 (N_4626,N_4314,N_4077);
nand U4627 (N_4627,N_4430,N_4247);
or U4628 (N_4628,N_4334,N_4121);
xor U4629 (N_4629,N_4420,N_4350);
xnor U4630 (N_4630,N_4086,N_4036);
or U4631 (N_4631,N_4022,N_4358);
or U4632 (N_4632,N_4153,N_4214);
or U4633 (N_4633,N_4472,N_4015);
xnor U4634 (N_4634,N_4185,N_4382);
xnor U4635 (N_4635,N_4257,N_4125);
and U4636 (N_4636,N_4337,N_4386);
and U4637 (N_4637,N_4116,N_4380);
nand U4638 (N_4638,N_4321,N_4356);
or U4639 (N_4639,N_4089,N_4394);
nor U4640 (N_4640,N_4034,N_4391);
nand U4641 (N_4641,N_4242,N_4483);
or U4642 (N_4642,N_4285,N_4295);
nand U4643 (N_4643,N_4001,N_4041);
nand U4644 (N_4644,N_4181,N_4074);
xnor U4645 (N_4645,N_4319,N_4345);
xnor U4646 (N_4646,N_4423,N_4139);
nor U4647 (N_4647,N_4373,N_4232);
nand U4648 (N_4648,N_4443,N_4169);
and U4649 (N_4649,N_4390,N_4442);
nand U4650 (N_4650,N_4262,N_4409);
and U4651 (N_4651,N_4372,N_4209);
or U4652 (N_4652,N_4312,N_4210);
or U4653 (N_4653,N_4164,N_4355);
xor U4654 (N_4654,N_4392,N_4166);
nand U4655 (N_4655,N_4406,N_4225);
nor U4656 (N_4656,N_4375,N_4146);
nand U4657 (N_4657,N_4251,N_4399);
or U4658 (N_4658,N_4174,N_4027);
and U4659 (N_4659,N_4246,N_4299);
nand U4660 (N_4660,N_4320,N_4189);
xnor U4661 (N_4661,N_4106,N_4330);
xnor U4662 (N_4662,N_4075,N_4045);
nand U4663 (N_4663,N_4308,N_4271);
nand U4664 (N_4664,N_4014,N_4118);
nor U4665 (N_4665,N_4469,N_4311);
nand U4666 (N_4666,N_4131,N_4338);
or U4667 (N_4667,N_4431,N_4466);
or U4668 (N_4668,N_4003,N_4403);
nand U4669 (N_4669,N_4385,N_4322);
and U4670 (N_4670,N_4078,N_4471);
nor U4671 (N_4671,N_4379,N_4091);
xor U4672 (N_4672,N_4452,N_4095);
nand U4673 (N_4673,N_4460,N_4294);
and U4674 (N_4674,N_4445,N_4485);
nor U4675 (N_4675,N_4424,N_4365);
nor U4676 (N_4676,N_4196,N_4063);
xor U4677 (N_4677,N_4165,N_4341);
nor U4678 (N_4678,N_4478,N_4303);
and U4679 (N_4679,N_4428,N_4411);
xnor U4680 (N_4680,N_4160,N_4378);
nand U4681 (N_4681,N_4177,N_4206);
and U4682 (N_4682,N_4289,N_4110);
and U4683 (N_4683,N_4192,N_4393);
and U4684 (N_4684,N_4427,N_4010);
xor U4685 (N_4685,N_4044,N_4111);
and U4686 (N_4686,N_4269,N_4444);
xnor U4687 (N_4687,N_4451,N_4492);
or U4688 (N_4688,N_4021,N_4254);
xnor U4689 (N_4689,N_4098,N_4002);
or U4690 (N_4690,N_4218,N_4199);
and U4691 (N_4691,N_4470,N_4304);
xnor U4692 (N_4692,N_4006,N_4193);
nand U4693 (N_4693,N_4140,N_4211);
nand U4694 (N_4694,N_4495,N_4088);
or U4695 (N_4695,N_4241,N_4429);
and U4696 (N_4696,N_4172,N_4024);
xnor U4697 (N_4697,N_4256,N_4462);
and U4698 (N_4698,N_4180,N_4159);
nand U4699 (N_4699,N_4109,N_4076);
and U4700 (N_4700,N_4449,N_4134);
xnor U4701 (N_4701,N_4018,N_4481);
nand U4702 (N_4702,N_4461,N_4217);
and U4703 (N_4703,N_4342,N_4057);
and U4704 (N_4704,N_4457,N_4013);
nand U4705 (N_4705,N_4426,N_4113);
nor U4706 (N_4706,N_4432,N_4440);
nor U4707 (N_4707,N_4128,N_4279);
nand U4708 (N_4708,N_4491,N_4353);
nand U4709 (N_4709,N_4318,N_4083);
and U4710 (N_4710,N_4197,N_4348);
or U4711 (N_4711,N_4331,N_4143);
nor U4712 (N_4712,N_4435,N_4187);
xnor U4713 (N_4713,N_4410,N_4418);
nand U4714 (N_4714,N_4240,N_4364);
or U4715 (N_4715,N_4046,N_4494);
nor U4716 (N_4716,N_4336,N_4144);
xor U4717 (N_4717,N_4447,N_4052);
xor U4718 (N_4718,N_4229,N_4438);
nor U4719 (N_4719,N_4306,N_4127);
or U4720 (N_4720,N_4145,N_4129);
nand U4721 (N_4721,N_4259,N_4042);
or U4722 (N_4722,N_4253,N_4371);
nand U4723 (N_4723,N_4272,N_4207);
and U4724 (N_4724,N_4248,N_4141);
nor U4725 (N_4725,N_4357,N_4275);
or U4726 (N_4726,N_4405,N_4493);
and U4727 (N_4727,N_4280,N_4233);
nand U4728 (N_4728,N_4149,N_4173);
and U4729 (N_4729,N_4473,N_4459);
xor U4730 (N_4730,N_4361,N_4255);
or U4731 (N_4731,N_4065,N_4344);
or U4732 (N_4732,N_4081,N_4056);
or U4733 (N_4733,N_4049,N_4383);
and U4734 (N_4734,N_4349,N_4048);
nor U4735 (N_4735,N_4245,N_4186);
nand U4736 (N_4736,N_4307,N_4362);
or U4737 (N_4737,N_4260,N_4136);
and U4738 (N_4738,N_4194,N_4408);
or U4739 (N_4739,N_4112,N_4064);
or U4740 (N_4740,N_4168,N_4099);
xor U4741 (N_4741,N_4009,N_4104);
xnor U4742 (N_4742,N_4004,N_4422);
xnor U4743 (N_4743,N_4363,N_4200);
and U4744 (N_4744,N_4250,N_4092);
nand U4745 (N_4745,N_4213,N_4488);
nor U4746 (N_4746,N_4019,N_4490);
nand U4747 (N_4747,N_4486,N_4264);
xnor U4748 (N_4748,N_4467,N_4370);
nor U4749 (N_4749,N_4441,N_4220);
nor U4750 (N_4750,N_4370,N_4173);
or U4751 (N_4751,N_4469,N_4438);
nor U4752 (N_4752,N_4200,N_4321);
xnor U4753 (N_4753,N_4317,N_4266);
xor U4754 (N_4754,N_4051,N_4413);
and U4755 (N_4755,N_4088,N_4302);
and U4756 (N_4756,N_4012,N_4279);
and U4757 (N_4757,N_4454,N_4002);
nor U4758 (N_4758,N_4459,N_4147);
nor U4759 (N_4759,N_4393,N_4223);
and U4760 (N_4760,N_4439,N_4044);
and U4761 (N_4761,N_4224,N_4412);
nand U4762 (N_4762,N_4235,N_4050);
and U4763 (N_4763,N_4172,N_4035);
nand U4764 (N_4764,N_4072,N_4200);
nand U4765 (N_4765,N_4143,N_4163);
nand U4766 (N_4766,N_4432,N_4448);
xnor U4767 (N_4767,N_4010,N_4496);
and U4768 (N_4768,N_4004,N_4076);
or U4769 (N_4769,N_4311,N_4232);
or U4770 (N_4770,N_4219,N_4034);
nor U4771 (N_4771,N_4399,N_4216);
nor U4772 (N_4772,N_4490,N_4031);
nand U4773 (N_4773,N_4211,N_4417);
nor U4774 (N_4774,N_4227,N_4456);
and U4775 (N_4775,N_4334,N_4226);
and U4776 (N_4776,N_4422,N_4362);
nor U4777 (N_4777,N_4236,N_4349);
xor U4778 (N_4778,N_4163,N_4016);
and U4779 (N_4779,N_4327,N_4426);
nor U4780 (N_4780,N_4434,N_4213);
and U4781 (N_4781,N_4495,N_4320);
and U4782 (N_4782,N_4429,N_4075);
and U4783 (N_4783,N_4332,N_4115);
or U4784 (N_4784,N_4214,N_4165);
nand U4785 (N_4785,N_4382,N_4124);
xnor U4786 (N_4786,N_4132,N_4423);
and U4787 (N_4787,N_4467,N_4340);
xnor U4788 (N_4788,N_4213,N_4266);
nor U4789 (N_4789,N_4293,N_4107);
xnor U4790 (N_4790,N_4041,N_4386);
nor U4791 (N_4791,N_4117,N_4438);
and U4792 (N_4792,N_4294,N_4018);
nor U4793 (N_4793,N_4233,N_4153);
nand U4794 (N_4794,N_4441,N_4474);
nor U4795 (N_4795,N_4341,N_4216);
or U4796 (N_4796,N_4123,N_4033);
xor U4797 (N_4797,N_4376,N_4395);
and U4798 (N_4798,N_4094,N_4175);
or U4799 (N_4799,N_4202,N_4053);
xnor U4800 (N_4800,N_4461,N_4121);
nor U4801 (N_4801,N_4234,N_4158);
and U4802 (N_4802,N_4036,N_4399);
nand U4803 (N_4803,N_4121,N_4244);
nor U4804 (N_4804,N_4311,N_4259);
nand U4805 (N_4805,N_4327,N_4494);
xnor U4806 (N_4806,N_4196,N_4047);
xor U4807 (N_4807,N_4033,N_4267);
xor U4808 (N_4808,N_4020,N_4201);
nor U4809 (N_4809,N_4086,N_4437);
xnor U4810 (N_4810,N_4466,N_4273);
or U4811 (N_4811,N_4316,N_4326);
and U4812 (N_4812,N_4097,N_4060);
or U4813 (N_4813,N_4422,N_4441);
xor U4814 (N_4814,N_4455,N_4048);
or U4815 (N_4815,N_4088,N_4331);
xnor U4816 (N_4816,N_4254,N_4132);
and U4817 (N_4817,N_4311,N_4173);
nand U4818 (N_4818,N_4355,N_4167);
nor U4819 (N_4819,N_4101,N_4307);
or U4820 (N_4820,N_4369,N_4211);
nor U4821 (N_4821,N_4499,N_4323);
or U4822 (N_4822,N_4316,N_4378);
xor U4823 (N_4823,N_4141,N_4013);
nor U4824 (N_4824,N_4340,N_4457);
and U4825 (N_4825,N_4106,N_4005);
nor U4826 (N_4826,N_4332,N_4220);
or U4827 (N_4827,N_4426,N_4466);
and U4828 (N_4828,N_4242,N_4377);
xnor U4829 (N_4829,N_4058,N_4228);
xnor U4830 (N_4830,N_4087,N_4082);
xnor U4831 (N_4831,N_4432,N_4399);
nor U4832 (N_4832,N_4286,N_4174);
nand U4833 (N_4833,N_4495,N_4254);
or U4834 (N_4834,N_4144,N_4147);
nor U4835 (N_4835,N_4284,N_4373);
nand U4836 (N_4836,N_4497,N_4170);
and U4837 (N_4837,N_4018,N_4420);
nor U4838 (N_4838,N_4087,N_4330);
nor U4839 (N_4839,N_4223,N_4208);
or U4840 (N_4840,N_4318,N_4452);
nor U4841 (N_4841,N_4062,N_4048);
or U4842 (N_4842,N_4378,N_4219);
or U4843 (N_4843,N_4018,N_4328);
nor U4844 (N_4844,N_4225,N_4299);
xor U4845 (N_4845,N_4019,N_4452);
nand U4846 (N_4846,N_4069,N_4362);
xor U4847 (N_4847,N_4366,N_4104);
nand U4848 (N_4848,N_4151,N_4002);
nand U4849 (N_4849,N_4266,N_4396);
and U4850 (N_4850,N_4217,N_4036);
xor U4851 (N_4851,N_4106,N_4455);
xor U4852 (N_4852,N_4349,N_4238);
or U4853 (N_4853,N_4359,N_4120);
nand U4854 (N_4854,N_4230,N_4399);
nand U4855 (N_4855,N_4070,N_4364);
and U4856 (N_4856,N_4218,N_4054);
and U4857 (N_4857,N_4031,N_4317);
and U4858 (N_4858,N_4457,N_4085);
xnor U4859 (N_4859,N_4205,N_4315);
nor U4860 (N_4860,N_4300,N_4426);
nor U4861 (N_4861,N_4310,N_4225);
nand U4862 (N_4862,N_4257,N_4235);
xnor U4863 (N_4863,N_4495,N_4065);
or U4864 (N_4864,N_4214,N_4060);
xor U4865 (N_4865,N_4429,N_4407);
and U4866 (N_4866,N_4140,N_4463);
nand U4867 (N_4867,N_4064,N_4157);
and U4868 (N_4868,N_4315,N_4248);
xnor U4869 (N_4869,N_4080,N_4241);
xnor U4870 (N_4870,N_4337,N_4293);
nand U4871 (N_4871,N_4483,N_4118);
nand U4872 (N_4872,N_4017,N_4312);
and U4873 (N_4873,N_4444,N_4021);
nand U4874 (N_4874,N_4156,N_4488);
nor U4875 (N_4875,N_4427,N_4342);
nand U4876 (N_4876,N_4281,N_4360);
nor U4877 (N_4877,N_4094,N_4169);
or U4878 (N_4878,N_4450,N_4380);
xnor U4879 (N_4879,N_4449,N_4413);
or U4880 (N_4880,N_4117,N_4394);
and U4881 (N_4881,N_4461,N_4466);
and U4882 (N_4882,N_4402,N_4249);
nand U4883 (N_4883,N_4490,N_4388);
and U4884 (N_4884,N_4496,N_4443);
xor U4885 (N_4885,N_4366,N_4364);
nor U4886 (N_4886,N_4196,N_4176);
xor U4887 (N_4887,N_4026,N_4253);
nor U4888 (N_4888,N_4281,N_4010);
nor U4889 (N_4889,N_4354,N_4218);
and U4890 (N_4890,N_4264,N_4291);
xnor U4891 (N_4891,N_4360,N_4278);
xor U4892 (N_4892,N_4289,N_4467);
or U4893 (N_4893,N_4083,N_4056);
xnor U4894 (N_4894,N_4135,N_4361);
and U4895 (N_4895,N_4247,N_4054);
xnor U4896 (N_4896,N_4372,N_4422);
nor U4897 (N_4897,N_4040,N_4003);
nand U4898 (N_4898,N_4095,N_4257);
nor U4899 (N_4899,N_4446,N_4333);
nand U4900 (N_4900,N_4409,N_4246);
xnor U4901 (N_4901,N_4234,N_4315);
and U4902 (N_4902,N_4157,N_4348);
nor U4903 (N_4903,N_4289,N_4497);
xnor U4904 (N_4904,N_4178,N_4136);
or U4905 (N_4905,N_4311,N_4175);
xnor U4906 (N_4906,N_4471,N_4485);
and U4907 (N_4907,N_4141,N_4397);
and U4908 (N_4908,N_4262,N_4269);
or U4909 (N_4909,N_4058,N_4193);
nand U4910 (N_4910,N_4481,N_4317);
and U4911 (N_4911,N_4285,N_4173);
or U4912 (N_4912,N_4097,N_4192);
or U4913 (N_4913,N_4455,N_4255);
xnor U4914 (N_4914,N_4104,N_4043);
xnor U4915 (N_4915,N_4144,N_4033);
or U4916 (N_4916,N_4299,N_4043);
nand U4917 (N_4917,N_4262,N_4060);
and U4918 (N_4918,N_4069,N_4074);
xnor U4919 (N_4919,N_4371,N_4230);
nand U4920 (N_4920,N_4062,N_4488);
xnor U4921 (N_4921,N_4386,N_4488);
or U4922 (N_4922,N_4132,N_4273);
and U4923 (N_4923,N_4396,N_4081);
and U4924 (N_4924,N_4039,N_4020);
or U4925 (N_4925,N_4176,N_4229);
nor U4926 (N_4926,N_4443,N_4450);
and U4927 (N_4927,N_4290,N_4037);
nand U4928 (N_4928,N_4380,N_4157);
nand U4929 (N_4929,N_4153,N_4032);
nand U4930 (N_4930,N_4483,N_4163);
xnor U4931 (N_4931,N_4271,N_4080);
and U4932 (N_4932,N_4282,N_4144);
nand U4933 (N_4933,N_4235,N_4175);
nand U4934 (N_4934,N_4315,N_4161);
and U4935 (N_4935,N_4163,N_4338);
xor U4936 (N_4936,N_4408,N_4490);
and U4937 (N_4937,N_4397,N_4401);
or U4938 (N_4938,N_4375,N_4198);
nor U4939 (N_4939,N_4334,N_4376);
and U4940 (N_4940,N_4419,N_4457);
xnor U4941 (N_4941,N_4216,N_4035);
nand U4942 (N_4942,N_4424,N_4116);
nor U4943 (N_4943,N_4469,N_4282);
nor U4944 (N_4944,N_4378,N_4369);
nor U4945 (N_4945,N_4417,N_4039);
nor U4946 (N_4946,N_4288,N_4293);
and U4947 (N_4947,N_4094,N_4301);
nor U4948 (N_4948,N_4354,N_4498);
or U4949 (N_4949,N_4358,N_4436);
and U4950 (N_4950,N_4125,N_4208);
nor U4951 (N_4951,N_4258,N_4295);
or U4952 (N_4952,N_4420,N_4416);
and U4953 (N_4953,N_4303,N_4096);
or U4954 (N_4954,N_4220,N_4324);
xor U4955 (N_4955,N_4152,N_4001);
xor U4956 (N_4956,N_4375,N_4004);
or U4957 (N_4957,N_4025,N_4037);
and U4958 (N_4958,N_4384,N_4262);
or U4959 (N_4959,N_4200,N_4214);
xor U4960 (N_4960,N_4215,N_4364);
xnor U4961 (N_4961,N_4260,N_4492);
xnor U4962 (N_4962,N_4058,N_4439);
nor U4963 (N_4963,N_4139,N_4084);
and U4964 (N_4964,N_4199,N_4373);
nor U4965 (N_4965,N_4316,N_4180);
nor U4966 (N_4966,N_4435,N_4036);
xnor U4967 (N_4967,N_4336,N_4271);
nor U4968 (N_4968,N_4404,N_4266);
nor U4969 (N_4969,N_4407,N_4199);
xnor U4970 (N_4970,N_4195,N_4240);
or U4971 (N_4971,N_4170,N_4300);
and U4972 (N_4972,N_4336,N_4185);
nand U4973 (N_4973,N_4159,N_4347);
xnor U4974 (N_4974,N_4072,N_4001);
and U4975 (N_4975,N_4231,N_4236);
xnor U4976 (N_4976,N_4216,N_4490);
nand U4977 (N_4977,N_4440,N_4138);
nand U4978 (N_4978,N_4283,N_4174);
or U4979 (N_4979,N_4279,N_4323);
xor U4980 (N_4980,N_4423,N_4299);
nand U4981 (N_4981,N_4486,N_4382);
nor U4982 (N_4982,N_4229,N_4347);
nor U4983 (N_4983,N_4244,N_4469);
nor U4984 (N_4984,N_4031,N_4103);
nor U4985 (N_4985,N_4266,N_4466);
nor U4986 (N_4986,N_4315,N_4472);
nor U4987 (N_4987,N_4399,N_4473);
xnor U4988 (N_4988,N_4038,N_4018);
nand U4989 (N_4989,N_4370,N_4289);
nor U4990 (N_4990,N_4385,N_4119);
nor U4991 (N_4991,N_4080,N_4351);
and U4992 (N_4992,N_4139,N_4325);
or U4993 (N_4993,N_4215,N_4449);
and U4994 (N_4994,N_4302,N_4396);
or U4995 (N_4995,N_4077,N_4206);
nand U4996 (N_4996,N_4040,N_4305);
nand U4997 (N_4997,N_4244,N_4158);
or U4998 (N_4998,N_4474,N_4159);
nor U4999 (N_4999,N_4162,N_4079);
xnor U5000 (N_5000,N_4784,N_4979);
nand U5001 (N_5001,N_4949,N_4975);
and U5002 (N_5002,N_4615,N_4556);
or U5003 (N_5003,N_4922,N_4779);
and U5004 (N_5004,N_4725,N_4758);
nand U5005 (N_5005,N_4567,N_4551);
or U5006 (N_5006,N_4711,N_4673);
xor U5007 (N_5007,N_4781,N_4601);
nand U5008 (N_5008,N_4737,N_4749);
nor U5009 (N_5009,N_4943,N_4706);
nand U5010 (N_5010,N_4665,N_4692);
or U5011 (N_5011,N_4807,N_4533);
or U5012 (N_5012,N_4868,N_4521);
or U5013 (N_5013,N_4919,N_4677);
nor U5014 (N_5014,N_4759,N_4780);
nor U5015 (N_5015,N_4789,N_4592);
and U5016 (N_5016,N_4757,N_4653);
nand U5017 (N_5017,N_4877,N_4596);
and U5018 (N_5018,N_4838,N_4873);
xor U5019 (N_5019,N_4754,N_4654);
xor U5020 (N_5020,N_4538,N_4973);
xor U5021 (N_5021,N_4762,N_4717);
nand U5022 (N_5022,N_4884,N_4516);
nor U5023 (N_5023,N_4980,N_4597);
nand U5024 (N_5024,N_4774,N_4995);
xnor U5025 (N_5025,N_4619,N_4939);
nand U5026 (N_5026,N_4520,N_4502);
xor U5027 (N_5027,N_4608,N_4766);
or U5028 (N_5028,N_4964,N_4863);
xnor U5029 (N_5029,N_4823,N_4934);
xnor U5030 (N_5030,N_4933,N_4657);
and U5031 (N_5031,N_4954,N_4517);
or U5032 (N_5032,N_4595,N_4890);
and U5033 (N_5033,N_4746,N_4817);
nor U5034 (N_5034,N_4843,N_4658);
or U5035 (N_5035,N_4745,N_4947);
nor U5036 (N_5036,N_4839,N_4829);
nor U5037 (N_5037,N_4752,N_4786);
or U5038 (N_5038,N_4887,N_4756);
and U5039 (N_5039,N_4664,N_4881);
xnor U5040 (N_5040,N_4531,N_4590);
nor U5041 (N_5041,N_4514,N_4747);
or U5042 (N_5042,N_4697,N_4679);
and U5043 (N_5043,N_4908,N_4764);
nor U5044 (N_5044,N_4668,N_4699);
or U5045 (N_5045,N_4965,N_4661);
and U5046 (N_5046,N_4687,N_4804);
nor U5047 (N_5047,N_4988,N_4994);
nor U5048 (N_5048,N_4923,N_4989);
nand U5049 (N_5049,N_4946,N_4820);
nand U5050 (N_5050,N_4510,N_4961);
and U5051 (N_5051,N_4802,N_4631);
nor U5052 (N_5052,N_4584,N_4501);
xor U5053 (N_5053,N_4869,N_4778);
and U5054 (N_5054,N_4945,N_4573);
xor U5055 (N_5055,N_4856,N_4633);
and U5056 (N_5056,N_4571,N_4763);
or U5057 (N_5057,N_4893,N_4587);
nand U5058 (N_5058,N_4998,N_4637);
and U5059 (N_5059,N_4635,N_4907);
nand U5060 (N_5060,N_4912,N_4525);
nor U5061 (N_5061,N_4710,N_4899);
or U5062 (N_5062,N_4667,N_4638);
and U5063 (N_5063,N_4996,N_4850);
nor U5064 (N_5064,N_4546,N_4929);
nor U5065 (N_5065,N_4519,N_4643);
or U5066 (N_5066,N_4917,N_4876);
nor U5067 (N_5067,N_4663,N_4523);
nand U5068 (N_5068,N_4532,N_4705);
xor U5069 (N_5069,N_4897,N_4901);
or U5070 (N_5070,N_4834,N_4669);
and U5071 (N_5071,N_4632,N_4909);
and U5072 (N_5072,N_4888,N_4844);
nand U5073 (N_5073,N_4809,N_4575);
and U5074 (N_5074,N_4832,N_4801);
or U5075 (N_5075,N_4741,N_4526);
nand U5076 (N_5076,N_4736,N_4915);
xnor U5077 (N_5077,N_4629,N_4794);
or U5078 (N_5078,N_4625,N_4616);
nand U5079 (N_5079,N_4788,N_4713);
nand U5080 (N_5080,N_4729,N_4626);
xnor U5081 (N_5081,N_4981,N_4606);
and U5082 (N_5082,N_4591,N_4544);
xnor U5083 (N_5083,N_4530,N_4503);
and U5084 (N_5084,N_4845,N_4603);
and U5085 (N_5085,N_4542,N_4722);
or U5086 (N_5086,N_4560,N_4925);
or U5087 (N_5087,N_4636,N_4730);
xor U5088 (N_5088,N_4536,N_4750);
xnor U5089 (N_5089,N_4685,N_4874);
nand U5090 (N_5090,N_4641,N_4822);
or U5091 (N_5091,N_4936,N_4691);
or U5092 (N_5092,N_4914,N_4642);
and U5093 (N_5093,N_4892,N_4751);
xor U5094 (N_5094,N_4840,N_4900);
or U5095 (N_5095,N_4977,N_4680);
xnor U5096 (N_5096,N_4739,N_4805);
xnor U5097 (N_5097,N_4671,N_4703);
and U5098 (N_5098,N_4707,N_4851);
nor U5099 (N_5099,N_4921,N_4612);
xnor U5100 (N_5100,N_4728,N_4513);
and U5101 (N_5101,N_4708,N_4785);
or U5102 (N_5102,N_4617,N_4806);
xnor U5103 (N_5103,N_4557,N_4767);
or U5104 (N_5104,N_4861,N_4647);
nor U5105 (N_5105,N_4846,N_4581);
nor U5106 (N_5106,N_4618,N_4795);
nor U5107 (N_5107,N_4716,N_4527);
or U5108 (N_5108,N_4955,N_4579);
and U5109 (N_5109,N_4660,N_4704);
nor U5110 (N_5110,N_4753,N_4734);
and U5111 (N_5111,N_4537,N_4937);
xor U5112 (N_5112,N_4515,N_4920);
nor U5113 (N_5113,N_4534,N_4572);
nor U5114 (N_5114,N_4577,N_4570);
xor U5115 (N_5115,N_4622,N_4718);
or U5116 (N_5116,N_4999,N_4755);
nor U5117 (N_5117,N_4621,N_4623);
or U5118 (N_5118,N_4549,N_4672);
or U5119 (N_5119,N_4506,N_4640);
nand U5120 (N_5120,N_4924,N_4870);
nor U5121 (N_5121,N_4528,N_4659);
nand U5122 (N_5122,N_4772,N_4656);
xor U5123 (N_5123,N_4848,N_4547);
or U5124 (N_5124,N_4613,N_4504);
or U5125 (N_5125,N_4889,N_4564);
xnor U5126 (N_5126,N_4720,N_4586);
nor U5127 (N_5127,N_4776,N_4858);
xor U5128 (N_5128,N_4942,N_4787);
and U5129 (N_5129,N_4676,N_4651);
nand U5130 (N_5130,N_4568,N_4896);
nand U5131 (N_5131,N_4849,N_4550);
or U5132 (N_5132,N_4593,N_4683);
and U5133 (N_5133,N_4953,N_4627);
and U5134 (N_5134,N_4831,N_4648);
nand U5135 (N_5135,N_4866,N_4916);
nand U5136 (N_5136,N_4803,N_4727);
or U5137 (N_5137,N_4562,N_4652);
nor U5138 (N_5138,N_4948,N_4726);
xnor U5139 (N_5139,N_4970,N_4518);
nor U5140 (N_5140,N_4681,N_4983);
nand U5141 (N_5141,N_4715,N_4552);
and U5142 (N_5142,N_4771,N_4740);
nand U5143 (N_5143,N_4927,N_4796);
nor U5144 (N_5144,N_4854,N_4875);
and U5145 (N_5145,N_4940,N_4976);
and U5146 (N_5146,N_4952,N_4935);
nor U5147 (N_5147,N_4860,N_4855);
nor U5148 (N_5148,N_4529,N_4878);
and U5149 (N_5149,N_4793,N_4960);
xor U5150 (N_5150,N_4524,N_4662);
nor U5151 (N_5151,N_4565,N_4993);
nand U5152 (N_5152,N_4959,N_4545);
or U5153 (N_5153,N_4733,N_4997);
or U5154 (N_5154,N_4598,N_4963);
or U5155 (N_5155,N_4882,N_4775);
or U5156 (N_5156,N_4956,N_4992);
xnor U5157 (N_5157,N_4972,N_4968);
xnor U5158 (N_5158,N_4883,N_4694);
nor U5159 (N_5159,N_4903,N_4828);
or U5160 (N_5160,N_4974,N_4902);
and U5161 (N_5161,N_4987,N_4885);
xor U5162 (N_5162,N_4600,N_4712);
or U5163 (N_5163,N_4906,N_4773);
and U5164 (N_5164,N_4624,N_4815);
or U5165 (N_5165,N_4872,N_4769);
or U5166 (N_5166,N_4693,N_4821);
or U5167 (N_5167,N_4941,N_4599);
nor U5168 (N_5168,N_4792,N_4926);
and U5169 (N_5169,N_4743,N_4814);
xnor U5170 (N_5170,N_4958,N_4871);
or U5171 (N_5171,N_4790,N_4583);
or U5172 (N_5172,N_4835,N_4985);
xnor U5173 (N_5173,N_4696,N_4990);
nand U5174 (N_5174,N_4826,N_4594);
or U5175 (N_5175,N_4678,N_4830);
nand U5176 (N_5176,N_4701,N_4978);
nor U5177 (N_5177,N_4818,N_4798);
or U5178 (N_5178,N_4837,N_4825);
or U5179 (N_5179,N_4799,N_4512);
and U5180 (N_5180,N_4862,N_4604);
nor U5181 (N_5181,N_4645,N_4841);
or U5182 (N_5182,N_4724,N_4555);
nor U5183 (N_5183,N_4723,N_4675);
or U5184 (N_5184,N_4865,N_4554);
nand U5185 (N_5185,N_4760,N_4607);
nor U5186 (N_5186,N_4931,N_4966);
xnor U5187 (N_5187,N_4684,N_4852);
xnor U5188 (N_5188,N_4833,N_4700);
nor U5189 (N_5189,N_4742,N_4649);
nor U5190 (N_5190,N_4614,N_4650);
nand U5191 (N_5191,N_4836,N_4569);
or U5192 (N_5192,N_4732,N_4859);
or U5193 (N_5193,N_4628,N_4951);
xnor U5194 (N_5194,N_4864,N_4574);
and U5195 (N_5195,N_4508,N_4655);
nor U5196 (N_5196,N_4904,N_4895);
nand U5197 (N_5197,N_4811,N_4761);
nor U5198 (N_5198,N_4563,N_4950);
and U5199 (N_5199,N_4507,N_4509);
nor U5200 (N_5200,N_4605,N_4553);
and U5201 (N_5201,N_4689,N_4886);
xnor U5202 (N_5202,N_4777,N_4666);
nor U5203 (N_5203,N_4646,N_4842);
or U5204 (N_5204,N_4827,N_4630);
nand U5205 (N_5205,N_4932,N_4539);
nor U5206 (N_5206,N_4602,N_4611);
nand U5207 (N_5207,N_4561,N_4748);
nand U5208 (N_5208,N_4690,N_4971);
nand U5209 (N_5209,N_4644,N_4731);
and U5210 (N_5210,N_4957,N_4735);
nor U5211 (N_5211,N_4911,N_4721);
xor U5212 (N_5212,N_4918,N_4610);
xor U5213 (N_5213,N_4797,N_4738);
and U5214 (N_5214,N_4580,N_4558);
nor U5215 (N_5215,N_4910,N_4576);
or U5216 (N_5216,N_4824,N_4800);
and U5217 (N_5217,N_4810,N_4535);
nand U5218 (N_5218,N_4894,N_4744);
and U5219 (N_5219,N_4944,N_4791);
and U5220 (N_5220,N_4768,N_4813);
or U5221 (N_5221,N_4578,N_4765);
nor U5222 (N_5222,N_4898,N_4609);
nor U5223 (N_5223,N_4709,N_4857);
xor U5224 (N_5224,N_4688,N_4522);
xor U5225 (N_5225,N_4770,N_4543);
or U5226 (N_5226,N_4695,N_4670);
nor U5227 (N_5227,N_4853,N_4682);
xnor U5228 (N_5228,N_4620,N_4674);
nand U5229 (N_5229,N_4566,N_4816);
nor U5230 (N_5230,N_4812,N_4541);
or U5231 (N_5231,N_4982,N_4930);
or U5232 (N_5232,N_4559,N_4808);
nor U5233 (N_5233,N_4548,N_4938);
nor U5234 (N_5234,N_4500,N_4714);
and U5235 (N_5235,N_4891,N_4589);
xor U5236 (N_5236,N_4969,N_4686);
and U5237 (N_5237,N_4540,N_4867);
xor U5238 (N_5238,N_4991,N_4880);
and U5239 (N_5239,N_4582,N_4585);
nor U5240 (N_5240,N_4782,N_4962);
and U5241 (N_5241,N_4783,N_4588);
and U5242 (N_5242,N_4511,N_4719);
xnor U5243 (N_5243,N_4984,N_4847);
and U5244 (N_5244,N_4905,N_4928);
xnor U5245 (N_5245,N_4505,N_4698);
and U5246 (N_5246,N_4967,N_4879);
xnor U5247 (N_5247,N_4986,N_4634);
or U5248 (N_5248,N_4819,N_4702);
or U5249 (N_5249,N_4913,N_4639);
or U5250 (N_5250,N_4749,N_4992);
or U5251 (N_5251,N_4719,N_4849);
nor U5252 (N_5252,N_4786,N_4990);
and U5253 (N_5253,N_4594,N_4974);
nand U5254 (N_5254,N_4889,N_4981);
nor U5255 (N_5255,N_4683,N_4867);
nand U5256 (N_5256,N_4919,N_4921);
and U5257 (N_5257,N_4519,N_4772);
nor U5258 (N_5258,N_4802,N_4856);
nand U5259 (N_5259,N_4901,N_4641);
or U5260 (N_5260,N_4644,N_4988);
or U5261 (N_5261,N_4749,N_4819);
or U5262 (N_5262,N_4678,N_4875);
or U5263 (N_5263,N_4546,N_4631);
xnor U5264 (N_5264,N_4528,N_4565);
nand U5265 (N_5265,N_4884,N_4999);
nor U5266 (N_5266,N_4681,N_4790);
nor U5267 (N_5267,N_4981,N_4962);
or U5268 (N_5268,N_4738,N_4895);
nand U5269 (N_5269,N_4791,N_4882);
nor U5270 (N_5270,N_4878,N_4990);
and U5271 (N_5271,N_4730,N_4998);
xor U5272 (N_5272,N_4736,N_4943);
and U5273 (N_5273,N_4736,N_4782);
nand U5274 (N_5274,N_4727,N_4602);
nand U5275 (N_5275,N_4912,N_4510);
xnor U5276 (N_5276,N_4995,N_4764);
and U5277 (N_5277,N_4854,N_4836);
xnor U5278 (N_5278,N_4975,N_4558);
or U5279 (N_5279,N_4721,N_4629);
or U5280 (N_5280,N_4971,N_4838);
nand U5281 (N_5281,N_4705,N_4879);
nand U5282 (N_5282,N_4738,N_4820);
or U5283 (N_5283,N_4904,N_4833);
nor U5284 (N_5284,N_4863,N_4722);
or U5285 (N_5285,N_4999,N_4726);
nand U5286 (N_5286,N_4523,N_4660);
nand U5287 (N_5287,N_4873,N_4654);
xor U5288 (N_5288,N_4909,N_4886);
nand U5289 (N_5289,N_4547,N_4944);
nor U5290 (N_5290,N_4860,N_4603);
or U5291 (N_5291,N_4568,N_4730);
or U5292 (N_5292,N_4782,N_4627);
and U5293 (N_5293,N_4653,N_4508);
xor U5294 (N_5294,N_4766,N_4676);
nor U5295 (N_5295,N_4865,N_4956);
nor U5296 (N_5296,N_4866,N_4540);
and U5297 (N_5297,N_4922,N_4732);
and U5298 (N_5298,N_4802,N_4832);
xnor U5299 (N_5299,N_4915,N_4892);
nor U5300 (N_5300,N_4931,N_4720);
nand U5301 (N_5301,N_4774,N_4614);
or U5302 (N_5302,N_4651,N_4587);
xor U5303 (N_5303,N_4855,N_4652);
nand U5304 (N_5304,N_4540,N_4504);
nor U5305 (N_5305,N_4750,N_4947);
nor U5306 (N_5306,N_4895,N_4560);
nand U5307 (N_5307,N_4839,N_4614);
or U5308 (N_5308,N_4795,N_4802);
nor U5309 (N_5309,N_4709,N_4892);
xnor U5310 (N_5310,N_4742,N_4682);
nand U5311 (N_5311,N_4519,N_4675);
nand U5312 (N_5312,N_4940,N_4932);
nor U5313 (N_5313,N_4592,N_4841);
nand U5314 (N_5314,N_4701,N_4681);
nor U5315 (N_5315,N_4542,N_4603);
and U5316 (N_5316,N_4512,N_4680);
and U5317 (N_5317,N_4722,N_4690);
xor U5318 (N_5318,N_4530,N_4558);
nor U5319 (N_5319,N_4882,N_4658);
and U5320 (N_5320,N_4600,N_4993);
nand U5321 (N_5321,N_4848,N_4826);
or U5322 (N_5322,N_4780,N_4660);
and U5323 (N_5323,N_4640,N_4849);
and U5324 (N_5324,N_4543,N_4970);
nor U5325 (N_5325,N_4911,N_4864);
and U5326 (N_5326,N_4764,N_4847);
or U5327 (N_5327,N_4868,N_4650);
or U5328 (N_5328,N_4731,N_4604);
nand U5329 (N_5329,N_4692,N_4527);
nand U5330 (N_5330,N_4863,N_4690);
nand U5331 (N_5331,N_4630,N_4983);
xnor U5332 (N_5332,N_4862,N_4897);
nand U5333 (N_5333,N_4805,N_4939);
nor U5334 (N_5334,N_4631,N_4585);
xor U5335 (N_5335,N_4715,N_4525);
and U5336 (N_5336,N_4733,N_4684);
and U5337 (N_5337,N_4680,N_4572);
xor U5338 (N_5338,N_4755,N_4619);
nor U5339 (N_5339,N_4852,N_4651);
nor U5340 (N_5340,N_4973,N_4505);
xnor U5341 (N_5341,N_4527,N_4624);
nor U5342 (N_5342,N_4707,N_4890);
nand U5343 (N_5343,N_4555,N_4533);
or U5344 (N_5344,N_4713,N_4550);
or U5345 (N_5345,N_4574,N_4978);
xor U5346 (N_5346,N_4721,N_4898);
xnor U5347 (N_5347,N_4710,N_4564);
or U5348 (N_5348,N_4987,N_4994);
nand U5349 (N_5349,N_4846,N_4573);
or U5350 (N_5350,N_4892,N_4546);
and U5351 (N_5351,N_4766,N_4982);
nor U5352 (N_5352,N_4585,N_4559);
xor U5353 (N_5353,N_4603,N_4859);
nand U5354 (N_5354,N_4830,N_4862);
and U5355 (N_5355,N_4672,N_4899);
and U5356 (N_5356,N_4851,N_4781);
xor U5357 (N_5357,N_4978,N_4915);
or U5358 (N_5358,N_4508,N_4602);
and U5359 (N_5359,N_4830,N_4604);
nor U5360 (N_5360,N_4678,N_4933);
xor U5361 (N_5361,N_4660,N_4927);
nor U5362 (N_5362,N_4980,N_4605);
or U5363 (N_5363,N_4952,N_4566);
nand U5364 (N_5364,N_4858,N_4892);
or U5365 (N_5365,N_4617,N_4849);
nand U5366 (N_5366,N_4770,N_4959);
and U5367 (N_5367,N_4643,N_4535);
nor U5368 (N_5368,N_4547,N_4610);
and U5369 (N_5369,N_4799,N_4826);
or U5370 (N_5370,N_4886,N_4977);
xor U5371 (N_5371,N_4947,N_4897);
nor U5372 (N_5372,N_4548,N_4806);
xnor U5373 (N_5373,N_4965,N_4621);
nand U5374 (N_5374,N_4997,N_4823);
and U5375 (N_5375,N_4995,N_4745);
xor U5376 (N_5376,N_4888,N_4714);
nor U5377 (N_5377,N_4974,N_4909);
or U5378 (N_5378,N_4931,N_4579);
or U5379 (N_5379,N_4607,N_4941);
and U5380 (N_5380,N_4672,N_4677);
and U5381 (N_5381,N_4578,N_4597);
nand U5382 (N_5382,N_4911,N_4601);
or U5383 (N_5383,N_4688,N_4656);
or U5384 (N_5384,N_4862,N_4740);
and U5385 (N_5385,N_4546,N_4937);
xor U5386 (N_5386,N_4555,N_4918);
or U5387 (N_5387,N_4620,N_4610);
nand U5388 (N_5388,N_4885,N_4860);
nor U5389 (N_5389,N_4714,N_4767);
nor U5390 (N_5390,N_4772,N_4592);
nand U5391 (N_5391,N_4894,N_4582);
xor U5392 (N_5392,N_4818,N_4715);
or U5393 (N_5393,N_4956,N_4571);
nor U5394 (N_5394,N_4760,N_4638);
or U5395 (N_5395,N_4582,N_4802);
xor U5396 (N_5396,N_4816,N_4511);
or U5397 (N_5397,N_4895,N_4864);
xnor U5398 (N_5398,N_4898,N_4846);
nand U5399 (N_5399,N_4968,N_4596);
xor U5400 (N_5400,N_4641,N_4897);
and U5401 (N_5401,N_4529,N_4816);
and U5402 (N_5402,N_4540,N_4849);
xnor U5403 (N_5403,N_4679,N_4988);
nor U5404 (N_5404,N_4721,N_4514);
xor U5405 (N_5405,N_4720,N_4593);
or U5406 (N_5406,N_4628,N_4748);
nand U5407 (N_5407,N_4687,N_4960);
xor U5408 (N_5408,N_4600,N_4812);
or U5409 (N_5409,N_4915,N_4747);
xnor U5410 (N_5410,N_4566,N_4514);
nor U5411 (N_5411,N_4883,N_4568);
nand U5412 (N_5412,N_4818,N_4979);
nand U5413 (N_5413,N_4818,N_4850);
nor U5414 (N_5414,N_4592,N_4676);
and U5415 (N_5415,N_4629,N_4714);
nand U5416 (N_5416,N_4602,N_4643);
or U5417 (N_5417,N_4608,N_4925);
or U5418 (N_5418,N_4879,N_4805);
or U5419 (N_5419,N_4692,N_4771);
xor U5420 (N_5420,N_4986,N_4953);
xnor U5421 (N_5421,N_4914,N_4501);
nand U5422 (N_5422,N_4775,N_4992);
nand U5423 (N_5423,N_4839,N_4660);
nand U5424 (N_5424,N_4748,N_4601);
or U5425 (N_5425,N_4525,N_4798);
nor U5426 (N_5426,N_4667,N_4754);
and U5427 (N_5427,N_4980,N_4793);
or U5428 (N_5428,N_4668,N_4763);
or U5429 (N_5429,N_4668,N_4877);
xor U5430 (N_5430,N_4702,N_4824);
nand U5431 (N_5431,N_4898,N_4605);
and U5432 (N_5432,N_4513,N_4800);
or U5433 (N_5433,N_4518,N_4862);
nor U5434 (N_5434,N_4886,N_4887);
nor U5435 (N_5435,N_4983,N_4501);
or U5436 (N_5436,N_4668,N_4986);
nor U5437 (N_5437,N_4940,N_4876);
nand U5438 (N_5438,N_4966,N_4734);
nor U5439 (N_5439,N_4641,N_4922);
xnor U5440 (N_5440,N_4927,N_4500);
nand U5441 (N_5441,N_4655,N_4607);
xor U5442 (N_5442,N_4781,N_4555);
nor U5443 (N_5443,N_4890,N_4979);
and U5444 (N_5444,N_4646,N_4759);
and U5445 (N_5445,N_4993,N_4954);
and U5446 (N_5446,N_4834,N_4636);
nor U5447 (N_5447,N_4831,N_4833);
nand U5448 (N_5448,N_4942,N_4717);
and U5449 (N_5449,N_4539,N_4674);
nor U5450 (N_5450,N_4986,N_4584);
xor U5451 (N_5451,N_4771,N_4981);
or U5452 (N_5452,N_4502,N_4988);
nor U5453 (N_5453,N_4674,N_4550);
nand U5454 (N_5454,N_4569,N_4789);
nand U5455 (N_5455,N_4678,N_4763);
or U5456 (N_5456,N_4829,N_4920);
and U5457 (N_5457,N_4814,N_4514);
nor U5458 (N_5458,N_4871,N_4600);
nand U5459 (N_5459,N_4637,N_4764);
and U5460 (N_5460,N_4649,N_4971);
and U5461 (N_5461,N_4720,N_4505);
or U5462 (N_5462,N_4589,N_4663);
xor U5463 (N_5463,N_4779,N_4785);
nor U5464 (N_5464,N_4900,N_4830);
nor U5465 (N_5465,N_4651,N_4846);
nand U5466 (N_5466,N_4516,N_4773);
nand U5467 (N_5467,N_4695,N_4786);
xnor U5468 (N_5468,N_4958,N_4737);
or U5469 (N_5469,N_4628,N_4568);
nand U5470 (N_5470,N_4563,N_4884);
nor U5471 (N_5471,N_4615,N_4871);
nor U5472 (N_5472,N_4546,N_4914);
or U5473 (N_5473,N_4808,N_4641);
xnor U5474 (N_5474,N_4946,N_4843);
xnor U5475 (N_5475,N_4760,N_4689);
or U5476 (N_5476,N_4695,N_4563);
xor U5477 (N_5477,N_4628,N_4850);
xnor U5478 (N_5478,N_4700,N_4723);
xor U5479 (N_5479,N_4919,N_4546);
nand U5480 (N_5480,N_4941,N_4832);
and U5481 (N_5481,N_4880,N_4946);
nor U5482 (N_5482,N_4710,N_4750);
nor U5483 (N_5483,N_4510,N_4558);
or U5484 (N_5484,N_4723,N_4777);
or U5485 (N_5485,N_4647,N_4672);
or U5486 (N_5486,N_4841,N_4937);
and U5487 (N_5487,N_4593,N_4983);
xor U5488 (N_5488,N_4873,N_4783);
nor U5489 (N_5489,N_4669,N_4547);
nor U5490 (N_5490,N_4577,N_4516);
nor U5491 (N_5491,N_4980,N_4516);
or U5492 (N_5492,N_4800,N_4539);
xnor U5493 (N_5493,N_4874,N_4812);
nor U5494 (N_5494,N_4737,N_4778);
or U5495 (N_5495,N_4505,N_4901);
and U5496 (N_5496,N_4516,N_4519);
and U5497 (N_5497,N_4900,N_4954);
xnor U5498 (N_5498,N_4536,N_4550);
nor U5499 (N_5499,N_4614,N_4853);
xnor U5500 (N_5500,N_5331,N_5056);
or U5501 (N_5501,N_5475,N_5457);
and U5502 (N_5502,N_5008,N_5047);
xnor U5503 (N_5503,N_5435,N_5073);
or U5504 (N_5504,N_5308,N_5136);
nor U5505 (N_5505,N_5084,N_5251);
nand U5506 (N_5506,N_5454,N_5175);
xnor U5507 (N_5507,N_5300,N_5159);
xor U5508 (N_5508,N_5206,N_5348);
nor U5509 (N_5509,N_5384,N_5424);
xor U5510 (N_5510,N_5313,N_5123);
nor U5511 (N_5511,N_5138,N_5211);
and U5512 (N_5512,N_5403,N_5082);
nand U5513 (N_5513,N_5202,N_5328);
or U5514 (N_5514,N_5397,N_5061);
nor U5515 (N_5515,N_5385,N_5076);
nand U5516 (N_5516,N_5162,N_5189);
nor U5517 (N_5517,N_5223,N_5407);
xnor U5518 (N_5518,N_5441,N_5085);
xor U5519 (N_5519,N_5266,N_5222);
nor U5520 (N_5520,N_5366,N_5089);
nor U5521 (N_5521,N_5349,N_5421);
nand U5522 (N_5522,N_5121,N_5354);
nor U5523 (N_5523,N_5149,N_5039);
nor U5524 (N_5524,N_5356,N_5013);
or U5525 (N_5525,N_5399,N_5195);
and U5526 (N_5526,N_5321,N_5258);
xnor U5527 (N_5527,N_5074,N_5458);
or U5528 (N_5528,N_5370,N_5020);
or U5529 (N_5529,N_5193,N_5029);
and U5530 (N_5530,N_5323,N_5310);
xnor U5531 (N_5531,N_5271,N_5192);
nand U5532 (N_5532,N_5128,N_5405);
and U5533 (N_5533,N_5183,N_5163);
nand U5534 (N_5534,N_5104,N_5317);
nor U5535 (N_5535,N_5391,N_5048);
or U5536 (N_5536,N_5395,N_5040);
or U5537 (N_5537,N_5187,N_5083);
nand U5538 (N_5538,N_5101,N_5044);
nand U5539 (N_5539,N_5152,N_5248);
and U5540 (N_5540,N_5031,N_5135);
nor U5541 (N_5541,N_5446,N_5352);
nand U5542 (N_5542,N_5035,N_5282);
nand U5543 (N_5543,N_5332,N_5420);
xnor U5544 (N_5544,N_5108,N_5287);
nor U5545 (N_5545,N_5422,N_5151);
and U5546 (N_5546,N_5011,N_5296);
nand U5547 (N_5547,N_5176,N_5371);
and U5548 (N_5548,N_5463,N_5250);
and U5549 (N_5549,N_5431,N_5461);
nand U5550 (N_5550,N_5259,N_5239);
and U5551 (N_5551,N_5402,N_5179);
and U5552 (N_5552,N_5497,N_5148);
and U5553 (N_5553,N_5109,N_5276);
nor U5554 (N_5554,N_5460,N_5080);
and U5555 (N_5555,N_5156,N_5359);
xor U5556 (N_5556,N_5474,N_5233);
xor U5557 (N_5557,N_5380,N_5469);
and U5558 (N_5558,N_5488,N_5429);
nor U5559 (N_5559,N_5219,N_5462);
and U5560 (N_5560,N_5470,N_5477);
nand U5561 (N_5561,N_5117,N_5007);
nor U5562 (N_5562,N_5131,N_5476);
xor U5563 (N_5563,N_5303,N_5419);
nand U5564 (N_5564,N_5059,N_5180);
and U5565 (N_5565,N_5426,N_5245);
or U5566 (N_5566,N_5337,N_5344);
xnor U5567 (N_5567,N_5423,N_5122);
nor U5568 (N_5568,N_5124,N_5118);
or U5569 (N_5569,N_5342,N_5091);
nand U5570 (N_5570,N_5433,N_5097);
or U5571 (N_5571,N_5499,N_5267);
xor U5572 (N_5572,N_5238,N_5115);
nand U5573 (N_5573,N_5382,N_5137);
or U5574 (N_5574,N_5280,N_5291);
xnor U5575 (N_5575,N_5273,N_5191);
nand U5576 (N_5576,N_5498,N_5281);
nand U5577 (N_5577,N_5336,N_5496);
xnor U5578 (N_5578,N_5409,N_5357);
nor U5579 (N_5579,N_5075,N_5088);
and U5580 (N_5580,N_5350,N_5213);
and U5581 (N_5581,N_5042,N_5070);
or U5582 (N_5582,N_5130,N_5052);
and U5583 (N_5583,N_5066,N_5144);
and U5584 (N_5584,N_5404,N_5246);
nor U5585 (N_5585,N_5057,N_5335);
xnor U5586 (N_5586,N_5244,N_5270);
or U5587 (N_5587,N_5453,N_5069);
or U5588 (N_5588,N_5230,N_5120);
nor U5589 (N_5589,N_5025,N_5033);
and U5590 (N_5590,N_5418,N_5012);
nor U5591 (N_5591,N_5212,N_5214);
nand U5592 (N_5592,N_5171,N_5227);
nand U5593 (N_5593,N_5046,N_5347);
or U5594 (N_5594,N_5168,N_5215);
or U5595 (N_5595,N_5334,N_5298);
xor U5596 (N_5596,N_5071,N_5150);
nand U5597 (N_5597,N_5440,N_5134);
nor U5598 (N_5598,N_5002,N_5018);
or U5599 (N_5599,N_5217,N_5177);
and U5600 (N_5600,N_5229,N_5410);
xor U5601 (N_5601,N_5284,N_5480);
nor U5602 (N_5602,N_5486,N_5493);
xor U5603 (N_5603,N_5316,N_5448);
nand U5604 (N_5604,N_5314,N_5072);
xor U5605 (N_5605,N_5106,N_5203);
xor U5606 (N_5606,N_5079,N_5125);
or U5607 (N_5607,N_5093,N_5015);
nor U5608 (N_5608,N_5466,N_5096);
or U5609 (N_5609,N_5367,N_5145);
nand U5610 (N_5610,N_5484,N_5077);
or U5611 (N_5611,N_5318,N_5372);
xor U5612 (N_5612,N_5412,N_5110);
nand U5613 (N_5613,N_5197,N_5373);
nand U5614 (N_5614,N_5247,N_5165);
or U5615 (N_5615,N_5242,N_5041);
or U5616 (N_5616,N_5100,N_5050);
xnor U5617 (N_5617,N_5283,N_5343);
and U5618 (N_5618,N_5058,N_5028);
and U5619 (N_5619,N_5388,N_5140);
nand U5620 (N_5620,N_5322,N_5293);
nand U5621 (N_5621,N_5302,N_5139);
and U5622 (N_5622,N_5290,N_5026);
xor U5623 (N_5623,N_5174,N_5155);
and U5624 (N_5624,N_5425,N_5232);
and U5625 (N_5625,N_5414,N_5260);
or U5626 (N_5626,N_5051,N_5286);
nor U5627 (N_5627,N_5235,N_5309);
and U5628 (N_5628,N_5236,N_5451);
or U5629 (N_5629,N_5208,N_5173);
nor U5630 (N_5630,N_5369,N_5487);
xor U5631 (N_5631,N_5377,N_5167);
nor U5632 (N_5632,N_5274,N_5320);
nand U5633 (N_5633,N_5311,N_5434);
nor U5634 (N_5634,N_5494,N_5065);
nor U5635 (N_5635,N_5225,N_5439);
nand U5636 (N_5636,N_5182,N_5471);
nor U5637 (N_5637,N_5060,N_5416);
xor U5638 (N_5638,N_5216,N_5081);
nor U5639 (N_5639,N_5181,N_5201);
and U5640 (N_5640,N_5237,N_5262);
or U5641 (N_5641,N_5278,N_5301);
and U5642 (N_5642,N_5055,N_5408);
nand U5643 (N_5643,N_5030,N_5207);
nand U5644 (N_5644,N_5333,N_5447);
nand U5645 (N_5645,N_5263,N_5415);
nand U5646 (N_5646,N_5194,N_5036);
nor U5647 (N_5647,N_5492,N_5147);
or U5648 (N_5648,N_5143,N_5275);
and U5649 (N_5649,N_5024,N_5126);
and U5650 (N_5650,N_5034,N_5010);
nor U5651 (N_5651,N_5406,N_5022);
nand U5652 (N_5652,N_5456,N_5345);
and U5653 (N_5653,N_5430,N_5315);
xnor U5654 (N_5654,N_5205,N_5411);
and U5655 (N_5655,N_5053,N_5252);
nor U5656 (N_5656,N_5132,N_5285);
nor U5657 (N_5657,N_5129,N_5340);
nand U5658 (N_5658,N_5390,N_5043);
and U5659 (N_5659,N_5133,N_5325);
nand U5660 (N_5660,N_5054,N_5491);
xnor U5661 (N_5661,N_5188,N_5166);
and U5662 (N_5662,N_5383,N_5210);
or U5663 (N_5663,N_5063,N_5226);
nand U5664 (N_5664,N_5398,N_5319);
nand U5665 (N_5665,N_5221,N_5360);
xor U5666 (N_5666,N_5339,N_5127);
nor U5667 (N_5667,N_5114,N_5169);
nand U5668 (N_5668,N_5467,N_5363);
nand U5669 (N_5669,N_5170,N_5037);
xnor U5670 (N_5670,N_5307,N_5241);
nand U5671 (N_5671,N_5001,N_5160);
nor U5672 (N_5672,N_5358,N_5164);
xor U5673 (N_5673,N_5338,N_5396);
xor U5674 (N_5674,N_5468,N_5279);
and U5675 (N_5675,N_5378,N_5346);
and U5676 (N_5676,N_5087,N_5204);
xnor U5677 (N_5677,N_5142,N_5253);
and U5678 (N_5678,N_5107,N_5368);
and U5679 (N_5679,N_5449,N_5341);
nand U5680 (N_5680,N_5220,N_5218);
xor U5681 (N_5681,N_5436,N_5005);
and U5682 (N_5682,N_5090,N_5200);
or U5683 (N_5683,N_5393,N_5009);
nand U5684 (N_5684,N_5444,N_5428);
and U5685 (N_5685,N_5157,N_5224);
nor U5686 (N_5686,N_5269,N_5092);
and U5687 (N_5687,N_5495,N_5019);
or U5688 (N_5688,N_5400,N_5437);
and U5689 (N_5689,N_5254,N_5021);
or U5690 (N_5690,N_5361,N_5099);
nand U5691 (N_5691,N_5146,N_5261);
nand U5692 (N_5692,N_5016,N_5459);
or U5693 (N_5693,N_5199,N_5288);
nor U5694 (N_5694,N_5299,N_5153);
xor U5695 (N_5695,N_5249,N_5105);
xnor U5696 (N_5696,N_5038,N_5228);
nor U5697 (N_5697,N_5098,N_5374);
nand U5698 (N_5698,N_5489,N_5004);
nor U5699 (N_5699,N_5113,N_5478);
and U5700 (N_5700,N_5362,N_5443);
xor U5701 (N_5701,N_5243,N_5067);
xnor U5702 (N_5702,N_5234,N_5389);
xnor U5703 (N_5703,N_5394,N_5268);
xnor U5704 (N_5704,N_5032,N_5103);
or U5705 (N_5705,N_5294,N_5330);
and U5706 (N_5706,N_5094,N_5112);
nor U5707 (N_5707,N_5483,N_5184);
xor U5708 (N_5708,N_5095,N_5353);
nor U5709 (N_5709,N_5473,N_5161);
and U5710 (N_5710,N_5386,N_5329);
nand U5711 (N_5711,N_5265,N_5485);
and U5712 (N_5712,N_5379,N_5185);
and U5713 (N_5713,N_5027,N_5365);
nand U5714 (N_5714,N_5045,N_5141);
nor U5715 (N_5715,N_5376,N_5445);
nor U5716 (N_5716,N_5427,N_5375);
nand U5717 (N_5717,N_5006,N_5438);
xor U5718 (N_5718,N_5351,N_5064);
nor U5719 (N_5719,N_5327,N_5178);
xnor U5720 (N_5720,N_5240,N_5479);
xnor U5721 (N_5721,N_5387,N_5472);
nand U5722 (N_5722,N_5190,N_5464);
nand U5723 (N_5723,N_5003,N_5401);
nor U5724 (N_5724,N_5086,N_5014);
nand U5725 (N_5725,N_5102,N_5304);
xor U5726 (N_5726,N_5000,N_5417);
nand U5727 (N_5727,N_5272,N_5255);
and U5728 (N_5728,N_5306,N_5289);
and U5729 (N_5729,N_5381,N_5465);
or U5730 (N_5730,N_5119,N_5442);
nand U5731 (N_5731,N_5116,N_5324);
xnor U5732 (N_5732,N_5297,N_5062);
nor U5733 (N_5733,N_5209,N_5256);
and U5734 (N_5734,N_5312,N_5264);
and U5735 (N_5735,N_5482,N_5413);
nor U5736 (N_5736,N_5432,N_5305);
or U5737 (N_5737,N_5158,N_5111);
nor U5738 (N_5738,N_5292,N_5490);
nand U5739 (N_5739,N_5257,N_5049);
xor U5740 (N_5740,N_5172,N_5452);
xor U5741 (N_5741,N_5326,N_5295);
xor U5742 (N_5742,N_5023,N_5078);
or U5743 (N_5743,N_5198,N_5154);
or U5744 (N_5744,N_5392,N_5455);
nor U5745 (N_5745,N_5196,N_5355);
nor U5746 (N_5746,N_5231,N_5277);
nor U5747 (N_5747,N_5017,N_5481);
and U5748 (N_5748,N_5186,N_5364);
nor U5749 (N_5749,N_5068,N_5450);
nand U5750 (N_5750,N_5276,N_5495);
or U5751 (N_5751,N_5283,N_5269);
xor U5752 (N_5752,N_5074,N_5040);
nand U5753 (N_5753,N_5182,N_5073);
nor U5754 (N_5754,N_5138,N_5309);
and U5755 (N_5755,N_5109,N_5006);
or U5756 (N_5756,N_5244,N_5482);
or U5757 (N_5757,N_5396,N_5189);
nor U5758 (N_5758,N_5051,N_5170);
or U5759 (N_5759,N_5068,N_5353);
and U5760 (N_5760,N_5331,N_5493);
xnor U5761 (N_5761,N_5474,N_5217);
or U5762 (N_5762,N_5155,N_5267);
and U5763 (N_5763,N_5013,N_5190);
xnor U5764 (N_5764,N_5258,N_5157);
nand U5765 (N_5765,N_5180,N_5091);
and U5766 (N_5766,N_5048,N_5195);
nand U5767 (N_5767,N_5252,N_5103);
nor U5768 (N_5768,N_5030,N_5217);
and U5769 (N_5769,N_5052,N_5162);
or U5770 (N_5770,N_5424,N_5138);
or U5771 (N_5771,N_5111,N_5488);
nor U5772 (N_5772,N_5353,N_5261);
xor U5773 (N_5773,N_5026,N_5211);
and U5774 (N_5774,N_5351,N_5393);
and U5775 (N_5775,N_5178,N_5013);
and U5776 (N_5776,N_5417,N_5132);
nor U5777 (N_5777,N_5127,N_5324);
nor U5778 (N_5778,N_5116,N_5286);
nand U5779 (N_5779,N_5093,N_5162);
nand U5780 (N_5780,N_5054,N_5249);
or U5781 (N_5781,N_5458,N_5264);
xor U5782 (N_5782,N_5135,N_5335);
or U5783 (N_5783,N_5469,N_5379);
or U5784 (N_5784,N_5432,N_5157);
or U5785 (N_5785,N_5441,N_5201);
and U5786 (N_5786,N_5365,N_5055);
nand U5787 (N_5787,N_5252,N_5340);
nor U5788 (N_5788,N_5360,N_5282);
or U5789 (N_5789,N_5027,N_5244);
nand U5790 (N_5790,N_5227,N_5205);
or U5791 (N_5791,N_5209,N_5215);
and U5792 (N_5792,N_5370,N_5348);
xnor U5793 (N_5793,N_5492,N_5486);
or U5794 (N_5794,N_5411,N_5091);
nor U5795 (N_5795,N_5438,N_5367);
nor U5796 (N_5796,N_5150,N_5017);
nand U5797 (N_5797,N_5153,N_5143);
and U5798 (N_5798,N_5328,N_5438);
and U5799 (N_5799,N_5192,N_5118);
or U5800 (N_5800,N_5190,N_5469);
and U5801 (N_5801,N_5195,N_5166);
or U5802 (N_5802,N_5399,N_5025);
and U5803 (N_5803,N_5156,N_5228);
or U5804 (N_5804,N_5475,N_5043);
and U5805 (N_5805,N_5189,N_5176);
and U5806 (N_5806,N_5148,N_5313);
xor U5807 (N_5807,N_5004,N_5397);
or U5808 (N_5808,N_5470,N_5411);
nor U5809 (N_5809,N_5460,N_5286);
nand U5810 (N_5810,N_5127,N_5353);
or U5811 (N_5811,N_5343,N_5187);
xnor U5812 (N_5812,N_5093,N_5376);
nor U5813 (N_5813,N_5056,N_5369);
nor U5814 (N_5814,N_5437,N_5373);
or U5815 (N_5815,N_5252,N_5035);
and U5816 (N_5816,N_5380,N_5489);
xnor U5817 (N_5817,N_5373,N_5005);
and U5818 (N_5818,N_5173,N_5270);
xor U5819 (N_5819,N_5190,N_5444);
nor U5820 (N_5820,N_5336,N_5133);
xor U5821 (N_5821,N_5018,N_5341);
nand U5822 (N_5822,N_5045,N_5152);
xor U5823 (N_5823,N_5332,N_5494);
or U5824 (N_5824,N_5455,N_5287);
or U5825 (N_5825,N_5292,N_5119);
and U5826 (N_5826,N_5109,N_5191);
xnor U5827 (N_5827,N_5441,N_5115);
xor U5828 (N_5828,N_5421,N_5321);
xor U5829 (N_5829,N_5407,N_5153);
xor U5830 (N_5830,N_5291,N_5273);
xor U5831 (N_5831,N_5112,N_5414);
nand U5832 (N_5832,N_5278,N_5215);
nor U5833 (N_5833,N_5050,N_5059);
nor U5834 (N_5834,N_5296,N_5353);
or U5835 (N_5835,N_5092,N_5256);
or U5836 (N_5836,N_5036,N_5421);
and U5837 (N_5837,N_5157,N_5250);
nand U5838 (N_5838,N_5417,N_5034);
or U5839 (N_5839,N_5486,N_5434);
nor U5840 (N_5840,N_5296,N_5304);
nand U5841 (N_5841,N_5335,N_5028);
nand U5842 (N_5842,N_5410,N_5268);
and U5843 (N_5843,N_5335,N_5053);
xor U5844 (N_5844,N_5195,N_5321);
nand U5845 (N_5845,N_5161,N_5423);
nand U5846 (N_5846,N_5155,N_5226);
xor U5847 (N_5847,N_5303,N_5131);
or U5848 (N_5848,N_5147,N_5171);
nor U5849 (N_5849,N_5410,N_5119);
and U5850 (N_5850,N_5229,N_5240);
xor U5851 (N_5851,N_5333,N_5336);
or U5852 (N_5852,N_5375,N_5470);
nand U5853 (N_5853,N_5342,N_5152);
nor U5854 (N_5854,N_5398,N_5470);
nand U5855 (N_5855,N_5256,N_5407);
xor U5856 (N_5856,N_5000,N_5378);
xnor U5857 (N_5857,N_5034,N_5499);
and U5858 (N_5858,N_5437,N_5039);
or U5859 (N_5859,N_5357,N_5385);
xor U5860 (N_5860,N_5423,N_5146);
nor U5861 (N_5861,N_5469,N_5241);
nor U5862 (N_5862,N_5087,N_5297);
or U5863 (N_5863,N_5356,N_5345);
nor U5864 (N_5864,N_5178,N_5130);
and U5865 (N_5865,N_5136,N_5479);
or U5866 (N_5866,N_5325,N_5462);
nor U5867 (N_5867,N_5367,N_5272);
or U5868 (N_5868,N_5191,N_5141);
xor U5869 (N_5869,N_5446,N_5230);
or U5870 (N_5870,N_5315,N_5078);
and U5871 (N_5871,N_5239,N_5335);
xnor U5872 (N_5872,N_5451,N_5036);
or U5873 (N_5873,N_5133,N_5407);
or U5874 (N_5874,N_5457,N_5231);
and U5875 (N_5875,N_5143,N_5301);
nor U5876 (N_5876,N_5324,N_5254);
nor U5877 (N_5877,N_5065,N_5426);
nor U5878 (N_5878,N_5458,N_5200);
or U5879 (N_5879,N_5073,N_5258);
nor U5880 (N_5880,N_5333,N_5151);
or U5881 (N_5881,N_5325,N_5369);
nand U5882 (N_5882,N_5154,N_5182);
xnor U5883 (N_5883,N_5365,N_5428);
and U5884 (N_5884,N_5192,N_5140);
nand U5885 (N_5885,N_5170,N_5144);
and U5886 (N_5886,N_5469,N_5175);
nand U5887 (N_5887,N_5239,N_5461);
xor U5888 (N_5888,N_5425,N_5070);
nor U5889 (N_5889,N_5046,N_5382);
xor U5890 (N_5890,N_5130,N_5095);
xnor U5891 (N_5891,N_5325,N_5099);
or U5892 (N_5892,N_5016,N_5344);
and U5893 (N_5893,N_5125,N_5215);
nor U5894 (N_5894,N_5058,N_5387);
or U5895 (N_5895,N_5338,N_5491);
or U5896 (N_5896,N_5019,N_5330);
nand U5897 (N_5897,N_5198,N_5300);
or U5898 (N_5898,N_5484,N_5082);
nand U5899 (N_5899,N_5398,N_5158);
nand U5900 (N_5900,N_5416,N_5390);
and U5901 (N_5901,N_5473,N_5456);
and U5902 (N_5902,N_5200,N_5375);
nand U5903 (N_5903,N_5182,N_5432);
and U5904 (N_5904,N_5193,N_5150);
or U5905 (N_5905,N_5404,N_5046);
and U5906 (N_5906,N_5194,N_5416);
or U5907 (N_5907,N_5315,N_5147);
and U5908 (N_5908,N_5085,N_5277);
nand U5909 (N_5909,N_5213,N_5064);
or U5910 (N_5910,N_5207,N_5231);
or U5911 (N_5911,N_5363,N_5498);
or U5912 (N_5912,N_5465,N_5018);
and U5913 (N_5913,N_5213,N_5280);
xnor U5914 (N_5914,N_5464,N_5033);
xnor U5915 (N_5915,N_5078,N_5464);
xnor U5916 (N_5916,N_5371,N_5292);
or U5917 (N_5917,N_5326,N_5213);
nor U5918 (N_5918,N_5460,N_5320);
or U5919 (N_5919,N_5496,N_5315);
xor U5920 (N_5920,N_5105,N_5174);
nand U5921 (N_5921,N_5026,N_5340);
nand U5922 (N_5922,N_5033,N_5498);
nand U5923 (N_5923,N_5434,N_5210);
and U5924 (N_5924,N_5078,N_5299);
nor U5925 (N_5925,N_5084,N_5057);
nand U5926 (N_5926,N_5279,N_5246);
xor U5927 (N_5927,N_5441,N_5154);
nor U5928 (N_5928,N_5145,N_5187);
xor U5929 (N_5929,N_5259,N_5033);
nand U5930 (N_5930,N_5433,N_5435);
and U5931 (N_5931,N_5403,N_5339);
or U5932 (N_5932,N_5491,N_5117);
or U5933 (N_5933,N_5329,N_5077);
or U5934 (N_5934,N_5299,N_5280);
or U5935 (N_5935,N_5273,N_5131);
and U5936 (N_5936,N_5039,N_5297);
xnor U5937 (N_5937,N_5040,N_5032);
or U5938 (N_5938,N_5237,N_5334);
nor U5939 (N_5939,N_5222,N_5462);
xnor U5940 (N_5940,N_5090,N_5023);
nor U5941 (N_5941,N_5191,N_5144);
and U5942 (N_5942,N_5075,N_5430);
and U5943 (N_5943,N_5023,N_5225);
nand U5944 (N_5944,N_5260,N_5433);
and U5945 (N_5945,N_5477,N_5300);
and U5946 (N_5946,N_5179,N_5141);
and U5947 (N_5947,N_5257,N_5137);
and U5948 (N_5948,N_5227,N_5496);
nor U5949 (N_5949,N_5238,N_5430);
nor U5950 (N_5950,N_5434,N_5363);
nor U5951 (N_5951,N_5379,N_5472);
and U5952 (N_5952,N_5281,N_5114);
nand U5953 (N_5953,N_5188,N_5302);
xor U5954 (N_5954,N_5252,N_5207);
or U5955 (N_5955,N_5271,N_5012);
xor U5956 (N_5956,N_5311,N_5147);
and U5957 (N_5957,N_5323,N_5096);
nor U5958 (N_5958,N_5096,N_5239);
xnor U5959 (N_5959,N_5134,N_5066);
xnor U5960 (N_5960,N_5436,N_5393);
nor U5961 (N_5961,N_5310,N_5053);
and U5962 (N_5962,N_5298,N_5287);
and U5963 (N_5963,N_5196,N_5294);
xor U5964 (N_5964,N_5436,N_5197);
xnor U5965 (N_5965,N_5462,N_5133);
xor U5966 (N_5966,N_5075,N_5061);
nand U5967 (N_5967,N_5019,N_5290);
nand U5968 (N_5968,N_5068,N_5495);
nor U5969 (N_5969,N_5491,N_5027);
xor U5970 (N_5970,N_5398,N_5466);
or U5971 (N_5971,N_5308,N_5001);
or U5972 (N_5972,N_5400,N_5446);
nor U5973 (N_5973,N_5168,N_5101);
or U5974 (N_5974,N_5108,N_5400);
xnor U5975 (N_5975,N_5013,N_5419);
nand U5976 (N_5976,N_5181,N_5112);
nor U5977 (N_5977,N_5042,N_5134);
xor U5978 (N_5978,N_5346,N_5034);
nor U5979 (N_5979,N_5055,N_5313);
nand U5980 (N_5980,N_5396,N_5381);
and U5981 (N_5981,N_5358,N_5360);
and U5982 (N_5982,N_5482,N_5028);
or U5983 (N_5983,N_5495,N_5013);
nand U5984 (N_5984,N_5374,N_5031);
nor U5985 (N_5985,N_5256,N_5415);
nand U5986 (N_5986,N_5456,N_5290);
nor U5987 (N_5987,N_5047,N_5182);
or U5988 (N_5988,N_5300,N_5004);
or U5989 (N_5989,N_5204,N_5086);
and U5990 (N_5990,N_5210,N_5094);
or U5991 (N_5991,N_5059,N_5194);
or U5992 (N_5992,N_5044,N_5332);
or U5993 (N_5993,N_5048,N_5005);
or U5994 (N_5994,N_5009,N_5118);
nand U5995 (N_5995,N_5158,N_5439);
xor U5996 (N_5996,N_5435,N_5087);
and U5997 (N_5997,N_5071,N_5422);
or U5998 (N_5998,N_5231,N_5370);
nor U5999 (N_5999,N_5012,N_5299);
nor U6000 (N_6000,N_5786,N_5704);
or U6001 (N_6001,N_5512,N_5524);
nor U6002 (N_6002,N_5963,N_5563);
and U6003 (N_6003,N_5811,N_5867);
or U6004 (N_6004,N_5924,N_5598);
or U6005 (N_6005,N_5666,N_5604);
nand U6006 (N_6006,N_5667,N_5987);
and U6007 (N_6007,N_5925,N_5671);
or U6008 (N_6008,N_5640,N_5908);
or U6009 (N_6009,N_5892,N_5961);
and U6010 (N_6010,N_5968,N_5787);
and U6011 (N_6011,N_5834,N_5506);
or U6012 (N_6012,N_5941,N_5803);
xnor U6013 (N_6013,N_5639,N_5986);
xor U6014 (N_6014,N_5675,N_5656);
nor U6015 (N_6015,N_5958,N_5648);
and U6016 (N_6016,N_5757,N_5553);
nand U6017 (N_6017,N_5505,N_5678);
and U6018 (N_6018,N_5770,N_5607);
xnor U6019 (N_6019,N_5875,N_5818);
and U6020 (N_6020,N_5830,N_5694);
nand U6021 (N_6021,N_5647,N_5576);
or U6022 (N_6022,N_5765,N_5882);
nor U6023 (N_6023,N_5885,N_5521);
xnor U6024 (N_6024,N_5832,N_5580);
or U6025 (N_6025,N_5767,N_5546);
xnor U6026 (N_6026,N_5616,N_5964);
xnor U6027 (N_6027,N_5884,N_5582);
nor U6028 (N_6028,N_5862,N_5898);
xor U6029 (N_6029,N_5539,N_5680);
nand U6030 (N_6030,N_5936,N_5500);
xor U6031 (N_6031,N_5516,N_5703);
nor U6032 (N_6032,N_5706,N_5802);
and U6033 (N_6033,N_5722,N_5838);
or U6034 (N_6034,N_5782,N_5552);
nor U6035 (N_6035,N_5890,N_5816);
or U6036 (N_6036,N_5612,N_5744);
xor U6037 (N_6037,N_5940,N_5550);
or U6038 (N_6038,N_5949,N_5798);
xnor U6039 (N_6039,N_5724,N_5950);
nor U6040 (N_6040,N_5689,N_5507);
and U6041 (N_6041,N_5651,N_5823);
nand U6042 (N_6042,N_5778,N_5502);
nand U6043 (N_6043,N_5855,N_5526);
xnor U6044 (N_6044,N_5727,N_5754);
nand U6045 (N_6045,N_5808,N_5942);
and U6046 (N_6046,N_5641,N_5791);
xnor U6047 (N_6047,N_5804,N_5827);
nor U6048 (N_6048,N_5794,N_5980);
nand U6049 (N_6049,N_5899,N_5917);
nand U6050 (N_6050,N_5895,N_5870);
xor U6051 (N_6051,N_5685,N_5698);
nor U6052 (N_6052,N_5509,N_5849);
nand U6053 (N_6053,N_5708,N_5932);
nor U6054 (N_6054,N_5730,N_5565);
or U6055 (N_6055,N_5726,N_5902);
nand U6056 (N_6056,N_5764,N_5945);
xor U6057 (N_6057,N_5682,N_5531);
nor U6058 (N_6058,N_5982,N_5904);
or U6059 (N_6059,N_5971,N_5631);
xor U6060 (N_6060,N_5959,N_5906);
nand U6061 (N_6061,N_5714,N_5723);
xnor U6062 (N_6062,N_5985,N_5688);
nor U6063 (N_6063,N_5807,N_5579);
nor U6064 (N_6064,N_5934,N_5707);
nor U6065 (N_6065,N_5684,N_5621);
or U6066 (N_6066,N_5900,N_5789);
xnor U6067 (N_6067,N_5594,N_5777);
nor U6068 (N_6068,N_5881,N_5624);
nand U6069 (N_6069,N_5872,N_5545);
nand U6070 (N_6070,N_5728,N_5756);
nand U6071 (N_6071,N_5812,N_5622);
and U6072 (N_6072,N_5913,N_5837);
or U6073 (N_6073,N_5790,N_5847);
and U6074 (N_6074,N_5608,N_5910);
nand U6075 (N_6075,N_5646,N_5976);
xor U6076 (N_6076,N_5712,N_5629);
nand U6077 (N_6077,N_5541,N_5610);
nand U6078 (N_6078,N_5783,N_5909);
or U6079 (N_6079,N_5713,N_5876);
xnor U6080 (N_6080,N_5717,N_5508);
nand U6081 (N_6081,N_5916,N_5681);
nor U6082 (N_6082,N_5861,N_5831);
nor U6083 (N_6083,N_5519,N_5788);
nor U6084 (N_6084,N_5809,N_5795);
nand U6085 (N_6085,N_5729,N_5822);
nor U6086 (N_6086,N_5709,N_5522);
xor U6087 (N_6087,N_5634,N_5653);
nand U6088 (N_6088,N_5743,N_5753);
xor U6089 (N_6089,N_5567,N_5981);
or U6090 (N_6090,N_5623,N_5548);
nor U6091 (N_6091,N_5915,N_5746);
nor U6092 (N_6092,N_5762,N_5953);
xor U6093 (N_6093,N_5537,N_5679);
nor U6094 (N_6094,N_5814,N_5673);
xor U6095 (N_6095,N_5735,N_5990);
nand U6096 (N_6096,N_5926,N_5905);
nor U6097 (N_6097,N_5829,N_5805);
nor U6098 (N_6098,N_5701,N_5687);
or U6099 (N_6099,N_5853,N_5815);
nand U6100 (N_6100,N_5768,N_5935);
or U6101 (N_6101,N_5965,N_5585);
nor U6102 (N_6102,N_5600,N_5865);
nand U6103 (N_6103,N_5590,N_5931);
and U6104 (N_6104,N_5535,N_5650);
xor U6105 (N_6105,N_5561,N_5760);
and U6106 (N_6106,N_5530,N_5578);
or U6107 (N_6107,N_5896,N_5742);
and U6108 (N_6108,N_5668,N_5903);
and U6109 (N_6109,N_5967,N_5540);
or U6110 (N_6110,N_5683,N_5700);
and U6111 (N_6111,N_5752,N_5996);
nand U6112 (N_6112,N_5891,N_5711);
nor U6113 (N_6113,N_5715,N_5551);
xor U6114 (N_6114,N_5674,N_5588);
xor U6115 (N_6115,N_5843,N_5658);
xor U6116 (N_6116,N_5605,N_5549);
xnor U6117 (N_6117,N_5560,N_5930);
nand U6118 (N_6118,N_5532,N_5574);
and U6119 (N_6119,N_5997,N_5810);
nor U6120 (N_6120,N_5611,N_5763);
or U6121 (N_6121,N_5866,N_5973);
xor U6122 (N_6122,N_5873,N_5970);
and U6123 (N_6123,N_5864,N_5796);
and U6124 (N_6124,N_5785,N_5586);
and U6125 (N_6125,N_5557,N_5773);
or U6126 (N_6126,N_5920,N_5633);
and U6127 (N_6127,N_5797,N_5665);
or U6128 (N_6128,N_5569,N_5937);
or U6129 (N_6129,N_5625,N_5840);
nand U6130 (N_6130,N_5741,N_5676);
or U6131 (N_6131,N_5564,N_5523);
and U6132 (N_6132,N_5793,N_5856);
xnor U6133 (N_6133,N_5533,N_5734);
and U6134 (N_6134,N_5589,N_5609);
nand U6135 (N_6135,N_5614,N_5771);
nor U6136 (N_6136,N_5852,N_5897);
nand U6137 (N_6137,N_5591,N_5697);
nor U6138 (N_6138,N_5740,N_5543);
and U6139 (N_6139,N_5806,N_5846);
xnor U6140 (N_6140,N_5739,N_5718);
and U6141 (N_6141,N_5946,N_5755);
and U6142 (N_6142,N_5517,N_5725);
nor U6143 (N_6143,N_5692,N_5738);
nand U6144 (N_6144,N_5603,N_5780);
xnor U6145 (N_6145,N_5836,N_5649);
nor U6146 (N_6146,N_5962,N_5869);
or U6147 (N_6147,N_5800,N_5766);
nor U6148 (N_6148,N_5593,N_5716);
nand U6149 (N_6149,N_5630,N_5581);
nand U6150 (N_6150,N_5660,N_5690);
nand U6151 (N_6151,N_5880,N_5907);
xor U6152 (N_6152,N_5599,N_5542);
or U6153 (N_6153,N_5914,N_5955);
xnor U6154 (N_6154,N_5878,N_5637);
xnor U6155 (N_6155,N_5960,N_5994);
nor U6156 (N_6156,N_5799,N_5828);
or U6157 (N_6157,N_5943,N_5670);
or U6158 (N_6158,N_5922,N_5558);
and U6159 (N_6159,N_5613,N_5520);
nand U6160 (N_6160,N_5559,N_5615);
and U6161 (N_6161,N_5825,N_5860);
and U6162 (N_6162,N_5669,N_5619);
xnor U6163 (N_6163,N_5995,N_5721);
xor U6164 (N_6164,N_5720,N_5759);
or U6165 (N_6165,N_5501,N_5868);
and U6166 (N_6166,N_5606,N_5748);
and U6167 (N_6167,N_5538,N_5951);
or U6168 (N_6168,N_5626,N_5632);
or U6169 (N_6169,N_5732,N_5979);
or U6170 (N_6170,N_5877,N_5528);
xnor U6171 (N_6171,N_5652,N_5657);
nor U6172 (N_6172,N_5597,N_5525);
or U6173 (N_6173,N_5779,N_5655);
and U6174 (N_6174,N_5912,N_5643);
or U6175 (N_6175,N_5894,N_5555);
and U6176 (N_6176,N_5737,N_5601);
or U6177 (N_6177,N_5554,N_5989);
or U6178 (N_6178,N_5664,N_5845);
and U6179 (N_6179,N_5999,N_5850);
nand U6180 (N_6180,N_5929,N_5644);
nor U6181 (N_6181,N_5954,N_5772);
nor U6182 (N_6182,N_5693,N_5957);
or U6183 (N_6183,N_5663,N_5817);
nand U6184 (N_6184,N_5504,N_5536);
or U6185 (N_6185,N_5848,N_5889);
nor U6186 (N_6186,N_5747,N_5696);
xor U6187 (N_6187,N_5736,N_5901);
and U6188 (N_6188,N_5705,N_5887);
nor U6189 (N_6189,N_5769,N_5577);
or U6190 (N_6190,N_5514,N_5571);
or U6191 (N_6191,N_5731,N_5833);
xor U6192 (N_6192,N_5749,N_5515);
nand U6193 (N_6193,N_5911,N_5819);
nand U6194 (N_6194,N_5928,N_5984);
or U6195 (N_6195,N_5854,N_5662);
nand U6196 (N_6196,N_5863,N_5774);
or U6197 (N_6197,N_5826,N_5975);
nor U6198 (N_6198,N_5570,N_5992);
nor U6199 (N_6199,N_5627,N_5851);
nand U6200 (N_6200,N_5620,N_5886);
nand U6201 (N_6201,N_5839,N_5820);
nand U6202 (N_6202,N_5801,N_5733);
or U6203 (N_6203,N_5952,N_5991);
nor U6204 (N_6204,N_5792,N_5584);
xnor U6205 (N_6205,N_5587,N_5510);
and U6206 (N_6206,N_5672,N_5842);
nand U6207 (N_6207,N_5874,N_5919);
nand U6208 (N_6208,N_5661,N_5617);
nand U6209 (N_6209,N_5939,N_5921);
nand U6210 (N_6210,N_5947,N_5974);
nand U6211 (N_6211,N_5927,N_5978);
nand U6212 (N_6212,N_5998,N_5750);
nor U6213 (N_6213,N_5977,N_5858);
xor U6214 (N_6214,N_5879,N_5654);
and U6215 (N_6215,N_5710,N_5602);
nand U6216 (N_6216,N_5691,N_5751);
or U6217 (N_6217,N_5595,N_5758);
nor U6218 (N_6218,N_5642,N_5956);
or U6219 (N_6219,N_5871,N_5699);
nand U6220 (N_6220,N_5993,N_5966);
or U6221 (N_6221,N_5572,N_5969);
nor U6222 (N_6222,N_5659,N_5888);
nor U6223 (N_6223,N_5562,N_5583);
nand U6224 (N_6224,N_5781,N_5635);
nor U6225 (N_6225,N_5547,N_5841);
nand U6226 (N_6226,N_5859,N_5776);
and U6227 (N_6227,N_5972,N_5566);
nor U6228 (N_6228,N_5628,N_5592);
and U6229 (N_6229,N_5518,N_5784);
xnor U6230 (N_6230,N_5775,N_5702);
xnor U6231 (N_6231,N_5645,N_5824);
nand U6232 (N_6232,N_5933,N_5618);
nor U6233 (N_6233,N_5638,N_5948);
nor U6234 (N_6234,N_5527,N_5983);
nor U6235 (N_6235,N_5556,N_5568);
nand U6236 (N_6236,N_5677,N_5695);
nor U6237 (N_6237,N_5529,N_5883);
and U6238 (N_6238,N_5686,N_5944);
nand U6239 (N_6239,N_5761,N_5857);
nand U6240 (N_6240,N_5893,N_5636);
or U6241 (N_6241,N_5719,N_5573);
nor U6242 (N_6242,N_5835,N_5821);
or U6243 (N_6243,N_5844,N_5534);
nand U6244 (N_6244,N_5503,N_5513);
nand U6245 (N_6245,N_5918,N_5544);
nor U6246 (N_6246,N_5575,N_5596);
nor U6247 (N_6247,N_5511,N_5938);
or U6248 (N_6248,N_5745,N_5813);
nor U6249 (N_6249,N_5988,N_5923);
nand U6250 (N_6250,N_5946,N_5753);
xor U6251 (N_6251,N_5709,N_5993);
and U6252 (N_6252,N_5745,N_5853);
or U6253 (N_6253,N_5862,N_5804);
or U6254 (N_6254,N_5791,N_5670);
or U6255 (N_6255,N_5521,N_5897);
xor U6256 (N_6256,N_5890,N_5824);
and U6257 (N_6257,N_5607,N_5949);
and U6258 (N_6258,N_5949,N_5801);
nand U6259 (N_6259,N_5976,N_5529);
or U6260 (N_6260,N_5600,N_5859);
xor U6261 (N_6261,N_5881,N_5591);
or U6262 (N_6262,N_5572,N_5592);
and U6263 (N_6263,N_5596,N_5776);
and U6264 (N_6264,N_5995,N_5860);
or U6265 (N_6265,N_5614,N_5992);
xor U6266 (N_6266,N_5678,N_5641);
nor U6267 (N_6267,N_5567,N_5686);
xnor U6268 (N_6268,N_5707,N_5970);
nand U6269 (N_6269,N_5667,N_5803);
and U6270 (N_6270,N_5635,N_5520);
nand U6271 (N_6271,N_5723,N_5855);
or U6272 (N_6272,N_5559,N_5732);
nor U6273 (N_6273,N_5732,N_5534);
xor U6274 (N_6274,N_5514,N_5612);
or U6275 (N_6275,N_5767,N_5534);
nor U6276 (N_6276,N_5756,N_5808);
or U6277 (N_6277,N_5592,N_5811);
or U6278 (N_6278,N_5673,N_5630);
or U6279 (N_6279,N_5972,N_5821);
and U6280 (N_6280,N_5750,N_5596);
or U6281 (N_6281,N_5876,N_5549);
and U6282 (N_6282,N_5507,N_5505);
and U6283 (N_6283,N_5660,N_5981);
xnor U6284 (N_6284,N_5845,N_5506);
xnor U6285 (N_6285,N_5675,N_5867);
nor U6286 (N_6286,N_5775,N_5721);
xnor U6287 (N_6287,N_5935,N_5934);
and U6288 (N_6288,N_5634,N_5794);
nand U6289 (N_6289,N_5966,N_5956);
nand U6290 (N_6290,N_5526,N_5606);
and U6291 (N_6291,N_5709,N_5902);
nand U6292 (N_6292,N_5790,N_5551);
nor U6293 (N_6293,N_5600,N_5793);
xnor U6294 (N_6294,N_5659,N_5865);
nor U6295 (N_6295,N_5533,N_5763);
and U6296 (N_6296,N_5683,N_5713);
nor U6297 (N_6297,N_5620,N_5529);
nor U6298 (N_6298,N_5998,N_5586);
xor U6299 (N_6299,N_5617,N_5646);
and U6300 (N_6300,N_5731,N_5561);
or U6301 (N_6301,N_5550,N_5787);
xor U6302 (N_6302,N_5836,N_5639);
and U6303 (N_6303,N_5574,N_5776);
nand U6304 (N_6304,N_5568,N_5711);
and U6305 (N_6305,N_5845,N_5990);
nand U6306 (N_6306,N_5884,N_5871);
nand U6307 (N_6307,N_5789,N_5807);
and U6308 (N_6308,N_5702,N_5670);
nand U6309 (N_6309,N_5806,N_5769);
xnor U6310 (N_6310,N_5581,N_5719);
nand U6311 (N_6311,N_5536,N_5842);
and U6312 (N_6312,N_5583,N_5906);
and U6313 (N_6313,N_5519,N_5711);
nor U6314 (N_6314,N_5568,N_5691);
xor U6315 (N_6315,N_5866,N_5855);
xnor U6316 (N_6316,N_5972,N_5636);
nand U6317 (N_6317,N_5735,N_5780);
xor U6318 (N_6318,N_5606,N_5618);
or U6319 (N_6319,N_5851,N_5633);
nor U6320 (N_6320,N_5519,N_5932);
and U6321 (N_6321,N_5569,N_5686);
nor U6322 (N_6322,N_5535,N_5670);
xnor U6323 (N_6323,N_5521,N_5649);
and U6324 (N_6324,N_5820,N_5874);
xor U6325 (N_6325,N_5736,N_5546);
or U6326 (N_6326,N_5780,N_5632);
nand U6327 (N_6327,N_5633,N_5570);
xnor U6328 (N_6328,N_5609,N_5754);
or U6329 (N_6329,N_5524,N_5875);
xor U6330 (N_6330,N_5681,N_5960);
nor U6331 (N_6331,N_5634,N_5603);
xor U6332 (N_6332,N_5696,N_5773);
nand U6333 (N_6333,N_5594,N_5869);
nand U6334 (N_6334,N_5965,N_5603);
nand U6335 (N_6335,N_5645,N_5558);
nor U6336 (N_6336,N_5596,N_5692);
or U6337 (N_6337,N_5902,N_5830);
nand U6338 (N_6338,N_5801,N_5701);
nand U6339 (N_6339,N_5884,N_5623);
or U6340 (N_6340,N_5545,N_5787);
xor U6341 (N_6341,N_5549,N_5723);
xor U6342 (N_6342,N_5994,N_5910);
xor U6343 (N_6343,N_5991,N_5995);
or U6344 (N_6344,N_5934,N_5700);
nor U6345 (N_6345,N_5908,N_5810);
nor U6346 (N_6346,N_5639,N_5587);
nor U6347 (N_6347,N_5591,N_5580);
xnor U6348 (N_6348,N_5809,N_5783);
nand U6349 (N_6349,N_5770,N_5611);
and U6350 (N_6350,N_5536,N_5778);
or U6351 (N_6351,N_5627,N_5520);
nand U6352 (N_6352,N_5741,N_5695);
nand U6353 (N_6353,N_5962,N_5519);
xor U6354 (N_6354,N_5560,N_5730);
and U6355 (N_6355,N_5962,N_5532);
or U6356 (N_6356,N_5789,N_5671);
xor U6357 (N_6357,N_5552,N_5841);
nand U6358 (N_6358,N_5527,N_5696);
and U6359 (N_6359,N_5917,N_5619);
xnor U6360 (N_6360,N_5533,N_5514);
nor U6361 (N_6361,N_5874,N_5965);
or U6362 (N_6362,N_5508,N_5934);
nand U6363 (N_6363,N_5650,N_5777);
xor U6364 (N_6364,N_5759,N_5557);
nand U6365 (N_6365,N_5844,N_5653);
nor U6366 (N_6366,N_5725,N_5873);
nand U6367 (N_6367,N_5666,N_5738);
nand U6368 (N_6368,N_5837,N_5826);
or U6369 (N_6369,N_5687,N_5613);
nand U6370 (N_6370,N_5620,N_5524);
and U6371 (N_6371,N_5563,N_5513);
nand U6372 (N_6372,N_5769,N_5903);
nor U6373 (N_6373,N_5926,N_5956);
or U6374 (N_6374,N_5739,N_5616);
or U6375 (N_6375,N_5844,N_5669);
or U6376 (N_6376,N_5852,N_5647);
nor U6377 (N_6377,N_5587,N_5707);
nand U6378 (N_6378,N_5916,N_5619);
and U6379 (N_6379,N_5695,N_5610);
nand U6380 (N_6380,N_5792,N_5838);
or U6381 (N_6381,N_5682,N_5701);
or U6382 (N_6382,N_5593,N_5533);
nand U6383 (N_6383,N_5870,N_5621);
xor U6384 (N_6384,N_5658,N_5577);
nand U6385 (N_6385,N_5585,N_5605);
or U6386 (N_6386,N_5940,N_5782);
and U6387 (N_6387,N_5706,N_5753);
nand U6388 (N_6388,N_5555,N_5969);
or U6389 (N_6389,N_5585,N_5547);
xnor U6390 (N_6390,N_5762,N_5826);
xor U6391 (N_6391,N_5676,N_5906);
nand U6392 (N_6392,N_5640,N_5629);
and U6393 (N_6393,N_5866,N_5653);
nor U6394 (N_6394,N_5548,N_5904);
or U6395 (N_6395,N_5547,N_5827);
nand U6396 (N_6396,N_5823,N_5502);
or U6397 (N_6397,N_5782,N_5673);
nor U6398 (N_6398,N_5575,N_5878);
nand U6399 (N_6399,N_5540,N_5787);
nor U6400 (N_6400,N_5675,N_5913);
nor U6401 (N_6401,N_5993,N_5914);
and U6402 (N_6402,N_5986,N_5782);
and U6403 (N_6403,N_5960,N_5757);
nand U6404 (N_6404,N_5621,N_5958);
nor U6405 (N_6405,N_5959,N_5609);
or U6406 (N_6406,N_5984,N_5840);
nor U6407 (N_6407,N_5974,N_5831);
nand U6408 (N_6408,N_5528,N_5586);
nand U6409 (N_6409,N_5875,N_5866);
and U6410 (N_6410,N_5742,N_5653);
and U6411 (N_6411,N_5796,N_5834);
or U6412 (N_6412,N_5725,N_5992);
xnor U6413 (N_6413,N_5698,N_5972);
or U6414 (N_6414,N_5615,N_5992);
or U6415 (N_6415,N_5753,N_5908);
nor U6416 (N_6416,N_5520,N_5973);
nand U6417 (N_6417,N_5926,N_5566);
nor U6418 (N_6418,N_5764,N_5532);
nor U6419 (N_6419,N_5723,N_5986);
or U6420 (N_6420,N_5517,N_5978);
and U6421 (N_6421,N_5927,N_5622);
xor U6422 (N_6422,N_5956,N_5570);
or U6423 (N_6423,N_5833,N_5584);
nor U6424 (N_6424,N_5595,N_5726);
nand U6425 (N_6425,N_5860,N_5844);
or U6426 (N_6426,N_5728,N_5733);
nor U6427 (N_6427,N_5632,N_5505);
xor U6428 (N_6428,N_5892,N_5905);
nand U6429 (N_6429,N_5960,N_5724);
xnor U6430 (N_6430,N_5559,N_5554);
or U6431 (N_6431,N_5889,N_5749);
or U6432 (N_6432,N_5630,N_5650);
nand U6433 (N_6433,N_5715,N_5632);
nor U6434 (N_6434,N_5540,N_5997);
and U6435 (N_6435,N_5820,N_5854);
xor U6436 (N_6436,N_5855,N_5934);
nand U6437 (N_6437,N_5972,N_5764);
nor U6438 (N_6438,N_5988,N_5530);
or U6439 (N_6439,N_5519,N_5921);
nand U6440 (N_6440,N_5715,N_5566);
nor U6441 (N_6441,N_5569,N_5528);
or U6442 (N_6442,N_5775,N_5546);
or U6443 (N_6443,N_5682,N_5510);
nand U6444 (N_6444,N_5985,N_5832);
nor U6445 (N_6445,N_5922,N_5673);
and U6446 (N_6446,N_5682,N_5518);
or U6447 (N_6447,N_5543,N_5588);
nand U6448 (N_6448,N_5550,N_5833);
nor U6449 (N_6449,N_5852,N_5963);
or U6450 (N_6450,N_5836,N_5928);
xor U6451 (N_6451,N_5829,N_5510);
xnor U6452 (N_6452,N_5738,N_5755);
and U6453 (N_6453,N_5668,N_5854);
and U6454 (N_6454,N_5716,N_5767);
nor U6455 (N_6455,N_5772,N_5709);
and U6456 (N_6456,N_5629,N_5979);
or U6457 (N_6457,N_5721,N_5852);
xnor U6458 (N_6458,N_5804,N_5882);
and U6459 (N_6459,N_5841,N_5641);
or U6460 (N_6460,N_5815,N_5854);
nor U6461 (N_6461,N_5941,N_5892);
and U6462 (N_6462,N_5937,N_5578);
or U6463 (N_6463,N_5900,N_5669);
xor U6464 (N_6464,N_5654,N_5975);
or U6465 (N_6465,N_5514,N_5719);
or U6466 (N_6466,N_5816,N_5725);
or U6467 (N_6467,N_5598,N_5863);
or U6468 (N_6468,N_5665,N_5766);
nor U6469 (N_6469,N_5903,N_5647);
xor U6470 (N_6470,N_5852,N_5851);
xnor U6471 (N_6471,N_5654,N_5998);
nand U6472 (N_6472,N_5638,N_5763);
xor U6473 (N_6473,N_5959,N_5933);
nor U6474 (N_6474,N_5981,N_5522);
nand U6475 (N_6475,N_5852,N_5774);
or U6476 (N_6476,N_5975,N_5762);
or U6477 (N_6477,N_5764,N_5503);
and U6478 (N_6478,N_5752,N_5883);
nor U6479 (N_6479,N_5998,N_5719);
nor U6480 (N_6480,N_5624,N_5585);
and U6481 (N_6481,N_5942,N_5757);
xor U6482 (N_6482,N_5822,N_5539);
and U6483 (N_6483,N_5780,N_5838);
and U6484 (N_6484,N_5546,N_5961);
xnor U6485 (N_6485,N_5989,N_5602);
or U6486 (N_6486,N_5871,N_5912);
or U6487 (N_6487,N_5710,N_5981);
nor U6488 (N_6488,N_5989,N_5794);
nand U6489 (N_6489,N_5669,N_5575);
or U6490 (N_6490,N_5621,N_5991);
nor U6491 (N_6491,N_5949,N_5796);
nand U6492 (N_6492,N_5862,N_5521);
or U6493 (N_6493,N_5740,N_5847);
xor U6494 (N_6494,N_5816,N_5747);
and U6495 (N_6495,N_5642,N_5831);
or U6496 (N_6496,N_5583,N_5675);
nand U6497 (N_6497,N_5500,N_5784);
or U6498 (N_6498,N_5802,N_5738);
xor U6499 (N_6499,N_5970,N_5860);
xnor U6500 (N_6500,N_6170,N_6205);
nor U6501 (N_6501,N_6386,N_6220);
and U6502 (N_6502,N_6338,N_6060);
nor U6503 (N_6503,N_6106,N_6454);
xnor U6504 (N_6504,N_6270,N_6400);
nor U6505 (N_6505,N_6376,N_6112);
and U6506 (N_6506,N_6153,N_6159);
or U6507 (N_6507,N_6490,N_6459);
nor U6508 (N_6508,N_6033,N_6450);
nand U6509 (N_6509,N_6413,N_6453);
nand U6510 (N_6510,N_6421,N_6337);
or U6511 (N_6511,N_6438,N_6240);
nor U6512 (N_6512,N_6175,N_6384);
and U6513 (N_6513,N_6061,N_6396);
and U6514 (N_6514,N_6293,N_6040);
nor U6515 (N_6515,N_6072,N_6285);
xor U6516 (N_6516,N_6388,N_6404);
nor U6517 (N_6517,N_6176,N_6377);
or U6518 (N_6518,N_6474,N_6251);
xnor U6519 (N_6519,N_6158,N_6408);
or U6520 (N_6520,N_6050,N_6335);
nand U6521 (N_6521,N_6369,N_6044);
nor U6522 (N_6522,N_6314,N_6137);
nand U6523 (N_6523,N_6020,N_6464);
nand U6524 (N_6524,N_6218,N_6317);
nor U6525 (N_6525,N_6245,N_6009);
or U6526 (N_6526,N_6300,N_6206);
or U6527 (N_6527,N_6208,N_6244);
xor U6528 (N_6528,N_6344,N_6414);
or U6529 (N_6529,N_6423,N_6179);
nand U6530 (N_6530,N_6315,N_6046);
or U6531 (N_6531,N_6417,N_6307);
nor U6532 (N_6532,N_6177,N_6378);
nand U6533 (N_6533,N_6134,N_6135);
nor U6534 (N_6534,N_6447,N_6083);
nand U6535 (N_6535,N_6405,N_6120);
nor U6536 (N_6536,N_6019,N_6368);
or U6537 (N_6537,N_6157,N_6451);
nand U6538 (N_6538,N_6483,N_6036);
nor U6539 (N_6539,N_6362,N_6077);
or U6540 (N_6540,N_6457,N_6006);
xnor U6541 (N_6541,N_6074,N_6243);
nor U6542 (N_6542,N_6139,N_6445);
and U6543 (N_6543,N_6308,N_6233);
xnor U6544 (N_6544,N_6493,N_6041);
xnor U6545 (N_6545,N_6299,N_6099);
xnor U6546 (N_6546,N_6105,N_6221);
and U6547 (N_6547,N_6320,N_6318);
xnor U6548 (N_6548,N_6169,N_6427);
xor U6549 (N_6549,N_6316,N_6002);
and U6550 (N_6550,N_6121,N_6382);
nor U6551 (N_6551,N_6183,N_6097);
xnor U6552 (N_6552,N_6212,N_6489);
and U6553 (N_6553,N_6287,N_6387);
or U6554 (N_6554,N_6096,N_6101);
nor U6555 (N_6555,N_6323,N_6154);
nand U6556 (N_6556,N_6406,N_6273);
nand U6557 (N_6557,N_6392,N_6381);
nand U6558 (N_6558,N_6425,N_6086);
nor U6559 (N_6559,N_6032,N_6108);
and U6560 (N_6560,N_6194,N_6217);
nand U6561 (N_6561,N_6491,N_6255);
or U6562 (N_6562,N_6286,N_6012);
xor U6563 (N_6563,N_6219,N_6042);
or U6564 (N_6564,N_6391,N_6264);
xor U6565 (N_6565,N_6340,N_6082);
or U6566 (N_6566,N_6399,N_6262);
nor U6567 (N_6567,N_6276,N_6141);
xor U6568 (N_6568,N_6089,N_6258);
nor U6569 (N_6569,N_6215,N_6067);
nand U6570 (N_6570,N_6346,N_6347);
nor U6571 (N_6571,N_6052,N_6291);
xnor U6572 (N_6572,N_6011,N_6229);
nor U6573 (N_6573,N_6479,N_6203);
or U6574 (N_6574,N_6094,N_6225);
nand U6575 (N_6575,N_6207,N_6301);
and U6576 (N_6576,N_6448,N_6186);
nor U6577 (N_6577,N_6172,N_6202);
and U6578 (N_6578,N_6100,N_6075);
or U6579 (N_6579,N_6003,N_6305);
or U6580 (N_6580,N_6357,N_6265);
and U6581 (N_6581,N_6419,N_6263);
or U6582 (N_6582,N_6260,N_6237);
nand U6583 (N_6583,N_6222,N_6339);
xnor U6584 (N_6584,N_6071,N_6107);
nand U6585 (N_6585,N_6185,N_6336);
xnor U6586 (N_6586,N_6252,N_6268);
xor U6587 (N_6587,N_6168,N_6138);
nand U6588 (N_6588,N_6480,N_6295);
xor U6589 (N_6589,N_6238,N_6296);
nor U6590 (N_6590,N_6443,N_6472);
and U6591 (N_6591,N_6231,N_6038);
nor U6592 (N_6592,N_6239,N_6210);
and U6593 (N_6593,N_6224,N_6005);
nand U6594 (N_6594,N_6484,N_6250);
nand U6595 (N_6595,N_6469,N_6078);
xor U6596 (N_6596,N_6156,N_6363);
nand U6597 (N_6597,N_6364,N_6371);
and U6598 (N_6598,N_6351,N_6193);
and U6599 (N_6599,N_6066,N_6249);
nand U6600 (N_6600,N_6087,N_6465);
xnor U6601 (N_6601,N_6290,N_6113);
nand U6602 (N_6602,N_6434,N_6494);
nor U6603 (N_6603,N_6393,N_6298);
nand U6604 (N_6604,N_6487,N_6282);
and U6605 (N_6605,N_6467,N_6326);
or U6606 (N_6606,N_6345,N_6014);
nor U6607 (N_6607,N_6095,N_6349);
or U6608 (N_6608,N_6028,N_6160);
nand U6609 (N_6609,N_6354,N_6063);
or U6610 (N_6610,N_6155,N_6246);
nor U6611 (N_6611,N_6361,N_6182);
nor U6612 (N_6612,N_6328,N_6021);
and U6613 (N_6613,N_6166,N_6189);
and U6614 (N_6614,N_6482,N_6211);
nor U6615 (N_6615,N_6178,N_6279);
or U6616 (N_6616,N_6247,N_6394);
nor U6617 (N_6617,N_6327,N_6149);
and U6618 (N_6618,N_6267,N_6226);
and U6619 (N_6619,N_6277,N_6288);
or U6620 (N_6620,N_6254,N_6026);
nand U6621 (N_6621,N_6410,N_6111);
and U6622 (N_6622,N_6025,N_6248);
and U6623 (N_6623,N_6214,N_6034);
or U6624 (N_6624,N_6365,N_6131);
or U6625 (N_6625,N_6147,N_6124);
or U6626 (N_6626,N_6426,N_6302);
or U6627 (N_6627,N_6356,N_6303);
xnor U6628 (N_6628,N_6462,N_6115);
or U6629 (N_6629,N_6043,N_6125);
nand U6630 (N_6630,N_6098,N_6440);
xnor U6631 (N_6631,N_6027,N_6397);
nand U6632 (N_6632,N_6016,N_6059);
nand U6633 (N_6633,N_6281,N_6306);
nand U6634 (N_6634,N_6437,N_6433);
nor U6635 (N_6635,N_6353,N_6294);
nor U6636 (N_6636,N_6054,N_6085);
nor U6637 (N_6637,N_6280,N_6039);
nor U6638 (N_6638,N_6004,N_6379);
xnor U6639 (N_6639,N_6058,N_6062);
nor U6640 (N_6640,N_6242,N_6259);
nor U6641 (N_6641,N_6374,N_6133);
nor U6642 (N_6642,N_6411,N_6236);
xnor U6643 (N_6643,N_6056,N_6395);
nor U6644 (N_6644,N_6496,N_6123);
nand U6645 (N_6645,N_6477,N_6117);
nor U6646 (N_6646,N_6495,N_6190);
and U6647 (N_6647,N_6241,N_6102);
nor U6648 (N_6648,N_6209,N_6136);
or U6649 (N_6649,N_6430,N_6227);
xor U6650 (N_6650,N_6180,N_6035);
xor U6651 (N_6651,N_6455,N_6162);
or U6652 (N_6652,N_6367,N_6142);
nor U6653 (N_6653,N_6132,N_6412);
and U6654 (N_6654,N_6171,N_6080);
nor U6655 (N_6655,N_6128,N_6010);
or U6656 (N_6656,N_6278,N_6081);
nand U6657 (N_6657,N_6029,N_6053);
and U6658 (N_6658,N_6311,N_6272);
and U6659 (N_6659,N_6390,N_6069);
and U6660 (N_6660,N_6380,N_6199);
nand U6661 (N_6661,N_6332,N_6329);
xor U6662 (N_6662,N_6116,N_6372);
xnor U6663 (N_6663,N_6140,N_6184);
or U6664 (N_6664,N_6070,N_6045);
or U6665 (N_6665,N_6325,N_6119);
xor U6666 (N_6666,N_6065,N_6449);
or U6667 (N_6667,N_6313,N_6271);
nand U6668 (N_6668,N_6073,N_6167);
or U6669 (N_6669,N_6018,N_6321);
and U6670 (N_6670,N_6331,N_6144);
nor U6671 (N_6671,N_6151,N_6103);
or U6672 (N_6672,N_6358,N_6261);
or U6673 (N_6673,N_6407,N_6256);
nand U6674 (N_6674,N_6463,N_6492);
nand U6675 (N_6675,N_6352,N_6173);
xnor U6676 (N_6676,N_6422,N_6235);
xnor U6677 (N_6677,N_6370,N_6476);
xor U6678 (N_6678,N_6499,N_6359);
nor U6679 (N_6679,N_6130,N_6230);
xnor U6680 (N_6680,N_6297,N_6442);
or U6681 (N_6681,N_6275,N_6164);
and U6682 (N_6682,N_6234,N_6401);
or U6683 (N_6683,N_6109,N_6415);
xnor U6684 (N_6684,N_6037,N_6228);
xnor U6685 (N_6685,N_6441,N_6129);
nand U6686 (N_6686,N_6030,N_6204);
or U6687 (N_6687,N_6418,N_6047);
nand U6688 (N_6688,N_6200,N_6497);
and U6689 (N_6689,N_6051,N_6334);
or U6690 (N_6690,N_6192,N_6283);
nand U6691 (N_6691,N_6452,N_6486);
or U6692 (N_6692,N_6289,N_6092);
nand U6693 (N_6693,N_6429,N_6017);
xor U6694 (N_6694,N_6161,N_6436);
and U6695 (N_6695,N_6064,N_6284);
nand U6696 (N_6696,N_6481,N_6145);
or U6697 (N_6697,N_6090,N_6439);
or U6698 (N_6698,N_6084,N_6000);
nand U6699 (N_6699,N_6428,N_6118);
nor U6700 (N_6700,N_6435,N_6188);
or U6701 (N_6701,N_6324,N_6485);
xnor U6702 (N_6702,N_6126,N_6104);
and U6703 (N_6703,N_6431,N_6383);
xor U6704 (N_6704,N_6389,N_6091);
or U6705 (N_6705,N_6402,N_6478);
nand U6706 (N_6706,N_6165,N_6048);
nand U6707 (N_6707,N_6488,N_6322);
nor U6708 (N_6708,N_6456,N_6470);
nand U6709 (N_6709,N_6163,N_6055);
nand U6710 (N_6710,N_6187,N_6350);
xnor U6711 (N_6711,N_6348,N_6355);
nand U6712 (N_6712,N_6181,N_6057);
nand U6713 (N_6713,N_6253,N_6023);
nor U6714 (N_6714,N_6013,N_6198);
and U6715 (N_6715,N_6174,N_6269);
nand U6716 (N_6716,N_6446,N_6197);
nand U6717 (N_6717,N_6498,N_6143);
nand U6718 (N_6718,N_6385,N_6444);
nor U6719 (N_6719,N_6424,N_6148);
or U6720 (N_6720,N_6319,N_6150);
xnor U6721 (N_6721,N_6232,N_6460);
or U6722 (N_6722,N_6398,N_6432);
nand U6723 (N_6723,N_6146,N_6152);
and U6724 (N_6724,N_6360,N_6195);
xnor U6725 (N_6725,N_6088,N_6015);
and U6726 (N_6726,N_6274,N_6373);
nand U6727 (N_6727,N_6471,N_6416);
or U6728 (N_6728,N_6473,N_6366);
nor U6729 (N_6729,N_6223,N_6409);
nor U6730 (N_6730,N_6341,N_6466);
or U6731 (N_6731,N_6213,N_6342);
nor U6732 (N_6732,N_6312,N_6110);
xnor U6733 (N_6733,N_6022,N_6266);
nor U6734 (N_6734,N_6304,N_6093);
or U6735 (N_6735,N_6257,N_6375);
xnor U6736 (N_6736,N_6333,N_6403);
xor U6737 (N_6737,N_6475,N_6458);
nand U6738 (N_6738,N_6201,N_6196);
and U6739 (N_6739,N_6127,N_6008);
nor U6740 (N_6740,N_6309,N_6024);
xor U6741 (N_6741,N_6310,N_6191);
xnor U6742 (N_6742,N_6216,N_6330);
nand U6743 (N_6743,N_6049,N_6343);
xnor U6744 (N_6744,N_6068,N_6076);
xor U6745 (N_6745,N_6079,N_6122);
xor U6746 (N_6746,N_6292,N_6468);
nor U6747 (N_6747,N_6461,N_6420);
nor U6748 (N_6748,N_6114,N_6001);
nand U6749 (N_6749,N_6031,N_6007);
nor U6750 (N_6750,N_6256,N_6493);
xnor U6751 (N_6751,N_6348,N_6295);
nor U6752 (N_6752,N_6283,N_6393);
or U6753 (N_6753,N_6151,N_6399);
or U6754 (N_6754,N_6456,N_6210);
nor U6755 (N_6755,N_6293,N_6085);
or U6756 (N_6756,N_6146,N_6371);
or U6757 (N_6757,N_6469,N_6345);
xnor U6758 (N_6758,N_6172,N_6068);
xnor U6759 (N_6759,N_6200,N_6381);
nand U6760 (N_6760,N_6155,N_6283);
xor U6761 (N_6761,N_6050,N_6463);
or U6762 (N_6762,N_6389,N_6018);
nor U6763 (N_6763,N_6460,N_6340);
nand U6764 (N_6764,N_6089,N_6002);
or U6765 (N_6765,N_6439,N_6242);
or U6766 (N_6766,N_6234,N_6336);
nand U6767 (N_6767,N_6264,N_6412);
or U6768 (N_6768,N_6249,N_6297);
and U6769 (N_6769,N_6121,N_6256);
or U6770 (N_6770,N_6046,N_6025);
nor U6771 (N_6771,N_6234,N_6125);
nand U6772 (N_6772,N_6077,N_6472);
nor U6773 (N_6773,N_6091,N_6054);
or U6774 (N_6774,N_6393,N_6008);
and U6775 (N_6775,N_6105,N_6347);
nor U6776 (N_6776,N_6266,N_6438);
xor U6777 (N_6777,N_6489,N_6349);
nand U6778 (N_6778,N_6242,N_6306);
and U6779 (N_6779,N_6336,N_6005);
and U6780 (N_6780,N_6203,N_6464);
nand U6781 (N_6781,N_6195,N_6499);
and U6782 (N_6782,N_6267,N_6386);
or U6783 (N_6783,N_6330,N_6335);
xor U6784 (N_6784,N_6107,N_6122);
or U6785 (N_6785,N_6469,N_6193);
or U6786 (N_6786,N_6258,N_6086);
xnor U6787 (N_6787,N_6264,N_6437);
xor U6788 (N_6788,N_6224,N_6080);
nand U6789 (N_6789,N_6234,N_6074);
xor U6790 (N_6790,N_6192,N_6411);
nand U6791 (N_6791,N_6227,N_6399);
xor U6792 (N_6792,N_6223,N_6029);
or U6793 (N_6793,N_6261,N_6458);
and U6794 (N_6794,N_6359,N_6381);
or U6795 (N_6795,N_6260,N_6490);
or U6796 (N_6796,N_6293,N_6308);
nand U6797 (N_6797,N_6122,N_6046);
or U6798 (N_6798,N_6130,N_6170);
or U6799 (N_6799,N_6020,N_6322);
and U6800 (N_6800,N_6147,N_6250);
xnor U6801 (N_6801,N_6047,N_6116);
xnor U6802 (N_6802,N_6282,N_6204);
and U6803 (N_6803,N_6142,N_6429);
xnor U6804 (N_6804,N_6228,N_6436);
nor U6805 (N_6805,N_6097,N_6408);
xnor U6806 (N_6806,N_6426,N_6022);
or U6807 (N_6807,N_6190,N_6209);
nor U6808 (N_6808,N_6334,N_6147);
xor U6809 (N_6809,N_6427,N_6152);
and U6810 (N_6810,N_6147,N_6388);
or U6811 (N_6811,N_6239,N_6456);
nor U6812 (N_6812,N_6057,N_6104);
nor U6813 (N_6813,N_6232,N_6287);
xnor U6814 (N_6814,N_6425,N_6431);
and U6815 (N_6815,N_6320,N_6362);
nand U6816 (N_6816,N_6409,N_6114);
or U6817 (N_6817,N_6141,N_6494);
or U6818 (N_6818,N_6198,N_6110);
and U6819 (N_6819,N_6164,N_6000);
or U6820 (N_6820,N_6311,N_6187);
nand U6821 (N_6821,N_6327,N_6035);
nand U6822 (N_6822,N_6233,N_6386);
or U6823 (N_6823,N_6244,N_6022);
nand U6824 (N_6824,N_6454,N_6431);
and U6825 (N_6825,N_6052,N_6101);
xnor U6826 (N_6826,N_6413,N_6298);
xnor U6827 (N_6827,N_6066,N_6187);
or U6828 (N_6828,N_6138,N_6319);
or U6829 (N_6829,N_6392,N_6041);
or U6830 (N_6830,N_6034,N_6479);
nand U6831 (N_6831,N_6136,N_6034);
nand U6832 (N_6832,N_6475,N_6080);
xor U6833 (N_6833,N_6265,N_6295);
xor U6834 (N_6834,N_6375,N_6294);
nand U6835 (N_6835,N_6284,N_6287);
or U6836 (N_6836,N_6319,N_6125);
or U6837 (N_6837,N_6290,N_6436);
nand U6838 (N_6838,N_6154,N_6162);
and U6839 (N_6839,N_6178,N_6027);
nor U6840 (N_6840,N_6121,N_6162);
and U6841 (N_6841,N_6108,N_6085);
nor U6842 (N_6842,N_6470,N_6432);
nor U6843 (N_6843,N_6412,N_6088);
or U6844 (N_6844,N_6016,N_6092);
and U6845 (N_6845,N_6033,N_6120);
and U6846 (N_6846,N_6330,N_6082);
nand U6847 (N_6847,N_6186,N_6091);
and U6848 (N_6848,N_6178,N_6433);
xor U6849 (N_6849,N_6023,N_6283);
or U6850 (N_6850,N_6469,N_6431);
nand U6851 (N_6851,N_6473,N_6094);
or U6852 (N_6852,N_6181,N_6480);
and U6853 (N_6853,N_6098,N_6339);
xnor U6854 (N_6854,N_6480,N_6373);
nor U6855 (N_6855,N_6483,N_6277);
xnor U6856 (N_6856,N_6018,N_6107);
nor U6857 (N_6857,N_6013,N_6355);
nand U6858 (N_6858,N_6436,N_6409);
and U6859 (N_6859,N_6373,N_6471);
and U6860 (N_6860,N_6179,N_6366);
nand U6861 (N_6861,N_6373,N_6295);
nor U6862 (N_6862,N_6257,N_6318);
nand U6863 (N_6863,N_6155,N_6334);
or U6864 (N_6864,N_6013,N_6031);
nor U6865 (N_6865,N_6274,N_6119);
nand U6866 (N_6866,N_6243,N_6099);
xnor U6867 (N_6867,N_6491,N_6379);
nor U6868 (N_6868,N_6072,N_6014);
and U6869 (N_6869,N_6383,N_6437);
nor U6870 (N_6870,N_6065,N_6091);
and U6871 (N_6871,N_6438,N_6279);
nor U6872 (N_6872,N_6459,N_6257);
nand U6873 (N_6873,N_6388,N_6208);
or U6874 (N_6874,N_6306,N_6084);
and U6875 (N_6875,N_6256,N_6464);
or U6876 (N_6876,N_6309,N_6281);
or U6877 (N_6877,N_6321,N_6392);
or U6878 (N_6878,N_6340,N_6093);
xnor U6879 (N_6879,N_6379,N_6425);
or U6880 (N_6880,N_6286,N_6324);
xor U6881 (N_6881,N_6255,N_6381);
and U6882 (N_6882,N_6143,N_6094);
nor U6883 (N_6883,N_6123,N_6061);
xnor U6884 (N_6884,N_6238,N_6106);
nand U6885 (N_6885,N_6061,N_6381);
nor U6886 (N_6886,N_6297,N_6140);
or U6887 (N_6887,N_6216,N_6341);
xor U6888 (N_6888,N_6415,N_6125);
xnor U6889 (N_6889,N_6112,N_6324);
or U6890 (N_6890,N_6097,N_6384);
or U6891 (N_6891,N_6301,N_6055);
nand U6892 (N_6892,N_6234,N_6210);
and U6893 (N_6893,N_6437,N_6033);
xor U6894 (N_6894,N_6065,N_6358);
and U6895 (N_6895,N_6420,N_6403);
nor U6896 (N_6896,N_6385,N_6413);
and U6897 (N_6897,N_6407,N_6465);
xnor U6898 (N_6898,N_6080,N_6083);
and U6899 (N_6899,N_6414,N_6053);
nand U6900 (N_6900,N_6162,N_6416);
nor U6901 (N_6901,N_6281,N_6431);
and U6902 (N_6902,N_6320,N_6389);
and U6903 (N_6903,N_6007,N_6440);
xor U6904 (N_6904,N_6321,N_6261);
and U6905 (N_6905,N_6210,N_6439);
nand U6906 (N_6906,N_6123,N_6058);
nor U6907 (N_6907,N_6263,N_6411);
and U6908 (N_6908,N_6145,N_6172);
nand U6909 (N_6909,N_6216,N_6032);
nor U6910 (N_6910,N_6287,N_6188);
nand U6911 (N_6911,N_6233,N_6370);
and U6912 (N_6912,N_6405,N_6132);
or U6913 (N_6913,N_6273,N_6159);
nand U6914 (N_6914,N_6131,N_6144);
nor U6915 (N_6915,N_6392,N_6318);
xnor U6916 (N_6916,N_6235,N_6188);
nand U6917 (N_6917,N_6357,N_6376);
or U6918 (N_6918,N_6141,N_6213);
xnor U6919 (N_6919,N_6172,N_6348);
xnor U6920 (N_6920,N_6498,N_6337);
nand U6921 (N_6921,N_6133,N_6309);
nand U6922 (N_6922,N_6019,N_6198);
nor U6923 (N_6923,N_6051,N_6166);
nor U6924 (N_6924,N_6373,N_6075);
and U6925 (N_6925,N_6207,N_6433);
xnor U6926 (N_6926,N_6317,N_6230);
or U6927 (N_6927,N_6102,N_6131);
xnor U6928 (N_6928,N_6252,N_6332);
xor U6929 (N_6929,N_6396,N_6388);
nor U6930 (N_6930,N_6051,N_6340);
nand U6931 (N_6931,N_6145,N_6243);
and U6932 (N_6932,N_6418,N_6478);
xor U6933 (N_6933,N_6400,N_6122);
nor U6934 (N_6934,N_6353,N_6325);
nand U6935 (N_6935,N_6496,N_6227);
nor U6936 (N_6936,N_6315,N_6112);
nor U6937 (N_6937,N_6252,N_6056);
xor U6938 (N_6938,N_6277,N_6116);
and U6939 (N_6939,N_6051,N_6196);
and U6940 (N_6940,N_6085,N_6245);
nor U6941 (N_6941,N_6465,N_6132);
nor U6942 (N_6942,N_6271,N_6224);
xor U6943 (N_6943,N_6437,N_6428);
or U6944 (N_6944,N_6405,N_6279);
or U6945 (N_6945,N_6130,N_6428);
or U6946 (N_6946,N_6169,N_6311);
xor U6947 (N_6947,N_6019,N_6109);
nor U6948 (N_6948,N_6173,N_6360);
nor U6949 (N_6949,N_6427,N_6035);
nand U6950 (N_6950,N_6459,N_6050);
or U6951 (N_6951,N_6301,N_6216);
nor U6952 (N_6952,N_6482,N_6423);
nor U6953 (N_6953,N_6243,N_6395);
xor U6954 (N_6954,N_6251,N_6400);
xnor U6955 (N_6955,N_6130,N_6316);
nand U6956 (N_6956,N_6081,N_6235);
and U6957 (N_6957,N_6483,N_6306);
and U6958 (N_6958,N_6111,N_6461);
and U6959 (N_6959,N_6098,N_6176);
or U6960 (N_6960,N_6101,N_6044);
xor U6961 (N_6961,N_6177,N_6200);
or U6962 (N_6962,N_6447,N_6008);
nor U6963 (N_6963,N_6006,N_6202);
or U6964 (N_6964,N_6428,N_6044);
nand U6965 (N_6965,N_6299,N_6238);
and U6966 (N_6966,N_6097,N_6210);
and U6967 (N_6967,N_6012,N_6335);
nand U6968 (N_6968,N_6271,N_6033);
xnor U6969 (N_6969,N_6082,N_6004);
xor U6970 (N_6970,N_6131,N_6202);
or U6971 (N_6971,N_6383,N_6211);
xor U6972 (N_6972,N_6122,N_6307);
nor U6973 (N_6973,N_6484,N_6178);
nor U6974 (N_6974,N_6388,N_6228);
nor U6975 (N_6975,N_6306,N_6136);
and U6976 (N_6976,N_6218,N_6299);
nand U6977 (N_6977,N_6017,N_6203);
xor U6978 (N_6978,N_6220,N_6378);
nand U6979 (N_6979,N_6421,N_6137);
xnor U6980 (N_6980,N_6329,N_6086);
nand U6981 (N_6981,N_6364,N_6110);
nor U6982 (N_6982,N_6190,N_6035);
nand U6983 (N_6983,N_6315,N_6001);
nor U6984 (N_6984,N_6033,N_6127);
nor U6985 (N_6985,N_6237,N_6438);
xor U6986 (N_6986,N_6096,N_6111);
xor U6987 (N_6987,N_6458,N_6023);
and U6988 (N_6988,N_6419,N_6340);
or U6989 (N_6989,N_6232,N_6247);
and U6990 (N_6990,N_6303,N_6261);
or U6991 (N_6991,N_6211,N_6270);
nor U6992 (N_6992,N_6198,N_6150);
xor U6993 (N_6993,N_6049,N_6331);
xnor U6994 (N_6994,N_6388,N_6296);
nor U6995 (N_6995,N_6320,N_6018);
nor U6996 (N_6996,N_6433,N_6310);
nand U6997 (N_6997,N_6292,N_6282);
or U6998 (N_6998,N_6104,N_6287);
nor U6999 (N_6999,N_6186,N_6222);
or U7000 (N_7000,N_6826,N_6971);
or U7001 (N_7001,N_6721,N_6818);
or U7002 (N_7002,N_6501,N_6705);
nor U7003 (N_7003,N_6875,N_6576);
xnor U7004 (N_7004,N_6665,N_6512);
xnor U7005 (N_7005,N_6733,N_6638);
or U7006 (N_7006,N_6860,N_6792);
and U7007 (N_7007,N_6752,N_6551);
nor U7008 (N_7008,N_6523,N_6850);
and U7009 (N_7009,N_6659,N_6834);
nor U7010 (N_7010,N_6714,N_6653);
and U7011 (N_7011,N_6704,N_6902);
or U7012 (N_7012,N_6662,N_6587);
xnor U7013 (N_7013,N_6696,N_6967);
or U7014 (N_7014,N_6647,N_6825);
nor U7015 (N_7015,N_6539,N_6796);
xnor U7016 (N_7016,N_6553,N_6962);
nand U7017 (N_7017,N_6734,N_6869);
or U7018 (N_7018,N_6595,N_6813);
and U7019 (N_7019,N_6511,N_6642);
and U7020 (N_7020,N_6697,N_6560);
and U7021 (N_7021,N_6926,N_6858);
nor U7022 (N_7022,N_6801,N_6631);
xnor U7023 (N_7023,N_6531,N_6703);
nand U7024 (N_7024,N_6740,N_6984);
and U7025 (N_7025,N_6570,N_6888);
xnor U7026 (N_7026,N_6824,N_6938);
nand U7027 (N_7027,N_6520,N_6775);
and U7028 (N_7028,N_6500,N_6545);
and U7029 (N_7029,N_6528,N_6953);
nand U7030 (N_7030,N_6514,N_6903);
xnor U7031 (N_7031,N_6982,N_6954);
nor U7032 (N_7032,N_6744,N_6836);
or U7033 (N_7033,N_6683,N_6550);
nand U7034 (N_7034,N_6717,N_6678);
nor U7035 (N_7035,N_6767,N_6680);
or U7036 (N_7036,N_6980,N_6592);
nand U7037 (N_7037,N_6513,N_6709);
xnor U7038 (N_7038,N_6863,N_6547);
nor U7039 (N_7039,N_6932,N_6636);
nor U7040 (N_7040,N_6632,N_6772);
nor U7041 (N_7041,N_6666,N_6517);
nor U7042 (N_7042,N_6761,N_6784);
xnor U7043 (N_7043,N_6635,N_6920);
xor U7044 (N_7044,N_6838,N_6710);
xnor U7045 (N_7045,N_6786,N_6798);
and U7046 (N_7046,N_6942,N_6948);
nand U7047 (N_7047,N_6605,N_6625);
xor U7048 (N_7048,N_6506,N_6979);
nand U7049 (N_7049,N_6994,N_6685);
or U7050 (N_7050,N_6541,N_6987);
nor U7051 (N_7051,N_6711,N_6886);
xor U7052 (N_7052,N_6943,N_6731);
nand U7053 (N_7053,N_6606,N_6654);
and U7054 (N_7054,N_6743,N_6961);
nor U7055 (N_7055,N_6530,N_6695);
xnor U7056 (N_7056,N_6811,N_6781);
nor U7057 (N_7057,N_6591,N_6751);
xor U7058 (N_7058,N_6660,N_6882);
and U7059 (N_7059,N_6768,N_6873);
and U7060 (N_7060,N_6968,N_6815);
nor U7061 (N_7061,N_6610,N_6912);
nand U7062 (N_7062,N_6684,N_6600);
or U7063 (N_7063,N_6527,N_6544);
or U7064 (N_7064,N_6599,N_6956);
nor U7065 (N_7065,N_6965,N_6650);
or U7066 (N_7066,N_6681,N_6661);
xor U7067 (N_7067,N_6603,N_6640);
or U7068 (N_7068,N_6742,N_6622);
xor U7069 (N_7069,N_6508,N_6891);
xnor U7070 (N_7070,N_6549,N_6657);
or U7071 (N_7071,N_6791,N_6690);
xnor U7072 (N_7072,N_6713,N_6829);
and U7073 (N_7073,N_6876,N_6516);
nand U7074 (N_7074,N_6578,N_6619);
xor U7075 (N_7075,N_6628,N_6581);
and U7076 (N_7076,N_6773,N_6613);
and U7077 (N_7077,N_6735,N_6522);
nand U7078 (N_7078,N_6941,N_6974);
xnor U7079 (N_7079,N_6676,N_6828);
nand U7080 (N_7080,N_6701,N_6723);
nor U7081 (N_7081,N_6799,N_6669);
xor U7082 (N_7082,N_6831,N_6585);
nand U7083 (N_7083,N_6845,N_6679);
nor U7084 (N_7084,N_6716,N_6552);
and U7085 (N_7085,N_6857,N_6614);
nor U7086 (N_7086,N_6533,N_6901);
or U7087 (N_7087,N_6852,N_6839);
or U7088 (N_7088,N_6866,N_6870);
or U7089 (N_7089,N_6949,N_6986);
xnor U7090 (N_7090,N_6577,N_6687);
xnor U7091 (N_7091,N_6846,N_6893);
or U7092 (N_7092,N_6970,N_6787);
nand U7093 (N_7093,N_6859,N_6726);
and U7094 (N_7094,N_6575,N_6981);
nand U7095 (N_7095,N_6915,N_6564);
nand U7096 (N_7096,N_6612,N_6992);
or U7097 (N_7097,N_6817,N_6651);
or U7098 (N_7098,N_6567,N_6972);
or U7099 (N_7099,N_6918,N_6675);
and U7100 (N_7100,N_6837,N_6874);
or U7101 (N_7101,N_6593,N_6853);
and U7102 (N_7102,N_6722,N_6770);
or U7103 (N_7103,N_6788,N_6579);
nor U7104 (N_7104,N_6790,N_6805);
and U7105 (N_7105,N_6691,N_6963);
xnor U7106 (N_7106,N_6867,N_6955);
nor U7107 (N_7107,N_6518,N_6785);
and U7108 (N_7108,N_6999,N_6643);
xnor U7109 (N_7109,N_6978,N_6618);
nand U7110 (N_7110,N_6559,N_6995);
xor U7111 (N_7111,N_6904,N_6928);
and U7112 (N_7112,N_6615,N_6849);
xnor U7113 (N_7113,N_6624,N_6923);
xnor U7114 (N_7114,N_6935,N_6626);
xnor U7115 (N_7115,N_6589,N_6692);
and U7116 (N_7116,N_6686,N_6765);
nor U7117 (N_7117,N_6543,N_6755);
nor U7118 (N_7118,N_6725,N_6871);
nor U7119 (N_7119,N_6515,N_6535);
and U7120 (N_7120,N_6645,N_6607);
and U7121 (N_7121,N_6909,N_6804);
xor U7122 (N_7122,N_6532,N_6538);
or U7123 (N_7123,N_6769,N_6969);
and U7124 (N_7124,N_6582,N_6729);
nand U7125 (N_7125,N_6759,N_6964);
and U7126 (N_7126,N_6843,N_6947);
xor U7127 (N_7127,N_6656,N_6644);
nor U7128 (N_7128,N_6749,N_6802);
and U7129 (N_7129,N_6602,N_6673);
nor U7130 (N_7130,N_6960,N_6993);
nand U7131 (N_7131,N_6563,N_6988);
or U7132 (N_7132,N_6504,N_6883);
and U7133 (N_7133,N_6919,N_6778);
nor U7134 (N_7134,N_6633,N_6668);
nand U7135 (N_7135,N_6914,N_6983);
xnor U7136 (N_7136,N_6823,N_6720);
xnor U7137 (N_7137,N_6921,N_6727);
or U7138 (N_7138,N_6944,N_6868);
or U7139 (N_7139,N_6899,N_6597);
and U7140 (N_7140,N_6763,N_6525);
or U7141 (N_7141,N_6865,N_6872);
nand U7142 (N_7142,N_6534,N_6739);
nand U7143 (N_7143,N_6639,N_6689);
and U7144 (N_7144,N_6677,N_6502);
nor U7145 (N_7145,N_6808,N_6841);
and U7146 (N_7146,N_6930,N_6598);
or U7147 (N_7147,N_6848,N_6833);
nor U7148 (N_7148,N_6996,N_6807);
nand U7149 (N_7149,N_6707,N_6616);
xor U7150 (N_7150,N_6572,N_6601);
nor U7151 (N_7151,N_6670,N_6569);
nor U7152 (N_7152,N_6950,N_6712);
nor U7153 (N_7153,N_6546,N_6561);
nor U7154 (N_7154,N_6574,N_6596);
and U7155 (N_7155,N_6728,N_6881);
or U7156 (N_7156,N_6795,N_6861);
nor U7157 (N_7157,N_6896,N_6758);
xnor U7158 (N_7158,N_6966,N_6537);
and U7159 (N_7159,N_6764,N_6708);
and U7160 (N_7160,N_6766,N_6706);
nand U7161 (N_7161,N_6900,N_6776);
nor U7162 (N_7162,N_6975,N_6946);
and U7163 (N_7163,N_6905,N_6976);
and U7164 (N_7164,N_6732,N_6736);
and U7165 (N_7165,N_6910,N_6936);
and U7166 (N_7166,N_6663,N_6864);
or U7167 (N_7167,N_6648,N_6630);
and U7168 (N_7168,N_6789,N_6604);
xnor U7169 (N_7169,N_6977,N_6998);
xor U7170 (N_7170,N_6620,N_6895);
xnor U7171 (N_7171,N_6794,N_6973);
nand U7172 (N_7172,N_6519,N_6526);
xor U7173 (N_7173,N_6753,N_6568);
or U7174 (N_7174,N_6617,N_6990);
nor U7175 (N_7175,N_6884,N_6851);
nand U7176 (N_7176,N_6608,N_6760);
or U7177 (N_7177,N_6814,N_6637);
nand U7178 (N_7178,N_6952,N_6951);
and U7179 (N_7179,N_6844,N_6566);
and U7180 (N_7180,N_6822,N_6590);
or U7181 (N_7181,N_6957,N_6584);
or U7182 (N_7182,N_6842,N_6509);
nor U7183 (N_7183,N_6611,N_6929);
or U7184 (N_7184,N_6819,N_6827);
xor U7185 (N_7185,N_6594,N_6922);
nor U7186 (N_7186,N_6702,N_6820);
xnor U7187 (N_7187,N_6885,N_6521);
nand U7188 (N_7188,N_6649,N_6989);
nor U7189 (N_7189,N_6991,N_6854);
xnor U7190 (N_7190,N_6718,N_6583);
nand U7191 (N_7191,N_6627,N_6586);
xnor U7192 (N_7192,N_6750,N_6667);
and U7193 (N_7193,N_6658,N_6931);
nand U7194 (N_7194,N_6693,N_6985);
xor U7195 (N_7195,N_6933,N_6894);
or U7196 (N_7196,N_6803,N_6892);
nor U7197 (N_7197,N_6925,N_6745);
nor U7198 (N_7198,N_6821,N_6571);
xnor U7199 (N_7199,N_6746,N_6507);
nand U7200 (N_7200,N_6937,N_6629);
nand U7201 (N_7201,N_6641,N_6906);
nor U7202 (N_7202,N_6877,N_6783);
nor U7203 (N_7203,N_6800,N_6505);
xnor U7204 (N_7204,N_6682,N_6847);
nor U7205 (N_7205,N_6655,N_6540);
xnor U7206 (N_7206,N_6939,N_6565);
nand U7207 (N_7207,N_6555,N_6699);
xnor U7208 (N_7208,N_6588,N_6878);
xnor U7209 (N_7209,N_6810,N_6958);
or U7210 (N_7210,N_6510,N_6782);
nand U7211 (N_7211,N_6672,N_6634);
or U7212 (N_7212,N_6835,N_6940);
nand U7213 (N_7213,N_6548,N_6806);
nor U7214 (N_7214,N_6694,N_6879);
nor U7215 (N_7215,N_6907,N_6777);
nand U7216 (N_7216,N_6913,N_6945);
xor U7217 (N_7217,N_6959,N_6908);
or U7218 (N_7218,N_6927,N_6719);
or U7219 (N_7219,N_6609,N_6880);
or U7220 (N_7220,N_6780,N_6862);
nand U7221 (N_7221,N_6897,N_6674);
xnor U7222 (N_7222,N_6779,N_6747);
nand U7223 (N_7223,N_6797,N_6646);
or U7224 (N_7224,N_6887,N_6856);
nor U7225 (N_7225,N_6754,N_6832);
nand U7226 (N_7226,N_6700,N_6557);
xnor U7227 (N_7227,N_6889,N_6997);
nand U7228 (N_7228,N_6724,N_6580);
nor U7229 (N_7229,N_6890,N_6793);
or U7230 (N_7230,N_6688,N_6558);
nor U7231 (N_7231,N_6698,N_6830);
or U7232 (N_7232,N_6529,N_6737);
nor U7233 (N_7233,N_6573,N_6542);
or U7234 (N_7234,N_6812,N_6738);
nand U7235 (N_7235,N_6730,N_6809);
nand U7236 (N_7236,N_6756,N_6934);
nor U7237 (N_7237,N_6623,N_6774);
or U7238 (N_7238,N_6762,N_6911);
and U7239 (N_7239,N_6556,N_6652);
or U7240 (N_7240,N_6757,N_6916);
nand U7241 (N_7241,N_6536,N_6748);
nor U7242 (N_7242,N_6917,N_6741);
or U7243 (N_7243,N_6554,N_6562);
xor U7244 (N_7244,N_6671,N_6816);
and U7245 (N_7245,N_6771,N_6855);
and U7246 (N_7246,N_6924,N_6503);
nor U7247 (N_7247,N_6621,N_6715);
nand U7248 (N_7248,N_6840,N_6664);
nand U7249 (N_7249,N_6524,N_6898);
or U7250 (N_7250,N_6853,N_6705);
nor U7251 (N_7251,N_6863,N_6638);
xnor U7252 (N_7252,N_6525,N_6734);
or U7253 (N_7253,N_6785,N_6874);
xor U7254 (N_7254,N_6557,N_6915);
xor U7255 (N_7255,N_6510,N_6754);
nor U7256 (N_7256,N_6995,N_6708);
and U7257 (N_7257,N_6794,N_6987);
nor U7258 (N_7258,N_6754,N_6585);
and U7259 (N_7259,N_6825,N_6828);
nor U7260 (N_7260,N_6813,N_6516);
or U7261 (N_7261,N_6882,N_6953);
or U7262 (N_7262,N_6761,N_6866);
and U7263 (N_7263,N_6914,N_6902);
nor U7264 (N_7264,N_6620,N_6592);
nor U7265 (N_7265,N_6709,N_6827);
nor U7266 (N_7266,N_6509,N_6753);
xnor U7267 (N_7267,N_6840,N_6541);
nand U7268 (N_7268,N_6511,N_6755);
nand U7269 (N_7269,N_6689,N_6611);
and U7270 (N_7270,N_6725,N_6642);
and U7271 (N_7271,N_6866,N_6503);
nand U7272 (N_7272,N_6771,N_6763);
or U7273 (N_7273,N_6598,N_6548);
xor U7274 (N_7274,N_6633,N_6588);
xor U7275 (N_7275,N_6521,N_6666);
nor U7276 (N_7276,N_6745,N_6764);
or U7277 (N_7277,N_6838,N_6917);
nand U7278 (N_7278,N_6571,N_6693);
nand U7279 (N_7279,N_6849,N_6783);
and U7280 (N_7280,N_6931,N_6983);
nand U7281 (N_7281,N_6523,N_6792);
xor U7282 (N_7282,N_6519,N_6755);
xor U7283 (N_7283,N_6526,N_6762);
nand U7284 (N_7284,N_6584,N_6790);
or U7285 (N_7285,N_6836,N_6596);
nor U7286 (N_7286,N_6552,N_6651);
nand U7287 (N_7287,N_6945,N_6806);
and U7288 (N_7288,N_6603,N_6692);
or U7289 (N_7289,N_6875,N_6699);
or U7290 (N_7290,N_6783,N_6992);
nor U7291 (N_7291,N_6982,N_6909);
and U7292 (N_7292,N_6604,N_6630);
nor U7293 (N_7293,N_6841,N_6674);
xnor U7294 (N_7294,N_6795,N_6516);
xnor U7295 (N_7295,N_6501,N_6533);
nor U7296 (N_7296,N_6652,N_6664);
and U7297 (N_7297,N_6788,N_6754);
nor U7298 (N_7298,N_6753,N_6561);
xnor U7299 (N_7299,N_6738,N_6839);
and U7300 (N_7300,N_6516,N_6978);
and U7301 (N_7301,N_6765,N_6952);
xnor U7302 (N_7302,N_6542,N_6980);
xor U7303 (N_7303,N_6775,N_6535);
nand U7304 (N_7304,N_6885,N_6692);
xnor U7305 (N_7305,N_6839,N_6717);
or U7306 (N_7306,N_6981,N_6855);
and U7307 (N_7307,N_6930,N_6500);
and U7308 (N_7308,N_6985,N_6960);
xor U7309 (N_7309,N_6609,N_6548);
nand U7310 (N_7310,N_6915,N_6599);
or U7311 (N_7311,N_6760,N_6952);
or U7312 (N_7312,N_6541,N_6878);
or U7313 (N_7313,N_6893,N_6632);
nand U7314 (N_7314,N_6648,N_6710);
nand U7315 (N_7315,N_6859,N_6655);
nor U7316 (N_7316,N_6639,N_6910);
and U7317 (N_7317,N_6952,N_6977);
and U7318 (N_7318,N_6745,N_6801);
or U7319 (N_7319,N_6668,N_6750);
nand U7320 (N_7320,N_6708,N_6609);
and U7321 (N_7321,N_6537,N_6521);
xor U7322 (N_7322,N_6978,N_6576);
nor U7323 (N_7323,N_6616,N_6855);
nand U7324 (N_7324,N_6679,N_6574);
nand U7325 (N_7325,N_6854,N_6627);
nand U7326 (N_7326,N_6633,N_6650);
and U7327 (N_7327,N_6603,N_6531);
nand U7328 (N_7328,N_6770,N_6708);
nand U7329 (N_7329,N_6640,N_6751);
and U7330 (N_7330,N_6936,N_6626);
xor U7331 (N_7331,N_6540,N_6944);
xor U7332 (N_7332,N_6915,N_6595);
nor U7333 (N_7333,N_6719,N_6867);
nor U7334 (N_7334,N_6591,N_6894);
and U7335 (N_7335,N_6502,N_6876);
nand U7336 (N_7336,N_6971,N_6816);
xnor U7337 (N_7337,N_6743,N_6510);
or U7338 (N_7338,N_6986,N_6583);
nor U7339 (N_7339,N_6795,N_6742);
nor U7340 (N_7340,N_6738,N_6907);
xnor U7341 (N_7341,N_6852,N_6563);
or U7342 (N_7342,N_6801,N_6800);
nand U7343 (N_7343,N_6945,N_6524);
or U7344 (N_7344,N_6699,N_6916);
or U7345 (N_7345,N_6503,N_6645);
or U7346 (N_7346,N_6691,N_6720);
and U7347 (N_7347,N_6938,N_6751);
nand U7348 (N_7348,N_6527,N_6967);
and U7349 (N_7349,N_6706,N_6700);
and U7350 (N_7350,N_6512,N_6893);
nor U7351 (N_7351,N_6782,N_6872);
nor U7352 (N_7352,N_6683,N_6626);
nor U7353 (N_7353,N_6784,N_6889);
nand U7354 (N_7354,N_6937,N_6990);
and U7355 (N_7355,N_6956,N_6778);
nor U7356 (N_7356,N_6813,N_6893);
and U7357 (N_7357,N_6825,N_6706);
xnor U7358 (N_7358,N_6751,N_6771);
and U7359 (N_7359,N_6621,N_6675);
nor U7360 (N_7360,N_6551,N_6915);
nor U7361 (N_7361,N_6730,N_6878);
or U7362 (N_7362,N_6605,N_6943);
xnor U7363 (N_7363,N_6792,N_6929);
or U7364 (N_7364,N_6629,N_6570);
nor U7365 (N_7365,N_6871,N_6988);
and U7366 (N_7366,N_6524,N_6664);
or U7367 (N_7367,N_6572,N_6851);
nor U7368 (N_7368,N_6689,N_6959);
or U7369 (N_7369,N_6948,N_6888);
nor U7370 (N_7370,N_6584,N_6742);
xnor U7371 (N_7371,N_6886,N_6960);
nand U7372 (N_7372,N_6842,N_6864);
nand U7373 (N_7373,N_6667,N_6763);
and U7374 (N_7374,N_6737,N_6890);
nand U7375 (N_7375,N_6871,N_6524);
nand U7376 (N_7376,N_6794,N_6863);
nand U7377 (N_7377,N_6729,N_6584);
and U7378 (N_7378,N_6752,N_6738);
xor U7379 (N_7379,N_6858,N_6919);
nor U7380 (N_7380,N_6986,N_6513);
nand U7381 (N_7381,N_6711,N_6682);
nand U7382 (N_7382,N_6809,N_6734);
or U7383 (N_7383,N_6654,N_6599);
and U7384 (N_7384,N_6807,N_6582);
xor U7385 (N_7385,N_6975,N_6668);
nor U7386 (N_7386,N_6709,N_6511);
and U7387 (N_7387,N_6755,N_6571);
nor U7388 (N_7388,N_6578,N_6514);
or U7389 (N_7389,N_6673,N_6613);
xnor U7390 (N_7390,N_6898,N_6865);
or U7391 (N_7391,N_6728,N_6913);
and U7392 (N_7392,N_6847,N_6524);
nand U7393 (N_7393,N_6533,N_6580);
nand U7394 (N_7394,N_6809,N_6625);
or U7395 (N_7395,N_6656,N_6990);
nand U7396 (N_7396,N_6992,N_6848);
or U7397 (N_7397,N_6777,N_6667);
or U7398 (N_7398,N_6740,N_6727);
or U7399 (N_7399,N_6594,N_6909);
xnor U7400 (N_7400,N_6709,N_6748);
or U7401 (N_7401,N_6650,N_6913);
nand U7402 (N_7402,N_6887,N_6574);
and U7403 (N_7403,N_6987,N_6959);
and U7404 (N_7404,N_6848,N_6595);
xnor U7405 (N_7405,N_6911,N_6993);
and U7406 (N_7406,N_6576,N_6868);
nor U7407 (N_7407,N_6503,N_6884);
nand U7408 (N_7408,N_6563,N_6771);
nand U7409 (N_7409,N_6800,N_6779);
xnor U7410 (N_7410,N_6754,N_6628);
xnor U7411 (N_7411,N_6527,N_6911);
and U7412 (N_7412,N_6693,N_6668);
nand U7413 (N_7413,N_6562,N_6948);
or U7414 (N_7414,N_6745,N_6859);
nand U7415 (N_7415,N_6637,N_6878);
or U7416 (N_7416,N_6605,N_6717);
xor U7417 (N_7417,N_6580,N_6942);
nand U7418 (N_7418,N_6622,N_6512);
and U7419 (N_7419,N_6903,N_6599);
nand U7420 (N_7420,N_6766,N_6741);
nand U7421 (N_7421,N_6710,N_6593);
and U7422 (N_7422,N_6702,N_6650);
and U7423 (N_7423,N_6746,N_6546);
or U7424 (N_7424,N_6851,N_6780);
xnor U7425 (N_7425,N_6801,N_6752);
nor U7426 (N_7426,N_6895,N_6585);
nor U7427 (N_7427,N_6874,N_6525);
xor U7428 (N_7428,N_6808,N_6777);
nand U7429 (N_7429,N_6552,N_6942);
xor U7430 (N_7430,N_6915,N_6618);
xor U7431 (N_7431,N_6540,N_6608);
nor U7432 (N_7432,N_6542,N_6650);
and U7433 (N_7433,N_6676,N_6786);
nor U7434 (N_7434,N_6599,N_6827);
nand U7435 (N_7435,N_6656,N_6864);
or U7436 (N_7436,N_6698,N_6712);
nand U7437 (N_7437,N_6539,N_6705);
nand U7438 (N_7438,N_6987,N_6801);
or U7439 (N_7439,N_6850,N_6680);
nand U7440 (N_7440,N_6571,N_6777);
nand U7441 (N_7441,N_6784,N_6688);
xnor U7442 (N_7442,N_6775,N_6969);
nand U7443 (N_7443,N_6543,N_6620);
nor U7444 (N_7444,N_6834,N_6906);
xnor U7445 (N_7445,N_6682,N_6569);
and U7446 (N_7446,N_6854,N_6712);
or U7447 (N_7447,N_6531,N_6587);
or U7448 (N_7448,N_6825,N_6905);
or U7449 (N_7449,N_6756,N_6603);
and U7450 (N_7450,N_6871,N_6615);
xor U7451 (N_7451,N_6940,N_6929);
nand U7452 (N_7452,N_6594,N_6507);
and U7453 (N_7453,N_6878,N_6610);
nand U7454 (N_7454,N_6743,N_6643);
xnor U7455 (N_7455,N_6990,N_6991);
nor U7456 (N_7456,N_6908,N_6730);
xor U7457 (N_7457,N_6721,N_6628);
nor U7458 (N_7458,N_6570,N_6514);
or U7459 (N_7459,N_6936,N_6787);
and U7460 (N_7460,N_6581,N_6545);
nand U7461 (N_7461,N_6518,N_6558);
xor U7462 (N_7462,N_6674,N_6584);
nand U7463 (N_7463,N_6608,N_6750);
and U7464 (N_7464,N_6853,N_6632);
or U7465 (N_7465,N_6672,N_6561);
and U7466 (N_7466,N_6746,N_6942);
nor U7467 (N_7467,N_6608,N_6552);
and U7468 (N_7468,N_6866,N_6782);
xnor U7469 (N_7469,N_6863,N_6821);
xor U7470 (N_7470,N_6683,N_6846);
and U7471 (N_7471,N_6629,N_6950);
nor U7472 (N_7472,N_6813,N_6536);
and U7473 (N_7473,N_6821,N_6990);
nand U7474 (N_7474,N_6762,N_6676);
nand U7475 (N_7475,N_6818,N_6581);
and U7476 (N_7476,N_6547,N_6730);
nor U7477 (N_7477,N_6635,N_6637);
or U7478 (N_7478,N_6793,N_6700);
or U7479 (N_7479,N_6502,N_6946);
nor U7480 (N_7480,N_6691,N_6611);
nand U7481 (N_7481,N_6654,N_6825);
nor U7482 (N_7482,N_6831,N_6659);
nand U7483 (N_7483,N_6876,N_6869);
xor U7484 (N_7484,N_6506,N_6866);
xor U7485 (N_7485,N_6781,N_6608);
xnor U7486 (N_7486,N_6532,N_6519);
nor U7487 (N_7487,N_6778,N_6782);
nand U7488 (N_7488,N_6751,N_6851);
nand U7489 (N_7489,N_6829,N_6551);
nand U7490 (N_7490,N_6517,N_6779);
nor U7491 (N_7491,N_6922,N_6718);
nand U7492 (N_7492,N_6754,N_6867);
nand U7493 (N_7493,N_6940,N_6936);
nand U7494 (N_7494,N_6520,N_6579);
nand U7495 (N_7495,N_6843,N_6937);
and U7496 (N_7496,N_6708,N_6988);
or U7497 (N_7497,N_6796,N_6574);
and U7498 (N_7498,N_6968,N_6912);
nand U7499 (N_7499,N_6764,N_6853);
xnor U7500 (N_7500,N_7097,N_7420);
nand U7501 (N_7501,N_7474,N_7424);
nor U7502 (N_7502,N_7089,N_7461);
nor U7503 (N_7503,N_7046,N_7333);
xnor U7504 (N_7504,N_7217,N_7106);
or U7505 (N_7505,N_7235,N_7225);
or U7506 (N_7506,N_7329,N_7100);
and U7507 (N_7507,N_7445,N_7468);
and U7508 (N_7508,N_7363,N_7198);
xor U7509 (N_7509,N_7218,N_7421);
nor U7510 (N_7510,N_7381,N_7079);
nor U7511 (N_7511,N_7268,N_7232);
nand U7512 (N_7512,N_7016,N_7024);
and U7513 (N_7513,N_7012,N_7127);
nor U7514 (N_7514,N_7011,N_7414);
xnor U7515 (N_7515,N_7365,N_7297);
xnor U7516 (N_7516,N_7241,N_7350);
or U7517 (N_7517,N_7063,N_7141);
nor U7518 (N_7518,N_7035,N_7344);
and U7519 (N_7519,N_7007,N_7384);
or U7520 (N_7520,N_7243,N_7376);
nor U7521 (N_7521,N_7234,N_7316);
and U7522 (N_7522,N_7188,N_7299);
and U7523 (N_7523,N_7306,N_7361);
nand U7524 (N_7524,N_7454,N_7162);
nor U7525 (N_7525,N_7419,N_7111);
nor U7526 (N_7526,N_7457,N_7207);
and U7527 (N_7527,N_7489,N_7137);
and U7528 (N_7528,N_7266,N_7170);
nand U7529 (N_7529,N_7041,N_7481);
or U7530 (N_7530,N_7403,N_7044);
xor U7531 (N_7531,N_7184,N_7324);
nand U7532 (N_7532,N_7005,N_7321);
or U7533 (N_7533,N_7471,N_7173);
and U7534 (N_7534,N_7150,N_7402);
xnor U7535 (N_7535,N_7259,N_7408);
nor U7536 (N_7536,N_7183,N_7497);
nor U7537 (N_7537,N_7032,N_7288);
xor U7538 (N_7538,N_7023,N_7199);
and U7539 (N_7539,N_7309,N_7144);
nand U7540 (N_7540,N_7192,N_7233);
nand U7541 (N_7541,N_7135,N_7278);
xnor U7542 (N_7542,N_7284,N_7227);
or U7543 (N_7543,N_7015,N_7081);
nand U7544 (N_7544,N_7283,N_7053);
and U7545 (N_7545,N_7047,N_7318);
nor U7546 (N_7546,N_7054,N_7033);
nor U7547 (N_7547,N_7138,N_7108);
nor U7548 (N_7548,N_7061,N_7436);
or U7549 (N_7549,N_7102,N_7274);
and U7550 (N_7550,N_7343,N_7431);
or U7551 (N_7551,N_7031,N_7267);
or U7552 (N_7552,N_7496,N_7475);
and U7553 (N_7553,N_7362,N_7096);
and U7554 (N_7554,N_7349,N_7050);
nor U7555 (N_7555,N_7179,N_7224);
nor U7556 (N_7556,N_7252,N_7312);
xnor U7557 (N_7557,N_7494,N_7051);
or U7558 (N_7558,N_7104,N_7302);
xnor U7559 (N_7559,N_7466,N_7294);
nor U7560 (N_7560,N_7404,N_7129);
or U7561 (N_7561,N_7480,N_7270);
xnor U7562 (N_7562,N_7107,N_7231);
or U7563 (N_7563,N_7222,N_7401);
nand U7564 (N_7564,N_7341,N_7038);
nor U7565 (N_7565,N_7352,N_7470);
nor U7566 (N_7566,N_7388,N_7413);
nand U7567 (N_7567,N_7258,N_7136);
xnor U7568 (N_7568,N_7269,N_7029);
or U7569 (N_7569,N_7479,N_7206);
or U7570 (N_7570,N_7189,N_7290);
or U7571 (N_7571,N_7262,N_7340);
or U7572 (N_7572,N_7392,N_7186);
and U7573 (N_7573,N_7026,N_7337);
nand U7574 (N_7574,N_7415,N_7453);
or U7575 (N_7575,N_7490,N_7220);
xor U7576 (N_7576,N_7301,N_7171);
nand U7577 (N_7577,N_7034,N_7372);
or U7578 (N_7578,N_7084,N_7209);
nand U7579 (N_7579,N_7037,N_7158);
nor U7580 (N_7580,N_7025,N_7257);
xnor U7581 (N_7581,N_7467,N_7131);
xor U7582 (N_7582,N_7169,N_7182);
xnor U7583 (N_7583,N_7152,N_7397);
and U7584 (N_7584,N_7027,N_7293);
xnor U7585 (N_7585,N_7326,N_7200);
or U7586 (N_7586,N_7380,N_7210);
and U7587 (N_7587,N_7400,N_7078);
and U7588 (N_7588,N_7006,N_7282);
or U7589 (N_7589,N_7382,N_7425);
and U7590 (N_7590,N_7263,N_7331);
or U7591 (N_7591,N_7391,N_7409);
nand U7592 (N_7592,N_7036,N_7369);
nand U7593 (N_7593,N_7004,N_7354);
nor U7594 (N_7594,N_7459,N_7020);
nor U7595 (N_7595,N_7332,N_7458);
nor U7596 (N_7596,N_7101,N_7310);
nand U7597 (N_7597,N_7307,N_7132);
nor U7598 (N_7598,N_7239,N_7143);
or U7599 (N_7599,N_7389,N_7378);
xor U7600 (N_7600,N_7160,N_7010);
nor U7601 (N_7601,N_7456,N_7056);
or U7602 (N_7602,N_7219,N_7336);
xor U7603 (N_7603,N_7465,N_7422);
xor U7604 (N_7604,N_7040,N_7066);
nor U7605 (N_7605,N_7493,N_7203);
and U7606 (N_7606,N_7237,N_7303);
nor U7607 (N_7607,N_7157,N_7075);
and U7608 (N_7608,N_7115,N_7483);
and U7609 (N_7609,N_7077,N_7142);
nor U7610 (N_7610,N_7279,N_7292);
xor U7611 (N_7611,N_7229,N_7165);
nor U7612 (N_7612,N_7426,N_7215);
xor U7613 (N_7613,N_7298,N_7126);
or U7614 (N_7614,N_7407,N_7285);
nand U7615 (N_7615,N_7476,N_7342);
and U7616 (N_7616,N_7065,N_7484);
nand U7617 (N_7617,N_7289,N_7181);
nand U7618 (N_7618,N_7260,N_7472);
nand U7619 (N_7619,N_7069,N_7118);
nand U7620 (N_7620,N_7121,N_7488);
and U7621 (N_7621,N_7264,N_7449);
nor U7622 (N_7622,N_7139,N_7327);
nand U7623 (N_7623,N_7338,N_7021);
nor U7624 (N_7624,N_7256,N_7335);
or U7625 (N_7625,N_7120,N_7228);
or U7626 (N_7626,N_7370,N_7473);
and U7627 (N_7627,N_7296,N_7076);
and U7628 (N_7628,N_7112,N_7379);
and U7629 (N_7629,N_7175,N_7067);
xor U7630 (N_7630,N_7367,N_7482);
nor U7631 (N_7631,N_7442,N_7113);
xnor U7632 (N_7632,N_7048,N_7399);
nor U7633 (N_7633,N_7491,N_7154);
nor U7634 (N_7634,N_7248,N_7276);
and U7635 (N_7635,N_7022,N_7002);
xor U7636 (N_7636,N_7052,N_7122);
nand U7637 (N_7637,N_7433,N_7230);
nor U7638 (N_7638,N_7202,N_7371);
nor U7639 (N_7639,N_7452,N_7167);
and U7640 (N_7640,N_7000,N_7242);
or U7641 (N_7641,N_7213,N_7130);
xor U7642 (N_7642,N_7319,N_7085);
or U7643 (N_7643,N_7398,N_7134);
and U7644 (N_7644,N_7357,N_7273);
and U7645 (N_7645,N_7383,N_7441);
nand U7646 (N_7646,N_7114,N_7455);
and U7647 (N_7647,N_7148,N_7345);
or U7648 (N_7648,N_7416,N_7091);
and U7649 (N_7649,N_7092,N_7166);
or U7650 (N_7650,N_7325,N_7396);
xnor U7651 (N_7651,N_7185,N_7255);
xnor U7652 (N_7652,N_7393,N_7071);
and U7653 (N_7653,N_7486,N_7430);
xor U7654 (N_7654,N_7295,N_7174);
nand U7655 (N_7655,N_7261,N_7105);
or U7656 (N_7656,N_7275,N_7238);
nor U7657 (N_7657,N_7440,N_7447);
and U7658 (N_7658,N_7394,N_7250);
and U7659 (N_7659,N_7159,N_7265);
and U7660 (N_7660,N_7145,N_7322);
and U7661 (N_7661,N_7197,N_7323);
and U7662 (N_7662,N_7348,N_7423);
nor U7663 (N_7663,N_7030,N_7249);
nor U7664 (N_7664,N_7001,N_7055);
nand U7665 (N_7665,N_7088,N_7064);
or U7666 (N_7666,N_7281,N_7246);
nand U7667 (N_7667,N_7049,N_7245);
or U7668 (N_7668,N_7446,N_7003);
and U7669 (N_7669,N_7103,N_7417);
nor U7670 (N_7670,N_7314,N_7221);
nor U7671 (N_7671,N_7043,N_7271);
and U7672 (N_7672,N_7018,N_7353);
or U7673 (N_7673,N_7028,N_7039);
nand U7674 (N_7674,N_7057,N_7315);
nor U7675 (N_7675,N_7254,N_7180);
and U7676 (N_7676,N_7240,N_7499);
and U7677 (N_7677,N_7305,N_7435);
nand U7678 (N_7678,N_7072,N_7082);
and U7679 (N_7679,N_7042,N_7487);
nand U7680 (N_7680,N_7008,N_7177);
nor U7681 (N_7681,N_7161,N_7410);
nor U7682 (N_7682,N_7311,N_7469);
nand U7683 (N_7683,N_7412,N_7187);
nor U7684 (N_7684,N_7247,N_7133);
and U7685 (N_7685,N_7201,N_7313);
nand U7686 (N_7686,N_7385,N_7366);
or U7687 (N_7687,N_7244,N_7405);
nor U7688 (N_7688,N_7411,N_7060);
xnor U7689 (N_7689,N_7094,N_7444);
and U7690 (N_7690,N_7176,N_7156);
nand U7691 (N_7691,N_7045,N_7390);
and U7692 (N_7692,N_7432,N_7375);
or U7693 (N_7693,N_7147,N_7339);
or U7694 (N_7694,N_7070,N_7226);
nor U7695 (N_7695,N_7355,N_7287);
xor U7696 (N_7696,N_7168,N_7073);
and U7697 (N_7697,N_7485,N_7429);
and U7698 (N_7698,N_7330,N_7058);
and U7699 (N_7699,N_7163,N_7317);
nor U7700 (N_7700,N_7328,N_7277);
and U7701 (N_7701,N_7110,N_7208);
and U7702 (N_7702,N_7172,N_7448);
nor U7703 (N_7703,N_7216,N_7194);
or U7704 (N_7704,N_7346,N_7211);
and U7705 (N_7705,N_7193,N_7368);
and U7706 (N_7706,N_7223,N_7438);
nand U7707 (N_7707,N_7212,N_7300);
or U7708 (N_7708,N_7427,N_7359);
nand U7709 (N_7709,N_7109,N_7117);
nor U7710 (N_7710,N_7356,N_7308);
nor U7711 (N_7711,N_7498,N_7347);
or U7712 (N_7712,N_7095,N_7286);
nand U7713 (N_7713,N_7334,N_7406);
nand U7714 (N_7714,N_7386,N_7164);
nand U7715 (N_7715,N_7123,N_7495);
or U7716 (N_7716,N_7304,N_7291);
nand U7717 (N_7717,N_7450,N_7253);
nand U7718 (N_7718,N_7418,N_7387);
xnor U7719 (N_7719,N_7477,N_7351);
nor U7720 (N_7720,N_7214,N_7395);
nor U7721 (N_7721,N_7492,N_7451);
and U7722 (N_7722,N_7320,N_7178);
nor U7723 (N_7723,N_7140,N_7153);
and U7724 (N_7724,N_7478,N_7464);
nand U7725 (N_7725,N_7195,N_7093);
nor U7726 (N_7726,N_7125,N_7128);
or U7727 (N_7727,N_7374,N_7205);
nor U7728 (N_7728,N_7191,N_7009);
or U7729 (N_7729,N_7062,N_7149);
nor U7730 (N_7730,N_7116,N_7014);
xnor U7731 (N_7731,N_7155,N_7090);
nor U7732 (N_7732,N_7099,N_7080);
xor U7733 (N_7733,N_7434,N_7068);
nand U7734 (N_7734,N_7462,N_7013);
nand U7735 (N_7735,N_7017,N_7272);
nand U7736 (N_7736,N_7019,N_7196);
and U7737 (N_7737,N_7059,N_7074);
xnor U7738 (N_7738,N_7460,N_7204);
nor U7739 (N_7739,N_7358,N_7437);
nor U7740 (N_7740,N_7443,N_7280);
or U7741 (N_7741,N_7428,N_7463);
xnor U7742 (N_7742,N_7377,N_7151);
nor U7743 (N_7743,N_7373,N_7098);
nand U7744 (N_7744,N_7119,N_7086);
and U7745 (N_7745,N_7364,N_7083);
nor U7746 (N_7746,N_7236,N_7087);
and U7747 (N_7747,N_7439,N_7190);
or U7748 (N_7748,N_7251,N_7146);
and U7749 (N_7749,N_7124,N_7360);
nor U7750 (N_7750,N_7031,N_7487);
and U7751 (N_7751,N_7165,N_7357);
or U7752 (N_7752,N_7185,N_7008);
xor U7753 (N_7753,N_7254,N_7080);
and U7754 (N_7754,N_7196,N_7366);
or U7755 (N_7755,N_7229,N_7375);
and U7756 (N_7756,N_7464,N_7399);
xnor U7757 (N_7757,N_7293,N_7133);
or U7758 (N_7758,N_7131,N_7282);
or U7759 (N_7759,N_7408,N_7282);
nand U7760 (N_7760,N_7056,N_7213);
or U7761 (N_7761,N_7170,N_7314);
or U7762 (N_7762,N_7015,N_7193);
and U7763 (N_7763,N_7218,N_7209);
and U7764 (N_7764,N_7459,N_7371);
nand U7765 (N_7765,N_7294,N_7490);
nand U7766 (N_7766,N_7243,N_7227);
or U7767 (N_7767,N_7494,N_7358);
and U7768 (N_7768,N_7485,N_7065);
xor U7769 (N_7769,N_7271,N_7470);
nand U7770 (N_7770,N_7470,N_7267);
nand U7771 (N_7771,N_7290,N_7066);
xor U7772 (N_7772,N_7029,N_7307);
or U7773 (N_7773,N_7436,N_7060);
and U7774 (N_7774,N_7439,N_7265);
xor U7775 (N_7775,N_7424,N_7202);
nor U7776 (N_7776,N_7476,N_7132);
nor U7777 (N_7777,N_7320,N_7405);
xnor U7778 (N_7778,N_7464,N_7113);
nor U7779 (N_7779,N_7186,N_7288);
nand U7780 (N_7780,N_7036,N_7465);
nor U7781 (N_7781,N_7451,N_7057);
or U7782 (N_7782,N_7087,N_7223);
or U7783 (N_7783,N_7325,N_7094);
nand U7784 (N_7784,N_7413,N_7468);
nor U7785 (N_7785,N_7481,N_7426);
xnor U7786 (N_7786,N_7040,N_7031);
nand U7787 (N_7787,N_7283,N_7284);
and U7788 (N_7788,N_7263,N_7267);
xor U7789 (N_7789,N_7201,N_7191);
nand U7790 (N_7790,N_7446,N_7030);
xor U7791 (N_7791,N_7266,N_7186);
xor U7792 (N_7792,N_7086,N_7184);
or U7793 (N_7793,N_7410,N_7436);
and U7794 (N_7794,N_7086,N_7353);
and U7795 (N_7795,N_7421,N_7054);
and U7796 (N_7796,N_7339,N_7122);
xor U7797 (N_7797,N_7227,N_7144);
xor U7798 (N_7798,N_7127,N_7147);
and U7799 (N_7799,N_7494,N_7417);
or U7800 (N_7800,N_7087,N_7416);
or U7801 (N_7801,N_7369,N_7389);
nand U7802 (N_7802,N_7157,N_7042);
or U7803 (N_7803,N_7214,N_7021);
or U7804 (N_7804,N_7125,N_7444);
nor U7805 (N_7805,N_7025,N_7140);
or U7806 (N_7806,N_7320,N_7437);
or U7807 (N_7807,N_7088,N_7371);
and U7808 (N_7808,N_7414,N_7443);
nand U7809 (N_7809,N_7255,N_7032);
or U7810 (N_7810,N_7065,N_7433);
nor U7811 (N_7811,N_7223,N_7058);
or U7812 (N_7812,N_7382,N_7149);
xor U7813 (N_7813,N_7354,N_7204);
nor U7814 (N_7814,N_7385,N_7113);
or U7815 (N_7815,N_7346,N_7319);
xnor U7816 (N_7816,N_7469,N_7353);
nor U7817 (N_7817,N_7125,N_7144);
xor U7818 (N_7818,N_7063,N_7240);
xor U7819 (N_7819,N_7015,N_7285);
xor U7820 (N_7820,N_7438,N_7066);
xnor U7821 (N_7821,N_7270,N_7257);
nor U7822 (N_7822,N_7310,N_7472);
xor U7823 (N_7823,N_7356,N_7269);
and U7824 (N_7824,N_7291,N_7179);
nor U7825 (N_7825,N_7089,N_7122);
nor U7826 (N_7826,N_7321,N_7400);
or U7827 (N_7827,N_7307,N_7000);
or U7828 (N_7828,N_7010,N_7277);
nor U7829 (N_7829,N_7390,N_7468);
and U7830 (N_7830,N_7329,N_7095);
nand U7831 (N_7831,N_7343,N_7057);
or U7832 (N_7832,N_7320,N_7078);
xnor U7833 (N_7833,N_7048,N_7067);
xnor U7834 (N_7834,N_7305,N_7273);
nor U7835 (N_7835,N_7079,N_7330);
and U7836 (N_7836,N_7481,N_7050);
nand U7837 (N_7837,N_7363,N_7100);
or U7838 (N_7838,N_7133,N_7107);
nand U7839 (N_7839,N_7421,N_7286);
nor U7840 (N_7840,N_7050,N_7450);
and U7841 (N_7841,N_7407,N_7263);
xor U7842 (N_7842,N_7001,N_7339);
nor U7843 (N_7843,N_7027,N_7436);
nand U7844 (N_7844,N_7036,N_7185);
nand U7845 (N_7845,N_7440,N_7039);
and U7846 (N_7846,N_7158,N_7060);
or U7847 (N_7847,N_7286,N_7389);
and U7848 (N_7848,N_7403,N_7153);
nand U7849 (N_7849,N_7105,N_7446);
or U7850 (N_7850,N_7010,N_7196);
or U7851 (N_7851,N_7468,N_7459);
nand U7852 (N_7852,N_7327,N_7188);
nor U7853 (N_7853,N_7370,N_7235);
nor U7854 (N_7854,N_7112,N_7002);
xor U7855 (N_7855,N_7496,N_7454);
nor U7856 (N_7856,N_7036,N_7454);
xnor U7857 (N_7857,N_7144,N_7497);
xor U7858 (N_7858,N_7452,N_7062);
nor U7859 (N_7859,N_7084,N_7358);
xor U7860 (N_7860,N_7352,N_7073);
xnor U7861 (N_7861,N_7287,N_7302);
xor U7862 (N_7862,N_7366,N_7271);
and U7863 (N_7863,N_7475,N_7176);
or U7864 (N_7864,N_7450,N_7110);
or U7865 (N_7865,N_7316,N_7172);
or U7866 (N_7866,N_7119,N_7020);
nand U7867 (N_7867,N_7059,N_7274);
nor U7868 (N_7868,N_7228,N_7229);
xor U7869 (N_7869,N_7432,N_7385);
and U7870 (N_7870,N_7088,N_7194);
xor U7871 (N_7871,N_7435,N_7239);
and U7872 (N_7872,N_7287,N_7384);
or U7873 (N_7873,N_7230,N_7117);
and U7874 (N_7874,N_7412,N_7249);
xnor U7875 (N_7875,N_7391,N_7302);
nor U7876 (N_7876,N_7453,N_7188);
and U7877 (N_7877,N_7274,N_7131);
and U7878 (N_7878,N_7115,N_7005);
nand U7879 (N_7879,N_7188,N_7093);
and U7880 (N_7880,N_7453,N_7080);
nand U7881 (N_7881,N_7074,N_7000);
or U7882 (N_7882,N_7237,N_7306);
and U7883 (N_7883,N_7050,N_7375);
or U7884 (N_7884,N_7041,N_7166);
xor U7885 (N_7885,N_7073,N_7011);
xnor U7886 (N_7886,N_7481,N_7472);
xor U7887 (N_7887,N_7249,N_7286);
or U7888 (N_7888,N_7479,N_7436);
or U7889 (N_7889,N_7076,N_7065);
or U7890 (N_7890,N_7277,N_7360);
xor U7891 (N_7891,N_7447,N_7083);
nand U7892 (N_7892,N_7137,N_7063);
or U7893 (N_7893,N_7087,N_7482);
and U7894 (N_7894,N_7180,N_7492);
and U7895 (N_7895,N_7171,N_7310);
and U7896 (N_7896,N_7044,N_7442);
nor U7897 (N_7897,N_7292,N_7434);
or U7898 (N_7898,N_7133,N_7353);
or U7899 (N_7899,N_7475,N_7300);
xnor U7900 (N_7900,N_7032,N_7218);
nor U7901 (N_7901,N_7037,N_7402);
nor U7902 (N_7902,N_7246,N_7454);
or U7903 (N_7903,N_7155,N_7003);
nand U7904 (N_7904,N_7467,N_7227);
and U7905 (N_7905,N_7074,N_7262);
nor U7906 (N_7906,N_7275,N_7039);
xor U7907 (N_7907,N_7070,N_7407);
nor U7908 (N_7908,N_7378,N_7090);
xor U7909 (N_7909,N_7490,N_7429);
and U7910 (N_7910,N_7379,N_7186);
xnor U7911 (N_7911,N_7071,N_7218);
xor U7912 (N_7912,N_7020,N_7016);
and U7913 (N_7913,N_7075,N_7067);
and U7914 (N_7914,N_7046,N_7267);
and U7915 (N_7915,N_7480,N_7223);
xnor U7916 (N_7916,N_7169,N_7426);
nand U7917 (N_7917,N_7098,N_7267);
nand U7918 (N_7918,N_7284,N_7073);
and U7919 (N_7919,N_7431,N_7181);
or U7920 (N_7920,N_7470,N_7350);
or U7921 (N_7921,N_7445,N_7248);
xor U7922 (N_7922,N_7238,N_7377);
xor U7923 (N_7923,N_7130,N_7192);
or U7924 (N_7924,N_7279,N_7233);
nand U7925 (N_7925,N_7374,N_7340);
xor U7926 (N_7926,N_7273,N_7497);
nor U7927 (N_7927,N_7365,N_7047);
and U7928 (N_7928,N_7495,N_7017);
nand U7929 (N_7929,N_7311,N_7387);
nand U7930 (N_7930,N_7281,N_7449);
or U7931 (N_7931,N_7063,N_7203);
or U7932 (N_7932,N_7466,N_7133);
or U7933 (N_7933,N_7393,N_7477);
nor U7934 (N_7934,N_7484,N_7188);
or U7935 (N_7935,N_7167,N_7428);
nand U7936 (N_7936,N_7356,N_7396);
nor U7937 (N_7937,N_7017,N_7273);
and U7938 (N_7938,N_7456,N_7026);
or U7939 (N_7939,N_7498,N_7332);
xor U7940 (N_7940,N_7039,N_7062);
xnor U7941 (N_7941,N_7173,N_7427);
or U7942 (N_7942,N_7236,N_7093);
nand U7943 (N_7943,N_7124,N_7115);
and U7944 (N_7944,N_7187,N_7122);
nor U7945 (N_7945,N_7245,N_7260);
nor U7946 (N_7946,N_7053,N_7330);
nor U7947 (N_7947,N_7375,N_7319);
nor U7948 (N_7948,N_7087,N_7188);
nor U7949 (N_7949,N_7365,N_7101);
or U7950 (N_7950,N_7204,N_7073);
and U7951 (N_7951,N_7407,N_7468);
and U7952 (N_7952,N_7292,N_7395);
nand U7953 (N_7953,N_7069,N_7003);
xor U7954 (N_7954,N_7368,N_7152);
and U7955 (N_7955,N_7164,N_7418);
nor U7956 (N_7956,N_7309,N_7272);
nor U7957 (N_7957,N_7156,N_7400);
or U7958 (N_7958,N_7326,N_7053);
nor U7959 (N_7959,N_7171,N_7166);
xnor U7960 (N_7960,N_7102,N_7215);
or U7961 (N_7961,N_7400,N_7188);
or U7962 (N_7962,N_7421,N_7030);
or U7963 (N_7963,N_7292,N_7368);
and U7964 (N_7964,N_7038,N_7171);
xor U7965 (N_7965,N_7452,N_7491);
xnor U7966 (N_7966,N_7192,N_7364);
or U7967 (N_7967,N_7303,N_7340);
or U7968 (N_7968,N_7460,N_7379);
xor U7969 (N_7969,N_7457,N_7403);
nor U7970 (N_7970,N_7364,N_7302);
nand U7971 (N_7971,N_7335,N_7364);
xor U7972 (N_7972,N_7000,N_7293);
and U7973 (N_7973,N_7313,N_7164);
nand U7974 (N_7974,N_7115,N_7059);
nand U7975 (N_7975,N_7289,N_7174);
xnor U7976 (N_7976,N_7104,N_7195);
nor U7977 (N_7977,N_7406,N_7217);
and U7978 (N_7978,N_7042,N_7234);
and U7979 (N_7979,N_7145,N_7480);
nand U7980 (N_7980,N_7363,N_7454);
nand U7981 (N_7981,N_7303,N_7250);
xnor U7982 (N_7982,N_7087,N_7312);
xnor U7983 (N_7983,N_7074,N_7359);
and U7984 (N_7984,N_7211,N_7442);
or U7985 (N_7985,N_7084,N_7194);
nand U7986 (N_7986,N_7458,N_7422);
and U7987 (N_7987,N_7242,N_7233);
xnor U7988 (N_7988,N_7404,N_7017);
and U7989 (N_7989,N_7242,N_7162);
xnor U7990 (N_7990,N_7273,N_7342);
nand U7991 (N_7991,N_7405,N_7349);
nand U7992 (N_7992,N_7310,N_7482);
or U7993 (N_7993,N_7316,N_7470);
nor U7994 (N_7994,N_7400,N_7323);
nand U7995 (N_7995,N_7377,N_7000);
or U7996 (N_7996,N_7385,N_7078);
nor U7997 (N_7997,N_7220,N_7016);
nand U7998 (N_7998,N_7082,N_7299);
or U7999 (N_7999,N_7126,N_7160);
or U8000 (N_8000,N_7958,N_7763);
nor U8001 (N_8001,N_7922,N_7657);
and U8002 (N_8002,N_7955,N_7656);
xnor U8003 (N_8003,N_7533,N_7778);
or U8004 (N_8004,N_7721,N_7770);
xor U8005 (N_8005,N_7799,N_7658);
xnor U8006 (N_8006,N_7804,N_7758);
and U8007 (N_8007,N_7748,N_7983);
or U8008 (N_8008,N_7891,N_7565);
and U8009 (N_8009,N_7628,N_7764);
and U8010 (N_8010,N_7601,N_7619);
nor U8011 (N_8011,N_7775,N_7986);
or U8012 (N_8012,N_7609,N_7696);
nand U8013 (N_8013,N_7845,N_7887);
xor U8014 (N_8014,N_7669,N_7627);
or U8015 (N_8015,N_7898,N_7724);
or U8016 (N_8016,N_7671,N_7596);
nor U8017 (N_8017,N_7947,N_7713);
nor U8018 (N_8018,N_7966,N_7868);
nor U8019 (N_8019,N_7807,N_7733);
nor U8020 (N_8020,N_7528,N_7766);
nand U8021 (N_8021,N_7895,N_7684);
xor U8022 (N_8022,N_7916,N_7925);
or U8023 (N_8023,N_7964,N_7701);
xnor U8024 (N_8024,N_7641,N_7811);
nor U8025 (N_8025,N_7662,N_7755);
and U8026 (N_8026,N_7754,N_7564);
and U8027 (N_8027,N_7537,N_7783);
xnor U8028 (N_8028,N_7938,N_7523);
nand U8029 (N_8029,N_7995,N_7718);
and U8030 (N_8030,N_7526,N_7976);
and U8031 (N_8031,N_7560,N_7607);
nand U8032 (N_8032,N_7962,N_7844);
nor U8033 (N_8033,N_7604,N_7728);
and U8034 (N_8034,N_7625,N_7683);
and U8035 (N_8035,N_7984,N_7871);
or U8036 (N_8036,N_7990,N_7589);
or U8037 (N_8037,N_7847,N_7531);
or U8038 (N_8038,N_7644,N_7579);
or U8039 (N_8039,N_7914,N_7681);
nand U8040 (N_8040,N_7997,N_7841);
or U8041 (N_8041,N_7889,N_7586);
xnor U8042 (N_8042,N_7636,N_7720);
or U8043 (N_8043,N_7854,N_7591);
and U8044 (N_8044,N_7902,N_7682);
nor U8045 (N_8045,N_7869,N_7812);
or U8046 (N_8046,N_7858,N_7928);
nor U8047 (N_8047,N_7842,N_7524);
or U8048 (N_8048,N_7632,N_7943);
or U8049 (N_8049,N_7855,N_7687);
or U8050 (N_8050,N_7796,N_7715);
xor U8051 (N_8051,N_7837,N_7660);
and U8052 (N_8052,N_7861,N_7939);
nand U8053 (N_8053,N_7952,N_7985);
nor U8054 (N_8054,N_7832,N_7708);
nor U8055 (N_8055,N_7706,N_7890);
nand U8056 (N_8056,N_7867,N_7782);
nand U8057 (N_8057,N_7940,N_7882);
and U8058 (N_8058,N_7639,N_7840);
and U8059 (N_8059,N_7774,N_7618);
nor U8060 (N_8060,N_7529,N_7870);
nand U8061 (N_8061,N_7633,N_7768);
nand U8062 (N_8062,N_7810,N_7582);
nand U8063 (N_8063,N_7572,N_7828);
or U8064 (N_8064,N_7592,N_7742);
or U8065 (N_8065,N_7675,N_7825);
nor U8066 (N_8066,N_7703,N_7593);
nand U8067 (N_8067,N_7900,N_7667);
nand U8068 (N_8068,N_7920,N_7773);
or U8069 (N_8069,N_7629,N_7926);
or U8070 (N_8070,N_7583,N_7835);
or U8071 (N_8071,N_7747,N_7602);
nor U8072 (N_8072,N_7600,N_7500);
or U8073 (N_8073,N_7885,N_7893);
nor U8074 (N_8074,N_7874,N_7884);
and U8075 (N_8075,N_7935,N_7970);
and U8076 (N_8076,N_7559,N_7829);
nand U8077 (N_8077,N_7875,N_7744);
nand U8078 (N_8078,N_7651,N_7505);
and U8079 (N_8079,N_7663,N_7954);
nor U8080 (N_8080,N_7692,N_7553);
or U8081 (N_8081,N_7843,N_7848);
xor U8082 (N_8082,N_7732,N_7557);
xor U8083 (N_8083,N_7784,N_7833);
nor U8084 (N_8084,N_7992,N_7597);
nor U8085 (N_8085,N_7679,N_7739);
nand U8086 (N_8086,N_7963,N_7862);
nor U8087 (N_8087,N_7736,N_7624);
or U8088 (N_8088,N_7856,N_7513);
nand U8089 (N_8089,N_7896,N_7769);
and U8090 (N_8090,N_7697,N_7622);
xnor U8091 (N_8091,N_7717,N_7948);
nor U8092 (N_8092,N_7913,N_7876);
or U8093 (N_8093,N_7652,N_7959);
xor U8094 (N_8094,N_7821,N_7551);
or U8095 (N_8095,N_7637,N_7780);
nor U8096 (N_8096,N_7897,N_7611);
xnor U8097 (N_8097,N_7568,N_7555);
nor U8098 (N_8098,N_7719,N_7688);
xnor U8099 (N_8099,N_7788,N_7511);
or U8100 (N_8100,N_7594,N_7953);
nand U8101 (N_8101,N_7677,N_7826);
xor U8102 (N_8102,N_7509,N_7908);
nand U8103 (N_8103,N_7647,N_7806);
nand U8104 (N_8104,N_7642,N_7886);
nand U8105 (N_8105,N_7792,N_7950);
xnor U8106 (N_8106,N_7814,N_7571);
nor U8107 (N_8107,N_7921,N_7978);
nor U8108 (N_8108,N_7694,N_7534);
nor U8109 (N_8109,N_7653,N_7960);
and U8110 (N_8110,N_7504,N_7936);
or U8111 (N_8111,N_7573,N_7542);
xor U8112 (N_8112,N_7535,N_7779);
or U8113 (N_8113,N_7888,N_7543);
xor U8114 (N_8114,N_7574,N_7680);
nor U8115 (N_8115,N_7693,N_7975);
or U8116 (N_8116,N_7909,N_7819);
nand U8117 (N_8117,N_7516,N_7723);
xnor U8118 (N_8118,N_7530,N_7836);
xor U8119 (N_8119,N_7969,N_7989);
nand U8120 (N_8120,N_7654,N_7793);
or U8121 (N_8121,N_7743,N_7917);
or U8122 (N_8122,N_7585,N_7631);
or U8123 (N_8123,N_7704,N_7546);
nor U8124 (N_8124,N_7690,N_7612);
or U8125 (N_8125,N_7981,N_7570);
or U8126 (N_8126,N_7839,N_7621);
or U8127 (N_8127,N_7588,N_7772);
xnor U8128 (N_8128,N_7857,N_7664);
xor U8129 (N_8129,N_7991,N_7711);
and U8130 (N_8130,N_7967,N_7761);
nor U8131 (N_8131,N_7831,N_7577);
nor U8132 (N_8132,N_7725,N_7980);
and U8133 (N_8133,N_7562,N_7918);
nor U8134 (N_8134,N_7808,N_7613);
or U8135 (N_8135,N_7581,N_7522);
and U8136 (N_8136,N_7595,N_7749);
nand U8137 (N_8137,N_7503,N_7757);
and U8138 (N_8138,N_7903,N_7996);
nor U8139 (N_8139,N_7659,N_7700);
xnor U8140 (N_8140,N_7547,N_7813);
nor U8141 (N_8141,N_7982,N_7698);
or U8142 (N_8142,N_7797,N_7883);
xnor U8143 (N_8143,N_7751,N_7750);
nor U8144 (N_8144,N_7899,N_7666);
nand U8145 (N_8145,N_7638,N_7853);
and U8146 (N_8146,N_7605,N_7809);
or U8147 (N_8147,N_7735,N_7881);
nand U8148 (N_8148,N_7803,N_7942);
and U8149 (N_8149,N_7575,N_7510);
or U8150 (N_8150,N_7822,N_7923);
or U8151 (N_8151,N_7635,N_7536);
xor U8152 (N_8152,N_7860,N_7722);
nand U8153 (N_8153,N_7645,N_7610);
nor U8154 (N_8154,N_7762,N_7599);
nor U8155 (N_8155,N_7643,N_7740);
nor U8156 (N_8156,N_7506,N_7834);
nor U8157 (N_8157,N_7608,N_7924);
nand U8158 (N_8158,N_7872,N_7702);
nand U8159 (N_8159,N_7672,N_7771);
nor U8160 (N_8160,N_7691,N_7576);
nor U8161 (N_8161,N_7616,N_7512);
or U8162 (N_8162,N_7539,N_7998);
xnor U8163 (N_8163,N_7846,N_7630);
nand U8164 (N_8164,N_7729,N_7668);
or U8165 (N_8165,N_7805,N_7518);
nand U8166 (N_8166,N_7752,N_7710);
nand U8167 (N_8167,N_7907,N_7532);
and U8168 (N_8168,N_7606,N_7765);
or U8169 (N_8169,N_7864,N_7695);
xnor U8170 (N_8170,N_7946,N_7877);
and U8171 (N_8171,N_7879,N_7915);
or U8172 (N_8172,N_7930,N_7540);
and U8173 (N_8173,N_7927,N_7988);
nor U8174 (N_8174,N_7714,N_7971);
or U8175 (N_8175,N_7767,N_7745);
and U8176 (N_8176,N_7649,N_7911);
xnor U8177 (N_8177,N_7965,N_7919);
nor U8178 (N_8178,N_7521,N_7685);
and U8179 (N_8179,N_7686,N_7678);
and U8180 (N_8180,N_7567,N_7705);
nor U8181 (N_8181,N_7515,N_7646);
xnor U8182 (N_8182,N_7738,N_7957);
xor U8183 (N_8183,N_7552,N_7554);
nor U8184 (N_8184,N_7852,N_7712);
or U8185 (N_8185,N_7508,N_7756);
xnor U8186 (N_8186,N_7781,N_7820);
nand U8187 (N_8187,N_7838,N_7650);
xnor U8188 (N_8188,N_7906,N_7801);
and U8189 (N_8189,N_7785,N_7753);
and U8190 (N_8190,N_7626,N_7640);
and U8191 (N_8191,N_7727,N_7961);
and U8192 (N_8192,N_7910,N_7556);
or U8193 (N_8193,N_7731,N_7746);
and U8194 (N_8194,N_7949,N_7550);
nand U8195 (N_8195,N_7561,N_7791);
or U8196 (N_8196,N_7865,N_7620);
nor U8197 (N_8197,N_7502,N_7979);
nor U8198 (N_8198,N_7880,N_7507);
and U8199 (N_8199,N_7514,N_7674);
nand U8200 (N_8200,N_7587,N_7993);
nand U8201 (N_8201,N_7972,N_7905);
nand U8202 (N_8202,N_7544,N_7863);
nand U8203 (N_8203,N_7818,N_7665);
nor U8204 (N_8204,N_7517,N_7802);
nand U8205 (N_8205,N_7933,N_7634);
nor U8206 (N_8206,N_7878,N_7563);
xor U8207 (N_8207,N_7707,N_7789);
nor U8208 (N_8208,N_7937,N_7859);
nor U8209 (N_8209,N_7538,N_7527);
nor U8210 (N_8210,N_7850,N_7790);
or U8211 (N_8211,N_7968,N_7987);
nor U8212 (N_8212,N_7892,N_7932);
or U8213 (N_8213,N_7520,N_7541);
nor U8214 (N_8214,N_7670,N_7974);
nand U8215 (N_8215,N_7584,N_7615);
or U8216 (N_8216,N_7734,N_7759);
or U8217 (N_8217,N_7912,N_7548);
nor U8218 (N_8218,N_7929,N_7944);
nor U8219 (N_8219,N_7873,N_7815);
nand U8220 (N_8220,N_7777,N_7798);
nor U8221 (N_8221,N_7590,N_7578);
xnor U8222 (N_8222,N_7941,N_7676);
or U8223 (N_8223,N_7786,N_7566);
nor U8224 (N_8224,N_7956,N_7730);
nor U8225 (N_8225,N_7977,N_7824);
or U8226 (N_8226,N_7617,N_7994);
xnor U8227 (N_8227,N_7549,N_7525);
and U8228 (N_8228,N_7951,N_7741);
nor U8229 (N_8229,N_7849,N_7699);
nor U8230 (N_8230,N_7737,N_7904);
nand U8231 (N_8231,N_7931,N_7501);
or U8232 (N_8232,N_7661,N_7519);
nor U8233 (N_8233,N_7603,N_7973);
nor U8234 (N_8234,N_7614,N_7851);
nand U8235 (N_8235,N_7794,N_7623);
and U8236 (N_8236,N_7569,N_7866);
xor U8237 (N_8237,N_7817,N_7558);
nand U8238 (N_8238,N_7894,N_7598);
and U8239 (N_8239,N_7689,N_7945);
or U8240 (N_8240,N_7655,N_7673);
nand U8241 (N_8241,N_7901,N_7648);
nand U8242 (N_8242,N_7830,N_7795);
nor U8243 (N_8243,N_7823,N_7716);
and U8244 (N_8244,N_7800,N_7816);
and U8245 (N_8245,N_7999,N_7760);
and U8246 (N_8246,N_7580,N_7545);
xor U8247 (N_8247,N_7827,N_7787);
or U8248 (N_8248,N_7776,N_7934);
nor U8249 (N_8249,N_7726,N_7709);
xnor U8250 (N_8250,N_7985,N_7600);
and U8251 (N_8251,N_7904,N_7933);
nor U8252 (N_8252,N_7891,N_7743);
nand U8253 (N_8253,N_7511,N_7823);
nor U8254 (N_8254,N_7968,N_7783);
nand U8255 (N_8255,N_7611,N_7916);
or U8256 (N_8256,N_7822,N_7604);
xor U8257 (N_8257,N_7848,N_7696);
and U8258 (N_8258,N_7746,N_7824);
nand U8259 (N_8259,N_7897,N_7816);
and U8260 (N_8260,N_7846,N_7751);
nand U8261 (N_8261,N_7732,N_7837);
and U8262 (N_8262,N_7828,N_7732);
nand U8263 (N_8263,N_7843,N_7791);
and U8264 (N_8264,N_7542,N_7850);
nand U8265 (N_8265,N_7544,N_7993);
or U8266 (N_8266,N_7832,N_7954);
or U8267 (N_8267,N_7919,N_7691);
or U8268 (N_8268,N_7554,N_7900);
nor U8269 (N_8269,N_7962,N_7876);
and U8270 (N_8270,N_7904,N_7602);
xor U8271 (N_8271,N_7569,N_7566);
xor U8272 (N_8272,N_7853,N_7962);
and U8273 (N_8273,N_7762,N_7910);
nand U8274 (N_8274,N_7822,N_7506);
xnor U8275 (N_8275,N_7542,N_7570);
nand U8276 (N_8276,N_7582,N_7982);
xnor U8277 (N_8277,N_7872,N_7880);
xor U8278 (N_8278,N_7713,N_7588);
or U8279 (N_8279,N_7919,N_7546);
nor U8280 (N_8280,N_7832,N_7727);
nor U8281 (N_8281,N_7818,N_7895);
nand U8282 (N_8282,N_7692,N_7859);
or U8283 (N_8283,N_7504,N_7907);
xor U8284 (N_8284,N_7619,N_7533);
nand U8285 (N_8285,N_7874,N_7554);
nand U8286 (N_8286,N_7997,N_7874);
nand U8287 (N_8287,N_7851,N_7649);
and U8288 (N_8288,N_7843,N_7908);
and U8289 (N_8289,N_7723,N_7576);
nand U8290 (N_8290,N_7605,N_7616);
nand U8291 (N_8291,N_7881,N_7653);
and U8292 (N_8292,N_7686,N_7672);
nand U8293 (N_8293,N_7960,N_7936);
xnor U8294 (N_8294,N_7943,N_7588);
or U8295 (N_8295,N_7765,N_7908);
nand U8296 (N_8296,N_7616,N_7886);
xnor U8297 (N_8297,N_7845,N_7768);
nand U8298 (N_8298,N_7933,N_7608);
nand U8299 (N_8299,N_7695,N_7595);
nand U8300 (N_8300,N_7880,N_7548);
nand U8301 (N_8301,N_7826,N_7608);
nor U8302 (N_8302,N_7674,N_7529);
nor U8303 (N_8303,N_7779,N_7866);
or U8304 (N_8304,N_7945,N_7539);
or U8305 (N_8305,N_7748,N_7772);
xnor U8306 (N_8306,N_7561,N_7534);
nor U8307 (N_8307,N_7925,N_7594);
nor U8308 (N_8308,N_7804,N_7787);
or U8309 (N_8309,N_7943,N_7713);
nand U8310 (N_8310,N_7883,N_7972);
or U8311 (N_8311,N_7608,N_7866);
or U8312 (N_8312,N_7921,N_7746);
nor U8313 (N_8313,N_7647,N_7876);
or U8314 (N_8314,N_7533,N_7639);
xnor U8315 (N_8315,N_7714,N_7886);
nand U8316 (N_8316,N_7564,N_7846);
nand U8317 (N_8317,N_7589,N_7669);
or U8318 (N_8318,N_7706,N_7919);
and U8319 (N_8319,N_7961,N_7505);
and U8320 (N_8320,N_7667,N_7526);
nor U8321 (N_8321,N_7784,N_7691);
or U8322 (N_8322,N_7966,N_7830);
or U8323 (N_8323,N_7543,N_7771);
nor U8324 (N_8324,N_7704,N_7727);
xor U8325 (N_8325,N_7813,N_7730);
nand U8326 (N_8326,N_7573,N_7544);
and U8327 (N_8327,N_7619,N_7807);
nor U8328 (N_8328,N_7541,N_7745);
xnor U8329 (N_8329,N_7891,N_7835);
xor U8330 (N_8330,N_7765,N_7928);
or U8331 (N_8331,N_7703,N_7807);
nor U8332 (N_8332,N_7992,N_7516);
or U8333 (N_8333,N_7869,N_7805);
nor U8334 (N_8334,N_7833,N_7574);
and U8335 (N_8335,N_7613,N_7862);
nor U8336 (N_8336,N_7692,N_7749);
and U8337 (N_8337,N_7667,N_7500);
xor U8338 (N_8338,N_7925,N_7850);
or U8339 (N_8339,N_7764,N_7700);
or U8340 (N_8340,N_7636,N_7718);
or U8341 (N_8341,N_7799,N_7955);
and U8342 (N_8342,N_7659,N_7766);
nand U8343 (N_8343,N_7609,N_7506);
nand U8344 (N_8344,N_7730,N_7888);
and U8345 (N_8345,N_7955,N_7655);
and U8346 (N_8346,N_7679,N_7507);
nor U8347 (N_8347,N_7594,N_7770);
nor U8348 (N_8348,N_7523,N_7845);
nor U8349 (N_8349,N_7534,N_7775);
nand U8350 (N_8350,N_7759,N_7968);
and U8351 (N_8351,N_7882,N_7611);
nand U8352 (N_8352,N_7577,N_7729);
xor U8353 (N_8353,N_7738,N_7830);
or U8354 (N_8354,N_7881,N_7984);
xnor U8355 (N_8355,N_7631,N_7786);
xor U8356 (N_8356,N_7743,N_7826);
xor U8357 (N_8357,N_7882,N_7802);
and U8358 (N_8358,N_7606,N_7558);
xnor U8359 (N_8359,N_7992,N_7987);
xor U8360 (N_8360,N_7608,N_7945);
nor U8361 (N_8361,N_7959,N_7562);
nand U8362 (N_8362,N_7631,N_7850);
xnor U8363 (N_8363,N_7521,N_7665);
nor U8364 (N_8364,N_7629,N_7734);
nand U8365 (N_8365,N_7778,N_7717);
xnor U8366 (N_8366,N_7847,N_7611);
xnor U8367 (N_8367,N_7503,N_7928);
xnor U8368 (N_8368,N_7763,N_7658);
xnor U8369 (N_8369,N_7915,N_7820);
and U8370 (N_8370,N_7837,N_7939);
and U8371 (N_8371,N_7796,N_7552);
and U8372 (N_8372,N_7558,N_7873);
or U8373 (N_8373,N_7549,N_7821);
or U8374 (N_8374,N_7988,N_7530);
or U8375 (N_8375,N_7732,N_7723);
nor U8376 (N_8376,N_7654,N_7807);
and U8377 (N_8377,N_7519,N_7566);
and U8378 (N_8378,N_7649,N_7591);
xor U8379 (N_8379,N_7578,N_7797);
or U8380 (N_8380,N_7891,N_7583);
nand U8381 (N_8381,N_7652,N_7867);
xnor U8382 (N_8382,N_7793,N_7717);
or U8383 (N_8383,N_7881,N_7747);
xnor U8384 (N_8384,N_7792,N_7898);
nor U8385 (N_8385,N_7523,N_7760);
and U8386 (N_8386,N_7729,N_7672);
xnor U8387 (N_8387,N_7983,N_7917);
nor U8388 (N_8388,N_7930,N_7820);
and U8389 (N_8389,N_7810,N_7910);
and U8390 (N_8390,N_7902,N_7773);
or U8391 (N_8391,N_7590,N_7838);
nor U8392 (N_8392,N_7805,N_7715);
and U8393 (N_8393,N_7782,N_7614);
or U8394 (N_8394,N_7663,N_7720);
nand U8395 (N_8395,N_7644,N_7622);
or U8396 (N_8396,N_7549,N_7531);
nor U8397 (N_8397,N_7840,N_7903);
or U8398 (N_8398,N_7616,N_7692);
and U8399 (N_8399,N_7780,N_7842);
xnor U8400 (N_8400,N_7801,N_7722);
xor U8401 (N_8401,N_7556,N_7836);
or U8402 (N_8402,N_7695,N_7749);
or U8403 (N_8403,N_7644,N_7506);
or U8404 (N_8404,N_7700,N_7849);
nand U8405 (N_8405,N_7531,N_7522);
and U8406 (N_8406,N_7858,N_7872);
or U8407 (N_8407,N_7904,N_7567);
and U8408 (N_8408,N_7721,N_7960);
and U8409 (N_8409,N_7841,N_7823);
nand U8410 (N_8410,N_7613,N_7567);
and U8411 (N_8411,N_7671,N_7986);
or U8412 (N_8412,N_7695,N_7786);
nor U8413 (N_8413,N_7555,N_7871);
or U8414 (N_8414,N_7830,N_7667);
nand U8415 (N_8415,N_7784,N_7528);
nor U8416 (N_8416,N_7584,N_7518);
nand U8417 (N_8417,N_7570,N_7596);
and U8418 (N_8418,N_7732,N_7727);
xor U8419 (N_8419,N_7906,N_7904);
nand U8420 (N_8420,N_7829,N_7766);
or U8421 (N_8421,N_7655,N_7681);
or U8422 (N_8422,N_7870,N_7899);
or U8423 (N_8423,N_7726,N_7581);
nand U8424 (N_8424,N_7501,N_7769);
and U8425 (N_8425,N_7838,N_7906);
nor U8426 (N_8426,N_7537,N_7634);
nand U8427 (N_8427,N_7915,N_7587);
xor U8428 (N_8428,N_7911,N_7755);
nor U8429 (N_8429,N_7829,N_7546);
and U8430 (N_8430,N_7731,N_7562);
or U8431 (N_8431,N_7849,N_7734);
or U8432 (N_8432,N_7966,N_7781);
and U8433 (N_8433,N_7832,N_7740);
nor U8434 (N_8434,N_7744,N_7918);
nor U8435 (N_8435,N_7704,N_7600);
xnor U8436 (N_8436,N_7728,N_7610);
and U8437 (N_8437,N_7857,N_7718);
and U8438 (N_8438,N_7520,N_7606);
and U8439 (N_8439,N_7906,N_7705);
and U8440 (N_8440,N_7739,N_7975);
nand U8441 (N_8441,N_7678,N_7828);
nand U8442 (N_8442,N_7710,N_7775);
and U8443 (N_8443,N_7788,N_7882);
nand U8444 (N_8444,N_7678,N_7919);
or U8445 (N_8445,N_7761,N_7789);
or U8446 (N_8446,N_7729,N_7883);
or U8447 (N_8447,N_7944,N_7531);
nand U8448 (N_8448,N_7887,N_7546);
or U8449 (N_8449,N_7583,N_7915);
or U8450 (N_8450,N_7575,N_7552);
nor U8451 (N_8451,N_7812,N_7553);
and U8452 (N_8452,N_7861,N_7966);
or U8453 (N_8453,N_7513,N_7871);
nand U8454 (N_8454,N_7547,N_7713);
and U8455 (N_8455,N_7655,N_7869);
nor U8456 (N_8456,N_7545,N_7944);
nor U8457 (N_8457,N_7823,N_7628);
or U8458 (N_8458,N_7799,N_7642);
and U8459 (N_8459,N_7977,N_7701);
nor U8460 (N_8460,N_7923,N_7882);
nand U8461 (N_8461,N_7788,N_7845);
or U8462 (N_8462,N_7556,N_7948);
and U8463 (N_8463,N_7808,N_7643);
and U8464 (N_8464,N_7983,N_7615);
nand U8465 (N_8465,N_7659,N_7988);
nand U8466 (N_8466,N_7631,N_7976);
or U8467 (N_8467,N_7510,N_7613);
xnor U8468 (N_8468,N_7986,N_7668);
and U8469 (N_8469,N_7998,N_7934);
and U8470 (N_8470,N_7781,N_7687);
and U8471 (N_8471,N_7787,N_7779);
and U8472 (N_8472,N_7807,N_7802);
xor U8473 (N_8473,N_7899,N_7887);
nand U8474 (N_8474,N_7880,N_7827);
or U8475 (N_8475,N_7528,N_7749);
and U8476 (N_8476,N_7892,N_7798);
or U8477 (N_8477,N_7545,N_7512);
nand U8478 (N_8478,N_7610,N_7854);
or U8479 (N_8479,N_7927,N_7937);
xnor U8480 (N_8480,N_7902,N_7917);
or U8481 (N_8481,N_7769,N_7548);
and U8482 (N_8482,N_7574,N_7915);
nand U8483 (N_8483,N_7685,N_7795);
nor U8484 (N_8484,N_7692,N_7945);
or U8485 (N_8485,N_7691,N_7850);
or U8486 (N_8486,N_7679,N_7740);
and U8487 (N_8487,N_7852,N_7978);
or U8488 (N_8488,N_7900,N_7999);
nor U8489 (N_8489,N_7809,N_7983);
or U8490 (N_8490,N_7909,N_7600);
xnor U8491 (N_8491,N_7745,N_7823);
nand U8492 (N_8492,N_7650,N_7601);
xnor U8493 (N_8493,N_7834,N_7582);
and U8494 (N_8494,N_7502,N_7985);
or U8495 (N_8495,N_7807,N_7595);
and U8496 (N_8496,N_7764,N_7788);
xnor U8497 (N_8497,N_7730,N_7983);
xnor U8498 (N_8498,N_7984,N_7831);
or U8499 (N_8499,N_7545,N_7916);
nand U8500 (N_8500,N_8291,N_8364);
nand U8501 (N_8501,N_8160,N_8258);
nor U8502 (N_8502,N_8400,N_8385);
xor U8503 (N_8503,N_8222,N_8138);
or U8504 (N_8504,N_8271,N_8351);
nor U8505 (N_8505,N_8215,N_8495);
xnor U8506 (N_8506,N_8022,N_8113);
nor U8507 (N_8507,N_8116,N_8050);
nor U8508 (N_8508,N_8273,N_8319);
and U8509 (N_8509,N_8217,N_8392);
or U8510 (N_8510,N_8081,N_8092);
or U8511 (N_8511,N_8387,N_8309);
nor U8512 (N_8512,N_8410,N_8482);
xnor U8513 (N_8513,N_8338,N_8292);
xnor U8514 (N_8514,N_8356,N_8213);
xor U8515 (N_8515,N_8305,N_8150);
or U8516 (N_8516,N_8268,N_8257);
nor U8517 (N_8517,N_8123,N_8151);
or U8518 (N_8518,N_8036,N_8287);
xnor U8519 (N_8519,N_8360,N_8326);
and U8520 (N_8520,N_8183,N_8030);
xor U8521 (N_8521,N_8432,N_8467);
nor U8522 (N_8522,N_8401,N_8494);
nand U8523 (N_8523,N_8015,N_8005);
nand U8524 (N_8524,N_8203,N_8204);
nand U8525 (N_8525,N_8358,N_8155);
and U8526 (N_8526,N_8377,N_8145);
nor U8527 (N_8527,N_8297,N_8043);
and U8528 (N_8528,N_8199,N_8352);
nand U8529 (N_8529,N_8454,N_8422);
nand U8530 (N_8530,N_8394,N_8375);
or U8531 (N_8531,N_8411,N_8052);
xor U8532 (N_8532,N_8485,N_8069);
xor U8533 (N_8533,N_8206,N_8107);
nor U8534 (N_8534,N_8104,N_8282);
nand U8535 (N_8535,N_8135,N_8261);
nand U8536 (N_8536,N_8314,N_8103);
and U8537 (N_8537,N_8253,N_8339);
xnor U8538 (N_8538,N_8279,N_8429);
or U8539 (N_8539,N_8265,N_8168);
nand U8540 (N_8540,N_8404,N_8438);
or U8541 (N_8541,N_8105,N_8070);
nand U8542 (N_8542,N_8235,N_8472);
nand U8543 (N_8543,N_8493,N_8024);
nor U8544 (N_8544,N_8062,N_8446);
and U8545 (N_8545,N_8254,N_8252);
nand U8546 (N_8546,N_8491,N_8376);
nor U8547 (N_8547,N_8322,N_8018);
or U8548 (N_8548,N_8255,N_8437);
xor U8549 (N_8549,N_8014,N_8124);
xor U8550 (N_8550,N_8122,N_8011);
and U8551 (N_8551,N_8250,N_8097);
and U8552 (N_8552,N_8276,N_8185);
xor U8553 (N_8553,N_8205,N_8266);
nor U8554 (N_8554,N_8051,N_8263);
nand U8555 (N_8555,N_8108,N_8238);
and U8556 (N_8556,N_8397,N_8285);
xor U8557 (N_8557,N_8182,N_8269);
nand U8558 (N_8558,N_8281,N_8186);
nand U8559 (N_8559,N_8169,N_8148);
nand U8560 (N_8560,N_8329,N_8361);
xor U8561 (N_8561,N_8100,N_8114);
xnor U8562 (N_8562,N_8398,N_8020);
nand U8563 (N_8563,N_8045,N_8307);
and U8564 (N_8564,N_8165,N_8334);
xor U8565 (N_8565,N_8032,N_8000);
and U8566 (N_8566,N_8303,N_8037);
nor U8567 (N_8567,N_8370,N_8126);
xnor U8568 (N_8568,N_8301,N_8059);
and U8569 (N_8569,N_8463,N_8178);
or U8570 (N_8570,N_8068,N_8080);
nand U8571 (N_8571,N_8284,N_8106);
or U8572 (N_8572,N_8099,N_8171);
or U8573 (N_8573,N_8187,N_8146);
nor U8574 (N_8574,N_8140,N_8378);
and U8575 (N_8575,N_8402,N_8490);
nor U8576 (N_8576,N_8328,N_8053);
nand U8577 (N_8577,N_8308,N_8181);
nor U8578 (N_8578,N_8009,N_8101);
nor U8579 (N_8579,N_8312,N_8163);
xnor U8580 (N_8580,N_8419,N_8465);
nor U8581 (N_8581,N_8211,N_8445);
or U8582 (N_8582,N_8343,N_8336);
xor U8583 (N_8583,N_8086,N_8142);
nand U8584 (N_8584,N_8195,N_8440);
nor U8585 (N_8585,N_8486,N_8412);
xor U8586 (N_8586,N_8335,N_8063);
xnor U8587 (N_8587,N_8190,N_8324);
or U8588 (N_8588,N_8026,N_8479);
nor U8589 (N_8589,N_8028,N_8202);
and U8590 (N_8590,N_8089,N_8004);
nor U8591 (N_8591,N_8354,N_8434);
nor U8592 (N_8592,N_8363,N_8112);
or U8593 (N_8593,N_8492,N_8128);
or U8594 (N_8594,N_8272,N_8316);
and U8595 (N_8595,N_8407,N_8427);
xor U8596 (N_8596,N_8221,N_8460);
nor U8597 (N_8597,N_8001,N_8130);
and U8598 (N_8598,N_8212,N_8289);
nand U8599 (N_8599,N_8313,N_8477);
and U8600 (N_8600,N_8264,N_8321);
xor U8601 (N_8601,N_8158,N_8295);
or U8602 (N_8602,N_8139,N_8457);
nand U8603 (N_8603,N_8210,N_8172);
and U8604 (N_8604,N_8023,N_8164);
or U8605 (N_8605,N_8323,N_8173);
nor U8606 (N_8606,N_8236,N_8248);
or U8607 (N_8607,N_8056,N_8071);
and U8608 (N_8608,N_8391,N_8499);
nor U8609 (N_8609,N_8484,N_8161);
nor U8610 (N_8610,N_8175,N_8027);
nand U8611 (N_8611,N_8405,N_8403);
nand U8612 (N_8612,N_8047,N_8380);
nor U8613 (N_8613,N_8331,N_8017);
xnor U8614 (N_8614,N_8159,N_8251);
xnor U8615 (N_8615,N_8325,N_8474);
or U8616 (N_8616,N_8156,N_8357);
nand U8617 (N_8617,N_8218,N_8274);
or U8618 (N_8618,N_8353,N_8332);
and U8619 (N_8619,N_8125,N_8077);
xnor U8620 (N_8620,N_8283,N_8049);
nor U8621 (N_8621,N_8483,N_8421);
nand U8622 (N_8622,N_8249,N_8079);
or U8623 (N_8623,N_8216,N_8367);
nand U8624 (N_8624,N_8451,N_8180);
or U8625 (N_8625,N_8496,N_8153);
nand U8626 (N_8626,N_8388,N_8386);
and U8627 (N_8627,N_8447,N_8428);
nor U8628 (N_8628,N_8290,N_8245);
nand U8629 (N_8629,N_8072,N_8455);
xnor U8630 (N_8630,N_8476,N_8228);
nand U8631 (N_8631,N_8346,N_8021);
nor U8632 (N_8632,N_8144,N_8433);
and U8633 (N_8633,N_8085,N_8067);
and U8634 (N_8634,N_8008,N_8372);
nor U8635 (N_8635,N_8132,N_8176);
xnor U8636 (N_8636,N_8487,N_8298);
nor U8637 (N_8637,N_8340,N_8296);
nand U8638 (N_8638,N_8087,N_8311);
and U8639 (N_8639,N_8304,N_8119);
nand U8640 (N_8640,N_8090,N_8083);
and U8641 (N_8641,N_8461,N_8420);
nor U8642 (N_8642,N_8209,N_8064);
and U8643 (N_8643,N_8136,N_8439);
and U8644 (N_8644,N_8365,N_8031);
xor U8645 (N_8645,N_8054,N_8111);
nand U8646 (N_8646,N_8348,N_8393);
xor U8647 (N_8647,N_8147,N_8016);
and U8648 (N_8648,N_8430,N_8157);
nand U8649 (N_8649,N_8078,N_8044);
nor U8650 (N_8650,N_8371,N_8344);
nand U8651 (N_8651,N_8260,N_8013);
or U8652 (N_8652,N_8224,N_8462);
nand U8653 (N_8653,N_8489,N_8154);
nor U8654 (N_8654,N_8207,N_8057);
nand U8655 (N_8655,N_8425,N_8456);
or U8656 (N_8656,N_8241,N_8424);
or U8657 (N_8657,N_8058,N_8127);
and U8658 (N_8658,N_8368,N_8450);
nor U8659 (N_8659,N_8184,N_8098);
nor U8660 (N_8660,N_8219,N_8464);
nor U8661 (N_8661,N_8441,N_8470);
or U8662 (N_8662,N_8243,N_8196);
or U8663 (N_8663,N_8042,N_8449);
and U8664 (N_8664,N_8084,N_8347);
or U8665 (N_8665,N_8019,N_8345);
and U8666 (N_8666,N_8468,N_8229);
nor U8667 (N_8667,N_8166,N_8442);
or U8668 (N_8668,N_8436,N_8234);
nand U8669 (N_8669,N_8162,N_8231);
or U8670 (N_8670,N_8133,N_8208);
or U8671 (N_8671,N_8034,N_8118);
nand U8672 (N_8672,N_8406,N_8362);
and U8673 (N_8673,N_8369,N_8395);
and U8674 (N_8674,N_8137,N_8275);
nand U8675 (N_8675,N_8115,N_8244);
xor U8676 (N_8676,N_8038,N_8060);
xnor U8677 (N_8677,N_8342,N_8179);
nand U8678 (N_8678,N_8220,N_8239);
nor U8679 (N_8679,N_8223,N_8414);
nand U8680 (N_8680,N_8143,N_8498);
and U8681 (N_8681,N_8390,N_8189);
or U8682 (N_8682,N_8277,N_8010);
nor U8683 (N_8683,N_8227,N_8497);
nand U8684 (N_8684,N_8481,N_8444);
xor U8685 (N_8685,N_8233,N_8214);
xnor U8686 (N_8686,N_8413,N_8330);
nand U8687 (N_8687,N_8041,N_8471);
nor U8688 (N_8688,N_8006,N_8374);
xnor U8689 (N_8689,N_8102,N_8299);
xnor U8690 (N_8690,N_8240,N_8192);
nor U8691 (N_8691,N_8046,N_8093);
and U8692 (N_8692,N_8035,N_8306);
xor U8693 (N_8693,N_8418,N_8431);
nand U8694 (N_8694,N_8278,N_8055);
or U8695 (N_8695,N_8256,N_8327);
nand U8696 (N_8696,N_8315,N_8423);
or U8697 (N_8697,N_8293,N_8480);
xnor U8698 (N_8698,N_8452,N_8318);
xnor U8699 (N_8699,N_8094,N_8366);
and U8700 (N_8700,N_8134,N_8225);
nor U8701 (N_8701,N_8488,N_8170);
nand U8702 (N_8702,N_8040,N_8141);
or U8703 (N_8703,N_8262,N_8478);
xor U8704 (N_8704,N_8242,N_8076);
or U8705 (N_8705,N_8226,N_8232);
nand U8706 (N_8706,N_8458,N_8310);
xor U8707 (N_8707,N_8129,N_8095);
xor U8708 (N_8708,N_8201,N_8191);
nand U8709 (N_8709,N_8435,N_8389);
or U8710 (N_8710,N_8443,N_8174);
or U8711 (N_8711,N_8198,N_8003);
nor U8712 (N_8712,N_8025,N_8197);
and U8713 (N_8713,N_8259,N_8088);
nor U8714 (N_8714,N_8409,N_8333);
or U8715 (N_8715,N_8396,N_8317);
nand U8716 (N_8716,N_8373,N_8012);
nand U8717 (N_8717,N_8300,N_8383);
nor U8718 (N_8718,N_8152,N_8475);
nand U8719 (N_8719,N_8075,N_8074);
xor U8720 (N_8720,N_8466,N_8247);
nor U8721 (N_8721,N_8417,N_8415);
nand U8722 (N_8722,N_8048,N_8381);
xnor U8723 (N_8723,N_8473,N_8121);
nor U8724 (N_8724,N_8110,N_8448);
and U8725 (N_8725,N_8302,N_8061);
nor U8726 (N_8726,N_8073,N_8007);
nand U8727 (N_8727,N_8355,N_8091);
and U8728 (N_8728,N_8453,N_8426);
xor U8729 (N_8729,N_8270,N_8131);
nand U8730 (N_8730,N_8349,N_8200);
nor U8731 (N_8731,N_8350,N_8359);
nand U8732 (N_8732,N_8416,N_8029);
nor U8733 (N_8733,N_8194,N_8337);
nor U8734 (N_8734,N_8379,N_8288);
or U8735 (N_8735,N_8177,N_8246);
or U8736 (N_8736,N_8237,N_8033);
nand U8737 (N_8737,N_8167,N_8280);
nand U8738 (N_8738,N_8066,N_8384);
xor U8739 (N_8739,N_8408,N_8120);
nand U8740 (N_8740,N_8459,N_8320);
or U8741 (N_8741,N_8117,N_8109);
nor U8742 (N_8742,N_8082,N_8065);
xnor U8743 (N_8743,N_8096,N_8039);
nand U8744 (N_8744,N_8399,N_8469);
or U8745 (N_8745,N_8193,N_8230);
nand U8746 (N_8746,N_8002,N_8286);
or U8747 (N_8747,N_8188,N_8267);
or U8748 (N_8748,N_8149,N_8341);
or U8749 (N_8749,N_8382,N_8294);
or U8750 (N_8750,N_8450,N_8022);
xor U8751 (N_8751,N_8100,N_8016);
xor U8752 (N_8752,N_8332,N_8215);
xnor U8753 (N_8753,N_8129,N_8343);
or U8754 (N_8754,N_8431,N_8087);
nand U8755 (N_8755,N_8054,N_8397);
nor U8756 (N_8756,N_8261,N_8004);
and U8757 (N_8757,N_8135,N_8356);
xnor U8758 (N_8758,N_8082,N_8339);
nand U8759 (N_8759,N_8191,N_8063);
nor U8760 (N_8760,N_8300,N_8043);
and U8761 (N_8761,N_8291,N_8186);
and U8762 (N_8762,N_8002,N_8410);
and U8763 (N_8763,N_8476,N_8312);
and U8764 (N_8764,N_8460,N_8125);
xnor U8765 (N_8765,N_8160,N_8136);
nor U8766 (N_8766,N_8045,N_8406);
and U8767 (N_8767,N_8263,N_8306);
or U8768 (N_8768,N_8384,N_8366);
or U8769 (N_8769,N_8209,N_8007);
xnor U8770 (N_8770,N_8333,N_8158);
xnor U8771 (N_8771,N_8261,N_8131);
nand U8772 (N_8772,N_8202,N_8470);
and U8773 (N_8773,N_8040,N_8402);
and U8774 (N_8774,N_8488,N_8095);
and U8775 (N_8775,N_8440,N_8174);
nand U8776 (N_8776,N_8343,N_8323);
nor U8777 (N_8777,N_8330,N_8099);
or U8778 (N_8778,N_8457,N_8371);
and U8779 (N_8779,N_8197,N_8055);
nor U8780 (N_8780,N_8479,N_8348);
xor U8781 (N_8781,N_8319,N_8012);
nor U8782 (N_8782,N_8205,N_8166);
and U8783 (N_8783,N_8224,N_8148);
nor U8784 (N_8784,N_8147,N_8445);
and U8785 (N_8785,N_8428,N_8096);
nor U8786 (N_8786,N_8348,N_8347);
nand U8787 (N_8787,N_8010,N_8189);
or U8788 (N_8788,N_8019,N_8091);
xor U8789 (N_8789,N_8123,N_8313);
nor U8790 (N_8790,N_8435,N_8442);
and U8791 (N_8791,N_8260,N_8100);
nor U8792 (N_8792,N_8269,N_8263);
and U8793 (N_8793,N_8181,N_8070);
xnor U8794 (N_8794,N_8148,N_8290);
or U8795 (N_8795,N_8427,N_8029);
xor U8796 (N_8796,N_8401,N_8013);
nand U8797 (N_8797,N_8323,N_8167);
nor U8798 (N_8798,N_8445,N_8112);
and U8799 (N_8799,N_8430,N_8366);
and U8800 (N_8800,N_8231,N_8212);
xnor U8801 (N_8801,N_8297,N_8460);
nor U8802 (N_8802,N_8204,N_8047);
and U8803 (N_8803,N_8355,N_8456);
nor U8804 (N_8804,N_8238,N_8356);
xor U8805 (N_8805,N_8190,N_8262);
nor U8806 (N_8806,N_8434,N_8383);
nor U8807 (N_8807,N_8114,N_8343);
or U8808 (N_8808,N_8262,N_8312);
nand U8809 (N_8809,N_8106,N_8252);
and U8810 (N_8810,N_8392,N_8130);
and U8811 (N_8811,N_8148,N_8090);
or U8812 (N_8812,N_8387,N_8487);
xor U8813 (N_8813,N_8125,N_8273);
nand U8814 (N_8814,N_8399,N_8316);
or U8815 (N_8815,N_8432,N_8015);
and U8816 (N_8816,N_8392,N_8044);
nor U8817 (N_8817,N_8220,N_8029);
and U8818 (N_8818,N_8478,N_8466);
or U8819 (N_8819,N_8373,N_8121);
nor U8820 (N_8820,N_8414,N_8471);
and U8821 (N_8821,N_8426,N_8364);
nor U8822 (N_8822,N_8114,N_8366);
nand U8823 (N_8823,N_8169,N_8097);
or U8824 (N_8824,N_8197,N_8429);
xnor U8825 (N_8825,N_8317,N_8128);
xnor U8826 (N_8826,N_8390,N_8314);
nand U8827 (N_8827,N_8233,N_8046);
nor U8828 (N_8828,N_8461,N_8364);
nand U8829 (N_8829,N_8254,N_8386);
or U8830 (N_8830,N_8445,N_8284);
or U8831 (N_8831,N_8122,N_8460);
nor U8832 (N_8832,N_8494,N_8235);
nor U8833 (N_8833,N_8352,N_8007);
and U8834 (N_8834,N_8444,N_8300);
xnor U8835 (N_8835,N_8133,N_8255);
and U8836 (N_8836,N_8079,N_8398);
or U8837 (N_8837,N_8277,N_8242);
nand U8838 (N_8838,N_8323,N_8116);
nor U8839 (N_8839,N_8142,N_8166);
nor U8840 (N_8840,N_8282,N_8322);
nor U8841 (N_8841,N_8284,N_8094);
or U8842 (N_8842,N_8146,N_8078);
nand U8843 (N_8843,N_8059,N_8038);
nand U8844 (N_8844,N_8187,N_8008);
xor U8845 (N_8845,N_8215,N_8136);
xnor U8846 (N_8846,N_8109,N_8484);
xnor U8847 (N_8847,N_8242,N_8056);
or U8848 (N_8848,N_8227,N_8354);
xnor U8849 (N_8849,N_8138,N_8116);
nor U8850 (N_8850,N_8211,N_8115);
nand U8851 (N_8851,N_8434,N_8473);
or U8852 (N_8852,N_8331,N_8007);
nor U8853 (N_8853,N_8310,N_8268);
nand U8854 (N_8854,N_8286,N_8199);
and U8855 (N_8855,N_8139,N_8281);
nand U8856 (N_8856,N_8105,N_8033);
or U8857 (N_8857,N_8181,N_8261);
or U8858 (N_8858,N_8085,N_8080);
xnor U8859 (N_8859,N_8071,N_8024);
nand U8860 (N_8860,N_8484,N_8074);
nand U8861 (N_8861,N_8420,N_8011);
and U8862 (N_8862,N_8242,N_8251);
nand U8863 (N_8863,N_8291,N_8413);
and U8864 (N_8864,N_8342,N_8434);
nand U8865 (N_8865,N_8013,N_8169);
xnor U8866 (N_8866,N_8255,N_8078);
xor U8867 (N_8867,N_8391,N_8073);
nand U8868 (N_8868,N_8016,N_8238);
nor U8869 (N_8869,N_8356,N_8101);
and U8870 (N_8870,N_8076,N_8137);
nor U8871 (N_8871,N_8070,N_8454);
or U8872 (N_8872,N_8038,N_8029);
nor U8873 (N_8873,N_8284,N_8299);
xnor U8874 (N_8874,N_8196,N_8192);
xnor U8875 (N_8875,N_8492,N_8345);
or U8876 (N_8876,N_8454,N_8429);
nand U8877 (N_8877,N_8056,N_8293);
and U8878 (N_8878,N_8187,N_8004);
xor U8879 (N_8879,N_8384,N_8172);
xnor U8880 (N_8880,N_8080,N_8154);
nand U8881 (N_8881,N_8221,N_8491);
and U8882 (N_8882,N_8036,N_8317);
or U8883 (N_8883,N_8413,N_8455);
or U8884 (N_8884,N_8310,N_8474);
nor U8885 (N_8885,N_8183,N_8442);
and U8886 (N_8886,N_8298,N_8430);
xor U8887 (N_8887,N_8489,N_8336);
nor U8888 (N_8888,N_8114,N_8279);
nand U8889 (N_8889,N_8207,N_8487);
nand U8890 (N_8890,N_8374,N_8205);
nand U8891 (N_8891,N_8374,N_8488);
xnor U8892 (N_8892,N_8331,N_8144);
and U8893 (N_8893,N_8428,N_8460);
nand U8894 (N_8894,N_8371,N_8289);
or U8895 (N_8895,N_8466,N_8127);
and U8896 (N_8896,N_8059,N_8171);
and U8897 (N_8897,N_8492,N_8327);
nor U8898 (N_8898,N_8206,N_8062);
and U8899 (N_8899,N_8143,N_8229);
nor U8900 (N_8900,N_8226,N_8021);
nor U8901 (N_8901,N_8000,N_8077);
xor U8902 (N_8902,N_8197,N_8347);
xor U8903 (N_8903,N_8472,N_8467);
or U8904 (N_8904,N_8368,N_8326);
xnor U8905 (N_8905,N_8388,N_8108);
and U8906 (N_8906,N_8143,N_8427);
or U8907 (N_8907,N_8340,N_8000);
nand U8908 (N_8908,N_8007,N_8335);
or U8909 (N_8909,N_8281,N_8133);
xor U8910 (N_8910,N_8181,N_8117);
and U8911 (N_8911,N_8054,N_8052);
nor U8912 (N_8912,N_8084,N_8095);
nor U8913 (N_8913,N_8222,N_8179);
nor U8914 (N_8914,N_8180,N_8238);
nor U8915 (N_8915,N_8291,N_8194);
nor U8916 (N_8916,N_8335,N_8192);
or U8917 (N_8917,N_8432,N_8047);
nor U8918 (N_8918,N_8025,N_8468);
nand U8919 (N_8919,N_8349,N_8143);
and U8920 (N_8920,N_8342,N_8214);
xor U8921 (N_8921,N_8419,N_8367);
xnor U8922 (N_8922,N_8240,N_8440);
xor U8923 (N_8923,N_8279,N_8207);
nand U8924 (N_8924,N_8221,N_8368);
and U8925 (N_8925,N_8340,N_8368);
xnor U8926 (N_8926,N_8091,N_8295);
xor U8927 (N_8927,N_8049,N_8464);
or U8928 (N_8928,N_8201,N_8452);
and U8929 (N_8929,N_8248,N_8028);
or U8930 (N_8930,N_8447,N_8478);
nand U8931 (N_8931,N_8315,N_8101);
nor U8932 (N_8932,N_8419,N_8324);
nand U8933 (N_8933,N_8076,N_8244);
nor U8934 (N_8934,N_8004,N_8077);
or U8935 (N_8935,N_8471,N_8205);
xor U8936 (N_8936,N_8308,N_8354);
nand U8937 (N_8937,N_8154,N_8250);
xnor U8938 (N_8938,N_8359,N_8322);
nand U8939 (N_8939,N_8007,N_8407);
or U8940 (N_8940,N_8187,N_8463);
nand U8941 (N_8941,N_8001,N_8260);
nand U8942 (N_8942,N_8363,N_8272);
nor U8943 (N_8943,N_8204,N_8449);
nand U8944 (N_8944,N_8328,N_8250);
or U8945 (N_8945,N_8028,N_8157);
nand U8946 (N_8946,N_8313,N_8218);
and U8947 (N_8947,N_8405,N_8080);
xnor U8948 (N_8948,N_8373,N_8403);
or U8949 (N_8949,N_8146,N_8199);
nor U8950 (N_8950,N_8401,N_8323);
xor U8951 (N_8951,N_8112,N_8057);
xnor U8952 (N_8952,N_8104,N_8322);
xor U8953 (N_8953,N_8449,N_8443);
nand U8954 (N_8954,N_8116,N_8202);
nor U8955 (N_8955,N_8078,N_8170);
nor U8956 (N_8956,N_8454,N_8336);
xnor U8957 (N_8957,N_8302,N_8354);
or U8958 (N_8958,N_8314,N_8107);
nand U8959 (N_8959,N_8352,N_8457);
or U8960 (N_8960,N_8117,N_8314);
and U8961 (N_8961,N_8037,N_8008);
nor U8962 (N_8962,N_8043,N_8131);
or U8963 (N_8963,N_8297,N_8368);
nor U8964 (N_8964,N_8269,N_8369);
nor U8965 (N_8965,N_8385,N_8484);
or U8966 (N_8966,N_8037,N_8336);
and U8967 (N_8967,N_8466,N_8406);
or U8968 (N_8968,N_8177,N_8271);
xnor U8969 (N_8969,N_8064,N_8226);
and U8970 (N_8970,N_8215,N_8480);
or U8971 (N_8971,N_8434,N_8176);
nand U8972 (N_8972,N_8395,N_8387);
xnor U8973 (N_8973,N_8482,N_8290);
nor U8974 (N_8974,N_8123,N_8041);
or U8975 (N_8975,N_8150,N_8041);
nor U8976 (N_8976,N_8417,N_8054);
nor U8977 (N_8977,N_8336,N_8232);
nor U8978 (N_8978,N_8057,N_8048);
xnor U8979 (N_8979,N_8423,N_8257);
nand U8980 (N_8980,N_8179,N_8186);
xnor U8981 (N_8981,N_8019,N_8233);
or U8982 (N_8982,N_8008,N_8146);
xor U8983 (N_8983,N_8389,N_8177);
xnor U8984 (N_8984,N_8158,N_8419);
xor U8985 (N_8985,N_8360,N_8021);
or U8986 (N_8986,N_8077,N_8486);
nand U8987 (N_8987,N_8334,N_8205);
nand U8988 (N_8988,N_8087,N_8337);
or U8989 (N_8989,N_8434,N_8421);
or U8990 (N_8990,N_8331,N_8406);
and U8991 (N_8991,N_8225,N_8471);
nand U8992 (N_8992,N_8003,N_8220);
and U8993 (N_8993,N_8112,N_8437);
or U8994 (N_8994,N_8208,N_8058);
nor U8995 (N_8995,N_8022,N_8354);
or U8996 (N_8996,N_8294,N_8197);
and U8997 (N_8997,N_8273,N_8477);
xnor U8998 (N_8998,N_8420,N_8053);
nor U8999 (N_8999,N_8016,N_8256);
or U9000 (N_9000,N_8929,N_8616);
and U9001 (N_9001,N_8515,N_8601);
nor U9002 (N_9002,N_8844,N_8747);
and U9003 (N_9003,N_8773,N_8996);
nor U9004 (N_9004,N_8905,N_8592);
and U9005 (N_9005,N_8866,N_8578);
xnor U9006 (N_9006,N_8897,N_8672);
nand U9007 (N_9007,N_8914,N_8626);
or U9008 (N_9008,N_8508,N_8685);
xnor U9009 (N_9009,N_8661,N_8957);
nand U9010 (N_9010,N_8721,N_8554);
xnor U9011 (N_9011,N_8575,N_8528);
and U9012 (N_9012,N_8899,N_8795);
and U9013 (N_9013,N_8633,N_8945);
nor U9014 (N_9014,N_8551,N_8989);
or U9015 (N_9015,N_8739,N_8911);
or U9016 (N_9016,N_8703,N_8712);
nand U9017 (N_9017,N_8780,N_8698);
xor U9018 (N_9018,N_8558,N_8852);
nand U9019 (N_9019,N_8519,N_8790);
nor U9020 (N_9020,N_8699,N_8867);
xnor U9021 (N_9021,N_8850,N_8845);
and U9022 (N_9022,N_8752,N_8724);
and U9023 (N_9023,N_8847,N_8667);
or U9024 (N_9024,N_8700,N_8588);
nor U9025 (N_9025,N_8875,N_8798);
xnor U9026 (N_9026,N_8876,N_8716);
and U9027 (N_9027,N_8769,N_8599);
nand U9028 (N_9028,N_8561,N_8512);
and U9029 (N_9029,N_8978,N_8931);
nand U9030 (N_9030,N_8538,N_8808);
and U9031 (N_9031,N_8797,N_8745);
nor U9032 (N_9032,N_8654,N_8776);
or U9033 (N_9033,N_8630,N_8854);
and U9034 (N_9034,N_8803,N_8536);
nor U9035 (N_9035,N_8783,N_8546);
nand U9036 (N_9036,N_8657,N_8974);
or U9037 (N_9037,N_8816,N_8821);
or U9038 (N_9038,N_8734,N_8927);
nor U9039 (N_9039,N_8761,N_8740);
and U9040 (N_9040,N_8620,N_8925);
xnor U9041 (N_9041,N_8799,N_8506);
or U9042 (N_9042,N_8713,N_8617);
or U9043 (N_9043,N_8636,N_8812);
or U9044 (N_9044,N_8909,N_8873);
and U9045 (N_9045,N_8789,N_8757);
nand U9046 (N_9046,N_8582,N_8600);
nor U9047 (N_9047,N_8933,N_8590);
nand U9048 (N_9048,N_8612,N_8597);
and U9049 (N_9049,N_8665,N_8853);
or U9050 (N_9050,N_8809,N_8946);
or U9051 (N_9051,N_8969,N_8882);
nand U9052 (N_9052,N_8874,N_8842);
and U9053 (N_9053,N_8505,N_8580);
nand U9054 (N_9054,N_8901,N_8749);
and U9055 (N_9055,N_8823,N_8912);
nor U9056 (N_9056,N_8513,N_8678);
and U9057 (N_9057,N_8598,N_8942);
and U9058 (N_9058,N_8687,N_8555);
and U9059 (N_9059,N_8963,N_8841);
nor U9060 (N_9060,N_8501,N_8768);
nor U9061 (N_9061,N_8619,N_8744);
xor U9062 (N_9062,N_8675,N_8576);
and U9063 (N_9063,N_8604,N_8522);
and U9064 (N_9064,N_8581,N_8574);
or U9065 (N_9065,N_8503,N_8863);
and U9066 (N_9066,N_8613,N_8741);
and U9067 (N_9067,N_8688,N_8804);
or U9068 (N_9068,N_8562,N_8702);
xor U9069 (N_9069,N_8608,N_8651);
nand U9070 (N_9070,N_8788,N_8579);
nand U9071 (N_9071,N_8550,N_8738);
nor U9072 (N_9072,N_8791,N_8924);
and U9073 (N_9073,N_8877,N_8614);
xor U9074 (N_9074,N_8603,N_8885);
xnor U9075 (N_9075,N_8895,N_8966);
or U9076 (N_9076,N_8694,N_8908);
or U9077 (N_9077,N_8610,N_8627);
and U9078 (N_9078,N_8870,N_8697);
and U9079 (N_9079,N_8922,N_8971);
xnor U9080 (N_9080,N_8767,N_8746);
nand U9081 (N_9081,N_8583,N_8527);
or U9082 (N_9082,N_8709,N_8858);
nor U9083 (N_9083,N_8883,N_8953);
nand U9084 (N_9084,N_8671,N_8985);
nand U9085 (N_9085,N_8997,N_8572);
xor U9086 (N_9086,N_8585,N_8526);
or U9087 (N_9087,N_8851,N_8930);
nor U9088 (N_9088,N_8535,N_8939);
and U9089 (N_9089,N_8820,N_8892);
nor U9090 (N_9090,N_8846,N_8557);
nor U9091 (N_9091,N_8840,N_8765);
and U9092 (N_9092,N_8544,N_8862);
nor U9093 (N_9093,N_8750,N_8838);
nor U9094 (N_9094,N_8988,N_8920);
xor U9095 (N_9095,N_8631,N_8782);
or U9096 (N_9096,N_8577,N_8861);
and U9097 (N_9097,N_8753,N_8928);
or U9098 (N_9098,N_8891,N_8679);
nor U9099 (N_9099,N_8692,N_8518);
and U9100 (N_9100,N_8507,N_8943);
or U9101 (N_9101,N_8637,N_8806);
nor U9102 (N_9102,N_8715,N_8980);
nor U9103 (N_9103,N_8961,N_8542);
or U9104 (N_9104,N_8981,N_8775);
or U9105 (N_9105,N_8849,N_8817);
xnor U9106 (N_9106,N_8811,N_8570);
nand U9107 (N_9107,N_8986,N_8962);
and U9108 (N_9108,N_8832,N_8856);
xnor U9109 (N_9109,N_8548,N_8990);
and U9110 (N_9110,N_8831,N_8947);
xnor U9111 (N_9111,N_8514,N_8500);
or U9112 (N_9112,N_8830,N_8762);
nand U9113 (N_9113,N_8763,N_8565);
xor U9114 (N_9114,N_8733,N_8725);
xor U9115 (N_9115,N_8711,N_8984);
and U9116 (N_9116,N_8516,N_8975);
nand U9117 (N_9117,N_8859,N_8921);
and U9118 (N_9118,N_8607,N_8824);
nor U9119 (N_9119,N_8683,N_8991);
nor U9120 (N_9120,N_8737,N_8609);
nor U9121 (N_9121,N_8802,N_8728);
or U9122 (N_9122,N_8673,N_8926);
and U9123 (N_9123,N_8903,N_8556);
or U9124 (N_9124,N_8954,N_8605);
nor U9125 (N_9125,N_8913,N_8509);
xor U9126 (N_9126,N_8755,N_8960);
nand U9127 (N_9127,N_8999,N_8525);
xnor U9128 (N_9128,N_8646,N_8615);
nand U9129 (N_9129,N_8731,N_8635);
nand U9130 (N_9130,N_8800,N_8676);
or U9131 (N_9131,N_8693,N_8958);
or U9132 (N_9132,N_8801,N_8826);
nor U9133 (N_9133,N_8704,N_8602);
or U9134 (N_9134,N_8829,N_8611);
or U9135 (N_9135,N_8622,N_8568);
xnor U9136 (N_9136,N_8596,N_8815);
xnor U9137 (N_9137,N_8569,N_8906);
or U9138 (N_9138,N_8643,N_8900);
and U9139 (N_9139,N_8977,N_8793);
and U9140 (N_9140,N_8835,N_8560);
and U9141 (N_9141,N_8502,N_8720);
xnor U9142 (N_9142,N_8872,N_8543);
or U9143 (N_9143,N_8530,N_8904);
or U9144 (N_9144,N_8691,N_8878);
nor U9145 (N_9145,N_8726,N_8653);
nor U9146 (N_9146,N_8994,N_8855);
or U9147 (N_9147,N_8881,N_8666);
and U9148 (N_9148,N_8706,N_8591);
nand U9149 (N_9149,N_8656,N_8638);
xor U9150 (N_9150,N_8756,N_8718);
nand U9151 (N_9151,N_8774,N_8668);
nand U9152 (N_9152,N_8982,N_8649);
and U9153 (N_9153,N_8735,N_8549);
nor U9154 (N_9154,N_8955,N_8717);
xnor U9155 (N_9155,N_8584,N_8968);
xor U9156 (N_9156,N_8664,N_8690);
or U9157 (N_9157,N_8972,N_8524);
and U9158 (N_9158,N_8659,N_8836);
nand U9159 (N_9159,N_8595,N_8934);
xnor U9160 (N_9160,N_8952,N_8979);
nand U9161 (N_9161,N_8837,N_8537);
nor U9162 (N_9162,N_8677,N_8710);
and U9163 (N_9163,N_8825,N_8792);
nor U9164 (N_9164,N_8736,N_8540);
xnor U9165 (N_9165,N_8937,N_8794);
xnor U9166 (N_9166,N_8628,N_8786);
xnor U9167 (N_9167,N_8684,N_8917);
nor U9168 (N_9168,N_8839,N_8886);
and U9169 (N_9169,N_8587,N_8935);
and U9170 (N_9170,N_8686,N_8833);
nor U9171 (N_9171,N_8814,N_8669);
xor U9172 (N_9172,N_8510,N_8632);
nor U9173 (N_9173,N_8751,N_8564);
nand U9174 (N_9174,N_8967,N_8992);
xor U9175 (N_9175,N_8828,N_8534);
nand U9176 (N_9176,N_8674,N_8918);
nand U9177 (N_9177,N_8818,N_8566);
or U9178 (N_9178,N_8662,N_8796);
nand U9179 (N_9179,N_8998,N_8707);
xnor U9180 (N_9180,N_8964,N_8655);
and U9181 (N_9181,N_8663,N_8742);
and U9182 (N_9182,N_8951,N_8898);
or U9183 (N_9183,N_8644,N_8956);
and U9184 (N_9184,N_8893,N_8680);
nand U9185 (N_9185,N_8642,N_8722);
xnor U9186 (N_9186,N_8865,N_8950);
nand U9187 (N_9187,N_8995,N_8910);
xor U9188 (N_9188,N_8521,N_8880);
nand U9189 (N_9189,N_8645,N_8593);
and U9190 (N_9190,N_8827,N_8573);
nand U9191 (N_9191,N_8729,N_8748);
or U9192 (N_9192,N_8948,N_8552);
xnor U9193 (N_9193,N_8860,N_8689);
xor U9194 (N_9194,N_8708,N_8976);
nor U9195 (N_9195,N_8959,N_8520);
or U9196 (N_9196,N_8625,N_8727);
xor U9197 (N_9197,N_8848,N_8743);
and U9198 (N_9198,N_8884,N_8965);
nand U9199 (N_9199,N_8621,N_8517);
xnor U9200 (N_9200,N_8887,N_8531);
or U9201 (N_9201,N_8888,N_8681);
nor U9202 (N_9202,N_8639,N_8629);
xor U9203 (N_9203,N_8779,N_8936);
xnor U9204 (N_9204,N_8696,N_8871);
and U9205 (N_9205,N_8787,N_8719);
nor U9206 (N_9206,N_8973,N_8819);
and U9207 (N_9207,N_8894,N_8529);
or U9208 (N_9208,N_8764,N_8563);
and U9209 (N_9209,N_8647,N_8547);
nand U9210 (N_9210,N_8784,N_8983);
nor U9211 (N_9211,N_8705,N_8523);
nor U9212 (N_9212,N_8869,N_8810);
xnor U9213 (N_9213,N_8940,N_8941);
and U9214 (N_9214,N_8567,N_8532);
and U9215 (N_9215,N_8640,N_8559);
and U9216 (N_9216,N_8533,N_8915);
xor U9217 (N_9217,N_8511,N_8944);
xnor U9218 (N_9218,N_8539,N_8623);
and U9219 (N_9219,N_8777,N_8778);
xor U9220 (N_9220,N_8732,N_8759);
xor U9221 (N_9221,N_8770,N_8658);
nand U9222 (N_9222,N_8993,N_8868);
xor U9223 (N_9223,N_8923,N_8670);
xor U9224 (N_9224,N_8586,N_8864);
xor U9225 (N_9225,N_8772,N_8754);
or U9226 (N_9226,N_8822,N_8634);
nor U9227 (N_9227,N_8807,N_8834);
and U9228 (N_9228,N_8594,N_8541);
or U9229 (N_9229,N_8902,N_8545);
nand U9230 (N_9230,N_8896,N_8624);
and U9231 (N_9231,N_8813,N_8890);
nor U9232 (N_9232,N_8571,N_8701);
and U9233 (N_9233,N_8618,N_8589);
xor U9234 (N_9234,N_8650,N_8652);
nor U9235 (N_9235,N_8641,N_8758);
nand U9236 (N_9236,N_8907,N_8682);
nor U9237 (N_9237,N_8760,N_8879);
nor U9238 (N_9238,N_8723,N_8771);
or U9239 (N_9239,N_8660,N_8606);
and U9240 (N_9240,N_8805,N_8843);
nor U9241 (N_9241,N_8730,N_8714);
xnor U9242 (N_9242,N_8932,N_8648);
or U9243 (N_9243,N_8766,N_8785);
xor U9244 (N_9244,N_8504,N_8949);
or U9245 (N_9245,N_8916,N_8695);
or U9246 (N_9246,N_8889,N_8938);
and U9247 (N_9247,N_8987,N_8857);
nor U9248 (N_9248,N_8919,N_8970);
xor U9249 (N_9249,N_8553,N_8781);
xnor U9250 (N_9250,N_8697,N_8951);
nand U9251 (N_9251,N_8540,N_8780);
nand U9252 (N_9252,N_8734,N_8588);
nor U9253 (N_9253,N_8879,N_8506);
and U9254 (N_9254,N_8508,N_8806);
xor U9255 (N_9255,N_8885,N_8596);
nor U9256 (N_9256,N_8608,N_8500);
nand U9257 (N_9257,N_8715,N_8749);
nor U9258 (N_9258,N_8624,N_8648);
xnor U9259 (N_9259,N_8540,N_8931);
nor U9260 (N_9260,N_8942,N_8825);
nor U9261 (N_9261,N_8951,N_8517);
xnor U9262 (N_9262,N_8523,N_8952);
xnor U9263 (N_9263,N_8773,N_8822);
and U9264 (N_9264,N_8806,N_8618);
xor U9265 (N_9265,N_8903,N_8886);
and U9266 (N_9266,N_8791,N_8509);
xor U9267 (N_9267,N_8864,N_8873);
nand U9268 (N_9268,N_8659,N_8620);
and U9269 (N_9269,N_8952,N_8939);
and U9270 (N_9270,N_8862,N_8655);
and U9271 (N_9271,N_8708,N_8566);
nor U9272 (N_9272,N_8606,N_8506);
nor U9273 (N_9273,N_8567,N_8960);
xnor U9274 (N_9274,N_8518,N_8819);
nor U9275 (N_9275,N_8689,N_8975);
nand U9276 (N_9276,N_8850,N_8889);
and U9277 (N_9277,N_8894,N_8789);
xor U9278 (N_9278,N_8943,N_8814);
nand U9279 (N_9279,N_8796,N_8745);
nand U9280 (N_9280,N_8626,N_8848);
or U9281 (N_9281,N_8977,N_8590);
and U9282 (N_9282,N_8609,N_8579);
nand U9283 (N_9283,N_8584,N_8886);
or U9284 (N_9284,N_8779,N_8751);
nor U9285 (N_9285,N_8792,N_8848);
nor U9286 (N_9286,N_8720,N_8591);
or U9287 (N_9287,N_8572,N_8651);
xnor U9288 (N_9288,N_8715,N_8852);
nand U9289 (N_9289,N_8998,N_8727);
or U9290 (N_9290,N_8910,N_8641);
or U9291 (N_9291,N_8520,N_8956);
nand U9292 (N_9292,N_8855,N_8718);
nand U9293 (N_9293,N_8734,N_8505);
or U9294 (N_9294,N_8649,N_8733);
nor U9295 (N_9295,N_8603,N_8607);
nor U9296 (N_9296,N_8811,N_8914);
nor U9297 (N_9297,N_8651,N_8916);
xnor U9298 (N_9298,N_8842,N_8834);
and U9299 (N_9299,N_8829,N_8599);
nand U9300 (N_9300,N_8971,N_8932);
nor U9301 (N_9301,N_8537,N_8505);
nor U9302 (N_9302,N_8568,N_8598);
or U9303 (N_9303,N_8909,N_8975);
nand U9304 (N_9304,N_8646,N_8617);
nand U9305 (N_9305,N_8881,N_8648);
nand U9306 (N_9306,N_8885,N_8962);
nor U9307 (N_9307,N_8874,N_8658);
nand U9308 (N_9308,N_8898,N_8574);
and U9309 (N_9309,N_8730,N_8843);
nand U9310 (N_9310,N_8892,N_8723);
xnor U9311 (N_9311,N_8740,N_8544);
and U9312 (N_9312,N_8964,N_8882);
or U9313 (N_9313,N_8748,N_8675);
nand U9314 (N_9314,N_8622,N_8546);
nand U9315 (N_9315,N_8811,N_8794);
or U9316 (N_9316,N_8866,N_8536);
nor U9317 (N_9317,N_8944,N_8906);
nand U9318 (N_9318,N_8970,N_8750);
nand U9319 (N_9319,N_8690,N_8917);
and U9320 (N_9320,N_8960,N_8824);
xor U9321 (N_9321,N_8737,N_8891);
or U9322 (N_9322,N_8762,N_8633);
or U9323 (N_9323,N_8669,N_8936);
nand U9324 (N_9324,N_8586,N_8968);
xnor U9325 (N_9325,N_8903,N_8976);
or U9326 (N_9326,N_8663,N_8628);
or U9327 (N_9327,N_8908,N_8819);
xnor U9328 (N_9328,N_8841,N_8948);
nor U9329 (N_9329,N_8905,N_8662);
nand U9330 (N_9330,N_8936,N_8518);
nand U9331 (N_9331,N_8519,N_8913);
and U9332 (N_9332,N_8784,N_8751);
nor U9333 (N_9333,N_8615,N_8696);
nand U9334 (N_9334,N_8822,N_8823);
nor U9335 (N_9335,N_8671,N_8730);
nor U9336 (N_9336,N_8710,N_8748);
xor U9337 (N_9337,N_8708,N_8629);
nand U9338 (N_9338,N_8721,N_8818);
xnor U9339 (N_9339,N_8808,N_8791);
xor U9340 (N_9340,N_8928,N_8772);
nand U9341 (N_9341,N_8624,N_8994);
or U9342 (N_9342,N_8658,N_8979);
and U9343 (N_9343,N_8874,N_8975);
or U9344 (N_9344,N_8991,N_8523);
and U9345 (N_9345,N_8547,N_8680);
and U9346 (N_9346,N_8915,N_8674);
nor U9347 (N_9347,N_8819,N_8615);
xor U9348 (N_9348,N_8998,N_8802);
nor U9349 (N_9349,N_8957,N_8550);
nor U9350 (N_9350,N_8946,N_8518);
xor U9351 (N_9351,N_8992,N_8556);
xnor U9352 (N_9352,N_8663,N_8517);
or U9353 (N_9353,N_8849,N_8823);
and U9354 (N_9354,N_8619,N_8964);
and U9355 (N_9355,N_8593,N_8506);
or U9356 (N_9356,N_8818,N_8511);
or U9357 (N_9357,N_8678,N_8814);
xnor U9358 (N_9358,N_8576,N_8846);
xnor U9359 (N_9359,N_8957,N_8542);
nor U9360 (N_9360,N_8705,N_8885);
and U9361 (N_9361,N_8693,N_8942);
and U9362 (N_9362,N_8559,N_8695);
nor U9363 (N_9363,N_8747,N_8820);
nand U9364 (N_9364,N_8695,N_8595);
nand U9365 (N_9365,N_8783,N_8842);
and U9366 (N_9366,N_8731,N_8693);
xor U9367 (N_9367,N_8698,N_8655);
or U9368 (N_9368,N_8798,N_8773);
xnor U9369 (N_9369,N_8597,N_8721);
nand U9370 (N_9370,N_8506,N_8997);
or U9371 (N_9371,N_8919,N_8826);
or U9372 (N_9372,N_8754,N_8833);
and U9373 (N_9373,N_8663,N_8527);
and U9374 (N_9374,N_8909,N_8981);
nand U9375 (N_9375,N_8738,N_8585);
or U9376 (N_9376,N_8992,N_8783);
xnor U9377 (N_9377,N_8781,N_8535);
and U9378 (N_9378,N_8612,N_8894);
xor U9379 (N_9379,N_8804,N_8571);
nor U9380 (N_9380,N_8627,N_8588);
nor U9381 (N_9381,N_8565,N_8609);
nor U9382 (N_9382,N_8583,N_8569);
nor U9383 (N_9383,N_8992,N_8980);
nand U9384 (N_9384,N_8540,N_8968);
nand U9385 (N_9385,N_8895,N_8981);
or U9386 (N_9386,N_8914,N_8758);
and U9387 (N_9387,N_8706,N_8896);
xor U9388 (N_9388,N_8684,N_8870);
and U9389 (N_9389,N_8747,N_8604);
nand U9390 (N_9390,N_8544,N_8640);
or U9391 (N_9391,N_8838,N_8841);
nand U9392 (N_9392,N_8625,N_8578);
and U9393 (N_9393,N_8940,N_8649);
nor U9394 (N_9394,N_8877,N_8988);
nand U9395 (N_9395,N_8992,N_8605);
xor U9396 (N_9396,N_8632,N_8990);
and U9397 (N_9397,N_8753,N_8703);
and U9398 (N_9398,N_8881,N_8725);
nor U9399 (N_9399,N_8731,N_8755);
nor U9400 (N_9400,N_8924,N_8684);
nand U9401 (N_9401,N_8508,N_8719);
or U9402 (N_9402,N_8666,N_8740);
xor U9403 (N_9403,N_8597,N_8984);
xor U9404 (N_9404,N_8702,N_8660);
nand U9405 (N_9405,N_8524,N_8758);
or U9406 (N_9406,N_8564,N_8838);
nand U9407 (N_9407,N_8738,N_8568);
and U9408 (N_9408,N_8650,N_8716);
xnor U9409 (N_9409,N_8717,N_8740);
nand U9410 (N_9410,N_8583,N_8657);
xnor U9411 (N_9411,N_8614,N_8562);
nand U9412 (N_9412,N_8903,N_8888);
and U9413 (N_9413,N_8809,N_8908);
nor U9414 (N_9414,N_8711,N_8803);
xor U9415 (N_9415,N_8584,N_8563);
xnor U9416 (N_9416,N_8589,N_8848);
nand U9417 (N_9417,N_8929,N_8603);
nand U9418 (N_9418,N_8572,N_8887);
xor U9419 (N_9419,N_8721,N_8694);
nor U9420 (N_9420,N_8518,N_8587);
and U9421 (N_9421,N_8551,N_8880);
and U9422 (N_9422,N_8701,N_8604);
nand U9423 (N_9423,N_8732,N_8794);
xnor U9424 (N_9424,N_8809,N_8651);
or U9425 (N_9425,N_8593,N_8798);
or U9426 (N_9426,N_8954,N_8940);
nand U9427 (N_9427,N_8893,N_8983);
or U9428 (N_9428,N_8635,N_8507);
and U9429 (N_9429,N_8561,N_8526);
and U9430 (N_9430,N_8986,N_8872);
xnor U9431 (N_9431,N_8691,N_8573);
nand U9432 (N_9432,N_8978,N_8691);
xnor U9433 (N_9433,N_8534,N_8640);
nand U9434 (N_9434,N_8842,N_8938);
nor U9435 (N_9435,N_8784,N_8670);
and U9436 (N_9436,N_8847,N_8572);
nor U9437 (N_9437,N_8963,N_8834);
nand U9438 (N_9438,N_8536,N_8806);
nand U9439 (N_9439,N_8540,N_8641);
and U9440 (N_9440,N_8920,N_8650);
and U9441 (N_9441,N_8563,N_8915);
nor U9442 (N_9442,N_8702,N_8779);
nor U9443 (N_9443,N_8794,N_8918);
nor U9444 (N_9444,N_8534,N_8959);
xor U9445 (N_9445,N_8792,N_8772);
xor U9446 (N_9446,N_8741,N_8606);
nor U9447 (N_9447,N_8835,N_8918);
and U9448 (N_9448,N_8782,N_8761);
xor U9449 (N_9449,N_8885,N_8683);
xnor U9450 (N_9450,N_8556,N_8690);
or U9451 (N_9451,N_8566,N_8737);
nor U9452 (N_9452,N_8899,N_8637);
nor U9453 (N_9453,N_8969,N_8913);
or U9454 (N_9454,N_8924,N_8586);
nor U9455 (N_9455,N_8719,N_8832);
nor U9456 (N_9456,N_8841,N_8997);
nand U9457 (N_9457,N_8522,N_8819);
or U9458 (N_9458,N_8956,N_8871);
xor U9459 (N_9459,N_8517,N_8659);
nor U9460 (N_9460,N_8913,N_8539);
nand U9461 (N_9461,N_8872,N_8813);
xnor U9462 (N_9462,N_8948,N_8501);
xor U9463 (N_9463,N_8857,N_8583);
or U9464 (N_9464,N_8676,N_8828);
nand U9465 (N_9465,N_8890,N_8606);
nor U9466 (N_9466,N_8695,N_8706);
xor U9467 (N_9467,N_8971,N_8567);
nand U9468 (N_9468,N_8752,N_8735);
nor U9469 (N_9469,N_8636,N_8795);
and U9470 (N_9470,N_8526,N_8640);
nand U9471 (N_9471,N_8749,N_8815);
xnor U9472 (N_9472,N_8639,N_8567);
nor U9473 (N_9473,N_8669,N_8783);
or U9474 (N_9474,N_8787,N_8764);
nand U9475 (N_9475,N_8861,N_8889);
or U9476 (N_9476,N_8640,N_8616);
nor U9477 (N_9477,N_8797,N_8767);
or U9478 (N_9478,N_8584,N_8786);
nor U9479 (N_9479,N_8659,N_8599);
nand U9480 (N_9480,N_8584,N_8944);
xor U9481 (N_9481,N_8806,N_8950);
nand U9482 (N_9482,N_8684,N_8520);
nor U9483 (N_9483,N_8675,N_8701);
nand U9484 (N_9484,N_8923,N_8998);
and U9485 (N_9485,N_8745,N_8695);
nand U9486 (N_9486,N_8777,N_8608);
or U9487 (N_9487,N_8591,N_8785);
nand U9488 (N_9488,N_8878,N_8533);
or U9489 (N_9489,N_8524,N_8681);
or U9490 (N_9490,N_8613,N_8628);
nand U9491 (N_9491,N_8512,N_8647);
nor U9492 (N_9492,N_8945,N_8678);
or U9493 (N_9493,N_8740,N_8756);
xnor U9494 (N_9494,N_8574,N_8967);
and U9495 (N_9495,N_8737,N_8840);
and U9496 (N_9496,N_8575,N_8798);
xnor U9497 (N_9497,N_8603,N_8756);
xor U9498 (N_9498,N_8752,N_8837);
and U9499 (N_9499,N_8855,N_8687);
xnor U9500 (N_9500,N_9132,N_9027);
nor U9501 (N_9501,N_9367,N_9135);
or U9502 (N_9502,N_9481,N_9474);
and U9503 (N_9503,N_9304,N_9083);
and U9504 (N_9504,N_9137,N_9016);
and U9505 (N_9505,N_9188,N_9281);
or U9506 (N_9506,N_9176,N_9112);
nand U9507 (N_9507,N_9371,N_9216);
nor U9508 (N_9508,N_9380,N_9094);
nor U9509 (N_9509,N_9357,N_9331);
nor U9510 (N_9510,N_9164,N_9383);
and U9511 (N_9511,N_9082,N_9059);
or U9512 (N_9512,N_9321,N_9064);
nand U9513 (N_9513,N_9084,N_9235);
nor U9514 (N_9514,N_9442,N_9422);
nor U9515 (N_9515,N_9229,N_9043);
nor U9516 (N_9516,N_9469,N_9300);
and U9517 (N_9517,N_9323,N_9073);
nor U9518 (N_9518,N_9149,N_9453);
xor U9519 (N_9519,N_9126,N_9069);
and U9520 (N_9520,N_9490,N_9253);
or U9521 (N_9521,N_9412,N_9088);
nand U9522 (N_9522,N_9291,N_9463);
and U9523 (N_9523,N_9386,N_9033);
nand U9524 (N_9524,N_9413,N_9382);
xnor U9525 (N_9525,N_9293,N_9133);
and U9526 (N_9526,N_9496,N_9232);
and U9527 (N_9527,N_9202,N_9451);
and U9528 (N_9528,N_9390,N_9272);
or U9529 (N_9529,N_9241,N_9044);
and U9530 (N_9530,N_9335,N_9428);
xor U9531 (N_9531,N_9226,N_9207);
xnor U9532 (N_9532,N_9103,N_9010);
and U9533 (N_9533,N_9396,N_9454);
nand U9534 (N_9534,N_9223,N_9434);
nand U9535 (N_9535,N_9320,N_9247);
and U9536 (N_9536,N_9147,N_9263);
and U9537 (N_9537,N_9204,N_9373);
nand U9538 (N_9538,N_9265,N_9210);
and U9539 (N_9539,N_9445,N_9089);
xor U9540 (N_9540,N_9462,N_9366);
or U9541 (N_9541,N_9198,N_9250);
and U9542 (N_9542,N_9234,N_9101);
xor U9543 (N_9543,N_9286,N_9116);
nor U9544 (N_9544,N_9276,N_9174);
nand U9545 (N_9545,N_9206,N_9045);
xor U9546 (N_9546,N_9260,N_9123);
nand U9547 (N_9547,N_9004,N_9273);
xnor U9548 (N_9548,N_9346,N_9003);
nor U9549 (N_9549,N_9047,N_9499);
nand U9550 (N_9550,N_9085,N_9289);
or U9551 (N_9551,N_9026,N_9056);
and U9552 (N_9552,N_9402,N_9217);
nand U9553 (N_9553,N_9065,N_9169);
or U9554 (N_9554,N_9430,N_9388);
xor U9555 (N_9555,N_9340,N_9185);
and U9556 (N_9556,N_9268,N_9087);
and U9557 (N_9557,N_9114,N_9076);
or U9558 (N_9558,N_9072,N_9316);
nand U9559 (N_9559,N_9024,N_9061);
or U9560 (N_9560,N_9324,N_9154);
xnor U9561 (N_9561,N_9029,N_9378);
and U9562 (N_9562,N_9048,N_9138);
nor U9563 (N_9563,N_9427,N_9086);
nand U9564 (N_9564,N_9470,N_9429);
and U9565 (N_9565,N_9444,N_9098);
and U9566 (N_9566,N_9079,N_9192);
or U9567 (N_9567,N_9242,N_9280);
and U9568 (N_9568,N_9482,N_9199);
nand U9569 (N_9569,N_9256,N_9160);
nor U9570 (N_9570,N_9053,N_9450);
nor U9571 (N_9571,N_9347,N_9358);
and U9572 (N_9572,N_9473,N_9224);
or U9573 (N_9573,N_9446,N_9140);
or U9574 (N_9574,N_9233,N_9020);
or U9575 (N_9575,N_9177,N_9001);
xor U9576 (N_9576,N_9353,N_9109);
nand U9577 (N_9577,N_9134,N_9285);
nor U9578 (N_9578,N_9136,N_9077);
nor U9579 (N_9579,N_9165,N_9187);
nor U9580 (N_9580,N_9262,N_9104);
and U9581 (N_9581,N_9051,N_9354);
nor U9582 (N_9582,N_9404,N_9037);
xnor U9583 (N_9583,N_9414,N_9194);
xnor U9584 (N_9584,N_9131,N_9180);
nor U9585 (N_9585,N_9157,N_9257);
and U9586 (N_9586,N_9017,N_9456);
or U9587 (N_9587,N_9363,N_9119);
nand U9588 (N_9588,N_9186,N_9407);
xor U9589 (N_9589,N_9118,N_9162);
or U9590 (N_9590,N_9307,N_9211);
nor U9591 (N_9591,N_9193,N_9183);
and U9592 (N_9592,N_9067,N_9200);
xor U9593 (N_9593,N_9326,N_9028);
nand U9594 (N_9594,N_9460,N_9095);
or U9595 (N_9595,N_9240,N_9171);
xor U9596 (N_9596,N_9345,N_9405);
nand U9597 (N_9597,N_9019,N_9343);
nor U9598 (N_9598,N_9419,N_9365);
nor U9599 (N_9599,N_9415,N_9361);
or U9600 (N_9600,N_9317,N_9392);
xnor U9601 (N_9601,N_9143,N_9355);
xor U9602 (N_9602,N_9055,N_9452);
xnor U9603 (N_9603,N_9274,N_9230);
or U9604 (N_9604,N_9021,N_9175);
nand U9605 (N_9605,N_9398,N_9002);
nor U9606 (N_9606,N_9493,N_9009);
nand U9607 (N_9607,N_9290,N_9052);
or U9608 (N_9608,N_9106,N_9038);
nand U9609 (N_9609,N_9041,N_9036);
nand U9610 (N_9610,N_9387,N_9178);
nor U9611 (N_9611,N_9278,N_9468);
nor U9612 (N_9612,N_9379,N_9014);
nand U9613 (N_9613,N_9225,N_9128);
or U9614 (N_9614,N_9333,N_9284);
nand U9615 (N_9615,N_9151,N_9011);
xor U9616 (N_9616,N_9237,N_9385);
nor U9617 (N_9617,N_9023,N_9349);
and U9618 (N_9618,N_9254,N_9492);
nor U9619 (N_9619,N_9218,N_9125);
nand U9620 (N_9620,N_9092,N_9472);
and U9621 (N_9621,N_9189,N_9288);
nor U9622 (N_9622,N_9375,N_9214);
and U9623 (N_9623,N_9337,N_9102);
or U9624 (N_9624,N_9115,N_9483);
nand U9625 (N_9625,N_9364,N_9018);
and U9626 (N_9626,N_9042,N_9251);
nand U9627 (N_9627,N_9093,N_9461);
and U9628 (N_9628,N_9113,N_9190);
and U9629 (N_9629,N_9105,N_9117);
xnor U9630 (N_9630,N_9158,N_9050);
or U9631 (N_9631,N_9341,N_9054);
nand U9632 (N_9632,N_9130,N_9269);
nor U9633 (N_9633,N_9301,N_9080);
or U9634 (N_9634,N_9219,N_9334);
or U9635 (N_9635,N_9479,N_9252);
and U9636 (N_9636,N_9172,N_9437);
xor U9637 (N_9637,N_9184,N_9314);
nand U9638 (N_9638,N_9152,N_9370);
nor U9639 (N_9639,N_9022,N_9145);
and U9640 (N_9640,N_9275,N_9328);
and U9641 (N_9641,N_9374,N_9410);
or U9642 (N_9642,N_9155,N_9330);
or U9643 (N_9643,N_9248,N_9013);
or U9644 (N_9644,N_9139,N_9231);
nor U9645 (N_9645,N_9447,N_9220);
xnor U9646 (N_9646,N_9426,N_9197);
and U9647 (N_9647,N_9008,N_9279);
nand U9648 (N_9648,N_9005,N_9025);
xnor U9649 (N_9649,N_9303,N_9411);
nor U9650 (N_9650,N_9270,N_9391);
and U9651 (N_9651,N_9039,N_9403);
xnor U9652 (N_9652,N_9352,N_9196);
nand U9653 (N_9653,N_9074,N_9163);
or U9654 (N_9654,N_9167,N_9243);
nand U9655 (N_9655,N_9322,N_9369);
nand U9656 (N_9656,N_9277,N_9215);
or U9657 (N_9657,N_9350,N_9209);
nor U9658 (N_9658,N_9338,N_9150);
xor U9659 (N_9659,N_9146,N_9295);
or U9660 (N_9660,N_9271,N_9212);
nor U9661 (N_9661,N_9015,N_9127);
and U9662 (N_9662,N_9332,N_9318);
and U9663 (N_9663,N_9467,N_9305);
or U9664 (N_9664,N_9181,N_9401);
nand U9665 (N_9665,N_9191,N_9182);
nand U9666 (N_9666,N_9108,N_9457);
or U9667 (N_9667,N_9173,N_9393);
xor U9668 (N_9668,N_9298,N_9416);
nand U9669 (N_9669,N_9432,N_9144);
xor U9670 (N_9670,N_9249,N_9170);
or U9671 (N_9671,N_9439,N_9486);
nand U9672 (N_9672,N_9299,N_9431);
or U9673 (N_9673,N_9075,N_9438);
or U9674 (N_9674,N_9208,N_9030);
nor U9675 (N_9675,N_9423,N_9397);
and U9676 (N_9676,N_9466,N_9062);
or U9677 (N_9677,N_9068,N_9287);
nand U9678 (N_9678,N_9421,N_9394);
or U9679 (N_9679,N_9296,N_9081);
nor U9680 (N_9680,N_9267,N_9478);
nor U9681 (N_9681,N_9161,N_9484);
xnor U9682 (N_9682,N_9205,N_9032);
or U9683 (N_9683,N_9377,N_9046);
nand U9684 (N_9684,N_9099,N_9362);
nor U9685 (N_9685,N_9063,N_9325);
and U9686 (N_9686,N_9049,N_9477);
nor U9687 (N_9687,N_9078,N_9148);
or U9688 (N_9688,N_9344,N_9306);
xnor U9689 (N_9689,N_9376,N_9097);
or U9690 (N_9690,N_9259,N_9327);
or U9691 (N_9691,N_9142,N_9000);
nand U9692 (N_9692,N_9107,N_9329);
xnor U9693 (N_9693,N_9308,N_9266);
nand U9694 (N_9694,N_9395,N_9264);
or U9695 (N_9695,N_9141,N_9381);
xnor U9696 (N_9696,N_9491,N_9400);
nor U9697 (N_9697,N_9201,N_9096);
nand U9698 (N_9698,N_9441,N_9443);
or U9699 (N_9699,N_9006,N_9489);
nand U9700 (N_9700,N_9058,N_9417);
nor U9701 (N_9701,N_9283,N_9485);
xor U9702 (N_9702,N_9040,N_9384);
nand U9703 (N_9703,N_9228,N_9292);
nand U9704 (N_9704,N_9465,N_9071);
nand U9705 (N_9705,N_9449,N_9475);
nor U9706 (N_9706,N_9471,N_9239);
nor U9707 (N_9707,N_9348,N_9246);
nor U9708 (N_9708,N_9455,N_9418);
nand U9709 (N_9709,N_9480,N_9124);
xor U9710 (N_9710,N_9121,N_9339);
nor U9711 (N_9711,N_9227,N_9244);
or U9712 (N_9712,N_9459,N_9360);
or U9713 (N_9713,N_9035,N_9356);
or U9714 (N_9714,N_9195,N_9458);
nand U9715 (N_9715,N_9309,N_9159);
and U9716 (N_9716,N_9359,N_9255);
and U9717 (N_9717,N_9122,N_9448);
nor U9718 (N_9718,N_9312,N_9297);
nand U9719 (N_9719,N_9464,N_9066);
nand U9720 (N_9720,N_9236,N_9261);
xor U9721 (N_9721,N_9222,N_9319);
or U9722 (N_9722,N_9245,N_9409);
and U9723 (N_9723,N_9420,N_9258);
xnor U9724 (N_9724,N_9111,N_9436);
xnor U9725 (N_9725,N_9408,N_9315);
xnor U9726 (N_9726,N_9336,N_9221);
xnor U9727 (N_9727,N_9091,N_9498);
nor U9728 (N_9728,N_9487,N_9168);
nor U9729 (N_9729,N_9031,N_9342);
and U9730 (N_9730,N_9153,N_9090);
and U9731 (N_9731,N_9476,N_9012);
or U9732 (N_9732,N_9488,N_9433);
nand U9733 (N_9733,N_9497,N_9213);
or U9734 (N_9734,N_9120,N_9057);
or U9735 (N_9735,N_9070,N_9399);
nor U9736 (N_9736,N_9389,N_9313);
xor U9737 (N_9737,N_9282,N_9310);
nor U9738 (N_9738,N_9179,N_9435);
and U9739 (N_9739,N_9129,N_9425);
and U9740 (N_9740,N_9495,N_9351);
or U9741 (N_9741,N_9494,N_9034);
and U9742 (N_9742,N_9203,N_9311);
xnor U9743 (N_9743,N_9424,N_9166);
xnor U9744 (N_9744,N_9368,N_9406);
nor U9745 (N_9745,N_9007,N_9302);
or U9746 (N_9746,N_9238,N_9372);
or U9747 (N_9747,N_9060,N_9294);
or U9748 (N_9748,N_9100,N_9156);
nand U9749 (N_9749,N_9440,N_9110);
nand U9750 (N_9750,N_9020,N_9079);
xor U9751 (N_9751,N_9458,N_9117);
and U9752 (N_9752,N_9179,N_9001);
and U9753 (N_9753,N_9075,N_9264);
xor U9754 (N_9754,N_9039,N_9385);
or U9755 (N_9755,N_9206,N_9384);
nand U9756 (N_9756,N_9422,N_9285);
xor U9757 (N_9757,N_9139,N_9148);
or U9758 (N_9758,N_9135,N_9070);
or U9759 (N_9759,N_9056,N_9316);
nand U9760 (N_9760,N_9496,N_9296);
xor U9761 (N_9761,N_9347,N_9156);
nand U9762 (N_9762,N_9023,N_9108);
or U9763 (N_9763,N_9202,N_9420);
or U9764 (N_9764,N_9392,N_9148);
nand U9765 (N_9765,N_9130,N_9483);
xnor U9766 (N_9766,N_9170,N_9272);
nor U9767 (N_9767,N_9233,N_9107);
or U9768 (N_9768,N_9104,N_9031);
or U9769 (N_9769,N_9492,N_9051);
or U9770 (N_9770,N_9109,N_9391);
nand U9771 (N_9771,N_9272,N_9202);
nand U9772 (N_9772,N_9271,N_9379);
nor U9773 (N_9773,N_9250,N_9187);
and U9774 (N_9774,N_9293,N_9209);
or U9775 (N_9775,N_9095,N_9332);
and U9776 (N_9776,N_9010,N_9376);
or U9777 (N_9777,N_9383,N_9328);
xor U9778 (N_9778,N_9170,N_9151);
and U9779 (N_9779,N_9225,N_9330);
nor U9780 (N_9780,N_9139,N_9007);
nand U9781 (N_9781,N_9328,N_9123);
xor U9782 (N_9782,N_9229,N_9037);
nor U9783 (N_9783,N_9184,N_9084);
or U9784 (N_9784,N_9423,N_9086);
xor U9785 (N_9785,N_9139,N_9221);
or U9786 (N_9786,N_9256,N_9466);
nand U9787 (N_9787,N_9461,N_9020);
and U9788 (N_9788,N_9341,N_9019);
nand U9789 (N_9789,N_9342,N_9441);
nand U9790 (N_9790,N_9015,N_9002);
and U9791 (N_9791,N_9274,N_9418);
nand U9792 (N_9792,N_9143,N_9199);
xnor U9793 (N_9793,N_9129,N_9219);
nand U9794 (N_9794,N_9107,N_9001);
or U9795 (N_9795,N_9066,N_9193);
xnor U9796 (N_9796,N_9458,N_9351);
nor U9797 (N_9797,N_9251,N_9300);
or U9798 (N_9798,N_9432,N_9411);
or U9799 (N_9799,N_9191,N_9468);
and U9800 (N_9800,N_9120,N_9466);
and U9801 (N_9801,N_9437,N_9443);
and U9802 (N_9802,N_9397,N_9154);
and U9803 (N_9803,N_9375,N_9382);
and U9804 (N_9804,N_9099,N_9465);
and U9805 (N_9805,N_9212,N_9138);
xor U9806 (N_9806,N_9011,N_9383);
and U9807 (N_9807,N_9216,N_9229);
or U9808 (N_9808,N_9221,N_9403);
or U9809 (N_9809,N_9449,N_9058);
nand U9810 (N_9810,N_9390,N_9326);
xnor U9811 (N_9811,N_9433,N_9210);
or U9812 (N_9812,N_9228,N_9034);
xnor U9813 (N_9813,N_9274,N_9461);
or U9814 (N_9814,N_9170,N_9487);
and U9815 (N_9815,N_9216,N_9436);
nor U9816 (N_9816,N_9020,N_9040);
nor U9817 (N_9817,N_9274,N_9182);
nor U9818 (N_9818,N_9063,N_9361);
xnor U9819 (N_9819,N_9308,N_9401);
nand U9820 (N_9820,N_9093,N_9082);
and U9821 (N_9821,N_9355,N_9415);
or U9822 (N_9822,N_9412,N_9433);
xor U9823 (N_9823,N_9175,N_9231);
xnor U9824 (N_9824,N_9197,N_9339);
and U9825 (N_9825,N_9153,N_9471);
nand U9826 (N_9826,N_9284,N_9022);
xor U9827 (N_9827,N_9112,N_9213);
nor U9828 (N_9828,N_9325,N_9194);
nand U9829 (N_9829,N_9232,N_9231);
xor U9830 (N_9830,N_9171,N_9131);
or U9831 (N_9831,N_9445,N_9381);
or U9832 (N_9832,N_9246,N_9393);
nor U9833 (N_9833,N_9479,N_9204);
nor U9834 (N_9834,N_9453,N_9338);
nand U9835 (N_9835,N_9122,N_9043);
xnor U9836 (N_9836,N_9387,N_9362);
xor U9837 (N_9837,N_9238,N_9380);
nand U9838 (N_9838,N_9493,N_9164);
xor U9839 (N_9839,N_9266,N_9286);
nand U9840 (N_9840,N_9454,N_9174);
nand U9841 (N_9841,N_9385,N_9005);
nor U9842 (N_9842,N_9218,N_9026);
xor U9843 (N_9843,N_9320,N_9362);
or U9844 (N_9844,N_9370,N_9378);
xor U9845 (N_9845,N_9080,N_9195);
nor U9846 (N_9846,N_9446,N_9034);
nor U9847 (N_9847,N_9249,N_9338);
or U9848 (N_9848,N_9336,N_9423);
and U9849 (N_9849,N_9326,N_9004);
and U9850 (N_9850,N_9497,N_9326);
nand U9851 (N_9851,N_9098,N_9182);
and U9852 (N_9852,N_9132,N_9248);
and U9853 (N_9853,N_9215,N_9388);
nor U9854 (N_9854,N_9280,N_9126);
or U9855 (N_9855,N_9330,N_9470);
or U9856 (N_9856,N_9012,N_9043);
and U9857 (N_9857,N_9094,N_9119);
nor U9858 (N_9858,N_9135,N_9482);
nand U9859 (N_9859,N_9487,N_9176);
nand U9860 (N_9860,N_9007,N_9161);
nor U9861 (N_9861,N_9391,N_9060);
nand U9862 (N_9862,N_9256,N_9362);
nor U9863 (N_9863,N_9463,N_9485);
nand U9864 (N_9864,N_9470,N_9127);
nand U9865 (N_9865,N_9044,N_9290);
nand U9866 (N_9866,N_9367,N_9269);
xor U9867 (N_9867,N_9349,N_9403);
or U9868 (N_9868,N_9272,N_9214);
or U9869 (N_9869,N_9237,N_9009);
or U9870 (N_9870,N_9277,N_9037);
and U9871 (N_9871,N_9115,N_9256);
nor U9872 (N_9872,N_9462,N_9142);
nand U9873 (N_9873,N_9246,N_9408);
nand U9874 (N_9874,N_9185,N_9337);
and U9875 (N_9875,N_9498,N_9052);
nor U9876 (N_9876,N_9277,N_9208);
nor U9877 (N_9877,N_9255,N_9183);
and U9878 (N_9878,N_9470,N_9366);
nor U9879 (N_9879,N_9153,N_9110);
xor U9880 (N_9880,N_9373,N_9230);
xnor U9881 (N_9881,N_9022,N_9375);
nor U9882 (N_9882,N_9493,N_9154);
nand U9883 (N_9883,N_9292,N_9065);
and U9884 (N_9884,N_9371,N_9093);
xor U9885 (N_9885,N_9419,N_9372);
nor U9886 (N_9886,N_9383,N_9249);
nor U9887 (N_9887,N_9351,N_9420);
and U9888 (N_9888,N_9221,N_9219);
xor U9889 (N_9889,N_9060,N_9420);
or U9890 (N_9890,N_9493,N_9340);
nor U9891 (N_9891,N_9035,N_9073);
nand U9892 (N_9892,N_9488,N_9201);
nand U9893 (N_9893,N_9155,N_9486);
nor U9894 (N_9894,N_9408,N_9496);
and U9895 (N_9895,N_9474,N_9296);
and U9896 (N_9896,N_9365,N_9033);
nand U9897 (N_9897,N_9048,N_9118);
nand U9898 (N_9898,N_9145,N_9254);
nor U9899 (N_9899,N_9049,N_9423);
nand U9900 (N_9900,N_9270,N_9478);
or U9901 (N_9901,N_9375,N_9033);
nor U9902 (N_9902,N_9405,N_9063);
or U9903 (N_9903,N_9087,N_9006);
or U9904 (N_9904,N_9296,N_9158);
or U9905 (N_9905,N_9382,N_9363);
nand U9906 (N_9906,N_9255,N_9228);
nand U9907 (N_9907,N_9236,N_9298);
or U9908 (N_9908,N_9201,N_9471);
and U9909 (N_9909,N_9159,N_9345);
nor U9910 (N_9910,N_9374,N_9454);
and U9911 (N_9911,N_9203,N_9144);
and U9912 (N_9912,N_9066,N_9173);
nand U9913 (N_9913,N_9477,N_9087);
xor U9914 (N_9914,N_9416,N_9463);
or U9915 (N_9915,N_9409,N_9319);
nand U9916 (N_9916,N_9468,N_9059);
xor U9917 (N_9917,N_9463,N_9492);
nor U9918 (N_9918,N_9210,N_9001);
nor U9919 (N_9919,N_9461,N_9009);
nand U9920 (N_9920,N_9090,N_9023);
xor U9921 (N_9921,N_9385,N_9348);
or U9922 (N_9922,N_9141,N_9052);
nand U9923 (N_9923,N_9318,N_9437);
nand U9924 (N_9924,N_9337,N_9075);
and U9925 (N_9925,N_9236,N_9421);
or U9926 (N_9926,N_9180,N_9139);
xnor U9927 (N_9927,N_9341,N_9422);
xnor U9928 (N_9928,N_9471,N_9484);
xor U9929 (N_9929,N_9084,N_9079);
nor U9930 (N_9930,N_9020,N_9253);
or U9931 (N_9931,N_9408,N_9260);
nor U9932 (N_9932,N_9252,N_9089);
and U9933 (N_9933,N_9145,N_9291);
and U9934 (N_9934,N_9042,N_9328);
xor U9935 (N_9935,N_9359,N_9165);
xnor U9936 (N_9936,N_9098,N_9409);
nand U9937 (N_9937,N_9189,N_9401);
xor U9938 (N_9938,N_9382,N_9071);
nand U9939 (N_9939,N_9340,N_9103);
nand U9940 (N_9940,N_9499,N_9401);
xor U9941 (N_9941,N_9426,N_9126);
nor U9942 (N_9942,N_9085,N_9178);
xor U9943 (N_9943,N_9496,N_9275);
and U9944 (N_9944,N_9436,N_9135);
or U9945 (N_9945,N_9465,N_9267);
nand U9946 (N_9946,N_9406,N_9011);
nand U9947 (N_9947,N_9162,N_9469);
or U9948 (N_9948,N_9071,N_9236);
nor U9949 (N_9949,N_9070,N_9063);
nor U9950 (N_9950,N_9067,N_9336);
or U9951 (N_9951,N_9429,N_9436);
nor U9952 (N_9952,N_9277,N_9467);
and U9953 (N_9953,N_9004,N_9212);
or U9954 (N_9954,N_9318,N_9084);
xor U9955 (N_9955,N_9380,N_9090);
nor U9956 (N_9956,N_9275,N_9348);
nand U9957 (N_9957,N_9323,N_9076);
xor U9958 (N_9958,N_9040,N_9412);
and U9959 (N_9959,N_9283,N_9129);
nand U9960 (N_9960,N_9399,N_9302);
xor U9961 (N_9961,N_9337,N_9018);
nor U9962 (N_9962,N_9413,N_9321);
or U9963 (N_9963,N_9060,N_9454);
xnor U9964 (N_9964,N_9153,N_9449);
and U9965 (N_9965,N_9186,N_9237);
xnor U9966 (N_9966,N_9447,N_9007);
nand U9967 (N_9967,N_9082,N_9090);
xor U9968 (N_9968,N_9001,N_9329);
or U9969 (N_9969,N_9330,N_9291);
or U9970 (N_9970,N_9263,N_9171);
and U9971 (N_9971,N_9218,N_9336);
and U9972 (N_9972,N_9470,N_9167);
and U9973 (N_9973,N_9428,N_9267);
xnor U9974 (N_9974,N_9288,N_9492);
and U9975 (N_9975,N_9468,N_9256);
or U9976 (N_9976,N_9291,N_9499);
and U9977 (N_9977,N_9468,N_9280);
nand U9978 (N_9978,N_9181,N_9245);
or U9979 (N_9979,N_9082,N_9067);
nor U9980 (N_9980,N_9213,N_9313);
xnor U9981 (N_9981,N_9465,N_9254);
nand U9982 (N_9982,N_9400,N_9268);
or U9983 (N_9983,N_9492,N_9039);
or U9984 (N_9984,N_9370,N_9029);
nand U9985 (N_9985,N_9432,N_9460);
nor U9986 (N_9986,N_9130,N_9253);
or U9987 (N_9987,N_9255,N_9046);
and U9988 (N_9988,N_9440,N_9003);
and U9989 (N_9989,N_9158,N_9308);
nand U9990 (N_9990,N_9055,N_9469);
and U9991 (N_9991,N_9407,N_9176);
xor U9992 (N_9992,N_9207,N_9048);
nor U9993 (N_9993,N_9248,N_9019);
nand U9994 (N_9994,N_9337,N_9489);
and U9995 (N_9995,N_9396,N_9110);
and U9996 (N_9996,N_9175,N_9214);
xor U9997 (N_9997,N_9273,N_9117);
nor U9998 (N_9998,N_9072,N_9043);
or U9999 (N_9999,N_9157,N_9169);
or U10000 (N_10000,N_9811,N_9955);
nor U10001 (N_10001,N_9965,N_9897);
nor U10002 (N_10002,N_9888,N_9751);
nand U10003 (N_10003,N_9749,N_9741);
or U10004 (N_10004,N_9640,N_9845);
nand U10005 (N_10005,N_9916,N_9667);
or U10006 (N_10006,N_9657,N_9935);
xnor U10007 (N_10007,N_9670,N_9874);
nor U10008 (N_10008,N_9701,N_9911);
nor U10009 (N_10009,N_9621,N_9922);
nand U10010 (N_10010,N_9954,N_9642);
nand U10011 (N_10011,N_9934,N_9942);
xnor U10012 (N_10012,N_9585,N_9549);
nor U10013 (N_10013,N_9509,N_9702);
or U10014 (N_10014,N_9545,N_9791);
nand U10015 (N_10015,N_9986,N_9512);
nor U10016 (N_10016,N_9528,N_9913);
nor U10017 (N_10017,N_9792,N_9574);
xnor U10018 (N_10018,N_9758,N_9678);
nor U10019 (N_10019,N_9788,N_9501);
or U10020 (N_10020,N_9736,N_9764);
and U10021 (N_10021,N_9853,N_9674);
xnor U10022 (N_10022,N_9914,N_9515);
nor U10023 (N_10023,N_9931,N_9752);
nand U10024 (N_10024,N_9819,N_9695);
or U10025 (N_10025,N_9614,N_9601);
nor U10026 (N_10026,N_9735,N_9883);
nor U10027 (N_10027,N_9840,N_9534);
xnor U10028 (N_10028,N_9952,N_9587);
nand U10029 (N_10029,N_9664,N_9576);
nand U10030 (N_10030,N_9979,N_9682);
nor U10031 (N_10031,N_9724,N_9833);
or U10032 (N_10032,N_9918,N_9849);
nor U10033 (N_10033,N_9600,N_9960);
xor U10034 (N_10034,N_9685,N_9522);
nand U10035 (N_10035,N_9963,N_9806);
and U10036 (N_10036,N_9930,N_9786);
or U10037 (N_10037,N_9705,N_9727);
nand U10038 (N_10038,N_9933,N_9805);
and U10039 (N_10039,N_9915,N_9793);
or U10040 (N_10040,N_9799,N_9946);
nand U10041 (N_10041,N_9629,N_9696);
or U10042 (N_10042,N_9530,N_9503);
xor U10043 (N_10043,N_9939,N_9851);
or U10044 (N_10044,N_9693,N_9532);
and U10045 (N_10045,N_9603,N_9710);
xnor U10046 (N_10046,N_9834,N_9763);
and U10047 (N_10047,N_9892,N_9541);
xnor U10048 (N_10048,N_9923,N_9513);
nor U10049 (N_10049,N_9783,N_9956);
and U10050 (N_10050,N_9533,N_9761);
xor U10051 (N_10051,N_9854,N_9604);
or U10052 (N_10052,N_9520,N_9597);
nor U10053 (N_10053,N_9653,N_9618);
nand U10054 (N_10054,N_9818,N_9999);
xnor U10055 (N_10055,N_9737,N_9624);
xor U10056 (N_10056,N_9686,N_9975);
and U10057 (N_10057,N_9639,N_9721);
and U10058 (N_10058,N_9738,N_9658);
nor U10059 (N_10059,N_9912,N_9767);
nand U10060 (N_10060,N_9745,N_9970);
and U10061 (N_10061,N_9998,N_9755);
or U10062 (N_10062,N_9714,N_9824);
xor U10063 (N_10063,N_9976,N_9798);
or U10064 (N_10064,N_9715,N_9837);
nor U10065 (N_10065,N_9890,N_9571);
nor U10066 (N_10066,N_9771,N_9876);
and U10067 (N_10067,N_9739,N_9831);
nor U10068 (N_10068,N_9562,N_9548);
nand U10069 (N_10069,N_9542,N_9974);
xnor U10070 (N_10070,N_9700,N_9568);
xnor U10071 (N_10071,N_9929,N_9633);
nand U10072 (N_10072,N_9590,N_9531);
xor U10073 (N_10073,N_9523,N_9740);
xnor U10074 (N_10074,N_9846,N_9602);
xnor U10075 (N_10075,N_9830,N_9619);
and U10076 (N_10076,N_9926,N_9723);
nor U10077 (N_10077,N_9638,N_9612);
nor U10078 (N_10078,N_9644,N_9932);
nor U10079 (N_10079,N_9921,N_9869);
and U10080 (N_10080,N_9617,N_9865);
xnor U10081 (N_10081,N_9748,N_9953);
or U10082 (N_10082,N_9726,N_9820);
nor U10083 (N_10083,N_9732,N_9719);
nand U10084 (N_10084,N_9539,N_9637);
or U10085 (N_10085,N_9866,N_9803);
xnor U10086 (N_10086,N_9776,N_9850);
nand U10087 (N_10087,N_9627,N_9887);
nor U10088 (N_10088,N_9675,N_9990);
or U10089 (N_10089,N_9943,N_9867);
and U10090 (N_10090,N_9949,N_9995);
nor U10091 (N_10091,N_9836,N_9645);
xnor U10092 (N_10092,N_9649,N_9839);
or U10093 (N_10093,N_9907,N_9804);
or U10094 (N_10094,N_9647,N_9608);
nor U10095 (N_10095,N_9742,N_9518);
nand U10096 (N_10096,N_9927,N_9648);
and U10097 (N_10097,N_9673,N_9757);
nand U10098 (N_10098,N_9625,N_9779);
and U10099 (N_10099,N_9588,N_9586);
xor U10100 (N_10100,N_9691,N_9709);
or U10101 (N_10101,N_9519,N_9605);
xnor U10102 (N_10102,N_9725,N_9558);
or U10103 (N_10103,N_9797,N_9718);
xor U10104 (N_10104,N_9623,N_9594);
nand U10105 (N_10105,N_9844,N_9772);
or U10106 (N_10106,N_9967,N_9762);
nor U10107 (N_10107,N_9988,N_9951);
nand U10108 (N_10108,N_9669,N_9575);
nand U10109 (N_10109,N_9861,N_9795);
and U10110 (N_10110,N_9920,N_9977);
nor U10111 (N_10111,N_9832,N_9596);
xor U10112 (N_10112,N_9753,N_9941);
nand U10113 (N_10113,N_9620,N_9769);
and U10114 (N_10114,N_9713,N_9925);
xnor U10115 (N_10115,N_9504,N_9547);
and U10116 (N_10116,N_9868,N_9997);
nand U10117 (N_10117,N_9668,N_9690);
or U10118 (N_10118,N_9982,N_9734);
xnor U10119 (N_10119,N_9641,N_9842);
nand U10120 (N_10120,N_9599,N_9557);
or U10121 (N_10121,N_9651,N_9527);
and U10122 (N_10122,N_9628,N_9631);
nor U10123 (N_10123,N_9801,N_9632);
and U10124 (N_10124,N_9903,N_9630);
or U10125 (N_10125,N_9744,N_9774);
and U10126 (N_10126,N_9650,N_9511);
nor U10127 (N_10127,N_9958,N_9676);
nor U10128 (N_10128,N_9589,N_9577);
xor U10129 (N_10129,N_9692,N_9784);
nor U10130 (N_10130,N_9505,N_9882);
nor U10131 (N_10131,N_9560,N_9857);
or U10132 (N_10132,N_9679,N_9889);
or U10133 (N_10133,N_9698,N_9961);
xnor U10134 (N_10134,N_9665,N_9583);
or U10135 (N_10135,N_9873,N_9856);
nand U10136 (N_10136,N_9556,N_9993);
nand U10137 (N_10137,N_9722,N_9613);
and U10138 (N_10138,N_9828,N_9694);
nor U10139 (N_10139,N_9591,N_9570);
xor U10140 (N_10140,N_9609,N_9582);
or U10141 (N_10141,N_9768,N_9672);
or U10142 (N_10142,N_9863,N_9728);
and U10143 (N_10143,N_9708,N_9860);
nand U10144 (N_10144,N_9981,N_9848);
xnor U10145 (N_10145,N_9712,N_9978);
nor U10146 (N_10146,N_9947,N_9950);
nand U10147 (N_10147,N_9537,N_9517);
nand U10148 (N_10148,N_9671,N_9689);
or U10149 (N_10149,N_9838,N_9827);
nor U10150 (N_10150,N_9969,N_9510);
and U10151 (N_10151,N_9810,N_9743);
or U10152 (N_10152,N_9782,N_9823);
nand U10153 (N_10153,N_9855,N_9566);
nor U10154 (N_10154,N_9524,N_9720);
xnor U10155 (N_10155,N_9937,N_9652);
or U10156 (N_10156,N_9529,N_9636);
nor U10157 (N_10157,N_9746,N_9731);
nand U10158 (N_10158,N_9521,N_9826);
nand U10159 (N_10159,N_9886,N_9663);
nand U10160 (N_10160,N_9567,N_9654);
xor U10161 (N_10161,N_9500,N_9870);
and U10162 (N_10162,N_9778,N_9610);
nor U10163 (N_10163,N_9777,N_9852);
nand U10164 (N_10164,N_9569,N_9506);
nor U10165 (N_10165,N_9626,N_9536);
xor U10166 (N_10166,N_9980,N_9551);
or U10167 (N_10167,N_9919,N_9507);
nand U10168 (N_10168,N_9972,N_9716);
nand U10169 (N_10169,N_9660,N_9508);
or U10170 (N_10170,N_9688,N_9787);
nand U10171 (N_10171,N_9606,N_9822);
and U10172 (N_10172,N_9991,N_9815);
nand U10173 (N_10173,N_9879,N_9634);
or U10174 (N_10174,N_9659,N_9580);
nor U10175 (N_10175,N_9550,N_9878);
or U10176 (N_10176,N_9514,N_9858);
or U10177 (N_10177,N_9994,N_9516);
or U10178 (N_10178,N_9829,N_9871);
nor U10179 (N_10179,N_9584,N_9661);
or U10180 (N_10180,N_9785,N_9796);
or U10181 (N_10181,N_9781,N_9872);
nor U10182 (N_10182,N_9502,N_9891);
nor U10183 (N_10183,N_9902,N_9711);
or U10184 (N_10184,N_9687,N_9572);
nor U10185 (N_10185,N_9877,N_9561);
nor U10186 (N_10186,N_9984,N_9756);
nand U10187 (N_10187,N_9717,N_9807);
nand U10188 (N_10188,N_9707,N_9940);
or U10189 (N_10189,N_9611,N_9593);
and U10190 (N_10190,N_9973,N_9526);
nand U10191 (N_10191,N_9592,N_9885);
or U10192 (N_10192,N_9643,N_9884);
nand U10193 (N_10193,N_9821,N_9555);
xnor U10194 (N_10194,N_9924,N_9864);
xor U10195 (N_10195,N_9546,N_9598);
or U10196 (N_10196,N_9908,N_9765);
or U10197 (N_10197,N_9750,N_9730);
and U10198 (N_10198,N_9699,N_9813);
or U10199 (N_10199,N_9944,N_9662);
or U10200 (N_10200,N_9968,N_9563);
and U10201 (N_10201,N_9697,N_9917);
or U10202 (N_10202,N_9565,N_9538);
xnor U10203 (N_10203,N_9835,N_9646);
nand U10204 (N_10204,N_9894,N_9959);
nand U10205 (N_10205,N_9904,N_9880);
nand U10206 (N_10206,N_9780,N_9683);
nor U10207 (N_10207,N_9881,N_9936);
and U10208 (N_10208,N_9684,N_9616);
and U10209 (N_10209,N_9800,N_9847);
xor U10210 (N_10210,N_9760,N_9553);
xnor U10211 (N_10211,N_9747,N_9680);
nor U10212 (N_10212,N_9816,N_9809);
and U10213 (N_10213,N_9910,N_9622);
nor U10214 (N_10214,N_9901,N_9775);
or U10215 (N_10215,N_9789,N_9770);
nand U10216 (N_10216,N_9573,N_9773);
nor U10217 (N_10217,N_9544,N_9825);
and U10218 (N_10218,N_9906,N_9564);
nand U10219 (N_10219,N_9595,N_9759);
nand U10220 (N_10220,N_9859,N_9615);
xor U10221 (N_10221,N_9579,N_9703);
nor U10222 (N_10222,N_9655,N_9656);
and U10223 (N_10223,N_9554,N_9983);
nor U10224 (N_10224,N_9559,N_9729);
or U10225 (N_10225,N_9987,N_9896);
xor U10226 (N_10226,N_9843,N_9841);
or U10227 (N_10227,N_9812,N_9964);
nor U10228 (N_10228,N_9754,N_9971);
xor U10229 (N_10229,N_9543,N_9957);
xnor U10230 (N_10230,N_9681,N_9966);
or U10231 (N_10231,N_9794,N_9875);
or U10232 (N_10232,N_9900,N_9704);
and U10233 (N_10233,N_9895,N_9535);
and U10234 (N_10234,N_9992,N_9607);
or U10235 (N_10235,N_9578,N_9581);
and U10236 (N_10236,N_9733,N_9893);
and U10237 (N_10237,N_9814,N_9706);
nand U10238 (N_10238,N_9666,N_9938);
nand U10239 (N_10239,N_9905,N_9909);
xnor U10240 (N_10240,N_9928,N_9802);
xnor U10241 (N_10241,N_9808,N_9948);
nor U10242 (N_10242,N_9945,N_9862);
nor U10243 (N_10243,N_9525,N_9996);
nor U10244 (N_10244,N_9635,N_9766);
or U10245 (N_10245,N_9899,N_9790);
nor U10246 (N_10246,N_9962,N_9677);
nor U10247 (N_10247,N_9817,N_9989);
and U10248 (N_10248,N_9898,N_9985);
or U10249 (N_10249,N_9540,N_9552);
nor U10250 (N_10250,N_9882,N_9759);
nor U10251 (N_10251,N_9694,N_9831);
or U10252 (N_10252,N_9595,N_9617);
nand U10253 (N_10253,N_9546,N_9869);
or U10254 (N_10254,N_9550,N_9963);
xor U10255 (N_10255,N_9726,N_9714);
or U10256 (N_10256,N_9626,N_9811);
xor U10257 (N_10257,N_9835,N_9720);
nor U10258 (N_10258,N_9585,N_9735);
and U10259 (N_10259,N_9808,N_9784);
or U10260 (N_10260,N_9789,N_9925);
or U10261 (N_10261,N_9677,N_9555);
or U10262 (N_10262,N_9768,N_9962);
or U10263 (N_10263,N_9901,N_9740);
and U10264 (N_10264,N_9639,N_9808);
and U10265 (N_10265,N_9966,N_9876);
xnor U10266 (N_10266,N_9631,N_9854);
xor U10267 (N_10267,N_9693,N_9918);
nor U10268 (N_10268,N_9597,N_9799);
or U10269 (N_10269,N_9784,N_9673);
xnor U10270 (N_10270,N_9879,N_9554);
xor U10271 (N_10271,N_9839,N_9972);
nand U10272 (N_10272,N_9672,N_9716);
and U10273 (N_10273,N_9502,N_9625);
xor U10274 (N_10274,N_9903,N_9580);
nand U10275 (N_10275,N_9527,N_9773);
nor U10276 (N_10276,N_9579,N_9637);
and U10277 (N_10277,N_9805,N_9902);
or U10278 (N_10278,N_9721,N_9934);
xnor U10279 (N_10279,N_9861,N_9716);
xor U10280 (N_10280,N_9814,N_9695);
or U10281 (N_10281,N_9661,N_9793);
nor U10282 (N_10282,N_9924,N_9754);
xnor U10283 (N_10283,N_9646,N_9869);
nor U10284 (N_10284,N_9827,N_9789);
xnor U10285 (N_10285,N_9946,N_9768);
or U10286 (N_10286,N_9621,N_9842);
nor U10287 (N_10287,N_9989,N_9532);
xor U10288 (N_10288,N_9762,N_9612);
nand U10289 (N_10289,N_9626,N_9994);
or U10290 (N_10290,N_9999,N_9780);
and U10291 (N_10291,N_9729,N_9749);
or U10292 (N_10292,N_9728,N_9975);
and U10293 (N_10293,N_9834,N_9693);
xnor U10294 (N_10294,N_9629,N_9943);
and U10295 (N_10295,N_9803,N_9865);
and U10296 (N_10296,N_9695,N_9515);
nand U10297 (N_10297,N_9620,N_9990);
nand U10298 (N_10298,N_9773,N_9685);
nand U10299 (N_10299,N_9791,N_9763);
xor U10300 (N_10300,N_9922,N_9992);
nand U10301 (N_10301,N_9817,N_9598);
and U10302 (N_10302,N_9570,N_9562);
and U10303 (N_10303,N_9673,N_9563);
nand U10304 (N_10304,N_9991,N_9570);
or U10305 (N_10305,N_9803,N_9905);
nand U10306 (N_10306,N_9801,N_9661);
nor U10307 (N_10307,N_9803,N_9718);
and U10308 (N_10308,N_9995,N_9516);
or U10309 (N_10309,N_9586,N_9869);
and U10310 (N_10310,N_9507,N_9855);
and U10311 (N_10311,N_9978,N_9791);
and U10312 (N_10312,N_9955,N_9506);
nor U10313 (N_10313,N_9688,N_9559);
nand U10314 (N_10314,N_9501,N_9572);
or U10315 (N_10315,N_9903,N_9760);
nor U10316 (N_10316,N_9755,N_9737);
nor U10317 (N_10317,N_9895,N_9746);
nand U10318 (N_10318,N_9973,N_9697);
and U10319 (N_10319,N_9932,N_9517);
or U10320 (N_10320,N_9866,N_9751);
nand U10321 (N_10321,N_9513,N_9783);
nor U10322 (N_10322,N_9975,N_9734);
xor U10323 (N_10323,N_9836,N_9560);
nand U10324 (N_10324,N_9709,N_9520);
and U10325 (N_10325,N_9610,N_9942);
and U10326 (N_10326,N_9755,N_9620);
xnor U10327 (N_10327,N_9729,N_9983);
nor U10328 (N_10328,N_9877,N_9627);
nand U10329 (N_10329,N_9875,N_9692);
nor U10330 (N_10330,N_9926,N_9790);
or U10331 (N_10331,N_9994,N_9556);
xnor U10332 (N_10332,N_9705,N_9564);
and U10333 (N_10333,N_9815,N_9587);
nor U10334 (N_10334,N_9873,N_9859);
or U10335 (N_10335,N_9924,N_9759);
xnor U10336 (N_10336,N_9583,N_9760);
xnor U10337 (N_10337,N_9602,N_9567);
and U10338 (N_10338,N_9880,N_9696);
or U10339 (N_10339,N_9655,N_9949);
nor U10340 (N_10340,N_9823,N_9853);
xor U10341 (N_10341,N_9503,N_9555);
nand U10342 (N_10342,N_9905,N_9702);
nand U10343 (N_10343,N_9508,N_9679);
nand U10344 (N_10344,N_9663,N_9939);
or U10345 (N_10345,N_9545,N_9928);
or U10346 (N_10346,N_9921,N_9616);
nor U10347 (N_10347,N_9742,N_9832);
or U10348 (N_10348,N_9780,N_9945);
xor U10349 (N_10349,N_9789,N_9800);
nand U10350 (N_10350,N_9786,N_9833);
or U10351 (N_10351,N_9692,N_9504);
nand U10352 (N_10352,N_9685,N_9741);
nor U10353 (N_10353,N_9815,N_9532);
nand U10354 (N_10354,N_9894,N_9939);
nand U10355 (N_10355,N_9677,N_9804);
or U10356 (N_10356,N_9642,N_9546);
nand U10357 (N_10357,N_9600,N_9691);
nand U10358 (N_10358,N_9770,N_9638);
nand U10359 (N_10359,N_9562,N_9959);
nand U10360 (N_10360,N_9892,N_9984);
or U10361 (N_10361,N_9957,N_9883);
nand U10362 (N_10362,N_9721,N_9534);
and U10363 (N_10363,N_9529,N_9895);
nand U10364 (N_10364,N_9992,N_9616);
nand U10365 (N_10365,N_9709,N_9949);
xor U10366 (N_10366,N_9665,N_9798);
or U10367 (N_10367,N_9825,N_9514);
xnor U10368 (N_10368,N_9866,N_9728);
nand U10369 (N_10369,N_9679,N_9998);
xor U10370 (N_10370,N_9818,N_9572);
nor U10371 (N_10371,N_9870,N_9985);
xnor U10372 (N_10372,N_9700,N_9811);
and U10373 (N_10373,N_9504,N_9611);
and U10374 (N_10374,N_9552,N_9517);
nand U10375 (N_10375,N_9996,N_9947);
xnor U10376 (N_10376,N_9637,N_9805);
or U10377 (N_10377,N_9629,N_9746);
and U10378 (N_10378,N_9631,N_9860);
xnor U10379 (N_10379,N_9548,N_9843);
nand U10380 (N_10380,N_9509,N_9556);
xor U10381 (N_10381,N_9977,N_9779);
nand U10382 (N_10382,N_9718,N_9730);
nand U10383 (N_10383,N_9527,N_9932);
nor U10384 (N_10384,N_9844,N_9975);
xnor U10385 (N_10385,N_9711,N_9846);
nor U10386 (N_10386,N_9824,N_9936);
nand U10387 (N_10387,N_9543,N_9734);
and U10388 (N_10388,N_9530,N_9608);
and U10389 (N_10389,N_9859,N_9703);
and U10390 (N_10390,N_9971,N_9713);
or U10391 (N_10391,N_9705,N_9574);
or U10392 (N_10392,N_9644,N_9710);
xor U10393 (N_10393,N_9910,N_9558);
and U10394 (N_10394,N_9558,N_9736);
nor U10395 (N_10395,N_9748,N_9838);
xnor U10396 (N_10396,N_9669,N_9692);
or U10397 (N_10397,N_9628,N_9856);
nand U10398 (N_10398,N_9821,N_9540);
or U10399 (N_10399,N_9517,N_9673);
xnor U10400 (N_10400,N_9750,N_9514);
nand U10401 (N_10401,N_9661,N_9818);
and U10402 (N_10402,N_9845,N_9720);
nor U10403 (N_10403,N_9829,N_9663);
xor U10404 (N_10404,N_9988,N_9881);
nand U10405 (N_10405,N_9822,N_9524);
xor U10406 (N_10406,N_9510,N_9735);
nor U10407 (N_10407,N_9759,N_9572);
xnor U10408 (N_10408,N_9905,N_9822);
nand U10409 (N_10409,N_9853,N_9972);
nor U10410 (N_10410,N_9657,N_9675);
nor U10411 (N_10411,N_9723,N_9833);
xnor U10412 (N_10412,N_9981,N_9878);
nand U10413 (N_10413,N_9684,N_9621);
or U10414 (N_10414,N_9904,N_9858);
or U10415 (N_10415,N_9573,N_9872);
nor U10416 (N_10416,N_9539,N_9618);
and U10417 (N_10417,N_9958,N_9906);
nand U10418 (N_10418,N_9811,N_9510);
or U10419 (N_10419,N_9842,N_9957);
xor U10420 (N_10420,N_9990,N_9766);
and U10421 (N_10421,N_9995,N_9828);
and U10422 (N_10422,N_9734,N_9884);
or U10423 (N_10423,N_9800,N_9946);
and U10424 (N_10424,N_9983,N_9914);
nand U10425 (N_10425,N_9995,N_9740);
nand U10426 (N_10426,N_9598,N_9867);
xor U10427 (N_10427,N_9620,N_9751);
nand U10428 (N_10428,N_9868,N_9508);
nand U10429 (N_10429,N_9641,N_9785);
xor U10430 (N_10430,N_9754,N_9767);
and U10431 (N_10431,N_9703,N_9610);
xnor U10432 (N_10432,N_9594,N_9933);
xnor U10433 (N_10433,N_9578,N_9849);
nand U10434 (N_10434,N_9600,N_9588);
nor U10435 (N_10435,N_9914,N_9901);
xnor U10436 (N_10436,N_9647,N_9761);
and U10437 (N_10437,N_9956,N_9550);
xnor U10438 (N_10438,N_9516,N_9791);
or U10439 (N_10439,N_9766,N_9754);
nor U10440 (N_10440,N_9980,N_9694);
and U10441 (N_10441,N_9532,N_9831);
and U10442 (N_10442,N_9643,N_9765);
nor U10443 (N_10443,N_9670,N_9613);
or U10444 (N_10444,N_9940,N_9938);
and U10445 (N_10445,N_9845,N_9923);
nor U10446 (N_10446,N_9923,N_9591);
nor U10447 (N_10447,N_9769,N_9624);
nand U10448 (N_10448,N_9705,N_9724);
nand U10449 (N_10449,N_9655,N_9958);
nor U10450 (N_10450,N_9946,N_9896);
or U10451 (N_10451,N_9694,N_9674);
nor U10452 (N_10452,N_9738,N_9707);
xor U10453 (N_10453,N_9650,N_9704);
xor U10454 (N_10454,N_9826,N_9992);
or U10455 (N_10455,N_9981,N_9822);
xnor U10456 (N_10456,N_9807,N_9862);
or U10457 (N_10457,N_9773,N_9615);
nand U10458 (N_10458,N_9591,N_9836);
nor U10459 (N_10459,N_9939,N_9815);
nand U10460 (N_10460,N_9884,N_9589);
xnor U10461 (N_10461,N_9891,N_9544);
and U10462 (N_10462,N_9682,N_9626);
and U10463 (N_10463,N_9808,N_9655);
nand U10464 (N_10464,N_9749,N_9609);
xnor U10465 (N_10465,N_9829,N_9924);
and U10466 (N_10466,N_9612,N_9567);
nand U10467 (N_10467,N_9940,N_9876);
xor U10468 (N_10468,N_9728,N_9956);
xor U10469 (N_10469,N_9514,N_9898);
or U10470 (N_10470,N_9803,N_9560);
nor U10471 (N_10471,N_9844,N_9637);
and U10472 (N_10472,N_9801,N_9947);
and U10473 (N_10473,N_9879,N_9585);
nor U10474 (N_10474,N_9824,N_9840);
or U10475 (N_10475,N_9865,N_9604);
nor U10476 (N_10476,N_9525,N_9802);
xnor U10477 (N_10477,N_9735,N_9830);
nor U10478 (N_10478,N_9561,N_9554);
nand U10479 (N_10479,N_9764,N_9557);
nand U10480 (N_10480,N_9992,N_9744);
nor U10481 (N_10481,N_9934,N_9549);
nand U10482 (N_10482,N_9873,N_9614);
xor U10483 (N_10483,N_9695,N_9963);
and U10484 (N_10484,N_9554,N_9730);
xnor U10485 (N_10485,N_9609,N_9731);
nor U10486 (N_10486,N_9569,N_9668);
nand U10487 (N_10487,N_9621,N_9872);
xnor U10488 (N_10488,N_9952,N_9609);
or U10489 (N_10489,N_9547,N_9698);
xor U10490 (N_10490,N_9504,N_9592);
and U10491 (N_10491,N_9535,N_9656);
and U10492 (N_10492,N_9559,N_9856);
and U10493 (N_10493,N_9950,N_9631);
xnor U10494 (N_10494,N_9908,N_9813);
nand U10495 (N_10495,N_9934,N_9969);
and U10496 (N_10496,N_9744,N_9693);
nor U10497 (N_10497,N_9652,N_9731);
xor U10498 (N_10498,N_9920,N_9788);
xnor U10499 (N_10499,N_9911,N_9813);
nand U10500 (N_10500,N_10391,N_10365);
xor U10501 (N_10501,N_10285,N_10149);
and U10502 (N_10502,N_10091,N_10114);
nand U10503 (N_10503,N_10394,N_10331);
xor U10504 (N_10504,N_10369,N_10171);
nand U10505 (N_10505,N_10252,N_10282);
nor U10506 (N_10506,N_10487,N_10130);
or U10507 (N_10507,N_10320,N_10306);
and U10508 (N_10508,N_10408,N_10090);
and U10509 (N_10509,N_10303,N_10450);
and U10510 (N_10510,N_10406,N_10194);
or U10511 (N_10511,N_10108,N_10440);
nor U10512 (N_10512,N_10368,N_10126);
nand U10513 (N_10513,N_10099,N_10201);
and U10514 (N_10514,N_10447,N_10380);
xnor U10515 (N_10515,N_10170,N_10029);
xnor U10516 (N_10516,N_10475,N_10421);
nor U10517 (N_10517,N_10094,N_10093);
xnor U10518 (N_10518,N_10212,N_10121);
xnor U10519 (N_10519,N_10134,N_10033);
nand U10520 (N_10520,N_10426,N_10110);
or U10521 (N_10521,N_10492,N_10417);
nand U10522 (N_10522,N_10240,N_10418);
and U10523 (N_10523,N_10480,N_10259);
and U10524 (N_10524,N_10453,N_10224);
or U10525 (N_10525,N_10222,N_10221);
and U10526 (N_10526,N_10032,N_10296);
nand U10527 (N_10527,N_10403,N_10359);
and U10528 (N_10528,N_10428,N_10400);
xnor U10529 (N_10529,N_10174,N_10405);
and U10530 (N_10530,N_10345,N_10059);
or U10531 (N_10531,N_10207,N_10189);
xnor U10532 (N_10532,N_10096,N_10107);
nand U10533 (N_10533,N_10324,N_10077);
and U10534 (N_10534,N_10347,N_10197);
or U10535 (N_10535,N_10407,N_10471);
nand U10536 (N_10536,N_10274,N_10276);
xor U10537 (N_10537,N_10131,N_10390);
nor U10538 (N_10538,N_10192,N_10250);
nand U10539 (N_10539,N_10488,N_10435);
or U10540 (N_10540,N_10294,N_10227);
and U10541 (N_10541,N_10313,N_10305);
and U10542 (N_10542,N_10361,N_10045);
nor U10543 (N_10543,N_10177,N_10000);
and U10544 (N_10544,N_10422,N_10003);
nor U10545 (N_10545,N_10217,N_10157);
nor U10546 (N_10546,N_10106,N_10196);
xor U10547 (N_10547,N_10145,N_10036);
nand U10548 (N_10548,N_10218,N_10229);
or U10549 (N_10549,N_10481,N_10413);
nor U10550 (N_10550,N_10261,N_10051);
nand U10551 (N_10551,N_10060,N_10239);
and U10552 (N_10552,N_10312,N_10138);
xnor U10553 (N_10553,N_10163,N_10358);
and U10554 (N_10554,N_10014,N_10223);
and U10555 (N_10555,N_10025,N_10436);
or U10556 (N_10556,N_10019,N_10010);
and U10557 (N_10557,N_10451,N_10314);
and U10558 (N_10558,N_10087,N_10387);
and U10559 (N_10559,N_10100,N_10468);
nand U10560 (N_10560,N_10042,N_10429);
nor U10561 (N_10561,N_10437,N_10442);
and U10562 (N_10562,N_10484,N_10257);
and U10563 (N_10563,N_10439,N_10225);
and U10564 (N_10564,N_10434,N_10216);
nand U10565 (N_10565,N_10123,N_10198);
and U10566 (N_10566,N_10136,N_10186);
xor U10567 (N_10567,N_10490,N_10443);
or U10568 (N_10568,N_10243,N_10351);
or U10569 (N_10569,N_10376,N_10325);
xnor U10570 (N_10570,N_10375,N_10291);
or U10571 (N_10571,N_10307,N_10273);
and U10572 (N_10572,N_10022,N_10255);
nand U10573 (N_10573,N_10004,N_10290);
nor U10574 (N_10574,N_10175,N_10353);
nor U10575 (N_10575,N_10113,N_10330);
nor U10576 (N_10576,N_10258,N_10178);
and U10577 (N_10577,N_10184,N_10112);
and U10578 (N_10578,N_10328,N_10310);
nand U10579 (N_10579,N_10052,N_10159);
nor U10580 (N_10580,N_10317,N_10166);
and U10581 (N_10581,N_10072,N_10287);
and U10582 (N_10582,N_10071,N_10173);
xnor U10583 (N_10583,N_10251,N_10206);
nor U10584 (N_10584,N_10367,N_10129);
or U10585 (N_10585,N_10152,N_10338);
xnor U10586 (N_10586,N_10247,N_10244);
nand U10587 (N_10587,N_10141,N_10050);
and U10588 (N_10588,N_10479,N_10409);
xor U10589 (N_10589,N_10055,N_10315);
nand U10590 (N_10590,N_10081,N_10069);
nand U10591 (N_10591,N_10279,N_10280);
nand U10592 (N_10592,N_10378,N_10160);
nand U10593 (N_10593,N_10013,N_10464);
nor U10594 (N_10594,N_10371,N_10483);
nand U10595 (N_10595,N_10078,N_10278);
nand U10596 (N_10596,N_10073,N_10344);
xor U10597 (N_10597,N_10309,N_10458);
xnor U10598 (N_10598,N_10153,N_10154);
nor U10599 (N_10599,N_10410,N_10180);
or U10600 (N_10600,N_10482,N_10208);
and U10601 (N_10601,N_10203,N_10193);
nand U10602 (N_10602,N_10476,N_10116);
or U10603 (N_10603,N_10363,N_10293);
nor U10604 (N_10604,N_10339,N_10117);
or U10605 (N_10605,N_10412,N_10416);
xnor U10606 (N_10606,N_10238,N_10377);
nor U10607 (N_10607,N_10139,N_10355);
nor U10608 (N_10608,N_10231,N_10028);
nand U10609 (N_10609,N_10397,N_10039);
xnor U10610 (N_10610,N_10414,N_10334);
or U10611 (N_10611,N_10191,N_10137);
nand U10612 (N_10612,N_10088,N_10089);
or U10613 (N_10613,N_10146,N_10142);
nor U10614 (N_10614,N_10404,N_10342);
or U10615 (N_10615,N_10057,N_10024);
nand U10616 (N_10616,N_10386,N_10053);
or U10617 (N_10617,N_10272,N_10133);
nor U10618 (N_10618,N_10232,N_10213);
nor U10619 (N_10619,N_10172,N_10444);
xnor U10620 (N_10620,N_10185,N_10187);
nand U10621 (N_10621,N_10283,N_10302);
or U10622 (N_10622,N_10493,N_10496);
xor U10623 (N_10623,N_10462,N_10002);
or U10624 (N_10624,N_10248,N_10054);
and U10625 (N_10625,N_10125,N_10379);
nor U10626 (N_10626,N_10155,N_10456);
nand U10627 (N_10627,N_10449,N_10372);
nor U10628 (N_10628,N_10230,N_10277);
nor U10629 (N_10629,N_10056,N_10271);
nand U10630 (N_10630,N_10388,N_10040);
nand U10631 (N_10631,N_10498,N_10064);
nand U10632 (N_10632,N_10084,N_10043);
xor U10633 (N_10633,N_10327,N_10009);
or U10634 (N_10634,N_10253,N_10499);
nand U10635 (N_10635,N_10161,N_10241);
nor U10636 (N_10636,N_10284,N_10485);
xor U10637 (N_10637,N_10046,N_10012);
or U10638 (N_10638,N_10176,N_10066);
and U10639 (N_10639,N_10415,N_10340);
nor U10640 (N_10640,N_10433,N_10061);
or U10641 (N_10641,N_10219,N_10199);
or U10642 (N_10642,N_10168,N_10079);
and U10643 (N_10643,N_10289,N_10349);
and U10644 (N_10644,N_10140,N_10200);
or U10645 (N_10645,N_10119,N_10427);
and U10646 (N_10646,N_10103,N_10211);
or U10647 (N_10647,N_10058,N_10445);
or U10648 (N_10648,N_10395,N_10370);
or U10649 (N_10649,N_10396,N_10144);
and U10650 (N_10650,N_10105,N_10038);
nor U10651 (N_10651,N_10182,N_10463);
nor U10652 (N_10652,N_10065,N_10169);
nand U10653 (N_10653,N_10011,N_10156);
nor U10654 (N_10654,N_10164,N_10343);
and U10655 (N_10655,N_10150,N_10335);
nand U10656 (N_10656,N_10362,N_10333);
and U10657 (N_10657,N_10266,N_10190);
nand U10658 (N_10658,N_10457,N_10023);
nor U10659 (N_10659,N_10383,N_10357);
xor U10660 (N_10660,N_10044,N_10419);
and U10661 (N_10661,N_10472,N_10195);
xor U10662 (N_10662,N_10062,N_10018);
xnor U10663 (N_10663,N_10308,N_10301);
and U10664 (N_10664,N_10494,N_10234);
nor U10665 (N_10665,N_10026,N_10295);
nand U10666 (N_10666,N_10249,N_10006);
nand U10667 (N_10667,N_10326,N_10111);
or U10668 (N_10668,N_10461,N_10473);
and U10669 (N_10669,N_10497,N_10034);
nor U10670 (N_10670,N_10148,N_10109);
or U10671 (N_10671,N_10214,N_10392);
and U10672 (N_10672,N_10478,N_10297);
nor U10673 (N_10673,N_10348,N_10101);
xor U10674 (N_10674,N_10288,N_10082);
xnor U10675 (N_10675,N_10228,N_10489);
nand U10676 (N_10676,N_10318,N_10031);
nand U10677 (N_10677,N_10454,N_10102);
xnor U10678 (N_10678,N_10430,N_10128);
and U10679 (N_10679,N_10469,N_10350);
nor U10680 (N_10680,N_10346,N_10432);
and U10681 (N_10681,N_10448,N_10298);
xor U10682 (N_10682,N_10423,N_10292);
nor U10683 (N_10683,N_10337,N_10226);
nand U10684 (N_10684,N_10167,N_10215);
xor U10685 (N_10685,N_10381,N_10354);
or U10686 (N_10686,N_10083,N_10188);
nand U10687 (N_10687,N_10235,N_10086);
nand U10688 (N_10688,N_10049,N_10459);
and U10689 (N_10689,N_10095,N_10321);
nor U10690 (N_10690,N_10202,N_10068);
xor U10691 (N_10691,N_10486,N_10098);
nand U10692 (N_10692,N_10151,N_10341);
nor U10693 (N_10693,N_10070,N_10384);
nor U10694 (N_10694,N_10382,N_10097);
nand U10695 (N_10695,N_10332,N_10204);
and U10696 (N_10696,N_10460,N_10329);
nand U10697 (N_10697,N_10270,N_10067);
and U10698 (N_10698,N_10263,N_10275);
or U10699 (N_10699,N_10356,N_10027);
nand U10700 (N_10700,N_10389,N_10304);
nor U10701 (N_10701,N_10385,N_10063);
nand U10702 (N_10702,N_10402,N_10474);
or U10703 (N_10703,N_10020,N_10092);
and U10704 (N_10704,N_10179,N_10048);
or U10705 (N_10705,N_10477,N_10075);
nor U10706 (N_10706,N_10135,N_10037);
and U10707 (N_10707,N_10124,N_10336);
xnor U10708 (N_10708,N_10431,N_10021);
nor U10709 (N_10709,N_10183,N_10267);
xor U10710 (N_10710,N_10316,N_10364);
xor U10711 (N_10711,N_10264,N_10262);
and U10712 (N_10712,N_10254,N_10017);
and U10713 (N_10713,N_10047,N_10181);
xnor U10714 (N_10714,N_10319,N_10165);
or U10715 (N_10715,N_10205,N_10246);
nor U10716 (N_10716,N_10076,N_10373);
xnor U10717 (N_10717,N_10452,N_10132);
and U10718 (N_10718,N_10007,N_10322);
nand U10719 (N_10719,N_10115,N_10242);
and U10720 (N_10720,N_10074,N_10005);
nor U10721 (N_10721,N_10420,N_10424);
xnor U10722 (N_10722,N_10158,N_10220);
nor U10723 (N_10723,N_10122,N_10120);
and U10724 (N_10724,N_10237,N_10491);
and U10725 (N_10725,N_10008,N_10085);
nor U10726 (N_10726,N_10233,N_10104);
and U10727 (N_10727,N_10467,N_10015);
nand U10728 (N_10728,N_10300,N_10127);
xor U10729 (N_10729,N_10016,N_10236);
nor U10730 (N_10730,N_10210,N_10398);
and U10731 (N_10731,N_10209,N_10281);
and U10732 (N_10732,N_10366,N_10256);
xnor U10733 (N_10733,N_10323,N_10495);
nand U10734 (N_10734,N_10299,N_10466);
or U10735 (N_10735,N_10441,N_10041);
nand U10736 (N_10736,N_10268,N_10399);
xnor U10737 (N_10737,N_10360,N_10446);
nand U10738 (N_10738,N_10352,N_10245);
or U10739 (N_10739,N_10260,N_10118);
nand U10740 (N_10740,N_10455,N_10470);
nand U10741 (N_10741,N_10393,N_10269);
and U10742 (N_10742,N_10374,N_10030);
and U10743 (N_10743,N_10401,N_10465);
or U10744 (N_10744,N_10438,N_10162);
and U10745 (N_10745,N_10286,N_10001);
nor U10746 (N_10746,N_10265,N_10311);
nor U10747 (N_10747,N_10080,N_10147);
and U10748 (N_10748,N_10035,N_10411);
nor U10749 (N_10749,N_10425,N_10143);
or U10750 (N_10750,N_10248,N_10134);
and U10751 (N_10751,N_10071,N_10013);
nor U10752 (N_10752,N_10185,N_10425);
nor U10753 (N_10753,N_10255,N_10167);
nor U10754 (N_10754,N_10362,N_10375);
or U10755 (N_10755,N_10376,N_10463);
xnor U10756 (N_10756,N_10030,N_10012);
xnor U10757 (N_10757,N_10120,N_10170);
xor U10758 (N_10758,N_10217,N_10137);
xor U10759 (N_10759,N_10038,N_10253);
or U10760 (N_10760,N_10282,N_10231);
nand U10761 (N_10761,N_10264,N_10385);
and U10762 (N_10762,N_10162,N_10196);
nand U10763 (N_10763,N_10484,N_10226);
nand U10764 (N_10764,N_10346,N_10467);
nor U10765 (N_10765,N_10318,N_10095);
or U10766 (N_10766,N_10424,N_10283);
or U10767 (N_10767,N_10313,N_10278);
nand U10768 (N_10768,N_10166,N_10105);
nor U10769 (N_10769,N_10179,N_10199);
or U10770 (N_10770,N_10407,N_10161);
or U10771 (N_10771,N_10028,N_10201);
nand U10772 (N_10772,N_10429,N_10460);
and U10773 (N_10773,N_10041,N_10248);
nand U10774 (N_10774,N_10122,N_10448);
nand U10775 (N_10775,N_10083,N_10236);
and U10776 (N_10776,N_10150,N_10426);
or U10777 (N_10777,N_10475,N_10330);
nand U10778 (N_10778,N_10435,N_10153);
nor U10779 (N_10779,N_10048,N_10311);
nor U10780 (N_10780,N_10414,N_10083);
and U10781 (N_10781,N_10133,N_10480);
and U10782 (N_10782,N_10422,N_10149);
xor U10783 (N_10783,N_10277,N_10394);
or U10784 (N_10784,N_10215,N_10261);
or U10785 (N_10785,N_10427,N_10357);
nor U10786 (N_10786,N_10136,N_10086);
and U10787 (N_10787,N_10214,N_10047);
nand U10788 (N_10788,N_10196,N_10117);
or U10789 (N_10789,N_10181,N_10332);
nor U10790 (N_10790,N_10334,N_10496);
nor U10791 (N_10791,N_10495,N_10409);
or U10792 (N_10792,N_10058,N_10421);
and U10793 (N_10793,N_10370,N_10063);
or U10794 (N_10794,N_10207,N_10086);
nor U10795 (N_10795,N_10142,N_10137);
and U10796 (N_10796,N_10397,N_10049);
nor U10797 (N_10797,N_10001,N_10278);
and U10798 (N_10798,N_10085,N_10055);
nor U10799 (N_10799,N_10244,N_10331);
and U10800 (N_10800,N_10127,N_10460);
nor U10801 (N_10801,N_10385,N_10279);
xnor U10802 (N_10802,N_10497,N_10158);
nand U10803 (N_10803,N_10249,N_10039);
and U10804 (N_10804,N_10210,N_10273);
nand U10805 (N_10805,N_10417,N_10488);
xor U10806 (N_10806,N_10390,N_10047);
and U10807 (N_10807,N_10006,N_10175);
xor U10808 (N_10808,N_10039,N_10109);
nor U10809 (N_10809,N_10136,N_10468);
xnor U10810 (N_10810,N_10072,N_10198);
xor U10811 (N_10811,N_10236,N_10106);
nor U10812 (N_10812,N_10031,N_10005);
nand U10813 (N_10813,N_10333,N_10358);
or U10814 (N_10814,N_10343,N_10190);
and U10815 (N_10815,N_10127,N_10165);
nand U10816 (N_10816,N_10234,N_10245);
nand U10817 (N_10817,N_10045,N_10366);
and U10818 (N_10818,N_10427,N_10465);
or U10819 (N_10819,N_10180,N_10123);
and U10820 (N_10820,N_10242,N_10221);
and U10821 (N_10821,N_10120,N_10326);
nor U10822 (N_10822,N_10399,N_10198);
nand U10823 (N_10823,N_10131,N_10210);
and U10824 (N_10824,N_10368,N_10389);
nand U10825 (N_10825,N_10479,N_10477);
or U10826 (N_10826,N_10186,N_10266);
and U10827 (N_10827,N_10490,N_10004);
nor U10828 (N_10828,N_10491,N_10184);
and U10829 (N_10829,N_10268,N_10264);
nor U10830 (N_10830,N_10169,N_10146);
xor U10831 (N_10831,N_10357,N_10142);
and U10832 (N_10832,N_10294,N_10312);
nand U10833 (N_10833,N_10403,N_10098);
nand U10834 (N_10834,N_10373,N_10341);
nand U10835 (N_10835,N_10120,N_10430);
and U10836 (N_10836,N_10245,N_10177);
nand U10837 (N_10837,N_10309,N_10091);
nand U10838 (N_10838,N_10032,N_10479);
xor U10839 (N_10839,N_10380,N_10007);
or U10840 (N_10840,N_10266,N_10112);
nor U10841 (N_10841,N_10096,N_10486);
nand U10842 (N_10842,N_10175,N_10009);
nand U10843 (N_10843,N_10103,N_10312);
and U10844 (N_10844,N_10037,N_10149);
nor U10845 (N_10845,N_10045,N_10092);
xnor U10846 (N_10846,N_10302,N_10041);
nor U10847 (N_10847,N_10395,N_10181);
and U10848 (N_10848,N_10367,N_10207);
xnor U10849 (N_10849,N_10246,N_10404);
or U10850 (N_10850,N_10297,N_10053);
nor U10851 (N_10851,N_10385,N_10078);
or U10852 (N_10852,N_10076,N_10009);
and U10853 (N_10853,N_10267,N_10059);
xnor U10854 (N_10854,N_10162,N_10419);
nor U10855 (N_10855,N_10230,N_10169);
nor U10856 (N_10856,N_10072,N_10153);
nor U10857 (N_10857,N_10258,N_10265);
nor U10858 (N_10858,N_10396,N_10482);
nand U10859 (N_10859,N_10011,N_10460);
or U10860 (N_10860,N_10017,N_10158);
nand U10861 (N_10861,N_10059,N_10470);
nor U10862 (N_10862,N_10436,N_10375);
xnor U10863 (N_10863,N_10152,N_10101);
and U10864 (N_10864,N_10395,N_10064);
and U10865 (N_10865,N_10343,N_10116);
and U10866 (N_10866,N_10278,N_10132);
xnor U10867 (N_10867,N_10183,N_10027);
nor U10868 (N_10868,N_10268,N_10183);
xor U10869 (N_10869,N_10461,N_10053);
or U10870 (N_10870,N_10370,N_10139);
nand U10871 (N_10871,N_10397,N_10151);
or U10872 (N_10872,N_10226,N_10051);
xor U10873 (N_10873,N_10303,N_10330);
xor U10874 (N_10874,N_10226,N_10208);
xnor U10875 (N_10875,N_10281,N_10117);
or U10876 (N_10876,N_10183,N_10460);
nor U10877 (N_10877,N_10330,N_10051);
nand U10878 (N_10878,N_10103,N_10170);
or U10879 (N_10879,N_10110,N_10231);
xnor U10880 (N_10880,N_10270,N_10169);
or U10881 (N_10881,N_10044,N_10346);
and U10882 (N_10882,N_10268,N_10178);
or U10883 (N_10883,N_10316,N_10106);
xnor U10884 (N_10884,N_10036,N_10169);
nor U10885 (N_10885,N_10144,N_10047);
nand U10886 (N_10886,N_10407,N_10455);
nor U10887 (N_10887,N_10259,N_10083);
or U10888 (N_10888,N_10406,N_10056);
and U10889 (N_10889,N_10459,N_10117);
xnor U10890 (N_10890,N_10264,N_10152);
or U10891 (N_10891,N_10192,N_10214);
nand U10892 (N_10892,N_10123,N_10007);
nand U10893 (N_10893,N_10208,N_10138);
nand U10894 (N_10894,N_10275,N_10495);
nand U10895 (N_10895,N_10206,N_10372);
xor U10896 (N_10896,N_10303,N_10135);
xor U10897 (N_10897,N_10358,N_10061);
and U10898 (N_10898,N_10375,N_10366);
xor U10899 (N_10899,N_10028,N_10430);
nor U10900 (N_10900,N_10402,N_10317);
nor U10901 (N_10901,N_10079,N_10074);
nand U10902 (N_10902,N_10416,N_10472);
xor U10903 (N_10903,N_10028,N_10194);
and U10904 (N_10904,N_10149,N_10116);
and U10905 (N_10905,N_10114,N_10293);
nor U10906 (N_10906,N_10348,N_10499);
and U10907 (N_10907,N_10361,N_10068);
nor U10908 (N_10908,N_10360,N_10277);
nand U10909 (N_10909,N_10217,N_10031);
nand U10910 (N_10910,N_10140,N_10416);
nand U10911 (N_10911,N_10420,N_10011);
or U10912 (N_10912,N_10085,N_10176);
or U10913 (N_10913,N_10399,N_10248);
and U10914 (N_10914,N_10047,N_10224);
xor U10915 (N_10915,N_10068,N_10079);
xor U10916 (N_10916,N_10278,N_10341);
nor U10917 (N_10917,N_10168,N_10403);
xnor U10918 (N_10918,N_10383,N_10143);
or U10919 (N_10919,N_10130,N_10341);
xor U10920 (N_10920,N_10069,N_10272);
or U10921 (N_10921,N_10003,N_10310);
nand U10922 (N_10922,N_10328,N_10002);
xnor U10923 (N_10923,N_10224,N_10360);
and U10924 (N_10924,N_10383,N_10486);
xnor U10925 (N_10925,N_10067,N_10210);
and U10926 (N_10926,N_10320,N_10281);
and U10927 (N_10927,N_10212,N_10036);
nand U10928 (N_10928,N_10112,N_10067);
xor U10929 (N_10929,N_10251,N_10428);
and U10930 (N_10930,N_10182,N_10366);
nor U10931 (N_10931,N_10150,N_10014);
and U10932 (N_10932,N_10342,N_10230);
and U10933 (N_10933,N_10173,N_10426);
xnor U10934 (N_10934,N_10444,N_10378);
and U10935 (N_10935,N_10338,N_10412);
and U10936 (N_10936,N_10190,N_10214);
nor U10937 (N_10937,N_10170,N_10469);
and U10938 (N_10938,N_10021,N_10294);
or U10939 (N_10939,N_10199,N_10370);
nor U10940 (N_10940,N_10163,N_10455);
nand U10941 (N_10941,N_10111,N_10419);
and U10942 (N_10942,N_10254,N_10323);
nor U10943 (N_10943,N_10407,N_10246);
and U10944 (N_10944,N_10208,N_10191);
nand U10945 (N_10945,N_10324,N_10032);
xor U10946 (N_10946,N_10433,N_10130);
nor U10947 (N_10947,N_10119,N_10313);
and U10948 (N_10948,N_10386,N_10283);
and U10949 (N_10949,N_10043,N_10377);
xnor U10950 (N_10950,N_10417,N_10370);
xor U10951 (N_10951,N_10185,N_10475);
nor U10952 (N_10952,N_10243,N_10327);
nor U10953 (N_10953,N_10352,N_10192);
or U10954 (N_10954,N_10489,N_10427);
or U10955 (N_10955,N_10159,N_10056);
nor U10956 (N_10956,N_10237,N_10016);
nor U10957 (N_10957,N_10038,N_10090);
and U10958 (N_10958,N_10088,N_10036);
xor U10959 (N_10959,N_10481,N_10393);
or U10960 (N_10960,N_10133,N_10048);
or U10961 (N_10961,N_10086,N_10309);
xnor U10962 (N_10962,N_10498,N_10134);
nor U10963 (N_10963,N_10387,N_10256);
xnor U10964 (N_10964,N_10291,N_10398);
or U10965 (N_10965,N_10453,N_10073);
and U10966 (N_10966,N_10289,N_10330);
and U10967 (N_10967,N_10342,N_10033);
nor U10968 (N_10968,N_10031,N_10238);
nand U10969 (N_10969,N_10492,N_10352);
nand U10970 (N_10970,N_10422,N_10466);
nand U10971 (N_10971,N_10457,N_10455);
nor U10972 (N_10972,N_10114,N_10050);
and U10973 (N_10973,N_10131,N_10473);
and U10974 (N_10974,N_10392,N_10201);
or U10975 (N_10975,N_10010,N_10119);
nand U10976 (N_10976,N_10356,N_10089);
nand U10977 (N_10977,N_10014,N_10347);
xor U10978 (N_10978,N_10146,N_10456);
nand U10979 (N_10979,N_10178,N_10193);
nand U10980 (N_10980,N_10323,N_10386);
nand U10981 (N_10981,N_10334,N_10069);
nor U10982 (N_10982,N_10047,N_10442);
or U10983 (N_10983,N_10475,N_10391);
nor U10984 (N_10984,N_10111,N_10280);
or U10985 (N_10985,N_10318,N_10199);
nor U10986 (N_10986,N_10270,N_10444);
nand U10987 (N_10987,N_10375,N_10117);
and U10988 (N_10988,N_10079,N_10003);
xor U10989 (N_10989,N_10177,N_10450);
nor U10990 (N_10990,N_10004,N_10439);
xor U10991 (N_10991,N_10118,N_10043);
or U10992 (N_10992,N_10266,N_10004);
and U10993 (N_10993,N_10155,N_10198);
nor U10994 (N_10994,N_10472,N_10123);
nand U10995 (N_10995,N_10155,N_10165);
nor U10996 (N_10996,N_10462,N_10387);
or U10997 (N_10997,N_10439,N_10269);
and U10998 (N_10998,N_10162,N_10133);
or U10999 (N_10999,N_10337,N_10400);
xnor U11000 (N_11000,N_10842,N_10509);
xnor U11001 (N_11001,N_10845,N_10899);
and U11002 (N_11002,N_10572,N_10979);
or U11003 (N_11003,N_10598,N_10906);
or U11004 (N_11004,N_10583,N_10679);
xnor U11005 (N_11005,N_10763,N_10794);
nand U11006 (N_11006,N_10862,N_10970);
or U11007 (N_11007,N_10852,N_10742);
or U11008 (N_11008,N_10769,N_10761);
xor U11009 (N_11009,N_10692,N_10615);
nand U11010 (N_11010,N_10659,N_10735);
and U11011 (N_11011,N_10560,N_10614);
nand U11012 (N_11012,N_10975,N_10526);
nand U11013 (N_11013,N_10789,N_10684);
or U11014 (N_11014,N_10767,N_10516);
and U11015 (N_11015,N_10506,N_10762);
and U11016 (N_11016,N_10559,N_10619);
nor U11017 (N_11017,N_10947,N_10775);
and U11018 (N_11018,N_10715,N_10960);
nor U11019 (N_11019,N_10942,N_10677);
nand U11020 (N_11020,N_10869,N_10626);
nand U11021 (N_11021,N_10901,N_10771);
xor U11022 (N_11022,N_10669,N_10853);
or U11023 (N_11023,N_10611,N_10877);
nand U11024 (N_11024,N_10688,N_10965);
and U11025 (N_11025,N_10702,N_10804);
or U11026 (N_11026,N_10689,N_10604);
xor U11027 (N_11027,N_10905,N_10579);
nand U11028 (N_11028,N_10838,N_10718);
nor U11029 (N_11029,N_10534,N_10897);
nor U11030 (N_11030,N_10703,N_10825);
xor U11031 (N_11031,N_10592,N_10632);
or U11032 (N_11032,N_10759,N_10800);
or U11033 (N_11033,N_10881,N_10891);
xor U11034 (N_11034,N_10671,N_10824);
or U11035 (N_11035,N_10991,N_10983);
or U11036 (N_11036,N_10541,N_10883);
or U11037 (N_11037,N_10680,N_10778);
nand U11038 (N_11038,N_10706,N_10610);
or U11039 (N_11039,N_10922,N_10525);
and U11040 (N_11040,N_10638,N_10840);
or U11041 (N_11041,N_10666,N_10907);
or U11042 (N_11042,N_10751,N_10788);
and U11043 (N_11043,N_10873,N_10744);
nor U11044 (N_11044,N_10773,N_10774);
and U11045 (N_11045,N_10756,N_10934);
xor U11046 (N_11046,N_10936,N_10507);
or U11047 (N_11047,N_10726,N_10729);
or U11048 (N_11048,N_10961,N_10861);
and U11049 (N_11049,N_10962,N_10605);
or U11050 (N_11050,N_10530,N_10843);
and U11051 (N_11051,N_10536,N_10567);
nor U11052 (N_11052,N_10935,N_10665);
or U11053 (N_11053,N_10676,N_10642);
and U11054 (N_11054,N_10557,N_10576);
nor U11055 (N_11055,N_10602,N_10958);
nand U11056 (N_11056,N_10972,N_10612);
and U11057 (N_11057,N_10870,N_10943);
nor U11058 (N_11058,N_10595,N_10953);
nor U11059 (N_11059,N_10667,N_10607);
or U11060 (N_11060,N_10816,N_10967);
nand U11061 (N_11061,N_10854,N_10799);
nand U11062 (N_11062,N_10549,N_10776);
nand U11063 (N_11063,N_10732,N_10987);
nand U11064 (N_11064,N_10821,N_10851);
or U11065 (N_11065,N_10832,N_10599);
nor U11066 (N_11066,N_10856,N_10911);
or U11067 (N_11067,N_10780,N_10639);
and U11068 (N_11068,N_10561,N_10948);
or U11069 (N_11069,N_10827,N_10848);
or U11070 (N_11070,N_10871,N_10920);
and U11071 (N_11071,N_10748,N_10888);
or U11072 (N_11072,N_10672,N_10551);
nor U11073 (N_11073,N_10834,N_10596);
nand U11074 (N_11074,N_10631,N_10741);
xnor U11075 (N_11075,N_10933,N_10555);
and U11076 (N_11076,N_10681,N_10841);
nor U11077 (N_11077,N_10685,N_10601);
or U11078 (N_11078,N_10621,N_10620);
xnor U11079 (N_11079,N_10652,N_10502);
nand U11080 (N_11080,N_10971,N_10650);
nor U11081 (N_11081,N_10819,N_10623);
or U11082 (N_11082,N_10553,N_10581);
nand U11083 (N_11083,N_10634,N_10939);
or U11084 (N_11084,N_10622,N_10700);
or U11085 (N_11085,N_10641,N_10575);
nor U11086 (N_11086,N_10932,N_10984);
xor U11087 (N_11087,N_10609,N_10670);
or U11088 (N_11088,N_10812,N_10828);
or U11089 (N_11089,N_10963,N_10616);
xnor U11090 (N_11090,N_10701,N_10929);
xnor U11091 (N_11091,N_10981,N_10790);
and U11092 (N_11092,N_10736,N_10591);
nor U11093 (N_11093,N_10938,N_10655);
and U11094 (N_11094,N_10783,N_10503);
nand U11095 (N_11095,N_10781,N_10895);
xnor U11096 (N_11096,N_10916,N_10528);
and U11097 (N_11097,N_10746,N_10860);
or U11098 (N_11098,N_10864,N_10578);
nand U11099 (N_11099,N_10768,N_10608);
nor U11100 (N_11100,N_10940,N_10535);
nor U11101 (N_11101,N_10894,N_10580);
nor U11102 (N_11102,N_10564,N_10945);
xor U11103 (N_11103,N_10857,N_10858);
nor U11104 (N_11104,N_10563,N_10833);
nand U11105 (N_11105,N_10887,N_10757);
xor U11106 (N_11106,N_10837,N_10802);
and U11107 (N_11107,N_10501,N_10500);
xor U11108 (N_11108,N_10784,N_10721);
nor U11109 (N_11109,N_10813,N_10879);
and U11110 (N_11110,N_10515,N_10570);
nor U11111 (N_11111,N_10914,N_10740);
and U11112 (N_11112,N_10946,N_10872);
nand U11113 (N_11113,N_10644,N_10649);
nand U11114 (N_11114,N_10654,N_10752);
nand U11115 (N_11115,N_10625,N_10973);
or U11116 (N_11116,N_10648,N_10547);
or U11117 (N_11117,N_10875,N_10537);
and U11118 (N_11118,N_10815,N_10898);
nor U11119 (N_11119,N_10797,N_10554);
and U11120 (N_11120,N_10782,N_10527);
xnor U11121 (N_11121,N_10931,N_10944);
xor U11122 (N_11122,N_10959,N_10545);
xor U11123 (N_11123,N_10588,N_10786);
nand U11124 (N_11124,N_10882,N_10719);
and U11125 (N_11125,N_10698,N_10846);
nor U11126 (N_11126,N_10678,N_10874);
nor U11127 (N_11127,N_10593,N_10558);
nand U11128 (N_11128,N_10635,N_10993);
xor U11129 (N_11129,N_10847,N_10806);
and U11130 (N_11130,N_10687,N_10704);
xor U11131 (N_11131,N_10992,N_10820);
nor U11132 (N_11132,N_10674,N_10976);
nand U11133 (N_11133,N_10660,N_10587);
or U11134 (N_11134,N_10517,N_10880);
nand U11135 (N_11135,N_10908,N_10540);
or U11136 (N_11136,N_10791,N_10831);
nand U11137 (N_11137,N_10533,N_10686);
or U11138 (N_11138,N_10747,N_10542);
or U11139 (N_11139,N_10629,N_10568);
xnor U11140 (N_11140,N_10653,N_10989);
xnor U11141 (N_11141,N_10966,N_10728);
and U11142 (N_11142,N_10628,N_10801);
xnor U11143 (N_11143,N_10921,N_10690);
and U11144 (N_11144,N_10705,N_10796);
or U11145 (N_11145,N_10569,N_10725);
nand U11146 (N_11146,N_10565,N_10717);
and U11147 (N_11147,N_10538,N_10531);
xor U11148 (N_11148,N_10520,N_10708);
xor U11149 (N_11149,N_10766,N_10618);
nand U11150 (N_11150,N_10900,N_10597);
nor U11151 (N_11151,N_10731,N_10519);
xnor U11152 (N_11152,N_10510,N_10859);
and U11153 (N_11153,N_10835,N_10624);
nand U11154 (N_11154,N_10556,N_10998);
xnor U11155 (N_11155,N_10903,N_10550);
or U11156 (N_11156,N_10863,N_10627);
xor U11157 (N_11157,N_10548,N_10904);
nor U11158 (N_11158,N_10829,N_10893);
xnor U11159 (N_11159,N_10941,N_10603);
xnor U11160 (N_11160,N_10518,N_10952);
and U11161 (N_11161,N_10892,N_10513);
nor U11162 (N_11162,N_10772,N_10600);
nand U11163 (N_11163,N_10886,N_10995);
and U11164 (N_11164,N_10977,N_10573);
xnor U11165 (N_11165,N_10954,N_10730);
nor U11166 (N_11166,N_10810,N_10696);
nor U11167 (N_11167,N_10613,N_10823);
and U11168 (N_11168,N_10969,N_10661);
and U11169 (N_11169,N_10571,N_10865);
nor U11170 (N_11170,N_10996,N_10915);
or U11171 (N_11171,N_10957,N_10878);
nor U11172 (N_11172,N_10805,N_10980);
and U11173 (N_11173,N_10523,N_10512);
or U11174 (N_11174,N_10755,N_10839);
and U11175 (N_11175,N_10694,N_10990);
xor U11176 (N_11176,N_10543,N_10733);
nand U11177 (N_11177,N_10814,N_10722);
or U11178 (N_11178,N_10978,N_10606);
and U11179 (N_11179,N_10584,N_10524);
and U11180 (N_11180,N_10912,N_10850);
and U11181 (N_11181,N_10988,N_10646);
xnor U11182 (N_11182,N_10785,N_10999);
nand U11183 (N_11183,N_10562,N_10675);
and U11184 (N_11184,N_10876,N_10918);
nand U11185 (N_11185,N_10727,N_10673);
xnor U11186 (N_11186,N_10657,N_10739);
nor U11187 (N_11187,N_10539,N_10822);
and U11188 (N_11188,N_10807,N_10884);
and U11189 (N_11189,N_10693,N_10633);
xnor U11190 (N_11190,N_10707,N_10811);
nand U11191 (N_11191,N_10712,N_10737);
xnor U11192 (N_11192,N_10713,N_10716);
xnor U11193 (N_11193,N_10949,N_10630);
xor U11194 (N_11194,N_10617,N_10855);
xor U11195 (N_11195,N_10511,N_10818);
xnor U11196 (N_11196,N_10695,N_10994);
nand U11197 (N_11197,N_10647,N_10985);
and U11198 (N_11198,N_10662,N_10777);
nor U11199 (N_11199,N_10928,N_10723);
xor U11200 (N_11200,N_10982,N_10795);
nor U11201 (N_11201,N_10809,N_10764);
nor U11202 (N_11202,N_10589,N_10508);
nand U11203 (N_11203,N_10817,N_10711);
nand U11204 (N_11204,N_10758,N_10925);
or U11205 (N_11205,N_10956,N_10779);
or U11206 (N_11206,N_10885,N_10724);
nor U11207 (N_11207,N_10913,N_10924);
nand U11208 (N_11208,N_10923,N_10643);
nand U11209 (N_11209,N_10836,N_10902);
or U11210 (N_11210,N_10504,N_10546);
nand U11211 (N_11211,N_10750,N_10826);
nand U11212 (N_11212,N_10699,N_10663);
nand U11213 (N_11213,N_10683,N_10866);
or U11214 (N_11214,N_10749,N_10574);
xor U11215 (N_11215,N_10594,N_10765);
nor U11216 (N_11216,N_10714,N_10552);
or U11217 (N_11217,N_10522,N_10968);
nand U11218 (N_11218,N_10745,N_10890);
nand U11219 (N_11219,N_10792,N_10682);
nand U11220 (N_11220,N_10521,N_10664);
and U11221 (N_11221,N_10734,N_10586);
xnor U11222 (N_11222,N_10636,N_10691);
or U11223 (N_11223,N_10710,N_10585);
and U11224 (N_11224,N_10656,N_10955);
nand U11225 (N_11225,N_10532,N_10808);
and U11226 (N_11226,N_10951,N_10770);
and U11227 (N_11227,N_10668,N_10830);
nor U11228 (N_11228,N_10997,N_10803);
and U11229 (N_11229,N_10910,N_10844);
nand U11230 (N_11230,N_10529,N_10919);
xnor U11231 (N_11231,N_10753,N_10787);
or U11232 (N_11232,N_10950,N_10909);
nand U11233 (N_11233,N_10658,N_10505);
nor U11234 (N_11234,N_10867,N_10974);
and U11235 (N_11235,N_10514,N_10640);
and U11236 (N_11236,N_10896,N_10793);
nand U11237 (N_11237,N_10582,N_10651);
or U11238 (N_11238,N_10937,N_10849);
xnor U11239 (N_11239,N_10889,N_10760);
xor U11240 (N_11240,N_10720,N_10964);
nand U11241 (N_11241,N_10926,N_10709);
xnor U11242 (N_11242,N_10927,N_10930);
and U11243 (N_11243,N_10577,N_10566);
and U11244 (N_11244,N_10798,N_10743);
nand U11245 (N_11245,N_10738,N_10754);
nand U11246 (N_11246,N_10590,N_10645);
xor U11247 (N_11247,N_10637,N_10697);
nand U11248 (N_11248,N_10544,N_10986);
and U11249 (N_11249,N_10917,N_10868);
and U11250 (N_11250,N_10794,N_10604);
and U11251 (N_11251,N_10956,N_10620);
nor U11252 (N_11252,N_10681,N_10788);
nand U11253 (N_11253,N_10876,N_10602);
and U11254 (N_11254,N_10726,N_10997);
nand U11255 (N_11255,N_10868,N_10743);
nand U11256 (N_11256,N_10936,N_10828);
nor U11257 (N_11257,N_10590,N_10627);
and U11258 (N_11258,N_10654,N_10876);
nand U11259 (N_11259,N_10842,N_10530);
nand U11260 (N_11260,N_10705,N_10910);
or U11261 (N_11261,N_10635,N_10765);
and U11262 (N_11262,N_10638,N_10715);
and U11263 (N_11263,N_10995,N_10917);
nor U11264 (N_11264,N_10756,N_10808);
or U11265 (N_11265,N_10935,N_10741);
nor U11266 (N_11266,N_10904,N_10739);
nand U11267 (N_11267,N_10795,N_10993);
or U11268 (N_11268,N_10973,N_10645);
nor U11269 (N_11269,N_10661,N_10744);
and U11270 (N_11270,N_10758,N_10555);
and U11271 (N_11271,N_10965,N_10934);
nand U11272 (N_11272,N_10604,N_10756);
and U11273 (N_11273,N_10522,N_10678);
or U11274 (N_11274,N_10684,N_10879);
nor U11275 (N_11275,N_10927,N_10751);
and U11276 (N_11276,N_10979,N_10600);
nand U11277 (N_11277,N_10899,N_10705);
xnor U11278 (N_11278,N_10534,N_10883);
or U11279 (N_11279,N_10959,N_10651);
and U11280 (N_11280,N_10691,N_10674);
xnor U11281 (N_11281,N_10961,N_10831);
nor U11282 (N_11282,N_10781,N_10875);
nor U11283 (N_11283,N_10712,N_10960);
and U11284 (N_11284,N_10596,N_10632);
nor U11285 (N_11285,N_10803,N_10762);
nor U11286 (N_11286,N_10754,N_10546);
nand U11287 (N_11287,N_10886,N_10582);
nand U11288 (N_11288,N_10625,N_10875);
nand U11289 (N_11289,N_10688,N_10669);
and U11290 (N_11290,N_10938,N_10960);
and U11291 (N_11291,N_10807,N_10864);
xor U11292 (N_11292,N_10559,N_10572);
nand U11293 (N_11293,N_10617,N_10760);
nand U11294 (N_11294,N_10808,N_10860);
or U11295 (N_11295,N_10995,N_10628);
nor U11296 (N_11296,N_10832,N_10866);
and U11297 (N_11297,N_10540,N_10819);
nand U11298 (N_11298,N_10954,N_10998);
or U11299 (N_11299,N_10930,N_10879);
or U11300 (N_11300,N_10810,N_10581);
nand U11301 (N_11301,N_10872,N_10798);
and U11302 (N_11302,N_10596,N_10946);
nand U11303 (N_11303,N_10576,N_10651);
and U11304 (N_11304,N_10526,N_10885);
xnor U11305 (N_11305,N_10693,N_10914);
nor U11306 (N_11306,N_10634,N_10990);
or U11307 (N_11307,N_10684,N_10968);
nand U11308 (N_11308,N_10946,N_10740);
and U11309 (N_11309,N_10527,N_10533);
nor U11310 (N_11310,N_10794,N_10655);
xnor U11311 (N_11311,N_10725,N_10756);
or U11312 (N_11312,N_10632,N_10646);
nand U11313 (N_11313,N_10930,N_10548);
nand U11314 (N_11314,N_10771,N_10988);
or U11315 (N_11315,N_10644,N_10875);
nor U11316 (N_11316,N_10756,N_10742);
nand U11317 (N_11317,N_10792,N_10607);
xor U11318 (N_11318,N_10855,N_10627);
or U11319 (N_11319,N_10613,N_10992);
nand U11320 (N_11320,N_10580,N_10886);
or U11321 (N_11321,N_10846,N_10752);
or U11322 (N_11322,N_10943,N_10795);
nor U11323 (N_11323,N_10676,N_10946);
xor U11324 (N_11324,N_10640,N_10910);
nor U11325 (N_11325,N_10861,N_10860);
and U11326 (N_11326,N_10935,N_10974);
nor U11327 (N_11327,N_10502,N_10546);
xnor U11328 (N_11328,N_10830,N_10532);
or U11329 (N_11329,N_10830,N_10938);
and U11330 (N_11330,N_10603,N_10773);
and U11331 (N_11331,N_10687,N_10942);
nor U11332 (N_11332,N_10696,N_10511);
nor U11333 (N_11333,N_10724,N_10565);
and U11334 (N_11334,N_10599,N_10654);
xnor U11335 (N_11335,N_10559,N_10757);
nor U11336 (N_11336,N_10866,N_10941);
xnor U11337 (N_11337,N_10661,N_10808);
xor U11338 (N_11338,N_10988,N_10900);
xnor U11339 (N_11339,N_10733,N_10682);
and U11340 (N_11340,N_10666,N_10799);
or U11341 (N_11341,N_10706,N_10953);
nand U11342 (N_11342,N_10645,N_10681);
and U11343 (N_11343,N_10993,N_10538);
nor U11344 (N_11344,N_10646,N_10913);
xnor U11345 (N_11345,N_10872,N_10653);
nor U11346 (N_11346,N_10949,N_10564);
or U11347 (N_11347,N_10555,N_10751);
nand U11348 (N_11348,N_10729,N_10859);
nand U11349 (N_11349,N_10728,N_10795);
nor U11350 (N_11350,N_10987,N_10639);
nor U11351 (N_11351,N_10571,N_10896);
xor U11352 (N_11352,N_10763,N_10577);
or U11353 (N_11353,N_10863,N_10517);
xnor U11354 (N_11354,N_10537,N_10585);
nand U11355 (N_11355,N_10599,N_10710);
nand U11356 (N_11356,N_10906,N_10777);
nor U11357 (N_11357,N_10553,N_10727);
nand U11358 (N_11358,N_10916,N_10788);
nor U11359 (N_11359,N_10563,N_10621);
or U11360 (N_11360,N_10962,N_10830);
or U11361 (N_11361,N_10591,N_10857);
and U11362 (N_11362,N_10838,N_10555);
or U11363 (N_11363,N_10660,N_10729);
and U11364 (N_11364,N_10707,N_10605);
xnor U11365 (N_11365,N_10912,N_10739);
nand U11366 (N_11366,N_10705,N_10708);
and U11367 (N_11367,N_10616,N_10905);
nand U11368 (N_11368,N_10959,N_10725);
xnor U11369 (N_11369,N_10967,N_10513);
xor U11370 (N_11370,N_10627,N_10940);
nand U11371 (N_11371,N_10824,N_10667);
nor U11372 (N_11372,N_10912,N_10501);
xnor U11373 (N_11373,N_10727,N_10644);
xnor U11374 (N_11374,N_10725,N_10646);
nand U11375 (N_11375,N_10728,N_10799);
xor U11376 (N_11376,N_10573,N_10965);
nor U11377 (N_11377,N_10860,N_10844);
and U11378 (N_11378,N_10708,N_10663);
and U11379 (N_11379,N_10699,N_10575);
nand U11380 (N_11380,N_10861,N_10854);
or U11381 (N_11381,N_10969,N_10915);
nand U11382 (N_11382,N_10951,N_10828);
nand U11383 (N_11383,N_10974,N_10552);
xnor U11384 (N_11384,N_10992,N_10605);
or U11385 (N_11385,N_10644,N_10759);
or U11386 (N_11386,N_10505,N_10728);
nor U11387 (N_11387,N_10767,N_10625);
nor U11388 (N_11388,N_10872,N_10527);
xor U11389 (N_11389,N_10581,N_10978);
and U11390 (N_11390,N_10561,N_10510);
nand U11391 (N_11391,N_10764,N_10676);
and U11392 (N_11392,N_10994,N_10945);
nand U11393 (N_11393,N_10798,N_10606);
nor U11394 (N_11394,N_10784,N_10990);
and U11395 (N_11395,N_10986,N_10985);
xnor U11396 (N_11396,N_10644,N_10900);
nand U11397 (N_11397,N_10694,N_10899);
or U11398 (N_11398,N_10793,N_10987);
nand U11399 (N_11399,N_10594,N_10981);
or U11400 (N_11400,N_10826,N_10516);
xor U11401 (N_11401,N_10704,N_10646);
and U11402 (N_11402,N_10899,N_10756);
xor U11403 (N_11403,N_10791,N_10611);
or U11404 (N_11404,N_10803,N_10821);
or U11405 (N_11405,N_10534,N_10662);
nor U11406 (N_11406,N_10519,N_10784);
nor U11407 (N_11407,N_10605,N_10806);
and U11408 (N_11408,N_10917,N_10690);
nor U11409 (N_11409,N_10809,N_10699);
nand U11410 (N_11410,N_10544,N_10938);
nand U11411 (N_11411,N_10841,N_10826);
or U11412 (N_11412,N_10890,N_10526);
or U11413 (N_11413,N_10708,N_10826);
and U11414 (N_11414,N_10789,N_10792);
or U11415 (N_11415,N_10791,N_10934);
nor U11416 (N_11416,N_10986,N_10803);
nor U11417 (N_11417,N_10781,N_10633);
and U11418 (N_11418,N_10872,N_10721);
xnor U11419 (N_11419,N_10648,N_10663);
and U11420 (N_11420,N_10910,N_10856);
xnor U11421 (N_11421,N_10755,N_10665);
and U11422 (N_11422,N_10847,N_10963);
nand U11423 (N_11423,N_10620,N_10886);
nand U11424 (N_11424,N_10826,N_10887);
and U11425 (N_11425,N_10628,N_10577);
nor U11426 (N_11426,N_10571,N_10603);
nor U11427 (N_11427,N_10573,N_10792);
and U11428 (N_11428,N_10976,N_10537);
and U11429 (N_11429,N_10613,N_10712);
and U11430 (N_11430,N_10874,N_10943);
nand U11431 (N_11431,N_10607,N_10666);
nand U11432 (N_11432,N_10609,N_10880);
xor U11433 (N_11433,N_10531,N_10902);
and U11434 (N_11434,N_10969,N_10834);
nand U11435 (N_11435,N_10623,N_10870);
and U11436 (N_11436,N_10761,N_10737);
and U11437 (N_11437,N_10635,N_10606);
xor U11438 (N_11438,N_10875,N_10563);
nor U11439 (N_11439,N_10624,N_10506);
nor U11440 (N_11440,N_10836,N_10690);
nor U11441 (N_11441,N_10578,N_10722);
nor U11442 (N_11442,N_10619,N_10577);
or U11443 (N_11443,N_10573,N_10732);
nand U11444 (N_11444,N_10637,N_10972);
nor U11445 (N_11445,N_10784,N_10568);
nand U11446 (N_11446,N_10744,N_10766);
nand U11447 (N_11447,N_10927,N_10924);
and U11448 (N_11448,N_10583,N_10707);
nand U11449 (N_11449,N_10553,N_10730);
nor U11450 (N_11450,N_10801,N_10823);
and U11451 (N_11451,N_10516,N_10844);
nand U11452 (N_11452,N_10576,N_10546);
xnor U11453 (N_11453,N_10810,N_10840);
or U11454 (N_11454,N_10833,N_10704);
xor U11455 (N_11455,N_10825,N_10890);
and U11456 (N_11456,N_10916,N_10721);
xnor U11457 (N_11457,N_10863,N_10932);
xor U11458 (N_11458,N_10704,N_10511);
xor U11459 (N_11459,N_10668,N_10719);
xor U11460 (N_11460,N_10962,N_10946);
or U11461 (N_11461,N_10534,N_10958);
and U11462 (N_11462,N_10511,N_10746);
nor U11463 (N_11463,N_10677,N_10521);
and U11464 (N_11464,N_10831,N_10833);
xor U11465 (N_11465,N_10721,N_10902);
or U11466 (N_11466,N_10510,N_10923);
xnor U11467 (N_11467,N_10711,N_10945);
and U11468 (N_11468,N_10808,N_10545);
and U11469 (N_11469,N_10615,N_10582);
nor U11470 (N_11470,N_10766,N_10578);
and U11471 (N_11471,N_10690,N_10502);
nor U11472 (N_11472,N_10860,N_10867);
xor U11473 (N_11473,N_10875,N_10585);
nor U11474 (N_11474,N_10546,N_10592);
nand U11475 (N_11475,N_10739,N_10874);
xor U11476 (N_11476,N_10869,N_10974);
or U11477 (N_11477,N_10899,N_10785);
nor U11478 (N_11478,N_10737,N_10984);
and U11479 (N_11479,N_10803,N_10996);
and U11480 (N_11480,N_10853,N_10751);
and U11481 (N_11481,N_10516,N_10861);
or U11482 (N_11482,N_10807,N_10652);
nor U11483 (N_11483,N_10565,N_10560);
nand U11484 (N_11484,N_10711,N_10900);
nor U11485 (N_11485,N_10512,N_10704);
nor U11486 (N_11486,N_10681,N_10594);
or U11487 (N_11487,N_10980,N_10921);
nand U11488 (N_11488,N_10614,N_10771);
nand U11489 (N_11489,N_10743,N_10860);
and U11490 (N_11490,N_10915,N_10698);
and U11491 (N_11491,N_10991,N_10585);
nand U11492 (N_11492,N_10556,N_10587);
and U11493 (N_11493,N_10806,N_10720);
and U11494 (N_11494,N_10749,N_10910);
nand U11495 (N_11495,N_10764,N_10507);
or U11496 (N_11496,N_10955,N_10660);
xnor U11497 (N_11497,N_10502,N_10510);
or U11498 (N_11498,N_10531,N_10661);
xor U11499 (N_11499,N_10802,N_10632);
or U11500 (N_11500,N_11112,N_11298);
or U11501 (N_11501,N_11049,N_11452);
or U11502 (N_11502,N_11394,N_11254);
or U11503 (N_11503,N_11231,N_11363);
or U11504 (N_11504,N_11270,N_11299);
nor U11505 (N_11505,N_11409,N_11309);
or U11506 (N_11506,N_11007,N_11288);
nand U11507 (N_11507,N_11241,N_11232);
xnor U11508 (N_11508,N_11424,N_11369);
or U11509 (N_11509,N_11017,N_11342);
xnor U11510 (N_11510,N_11258,N_11196);
nand U11511 (N_11511,N_11395,N_11066);
and U11512 (N_11512,N_11463,N_11084);
nand U11513 (N_11513,N_11466,N_11477);
nor U11514 (N_11514,N_11350,N_11286);
xnor U11515 (N_11515,N_11328,N_11485);
nor U11516 (N_11516,N_11287,N_11207);
and U11517 (N_11517,N_11190,N_11205);
or U11518 (N_11518,N_11300,N_11474);
and U11519 (N_11519,N_11406,N_11158);
nand U11520 (N_11520,N_11365,N_11386);
and U11521 (N_11521,N_11292,N_11398);
xnor U11522 (N_11522,N_11175,N_11295);
and U11523 (N_11523,N_11281,N_11070);
and U11524 (N_11524,N_11234,N_11100);
or U11525 (N_11525,N_11156,N_11255);
and U11526 (N_11526,N_11347,N_11054);
nor U11527 (N_11527,N_11097,N_11072);
or U11528 (N_11528,N_11227,N_11319);
or U11529 (N_11529,N_11191,N_11020);
nor U11530 (N_11530,N_11252,N_11229);
and U11531 (N_11531,N_11022,N_11348);
xor U11532 (N_11532,N_11098,N_11338);
or U11533 (N_11533,N_11310,N_11472);
or U11534 (N_11534,N_11060,N_11094);
xnor U11535 (N_11535,N_11499,N_11491);
nor U11536 (N_11536,N_11497,N_11460);
xnor U11537 (N_11537,N_11351,N_11023);
nand U11538 (N_11538,N_11279,N_11004);
nor U11539 (N_11539,N_11128,N_11178);
nand U11540 (N_11540,N_11462,N_11407);
nor U11541 (N_11541,N_11129,N_11396);
xnor U11542 (N_11542,N_11102,N_11036);
nor U11543 (N_11543,N_11177,N_11256);
or U11544 (N_11544,N_11385,N_11087);
nor U11545 (N_11545,N_11449,N_11275);
nand U11546 (N_11546,N_11209,N_11186);
nand U11547 (N_11547,N_11239,N_11495);
or U11548 (N_11548,N_11142,N_11290);
nor U11549 (N_11549,N_11431,N_11006);
and U11550 (N_11550,N_11088,N_11170);
or U11551 (N_11551,N_11243,N_11030);
nand U11552 (N_11552,N_11179,N_11195);
and U11553 (N_11553,N_11215,N_11494);
xor U11554 (N_11554,N_11492,N_11330);
and U11555 (N_11555,N_11135,N_11113);
and U11556 (N_11556,N_11235,N_11005);
or U11557 (N_11557,N_11289,N_11109);
or U11558 (N_11558,N_11050,N_11326);
nor U11559 (N_11559,N_11484,N_11206);
and U11560 (N_11560,N_11199,N_11151);
or U11561 (N_11561,N_11172,N_11306);
xor U11562 (N_11562,N_11317,N_11487);
xor U11563 (N_11563,N_11180,N_11169);
and U11564 (N_11564,N_11440,N_11481);
and U11565 (N_11565,N_11184,N_11391);
nand U11566 (N_11566,N_11273,N_11403);
and U11567 (N_11567,N_11435,N_11405);
or U11568 (N_11568,N_11046,N_11422);
or U11569 (N_11569,N_11441,N_11321);
nand U11570 (N_11570,N_11136,N_11305);
or U11571 (N_11571,N_11411,N_11019);
and U11572 (N_11572,N_11119,N_11436);
or U11573 (N_11573,N_11160,N_11442);
nand U11574 (N_11574,N_11304,N_11237);
nor U11575 (N_11575,N_11408,N_11147);
or U11576 (N_11576,N_11444,N_11498);
nor U11577 (N_11577,N_11220,N_11001);
nor U11578 (N_11578,N_11427,N_11111);
xor U11579 (N_11579,N_11473,N_11013);
xnor U11580 (N_11580,N_11373,N_11397);
nor U11581 (N_11581,N_11090,N_11134);
xor U11582 (N_11582,N_11432,N_11114);
nor U11583 (N_11583,N_11340,N_11312);
or U11584 (N_11584,N_11464,N_11371);
nand U11585 (N_11585,N_11166,N_11272);
nand U11586 (N_11586,N_11461,N_11382);
and U11587 (N_11587,N_11092,N_11245);
or U11588 (N_11588,N_11041,N_11390);
and U11589 (N_11589,N_11198,N_11325);
xor U11590 (N_11590,N_11341,N_11434);
or U11591 (N_11591,N_11155,N_11426);
or U11592 (N_11592,N_11327,N_11323);
nor U11593 (N_11593,N_11250,N_11193);
nand U11594 (N_11594,N_11257,N_11367);
or U11595 (N_11595,N_11116,N_11419);
or U11596 (N_11596,N_11459,N_11211);
nand U11597 (N_11597,N_11318,N_11366);
nor U11598 (N_11598,N_11354,N_11152);
or U11599 (N_11599,N_11058,N_11331);
and U11600 (N_11600,N_11133,N_11101);
xor U11601 (N_11601,N_11471,N_11031);
or U11602 (N_11602,N_11187,N_11453);
xor U11603 (N_11603,N_11271,N_11455);
nor U11604 (N_11604,N_11416,N_11131);
nand U11605 (N_11605,N_11439,N_11115);
xor U11606 (N_11606,N_11410,N_11110);
or U11607 (N_11607,N_11016,N_11430);
or U11608 (N_11608,N_11345,N_11073);
or U11609 (N_11609,N_11141,N_11042);
nand U11610 (N_11610,N_11470,N_11285);
or U11611 (N_11611,N_11238,N_11414);
nor U11612 (N_11612,N_11208,N_11105);
nor U11613 (N_11613,N_11081,N_11329);
xnor U11614 (N_11614,N_11037,N_11143);
nand U11615 (N_11615,N_11099,N_11139);
nand U11616 (N_11616,N_11266,N_11448);
nand U11617 (N_11617,N_11149,N_11138);
nand U11618 (N_11618,N_11322,N_11202);
nand U11619 (N_11619,N_11228,N_11320);
nor U11620 (N_11620,N_11248,N_11388);
xor U11621 (N_11621,N_11224,N_11137);
xnor U11622 (N_11622,N_11358,N_11075);
nand U11623 (N_11623,N_11264,N_11085);
or U11624 (N_11624,N_11417,N_11233);
nor U11625 (N_11625,N_11401,N_11200);
nand U11626 (N_11626,N_11118,N_11011);
nand U11627 (N_11627,N_11103,N_11026);
or U11628 (N_11628,N_11384,N_11475);
or U11629 (N_11629,N_11380,N_11337);
nor U11630 (N_11630,N_11402,N_11478);
and U11631 (N_11631,N_11488,N_11167);
xnor U11632 (N_11632,N_11324,N_11284);
nor U11633 (N_11633,N_11486,N_11443);
nor U11634 (N_11634,N_11123,N_11104);
nor U11635 (N_11635,N_11218,N_11379);
nor U11636 (N_11636,N_11413,N_11062);
and U11637 (N_11637,N_11376,N_11236);
nor U11638 (N_11638,N_11387,N_11389);
nand U11639 (N_11639,N_11009,N_11377);
nand U11640 (N_11640,N_11421,N_11428);
and U11641 (N_11641,N_11400,N_11045);
xnor U11642 (N_11642,N_11153,N_11311);
nor U11643 (N_11643,N_11213,N_11047);
and U11644 (N_11644,N_11165,N_11018);
or U11645 (N_11645,N_11032,N_11360);
nor U11646 (N_11646,N_11242,N_11127);
nand U11647 (N_11647,N_11126,N_11159);
nand U11648 (N_11648,N_11489,N_11483);
nor U11649 (N_11649,N_11185,N_11482);
nand U11650 (N_11650,N_11253,N_11124);
xor U11651 (N_11651,N_11450,N_11192);
nand U11652 (N_11652,N_11003,N_11044);
nand U11653 (N_11653,N_11121,N_11339);
nand U11654 (N_11654,N_11399,N_11189);
and U11655 (N_11655,N_11067,N_11313);
or U11656 (N_11656,N_11061,N_11425);
and U11657 (N_11657,N_11162,N_11146);
and U11658 (N_11658,N_11219,N_11000);
or U11659 (N_11659,N_11035,N_11040);
and U11660 (N_11660,N_11217,N_11336);
and U11661 (N_11661,N_11262,N_11423);
nor U11662 (N_11662,N_11274,N_11353);
and U11663 (N_11663,N_11161,N_11480);
and U11664 (N_11664,N_11157,N_11107);
or U11665 (N_11665,N_11445,N_11210);
nand U11666 (N_11666,N_11335,N_11294);
or U11667 (N_11667,N_11028,N_11469);
nand U11668 (N_11668,N_11034,N_11182);
nand U11669 (N_11669,N_11008,N_11203);
nor U11670 (N_11670,N_11333,N_11029);
xnor U11671 (N_11671,N_11214,N_11240);
nand U11672 (N_11672,N_11053,N_11267);
nor U11673 (N_11673,N_11490,N_11089);
or U11674 (N_11674,N_11154,N_11260);
nor U11675 (N_11675,N_11244,N_11144);
and U11676 (N_11676,N_11173,N_11392);
xnor U11677 (N_11677,N_11343,N_11457);
nor U11678 (N_11678,N_11280,N_11496);
xnor U11679 (N_11679,N_11226,N_11316);
xnor U11680 (N_11680,N_11375,N_11188);
or U11681 (N_11681,N_11171,N_11269);
or U11682 (N_11682,N_11130,N_11314);
or U11683 (N_11683,N_11117,N_11012);
xnor U11684 (N_11684,N_11212,N_11216);
and U11685 (N_11685,N_11378,N_11420);
nor U11686 (N_11686,N_11451,N_11263);
nor U11687 (N_11687,N_11438,N_11282);
and U11688 (N_11688,N_11194,N_11374);
nand U11689 (N_11689,N_11468,N_11251);
or U11690 (N_11690,N_11064,N_11145);
nor U11691 (N_11691,N_11043,N_11063);
xor U11692 (N_11692,N_11249,N_11176);
or U11693 (N_11693,N_11059,N_11412);
nand U11694 (N_11694,N_11204,N_11078);
xnor U11695 (N_11695,N_11148,N_11002);
nor U11696 (N_11696,N_11476,N_11021);
nor U11697 (N_11697,N_11164,N_11024);
xor U11698 (N_11698,N_11091,N_11296);
and U11699 (N_11699,N_11015,N_11247);
nand U11700 (N_11700,N_11381,N_11467);
nor U11701 (N_11701,N_11074,N_11181);
or U11702 (N_11702,N_11297,N_11418);
nor U11703 (N_11703,N_11068,N_11246);
nor U11704 (N_11704,N_11291,N_11458);
or U11705 (N_11705,N_11069,N_11307);
nor U11706 (N_11706,N_11225,N_11259);
and U11707 (N_11707,N_11276,N_11056);
or U11708 (N_11708,N_11076,N_11301);
nand U11709 (N_11709,N_11080,N_11261);
nor U11710 (N_11710,N_11393,N_11132);
and U11711 (N_11711,N_11071,N_11052);
or U11712 (N_11712,N_11222,N_11014);
xor U11713 (N_11713,N_11095,N_11352);
nor U11714 (N_11714,N_11346,N_11278);
nand U11715 (N_11715,N_11303,N_11163);
nor U11716 (N_11716,N_11221,N_11372);
nand U11717 (N_11717,N_11230,N_11283);
xnor U11718 (N_11718,N_11308,N_11361);
nor U11719 (N_11719,N_11174,N_11357);
nor U11720 (N_11720,N_11447,N_11010);
or U11721 (N_11721,N_11302,N_11106);
or U11722 (N_11722,N_11033,N_11082);
nor U11723 (N_11723,N_11027,N_11349);
nor U11724 (N_11724,N_11093,N_11083);
and U11725 (N_11725,N_11493,N_11446);
xor U11726 (N_11726,N_11140,N_11368);
and U11727 (N_11727,N_11150,N_11293);
and U11728 (N_11728,N_11429,N_11055);
xor U11729 (N_11729,N_11201,N_11415);
nand U11730 (N_11730,N_11079,N_11404);
and U11731 (N_11731,N_11362,N_11077);
or U11732 (N_11732,N_11086,N_11364);
nand U11733 (N_11733,N_11334,N_11265);
xor U11734 (N_11734,N_11356,N_11465);
or U11735 (N_11735,N_11120,N_11057);
or U11736 (N_11736,N_11051,N_11197);
or U11737 (N_11737,N_11108,N_11355);
xnor U11738 (N_11738,N_11437,N_11454);
or U11739 (N_11739,N_11370,N_11048);
nor U11740 (N_11740,N_11332,N_11065);
or U11741 (N_11741,N_11125,N_11315);
xnor U11742 (N_11742,N_11096,N_11025);
nor U11743 (N_11743,N_11039,N_11479);
nand U11744 (N_11744,N_11168,N_11383);
nand U11745 (N_11745,N_11038,N_11277);
and U11746 (N_11746,N_11344,N_11183);
nand U11747 (N_11747,N_11122,N_11359);
or U11748 (N_11748,N_11456,N_11433);
xor U11749 (N_11749,N_11223,N_11268);
nor U11750 (N_11750,N_11276,N_11179);
nand U11751 (N_11751,N_11088,N_11151);
and U11752 (N_11752,N_11123,N_11393);
nor U11753 (N_11753,N_11081,N_11077);
xor U11754 (N_11754,N_11167,N_11149);
or U11755 (N_11755,N_11484,N_11223);
xor U11756 (N_11756,N_11198,N_11494);
and U11757 (N_11757,N_11227,N_11192);
xor U11758 (N_11758,N_11226,N_11416);
xor U11759 (N_11759,N_11001,N_11151);
xor U11760 (N_11760,N_11312,N_11307);
nor U11761 (N_11761,N_11392,N_11353);
nor U11762 (N_11762,N_11448,N_11165);
nand U11763 (N_11763,N_11267,N_11407);
xnor U11764 (N_11764,N_11372,N_11186);
nor U11765 (N_11765,N_11215,N_11157);
or U11766 (N_11766,N_11162,N_11400);
and U11767 (N_11767,N_11013,N_11110);
nor U11768 (N_11768,N_11279,N_11117);
xnor U11769 (N_11769,N_11288,N_11212);
or U11770 (N_11770,N_11036,N_11303);
and U11771 (N_11771,N_11206,N_11129);
xor U11772 (N_11772,N_11200,N_11158);
nor U11773 (N_11773,N_11298,N_11370);
nor U11774 (N_11774,N_11181,N_11125);
and U11775 (N_11775,N_11095,N_11177);
and U11776 (N_11776,N_11410,N_11336);
xnor U11777 (N_11777,N_11494,N_11274);
nand U11778 (N_11778,N_11117,N_11240);
xnor U11779 (N_11779,N_11112,N_11497);
nand U11780 (N_11780,N_11205,N_11458);
and U11781 (N_11781,N_11399,N_11192);
and U11782 (N_11782,N_11480,N_11195);
xor U11783 (N_11783,N_11249,N_11066);
or U11784 (N_11784,N_11284,N_11018);
or U11785 (N_11785,N_11463,N_11494);
or U11786 (N_11786,N_11051,N_11396);
or U11787 (N_11787,N_11019,N_11110);
nor U11788 (N_11788,N_11268,N_11444);
and U11789 (N_11789,N_11402,N_11264);
and U11790 (N_11790,N_11042,N_11367);
xnor U11791 (N_11791,N_11484,N_11478);
xor U11792 (N_11792,N_11193,N_11071);
and U11793 (N_11793,N_11168,N_11127);
xor U11794 (N_11794,N_11385,N_11236);
xnor U11795 (N_11795,N_11284,N_11209);
xnor U11796 (N_11796,N_11135,N_11383);
and U11797 (N_11797,N_11485,N_11487);
or U11798 (N_11798,N_11179,N_11411);
or U11799 (N_11799,N_11211,N_11114);
and U11800 (N_11800,N_11036,N_11284);
xor U11801 (N_11801,N_11197,N_11376);
xor U11802 (N_11802,N_11065,N_11482);
or U11803 (N_11803,N_11001,N_11377);
and U11804 (N_11804,N_11490,N_11216);
and U11805 (N_11805,N_11344,N_11306);
nand U11806 (N_11806,N_11406,N_11063);
or U11807 (N_11807,N_11142,N_11287);
or U11808 (N_11808,N_11073,N_11397);
and U11809 (N_11809,N_11197,N_11390);
and U11810 (N_11810,N_11398,N_11162);
xor U11811 (N_11811,N_11047,N_11306);
xor U11812 (N_11812,N_11015,N_11394);
xor U11813 (N_11813,N_11104,N_11037);
nand U11814 (N_11814,N_11176,N_11046);
nor U11815 (N_11815,N_11081,N_11063);
nand U11816 (N_11816,N_11328,N_11479);
xnor U11817 (N_11817,N_11030,N_11337);
nand U11818 (N_11818,N_11177,N_11170);
xor U11819 (N_11819,N_11243,N_11302);
or U11820 (N_11820,N_11435,N_11234);
xnor U11821 (N_11821,N_11397,N_11049);
or U11822 (N_11822,N_11225,N_11471);
xnor U11823 (N_11823,N_11087,N_11349);
nor U11824 (N_11824,N_11197,N_11264);
xor U11825 (N_11825,N_11387,N_11325);
nand U11826 (N_11826,N_11333,N_11033);
nor U11827 (N_11827,N_11123,N_11358);
or U11828 (N_11828,N_11419,N_11160);
xnor U11829 (N_11829,N_11409,N_11043);
or U11830 (N_11830,N_11414,N_11150);
nor U11831 (N_11831,N_11187,N_11296);
xor U11832 (N_11832,N_11319,N_11360);
nand U11833 (N_11833,N_11263,N_11342);
and U11834 (N_11834,N_11398,N_11409);
nand U11835 (N_11835,N_11253,N_11458);
xor U11836 (N_11836,N_11322,N_11052);
or U11837 (N_11837,N_11004,N_11295);
or U11838 (N_11838,N_11027,N_11021);
xor U11839 (N_11839,N_11305,N_11431);
nor U11840 (N_11840,N_11442,N_11329);
or U11841 (N_11841,N_11054,N_11238);
nor U11842 (N_11842,N_11175,N_11357);
or U11843 (N_11843,N_11385,N_11435);
nor U11844 (N_11844,N_11142,N_11176);
nor U11845 (N_11845,N_11051,N_11125);
nand U11846 (N_11846,N_11486,N_11288);
nand U11847 (N_11847,N_11140,N_11170);
nor U11848 (N_11848,N_11246,N_11164);
nand U11849 (N_11849,N_11497,N_11248);
nand U11850 (N_11850,N_11396,N_11217);
and U11851 (N_11851,N_11463,N_11308);
or U11852 (N_11852,N_11115,N_11073);
and U11853 (N_11853,N_11375,N_11017);
xor U11854 (N_11854,N_11417,N_11465);
nand U11855 (N_11855,N_11459,N_11149);
nand U11856 (N_11856,N_11175,N_11434);
or U11857 (N_11857,N_11134,N_11117);
or U11858 (N_11858,N_11322,N_11177);
and U11859 (N_11859,N_11390,N_11404);
or U11860 (N_11860,N_11400,N_11476);
nor U11861 (N_11861,N_11278,N_11487);
nand U11862 (N_11862,N_11025,N_11042);
and U11863 (N_11863,N_11457,N_11280);
and U11864 (N_11864,N_11424,N_11216);
nand U11865 (N_11865,N_11202,N_11268);
and U11866 (N_11866,N_11351,N_11193);
xnor U11867 (N_11867,N_11070,N_11496);
xor U11868 (N_11868,N_11456,N_11190);
nor U11869 (N_11869,N_11424,N_11179);
nand U11870 (N_11870,N_11365,N_11287);
nand U11871 (N_11871,N_11362,N_11457);
or U11872 (N_11872,N_11020,N_11114);
or U11873 (N_11873,N_11427,N_11012);
nand U11874 (N_11874,N_11201,N_11313);
nand U11875 (N_11875,N_11408,N_11030);
nor U11876 (N_11876,N_11440,N_11371);
nand U11877 (N_11877,N_11232,N_11064);
xnor U11878 (N_11878,N_11465,N_11049);
or U11879 (N_11879,N_11164,N_11240);
xnor U11880 (N_11880,N_11013,N_11188);
or U11881 (N_11881,N_11352,N_11382);
and U11882 (N_11882,N_11453,N_11289);
nor U11883 (N_11883,N_11246,N_11433);
xnor U11884 (N_11884,N_11248,N_11218);
xnor U11885 (N_11885,N_11377,N_11269);
or U11886 (N_11886,N_11020,N_11401);
nand U11887 (N_11887,N_11204,N_11244);
xor U11888 (N_11888,N_11393,N_11160);
nor U11889 (N_11889,N_11045,N_11081);
nand U11890 (N_11890,N_11360,N_11113);
nor U11891 (N_11891,N_11388,N_11496);
and U11892 (N_11892,N_11475,N_11263);
nand U11893 (N_11893,N_11065,N_11477);
and U11894 (N_11894,N_11123,N_11458);
xnor U11895 (N_11895,N_11263,N_11249);
and U11896 (N_11896,N_11183,N_11028);
nor U11897 (N_11897,N_11338,N_11157);
nand U11898 (N_11898,N_11474,N_11248);
and U11899 (N_11899,N_11347,N_11484);
nor U11900 (N_11900,N_11153,N_11363);
nand U11901 (N_11901,N_11275,N_11306);
and U11902 (N_11902,N_11364,N_11456);
xor U11903 (N_11903,N_11075,N_11258);
xor U11904 (N_11904,N_11253,N_11489);
nand U11905 (N_11905,N_11274,N_11447);
xnor U11906 (N_11906,N_11235,N_11034);
nand U11907 (N_11907,N_11162,N_11467);
nor U11908 (N_11908,N_11308,N_11107);
nor U11909 (N_11909,N_11332,N_11131);
or U11910 (N_11910,N_11287,N_11325);
nor U11911 (N_11911,N_11226,N_11117);
xnor U11912 (N_11912,N_11324,N_11052);
nor U11913 (N_11913,N_11254,N_11045);
and U11914 (N_11914,N_11087,N_11090);
or U11915 (N_11915,N_11335,N_11375);
or U11916 (N_11916,N_11175,N_11280);
and U11917 (N_11917,N_11183,N_11061);
xor U11918 (N_11918,N_11172,N_11064);
nor U11919 (N_11919,N_11308,N_11039);
xnor U11920 (N_11920,N_11033,N_11335);
and U11921 (N_11921,N_11311,N_11155);
and U11922 (N_11922,N_11485,N_11361);
nor U11923 (N_11923,N_11263,N_11149);
and U11924 (N_11924,N_11498,N_11333);
xor U11925 (N_11925,N_11075,N_11107);
nor U11926 (N_11926,N_11260,N_11225);
and U11927 (N_11927,N_11217,N_11411);
xor U11928 (N_11928,N_11057,N_11143);
nor U11929 (N_11929,N_11307,N_11420);
nand U11930 (N_11930,N_11456,N_11225);
or U11931 (N_11931,N_11454,N_11498);
nor U11932 (N_11932,N_11101,N_11338);
nor U11933 (N_11933,N_11323,N_11452);
xnor U11934 (N_11934,N_11025,N_11171);
nor U11935 (N_11935,N_11139,N_11129);
nand U11936 (N_11936,N_11228,N_11415);
nand U11937 (N_11937,N_11245,N_11256);
nor U11938 (N_11938,N_11430,N_11182);
nor U11939 (N_11939,N_11427,N_11321);
nand U11940 (N_11940,N_11033,N_11289);
nand U11941 (N_11941,N_11338,N_11290);
nor U11942 (N_11942,N_11042,N_11252);
and U11943 (N_11943,N_11499,N_11126);
xnor U11944 (N_11944,N_11429,N_11118);
or U11945 (N_11945,N_11486,N_11274);
xnor U11946 (N_11946,N_11409,N_11271);
and U11947 (N_11947,N_11324,N_11128);
xor U11948 (N_11948,N_11103,N_11188);
and U11949 (N_11949,N_11451,N_11257);
xor U11950 (N_11950,N_11124,N_11382);
nor U11951 (N_11951,N_11321,N_11419);
nor U11952 (N_11952,N_11364,N_11067);
xor U11953 (N_11953,N_11148,N_11228);
xnor U11954 (N_11954,N_11494,N_11061);
nor U11955 (N_11955,N_11403,N_11390);
and U11956 (N_11956,N_11451,N_11370);
xor U11957 (N_11957,N_11043,N_11309);
nand U11958 (N_11958,N_11479,N_11238);
nor U11959 (N_11959,N_11401,N_11215);
xor U11960 (N_11960,N_11236,N_11401);
and U11961 (N_11961,N_11457,N_11065);
or U11962 (N_11962,N_11389,N_11261);
xnor U11963 (N_11963,N_11176,N_11203);
and U11964 (N_11964,N_11403,N_11456);
nor U11965 (N_11965,N_11190,N_11133);
xor U11966 (N_11966,N_11492,N_11487);
or U11967 (N_11967,N_11001,N_11235);
or U11968 (N_11968,N_11460,N_11476);
or U11969 (N_11969,N_11193,N_11424);
or U11970 (N_11970,N_11102,N_11360);
xor U11971 (N_11971,N_11362,N_11492);
nand U11972 (N_11972,N_11055,N_11143);
xor U11973 (N_11973,N_11034,N_11416);
and U11974 (N_11974,N_11280,N_11027);
or U11975 (N_11975,N_11463,N_11434);
nor U11976 (N_11976,N_11176,N_11155);
or U11977 (N_11977,N_11041,N_11000);
xor U11978 (N_11978,N_11333,N_11436);
or U11979 (N_11979,N_11334,N_11072);
xnor U11980 (N_11980,N_11344,N_11046);
or U11981 (N_11981,N_11211,N_11393);
xnor U11982 (N_11982,N_11264,N_11490);
and U11983 (N_11983,N_11084,N_11091);
nor U11984 (N_11984,N_11148,N_11251);
nand U11985 (N_11985,N_11436,N_11211);
nand U11986 (N_11986,N_11062,N_11300);
xnor U11987 (N_11987,N_11186,N_11417);
and U11988 (N_11988,N_11469,N_11423);
nand U11989 (N_11989,N_11310,N_11394);
or U11990 (N_11990,N_11267,N_11362);
nand U11991 (N_11991,N_11395,N_11468);
or U11992 (N_11992,N_11379,N_11135);
nand U11993 (N_11993,N_11174,N_11481);
nor U11994 (N_11994,N_11451,N_11387);
xor U11995 (N_11995,N_11078,N_11446);
and U11996 (N_11996,N_11026,N_11145);
xor U11997 (N_11997,N_11153,N_11049);
nor U11998 (N_11998,N_11342,N_11055);
and U11999 (N_11999,N_11158,N_11172);
xor U12000 (N_12000,N_11514,N_11531);
nor U12001 (N_12001,N_11976,N_11629);
or U12002 (N_12002,N_11769,N_11625);
nand U12003 (N_12003,N_11548,N_11800);
nor U12004 (N_12004,N_11960,N_11890);
nor U12005 (N_12005,N_11705,N_11693);
nor U12006 (N_12006,N_11538,N_11750);
nand U12007 (N_12007,N_11650,N_11738);
xor U12008 (N_12008,N_11661,N_11667);
or U12009 (N_12009,N_11555,N_11784);
or U12010 (N_12010,N_11528,N_11993);
xnor U12011 (N_12011,N_11745,N_11541);
nand U12012 (N_12012,N_11992,N_11668);
nor U12013 (N_12013,N_11512,N_11771);
nand U12014 (N_12014,N_11818,N_11766);
nand U12015 (N_12015,N_11967,N_11916);
xor U12016 (N_12016,N_11898,N_11713);
or U12017 (N_12017,N_11994,N_11982);
nand U12018 (N_12018,N_11809,N_11804);
nor U12019 (N_12019,N_11805,N_11588);
xnor U12020 (N_12020,N_11817,N_11795);
and U12021 (N_12021,N_11663,N_11664);
and U12022 (N_12022,N_11787,N_11697);
xnor U12023 (N_12023,N_11918,N_11732);
nand U12024 (N_12024,N_11507,N_11854);
or U12025 (N_12025,N_11843,N_11856);
nand U12026 (N_12026,N_11756,N_11792);
xnor U12027 (N_12027,N_11803,N_11691);
nor U12028 (N_12028,N_11682,N_11920);
nand U12029 (N_12029,N_11881,N_11814);
xor U12030 (N_12030,N_11883,N_11670);
nand U12031 (N_12031,N_11571,N_11755);
and U12032 (N_12032,N_11761,N_11717);
nor U12033 (N_12033,N_11719,N_11739);
or U12034 (N_12034,N_11645,N_11746);
and U12035 (N_12035,N_11515,N_11585);
nor U12036 (N_12036,N_11783,N_11500);
and U12037 (N_12037,N_11901,N_11698);
xor U12038 (N_12038,N_11654,N_11871);
nor U12039 (N_12039,N_11572,N_11943);
or U12040 (N_12040,N_11924,N_11927);
and U12041 (N_12041,N_11897,N_11812);
nand U12042 (N_12042,N_11742,N_11636);
or U12043 (N_12043,N_11895,N_11914);
nand U12044 (N_12044,N_11546,N_11708);
nor U12045 (N_12045,N_11974,N_11880);
nand U12046 (N_12046,N_11554,N_11600);
nand U12047 (N_12047,N_11839,N_11539);
or U12048 (N_12048,N_11613,N_11936);
xnor U12049 (N_12049,N_11928,N_11655);
nand U12050 (N_12050,N_11889,N_11774);
xor U12051 (N_12051,N_11775,N_11549);
or U12052 (N_12052,N_11882,N_11648);
nor U12053 (N_12053,N_11830,N_11999);
or U12054 (N_12054,N_11886,N_11751);
nand U12055 (N_12055,N_11521,N_11560);
nor U12056 (N_12056,N_11724,N_11503);
and U12057 (N_12057,N_11797,N_11847);
xor U12058 (N_12058,N_11574,N_11984);
xnor U12059 (N_12059,N_11913,N_11516);
or U12060 (N_12060,N_11911,N_11857);
xor U12061 (N_12061,N_11846,N_11811);
nor U12062 (N_12062,N_11540,N_11603);
nand U12063 (N_12063,N_11606,N_11729);
xor U12064 (N_12064,N_11653,N_11932);
nor U12065 (N_12065,N_11631,N_11799);
xor U12066 (N_12066,N_11707,N_11647);
and U12067 (N_12067,N_11835,N_11673);
nor U12068 (N_12068,N_11931,N_11619);
or U12069 (N_12069,N_11520,N_11782);
or U12070 (N_12070,N_11537,N_11923);
and U12071 (N_12071,N_11510,N_11626);
and U12072 (N_12072,N_11524,N_11747);
nor U12073 (N_12073,N_11872,N_11978);
and U12074 (N_12074,N_11988,N_11579);
nor U12075 (N_12075,N_11942,N_11852);
xor U12076 (N_12076,N_11547,N_11624);
and U12077 (N_12077,N_11837,N_11822);
nor U12078 (N_12078,N_11595,N_11940);
nor U12079 (N_12079,N_11831,N_11874);
xor U12080 (N_12080,N_11987,N_11824);
and U12081 (N_12081,N_11651,N_11778);
or U12082 (N_12082,N_11505,N_11656);
nor U12083 (N_12083,N_11760,N_11829);
xor U12084 (N_12084,N_11602,N_11679);
xnor U12085 (N_12085,N_11850,N_11963);
or U12086 (N_12086,N_11888,N_11855);
nor U12087 (N_12087,N_11637,N_11519);
and U12088 (N_12088,N_11687,N_11966);
nand U12089 (N_12089,N_11623,N_11870);
nand U12090 (N_12090,N_11813,N_11721);
and U12091 (N_12091,N_11965,N_11935);
nand U12092 (N_12092,N_11915,N_11532);
or U12093 (N_12093,N_11596,N_11744);
nand U12094 (N_12094,N_11973,N_11727);
xnor U12095 (N_12095,N_11710,N_11646);
and U12096 (N_12096,N_11536,N_11733);
and U12097 (N_12097,N_11815,N_11849);
and U12098 (N_12098,N_11734,N_11550);
and U12099 (N_12099,N_11950,N_11677);
or U12100 (N_12100,N_11525,N_11684);
and U12101 (N_12101,N_11564,N_11703);
and U12102 (N_12102,N_11757,N_11808);
nor U12103 (N_12103,N_11910,N_11568);
xor U12104 (N_12104,N_11802,N_11501);
nand U12105 (N_12105,N_11894,N_11580);
and U12106 (N_12106,N_11810,N_11930);
and U12107 (N_12107,N_11971,N_11925);
and U12108 (N_12108,N_11904,N_11832);
and U12109 (N_12109,N_11640,N_11630);
xnor U12110 (N_12110,N_11628,N_11907);
or U12111 (N_12111,N_11558,N_11544);
and U12112 (N_12112,N_11581,N_11590);
or U12113 (N_12113,N_11798,N_11593);
or U12114 (N_12114,N_11565,N_11542);
and U12115 (N_12115,N_11868,N_11662);
nor U12116 (N_12116,N_11686,N_11995);
and U12117 (N_12117,N_11641,N_11634);
or U12118 (N_12118,N_11678,N_11534);
xor U12119 (N_12119,N_11842,N_11591);
xnor U12120 (N_12120,N_11681,N_11582);
or U12121 (N_12121,N_11598,N_11526);
nor U12122 (N_12122,N_11644,N_11511);
or U12123 (N_12123,N_11617,N_11776);
or U12124 (N_12124,N_11529,N_11551);
xnor U12125 (N_12125,N_11700,N_11887);
xor U12126 (N_12126,N_11723,N_11779);
nor U12127 (N_12127,N_11658,N_11561);
xor U12128 (N_12128,N_11557,N_11860);
xnor U12129 (N_12129,N_11718,N_11577);
and U12130 (N_12130,N_11789,N_11917);
xor U12131 (N_12131,N_11906,N_11896);
and U12132 (N_12132,N_11938,N_11683);
nor U12133 (N_12133,N_11801,N_11922);
and U12134 (N_12134,N_11699,N_11608);
nor U12135 (N_12135,N_11562,N_11592);
xor U12136 (N_12136,N_11513,N_11676);
or U12137 (N_12137,N_11753,N_11711);
nand U12138 (N_12138,N_11875,N_11517);
and U12139 (N_12139,N_11688,N_11570);
nand U12140 (N_12140,N_11786,N_11749);
nand U12141 (N_12141,N_11956,N_11859);
nand U12142 (N_12142,N_11934,N_11566);
nand U12143 (N_12143,N_11618,N_11530);
nand U12144 (N_12144,N_11518,N_11702);
nand U12145 (N_12145,N_11998,N_11876);
xnor U12146 (N_12146,N_11861,N_11969);
or U12147 (N_12147,N_11765,N_11838);
or U12148 (N_12148,N_11780,N_11997);
and U12149 (N_12149,N_11704,N_11985);
and U12150 (N_12150,N_11899,N_11848);
and U12151 (N_12151,N_11652,N_11863);
nor U12152 (N_12152,N_11773,N_11902);
and U12153 (N_12153,N_11764,N_11639);
or U12154 (N_12154,N_11594,N_11671);
nor U12155 (N_12155,N_11825,N_11944);
nand U12156 (N_12156,N_11826,N_11845);
nand U12157 (N_12157,N_11844,N_11589);
nand U12158 (N_12158,N_11737,N_11772);
nor U12159 (N_12159,N_11919,N_11754);
xor U12160 (N_12160,N_11523,N_11725);
xor U12161 (N_12161,N_11941,N_11862);
nand U12162 (N_12162,N_11840,N_11605);
or U12163 (N_12163,N_11642,N_11615);
and U12164 (N_12164,N_11722,N_11567);
and U12165 (N_12165,N_11970,N_11948);
or U12166 (N_12166,N_11694,N_11946);
or U12167 (N_12167,N_11939,N_11949);
nor U12168 (N_12168,N_11977,N_11893);
and U12169 (N_12169,N_11643,N_11543);
nand U12170 (N_12170,N_11611,N_11533);
and U12171 (N_12171,N_11635,N_11945);
nand U12172 (N_12172,N_11716,N_11576);
nand U12173 (N_12173,N_11759,N_11584);
or U12174 (N_12174,N_11535,N_11884);
or U12175 (N_12175,N_11657,N_11569);
nand U12176 (N_12176,N_11864,N_11794);
nor U12177 (N_12177,N_11841,N_11865);
and U12178 (N_12178,N_11690,N_11877);
or U12179 (N_12179,N_11908,N_11912);
xnor U12180 (N_12180,N_11587,N_11921);
nor U12181 (N_12181,N_11672,N_11980);
nor U12182 (N_12182,N_11714,N_11731);
nor U12183 (N_12183,N_11506,N_11622);
nor U12184 (N_12184,N_11905,N_11752);
nand U12185 (N_12185,N_11762,N_11796);
nand U12186 (N_12186,N_11621,N_11763);
or U12187 (N_12187,N_11620,N_11701);
xor U12188 (N_12188,N_11954,N_11659);
nand U12189 (N_12189,N_11892,N_11819);
nand U12190 (N_12190,N_11720,N_11827);
and U12191 (N_12191,N_11614,N_11604);
xor U12192 (N_12192,N_11770,N_11959);
or U12193 (N_12193,N_11858,N_11586);
or U12194 (N_12194,N_11957,N_11785);
or U12195 (N_12195,N_11578,N_11768);
nor U12196 (N_12196,N_11575,N_11649);
nor U12197 (N_12197,N_11638,N_11715);
nand U12198 (N_12198,N_11929,N_11983);
xnor U12199 (N_12199,N_11748,N_11610);
or U12200 (N_12200,N_11573,N_11504);
or U12201 (N_12201,N_11979,N_11616);
or U12202 (N_12202,N_11736,N_11706);
and U12203 (N_12203,N_11597,N_11633);
nand U12204 (N_12204,N_11952,N_11806);
and U12205 (N_12205,N_11607,N_11527);
or U12206 (N_12206,N_11851,N_11730);
xnor U12207 (N_12207,N_11964,N_11879);
nand U12208 (N_12208,N_11758,N_11947);
or U12209 (N_12209,N_11728,N_11991);
and U12210 (N_12210,N_11583,N_11820);
nand U12211 (N_12211,N_11989,N_11961);
nand U12212 (N_12212,N_11689,N_11559);
nand U12213 (N_12213,N_11563,N_11828);
nor U12214 (N_12214,N_11692,N_11777);
nand U12215 (N_12215,N_11981,N_11834);
nand U12216 (N_12216,N_11674,N_11807);
and U12217 (N_12217,N_11869,N_11866);
and U12218 (N_12218,N_11781,N_11823);
and U12219 (N_12219,N_11972,N_11508);
nand U12220 (N_12220,N_11743,N_11509);
nand U12221 (N_12221,N_11788,N_11502);
nand U12222 (N_12222,N_11867,N_11675);
or U12223 (N_12223,N_11873,N_11986);
nor U12224 (N_12224,N_11685,N_11609);
or U12225 (N_12225,N_11996,N_11903);
or U12226 (N_12226,N_11990,N_11955);
nand U12227 (N_12227,N_11556,N_11660);
xor U12228 (N_12228,N_11933,N_11712);
nand U12229 (N_12229,N_11878,N_11836);
or U12230 (N_12230,N_11599,N_11666);
or U12231 (N_12231,N_11741,N_11695);
nand U12232 (N_12232,N_11909,N_11953);
nand U12233 (N_12233,N_11552,N_11891);
nand U12234 (N_12234,N_11627,N_11790);
and U12235 (N_12235,N_11735,N_11612);
nand U12236 (N_12236,N_11885,N_11726);
nand U12237 (N_12237,N_11522,N_11709);
and U12238 (N_12238,N_11975,N_11937);
nand U12239 (N_12239,N_11553,N_11968);
nor U12240 (N_12240,N_11962,N_11601);
and U12241 (N_12241,N_11632,N_11900);
or U12242 (N_12242,N_11791,N_11816);
nand U12243 (N_12243,N_11680,N_11696);
or U12244 (N_12244,N_11958,N_11665);
and U12245 (N_12245,N_11669,N_11853);
nand U12246 (N_12246,N_11793,N_11767);
or U12247 (N_12247,N_11740,N_11821);
nor U12248 (N_12248,N_11545,N_11951);
xor U12249 (N_12249,N_11926,N_11833);
and U12250 (N_12250,N_11660,N_11983);
nor U12251 (N_12251,N_11646,N_11871);
nor U12252 (N_12252,N_11785,N_11844);
nand U12253 (N_12253,N_11978,N_11651);
or U12254 (N_12254,N_11562,N_11972);
nand U12255 (N_12255,N_11516,N_11986);
or U12256 (N_12256,N_11674,N_11778);
xnor U12257 (N_12257,N_11701,N_11958);
or U12258 (N_12258,N_11882,N_11831);
or U12259 (N_12259,N_11706,N_11560);
or U12260 (N_12260,N_11606,N_11933);
and U12261 (N_12261,N_11957,N_11606);
nand U12262 (N_12262,N_11756,N_11619);
nor U12263 (N_12263,N_11871,N_11509);
or U12264 (N_12264,N_11871,N_11686);
xnor U12265 (N_12265,N_11588,N_11950);
nand U12266 (N_12266,N_11643,N_11686);
nand U12267 (N_12267,N_11874,N_11531);
xnor U12268 (N_12268,N_11945,N_11986);
and U12269 (N_12269,N_11993,N_11652);
nand U12270 (N_12270,N_11826,N_11509);
nor U12271 (N_12271,N_11886,N_11808);
and U12272 (N_12272,N_11729,N_11909);
and U12273 (N_12273,N_11938,N_11646);
or U12274 (N_12274,N_11959,N_11802);
xnor U12275 (N_12275,N_11841,N_11640);
xor U12276 (N_12276,N_11637,N_11960);
nor U12277 (N_12277,N_11854,N_11907);
and U12278 (N_12278,N_11528,N_11834);
nand U12279 (N_12279,N_11666,N_11765);
or U12280 (N_12280,N_11911,N_11761);
nor U12281 (N_12281,N_11722,N_11794);
and U12282 (N_12282,N_11821,N_11581);
nand U12283 (N_12283,N_11892,N_11587);
nand U12284 (N_12284,N_11942,N_11719);
or U12285 (N_12285,N_11797,N_11811);
or U12286 (N_12286,N_11788,N_11812);
nor U12287 (N_12287,N_11845,N_11795);
or U12288 (N_12288,N_11513,N_11541);
or U12289 (N_12289,N_11939,N_11510);
and U12290 (N_12290,N_11617,N_11637);
and U12291 (N_12291,N_11722,N_11882);
nor U12292 (N_12292,N_11662,N_11998);
or U12293 (N_12293,N_11776,N_11927);
nor U12294 (N_12294,N_11600,N_11951);
xor U12295 (N_12295,N_11588,N_11922);
or U12296 (N_12296,N_11511,N_11741);
nand U12297 (N_12297,N_11884,N_11893);
and U12298 (N_12298,N_11597,N_11956);
nor U12299 (N_12299,N_11840,N_11945);
and U12300 (N_12300,N_11775,N_11865);
xor U12301 (N_12301,N_11781,N_11876);
or U12302 (N_12302,N_11851,N_11517);
or U12303 (N_12303,N_11790,N_11987);
and U12304 (N_12304,N_11553,N_11692);
and U12305 (N_12305,N_11823,N_11961);
or U12306 (N_12306,N_11743,N_11983);
or U12307 (N_12307,N_11711,N_11528);
nand U12308 (N_12308,N_11569,N_11848);
xnor U12309 (N_12309,N_11736,N_11756);
nor U12310 (N_12310,N_11749,N_11882);
xor U12311 (N_12311,N_11629,N_11754);
xor U12312 (N_12312,N_11889,N_11772);
and U12313 (N_12313,N_11721,N_11891);
and U12314 (N_12314,N_11858,N_11525);
or U12315 (N_12315,N_11510,N_11529);
nand U12316 (N_12316,N_11603,N_11591);
and U12317 (N_12317,N_11560,N_11984);
and U12318 (N_12318,N_11954,N_11871);
or U12319 (N_12319,N_11635,N_11781);
or U12320 (N_12320,N_11999,N_11977);
nand U12321 (N_12321,N_11966,N_11683);
or U12322 (N_12322,N_11713,N_11597);
xnor U12323 (N_12323,N_11655,N_11519);
and U12324 (N_12324,N_11601,N_11594);
nand U12325 (N_12325,N_11975,N_11797);
nand U12326 (N_12326,N_11609,N_11785);
nor U12327 (N_12327,N_11791,N_11932);
and U12328 (N_12328,N_11997,N_11523);
xor U12329 (N_12329,N_11966,N_11558);
nand U12330 (N_12330,N_11742,N_11810);
or U12331 (N_12331,N_11605,N_11992);
or U12332 (N_12332,N_11770,N_11792);
nand U12333 (N_12333,N_11927,N_11632);
or U12334 (N_12334,N_11957,N_11737);
nand U12335 (N_12335,N_11510,N_11616);
or U12336 (N_12336,N_11625,N_11777);
xor U12337 (N_12337,N_11742,N_11717);
nand U12338 (N_12338,N_11762,N_11830);
nor U12339 (N_12339,N_11616,N_11731);
nor U12340 (N_12340,N_11630,N_11806);
or U12341 (N_12341,N_11597,N_11587);
or U12342 (N_12342,N_11661,N_11997);
nand U12343 (N_12343,N_11764,N_11931);
and U12344 (N_12344,N_11908,N_11797);
or U12345 (N_12345,N_11988,N_11962);
nor U12346 (N_12346,N_11614,N_11695);
nand U12347 (N_12347,N_11757,N_11619);
xnor U12348 (N_12348,N_11837,N_11970);
or U12349 (N_12349,N_11863,N_11627);
xor U12350 (N_12350,N_11609,N_11969);
nor U12351 (N_12351,N_11848,N_11826);
xnor U12352 (N_12352,N_11961,N_11986);
nor U12353 (N_12353,N_11823,N_11567);
xnor U12354 (N_12354,N_11821,N_11657);
nor U12355 (N_12355,N_11971,N_11603);
nor U12356 (N_12356,N_11918,N_11603);
or U12357 (N_12357,N_11974,N_11566);
xnor U12358 (N_12358,N_11934,N_11931);
nor U12359 (N_12359,N_11841,N_11592);
nor U12360 (N_12360,N_11509,N_11903);
nor U12361 (N_12361,N_11874,N_11919);
xnor U12362 (N_12362,N_11797,N_11994);
or U12363 (N_12363,N_11655,N_11755);
or U12364 (N_12364,N_11660,N_11641);
nand U12365 (N_12365,N_11546,N_11713);
nand U12366 (N_12366,N_11791,N_11684);
xnor U12367 (N_12367,N_11653,N_11651);
nand U12368 (N_12368,N_11846,N_11856);
xnor U12369 (N_12369,N_11710,N_11982);
nand U12370 (N_12370,N_11877,N_11935);
nor U12371 (N_12371,N_11882,N_11700);
nor U12372 (N_12372,N_11705,N_11509);
and U12373 (N_12373,N_11881,N_11722);
and U12374 (N_12374,N_11531,N_11984);
nor U12375 (N_12375,N_11507,N_11997);
xor U12376 (N_12376,N_11577,N_11534);
nor U12377 (N_12377,N_11675,N_11617);
nand U12378 (N_12378,N_11713,N_11921);
and U12379 (N_12379,N_11690,N_11673);
and U12380 (N_12380,N_11557,N_11637);
xor U12381 (N_12381,N_11718,N_11978);
nand U12382 (N_12382,N_11517,N_11631);
xnor U12383 (N_12383,N_11656,N_11686);
and U12384 (N_12384,N_11820,N_11633);
nand U12385 (N_12385,N_11995,N_11921);
or U12386 (N_12386,N_11904,N_11683);
or U12387 (N_12387,N_11684,N_11733);
and U12388 (N_12388,N_11816,N_11985);
and U12389 (N_12389,N_11926,N_11823);
nor U12390 (N_12390,N_11679,N_11575);
nand U12391 (N_12391,N_11580,N_11926);
nand U12392 (N_12392,N_11613,N_11573);
nor U12393 (N_12393,N_11626,N_11819);
nand U12394 (N_12394,N_11886,N_11999);
or U12395 (N_12395,N_11792,N_11871);
or U12396 (N_12396,N_11527,N_11917);
or U12397 (N_12397,N_11543,N_11776);
or U12398 (N_12398,N_11794,N_11648);
and U12399 (N_12399,N_11957,N_11956);
and U12400 (N_12400,N_11701,N_11799);
nor U12401 (N_12401,N_11953,N_11516);
nand U12402 (N_12402,N_11586,N_11934);
xor U12403 (N_12403,N_11715,N_11698);
nand U12404 (N_12404,N_11806,N_11626);
nand U12405 (N_12405,N_11836,N_11973);
xor U12406 (N_12406,N_11702,N_11879);
nor U12407 (N_12407,N_11888,N_11973);
nand U12408 (N_12408,N_11865,N_11507);
or U12409 (N_12409,N_11516,N_11590);
or U12410 (N_12410,N_11687,N_11523);
and U12411 (N_12411,N_11739,N_11701);
and U12412 (N_12412,N_11680,N_11571);
xor U12413 (N_12413,N_11659,N_11762);
nor U12414 (N_12414,N_11709,N_11959);
and U12415 (N_12415,N_11612,N_11698);
nand U12416 (N_12416,N_11717,N_11867);
and U12417 (N_12417,N_11907,N_11503);
or U12418 (N_12418,N_11833,N_11678);
and U12419 (N_12419,N_11915,N_11807);
nor U12420 (N_12420,N_11653,N_11709);
nor U12421 (N_12421,N_11530,N_11823);
nor U12422 (N_12422,N_11920,N_11516);
or U12423 (N_12423,N_11642,N_11965);
nand U12424 (N_12424,N_11783,N_11681);
and U12425 (N_12425,N_11862,N_11607);
xor U12426 (N_12426,N_11706,N_11760);
xor U12427 (N_12427,N_11923,N_11931);
nand U12428 (N_12428,N_11546,N_11940);
and U12429 (N_12429,N_11907,N_11597);
or U12430 (N_12430,N_11767,N_11557);
or U12431 (N_12431,N_11920,N_11730);
and U12432 (N_12432,N_11913,N_11922);
nor U12433 (N_12433,N_11561,N_11507);
or U12434 (N_12434,N_11963,N_11630);
or U12435 (N_12435,N_11829,N_11917);
or U12436 (N_12436,N_11642,N_11549);
nand U12437 (N_12437,N_11505,N_11709);
and U12438 (N_12438,N_11762,N_11637);
nor U12439 (N_12439,N_11828,N_11834);
nand U12440 (N_12440,N_11879,N_11747);
xor U12441 (N_12441,N_11917,N_11592);
and U12442 (N_12442,N_11956,N_11524);
nand U12443 (N_12443,N_11969,N_11860);
nor U12444 (N_12444,N_11676,N_11989);
and U12445 (N_12445,N_11568,N_11726);
or U12446 (N_12446,N_11949,N_11801);
nor U12447 (N_12447,N_11964,N_11623);
xnor U12448 (N_12448,N_11887,N_11582);
or U12449 (N_12449,N_11633,N_11628);
or U12450 (N_12450,N_11633,N_11595);
xor U12451 (N_12451,N_11682,N_11915);
nor U12452 (N_12452,N_11902,N_11760);
xor U12453 (N_12453,N_11780,N_11784);
xor U12454 (N_12454,N_11920,N_11699);
nand U12455 (N_12455,N_11884,N_11965);
nand U12456 (N_12456,N_11957,N_11671);
or U12457 (N_12457,N_11876,N_11970);
or U12458 (N_12458,N_11813,N_11826);
or U12459 (N_12459,N_11689,N_11737);
nand U12460 (N_12460,N_11982,N_11659);
nand U12461 (N_12461,N_11523,N_11701);
nand U12462 (N_12462,N_11915,N_11848);
nor U12463 (N_12463,N_11695,N_11768);
nand U12464 (N_12464,N_11584,N_11711);
and U12465 (N_12465,N_11500,N_11895);
nand U12466 (N_12466,N_11908,N_11800);
and U12467 (N_12467,N_11893,N_11907);
nor U12468 (N_12468,N_11609,N_11756);
xor U12469 (N_12469,N_11886,N_11843);
nor U12470 (N_12470,N_11916,N_11756);
and U12471 (N_12471,N_11811,N_11832);
or U12472 (N_12472,N_11607,N_11975);
and U12473 (N_12473,N_11991,N_11596);
and U12474 (N_12474,N_11730,N_11601);
and U12475 (N_12475,N_11646,N_11808);
and U12476 (N_12476,N_11680,N_11873);
or U12477 (N_12477,N_11945,N_11666);
nor U12478 (N_12478,N_11973,N_11500);
xnor U12479 (N_12479,N_11919,N_11932);
or U12480 (N_12480,N_11699,N_11523);
nand U12481 (N_12481,N_11833,N_11640);
or U12482 (N_12482,N_11864,N_11960);
xnor U12483 (N_12483,N_11977,N_11749);
or U12484 (N_12484,N_11920,N_11504);
xnor U12485 (N_12485,N_11776,N_11745);
nand U12486 (N_12486,N_11615,N_11515);
xor U12487 (N_12487,N_11934,N_11535);
xnor U12488 (N_12488,N_11951,N_11670);
nand U12489 (N_12489,N_11590,N_11787);
nor U12490 (N_12490,N_11580,N_11504);
nor U12491 (N_12491,N_11786,N_11935);
xor U12492 (N_12492,N_11725,N_11769);
or U12493 (N_12493,N_11694,N_11992);
and U12494 (N_12494,N_11759,N_11787);
nand U12495 (N_12495,N_11606,N_11884);
or U12496 (N_12496,N_11507,N_11696);
and U12497 (N_12497,N_11913,N_11566);
and U12498 (N_12498,N_11515,N_11663);
xnor U12499 (N_12499,N_11627,N_11537);
and U12500 (N_12500,N_12056,N_12170);
nor U12501 (N_12501,N_12120,N_12353);
and U12502 (N_12502,N_12036,N_12002);
nor U12503 (N_12503,N_12351,N_12319);
nor U12504 (N_12504,N_12160,N_12289);
and U12505 (N_12505,N_12206,N_12414);
nor U12506 (N_12506,N_12010,N_12122);
nand U12507 (N_12507,N_12069,N_12374);
nand U12508 (N_12508,N_12118,N_12349);
xor U12509 (N_12509,N_12078,N_12057);
nor U12510 (N_12510,N_12202,N_12434);
and U12511 (N_12511,N_12427,N_12464);
nand U12512 (N_12512,N_12014,N_12305);
or U12513 (N_12513,N_12108,N_12273);
nor U12514 (N_12514,N_12035,N_12176);
and U12515 (N_12515,N_12405,N_12342);
nor U12516 (N_12516,N_12263,N_12450);
and U12517 (N_12517,N_12456,N_12309);
and U12518 (N_12518,N_12300,N_12062);
or U12519 (N_12519,N_12214,N_12378);
and U12520 (N_12520,N_12210,N_12113);
nand U12521 (N_12521,N_12320,N_12334);
nand U12522 (N_12522,N_12071,N_12333);
nor U12523 (N_12523,N_12100,N_12163);
xor U12524 (N_12524,N_12147,N_12257);
nand U12525 (N_12525,N_12497,N_12087);
or U12526 (N_12526,N_12086,N_12447);
and U12527 (N_12527,N_12322,N_12045);
nand U12528 (N_12528,N_12271,N_12034);
or U12529 (N_12529,N_12357,N_12454);
or U12530 (N_12530,N_12261,N_12395);
nor U12531 (N_12531,N_12194,N_12294);
or U12532 (N_12532,N_12241,N_12193);
xor U12533 (N_12533,N_12117,N_12156);
nand U12534 (N_12534,N_12327,N_12407);
nand U12535 (N_12535,N_12252,N_12144);
and U12536 (N_12536,N_12483,N_12268);
xnor U12537 (N_12537,N_12188,N_12097);
and U12538 (N_12538,N_12204,N_12417);
nor U12539 (N_12539,N_12197,N_12164);
and U12540 (N_12540,N_12362,N_12475);
xnor U12541 (N_12541,N_12031,N_12138);
and U12542 (N_12542,N_12123,N_12481);
nand U12543 (N_12543,N_12020,N_12493);
or U12544 (N_12544,N_12077,N_12376);
nor U12545 (N_12545,N_12179,N_12452);
nand U12546 (N_12546,N_12393,N_12114);
nor U12547 (N_12547,N_12477,N_12006);
nand U12548 (N_12548,N_12043,N_12330);
or U12549 (N_12549,N_12404,N_12207);
nor U12550 (N_12550,N_12391,N_12367);
nor U12551 (N_12551,N_12083,N_12223);
xor U12552 (N_12552,N_12239,N_12266);
xor U12553 (N_12553,N_12005,N_12159);
xnor U12554 (N_12554,N_12458,N_12343);
nor U12555 (N_12555,N_12152,N_12496);
xnor U12556 (N_12556,N_12486,N_12172);
nand U12557 (N_12557,N_12396,N_12335);
and U12558 (N_12558,N_12431,N_12449);
nand U12559 (N_12559,N_12368,N_12121);
nor U12560 (N_12560,N_12430,N_12386);
and U12561 (N_12561,N_12130,N_12242);
nor U12562 (N_12562,N_12403,N_12480);
xnor U12563 (N_12563,N_12438,N_12093);
and U12564 (N_12564,N_12084,N_12004);
xnor U12565 (N_12565,N_12303,N_12279);
xor U12566 (N_12566,N_12366,N_12371);
or U12567 (N_12567,N_12253,N_12285);
xnor U12568 (N_12568,N_12418,N_12240);
and U12569 (N_12569,N_12324,N_12135);
nor U12570 (N_12570,N_12140,N_12401);
or U12571 (N_12571,N_12095,N_12375);
and U12572 (N_12572,N_12074,N_12192);
nand U12573 (N_12573,N_12054,N_12321);
xor U12574 (N_12574,N_12247,N_12316);
xnor U12575 (N_12575,N_12498,N_12021);
xor U12576 (N_12576,N_12165,N_12145);
nand U12577 (N_12577,N_12220,N_12415);
or U12578 (N_12578,N_12402,N_12384);
nand U12579 (N_12579,N_12103,N_12180);
nor U12580 (N_12580,N_12389,N_12030);
nor U12581 (N_12581,N_12262,N_12166);
and U12582 (N_12582,N_12275,N_12260);
nand U12583 (N_12583,N_12025,N_12090);
or U12584 (N_12584,N_12280,N_12420);
nand U12585 (N_12585,N_12104,N_12133);
nor U12586 (N_12586,N_12479,N_12162);
nand U12587 (N_12587,N_12015,N_12345);
nand U12588 (N_12588,N_12255,N_12284);
and U12589 (N_12589,N_12124,N_12151);
or U12590 (N_12590,N_12258,N_12428);
nand U12591 (N_12591,N_12238,N_12363);
and U12592 (N_12592,N_12058,N_12317);
or U12593 (N_12593,N_12463,N_12047);
and U12594 (N_12594,N_12492,N_12484);
xnor U12595 (N_12595,N_12033,N_12226);
nor U12596 (N_12596,N_12168,N_12313);
xnor U12597 (N_12597,N_12233,N_12296);
nand U12598 (N_12598,N_12178,N_12244);
xor U12599 (N_12599,N_12236,N_12471);
nor U12600 (N_12600,N_12485,N_12410);
and U12601 (N_12601,N_12329,N_12311);
nor U12602 (N_12602,N_12256,N_12196);
nor U12603 (N_12603,N_12198,N_12435);
xnor U12604 (N_12604,N_12234,N_12344);
nand U12605 (N_12605,N_12221,N_12409);
nand U12606 (N_12606,N_12302,N_12448);
or U12607 (N_12607,N_12356,N_12306);
nor U12608 (N_12608,N_12171,N_12237);
or U12609 (N_12609,N_12065,N_12219);
or U12610 (N_12610,N_12441,N_12044);
xor U12611 (N_12611,N_12457,N_12495);
and U12612 (N_12612,N_12169,N_12115);
nor U12613 (N_12613,N_12200,N_12332);
or U12614 (N_12614,N_12224,N_12099);
or U12615 (N_12615,N_12177,N_12009);
nor U12616 (N_12616,N_12397,N_12119);
xnor U12617 (N_12617,N_12143,N_12426);
or U12618 (N_12618,N_12232,N_12173);
nand U12619 (N_12619,N_12195,N_12024);
and U12620 (N_12620,N_12096,N_12336);
xnor U12621 (N_12621,N_12017,N_12229);
and U12622 (N_12622,N_12270,N_12128);
nor U12623 (N_12623,N_12080,N_12063);
and U12624 (N_12624,N_12429,N_12055);
or U12625 (N_12625,N_12149,N_12307);
nand U12626 (N_12626,N_12041,N_12433);
xor U12627 (N_12627,N_12411,N_12267);
or U12628 (N_12628,N_12412,N_12445);
xnor U12629 (N_12629,N_12107,N_12383);
nand U12630 (N_12630,N_12227,N_12315);
or U12631 (N_12631,N_12439,N_12432);
and U12632 (N_12632,N_12364,N_12372);
and U12633 (N_12633,N_12325,N_12476);
and U12634 (N_12634,N_12085,N_12116);
or U12635 (N_12635,N_12112,N_12436);
or U12636 (N_12636,N_12131,N_12191);
xor U12637 (N_12637,N_12174,N_12032);
xor U12638 (N_12638,N_12264,N_12478);
nand U12639 (N_12639,N_12146,N_12444);
nand U12640 (N_12640,N_12455,N_12148);
or U12641 (N_12641,N_12269,N_12385);
xor U12642 (N_12642,N_12295,N_12126);
or U12643 (N_12643,N_12377,N_12379);
nand U12644 (N_12644,N_12446,N_12487);
nor U12645 (N_12645,N_12167,N_12440);
or U12646 (N_12646,N_12408,N_12105);
and U12647 (N_12647,N_12283,N_12060);
xnor U12648 (N_12648,N_12380,N_12046);
or U12649 (N_12649,N_12026,N_12139);
nor U12650 (N_12650,N_12049,N_12051);
nand U12651 (N_12651,N_12340,N_12016);
nand U12652 (N_12652,N_12352,N_12155);
and U12653 (N_12653,N_12469,N_12066);
and U12654 (N_12654,N_12235,N_12109);
and U12655 (N_12655,N_12392,N_12423);
and U12656 (N_12656,N_12079,N_12474);
or U12657 (N_12657,N_12137,N_12212);
nor U12658 (N_12658,N_12248,N_12466);
or U12659 (N_12659,N_12072,N_12354);
nand U12660 (N_12660,N_12125,N_12075);
nand U12661 (N_12661,N_12413,N_12039);
xor U12662 (N_12662,N_12150,N_12259);
nand U12663 (N_12663,N_12136,N_12337);
or U12664 (N_12664,N_12157,N_12208);
xnor U12665 (N_12665,N_12184,N_12462);
nand U12666 (N_12666,N_12488,N_12175);
xor U12667 (N_12667,N_12050,N_12468);
or U12668 (N_12668,N_12365,N_12023);
nor U12669 (N_12669,N_12064,N_12281);
xor U12670 (N_12670,N_12355,N_12394);
nor U12671 (N_12671,N_12425,N_12491);
nor U12672 (N_12672,N_12076,N_12310);
or U12673 (N_12673,N_12048,N_12231);
and U12674 (N_12674,N_12298,N_12052);
nor U12675 (N_12675,N_12018,N_12102);
xnor U12676 (N_12676,N_12217,N_12091);
nor U12677 (N_12677,N_12028,N_12348);
or U12678 (N_12678,N_12001,N_12081);
xnor U12679 (N_12679,N_12350,N_12299);
nor U12680 (N_12680,N_12301,N_12019);
xnor U12681 (N_12681,N_12245,N_12061);
nor U12682 (N_12682,N_12465,N_12129);
or U12683 (N_12683,N_12092,N_12183);
nand U12684 (N_12684,N_12154,N_12181);
or U12685 (N_12685,N_12250,N_12489);
xor U12686 (N_12686,N_12461,N_12153);
xor U12687 (N_12687,N_12228,N_12098);
and U12688 (N_12688,N_12215,N_12276);
nand U12689 (N_12689,N_12007,N_12287);
or U12690 (N_12690,N_12088,N_12127);
nor U12691 (N_12691,N_12490,N_12225);
and U12692 (N_12692,N_12161,N_12040);
nand U12693 (N_12693,N_12453,N_12359);
and U12694 (N_12694,N_12459,N_12347);
nor U12695 (N_12695,N_12400,N_12089);
or U12696 (N_12696,N_12297,N_12361);
and U12697 (N_12697,N_12070,N_12027);
or U12698 (N_12698,N_12338,N_12388);
xor U12699 (N_12699,N_12370,N_12341);
xnor U12700 (N_12700,N_12387,N_12243);
or U12701 (N_12701,N_12042,N_12360);
and U12702 (N_12702,N_12277,N_12282);
xor U12703 (N_12703,N_12209,N_12187);
or U12704 (N_12704,N_12067,N_12059);
nor U12705 (N_12705,N_12470,N_12314);
and U12706 (N_12706,N_12358,N_12205);
and U12707 (N_12707,N_12422,N_12272);
and U12708 (N_12708,N_12201,N_12213);
and U12709 (N_12709,N_12499,N_12111);
or U12710 (N_12710,N_12211,N_12318);
xnor U12711 (N_12711,N_12011,N_12451);
nor U12712 (N_12712,N_12094,N_12460);
nand U12713 (N_12713,N_12421,N_12382);
xnor U12714 (N_12714,N_12186,N_12278);
xnor U12715 (N_12715,N_12199,N_12101);
xor U12716 (N_12716,N_12472,N_12399);
xnor U12717 (N_12717,N_12323,N_12251);
nand U12718 (N_12718,N_12290,N_12182);
or U12719 (N_12719,N_12189,N_12312);
or U12720 (N_12720,N_12082,N_12106);
nand U12721 (N_12721,N_12473,N_12142);
and U12722 (N_12722,N_12398,N_12346);
nor U12723 (N_12723,N_12286,N_12216);
and U12724 (N_12724,N_12293,N_12230);
xnor U12725 (N_12725,N_12373,N_12029);
nor U12726 (N_12726,N_12288,N_12158);
or U12727 (N_12727,N_12308,N_12406);
or U12728 (N_12728,N_12000,N_12482);
nor U12729 (N_12729,N_12274,N_12022);
nand U12730 (N_12730,N_12037,N_12190);
and U12731 (N_12731,N_12424,N_12218);
and U12732 (N_12732,N_12132,N_12328);
xnor U12733 (N_12733,N_12249,N_12437);
nand U12734 (N_12734,N_12339,N_12246);
or U12735 (N_12735,N_12008,N_12013);
or U12736 (N_12736,N_12265,N_12073);
nor U12737 (N_12737,N_12443,N_12416);
or U12738 (N_12738,N_12442,N_12141);
xnor U12739 (N_12739,N_12003,N_12012);
and U12740 (N_12740,N_12291,N_12369);
nand U12741 (N_12741,N_12053,N_12304);
xnor U12742 (N_12742,N_12134,N_12203);
and U12743 (N_12743,N_12292,N_12326);
nor U12744 (N_12744,N_12419,N_12110);
nor U12745 (N_12745,N_12068,N_12494);
xor U12746 (N_12746,N_12222,N_12185);
nor U12747 (N_12747,N_12038,N_12331);
nand U12748 (N_12748,N_12254,N_12390);
or U12749 (N_12749,N_12381,N_12467);
xor U12750 (N_12750,N_12162,N_12047);
nand U12751 (N_12751,N_12043,N_12364);
and U12752 (N_12752,N_12086,N_12193);
nor U12753 (N_12753,N_12060,N_12438);
nand U12754 (N_12754,N_12044,N_12249);
nand U12755 (N_12755,N_12351,N_12330);
and U12756 (N_12756,N_12350,N_12314);
and U12757 (N_12757,N_12204,N_12423);
and U12758 (N_12758,N_12066,N_12176);
or U12759 (N_12759,N_12181,N_12079);
and U12760 (N_12760,N_12203,N_12020);
nor U12761 (N_12761,N_12189,N_12296);
nor U12762 (N_12762,N_12375,N_12204);
or U12763 (N_12763,N_12205,N_12153);
nor U12764 (N_12764,N_12493,N_12034);
xor U12765 (N_12765,N_12161,N_12230);
or U12766 (N_12766,N_12276,N_12052);
xnor U12767 (N_12767,N_12145,N_12395);
nand U12768 (N_12768,N_12299,N_12108);
and U12769 (N_12769,N_12314,N_12169);
nand U12770 (N_12770,N_12479,N_12425);
xnor U12771 (N_12771,N_12084,N_12104);
or U12772 (N_12772,N_12291,N_12268);
or U12773 (N_12773,N_12419,N_12145);
xnor U12774 (N_12774,N_12468,N_12254);
nor U12775 (N_12775,N_12319,N_12248);
nand U12776 (N_12776,N_12123,N_12008);
or U12777 (N_12777,N_12459,N_12350);
nor U12778 (N_12778,N_12144,N_12433);
nor U12779 (N_12779,N_12325,N_12089);
and U12780 (N_12780,N_12370,N_12158);
xor U12781 (N_12781,N_12220,N_12317);
nand U12782 (N_12782,N_12443,N_12085);
or U12783 (N_12783,N_12480,N_12156);
nand U12784 (N_12784,N_12293,N_12371);
nand U12785 (N_12785,N_12033,N_12026);
or U12786 (N_12786,N_12084,N_12389);
or U12787 (N_12787,N_12388,N_12146);
nand U12788 (N_12788,N_12159,N_12248);
xnor U12789 (N_12789,N_12225,N_12389);
xor U12790 (N_12790,N_12022,N_12157);
nand U12791 (N_12791,N_12472,N_12066);
and U12792 (N_12792,N_12011,N_12136);
xor U12793 (N_12793,N_12368,N_12396);
and U12794 (N_12794,N_12438,N_12441);
nand U12795 (N_12795,N_12156,N_12099);
nand U12796 (N_12796,N_12125,N_12449);
xnor U12797 (N_12797,N_12195,N_12170);
and U12798 (N_12798,N_12075,N_12484);
or U12799 (N_12799,N_12394,N_12229);
and U12800 (N_12800,N_12376,N_12205);
nor U12801 (N_12801,N_12340,N_12296);
nor U12802 (N_12802,N_12359,N_12296);
and U12803 (N_12803,N_12193,N_12068);
or U12804 (N_12804,N_12314,N_12209);
or U12805 (N_12805,N_12384,N_12106);
and U12806 (N_12806,N_12387,N_12226);
nand U12807 (N_12807,N_12360,N_12462);
xor U12808 (N_12808,N_12445,N_12382);
nand U12809 (N_12809,N_12090,N_12139);
or U12810 (N_12810,N_12085,N_12454);
xor U12811 (N_12811,N_12359,N_12274);
and U12812 (N_12812,N_12271,N_12042);
nand U12813 (N_12813,N_12209,N_12355);
nand U12814 (N_12814,N_12012,N_12292);
or U12815 (N_12815,N_12447,N_12037);
nand U12816 (N_12816,N_12294,N_12041);
xnor U12817 (N_12817,N_12175,N_12363);
nor U12818 (N_12818,N_12300,N_12362);
nor U12819 (N_12819,N_12336,N_12148);
and U12820 (N_12820,N_12496,N_12313);
xnor U12821 (N_12821,N_12393,N_12097);
nand U12822 (N_12822,N_12243,N_12351);
nor U12823 (N_12823,N_12068,N_12251);
and U12824 (N_12824,N_12026,N_12330);
and U12825 (N_12825,N_12093,N_12028);
or U12826 (N_12826,N_12346,N_12033);
nor U12827 (N_12827,N_12265,N_12070);
nand U12828 (N_12828,N_12407,N_12091);
or U12829 (N_12829,N_12435,N_12117);
xor U12830 (N_12830,N_12275,N_12362);
nand U12831 (N_12831,N_12269,N_12163);
xnor U12832 (N_12832,N_12421,N_12379);
nand U12833 (N_12833,N_12420,N_12262);
xor U12834 (N_12834,N_12464,N_12362);
or U12835 (N_12835,N_12429,N_12054);
nor U12836 (N_12836,N_12216,N_12429);
and U12837 (N_12837,N_12480,N_12341);
and U12838 (N_12838,N_12160,N_12158);
nor U12839 (N_12839,N_12111,N_12452);
xnor U12840 (N_12840,N_12354,N_12022);
xnor U12841 (N_12841,N_12075,N_12239);
nand U12842 (N_12842,N_12494,N_12412);
and U12843 (N_12843,N_12475,N_12329);
xnor U12844 (N_12844,N_12112,N_12170);
xnor U12845 (N_12845,N_12142,N_12485);
nor U12846 (N_12846,N_12396,N_12131);
and U12847 (N_12847,N_12125,N_12264);
nand U12848 (N_12848,N_12459,N_12464);
xnor U12849 (N_12849,N_12431,N_12451);
xor U12850 (N_12850,N_12066,N_12089);
xor U12851 (N_12851,N_12088,N_12397);
and U12852 (N_12852,N_12348,N_12042);
or U12853 (N_12853,N_12300,N_12196);
or U12854 (N_12854,N_12137,N_12278);
or U12855 (N_12855,N_12165,N_12090);
or U12856 (N_12856,N_12359,N_12435);
or U12857 (N_12857,N_12491,N_12185);
and U12858 (N_12858,N_12237,N_12388);
xor U12859 (N_12859,N_12493,N_12498);
and U12860 (N_12860,N_12061,N_12410);
nor U12861 (N_12861,N_12331,N_12039);
or U12862 (N_12862,N_12083,N_12442);
or U12863 (N_12863,N_12398,N_12304);
nand U12864 (N_12864,N_12108,N_12017);
nor U12865 (N_12865,N_12240,N_12344);
nor U12866 (N_12866,N_12126,N_12330);
xor U12867 (N_12867,N_12471,N_12250);
xnor U12868 (N_12868,N_12389,N_12190);
or U12869 (N_12869,N_12489,N_12456);
xor U12870 (N_12870,N_12443,N_12330);
xnor U12871 (N_12871,N_12250,N_12499);
xnor U12872 (N_12872,N_12083,N_12278);
xor U12873 (N_12873,N_12073,N_12449);
nor U12874 (N_12874,N_12319,N_12142);
nand U12875 (N_12875,N_12124,N_12294);
xor U12876 (N_12876,N_12461,N_12413);
or U12877 (N_12877,N_12113,N_12311);
nor U12878 (N_12878,N_12164,N_12049);
xor U12879 (N_12879,N_12329,N_12319);
or U12880 (N_12880,N_12155,N_12350);
nor U12881 (N_12881,N_12021,N_12435);
or U12882 (N_12882,N_12260,N_12137);
nand U12883 (N_12883,N_12315,N_12414);
and U12884 (N_12884,N_12125,N_12215);
nand U12885 (N_12885,N_12041,N_12200);
and U12886 (N_12886,N_12044,N_12284);
nor U12887 (N_12887,N_12343,N_12473);
xnor U12888 (N_12888,N_12141,N_12090);
nor U12889 (N_12889,N_12349,N_12065);
nor U12890 (N_12890,N_12356,N_12091);
or U12891 (N_12891,N_12330,N_12312);
xor U12892 (N_12892,N_12483,N_12132);
xor U12893 (N_12893,N_12016,N_12276);
nor U12894 (N_12894,N_12205,N_12027);
xor U12895 (N_12895,N_12133,N_12335);
nor U12896 (N_12896,N_12134,N_12462);
nor U12897 (N_12897,N_12449,N_12286);
nand U12898 (N_12898,N_12189,N_12079);
nand U12899 (N_12899,N_12033,N_12063);
nor U12900 (N_12900,N_12332,N_12069);
xnor U12901 (N_12901,N_12174,N_12087);
nor U12902 (N_12902,N_12170,N_12458);
and U12903 (N_12903,N_12139,N_12361);
nor U12904 (N_12904,N_12400,N_12006);
nor U12905 (N_12905,N_12116,N_12065);
nand U12906 (N_12906,N_12269,N_12472);
nor U12907 (N_12907,N_12065,N_12462);
or U12908 (N_12908,N_12211,N_12314);
nor U12909 (N_12909,N_12477,N_12286);
nand U12910 (N_12910,N_12243,N_12141);
nor U12911 (N_12911,N_12230,N_12435);
nor U12912 (N_12912,N_12224,N_12404);
and U12913 (N_12913,N_12471,N_12184);
or U12914 (N_12914,N_12077,N_12038);
nor U12915 (N_12915,N_12149,N_12276);
or U12916 (N_12916,N_12190,N_12371);
xnor U12917 (N_12917,N_12048,N_12465);
and U12918 (N_12918,N_12319,N_12114);
nand U12919 (N_12919,N_12309,N_12405);
and U12920 (N_12920,N_12222,N_12127);
nor U12921 (N_12921,N_12309,N_12238);
xnor U12922 (N_12922,N_12080,N_12222);
or U12923 (N_12923,N_12248,N_12264);
nand U12924 (N_12924,N_12384,N_12141);
or U12925 (N_12925,N_12060,N_12416);
xnor U12926 (N_12926,N_12040,N_12419);
and U12927 (N_12927,N_12018,N_12015);
nand U12928 (N_12928,N_12251,N_12020);
xor U12929 (N_12929,N_12497,N_12013);
nor U12930 (N_12930,N_12389,N_12361);
xnor U12931 (N_12931,N_12397,N_12127);
nand U12932 (N_12932,N_12440,N_12208);
or U12933 (N_12933,N_12198,N_12441);
and U12934 (N_12934,N_12418,N_12064);
nand U12935 (N_12935,N_12475,N_12343);
or U12936 (N_12936,N_12480,N_12145);
or U12937 (N_12937,N_12073,N_12308);
nor U12938 (N_12938,N_12307,N_12442);
and U12939 (N_12939,N_12413,N_12147);
xor U12940 (N_12940,N_12138,N_12219);
or U12941 (N_12941,N_12453,N_12043);
nand U12942 (N_12942,N_12268,N_12290);
or U12943 (N_12943,N_12460,N_12317);
xnor U12944 (N_12944,N_12337,N_12022);
nand U12945 (N_12945,N_12009,N_12031);
nand U12946 (N_12946,N_12148,N_12384);
and U12947 (N_12947,N_12478,N_12240);
nand U12948 (N_12948,N_12407,N_12422);
or U12949 (N_12949,N_12054,N_12346);
nand U12950 (N_12950,N_12130,N_12138);
nor U12951 (N_12951,N_12232,N_12382);
xnor U12952 (N_12952,N_12132,N_12145);
nand U12953 (N_12953,N_12414,N_12342);
xnor U12954 (N_12954,N_12202,N_12293);
or U12955 (N_12955,N_12069,N_12082);
or U12956 (N_12956,N_12246,N_12209);
or U12957 (N_12957,N_12353,N_12327);
and U12958 (N_12958,N_12470,N_12143);
nor U12959 (N_12959,N_12269,N_12307);
xnor U12960 (N_12960,N_12040,N_12411);
nor U12961 (N_12961,N_12179,N_12321);
xor U12962 (N_12962,N_12257,N_12368);
and U12963 (N_12963,N_12037,N_12107);
nor U12964 (N_12964,N_12370,N_12282);
xor U12965 (N_12965,N_12345,N_12478);
nand U12966 (N_12966,N_12114,N_12469);
and U12967 (N_12967,N_12460,N_12283);
or U12968 (N_12968,N_12326,N_12323);
nor U12969 (N_12969,N_12049,N_12266);
and U12970 (N_12970,N_12298,N_12280);
nand U12971 (N_12971,N_12087,N_12399);
xor U12972 (N_12972,N_12310,N_12211);
or U12973 (N_12973,N_12002,N_12335);
xor U12974 (N_12974,N_12268,N_12187);
xor U12975 (N_12975,N_12215,N_12390);
and U12976 (N_12976,N_12136,N_12196);
or U12977 (N_12977,N_12338,N_12263);
nor U12978 (N_12978,N_12386,N_12456);
or U12979 (N_12979,N_12342,N_12226);
nand U12980 (N_12980,N_12365,N_12142);
nor U12981 (N_12981,N_12360,N_12451);
or U12982 (N_12982,N_12457,N_12480);
or U12983 (N_12983,N_12230,N_12364);
nor U12984 (N_12984,N_12323,N_12204);
nand U12985 (N_12985,N_12378,N_12064);
nand U12986 (N_12986,N_12450,N_12328);
nand U12987 (N_12987,N_12095,N_12055);
and U12988 (N_12988,N_12297,N_12415);
nor U12989 (N_12989,N_12408,N_12173);
or U12990 (N_12990,N_12093,N_12171);
xor U12991 (N_12991,N_12053,N_12485);
and U12992 (N_12992,N_12141,N_12146);
or U12993 (N_12993,N_12452,N_12445);
nor U12994 (N_12994,N_12205,N_12107);
or U12995 (N_12995,N_12468,N_12087);
nand U12996 (N_12996,N_12301,N_12264);
and U12997 (N_12997,N_12070,N_12445);
or U12998 (N_12998,N_12410,N_12190);
and U12999 (N_12999,N_12295,N_12188);
xor U13000 (N_13000,N_12829,N_12826);
or U13001 (N_13001,N_12947,N_12772);
or U13002 (N_13002,N_12588,N_12750);
xor U13003 (N_13003,N_12738,N_12878);
nor U13004 (N_13004,N_12566,N_12816);
nor U13005 (N_13005,N_12709,N_12877);
and U13006 (N_13006,N_12745,N_12714);
xnor U13007 (N_13007,N_12518,N_12621);
xor U13008 (N_13008,N_12847,N_12562);
and U13009 (N_13009,N_12648,N_12806);
or U13010 (N_13010,N_12994,N_12704);
and U13011 (N_13011,N_12602,N_12990);
nor U13012 (N_13012,N_12836,N_12611);
and U13013 (N_13013,N_12788,N_12778);
nand U13014 (N_13014,N_12871,N_12601);
nor U13015 (N_13015,N_12809,N_12755);
xor U13016 (N_13016,N_12657,N_12559);
or U13017 (N_13017,N_12623,N_12682);
nor U13018 (N_13018,N_12617,N_12692);
nor U13019 (N_13019,N_12673,N_12577);
nor U13020 (N_13020,N_12522,N_12606);
or U13021 (N_13021,N_12838,N_12919);
nand U13022 (N_13022,N_12550,N_12984);
xor U13023 (N_13023,N_12855,N_12681);
and U13024 (N_13024,N_12540,N_12767);
xor U13025 (N_13025,N_12624,N_12567);
nor U13026 (N_13026,N_12867,N_12728);
xor U13027 (N_13027,N_12554,N_12515);
nor U13028 (N_13028,N_12961,N_12907);
and U13029 (N_13029,N_12524,N_12687);
nor U13030 (N_13030,N_12944,N_12655);
xor U13031 (N_13031,N_12869,N_12979);
xnor U13032 (N_13032,N_12822,N_12744);
xnor U13033 (N_13033,N_12552,N_12993);
or U13034 (N_13034,N_12899,N_12946);
nor U13035 (N_13035,N_12995,N_12610);
nand U13036 (N_13036,N_12641,N_12991);
xor U13037 (N_13037,N_12781,N_12876);
or U13038 (N_13038,N_12960,N_12975);
nor U13039 (N_13039,N_12691,N_12951);
and U13040 (N_13040,N_12799,N_12743);
xnor U13041 (N_13041,N_12882,N_12690);
or U13042 (N_13042,N_12881,N_12708);
nand U13043 (N_13043,N_12604,N_12997);
nand U13044 (N_13044,N_12831,N_12773);
xnor U13045 (N_13045,N_12715,N_12915);
xnor U13046 (N_13046,N_12651,N_12584);
nor U13047 (N_13047,N_12563,N_12885);
and U13048 (N_13048,N_12790,N_12910);
nand U13049 (N_13049,N_12766,N_12627);
nor U13050 (N_13050,N_12520,N_12897);
nand U13051 (N_13051,N_12710,N_12747);
xnor U13052 (N_13052,N_12640,N_12635);
xor U13053 (N_13053,N_12940,N_12787);
xnor U13054 (N_13054,N_12535,N_12553);
or U13055 (N_13055,N_12542,N_12913);
nand U13056 (N_13056,N_12803,N_12865);
and U13057 (N_13057,N_12758,N_12805);
nor U13058 (N_13058,N_12544,N_12719);
xnor U13059 (N_13059,N_12683,N_12779);
nor U13060 (N_13060,N_12892,N_12536);
nor U13061 (N_13061,N_12506,N_12630);
xor U13062 (N_13062,N_12631,N_12762);
nand U13063 (N_13063,N_12634,N_12976);
nor U13064 (N_13064,N_12547,N_12771);
nand U13065 (N_13065,N_12924,N_12688);
xnor U13066 (N_13066,N_12653,N_12686);
nor U13067 (N_13067,N_12841,N_12693);
and U13068 (N_13068,N_12736,N_12797);
or U13069 (N_13069,N_12587,N_12902);
xor U13070 (N_13070,N_12864,N_12586);
nand U13071 (N_13071,N_12879,N_12849);
xnor U13072 (N_13072,N_12863,N_12917);
xnor U13073 (N_13073,N_12928,N_12903);
nand U13074 (N_13074,N_12672,N_12615);
and U13075 (N_13075,N_12723,N_12543);
or U13076 (N_13076,N_12721,N_12956);
nand U13077 (N_13077,N_12846,N_12854);
xor U13078 (N_13078,N_12858,N_12868);
or U13079 (N_13079,N_12717,N_12986);
nor U13080 (N_13080,N_12908,N_12894);
xnor U13081 (N_13081,N_12952,N_12861);
xor U13082 (N_13082,N_12784,N_12703);
or U13083 (N_13083,N_12911,N_12571);
nor U13084 (N_13084,N_12810,N_12546);
or U13085 (N_13085,N_12887,N_12938);
and U13086 (N_13086,N_12628,N_12666);
nor U13087 (N_13087,N_12914,N_12966);
or U13088 (N_13088,N_12740,N_12579);
xnor U13089 (N_13089,N_12950,N_12945);
xnor U13090 (N_13090,N_12503,N_12794);
nand U13091 (N_13091,N_12873,N_12848);
xnor U13092 (N_13092,N_12795,N_12982);
and U13093 (N_13093,N_12981,N_12501);
xnor U13094 (N_13094,N_12519,N_12551);
nor U13095 (N_13095,N_12517,N_12833);
nor U13096 (N_13096,N_12523,N_12815);
xor U13097 (N_13097,N_12886,N_12916);
or U13098 (N_13098,N_12942,N_12752);
xor U13099 (N_13099,N_12748,N_12510);
and U13100 (N_13100,N_12646,N_12680);
or U13101 (N_13101,N_12637,N_12801);
nor U13102 (N_13102,N_12605,N_12955);
nand U13103 (N_13103,N_12599,N_12880);
nand U13104 (N_13104,N_12670,N_12575);
nand U13105 (N_13105,N_12525,N_12711);
and U13106 (N_13106,N_12832,N_12972);
xnor U13107 (N_13107,N_12853,N_12576);
nand U13108 (N_13108,N_12500,N_12590);
nor U13109 (N_13109,N_12851,N_12812);
and U13110 (N_13110,N_12593,N_12514);
xnor U13111 (N_13111,N_12870,N_12732);
and U13112 (N_13112,N_12968,N_12607);
and U13113 (N_13113,N_12595,N_12565);
xnor U13114 (N_13114,N_12558,N_12701);
nor U13115 (N_13115,N_12927,N_12619);
and U13116 (N_13116,N_12932,N_12684);
nand U13117 (N_13117,N_12912,N_12931);
nand U13118 (N_13118,N_12729,N_12578);
nor U13119 (N_13119,N_12548,N_12645);
xnor U13120 (N_13120,N_12921,N_12639);
nand U13121 (N_13121,N_12937,N_12888);
or U13122 (N_13122,N_12786,N_12959);
nor U13123 (N_13123,N_12922,N_12753);
or U13124 (N_13124,N_12695,N_12782);
and U13125 (N_13125,N_12502,N_12652);
xnor U13126 (N_13126,N_12895,N_12793);
and U13127 (N_13127,N_12570,N_12574);
and U13128 (N_13128,N_12713,N_12970);
nand U13129 (N_13129,N_12900,N_12580);
nor U13130 (N_13130,N_12859,N_12532);
xnor U13131 (N_13131,N_12813,N_12739);
and U13132 (N_13132,N_12662,N_12700);
or U13133 (N_13133,N_12953,N_12834);
nand U13134 (N_13134,N_12776,N_12731);
nand U13135 (N_13135,N_12842,N_12596);
or U13136 (N_13136,N_12583,N_12933);
nand U13137 (N_13137,N_12702,N_12685);
nor U13138 (N_13138,N_12760,N_12513);
nor U13139 (N_13139,N_12789,N_12712);
and U13140 (N_13140,N_12845,N_12737);
nand U13141 (N_13141,N_12898,N_12971);
nor U13142 (N_13142,N_12835,N_12636);
or U13143 (N_13143,N_12527,N_12644);
or U13144 (N_13144,N_12706,N_12939);
or U13145 (N_13145,N_12891,N_12862);
xor U13146 (N_13146,N_12512,N_12957);
xor U13147 (N_13147,N_12850,N_12821);
and U13148 (N_13148,N_12622,N_12992);
nand U13149 (N_13149,N_12958,N_12973);
nor U13150 (N_13150,N_12844,N_12647);
and U13151 (N_13151,N_12720,N_12504);
or U13152 (N_13152,N_12671,N_12526);
or U13153 (N_13153,N_12726,N_12603);
nor U13154 (N_13154,N_12677,N_12597);
and U13155 (N_13155,N_12820,N_12564);
or U13156 (N_13156,N_12777,N_12727);
and U13157 (N_13157,N_12585,N_12965);
xnor U13158 (N_13158,N_12626,N_12507);
nor U13159 (N_13159,N_12722,N_12694);
and U13160 (N_13160,N_12591,N_12733);
or U13161 (N_13161,N_12904,N_12857);
xor U13162 (N_13162,N_12852,N_12757);
nor U13163 (N_13163,N_12807,N_12874);
xnor U13164 (N_13164,N_12998,N_12780);
and U13165 (N_13165,N_12906,N_12749);
xor U13166 (N_13166,N_12872,N_12901);
and U13167 (N_13167,N_12516,N_12632);
and U13168 (N_13168,N_12817,N_12661);
nand U13169 (N_13169,N_12676,N_12837);
nor U13170 (N_13170,N_12609,N_12734);
nor U13171 (N_13171,N_12770,N_12923);
or U13172 (N_13172,N_12556,N_12643);
and U13173 (N_13173,N_12980,N_12572);
nand U13174 (N_13174,N_12598,N_12533);
and U13175 (N_13175,N_12936,N_12557);
and U13176 (N_13176,N_12509,N_12808);
and U13177 (N_13177,N_12531,N_12746);
nand U13178 (N_13178,N_12920,N_12538);
or U13179 (N_13179,N_12941,N_12689);
nand U13180 (N_13180,N_12761,N_12905);
or U13181 (N_13181,N_12698,N_12716);
nor U13182 (N_13182,N_12742,N_12783);
xor U13183 (N_13183,N_12528,N_12560);
nand U13184 (N_13184,N_12629,N_12613);
or U13185 (N_13185,N_12718,N_12978);
nor U13186 (N_13186,N_12884,N_12568);
or U13187 (N_13187,N_12883,N_12592);
nand U13188 (N_13188,N_12823,N_12638);
xnor U13189 (N_13189,N_12875,N_12696);
and U13190 (N_13190,N_12893,N_12825);
nand U13191 (N_13191,N_12765,N_12511);
nand U13192 (N_13192,N_12963,N_12798);
nor U13193 (N_13193,N_12725,N_12660);
and U13194 (N_13194,N_12534,N_12561);
xor U13195 (N_13195,N_12785,N_12600);
and U13196 (N_13196,N_12530,N_12614);
nor U13197 (N_13197,N_12705,N_12549);
nand U13198 (N_13198,N_12792,N_12659);
nor U13199 (N_13199,N_12828,N_12811);
and U13200 (N_13200,N_12650,N_12667);
nand U13201 (N_13201,N_12843,N_12943);
nand U13202 (N_13202,N_12608,N_12663);
and U13203 (N_13203,N_12679,N_12707);
xor U13204 (N_13204,N_12999,N_12581);
or U13205 (N_13205,N_12537,N_12541);
xor U13206 (N_13206,N_12674,N_12800);
xor U13207 (N_13207,N_12804,N_12974);
or U13208 (N_13208,N_12830,N_12763);
or U13209 (N_13209,N_12529,N_12890);
or U13210 (N_13210,N_12935,N_12756);
nand U13211 (N_13211,N_12582,N_12678);
nand U13212 (N_13212,N_12969,N_12754);
or U13213 (N_13213,N_12896,N_12569);
and U13214 (N_13214,N_12618,N_12521);
nor U13215 (N_13215,N_12949,N_12989);
xor U13216 (N_13216,N_12764,N_12768);
or U13217 (N_13217,N_12866,N_12819);
nand U13218 (N_13218,N_12751,N_12818);
and U13219 (N_13219,N_12987,N_12625);
nand U13220 (N_13220,N_12697,N_12649);
xor U13221 (N_13221,N_12967,N_12730);
nor U13222 (N_13222,N_12508,N_12996);
nor U13223 (N_13223,N_12505,N_12934);
and U13224 (N_13224,N_12658,N_12669);
and U13225 (N_13225,N_12926,N_12918);
nor U13226 (N_13226,N_12664,N_12909);
nor U13227 (N_13227,N_12814,N_12769);
nor U13228 (N_13228,N_12964,N_12827);
and U13229 (N_13229,N_12735,N_12985);
nor U13230 (N_13230,N_12589,N_12620);
and U13231 (N_13231,N_12930,N_12759);
nand U13232 (N_13232,N_12983,N_12791);
nor U13233 (N_13233,N_12840,N_12962);
nand U13234 (N_13234,N_12545,N_12824);
and U13235 (N_13235,N_12612,N_12948);
nand U13236 (N_13236,N_12665,N_12539);
nand U13237 (N_13237,N_12668,N_12929);
and U13238 (N_13238,N_12796,N_12774);
or U13239 (N_13239,N_12954,N_12839);
and U13240 (N_13240,N_12860,N_12741);
xnor U13241 (N_13241,N_12724,N_12555);
nor U13242 (N_13242,N_12856,N_12616);
or U13243 (N_13243,N_12675,N_12775);
and U13244 (N_13244,N_12988,N_12977);
nor U13245 (N_13245,N_12802,N_12594);
nor U13246 (N_13246,N_12699,N_12642);
or U13247 (N_13247,N_12573,N_12656);
nor U13248 (N_13248,N_12889,N_12654);
or U13249 (N_13249,N_12925,N_12633);
and U13250 (N_13250,N_12898,N_12844);
xor U13251 (N_13251,N_12859,N_12821);
or U13252 (N_13252,N_12507,N_12638);
xnor U13253 (N_13253,N_12771,N_12609);
nand U13254 (N_13254,N_12560,N_12558);
nor U13255 (N_13255,N_12959,N_12668);
nand U13256 (N_13256,N_12965,N_12843);
nand U13257 (N_13257,N_12781,N_12866);
and U13258 (N_13258,N_12806,N_12734);
or U13259 (N_13259,N_12838,N_12512);
and U13260 (N_13260,N_12682,N_12770);
xor U13261 (N_13261,N_12666,N_12986);
nand U13262 (N_13262,N_12832,N_12656);
xor U13263 (N_13263,N_12959,N_12919);
nand U13264 (N_13264,N_12784,N_12943);
or U13265 (N_13265,N_12617,N_12859);
and U13266 (N_13266,N_12648,N_12687);
nand U13267 (N_13267,N_12707,N_12785);
and U13268 (N_13268,N_12944,N_12631);
or U13269 (N_13269,N_12684,N_12816);
or U13270 (N_13270,N_12693,N_12548);
or U13271 (N_13271,N_12556,N_12748);
xor U13272 (N_13272,N_12968,N_12580);
xnor U13273 (N_13273,N_12576,N_12694);
xor U13274 (N_13274,N_12548,N_12518);
and U13275 (N_13275,N_12746,N_12984);
and U13276 (N_13276,N_12576,N_12658);
nand U13277 (N_13277,N_12727,N_12813);
or U13278 (N_13278,N_12852,N_12756);
and U13279 (N_13279,N_12957,N_12862);
nor U13280 (N_13280,N_12637,N_12918);
nor U13281 (N_13281,N_12797,N_12881);
and U13282 (N_13282,N_12710,N_12716);
or U13283 (N_13283,N_12956,N_12876);
nor U13284 (N_13284,N_12894,N_12823);
xor U13285 (N_13285,N_12614,N_12508);
and U13286 (N_13286,N_12947,N_12518);
or U13287 (N_13287,N_12964,N_12689);
nand U13288 (N_13288,N_12655,N_12870);
nor U13289 (N_13289,N_12717,N_12706);
nand U13290 (N_13290,N_12922,N_12684);
and U13291 (N_13291,N_12867,N_12593);
nand U13292 (N_13292,N_12726,N_12652);
nor U13293 (N_13293,N_12655,N_12902);
or U13294 (N_13294,N_12733,N_12675);
and U13295 (N_13295,N_12854,N_12598);
nand U13296 (N_13296,N_12879,N_12745);
nand U13297 (N_13297,N_12907,N_12912);
and U13298 (N_13298,N_12534,N_12511);
nand U13299 (N_13299,N_12530,N_12797);
xnor U13300 (N_13300,N_12914,N_12811);
and U13301 (N_13301,N_12984,N_12798);
and U13302 (N_13302,N_12863,N_12827);
xnor U13303 (N_13303,N_12544,N_12725);
xnor U13304 (N_13304,N_12662,N_12817);
and U13305 (N_13305,N_12771,N_12892);
xor U13306 (N_13306,N_12665,N_12868);
or U13307 (N_13307,N_12785,N_12804);
and U13308 (N_13308,N_12956,N_12971);
nor U13309 (N_13309,N_12749,N_12579);
nand U13310 (N_13310,N_12519,N_12881);
xor U13311 (N_13311,N_12722,N_12716);
nand U13312 (N_13312,N_12927,N_12644);
nor U13313 (N_13313,N_12927,N_12570);
and U13314 (N_13314,N_12905,N_12972);
and U13315 (N_13315,N_12683,N_12845);
and U13316 (N_13316,N_12995,N_12999);
nor U13317 (N_13317,N_12651,N_12696);
or U13318 (N_13318,N_12764,N_12591);
and U13319 (N_13319,N_12830,N_12517);
or U13320 (N_13320,N_12666,N_12882);
nand U13321 (N_13321,N_12823,N_12729);
nand U13322 (N_13322,N_12782,N_12839);
nand U13323 (N_13323,N_12679,N_12650);
or U13324 (N_13324,N_12971,N_12770);
and U13325 (N_13325,N_12539,N_12797);
and U13326 (N_13326,N_12601,N_12521);
xor U13327 (N_13327,N_12767,N_12894);
nor U13328 (N_13328,N_12801,N_12511);
nand U13329 (N_13329,N_12752,N_12883);
xnor U13330 (N_13330,N_12932,N_12762);
xnor U13331 (N_13331,N_12705,N_12585);
nand U13332 (N_13332,N_12643,N_12516);
or U13333 (N_13333,N_12558,N_12539);
xnor U13334 (N_13334,N_12902,N_12535);
nand U13335 (N_13335,N_12589,N_12897);
or U13336 (N_13336,N_12755,N_12536);
xnor U13337 (N_13337,N_12632,N_12856);
or U13338 (N_13338,N_12765,N_12867);
nand U13339 (N_13339,N_12693,N_12978);
xor U13340 (N_13340,N_12827,N_12901);
xor U13341 (N_13341,N_12613,N_12793);
or U13342 (N_13342,N_12538,N_12979);
and U13343 (N_13343,N_12979,N_12779);
xnor U13344 (N_13344,N_12556,N_12651);
nand U13345 (N_13345,N_12822,N_12858);
nor U13346 (N_13346,N_12771,N_12821);
or U13347 (N_13347,N_12563,N_12775);
or U13348 (N_13348,N_12614,N_12945);
nor U13349 (N_13349,N_12611,N_12993);
and U13350 (N_13350,N_12669,N_12721);
nand U13351 (N_13351,N_12883,N_12873);
xnor U13352 (N_13352,N_12597,N_12962);
xnor U13353 (N_13353,N_12799,N_12961);
nor U13354 (N_13354,N_12760,N_12850);
and U13355 (N_13355,N_12889,N_12865);
and U13356 (N_13356,N_12525,N_12762);
or U13357 (N_13357,N_12552,N_12970);
and U13358 (N_13358,N_12848,N_12990);
and U13359 (N_13359,N_12505,N_12918);
xor U13360 (N_13360,N_12822,N_12798);
nor U13361 (N_13361,N_12968,N_12892);
nand U13362 (N_13362,N_12901,N_12641);
nand U13363 (N_13363,N_12716,N_12937);
and U13364 (N_13364,N_12655,N_12886);
and U13365 (N_13365,N_12875,N_12735);
or U13366 (N_13366,N_12752,N_12775);
or U13367 (N_13367,N_12847,N_12506);
nor U13368 (N_13368,N_12681,N_12527);
nor U13369 (N_13369,N_12870,N_12666);
xnor U13370 (N_13370,N_12664,N_12780);
or U13371 (N_13371,N_12582,N_12972);
nor U13372 (N_13372,N_12789,N_12823);
nor U13373 (N_13373,N_12972,N_12564);
and U13374 (N_13374,N_12803,N_12701);
nand U13375 (N_13375,N_12780,N_12602);
and U13376 (N_13376,N_12741,N_12981);
and U13377 (N_13377,N_12584,N_12965);
and U13378 (N_13378,N_12895,N_12569);
or U13379 (N_13379,N_12739,N_12602);
xor U13380 (N_13380,N_12814,N_12893);
xnor U13381 (N_13381,N_12986,N_12927);
nand U13382 (N_13382,N_12902,N_12869);
or U13383 (N_13383,N_12623,N_12616);
and U13384 (N_13384,N_12701,N_12654);
xor U13385 (N_13385,N_12837,N_12512);
xnor U13386 (N_13386,N_12528,N_12529);
xnor U13387 (N_13387,N_12855,N_12728);
or U13388 (N_13388,N_12602,N_12885);
or U13389 (N_13389,N_12642,N_12783);
nand U13390 (N_13390,N_12743,N_12949);
nor U13391 (N_13391,N_12836,N_12678);
or U13392 (N_13392,N_12585,N_12752);
and U13393 (N_13393,N_12943,N_12786);
nor U13394 (N_13394,N_12513,N_12998);
nand U13395 (N_13395,N_12621,N_12758);
and U13396 (N_13396,N_12840,N_12836);
or U13397 (N_13397,N_12585,N_12636);
or U13398 (N_13398,N_12694,N_12837);
xnor U13399 (N_13399,N_12775,N_12677);
and U13400 (N_13400,N_12657,N_12824);
nor U13401 (N_13401,N_12731,N_12511);
nand U13402 (N_13402,N_12659,N_12673);
and U13403 (N_13403,N_12619,N_12616);
nor U13404 (N_13404,N_12962,N_12624);
or U13405 (N_13405,N_12607,N_12894);
nor U13406 (N_13406,N_12585,N_12891);
or U13407 (N_13407,N_12507,N_12797);
and U13408 (N_13408,N_12720,N_12793);
nor U13409 (N_13409,N_12658,N_12789);
and U13410 (N_13410,N_12740,N_12595);
xnor U13411 (N_13411,N_12781,N_12962);
nand U13412 (N_13412,N_12733,N_12688);
xor U13413 (N_13413,N_12675,N_12735);
nand U13414 (N_13414,N_12804,N_12750);
nor U13415 (N_13415,N_12725,N_12614);
nand U13416 (N_13416,N_12585,N_12610);
nand U13417 (N_13417,N_12645,N_12555);
nand U13418 (N_13418,N_12865,N_12567);
xnor U13419 (N_13419,N_12819,N_12856);
xor U13420 (N_13420,N_12512,N_12971);
xor U13421 (N_13421,N_12859,N_12720);
and U13422 (N_13422,N_12776,N_12517);
xnor U13423 (N_13423,N_12553,N_12980);
and U13424 (N_13424,N_12758,N_12730);
nor U13425 (N_13425,N_12750,N_12853);
nor U13426 (N_13426,N_12588,N_12918);
nor U13427 (N_13427,N_12789,N_12854);
or U13428 (N_13428,N_12853,N_12545);
xor U13429 (N_13429,N_12712,N_12986);
and U13430 (N_13430,N_12651,N_12890);
or U13431 (N_13431,N_12994,N_12513);
or U13432 (N_13432,N_12659,N_12844);
xnor U13433 (N_13433,N_12893,N_12687);
and U13434 (N_13434,N_12960,N_12890);
or U13435 (N_13435,N_12692,N_12894);
and U13436 (N_13436,N_12853,N_12892);
nand U13437 (N_13437,N_12704,N_12714);
or U13438 (N_13438,N_12713,N_12564);
or U13439 (N_13439,N_12905,N_12553);
nand U13440 (N_13440,N_12536,N_12809);
nor U13441 (N_13441,N_12921,N_12595);
or U13442 (N_13442,N_12800,N_12938);
nor U13443 (N_13443,N_12590,N_12744);
or U13444 (N_13444,N_12577,N_12905);
xor U13445 (N_13445,N_12795,N_12671);
xor U13446 (N_13446,N_12508,N_12775);
xor U13447 (N_13447,N_12988,N_12576);
xor U13448 (N_13448,N_12993,N_12595);
and U13449 (N_13449,N_12572,N_12833);
nor U13450 (N_13450,N_12832,N_12927);
or U13451 (N_13451,N_12538,N_12862);
nand U13452 (N_13452,N_12938,N_12862);
xor U13453 (N_13453,N_12944,N_12667);
xor U13454 (N_13454,N_12807,N_12585);
and U13455 (N_13455,N_12701,N_12551);
or U13456 (N_13456,N_12881,N_12650);
and U13457 (N_13457,N_12906,N_12536);
nor U13458 (N_13458,N_12788,N_12883);
nor U13459 (N_13459,N_12581,N_12705);
or U13460 (N_13460,N_12661,N_12648);
and U13461 (N_13461,N_12929,N_12551);
and U13462 (N_13462,N_12862,N_12650);
and U13463 (N_13463,N_12891,N_12819);
or U13464 (N_13464,N_12635,N_12871);
nand U13465 (N_13465,N_12538,N_12524);
or U13466 (N_13466,N_12548,N_12827);
nor U13467 (N_13467,N_12582,N_12814);
xnor U13468 (N_13468,N_12946,N_12506);
and U13469 (N_13469,N_12561,N_12933);
or U13470 (N_13470,N_12595,N_12900);
and U13471 (N_13471,N_12630,N_12793);
and U13472 (N_13472,N_12598,N_12645);
or U13473 (N_13473,N_12523,N_12975);
nand U13474 (N_13474,N_12716,N_12666);
xor U13475 (N_13475,N_12915,N_12867);
nand U13476 (N_13476,N_12569,N_12932);
nand U13477 (N_13477,N_12914,N_12714);
and U13478 (N_13478,N_12615,N_12509);
xor U13479 (N_13479,N_12829,N_12531);
nand U13480 (N_13480,N_12691,N_12794);
nor U13481 (N_13481,N_12714,N_12715);
nand U13482 (N_13482,N_12693,N_12521);
xnor U13483 (N_13483,N_12785,N_12579);
and U13484 (N_13484,N_12975,N_12725);
xnor U13485 (N_13485,N_12514,N_12964);
nand U13486 (N_13486,N_12801,N_12986);
xor U13487 (N_13487,N_12699,N_12834);
and U13488 (N_13488,N_12712,N_12718);
xor U13489 (N_13489,N_12833,N_12646);
and U13490 (N_13490,N_12614,N_12738);
nor U13491 (N_13491,N_12785,N_12963);
and U13492 (N_13492,N_12746,N_12696);
nor U13493 (N_13493,N_12966,N_12963);
nor U13494 (N_13494,N_12838,N_12997);
xor U13495 (N_13495,N_12868,N_12594);
nor U13496 (N_13496,N_12986,N_12721);
or U13497 (N_13497,N_12701,N_12786);
nor U13498 (N_13498,N_12698,N_12501);
or U13499 (N_13499,N_12933,N_12666);
nand U13500 (N_13500,N_13219,N_13166);
xnor U13501 (N_13501,N_13373,N_13189);
and U13502 (N_13502,N_13042,N_13030);
nor U13503 (N_13503,N_13422,N_13286);
or U13504 (N_13504,N_13357,N_13162);
and U13505 (N_13505,N_13020,N_13003);
or U13506 (N_13506,N_13490,N_13266);
or U13507 (N_13507,N_13033,N_13330);
nand U13508 (N_13508,N_13382,N_13074);
nand U13509 (N_13509,N_13183,N_13334);
and U13510 (N_13510,N_13467,N_13368);
and U13511 (N_13511,N_13126,N_13326);
nor U13512 (N_13512,N_13083,N_13175);
nor U13513 (N_13513,N_13255,N_13433);
and U13514 (N_13514,N_13039,N_13023);
nand U13515 (N_13515,N_13131,N_13193);
xnor U13516 (N_13516,N_13116,N_13224);
nand U13517 (N_13517,N_13073,N_13497);
xor U13518 (N_13518,N_13237,N_13396);
or U13519 (N_13519,N_13135,N_13343);
or U13520 (N_13520,N_13350,N_13102);
xor U13521 (N_13521,N_13077,N_13208);
or U13522 (N_13522,N_13006,N_13066);
xnor U13523 (N_13523,N_13256,N_13246);
xor U13524 (N_13524,N_13276,N_13281);
or U13525 (N_13525,N_13241,N_13134);
nand U13526 (N_13526,N_13002,N_13488);
or U13527 (N_13527,N_13464,N_13097);
nand U13528 (N_13528,N_13137,N_13052);
and U13529 (N_13529,N_13474,N_13320);
xnor U13530 (N_13530,N_13265,N_13452);
nand U13531 (N_13531,N_13204,N_13218);
xnor U13532 (N_13532,N_13225,N_13104);
nand U13533 (N_13533,N_13412,N_13056);
nand U13534 (N_13534,N_13181,N_13348);
nor U13535 (N_13535,N_13191,N_13240);
and U13536 (N_13536,N_13391,N_13092);
nand U13537 (N_13537,N_13388,N_13115);
xor U13538 (N_13538,N_13302,N_13300);
or U13539 (N_13539,N_13378,N_13456);
nor U13540 (N_13540,N_13315,N_13366);
nand U13541 (N_13541,N_13428,N_13472);
and U13542 (N_13542,N_13211,N_13178);
or U13543 (N_13543,N_13340,N_13406);
and U13544 (N_13544,N_13027,N_13261);
nor U13545 (N_13545,N_13200,N_13125);
nor U13546 (N_13546,N_13132,N_13036);
or U13547 (N_13547,N_13417,N_13336);
nor U13548 (N_13548,N_13105,N_13057);
and U13549 (N_13549,N_13450,N_13195);
or U13550 (N_13550,N_13228,N_13419);
and U13551 (N_13551,N_13223,N_13100);
and U13552 (N_13552,N_13230,N_13446);
or U13553 (N_13553,N_13167,N_13038);
xor U13554 (N_13554,N_13093,N_13214);
and U13555 (N_13555,N_13453,N_13264);
nand U13556 (N_13556,N_13044,N_13114);
or U13557 (N_13557,N_13122,N_13227);
nor U13558 (N_13558,N_13411,N_13101);
nand U13559 (N_13559,N_13386,N_13408);
and U13560 (N_13560,N_13435,N_13476);
nand U13561 (N_13561,N_13064,N_13184);
and U13562 (N_13562,N_13109,N_13196);
nor U13563 (N_13563,N_13138,N_13233);
xnor U13564 (N_13564,N_13274,N_13098);
and U13565 (N_13565,N_13040,N_13113);
nor U13566 (N_13566,N_13017,N_13254);
xor U13567 (N_13567,N_13065,N_13094);
or U13568 (N_13568,N_13141,N_13048);
or U13569 (N_13569,N_13173,N_13339);
nand U13570 (N_13570,N_13427,N_13447);
or U13571 (N_13571,N_13229,N_13441);
nor U13572 (N_13572,N_13192,N_13130);
nand U13573 (N_13573,N_13164,N_13367);
nor U13574 (N_13574,N_13182,N_13213);
nor U13575 (N_13575,N_13426,N_13494);
or U13576 (N_13576,N_13272,N_13220);
xor U13577 (N_13577,N_13421,N_13055);
or U13578 (N_13578,N_13069,N_13331);
or U13579 (N_13579,N_13318,N_13215);
xor U13580 (N_13580,N_13163,N_13022);
and U13581 (N_13581,N_13153,N_13398);
or U13582 (N_13582,N_13086,N_13103);
or U13583 (N_13583,N_13176,N_13015);
or U13584 (N_13584,N_13142,N_13257);
and U13585 (N_13585,N_13159,N_13321);
nand U13586 (N_13586,N_13185,N_13448);
and U13587 (N_13587,N_13157,N_13053);
or U13588 (N_13588,N_13050,N_13404);
and U13589 (N_13589,N_13371,N_13080);
and U13590 (N_13590,N_13310,N_13444);
nor U13591 (N_13591,N_13025,N_13084);
nor U13592 (N_13592,N_13294,N_13370);
and U13593 (N_13593,N_13322,N_13091);
nand U13594 (N_13594,N_13385,N_13009);
or U13595 (N_13595,N_13059,N_13362);
nand U13596 (N_13596,N_13136,N_13271);
and U13597 (N_13597,N_13263,N_13262);
xnor U13598 (N_13598,N_13212,N_13041);
and U13599 (N_13599,N_13149,N_13127);
xor U13600 (N_13600,N_13324,N_13400);
nand U13601 (N_13601,N_13117,N_13155);
and U13602 (N_13602,N_13303,N_13121);
and U13603 (N_13603,N_13360,N_13244);
and U13604 (N_13604,N_13158,N_13110);
xor U13605 (N_13605,N_13221,N_13112);
and U13606 (N_13606,N_13222,N_13209);
or U13607 (N_13607,N_13111,N_13407);
or U13608 (N_13608,N_13005,N_13389);
nand U13609 (N_13609,N_13392,N_13235);
or U13610 (N_13610,N_13152,N_13304);
or U13611 (N_13611,N_13424,N_13416);
nor U13612 (N_13612,N_13377,N_13460);
xor U13613 (N_13613,N_13067,N_13409);
and U13614 (N_13614,N_13075,N_13353);
nand U13615 (N_13615,N_13096,N_13107);
nor U13616 (N_13616,N_13293,N_13455);
xor U13617 (N_13617,N_13365,N_13024);
nand U13618 (N_13618,N_13258,N_13451);
or U13619 (N_13619,N_13089,N_13190);
or U13620 (N_13620,N_13305,N_13418);
nor U13621 (N_13621,N_13147,N_13248);
xnor U13622 (N_13622,N_13429,N_13496);
and U13623 (N_13623,N_13280,N_13345);
xnor U13624 (N_13624,N_13432,N_13297);
xor U13625 (N_13625,N_13226,N_13313);
and U13626 (N_13626,N_13070,N_13465);
nand U13627 (N_13627,N_13168,N_13119);
or U13628 (N_13628,N_13380,N_13430);
and U13629 (N_13629,N_13442,N_13376);
nor U13630 (N_13630,N_13425,N_13410);
nand U13631 (N_13631,N_13043,N_13462);
nor U13632 (N_13632,N_13045,N_13128);
xor U13633 (N_13633,N_13449,N_13049);
nor U13634 (N_13634,N_13270,N_13437);
and U13635 (N_13635,N_13301,N_13277);
or U13636 (N_13636,N_13239,N_13351);
nor U13637 (N_13637,N_13471,N_13394);
nor U13638 (N_13638,N_13347,N_13046);
xnor U13639 (N_13639,N_13390,N_13150);
xor U13640 (N_13640,N_13354,N_13275);
nor U13641 (N_13641,N_13312,N_13217);
nor U13642 (N_13642,N_13018,N_13165);
nor U13643 (N_13643,N_13260,N_13259);
and U13644 (N_13644,N_13288,N_13188);
xnor U13645 (N_13645,N_13307,N_13061);
or U13646 (N_13646,N_13268,N_13478);
xor U13647 (N_13647,N_13319,N_13470);
or U13648 (N_13648,N_13387,N_13144);
and U13649 (N_13649,N_13361,N_13078);
and U13650 (N_13650,N_13201,N_13287);
or U13651 (N_13651,N_13363,N_13172);
or U13652 (N_13652,N_13123,N_13481);
nand U13653 (N_13653,N_13012,N_13072);
nor U13654 (N_13654,N_13440,N_13405);
or U13655 (N_13655,N_13458,N_13186);
nor U13656 (N_13656,N_13491,N_13037);
nand U13657 (N_13657,N_13384,N_13381);
xor U13658 (N_13658,N_13187,N_13352);
nand U13659 (N_13659,N_13311,N_13249);
or U13660 (N_13660,N_13206,N_13231);
nand U13661 (N_13661,N_13236,N_13194);
nor U13662 (N_13662,N_13431,N_13296);
nand U13663 (N_13663,N_13395,N_13068);
and U13664 (N_13664,N_13216,N_13011);
nand U13665 (N_13665,N_13001,N_13461);
and U13666 (N_13666,N_13129,N_13063);
and U13667 (N_13667,N_13285,N_13375);
or U13668 (N_13668,N_13156,N_13489);
xnor U13669 (N_13669,N_13328,N_13054);
and U13670 (N_13670,N_13468,N_13308);
nand U13671 (N_13671,N_13060,N_13358);
nor U13672 (N_13672,N_13014,N_13338);
nand U13673 (N_13673,N_13414,N_13314);
and U13674 (N_13674,N_13133,N_13087);
nand U13675 (N_13675,N_13309,N_13482);
nor U13676 (N_13676,N_13383,N_13180);
and U13677 (N_13677,N_13203,N_13306);
or U13678 (N_13678,N_13151,N_13483);
and U13679 (N_13679,N_13140,N_13359);
nand U13680 (N_13680,N_13459,N_13047);
nand U13681 (N_13681,N_13317,N_13160);
and U13682 (N_13682,N_13438,N_13238);
or U13683 (N_13683,N_13355,N_13245);
or U13684 (N_13684,N_13085,N_13493);
or U13685 (N_13685,N_13436,N_13013);
nor U13686 (N_13686,N_13028,N_13364);
nor U13687 (N_13687,N_13278,N_13034);
nand U13688 (N_13688,N_13327,N_13199);
and U13689 (N_13689,N_13492,N_13342);
xor U13690 (N_13690,N_13420,N_13253);
and U13691 (N_13691,N_13243,N_13332);
nand U13692 (N_13692,N_13487,N_13289);
or U13693 (N_13693,N_13171,N_13346);
nand U13694 (N_13694,N_13007,N_13403);
nor U13695 (N_13695,N_13008,N_13120);
and U13696 (N_13696,N_13273,N_13177);
or U13697 (N_13697,N_13369,N_13242);
nor U13698 (N_13698,N_13399,N_13466);
nor U13699 (N_13699,N_13250,N_13283);
nand U13700 (N_13700,N_13356,N_13210);
nor U13701 (N_13701,N_13207,N_13198);
nand U13702 (N_13702,N_13058,N_13004);
xnor U13703 (N_13703,N_13299,N_13082);
or U13704 (N_13704,N_13295,N_13484);
and U13705 (N_13705,N_13000,N_13393);
and U13706 (N_13706,N_13118,N_13349);
and U13707 (N_13707,N_13081,N_13251);
xnor U13708 (N_13708,N_13298,N_13415);
nand U13709 (N_13709,N_13090,N_13095);
or U13710 (N_13710,N_13071,N_13291);
nor U13711 (N_13711,N_13486,N_13413);
or U13712 (N_13712,N_13434,N_13205);
nor U13713 (N_13713,N_13010,N_13423);
and U13714 (N_13714,N_13202,N_13374);
and U13715 (N_13715,N_13076,N_13079);
xor U13716 (N_13716,N_13469,N_13401);
nand U13717 (N_13717,N_13341,N_13169);
and U13718 (N_13718,N_13143,N_13473);
xor U13719 (N_13719,N_13495,N_13179);
xnor U13720 (N_13720,N_13148,N_13443);
xnor U13721 (N_13721,N_13051,N_13232);
nand U13722 (N_13722,N_13267,N_13021);
xnor U13723 (N_13723,N_13284,N_13026);
xnor U13724 (N_13724,N_13019,N_13029);
xor U13725 (N_13725,N_13498,N_13139);
or U13726 (N_13726,N_13035,N_13479);
and U13727 (N_13727,N_13445,N_13279);
nand U13728 (N_13728,N_13154,N_13106);
and U13729 (N_13729,N_13234,N_13031);
xnor U13730 (N_13730,N_13323,N_13032);
and U13731 (N_13731,N_13475,N_13379);
xor U13732 (N_13732,N_13145,N_13170);
xnor U13733 (N_13733,N_13499,N_13335);
nor U13734 (N_13734,N_13316,N_13247);
or U13735 (N_13735,N_13457,N_13480);
nand U13736 (N_13736,N_13108,N_13088);
nand U13737 (N_13737,N_13329,N_13337);
xnor U13738 (N_13738,N_13402,N_13290);
and U13739 (N_13739,N_13062,N_13269);
nor U13740 (N_13740,N_13197,N_13485);
xor U13741 (N_13741,N_13282,N_13016);
nand U13742 (N_13742,N_13454,N_13333);
nand U13743 (N_13743,N_13344,N_13397);
xnor U13744 (N_13744,N_13099,N_13146);
xor U13745 (N_13745,N_13174,N_13325);
and U13746 (N_13746,N_13477,N_13161);
xnor U13747 (N_13747,N_13124,N_13252);
or U13748 (N_13748,N_13372,N_13292);
nand U13749 (N_13749,N_13439,N_13463);
nor U13750 (N_13750,N_13322,N_13306);
nor U13751 (N_13751,N_13030,N_13476);
nand U13752 (N_13752,N_13076,N_13301);
and U13753 (N_13753,N_13166,N_13161);
or U13754 (N_13754,N_13425,N_13400);
and U13755 (N_13755,N_13458,N_13448);
nand U13756 (N_13756,N_13249,N_13200);
and U13757 (N_13757,N_13477,N_13109);
nand U13758 (N_13758,N_13211,N_13427);
or U13759 (N_13759,N_13459,N_13347);
and U13760 (N_13760,N_13418,N_13255);
nor U13761 (N_13761,N_13359,N_13377);
nand U13762 (N_13762,N_13089,N_13119);
nor U13763 (N_13763,N_13208,N_13454);
and U13764 (N_13764,N_13197,N_13409);
or U13765 (N_13765,N_13095,N_13167);
xnor U13766 (N_13766,N_13433,N_13412);
or U13767 (N_13767,N_13220,N_13213);
nor U13768 (N_13768,N_13409,N_13460);
or U13769 (N_13769,N_13129,N_13001);
nor U13770 (N_13770,N_13390,N_13156);
xor U13771 (N_13771,N_13003,N_13225);
nor U13772 (N_13772,N_13491,N_13142);
nor U13773 (N_13773,N_13181,N_13356);
or U13774 (N_13774,N_13228,N_13144);
nand U13775 (N_13775,N_13383,N_13291);
xnor U13776 (N_13776,N_13129,N_13440);
xor U13777 (N_13777,N_13370,N_13236);
nand U13778 (N_13778,N_13428,N_13464);
nand U13779 (N_13779,N_13420,N_13173);
nand U13780 (N_13780,N_13078,N_13063);
nor U13781 (N_13781,N_13008,N_13012);
xor U13782 (N_13782,N_13374,N_13381);
and U13783 (N_13783,N_13042,N_13366);
nand U13784 (N_13784,N_13427,N_13218);
and U13785 (N_13785,N_13282,N_13345);
and U13786 (N_13786,N_13414,N_13189);
nand U13787 (N_13787,N_13221,N_13248);
nor U13788 (N_13788,N_13062,N_13027);
nand U13789 (N_13789,N_13300,N_13441);
xnor U13790 (N_13790,N_13331,N_13420);
and U13791 (N_13791,N_13158,N_13066);
or U13792 (N_13792,N_13167,N_13175);
nand U13793 (N_13793,N_13180,N_13133);
xnor U13794 (N_13794,N_13041,N_13215);
and U13795 (N_13795,N_13484,N_13319);
and U13796 (N_13796,N_13299,N_13262);
xor U13797 (N_13797,N_13349,N_13406);
and U13798 (N_13798,N_13320,N_13352);
and U13799 (N_13799,N_13103,N_13197);
and U13800 (N_13800,N_13340,N_13407);
or U13801 (N_13801,N_13190,N_13461);
nand U13802 (N_13802,N_13392,N_13078);
or U13803 (N_13803,N_13336,N_13234);
or U13804 (N_13804,N_13053,N_13003);
and U13805 (N_13805,N_13481,N_13009);
nand U13806 (N_13806,N_13108,N_13019);
nand U13807 (N_13807,N_13176,N_13017);
nand U13808 (N_13808,N_13047,N_13003);
or U13809 (N_13809,N_13161,N_13283);
and U13810 (N_13810,N_13057,N_13301);
xor U13811 (N_13811,N_13081,N_13357);
and U13812 (N_13812,N_13488,N_13122);
xor U13813 (N_13813,N_13047,N_13487);
and U13814 (N_13814,N_13170,N_13259);
nor U13815 (N_13815,N_13307,N_13350);
xnor U13816 (N_13816,N_13384,N_13007);
nor U13817 (N_13817,N_13045,N_13174);
xor U13818 (N_13818,N_13371,N_13195);
or U13819 (N_13819,N_13013,N_13360);
or U13820 (N_13820,N_13232,N_13034);
nor U13821 (N_13821,N_13383,N_13143);
or U13822 (N_13822,N_13142,N_13365);
nand U13823 (N_13823,N_13060,N_13091);
and U13824 (N_13824,N_13366,N_13494);
xnor U13825 (N_13825,N_13403,N_13092);
and U13826 (N_13826,N_13473,N_13262);
and U13827 (N_13827,N_13133,N_13232);
and U13828 (N_13828,N_13078,N_13257);
nand U13829 (N_13829,N_13005,N_13496);
xor U13830 (N_13830,N_13091,N_13407);
and U13831 (N_13831,N_13251,N_13381);
nor U13832 (N_13832,N_13153,N_13043);
xnor U13833 (N_13833,N_13242,N_13285);
nor U13834 (N_13834,N_13071,N_13128);
and U13835 (N_13835,N_13434,N_13068);
nand U13836 (N_13836,N_13188,N_13325);
xor U13837 (N_13837,N_13333,N_13018);
or U13838 (N_13838,N_13351,N_13290);
and U13839 (N_13839,N_13032,N_13482);
and U13840 (N_13840,N_13424,N_13188);
or U13841 (N_13841,N_13340,N_13353);
or U13842 (N_13842,N_13368,N_13095);
or U13843 (N_13843,N_13409,N_13209);
and U13844 (N_13844,N_13037,N_13395);
or U13845 (N_13845,N_13452,N_13350);
and U13846 (N_13846,N_13261,N_13472);
nor U13847 (N_13847,N_13365,N_13475);
nand U13848 (N_13848,N_13233,N_13107);
nor U13849 (N_13849,N_13042,N_13202);
or U13850 (N_13850,N_13133,N_13435);
nor U13851 (N_13851,N_13170,N_13338);
nor U13852 (N_13852,N_13103,N_13457);
nor U13853 (N_13853,N_13144,N_13484);
and U13854 (N_13854,N_13214,N_13484);
nor U13855 (N_13855,N_13346,N_13247);
and U13856 (N_13856,N_13358,N_13261);
or U13857 (N_13857,N_13403,N_13457);
or U13858 (N_13858,N_13100,N_13095);
nor U13859 (N_13859,N_13330,N_13026);
and U13860 (N_13860,N_13123,N_13132);
nor U13861 (N_13861,N_13300,N_13361);
or U13862 (N_13862,N_13331,N_13493);
nor U13863 (N_13863,N_13052,N_13014);
nor U13864 (N_13864,N_13297,N_13477);
xnor U13865 (N_13865,N_13370,N_13302);
or U13866 (N_13866,N_13463,N_13202);
or U13867 (N_13867,N_13459,N_13345);
and U13868 (N_13868,N_13196,N_13464);
nor U13869 (N_13869,N_13047,N_13470);
xnor U13870 (N_13870,N_13278,N_13297);
nor U13871 (N_13871,N_13184,N_13237);
xnor U13872 (N_13872,N_13419,N_13415);
and U13873 (N_13873,N_13225,N_13455);
nor U13874 (N_13874,N_13425,N_13023);
nor U13875 (N_13875,N_13433,N_13312);
xor U13876 (N_13876,N_13415,N_13489);
and U13877 (N_13877,N_13332,N_13167);
nand U13878 (N_13878,N_13144,N_13351);
or U13879 (N_13879,N_13370,N_13305);
xor U13880 (N_13880,N_13451,N_13458);
xnor U13881 (N_13881,N_13495,N_13397);
or U13882 (N_13882,N_13020,N_13469);
xor U13883 (N_13883,N_13123,N_13122);
and U13884 (N_13884,N_13385,N_13100);
nor U13885 (N_13885,N_13275,N_13407);
nand U13886 (N_13886,N_13361,N_13416);
or U13887 (N_13887,N_13288,N_13180);
nand U13888 (N_13888,N_13058,N_13017);
nand U13889 (N_13889,N_13199,N_13296);
nand U13890 (N_13890,N_13344,N_13104);
nor U13891 (N_13891,N_13184,N_13378);
and U13892 (N_13892,N_13162,N_13353);
xor U13893 (N_13893,N_13242,N_13458);
nand U13894 (N_13894,N_13411,N_13456);
nand U13895 (N_13895,N_13065,N_13237);
or U13896 (N_13896,N_13114,N_13196);
or U13897 (N_13897,N_13234,N_13427);
nor U13898 (N_13898,N_13074,N_13199);
nand U13899 (N_13899,N_13194,N_13412);
and U13900 (N_13900,N_13052,N_13027);
nand U13901 (N_13901,N_13245,N_13098);
and U13902 (N_13902,N_13485,N_13136);
nand U13903 (N_13903,N_13164,N_13047);
or U13904 (N_13904,N_13454,N_13083);
nand U13905 (N_13905,N_13190,N_13111);
xor U13906 (N_13906,N_13052,N_13012);
nor U13907 (N_13907,N_13379,N_13044);
nor U13908 (N_13908,N_13471,N_13094);
xnor U13909 (N_13909,N_13302,N_13359);
and U13910 (N_13910,N_13272,N_13362);
or U13911 (N_13911,N_13458,N_13153);
and U13912 (N_13912,N_13338,N_13451);
nand U13913 (N_13913,N_13296,N_13190);
nand U13914 (N_13914,N_13264,N_13010);
or U13915 (N_13915,N_13102,N_13479);
nand U13916 (N_13916,N_13225,N_13061);
or U13917 (N_13917,N_13460,N_13042);
nand U13918 (N_13918,N_13298,N_13048);
xnor U13919 (N_13919,N_13428,N_13037);
xor U13920 (N_13920,N_13380,N_13189);
and U13921 (N_13921,N_13433,N_13108);
nor U13922 (N_13922,N_13495,N_13463);
nand U13923 (N_13923,N_13062,N_13377);
or U13924 (N_13924,N_13198,N_13414);
and U13925 (N_13925,N_13155,N_13035);
nor U13926 (N_13926,N_13478,N_13078);
xnor U13927 (N_13927,N_13038,N_13156);
and U13928 (N_13928,N_13242,N_13035);
xor U13929 (N_13929,N_13438,N_13155);
and U13930 (N_13930,N_13419,N_13420);
or U13931 (N_13931,N_13132,N_13236);
xor U13932 (N_13932,N_13480,N_13193);
or U13933 (N_13933,N_13015,N_13459);
nor U13934 (N_13934,N_13392,N_13284);
or U13935 (N_13935,N_13271,N_13064);
nand U13936 (N_13936,N_13209,N_13382);
or U13937 (N_13937,N_13140,N_13005);
nor U13938 (N_13938,N_13229,N_13462);
or U13939 (N_13939,N_13315,N_13259);
xnor U13940 (N_13940,N_13163,N_13305);
nand U13941 (N_13941,N_13111,N_13212);
xor U13942 (N_13942,N_13429,N_13436);
xnor U13943 (N_13943,N_13173,N_13390);
xnor U13944 (N_13944,N_13286,N_13027);
xor U13945 (N_13945,N_13071,N_13257);
nor U13946 (N_13946,N_13177,N_13263);
or U13947 (N_13947,N_13078,N_13233);
nor U13948 (N_13948,N_13072,N_13161);
xor U13949 (N_13949,N_13309,N_13160);
nor U13950 (N_13950,N_13237,N_13098);
nor U13951 (N_13951,N_13030,N_13024);
and U13952 (N_13952,N_13019,N_13424);
and U13953 (N_13953,N_13153,N_13367);
nor U13954 (N_13954,N_13135,N_13222);
or U13955 (N_13955,N_13211,N_13194);
nand U13956 (N_13956,N_13426,N_13056);
and U13957 (N_13957,N_13468,N_13292);
and U13958 (N_13958,N_13209,N_13309);
nand U13959 (N_13959,N_13360,N_13385);
or U13960 (N_13960,N_13186,N_13415);
nor U13961 (N_13961,N_13003,N_13358);
and U13962 (N_13962,N_13354,N_13029);
and U13963 (N_13963,N_13003,N_13092);
and U13964 (N_13964,N_13400,N_13416);
nand U13965 (N_13965,N_13016,N_13198);
or U13966 (N_13966,N_13253,N_13314);
and U13967 (N_13967,N_13417,N_13378);
nor U13968 (N_13968,N_13063,N_13138);
nand U13969 (N_13969,N_13260,N_13480);
xnor U13970 (N_13970,N_13072,N_13376);
or U13971 (N_13971,N_13467,N_13444);
and U13972 (N_13972,N_13492,N_13346);
xor U13973 (N_13973,N_13225,N_13489);
and U13974 (N_13974,N_13499,N_13312);
xnor U13975 (N_13975,N_13047,N_13417);
nand U13976 (N_13976,N_13097,N_13433);
nor U13977 (N_13977,N_13247,N_13238);
or U13978 (N_13978,N_13196,N_13297);
nand U13979 (N_13979,N_13198,N_13144);
nor U13980 (N_13980,N_13403,N_13417);
or U13981 (N_13981,N_13101,N_13463);
nand U13982 (N_13982,N_13372,N_13137);
xor U13983 (N_13983,N_13326,N_13431);
nor U13984 (N_13984,N_13360,N_13322);
xnor U13985 (N_13985,N_13440,N_13121);
xnor U13986 (N_13986,N_13378,N_13327);
nor U13987 (N_13987,N_13167,N_13311);
or U13988 (N_13988,N_13219,N_13472);
or U13989 (N_13989,N_13167,N_13136);
xor U13990 (N_13990,N_13460,N_13407);
or U13991 (N_13991,N_13088,N_13410);
nand U13992 (N_13992,N_13350,N_13315);
or U13993 (N_13993,N_13220,N_13083);
xor U13994 (N_13994,N_13148,N_13122);
and U13995 (N_13995,N_13122,N_13287);
nand U13996 (N_13996,N_13335,N_13061);
xnor U13997 (N_13997,N_13025,N_13014);
or U13998 (N_13998,N_13248,N_13195);
or U13999 (N_13999,N_13466,N_13347);
nand U14000 (N_14000,N_13704,N_13559);
xor U14001 (N_14001,N_13977,N_13918);
nand U14002 (N_14002,N_13631,N_13660);
or U14003 (N_14003,N_13819,N_13715);
xor U14004 (N_14004,N_13993,N_13900);
or U14005 (N_14005,N_13769,N_13808);
nor U14006 (N_14006,N_13873,N_13696);
nor U14007 (N_14007,N_13664,N_13632);
xor U14008 (N_14008,N_13840,N_13941);
and U14009 (N_14009,N_13733,N_13770);
nor U14010 (N_14010,N_13590,N_13627);
nor U14011 (N_14011,N_13948,N_13556);
nand U14012 (N_14012,N_13915,N_13966);
nor U14013 (N_14013,N_13581,N_13899);
xor U14014 (N_14014,N_13884,N_13897);
nor U14015 (N_14015,N_13806,N_13766);
and U14016 (N_14016,N_13836,N_13751);
or U14017 (N_14017,N_13686,N_13894);
xnor U14018 (N_14018,N_13618,N_13600);
xor U14019 (N_14019,N_13591,N_13845);
xnor U14020 (N_14020,N_13516,N_13655);
and U14021 (N_14021,N_13519,N_13865);
or U14022 (N_14022,N_13677,N_13799);
and U14023 (N_14023,N_13526,N_13726);
nor U14024 (N_14024,N_13725,N_13574);
nand U14025 (N_14025,N_13714,N_13602);
or U14026 (N_14026,N_13752,N_13853);
nand U14027 (N_14027,N_13589,N_13886);
and U14028 (N_14028,N_13812,N_13976);
or U14029 (N_14029,N_13986,N_13832);
xor U14030 (N_14030,N_13956,N_13807);
or U14031 (N_14031,N_13640,N_13851);
nand U14032 (N_14032,N_13539,N_13579);
and U14033 (N_14033,N_13774,N_13713);
or U14034 (N_14034,N_13711,N_13735);
and U14035 (N_14035,N_13973,N_13916);
or U14036 (N_14036,N_13998,N_13626);
and U14037 (N_14037,N_13734,N_13944);
nor U14038 (N_14038,N_13820,N_13954);
nor U14039 (N_14039,N_13995,N_13773);
nor U14040 (N_14040,N_13505,N_13762);
nand U14041 (N_14041,N_13515,N_13763);
nor U14042 (N_14042,N_13864,N_13643);
nor U14043 (N_14043,N_13779,N_13546);
nor U14044 (N_14044,N_13800,N_13983);
or U14045 (N_14045,N_13937,N_13697);
and U14046 (N_14046,N_13789,N_13580);
and U14047 (N_14047,N_13549,N_13963);
nor U14048 (N_14048,N_13657,N_13501);
or U14049 (N_14049,N_13532,N_13710);
xnor U14050 (N_14050,N_13508,N_13658);
and U14051 (N_14051,N_13747,N_13652);
and U14052 (N_14052,N_13835,N_13616);
and U14053 (N_14053,N_13606,N_13518);
nand U14054 (N_14054,N_13538,N_13682);
nand U14055 (N_14055,N_13957,N_13745);
nand U14056 (N_14056,N_13996,N_13938);
nand U14057 (N_14057,N_13932,N_13582);
xor U14058 (N_14058,N_13622,N_13802);
and U14059 (N_14059,N_13716,N_13634);
nand U14060 (N_14060,N_13911,N_13533);
nand U14061 (N_14061,N_13862,N_13987);
xnor U14062 (N_14062,N_13568,N_13969);
xor U14063 (N_14063,N_13588,N_13831);
nand U14064 (N_14064,N_13841,N_13542);
and U14065 (N_14065,N_13702,N_13760);
nor U14066 (N_14066,N_13794,N_13690);
nand U14067 (N_14067,N_13666,N_13685);
or U14068 (N_14068,N_13687,N_13936);
nor U14069 (N_14069,N_13972,N_13815);
nand U14070 (N_14070,N_13651,N_13708);
nor U14071 (N_14071,N_13898,N_13950);
xnor U14072 (N_14072,N_13576,N_13573);
xor U14073 (N_14073,N_13824,N_13695);
or U14074 (N_14074,N_13537,N_13509);
nand U14075 (N_14075,N_13730,N_13585);
xnor U14076 (N_14076,N_13625,N_13759);
nor U14077 (N_14077,N_13684,N_13777);
and U14078 (N_14078,N_13907,N_13741);
and U14079 (N_14079,N_13903,N_13738);
and U14080 (N_14080,N_13617,N_13952);
nor U14081 (N_14081,N_13727,N_13951);
xor U14082 (N_14082,N_13883,N_13653);
xor U14083 (N_14083,N_13614,N_13829);
nand U14084 (N_14084,N_13927,N_13563);
or U14085 (N_14085,N_13707,N_13608);
xnor U14086 (N_14086,N_13848,N_13888);
and U14087 (N_14087,N_13648,N_13929);
and U14088 (N_14088,N_13558,N_13992);
nand U14089 (N_14089,N_13828,N_13749);
xor U14090 (N_14090,N_13717,N_13876);
and U14091 (N_14091,N_13858,N_13721);
or U14092 (N_14092,N_13594,N_13557);
or U14093 (N_14093,N_13723,N_13673);
nand U14094 (N_14094,N_13678,N_13659);
or U14095 (N_14095,N_13867,N_13786);
xnor U14096 (N_14096,N_13940,N_13822);
and U14097 (N_14097,N_13919,N_13795);
nor U14098 (N_14098,N_13587,N_13781);
xor U14099 (N_14099,N_13688,N_13758);
or U14100 (N_14100,N_13810,N_13880);
or U14101 (N_14101,N_13592,N_13562);
xor U14102 (N_14102,N_13661,N_13842);
nand U14103 (N_14103,N_13910,N_13837);
or U14104 (N_14104,N_13586,N_13968);
or U14105 (N_14105,N_13906,N_13826);
nor U14106 (N_14106,N_13544,N_13772);
nor U14107 (N_14107,N_13550,N_13679);
nor U14108 (N_14108,N_13896,N_13722);
nor U14109 (N_14109,N_13566,N_13583);
and U14110 (N_14110,N_13649,N_13870);
or U14111 (N_14111,N_13805,N_13584);
nand U14112 (N_14112,N_13512,N_13724);
xnor U14113 (N_14113,N_13732,N_13619);
xor U14114 (N_14114,N_13925,N_13784);
nand U14115 (N_14115,N_13520,N_13612);
nand U14116 (N_14116,N_13613,N_13570);
or U14117 (N_14117,N_13611,N_13645);
nand U14118 (N_14118,N_13671,N_13691);
nor U14119 (N_14119,N_13676,N_13924);
xor U14120 (N_14120,N_13525,N_13750);
nor U14121 (N_14121,N_13528,N_13877);
nor U14122 (N_14122,N_13793,N_13530);
xor U14123 (N_14123,N_13739,N_13680);
or U14124 (N_14124,N_13979,N_13788);
xor U14125 (N_14125,N_13737,N_13521);
nor U14126 (N_14126,N_13565,N_13912);
xor U14127 (N_14127,N_13889,N_13719);
or U14128 (N_14128,N_13668,N_13629);
or U14129 (N_14129,N_13596,N_13939);
or U14130 (N_14130,N_13798,N_13561);
nor U14131 (N_14131,N_13922,N_13635);
nor U14132 (N_14132,N_13895,N_13905);
nor U14133 (N_14133,N_13796,N_13644);
nand U14134 (N_14134,N_13693,N_13578);
nor U14135 (N_14135,N_13683,N_13637);
nand U14136 (N_14136,N_13534,N_13605);
nand U14137 (N_14137,N_13554,N_13999);
nand U14138 (N_14138,N_13630,N_13597);
xnor U14139 (N_14139,N_13931,N_13981);
nor U14140 (N_14140,N_13620,N_13847);
and U14141 (N_14141,N_13875,N_13731);
and U14142 (N_14142,N_13874,N_13933);
xnor U14143 (N_14143,N_13599,N_13672);
nor U14144 (N_14144,N_13609,N_13857);
xnor U14145 (N_14145,N_13775,N_13964);
and U14146 (N_14146,N_13830,N_13809);
and U14147 (N_14147,N_13949,N_13804);
nand U14148 (N_14148,N_13572,N_13982);
nand U14149 (N_14149,N_13641,N_13926);
nand U14150 (N_14150,N_13610,N_13548);
nor U14151 (N_14151,N_13890,N_13506);
nand U14152 (N_14152,N_13507,N_13856);
nor U14153 (N_14153,N_13628,N_13958);
xor U14154 (N_14154,N_13965,N_13720);
xnor U14155 (N_14155,N_13694,N_13813);
and U14156 (N_14156,N_13863,N_13959);
nand U14157 (N_14157,N_13689,N_13852);
nor U14158 (N_14158,N_13975,N_13878);
nor U14159 (N_14159,N_13881,N_13571);
nor U14160 (N_14160,N_13901,N_13791);
nor U14161 (N_14161,N_13553,N_13844);
nand U14162 (N_14162,N_13706,N_13754);
nor U14163 (N_14163,N_13990,N_13569);
or U14164 (N_14164,N_13768,N_13792);
xnor U14165 (N_14165,N_13882,N_13513);
nor U14166 (N_14166,N_13555,N_13838);
or U14167 (N_14167,N_13849,N_13543);
or U14168 (N_14168,N_13633,N_13756);
and U14169 (N_14169,N_13712,N_13598);
xor U14170 (N_14170,N_13892,N_13729);
nand U14171 (N_14171,N_13928,N_13943);
and U14172 (N_14172,N_13833,N_13980);
or U14173 (N_14173,N_13700,N_13891);
and U14174 (N_14174,N_13991,N_13934);
nor U14175 (N_14175,N_13913,N_13771);
xnor U14176 (N_14176,N_13701,N_13776);
or U14177 (N_14177,N_13642,N_13654);
and U14178 (N_14178,N_13960,N_13669);
nand U14179 (N_14179,N_13511,N_13879);
xor U14180 (N_14180,N_13709,N_13524);
or U14181 (N_14181,N_13967,N_13988);
xnor U14182 (N_14182,N_13665,N_13545);
nand U14183 (N_14183,N_13593,N_13855);
or U14184 (N_14184,N_13974,N_13904);
and U14185 (N_14185,N_13984,N_13601);
nand U14186 (N_14186,N_13947,N_13767);
nand U14187 (N_14187,N_13985,N_13790);
nor U14188 (N_14188,N_13502,N_13914);
or U14189 (N_14189,N_13503,N_13811);
xor U14190 (N_14190,N_13782,N_13510);
and U14191 (N_14191,N_13978,N_13761);
nor U14192 (N_14192,N_13698,N_13930);
nand U14193 (N_14193,N_13785,N_13667);
xnor U14194 (N_14194,N_13971,N_13755);
and U14195 (N_14195,N_13803,N_13753);
nor U14196 (N_14196,N_13869,N_13604);
nand U14197 (N_14197,N_13740,N_13923);
nor U14198 (N_14198,N_13868,N_13529);
nand U14199 (N_14199,N_13663,N_13577);
and U14200 (N_14200,N_13681,N_13765);
or U14201 (N_14201,N_13675,N_13962);
xor U14202 (N_14202,N_13670,N_13764);
or U14203 (N_14203,N_13860,N_13531);
nor U14204 (N_14204,N_13736,N_13551);
nor U14205 (N_14205,N_13744,N_13623);
nor U14206 (N_14206,N_13872,N_13825);
nor U14207 (N_14207,N_13994,N_13517);
and U14208 (N_14208,N_13834,N_13921);
and U14209 (N_14209,N_13780,N_13636);
and U14210 (N_14210,N_13607,N_13850);
nand U14211 (N_14211,N_13817,N_13742);
xnor U14212 (N_14212,N_13946,N_13603);
xor U14213 (N_14213,N_13567,N_13692);
nand U14214 (N_14214,N_13816,N_13522);
xnor U14215 (N_14215,N_13823,N_13646);
nand U14216 (N_14216,N_13902,N_13787);
nand U14217 (N_14217,N_13500,N_13656);
and U14218 (N_14218,N_13997,N_13818);
xnor U14219 (N_14219,N_13699,N_13674);
nor U14220 (N_14220,N_13564,N_13514);
nand U14221 (N_14221,N_13854,N_13718);
or U14222 (N_14222,N_13647,N_13871);
xor U14223 (N_14223,N_13859,N_13942);
nand U14224 (N_14224,N_13955,N_13703);
nand U14225 (N_14225,N_13535,N_13527);
nand U14226 (N_14226,N_13953,N_13861);
xor U14227 (N_14227,N_13827,N_13814);
or U14228 (N_14228,N_13908,N_13743);
and U14229 (N_14229,N_13547,N_13945);
nor U14230 (N_14230,N_13970,N_13650);
xor U14231 (N_14231,N_13887,N_13801);
or U14232 (N_14232,N_13504,N_13839);
nor U14233 (N_14233,N_13638,N_13893);
nor U14234 (N_14234,N_13961,N_13536);
nand U14235 (N_14235,N_13866,N_13920);
xnor U14236 (N_14236,N_13662,N_13705);
or U14237 (N_14237,N_13523,N_13885);
or U14238 (N_14238,N_13621,N_13778);
xor U14239 (N_14239,N_13540,N_13728);
nand U14240 (N_14240,N_13843,N_13846);
nand U14241 (N_14241,N_13797,N_13909);
xnor U14242 (N_14242,N_13541,N_13748);
and U14243 (N_14243,N_13917,N_13783);
and U14244 (N_14244,N_13560,N_13746);
nor U14245 (N_14245,N_13935,N_13624);
nand U14246 (N_14246,N_13989,N_13595);
and U14247 (N_14247,N_13552,N_13757);
xnor U14248 (N_14248,N_13639,N_13575);
and U14249 (N_14249,N_13821,N_13615);
nand U14250 (N_14250,N_13976,N_13856);
nand U14251 (N_14251,N_13668,N_13584);
or U14252 (N_14252,N_13821,N_13726);
nor U14253 (N_14253,N_13502,N_13583);
xnor U14254 (N_14254,N_13672,N_13971);
and U14255 (N_14255,N_13601,N_13559);
or U14256 (N_14256,N_13712,N_13996);
or U14257 (N_14257,N_13708,N_13919);
nand U14258 (N_14258,N_13911,N_13539);
nor U14259 (N_14259,N_13754,N_13524);
and U14260 (N_14260,N_13616,N_13697);
nor U14261 (N_14261,N_13722,N_13738);
nor U14262 (N_14262,N_13716,N_13896);
and U14263 (N_14263,N_13952,N_13858);
nand U14264 (N_14264,N_13782,N_13784);
nand U14265 (N_14265,N_13766,N_13665);
nand U14266 (N_14266,N_13699,N_13732);
xor U14267 (N_14267,N_13746,N_13626);
or U14268 (N_14268,N_13985,N_13836);
nor U14269 (N_14269,N_13894,N_13945);
nor U14270 (N_14270,N_13828,N_13928);
nor U14271 (N_14271,N_13797,N_13565);
nor U14272 (N_14272,N_13525,N_13900);
nand U14273 (N_14273,N_13649,N_13798);
and U14274 (N_14274,N_13799,N_13521);
nor U14275 (N_14275,N_13539,N_13626);
or U14276 (N_14276,N_13956,N_13827);
nor U14277 (N_14277,N_13986,N_13788);
nand U14278 (N_14278,N_13702,N_13608);
and U14279 (N_14279,N_13803,N_13549);
and U14280 (N_14280,N_13999,N_13700);
or U14281 (N_14281,N_13969,N_13523);
nand U14282 (N_14282,N_13567,N_13941);
and U14283 (N_14283,N_13696,N_13704);
nor U14284 (N_14284,N_13638,N_13944);
xor U14285 (N_14285,N_13899,N_13785);
nand U14286 (N_14286,N_13758,N_13722);
xnor U14287 (N_14287,N_13859,N_13521);
nor U14288 (N_14288,N_13672,N_13683);
nand U14289 (N_14289,N_13733,N_13695);
or U14290 (N_14290,N_13602,N_13514);
or U14291 (N_14291,N_13585,N_13522);
and U14292 (N_14292,N_13839,N_13645);
xor U14293 (N_14293,N_13553,N_13854);
or U14294 (N_14294,N_13847,N_13563);
or U14295 (N_14295,N_13949,N_13979);
or U14296 (N_14296,N_13922,N_13539);
and U14297 (N_14297,N_13659,N_13972);
nor U14298 (N_14298,N_13633,N_13503);
xor U14299 (N_14299,N_13882,N_13665);
nand U14300 (N_14300,N_13758,N_13753);
or U14301 (N_14301,N_13671,N_13580);
and U14302 (N_14302,N_13677,N_13862);
or U14303 (N_14303,N_13701,N_13666);
and U14304 (N_14304,N_13761,N_13658);
nor U14305 (N_14305,N_13670,N_13736);
xnor U14306 (N_14306,N_13637,N_13702);
and U14307 (N_14307,N_13716,N_13590);
or U14308 (N_14308,N_13736,N_13565);
and U14309 (N_14309,N_13939,N_13597);
xnor U14310 (N_14310,N_13727,N_13765);
and U14311 (N_14311,N_13806,N_13899);
xnor U14312 (N_14312,N_13780,N_13986);
nor U14313 (N_14313,N_13727,N_13614);
nand U14314 (N_14314,N_13588,N_13867);
or U14315 (N_14315,N_13525,N_13584);
nor U14316 (N_14316,N_13618,N_13523);
or U14317 (N_14317,N_13680,N_13963);
and U14318 (N_14318,N_13976,N_13868);
or U14319 (N_14319,N_13755,N_13851);
and U14320 (N_14320,N_13664,N_13714);
and U14321 (N_14321,N_13560,N_13738);
xor U14322 (N_14322,N_13617,N_13767);
xor U14323 (N_14323,N_13590,N_13598);
nor U14324 (N_14324,N_13601,N_13968);
nand U14325 (N_14325,N_13676,N_13579);
nor U14326 (N_14326,N_13909,N_13816);
nor U14327 (N_14327,N_13968,N_13521);
nor U14328 (N_14328,N_13508,N_13739);
or U14329 (N_14329,N_13610,N_13915);
and U14330 (N_14330,N_13804,N_13712);
nor U14331 (N_14331,N_13772,N_13871);
or U14332 (N_14332,N_13896,N_13878);
and U14333 (N_14333,N_13517,N_13847);
and U14334 (N_14334,N_13962,N_13829);
xor U14335 (N_14335,N_13506,N_13707);
and U14336 (N_14336,N_13768,N_13745);
nor U14337 (N_14337,N_13589,N_13985);
and U14338 (N_14338,N_13501,N_13954);
nor U14339 (N_14339,N_13675,N_13589);
or U14340 (N_14340,N_13946,N_13703);
xor U14341 (N_14341,N_13519,N_13504);
xnor U14342 (N_14342,N_13715,N_13728);
nand U14343 (N_14343,N_13810,N_13695);
xor U14344 (N_14344,N_13520,N_13598);
and U14345 (N_14345,N_13895,N_13886);
or U14346 (N_14346,N_13606,N_13622);
nand U14347 (N_14347,N_13600,N_13886);
nor U14348 (N_14348,N_13522,N_13620);
nor U14349 (N_14349,N_13840,N_13818);
nand U14350 (N_14350,N_13720,N_13855);
or U14351 (N_14351,N_13647,N_13930);
nand U14352 (N_14352,N_13742,N_13890);
xnor U14353 (N_14353,N_13525,N_13684);
or U14354 (N_14354,N_13572,N_13957);
nor U14355 (N_14355,N_13514,N_13818);
or U14356 (N_14356,N_13825,N_13569);
xnor U14357 (N_14357,N_13523,N_13896);
or U14358 (N_14358,N_13676,N_13567);
xnor U14359 (N_14359,N_13657,N_13555);
nand U14360 (N_14360,N_13876,N_13553);
nand U14361 (N_14361,N_13794,N_13641);
xnor U14362 (N_14362,N_13582,N_13686);
and U14363 (N_14363,N_13700,N_13889);
or U14364 (N_14364,N_13568,N_13909);
nand U14365 (N_14365,N_13700,N_13957);
nand U14366 (N_14366,N_13988,N_13849);
nand U14367 (N_14367,N_13802,N_13714);
and U14368 (N_14368,N_13650,N_13675);
nor U14369 (N_14369,N_13880,N_13846);
and U14370 (N_14370,N_13842,N_13804);
and U14371 (N_14371,N_13640,N_13674);
and U14372 (N_14372,N_13560,N_13523);
nor U14373 (N_14373,N_13566,N_13552);
xnor U14374 (N_14374,N_13881,N_13548);
nand U14375 (N_14375,N_13586,N_13564);
or U14376 (N_14376,N_13734,N_13739);
or U14377 (N_14377,N_13722,N_13564);
nand U14378 (N_14378,N_13768,N_13842);
xor U14379 (N_14379,N_13676,N_13798);
nor U14380 (N_14380,N_13981,N_13956);
nor U14381 (N_14381,N_13533,N_13786);
and U14382 (N_14382,N_13688,N_13614);
or U14383 (N_14383,N_13997,N_13574);
xnor U14384 (N_14384,N_13537,N_13583);
and U14385 (N_14385,N_13540,N_13645);
xor U14386 (N_14386,N_13811,N_13617);
or U14387 (N_14387,N_13634,N_13883);
nor U14388 (N_14388,N_13754,N_13587);
nand U14389 (N_14389,N_13761,N_13540);
nand U14390 (N_14390,N_13720,N_13550);
nand U14391 (N_14391,N_13699,N_13845);
xor U14392 (N_14392,N_13803,N_13952);
and U14393 (N_14393,N_13980,N_13656);
and U14394 (N_14394,N_13771,N_13682);
xnor U14395 (N_14395,N_13514,N_13832);
nand U14396 (N_14396,N_13772,N_13707);
nand U14397 (N_14397,N_13832,N_13665);
or U14398 (N_14398,N_13558,N_13652);
or U14399 (N_14399,N_13850,N_13688);
nor U14400 (N_14400,N_13632,N_13782);
and U14401 (N_14401,N_13994,N_13632);
xnor U14402 (N_14402,N_13992,N_13530);
and U14403 (N_14403,N_13830,N_13897);
nor U14404 (N_14404,N_13676,N_13915);
nor U14405 (N_14405,N_13851,N_13968);
nand U14406 (N_14406,N_13822,N_13561);
xnor U14407 (N_14407,N_13521,N_13570);
nand U14408 (N_14408,N_13547,N_13694);
xnor U14409 (N_14409,N_13896,N_13934);
nand U14410 (N_14410,N_13954,N_13625);
and U14411 (N_14411,N_13995,N_13801);
or U14412 (N_14412,N_13969,N_13601);
nor U14413 (N_14413,N_13701,N_13710);
and U14414 (N_14414,N_13747,N_13589);
nand U14415 (N_14415,N_13566,N_13567);
xnor U14416 (N_14416,N_13539,N_13871);
and U14417 (N_14417,N_13723,N_13707);
and U14418 (N_14418,N_13892,N_13787);
nand U14419 (N_14419,N_13685,N_13569);
xnor U14420 (N_14420,N_13874,N_13508);
and U14421 (N_14421,N_13562,N_13946);
xnor U14422 (N_14422,N_13527,N_13646);
xor U14423 (N_14423,N_13873,N_13816);
or U14424 (N_14424,N_13886,N_13722);
or U14425 (N_14425,N_13989,N_13673);
and U14426 (N_14426,N_13706,N_13864);
or U14427 (N_14427,N_13515,N_13873);
and U14428 (N_14428,N_13761,N_13888);
nand U14429 (N_14429,N_13841,N_13696);
xor U14430 (N_14430,N_13794,N_13875);
or U14431 (N_14431,N_13992,N_13977);
nor U14432 (N_14432,N_13688,N_13765);
or U14433 (N_14433,N_13655,N_13559);
and U14434 (N_14434,N_13520,N_13610);
xnor U14435 (N_14435,N_13859,N_13609);
and U14436 (N_14436,N_13598,N_13725);
nor U14437 (N_14437,N_13661,N_13879);
nand U14438 (N_14438,N_13961,N_13933);
or U14439 (N_14439,N_13657,N_13914);
nand U14440 (N_14440,N_13778,N_13951);
nand U14441 (N_14441,N_13872,N_13649);
nand U14442 (N_14442,N_13693,N_13500);
nor U14443 (N_14443,N_13851,N_13671);
xor U14444 (N_14444,N_13860,N_13858);
or U14445 (N_14445,N_13679,N_13653);
or U14446 (N_14446,N_13662,N_13946);
nor U14447 (N_14447,N_13629,N_13702);
or U14448 (N_14448,N_13886,N_13890);
xor U14449 (N_14449,N_13976,N_13942);
or U14450 (N_14450,N_13800,N_13790);
or U14451 (N_14451,N_13757,N_13516);
and U14452 (N_14452,N_13891,N_13781);
or U14453 (N_14453,N_13904,N_13999);
and U14454 (N_14454,N_13896,N_13979);
nor U14455 (N_14455,N_13735,N_13908);
nor U14456 (N_14456,N_13984,N_13728);
nand U14457 (N_14457,N_13980,N_13701);
nand U14458 (N_14458,N_13625,N_13872);
nand U14459 (N_14459,N_13828,N_13686);
and U14460 (N_14460,N_13542,N_13559);
or U14461 (N_14461,N_13597,N_13897);
xor U14462 (N_14462,N_13830,N_13956);
xor U14463 (N_14463,N_13692,N_13548);
nor U14464 (N_14464,N_13707,N_13511);
nor U14465 (N_14465,N_13714,N_13715);
nor U14466 (N_14466,N_13877,N_13594);
nor U14467 (N_14467,N_13725,N_13609);
or U14468 (N_14468,N_13876,N_13518);
xor U14469 (N_14469,N_13581,N_13500);
nor U14470 (N_14470,N_13958,N_13900);
or U14471 (N_14471,N_13705,N_13925);
or U14472 (N_14472,N_13746,N_13640);
nor U14473 (N_14473,N_13710,N_13929);
and U14474 (N_14474,N_13927,N_13885);
nand U14475 (N_14475,N_13590,N_13978);
or U14476 (N_14476,N_13866,N_13547);
and U14477 (N_14477,N_13632,N_13585);
nand U14478 (N_14478,N_13544,N_13612);
nor U14479 (N_14479,N_13563,N_13545);
nor U14480 (N_14480,N_13858,N_13989);
nand U14481 (N_14481,N_13957,N_13869);
nor U14482 (N_14482,N_13967,N_13605);
and U14483 (N_14483,N_13515,N_13689);
xnor U14484 (N_14484,N_13932,N_13925);
xnor U14485 (N_14485,N_13781,N_13660);
nor U14486 (N_14486,N_13576,N_13914);
nand U14487 (N_14487,N_13576,N_13907);
nor U14488 (N_14488,N_13997,N_13643);
and U14489 (N_14489,N_13884,N_13540);
nand U14490 (N_14490,N_13505,N_13968);
nand U14491 (N_14491,N_13926,N_13575);
nor U14492 (N_14492,N_13994,N_13962);
or U14493 (N_14493,N_13747,N_13704);
nand U14494 (N_14494,N_13845,N_13580);
nor U14495 (N_14495,N_13543,N_13562);
nand U14496 (N_14496,N_13565,N_13759);
nor U14497 (N_14497,N_13793,N_13936);
nand U14498 (N_14498,N_13850,N_13565);
nand U14499 (N_14499,N_13536,N_13844);
nand U14500 (N_14500,N_14196,N_14354);
xor U14501 (N_14501,N_14431,N_14271);
xor U14502 (N_14502,N_14363,N_14395);
nand U14503 (N_14503,N_14422,N_14236);
or U14504 (N_14504,N_14112,N_14106);
xnor U14505 (N_14505,N_14489,N_14254);
xnor U14506 (N_14506,N_14338,N_14324);
nand U14507 (N_14507,N_14207,N_14351);
xor U14508 (N_14508,N_14441,N_14307);
and U14509 (N_14509,N_14266,N_14358);
nor U14510 (N_14510,N_14239,N_14115);
nor U14511 (N_14511,N_14435,N_14326);
nor U14512 (N_14512,N_14290,N_14000);
or U14513 (N_14513,N_14490,N_14339);
xor U14514 (N_14514,N_14197,N_14301);
nand U14515 (N_14515,N_14285,N_14163);
nand U14516 (N_14516,N_14460,N_14274);
nand U14517 (N_14517,N_14204,N_14279);
nor U14518 (N_14518,N_14497,N_14401);
nand U14519 (N_14519,N_14015,N_14081);
and U14520 (N_14520,N_14117,N_14087);
or U14521 (N_14521,N_14437,N_14120);
xor U14522 (N_14522,N_14183,N_14073);
nor U14523 (N_14523,N_14213,N_14452);
xnor U14524 (N_14524,N_14461,N_14310);
or U14525 (N_14525,N_14295,N_14159);
nand U14526 (N_14526,N_14138,N_14165);
nor U14527 (N_14527,N_14039,N_14292);
or U14528 (N_14528,N_14424,N_14356);
or U14529 (N_14529,N_14051,N_14261);
nand U14530 (N_14530,N_14366,N_14203);
and U14531 (N_14531,N_14092,N_14294);
nor U14532 (N_14532,N_14030,N_14414);
or U14533 (N_14533,N_14089,N_14256);
xnor U14534 (N_14534,N_14355,N_14264);
nand U14535 (N_14535,N_14071,N_14245);
xnor U14536 (N_14536,N_14157,N_14387);
nor U14537 (N_14537,N_14146,N_14302);
and U14538 (N_14538,N_14369,N_14238);
nor U14539 (N_14539,N_14413,N_14468);
and U14540 (N_14540,N_14110,N_14291);
nor U14541 (N_14541,N_14058,N_14288);
and U14542 (N_14542,N_14373,N_14416);
nand U14543 (N_14543,N_14402,N_14017);
nor U14544 (N_14544,N_14091,N_14141);
nor U14545 (N_14545,N_14242,N_14477);
or U14546 (N_14546,N_14160,N_14020);
nand U14547 (N_14547,N_14080,N_14113);
nand U14548 (N_14548,N_14352,N_14337);
xor U14549 (N_14549,N_14098,N_14341);
or U14550 (N_14550,N_14144,N_14331);
nor U14551 (N_14551,N_14411,N_14140);
nor U14552 (N_14552,N_14483,N_14346);
and U14553 (N_14553,N_14170,N_14137);
nand U14554 (N_14554,N_14304,N_14225);
nor U14555 (N_14555,N_14206,N_14428);
xor U14556 (N_14556,N_14219,N_14066);
nor U14557 (N_14557,N_14313,N_14174);
xnor U14558 (N_14558,N_14485,N_14448);
or U14559 (N_14559,N_14190,N_14275);
or U14560 (N_14560,N_14166,N_14007);
xnor U14561 (N_14561,N_14226,N_14224);
and U14562 (N_14562,N_14014,N_14218);
and U14563 (N_14563,N_14364,N_14436);
nor U14564 (N_14564,N_14076,N_14316);
or U14565 (N_14565,N_14013,N_14379);
nor U14566 (N_14566,N_14357,N_14494);
xnor U14567 (N_14567,N_14067,N_14300);
or U14568 (N_14568,N_14037,N_14078);
nand U14569 (N_14569,N_14365,N_14367);
and U14570 (N_14570,N_14345,N_14398);
xor U14571 (N_14571,N_14147,N_14121);
nand U14572 (N_14572,N_14317,N_14488);
or U14573 (N_14573,N_14103,N_14195);
xor U14574 (N_14574,N_14096,N_14036);
nor U14575 (N_14575,N_14479,N_14077);
xor U14576 (N_14576,N_14168,N_14472);
xnor U14577 (N_14577,N_14027,N_14334);
and U14578 (N_14578,N_14045,N_14185);
nor U14579 (N_14579,N_14114,N_14247);
nand U14580 (N_14580,N_14393,N_14167);
xor U14581 (N_14581,N_14033,N_14131);
or U14582 (N_14582,N_14487,N_14056);
xor U14583 (N_14583,N_14377,N_14263);
and U14584 (N_14584,N_14212,N_14386);
or U14585 (N_14585,N_14123,N_14150);
nand U14586 (N_14586,N_14287,N_14122);
xor U14587 (N_14587,N_14199,N_14074);
nand U14588 (N_14588,N_14093,N_14278);
or U14589 (N_14589,N_14069,N_14068);
or U14590 (N_14590,N_14361,N_14409);
or U14591 (N_14591,N_14408,N_14156);
xnor U14592 (N_14592,N_14430,N_14025);
xnor U14593 (N_14593,N_14446,N_14153);
nand U14594 (N_14594,N_14133,N_14325);
nand U14595 (N_14595,N_14445,N_14423);
xnor U14596 (N_14596,N_14433,N_14396);
nand U14597 (N_14597,N_14223,N_14482);
xnor U14598 (N_14598,N_14250,N_14231);
or U14599 (N_14599,N_14155,N_14399);
nand U14600 (N_14600,N_14097,N_14029);
nand U14601 (N_14601,N_14297,N_14421);
nand U14602 (N_14602,N_14070,N_14440);
and U14603 (N_14603,N_14397,N_14130);
xor U14604 (N_14604,N_14032,N_14383);
and U14605 (N_14605,N_14062,N_14173);
xor U14606 (N_14606,N_14281,N_14273);
or U14607 (N_14607,N_14444,N_14205);
or U14608 (N_14608,N_14235,N_14178);
xnor U14609 (N_14609,N_14400,N_14450);
nor U14610 (N_14610,N_14349,N_14456);
or U14611 (N_14611,N_14284,N_14187);
and U14612 (N_14612,N_14362,N_14086);
xor U14613 (N_14613,N_14230,N_14127);
xor U14614 (N_14614,N_14063,N_14368);
nor U14615 (N_14615,N_14404,N_14006);
nor U14616 (N_14616,N_14001,N_14040);
nand U14617 (N_14617,N_14286,N_14403);
xor U14618 (N_14618,N_14289,N_14008);
xnor U14619 (N_14619,N_14049,N_14018);
and U14620 (N_14620,N_14299,N_14134);
nor U14621 (N_14621,N_14149,N_14493);
xnor U14622 (N_14622,N_14336,N_14449);
or U14623 (N_14623,N_14481,N_14272);
and U14624 (N_14624,N_14026,N_14139);
or U14625 (N_14625,N_14375,N_14392);
or U14626 (N_14626,N_14464,N_14151);
and U14627 (N_14627,N_14303,N_14312);
xnor U14628 (N_14628,N_14182,N_14003);
nand U14629 (N_14629,N_14405,N_14046);
nor U14630 (N_14630,N_14048,N_14469);
and U14631 (N_14631,N_14044,N_14038);
nor U14632 (N_14632,N_14220,N_14283);
xnor U14633 (N_14633,N_14463,N_14251);
nand U14634 (N_14634,N_14353,N_14010);
nand U14635 (N_14635,N_14216,N_14023);
or U14636 (N_14636,N_14330,N_14342);
and U14637 (N_14637,N_14109,N_14119);
and U14638 (N_14638,N_14169,N_14480);
xnor U14639 (N_14639,N_14360,N_14277);
and U14640 (N_14640,N_14496,N_14298);
and U14641 (N_14641,N_14060,N_14486);
or U14642 (N_14642,N_14466,N_14370);
nand U14643 (N_14643,N_14035,N_14154);
xnor U14644 (N_14644,N_14417,N_14193);
nor U14645 (N_14645,N_14255,N_14253);
xnor U14646 (N_14646,N_14012,N_14259);
nand U14647 (N_14647,N_14107,N_14410);
nor U14648 (N_14648,N_14495,N_14459);
or U14649 (N_14649,N_14455,N_14102);
xor U14650 (N_14650,N_14306,N_14427);
and U14651 (N_14651,N_14350,N_14391);
or U14652 (N_14652,N_14101,N_14432);
and U14653 (N_14653,N_14095,N_14234);
nor U14654 (N_14654,N_14210,N_14249);
nand U14655 (N_14655,N_14376,N_14343);
nand U14656 (N_14656,N_14308,N_14057);
nand U14657 (N_14657,N_14082,N_14378);
and U14658 (N_14658,N_14072,N_14471);
or U14659 (N_14659,N_14282,N_14004);
nor U14660 (N_14660,N_14053,N_14221);
or U14661 (N_14661,N_14229,N_14111);
xnor U14662 (N_14662,N_14333,N_14176);
or U14663 (N_14663,N_14108,N_14458);
and U14664 (N_14664,N_14269,N_14175);
and U14665 (N_14665,N_14415,N_14457);
nor U14666 (N_14666,N_14191,N_14055);
xnor U14667 (N_14667,N_14389,N_14258);
or U14668 (N_14668,N_14244,N_14246);
xor U14669 (N_14669,N_14009,N_14348);
nand U14670 (N_14670,N_14347,N_14498);
nand U14671 (N_14671,N_14184,N_14200);
xnor U14672 (N_14672,N_14188,N_14126);
nand U14673 (N_14673,N_14100,N_14328);
nand U14674 (N_14674,N_14314,N_14248);
nor U14675 (N_14675,N_14209,N_14124);
nor U14676 (N_14676,N_14390,N_14438);
and U14677 (N_14677,N_14474,N_14136);
nand U14678 (N_14678,N_14280,N_14252);
xnor U14679 (N_14679,N_14059,N_14181);
xor U14680 (N_14680,N_14104,N_14084);
or U14681 (N_14681,N_14262,N_14499);
or U14682 (N_14682,N_14233,N_14344);
and U14683 (N_14683,N_14476,N_14016);
or U14684 (N_14684,N_14443,N_14128);
and U14685 (N_14685,N_14359,N_14061);
and U14686 (N_14686,N_14478,N_14177);
nor U14687 (N_14687,N_14028,N_14371);
or U14688 (N_14688,N_14132,N_14142);
or U14689 (N_14689,N_14002,N_14276);
and U14690 (N_14690,N_14227,N_14215);
nor U14691 (N_14691,N_14434,N_14332);
xor U14692 (N_14692,N_14171,N_14083);
or U14693 (N_14693,N_14382,N_14462);
or U14694 (N_14694,N_14257,N_14047);
nand U14695 (N_14695,N_14412,N_14043);
nor U14696 (N_14696,N_14031,N_14473);
nor U14697 (N_14697,N_14315,N_14406);
and U14698 (N_14698,N_14372,N_14267);
or U14699 (N_14699,N_14237,N_14161);
nand U14700 (N_14700,N_14054,N_14322);
xor U14701 (N_14701,N_14075,N_14309);
and U14702 (N_14702,N_14208,N_14172);
and U14703 (N_14703,N_14129,N_14491);
or U14704 (N_14704,N_14320,N_14228);
nand U14705 (N_14705,N_14492,N_14327);
xor U14706 (N_14706,N_14042,N_14293);
nor U14707 (N_14707,N_14340,N_14394);
nor U14708 (N_14708,N_14214,N_14467);
xor U14709 (N_14709,N_14447,N_14011);
and U14710 (N_14710,N_14019,N_14268);
nor U14711 (N_14711,N_14374,N_14192);
nor U14712 (N_14712,N_14311,N_14194);
xnor U14713 (N_14713,N_14050,N_14270);
and U14714 (N_14714,N_14021,N_14380);
nor U14715 (N_14715,N_14381,N_14321);
nand U14716 (N_14716,N_14484,N_14202);
and U14717 (N_14717,N_14116,N_14426);
nor U14718 (N_14718,N_14085,N_14024);
and U14719 (N_14719,N_14319,N_14180);
and U14720 (N_14720,N_14454,N_14222);
nand U14721 (N_14721,N_14158,N_14419);
and U14722 (N_14722,N_14475,N_14041);
nand U14723 (N_14723,N_14198,N_14135);
xor U14724 (N_14724,N_14094,N_14145);
nand U14725 (N_14725,N_14052,N_14065);
xor U14726 (N_14726,N_14162,N_14453);
nor U14727 (N_14727,N_14470,N_14305);
nor U14728 (N_14728,N_14179,N_14451);
nand U14729 (N_14729,N_14323,N_14385);
nand U14730 (N_14730,N_14064,N_14240);
nor U14731 (N_14731,N_14211,N_14186);
xor U14732 (N_14732,N_14022,N_14425);
xor U14733 (N_14733,N_14034,N_14143);
and U14734 (N_14734,N_14241,N_14265);
or U14735 (N_14735,N_14335,N_14407);
nor U14736 (N_14736,N_14232,N_14105);
and U14737 (N_14737,N_14442,N_14099);
nor U14738 (N_14738,N_14152,N_14079);
or U14739 (N_14739,N_14189,N_14329);
and U14740 (N_14740,N_14118,N_14125);
and U14741 (N_14741,N_14088,N_14243);
or U14742 (N_14742,N_14148,N_14418);
nor U14743 (N_14743,N_14164,N_14429);
nor U14744 (N_14744,N_14388,N_14296);
and U14745 (N_14745,N_14439,N_14318);
or U14746 (N_14746,N_14384,N_14420);
nor U14747 (N_14747,N_14217,N_14260);
nand U14748 (N_14748,N_14090,N_14465);
and U14749 (N_14749,N_14201,N_14005);
nand U14750 (N_14750,N_14009,N_14037);
or U14751 (N_14751,N_14284,N_14476);
or U14752 (N_14752,N_14145,N_14455);
nand U14753 (N_14753,N_14490,N_14001);
xor U14754 (N_14754,N_14198,N_14275);
nand U14755 (N_14755,N_14360,N_14130);
nor U14756 (N_14756,N_14416,N_14078);
nand U14757 (N_14757,N_14312,N_14060);
or U14758 (N_14758,N_14215,N_14447);
nor U14759 (N_14759,N_14361,N_14166);
nor U14760 (N_14760,N_14018,N_14403);
nor U14761 (N_14761,N_14474,N_14441);
or U14762 (N_14762,N_14358,N_14142);
nor U14763 (N_14763,N_14372,N_14479);
xnor U14764 (N_14764,N_14249,N_14374);
or U14765 (N_14765,N_14496,N_14039);
or U14766 (N_14766,N_14472,N_14082);
nor U14767 (N_14767,N_14084,N_14282);
or U14768 (N_14768,N_14083,N_14146);
xor U14769 (N_14769,N_14461,N_14404);
and U14770 (N_14770,N_14058,N_14241);
or U14771 (N_14771,N_14366,N_14236);
or U14772 (N_14772,N_14027,N_14233);
and U14773 (N_14773,N_14113,N_14185);
or U14774 (N_14774,N_14252,N_14453);
and U14775 (N_14775,N_14491,N_14107);
or U14776 (N_14776,N_14132,N_14035);
nand U14777 (N_14777,N_14271,N_14083);
and U14778 (N_14778,N_14148,N_14472);
or U14779 (N_14779,N_14454,N_14394);
xnor U14780 (N_14780,N_14249,N_14246);
and U14781 (N_14781,N_14402,N_14126);
or U14782 (N_14782,N_14317,N_14038);
or U14783 (N_14783,N_14455,N_14465);
and U14784 (N_14784,N_14151,N_14481);
nand U14785 (N_14785,N_14026,N_14307);
nand U14786 (N_14786,N_14458,N_14121);
or U14787 (N_14787,N_14487,N_14472);
nor U14788 (N_14788,N_14279,N_14342);
and U14789 (N_14789,N_14341,N_14122);
nand U14790 (N_14790,N_14470,N_14454);
or U14791 (N_14791,N_14432,N_14271);
or U14792 (N_14792,N_14163,N_14151);
nor U14793 (N_14793,N_14272,N_14132);
nor U14794 (N_14794,N_14045,N_14218);
or U14795 (N_14795,N_14172,N_14352);
xor U14796 (N_14796,N_14296,N_14145);
and U14797 (N_14797,N_14072,N_14352);
nor U14798 (N_14798,N_14437,N_14455);
nand U14799 (N_14799,N_14074,N_14250);
xnor U14800 (N_14800,N_14211,N_14188);
xor U14801 (N_14801,N_14426,N_14017);
nand U14802 (N_14802,N_14351,N_14150);
or U14803 (N_14803,N_14299,N_14051);
nand U14804 (N_14804,N_14213,N_14234);
nor U14805 (N_14805,N_14271,N_14302);
and U14806 (N_14806,N_14104,N_14019);
nor U14807 (N_14807,N_14329,N_14164);
nor U14808 (N_14808,N_14281,N_14068);
nand U14809 (N_14809,N_14424,N_14105);
or U14810 (N_14810,N_14331,N_14047);
xnor U14811 (N_14811,N_14153,N_14404);
and U14812 (N_14812,N_14306,N_14167);
xnor U14813 (N_14813,N_14294,N_14106);
nor U14814 (N_14814,N_14485,N_14044);
nor U14815 (N_14815,N_14285,N_14242);
and U14816 (N_14816,N_14480,N_14261);
or U14817 (N_14817,N_14254,N_14008);
nand U14818 (N_14818,N_14315,N_14053);
nor U14819 (N_14819,N_14111,N_14306);
and U14820 (N_14820,N_14205,N_14283);
nor U14821 (N_14821,N_14153,N_14392);
xnor U14822 (N_14822,N_14221,N_14492);
nand U14823 (N_14823,N_14183,N_14097);
or U14824 (N_14824,N_14038,N_14292);
or U14825 (N_14825,N_14116,N_14210);
xnor U14826 (N_14826,N_14346,N_14043);
or U14827 (N_14827,N_14401,N_14063);
nand U14828 (N_14828,N_14164,N_14298);
or U14829 (N_14829,N_14133,N_14390);
and U14830 (N_14830,N_14493,N_14153);
nor U14831 (N_14831,N_14012,N_14331);
or U14832 (N_14832,N_14243,N_14387);
nand U14833 (N_14833,N_14369,N_14227);
or U14834 (N_14834,N_14276,N_14244);
nand U14835 (N_14835,N_14459,N_14284);
nand U14836 (N_14836,N_14084,N_14130);
or U14837 (N_14837,N_14051,N_14286);
and U14838 (N_14838,N_14038,N_14030);
and U14839 (N_14839,N_14333,N_14458);
nor U14840 (N_14840,N_14214,N_14230);
nand U14841 (N_14841,N_14154,N_14229);
xor U14842 (N_14842,N_14111,N_14031);
xnor U14843 (N_14843,N_14208,N_14311);
nand U14844 (N_14844,N_14345,N_14377);
xnor U14845 (N_14845,N_14263,N_14060);
nand U14846 (N_14846,N_14442,N_14195);
and U14847 (N_14847,N_14266,N_14466);
nor U14848 (N_14848,N_14401,N_14115);
nand U14849 (N_14849,N_14232,N_14158);
xor U14850 (N_14850,N_14122,N_14473);
or U14851 (N_14851,N_14031,N_14011);
xor U14852 (N_14852,N_14141,N_14131);
nor U14853 (N_14853,N_14270,N_14460);
and U14854 (N_14854,N_14193,N_14391);
nand U14855 (N_14855,N_14067,N_14170);
or U14856 (N_14856,N_14295,N_14484);
and U14857 (N_14857,N_14256,N_14010);
xor U14858 (N_14858,N_14314,N_14408);
nand U14859 (N_14859,N_14012,N_14124);
and U14860 (N_14860,N_14462,N_14021);
or U14861 (N_14861,N_14169,N_14419);
xnor U14862 (N_14862,N_14171,N_14186);
and U14863 (N_14863,N_14386,N_14003);
nor U14864 (N_14864,N_14345,N_14180);
xnor U14865 (N_14865,N_14462,N_14241);
xnor U14866 (N_14866,N_14186,N_14491);
nand U14867 (N_14867,N_14406,N_14029);
and U14868 (N_14868,N_14009,N_14343);
nand U14869 (N_14869,N_14231,N_14430);
and U14870 (N_14870,N_14078,N_14208);
nor U14871 (N_14871,N_14327,N_14457);
and U14872 (N_14872,N_14270,N_14216);
nand U14873 (N_14873,N_14373,N_14223);
or U14874 (N_14874,N_14107,N_14197);
xnor U14875 (N_14875,N_14220,N_14005);
xnor U14876 (N_14876,N_14036,N_14126);
nand U14877 (N_14877,N_14142,N_14498);
nor U14878 (N_14878,N_14253,N_14317);
nand U14879 (N_14879,N_14484,N_14007);
or U14880 (N_14880,N_14056,N_14229);
and U14881 (N_14881,N_14194,N_14289);
and U14882 (N_14882,N_14190,N_14413);
nand U14883 (N_14883,N_14014,N_14026);
and U14884 (N_14884,N_14328,N_14176);
nand U14885 (N_14885,N_14190,N_14132);
xnor U14886 (N_14886,N_14425,N_14059);
and U14887 (N_14887,N_14288,N_14045);
or U14888 (N_14888,N_14438,N_14245);
nand U14889 (N_14889,N_14011,N_14482);
xor U14890 (N_14890,N_14475,N_14119);
or U14891 (N_14891,N_14196,N_14195);
nand U14892 (N_14892,N_14477,N_14215);
nor U14893 (N_14893,N_14468,N_14260);
nand U14894 (N_14894,N_14460,N_14326);
xor U14895 (N_14895,N_14049,N_14470);
xor U14896 (N_14896,N_14098,N_14066);
nor U14897 (N_14897,N_14414,N_14175);
and U14898 (N_14898,N_14359,N_14433);
or U14899 (N_14899,N_14046,N_14048);
nor U14900 (N_14900,N_14111,N_14407);
and U14901 (N_14901,N_14138,N_14205);
and U14902 (N_14902,N_14490,N_14329);
xor U14903 (N_14903,N_14461,N_14355);
or U14904 (N_14904,N_14218,N_14445);
xnor U14905 (N_14905,N_14050,N_14319);
nor U14906 (N_14906,N_14434,N_14144);
nor U14907 (N_14907,N_14229,N_14474);
nand U14908 (N_14908,N_14092,N_14327);
nor U14909 (N_14909,N_14193,N_14055);
nand U14910 (N_14910,N_14140,N_14000);
nand U14911 (N_14911,N_14106,N_14066);
and U14912 (N_14912,N_14236,N_14281);
or U14913 (N_14913,N_14141,N_14092);
or U14914 (N_14914,N_14179,N_14309);
and U14915 (N_14915,N_14448,N_14353);
nor U14916 (N_14916,N_14338,N_14250);
or U14917 (N_14917,N_14202,N_14364);
nor U14918 (N_14918,N_14141,N_14307);
and U14919 (N_14919,N_14127,N_14152);
and U14920 (N_14920,N_14397,N_14495);
nor U14921 (N_14921,N_14312,N_14030);
nand U14922 (N_14922,N_14478,N_14453);
or U14923 (N_14923,N_14103,N_14141);
nor U14924 (N_14924,N_14290,N_14148);
nand U14925 (N_14925,N_14127,N_14098);
xnor U14926 (N_14926,N_14356,N_14087);
xor U14927 (N_14927,N_14076,N_14069);
nor U14928 (N_14928,N_14277,N_14191);
xnor U14929 (N_14929,N_14221,N_14383);
nand U14930 (N_14930,N_14105,N_14483);
or U14931 (N_14931,N_14250,N_14168);
xor U14932 (N_14932,N_14082,N_14312);
xnor U14933 (N_14933,N_14275,N_14037);
xnor U14934 (N_14934,N_14202,N_14195);
or U14935 (N_14935,N_14009,N_14308);
or U14936 (N_14936,N_14211,N_14448);
and U14937 (N_14937,N_14161,N_14462);
and U14938 (N_14938,N_14151,N_14224);
nand U14939 (N_14939,N_14213,N_14140);
nand U14940 (N_14940,N_14334,N_14241);
xnor U14941 (N_14941,N_14310,N_14316);
nor U14942 (N_14942,N_14244,N_14499);
nand U14943 (N_14943,N_14156,N_14231);
or U14944 (N_14944,N_14403,N_14023);
and U14945 (N_14945,N_14048,N_14429);
or U14946 (N_14946,N_14321,N_14232);
xnor U14947 (N_14947,N_14229,N_14432);
nor U14948 (N_14948,N_14067,N_14241);
xor U14949 (N_14949,N_14479,N_14317);
nor U14950 (N_14950,N_14254,N_14314);
nand U14951 (N_14951,N_14495,N_14329);
and U14952 (N_14952,N_14155,N_14352);
and U14953 (N_14953,N_14499,N_14196);
xor U14954 (N_14954,N_14387,N_14454);
and U14955 (N_14955,N_14092,N_14313);
xnor U14956 (N_14956,N_14261,N_14156);
xnor U14957 (N_14957,N_14051,N_14222);
and U14958 (N_14958,N_14076,N_14478);
or U14959 (N_14959,N_14020,N_14076);
and U14960 (N_14960,N_14091,N_14359);
nand U14961 (N_14961,N_14130,N_14396);
nand U14962 (N_14962,N_14364,N_14431);
xnor U14963 (N_14963,N_14101,N_14056);
xnor U14964 (N_14964,N_14250,N_14103);
nand U14965 (N_14965,N_14265,N_14416);
xor U14966 (N_14966,N_14307,N_14234);
xnor U14967 (N_14967,N_14371,N_14131);
and U14968 (N_14968,N_14221,N_14347);
nor U14969 (N_14969,N_14436,N_14459);
nor U14970 (N_14970,N_14062,N_14338);
nand U14971 (N_14971,N_14174,N_14119);
or U14972 (N_14972,N_14431,N_14031);
nor U14973 (N_14973,N_14431,N_14218);
or U14974 (N_14974,N_14144,N_14103);
and U14975 (N_14975,N_14368,N_14437);
nand U14976 (N_14976,N_14400,N_14119);
or U14977 (N_14977,N_14083,N_14414);
nor U14978 (N_14978,N_14484,N_14128);
or U14979 (N_14979,N_14482,N_14438);
nand U14980 (N_14980,N_14295,N_14066);
nand U14981 (N_14981,N_14458,N_14361);
or U14982 (N_14982,N_14271,N_14318);
or U14983 (N_14983,N_14281,N_14260);
nand U14984 (N_14984,N_14068,N_14383);
and U14985 (N_14985,N_14063,N_14267);
xor U14986 (N_14986,N_14355,N_14283);
or U14987 (N_14987,N_14339,N_14186);
or U14988 (N_14988,N_14188,N_14488);
xnor U14989 (N_14989,N_14388,N_14154);
or U14990 (N_14990,N_14199,N_14004);
nor U14991 (N_14991,N_14146,N_14010);
and U14992 (N_14992,N_14471,N_14329);
nor U14993 (N_14993,N_14046,N_14082);
and U14994 (N_14994,N_14432,N_14081);
or U14995 (N_14995,N_14277,N_14134);
or U14996 (N_14996,N_14494,N_14472);
nor U14997 (N_14997,N_14040,N_14202);
nand U14998 (N_14998,N_14047,N_14045);
nor U14999 (N_14999,N_14174,N_14275);
or U15000 (N_15000,N_14553,N_14878);
nand U15001 (N_15001,N_14538,N_14778);
and U15002 (N_15002,N_14913,N_14510);
and U15003 (N_15003,N_14663,N_14699);
nor U15004 (N_15004,N_14679,N_14896);
nor U15005 (N_15005,N_14862,N_14639);
nor U15006 (N_15006,N_14861,N_14695);
or U15007 (N_15007,N_14953,N_14536);
nor U15008 (N_15008,N_14543,N_14572);
and U15009 (N_15009,N_14783,N_14689);
and U15010 (N_15010,N_14566,N_14730);
nand U15011 (N_15011,N_14869,N_14844);
or U15012 (N_15012,N_14751,N_14902);
or U15013 (N_15013,N_14574,N_14777);
or U15014 (N_15014,N_14959,N_14788);
nor U15015 (N_15015,N_14764,N_14883);
nor U15016 (N_15016,N_14700,N_14993);
and U15017 (N_15017,N_14654,N_14938);
nor U15018 (N_15018,N_14604,N_14998);
and U15019 (N_15019,N_14534,N_14637);
and U15020 (N_15020,N_14602,N_14759);
nand U15021 (N_15021,N_14752,N_14592);
nor U15022 (N_15022,N_14780,N_14791);
xor U15023 (N_15023,N_14607,N_14640);
nor U15024 (N_15024,N_14939,N_14580);
and U15025 (N_15025,N_14564,N_14990);
and U15026 (N_15026,N_14765,N_14531);
nand U15027 (N_15027,N_14545,N_14682);
or U15028 (N_15028,N_14879,N_14694);
nand U15029 (N_15029,N_14641,N_14949);
nand U15030 (N_15030,N_14661,N_14827);
xor U15031 (N_15031,N_14808,N_14926);
and U15032 (N_15032,N_14519,N_14824);
or U15033 (N_15033,N_14756,N_14611);
nand U15034 (N_15034,N_14721,N_14810);
or U15035 (N_15035,N_14528,N_14658);
nand U15036 (N_15036,N_14979,N_14763);
nor U15037 (N_15037,N_14889,N_14985);
and U15038 (N_15038,N_14718,N_14908);
and U15039 (N_15039,N_14547,N_14933);
nand U15040 (N_15040,N_14505,N_14921);
nor U15041 (N_15041,N_14729,N_14923);
nor U15042 (N_15042,N_14669,N_14762);
or U15043 (N_15043,N_14606,N_14631);
or U15044 (N_15044,N_14868,N_14976);
xnor U15045 (N_15045,N_14743,N_14915);
nor U15046 (N_15046,N_14712,N_14713);
nand U15047 (N_15047,N_14825,N_14530);
and U15048 (N_15048,N_14533,N_14680);
and U15049 (N_15049,N_14821,N_14685);
and U15050 (N_15050,N_14974,N_14969);
and U15051 (N_15051,N_14683,N_14761);
nor U15052 (N_15052,N_14818,N_14942);
nand U15053 (N_15053,N_14556,N_14892);
nand U15054 (N_15054,N_14623,N_14583);
nand U15055 (N_15055,N_14850,N_14677);
xor U15056 (N_15056,N_14706,N_14906);
nand U15057 (N_15057,N_14571,N_14946);
and U15058 (N_15058,N_14829,N_14582);
or U15059 (N_15059,N_14613,N_14676);
xor U15060 (N_15060,N_14554,N_14831);
and U15061 (N_15061,N_14665,N_14684);
nand U15062 (N_15062,N_14912,N_14612);
or U15063 (N_15063,N_14725,N_14715);
nand U15064 (N_15064,N_14900,N_14708);
nor U15065 (N_15065,N_14941,N_14903);
and U15066 (N_15066,N_14872,N_14935);
xor U15067 (N_15067,N_14659,N_14595);
or U15068 (N_15068,N_14506,N_14773);
nor U15069 (N_15069,N_14522,N_14551);
nand U15070 (N_15070,N_14964,N_14717);
or U15071 (N_15071,N_14890,N_14855);
nand U15072 (N_15072,N_14688,N_14512);
nand U15073 (N_15073,N_14845,N_14738);
nand U15074 (N_15074,N_14875,N_14650);
or U15075 (N_15075,N_14884,N_14853);
nor U15076 (N_15076,N_14747,N_14815);
nor U15077 (N_15077,N_14877,N_14834);
and U15078 (N_15078,N_14876,N_14775);
nand U15079 (N_15079,N_14901,N_14995);
nor U15080 (N_15080,N_14922,N_14793);
and U15081 (N_15081,N_14958,N_14576);
and U15082 (N_15082,N_14568,N_14649);
xor U15083 (N_15083,N_14956,N_14806);
or U15084 (N_15084,N_14809,N_14513);
nand U15085 (N_15085,N_14776,N_14714);
xor U15086 (N_15086,N_14803,N_14916);
nor U15087 (N_15087,N_14696,N_14739);
or U15088 (N_15088,N_14924,N_14502);
nor U15089 (N_15089,N_14811,N_14526);
and U15090 (N_15090,N_14962,N_14929);
and U15091 (N_15091,N_14863,N_14873);
xnor U15092 (N_15092,N_14711,N_14973);
xor U15093 (N_15093,N_14947,N_14702);
nor U15094 (N_15094,N_14591,N_14521);
and U15095 (N_15095,N_14820,N_14804);
xor U15096 (N_15096,N_14828,N_14617);
xor U15097 (N_15097,N_14507,N_14629);
nor U15098 (N_15098,N_14544,N_14887);
nand U15099 (N_15099,N_14838,N_14609);
and U15100 (N_15100,N_14552,N_14523);
nand U15101 (N_15101,N_14532,N_14678);
and U15102 (N_15102,N_14529,N_14546);
or U15103 (N_15103,N_14894,N_14588);
or U15104 (N_15104,N_14646,N_14871);
or U15105 (N_15105,N_14686,N_14614);
or U15106 (N_15106,N_14563,N_14594);
and U15107 (N_15107,N_14636,N_14643);
nand U15108 (N_15108,N_14920,N_14874);
nand U15109 (N_15109,N_14832,N_14549);
nand U15110 (N_15110,N_14540,N_14570);
and U15111 (N_15111,N_14585,N_14774);
or U15112 (N_15112,N_14746,N_14726);
or U15113 (N_15113,N_14798,N_14977);
or U15114 (N_15114,N_14928,N_14535);
nor U15115 (N_15115,N_14660,N_14560);
or U15116 (N_15116,N_14899,N_14772);
and U15117 (N_15117,N_14737,N_14662);
nor U15118 (N_15118,N_14754,N_14504);
and U15119 (N_15119,N_14945,N_14885);
nor U15120 (N_15120,N_14794,N_14757);
nor U15121 (N_15121,N_14787,N_14517);
or U15122 (N_15122,N_14800,N_14734);
or U15123 (N_15123,N_14954,N_14710);
nor U15124 (N_15124,N_14723,N_14842);
and U15125 (N_15125,N_14657,N_14673);
and U15126 (N_15126,N_14701,N_14854);
or U15127 (N_15127,N_14625,N_14852);
or U15128 (N_15128,N_14860,N_14849);
or U15129 (N_15129,N_14719,N_14742);
nor U15130 (N_15130,N_14988,N_14681);
or U15131 (N_15131,N_14904,N_14830);
nor U15132 (N_15132,N_14771,N_14927);
or U15133 (N_15133,N_14652,N_14967);
xnor U15134 (N_15134,N_14603,N_14666);
nand U15135 (N_15135,N_14668,N_14596);
nor U15136 (N_15136,N_14720,N_14950);
nor U15137 (N_15137,N_14909,N_14630);
nor U15138 (N_15138,N_14575,N_14741);
nand U15139 (N_15139,N_14760,N_14981);
xor U15140 (N_15140,N_14848,N_14598);
nand U15141 (N_15141,N_14968,N_14870);
and U15142 (N_15142,N_14881,N_14687);
or U15143 (N_15143,N_14722,N_14664);
xor U15144 (N_15144,N_14690,N_14667);
nor U15145 (N_15145,N_14727,N_14886);
nor U15146 (N_15146,N_14785,N_14500);
or U15147 (N_15147,N_14621,N_14936);
xnor U15148 (N_15148,N_14655,N_14514);
and U15149 (N_15149,N_14907,N_14593);
nor U15150 (N_15150,N_14579,N_14561);
nand U15151 (N_15151,N_14578,N_14786);
nor U15152 (N_15152,N_14704,N_14557);
nand U15153 (N_15153,N_14618,N_14893);
and U15154 (N_15154,N_14565,N_14835);
nor U15155 (N_15155,N_14693,N_14980);
or U15156 (N_15156,N_14724,N_14731);
nand U15157 (N_15157,N_14882,N_14841);
nor U15158 (N_15158,N_14816,N_14697);
nand U15159 (N_15159,N_14635,N_14952);
nand U15160 (N_15160,N_14823,N_14846);
or U15161 (N_15161,N_14653,N_14638);
xor U15162 (N_15162,N_14840,N_14957);
nand U15163 (N_15163,N_14895,N_14856);
nand U15164 (N_15164,N_14897,N_14867);
nor U15165 (N_15165,N_14975,N_14991);
or U15166 (N_15166,N_14733,N_14511);
nand U15167 (N_15167,N_14509,N_14750);
nand U15168 (N_15168,N_14801,N_14632);
and U15169 (N_15169,N_14891,N_14698);
xor U15170 (N_15170,N_14753,N_14758);
nand U15171 (N_15171,N_14672,N_14642);
or U15172 (N_15172,N_14779,N_14930);
and U15173 (N_15173,N_14826,N_14501);
nand U15174 (N_15174,N_14911,N_14709);
and U15175 (N_15175,N_14971,N_14656);
nor U15176 (N_15176,N_14813,N_14802);
nand U15177 (N_15177,N_14864,N_14932);
or U15178 (N_15178,N_14955,N_14768);
and U15179 (N_15179,N_14518,N_14749);
nand U15180 (N_15180,N_14705,N_14624);
nand U15181 (N_15181,N_14986,N_14951);
nand U15182 (N_15182,N_14859,N_14965);
or U15183 (N_15183,N_14766,N_14542);
xor U15184 (N_15184,N_14740,N_14790);
nand U15185 (N_15185,N_14917,N_14931);
and U15186 (N_15186,N_14966,N_14847);
and U15187 (N_15187,N_14960,N_14888);
or U15188 (N_15188,N_14914,N_14516);
and U15189 (N_15189,N_14691,N_14910);
nor U15190 (N_15190,N_14515,N_14994);
or U15191 (N_15191,N_14807,N_14732);
or U15192 (N_15192,N_14628,N_14525);
and U15193 (N_15193,N_14999,N_14984);
nor U15194 (N_15194,N_14608,N_14537);
or U15195 (N_15195,N_14634,N_14944);
nor U15196 (N_15196,N_14992,N_14978);
or U15197 (N_15197,N_14918,N_14550);
or U15198 (N_15198,N_14796,N_14805);
and U15199 (N_15199,N_14674,N_14728);
nor U15200 (N_15200,N_14940,N_14548);
or U15201 (N_15201,N_14972,N_14937);
xor U15202 (N_15202,N_14586,N_14919);
xnor U15203 (N_15203,N_14851,N_14970);
xnor U15204 (N_15204,N_14735,N_14843);
xor U15205 (N_15205,N_14792,N_14997);
nand U15206 (N_15206,N_14627,N_14836);
nor U15207 (N_15207,N_14616,N_14648);
xnor U15208 (N_15208,N_14633,N_14541);
and U15209 (N_15209,N_14577,N_14716);
nor U15210 (N_15210,N_14782,N_14584);
nand U15211 (N_15211,N_14597,N_14934);
nor U15212 (N_15212,N_14527,N_14589);
nor U15213 (N_15213,N_14569,N_14814);
or U15214 (N_15214,N_14865,N_14620);
xnor U15215 (N_15215,N_14590,N_14619);
nand U15216 (N_15216,N_14989,N_14562);
nor U15217 (N_15217,N_14671,N_14622);
nor U15218 (N_15218,N_14670,N_14558);
nor U15219 (N_15219,N_14819,N_14898);
xnor U15220 (N_15220,N_14755,N_14797);
nor U15221 (N_15221,N_14744,N_14767);
nand U15222 (N_15222,N_14996,N_14839);
or U15223 (N_15223,N_14781,N_14795);
or U15224 (N_15224,N_14858,N_14605);
or U15225 (N_15225,N_14567,N_14880);
or U15226 (N_15226,N_14520,N_14905);
and U15227 (N_15227,N_14770,N_14703);
nor U15228 (N_15228,N_14539,N_14748);
or U15229 (N_15229,N_14987,N_14982);
nand U15230 (N_15230,N_14817,N_14857);
or U15231 (N_15231,N_14822,N_14837);
or U15232 (N_15232,N_14789,N_14581);
and U15233 (N_15233,N_14769,N_14692);
nor U15234 (N_15234,N_14508,N_14645);
or U15235 (N_15235,N_14925,N_14963);
xnor U15236 (N_15236,N_14524,N_14587);
nand U15237 (N_15237,N_14866,N_14745);
xor U15238 (N_15238,N_14833,N_14555);
or U15239 (N_15239,N_14647,N_14599);
xnor U15240 (N_15240,N_14503,N_14600);
and U15241 (N_15241,N_14983,N_14601);
or U15242 (N_15242,N_14943,N_14626);
xor U15243 (N_15243,N_14812,N_14675);
nor U15244 (N_15244,N_14799,N_14615);
or U15245 (N_15245,N_14573,N_14784);
and U15246 (N_15246,N_14559,N_14948);
or U15247 (N_15247,N_14736,N_14707);
and U15248 (N_15248,N_14644,N_14651);
or U15249 (N_15249,N_14610,N_14961);
or U15250 (N_15250,N_14707,N_14982);
nor U15251 (N_15251,N_14628,N_14638);
or U15252 (N_15252,N_14893,N_14558);
nor U15253 (N_15253,N_14852,N_14967);
nand U15254 (N_15254,N_14566,N_14771);
nand U15255 (N_15255,N_14588,N_14594);
xnor U15256 (N_15256,N_14817,N_14834);
nor U15257 (N_15257,N_14551,N_14826);
nor U15258 (N_15258,N_14525,N_14887);
and U15259 (N_15259,N_14643,N_14739);
nor U15260 (N_15260,N_14741,N_14862);
xor U15261 (N_15261,N_14745,N_14614);
nor U15262 (N_15262,N_14957,N_14931);
and U15263 (N_15263,N_14659,N_14520);
nor U15264 (N_15264,N_14639,N_14760);
xnor U15265 (N_15265,N_14528,N_14706);
nand U15266 (N_15266,N_14944,N_14750);
nand U15267 (N_15267,N_14563,N_14760);
or U15268 (N_15268,N_14914,N_14549);
xor U15269 (N_15269,N_14618,N_14779);
xnor U15270 (N_15270,N_14893,N_14938);
and U15271 (N_15271,N_14699,N_14971);
nor U15272 (N_15272,N_14943,N_14825);
nand U15273 (N_15273,N_14723,N_14939);
nand U15274 (N_15274,N_14786,N_14639);
nand U15275 (N_15275,N_14620,N_14875);
nand U15276 (N_15276,N_14785,N_14813);
nor U15277 (N_15277,N_14527,N_14627);
nor U15278 (N_15278,N_14812,N_14933);
nor U15279 (N_15279,N_14936,N_14954);
xnor U15280 (N_15280,N_14919,N_14754);
and U15281 (N_15281,N_14897,N_14835);
and U15282 (N_15282,N_14781,N_14638);
and U15283 (N_15283,N_14632,N_14636);
xor U15284 (N_15284,N_14800,N_14801);
xnor U15285 (N_15285,N_14640,N_14526);
and U15286 (N_15286,N_14977,N_14952);
nor U15287 (N_15287,N_14914,N_14581);
and U15288 (N_15288,N_14741,N_14557);
xor U15289 (N_15289,N_14832,N_14585);
nand U15290 (N_15290,N_14627,N_14737);
and U15291 (N_15291,N_14582,N_14975);
xnor U15292 (N_15292,N_14600,N_14734);
xnor U15293 (N_15293,N_14943,N_14572);
or U15294 (N_15294,N_14840,N_14609);
nor U15295 (N_15295,N_14639,N_14662);
nor U15296 (N_15296,N_14926,N_14940);
nor U15297 (N_15297,N_14642,N_14815);
nand U15298 (N_15298,N_14849,N_14597);
and U15299 (N_15299,N_14601,N_14643);
nand U15300 (N_15300,N_14673,N_14600);
xor U15301 (N_15301,N_14885,N_14704);
xor U15302 (N_15302,N_14547,N_14697);
xnor U15303 (N_15303,N_14650,N_14963);
xor U15304 (N_15304,N_14885,N_14809);
nor U15305 (N_15305,N_14907,N_14737);
and U15306 (N_15306,N_14965,N_14869);
and U15307 (N_15307,N_14892,N_14907);
xor U15308 (N_15308,N_14736,N_14864);
nand U15309 (N_15309,N_14835,N_14596);
nand U15310 (N_15310,N_14807,N_14533);
and U15311 (N_15311,N_14654,N_14622);
xnor U15312 (N_15312,N_14938,N_14510);
or U15313 (N_15313,N_14740,N_14709);
and U15314 (N_15314,N_14510,N_14940);
xor U15315 (N_15315,N_14850,N_14564);
nor U15316 (N_15316,N_14610,N_14920);
nand U15317 (N_15317,N_14738,N_14849);
xor U15318 (N_15318,N_14504,N_14934);
nor U15319 (N_15319,N_14564,N_14705);
nor U15320 (N_15320,N_14742,N_14908);
nor U15321 (N_15321,N_14635,N_14973);
or U15322 (N_15322,N_14582,N_14746);
and U15323 (N_15323,N_14781,N_14761);
or U15324 (N_15324,N_14937,N_14711);
nand U15325 (N_15325,N_14668,N_14833);
xnor U15326 (N_15326,N_14753,N_14772);
nor U15327 (N_15327,N_14583,N_14775);
xnor U15328 (N_15328,N_14680,N_14937);
or U15329 (N_15329,N_14986,N_14557);
and U15330 (N_15330,N_14615,N_14877);
nor U15331 (N_15331,N_14986,N_14846);
xnor U15332 (N_15332,N_14989,N_14877);
or U15333 (N_15333,N_14903,N_14514);
or U15334 (N_15334,N_14960,N_14950);
or U15335 (N_15335,N_14922,N_14866);
or U15336 (N_15336,N_14624,N_14870);
and U15337 (N_15337,N_14873,N_14791);
xnor U15338 (N_15338,N_14953,N_14737);
or U15339 (N_15339,N_14767,N_14880);
and U15340 (N_15340,N_14539,N_14717);
and U15341 (N_15341,N_14690,N_14518);
and U15342 (N_15342,N_14545,N_14998);
nor U15343 (N_15343,N_14550,N_14628);
nand U15344 (N_15344,N_14505,N_14561);
xnor U15345 (N_15345,N_14537,N_14632);
nand U15346 (N_15346,N_14886,N_14847);
xor U15347 (N_15347,N_14610,N_14740);
nand U15348 (N_15348,N_14590,N_14670);
or U15349 (N_15349,N_14543,N_14696);
nand U15350 (N_15350,N_14803,N_14771);
xor U15351 (N_15351,N_14534,N_14954);
xnor U15352 (N_15352,N_14628,N_14606);
nor U15353 (N_15353,N_14572,N_14938);
nand U15354 (N_15354,N_14737,N_14513);
nand U15355 (N_15355,N_14709,N_14923);
xnor U15356 (N_15356,N_14767,N_14690);
nand U15357 (N_15357,N_14618,N_14671);
nor U15358 (N_15358,N_14930,N_14858);
xor U15359 (N_15359,N_14929,N_14688);
and U15360 (N_15360,N_14500,N_14827);
nor U15361 (N_15361,N_14800,N_14959);
and U15362 (N_15362,N_14835,N_14797);
and U15363 (N_15363,N_14621,N_14637);
or U15364 (N_15364,N_14668,N_14547);
xnor U15365 (N_15365,N_14542,N_14822);
nand U15366 (N_15366,N_14931,N_14552);
or U15367 (N_15367,N_14542,N_14588);
xnor U15368 (N_15368,N_14999,N_14886);
or U15369 (N_15369,N_14723,N_14652);
nor U15370 (N_15370,N_14797,N_14596);
nand U15371 (N_15371,N_14746,N_14868);
and U15372 (N_15372,N_14865,N_14755);
xor U15373 (N_15373,N_14798,N_14897);
nand U15374 (N_15374,N_14594,N_14914);
nor U15375 (N_15375,N_14655,N_14704);
xor U15376 (N_15376,N_14970,N_14825);
xor U15377 (N_15377,N_14962,N_14507);
and U15378 (N_15378,N_14527,N_14984);
xor U15379 (N_15379,N_14623,N_14740);
xor U15380 (N_15380,N_14676,N_14627);
nand U15381 (N_15381,N_14751,N_14579);
or U15382 (N_15382,N_14717,N_14608);
nand U15383 (N_15383,N_14981,N_14511);
or U15384 (N_15384,N_14821,N_14776);
xor U15385 (N_15385,N_14718,N_14647);
nor U15386 (N_15386,N_14684,N_14640);
xor U15387 (N_15387,N_14554,N_14734);
nand U15388 (N_15388,N_14589,N_14762);
or U15389 (N_15389,N_14522,N_14825);
and U15390 (N_15390,N_14543,N_14776);
nor U15391 (N_15391,N_14819,N_14604);
nand U15392 (N_15392,N_14907,N_14872);
nor U15393 (N_15393,N_14537,N_14662);
or U15394 (N_15394,N_14715,N_14924);
or U15395 (N_15395,N_14955,N_14655);
xnor U15396 (N_15396,N_14759,N_14537);
xor U15397 (N_15397,N_14665,N_14954);
xnor U15398 (N_15398,N_14515,N_14707);
xor U15399 (N_15399,N_14820,N_14786);
nand U15400 (N_15400,N_14753,N_14802);
nand U15401 (N_15401,N_14926,N_14619);
and U15402 (N_15402,N_14831,N_14902);
and U15403 (N_15403,N_14514,N_14952);
and U15404 (N_15404,N_14724,N_14635);
or U15405 (N_15405,N_14805,N_14748);
or U15406 (N_15406,N_14570,N_14605);
or U15407 (N_15407,N_14635,N_14905);
nand U15408 (N_15408,N_14652,N_14903);
nor U15409 (N_15409,N_14894,N_14885);
nor U15410 (N_15410,N_14915,N_14741);
or U15411 (N_15411,N_14729,N_14723);
and U15412 (N_15412,N_14862,N_14817);
and U15413 (N_15413,N_14596,N_14772);
nor U15414 (N_15414,N_14811,N_14815);
or U15415 (N_15415,N_14882,N_14622);
nor U15416 (N_15416,N_14998,N_14781);
xnor U15417 (N_15417,N_14891,N_14941);
or U15418 (N_15418,N_14828,N_14734);
xor U15419 (N_15419,N_14627,N_14882);
nand U15420 (N_15420,N_14864,N_14807);
and U15421 (N_15421,N_14850,N_14605);
xnor U15422 (N_15422,N_14890,N_14672);
nand U15423 (N_15423,N_14513,N_14715);
nor U15424 (N_15424,N_14792,N_14692);
nand U15425 (N_15425,N_14503,N_14551);
xnor U15426 (N_15426,N_14725,N_14861);
or U15427 (N_15427,N_14737,N_14505);
and U15428 (N_15428,N_14997,N_14842);
and U15429 (N_15429,N_14863,N_14926);
nor U15430 (N_15430,N_14720,N_14619);
xor U15431 (N_15431,N_14648,N_14650);
nand U15432 (N_15432,N_14907,N_14599);
or U15433 (N_15433,N_14663,N_14853);
nand U15434 (N_15434,N_14527,N_14757);
or U15435 (N_15435,N_14868,N_14967);
nand U15436 (N_15436,N_14828,N_14537);
xor U15437 (N_15437,N_14751,N_14730);
nand U15438 (N_15438,N_14911,N_14538);
nand U15439 (N_15439,N_14606,N_14715);
nor U15440 (N_15440,N_14513,N_14573);
or U15441 (N_15441,N_14578,N_14656);
nand U15442 (N_15442,N_14651,N_14582);
xnor U15443 (N_15443,N_14701,N_14874);
nand U15444 (N_15444,N_14984,N_14590);
nand U15445 (N_15445,N_14851,N_14983);
xnor U15446 (N_15446,N_14593,N_14511);
nor U15447 (N_15447,N_14666,N_14902);
xnor U15448 (N_15448,N_14954,N_14912);
and U15449 (N_15449,N_14616,N_14873);
nand U15450 (N_15450,N_14589,N_14510);
xor U15451 (N_15451,N_14990,N_14602);
and U15452 (N_15452,N_14896,N_14998);
or U15453 (N_15453,N_14560,N_14687);
nor U15454 (N_15454,N_14996,N_14633);
xnor U15455 (N_15455,N_14705,N_14785);
and U15456 (N_15456,N_14692,N_14674);
or U15457 (N_15457,N_14951,N_14568);
and U15458 (N_15458,N_14737,N_14989);
nor U15459 (N_15459,N_14558,N_14996);
or U15460 (N_15460,N_14690,N_14959);
nand U15461 (N_15461,N_14743,N_14536);
nor U15462 (N_15462,N_14971,N_14994);
or U15463 (N_15463,N_14919,N_14745);
and U15464 (N_15464,N_14506,N_14772);
xnor U15465 (N_15465,N_14585,N_14633);
nor U15466 (N_15466,N_14878,N_14855);
xor U15467 (N_15467,N_14659,N_14948);
or U15468 (N_15468,N_14522,N_14661);
and U15469 (N_15469,N_14813,N_14603);
and U15470 (N_15470,N_14689,N_14674);
or U15471 (N_15471,N_14539,N_14508);
xor U15472 (N_15472,N_14532,N_14779);
and U15473 (N_15473,N_14545,N_14605);
or U15474 (N_15474,N_14836,N_14864);
nor U15475 (N_15475,N_14584,N_14614);
and U15476 (N_15476,N_14983,N_14911);
nor U15477 (N_15477,N_14979,N_14993);
nand U15478 (N_15478,N_14813,N_14614);
xnor U15479 (N_15479,N_14735,N_14801);
xnor U15480 (N_15480,N_14533,N_14529);
or U15481 (N_15481,N_14725,N_14665);
and U15482 (N_15482,N_14714,N_14778);
nor U15483 (N_15483,N_14880,N_14669);
and U15484 (N_15484,N_14602,N_14626);
and U15485 (N_15485,N_14684,N_14760);
nand U15486 (N_15486,N_14507,N_14662);
xor U15487 (N_15487,N_14983,N_14956);
or U15488 (N_15488,N_14680,N_14801);
and U15489 (N_15489,N_14801,N_14945);
nor U15490 (N_15490,N_14871,N_14777);
or U15491 (N_15491,N_14719,N_14522);
nand U15492 (N_15492,N_14874,N_14630);
nand U15493 (N_15493,N_14558,N_14576);
nor U15494 (N_15494,N_14510,N_14729);
xor U15495 (N_15495,N_14975,N_14636);
xor U15496 (N_15496,N_14536,N_14868);
xor U15497 (N_15497,N_14767,N_14897);
nand U15498 (N_15498,N_14716,N_14664);
and U15499 (N_15499,N_14520,N_14803);
nor U15500 (N_15500,N_15177,N_15014);
or U15501 (N_15501,N_15441,N_15237);
or U15502 (N_15502,N_15083,N_15216);
and U15503 (N_15503,N_15484,N_15469);
or U15504 (N_15504,N_15477,N_15282);
and U15505 (N_15505,N_15337,N_15463);
nor U15506 (N_15506,N_15331,N_15077);
xnor U15507 (N_15507,N_15189,N_15298);
nor U15508 (N_15508,N_15163,N_15111);
nor U15509 (N_15509,N_15359,N_15131);
nor U15510 (N_15510,N_15417,N_15062);
and U15511 (N_15511,N_15490,N_15200);
or U15512 (N_15512,N_15411,N_15385);
xnor U15513 (N_15513,N_15404,N_15425);
xnor U15514 (N_15514,N_15066,N_15136);
nand U15515 (N_15515,N_15160,N_15258);
nand U15516 (N_15516,N_15152,N_15130);
nor U15517 (N_15517,N_15384,N_15491);
nand U15518 (N_15518,N_15346,N_15156);
nor U15519 (N_15519,N_15195,N_15168);
or U15520 (N_15520,N_15045,N_15106);
nand U15521 (N_15521,N_15209,N_15080);
nor U15522 (N_15522,N_15095,N_15219);
or U15523 (N_15523,N_15462,N_15186);
xor U15524 (N_15524,N_15245,N_15496);
and U15525 (N_15525,N_15374,N_15357);
nor U15526 (N_15526,N_15064,N_15029);
or U15527 (N_15527,N_15344,N_15323);
and U15528 (N_15528,N_15220,N_15234);
xor U15529 (N_15529,N_15035,N_15386);
xnor U15530 (N_15530,N_15324,N_15471);
and U15531 (N_15531,N_15141,N_15101);
xor U15532 (N_15532,N_15159,N_15314);
nor U15533 (N_15533,N_15096,N_15086);
nand U15534 (N_15534,N_15443,N_15285);
nand U15535 (N_15535,N_15303,N_15199);
nand U15536 (N_15536,N_15482,N_15015);
nand U15537 (N_15537,N_15452,N_15218);
or U15538 (N_15538,N_15248,N_15224);
xnor U15539 (N_15539,N_15355,N_15495);
nor U15540 (N_15540,N_15435,N_15294);
xor U15541 (N_15541,N_15475,N_15065);
xnor U15542 (N_15542,N_15120,N_15124);
xnor U15543 (N_15543,N_15005,N_15138);
and U15544 (N_15544,N_15423,N_15320);
or U15545 (N_15545,N_15135,N_15094);
xor U15546 (N_15546,N_15287,N_15261);
or U15547 (N_15547,N_15307,N_15039);
nand U15548 (N_15548,N_15453,N_15302);
or U15549 (N_15549,N_15099,N_15273);
xor U15550 (N_15550,N_15157,N_15461);
nor U15551 (N_15551,N_15436,N_15191);
or U15552 (N_15552,N_15059,N_15254);
xnor U15553 (N_15553,N_15370,N_15037);
xor U15554 (N_15554,N_15052,N_15450);
nand U15555 (N_15555,N_15342,N_15444);
and U15556 (N_15556,N_15310,N_15176);
nor U15557 (N_15557,N_15119,N_15365);
nand U15558 (N_15558,N_15449,N_15033);
nor U15559 (N_15559,N_15115,N_15363);
xor U15560 (N_15560,N_15277,N_15356);
nand U15561 (N_15561,N_15414,N_15304);
nor U15562 (N_15562,N_15071,N_15420);
or U15563 (N_15563,N_15103,N_15421);
nand U15564 (N_15564,N_15088,N_15118);
or U15565 (N_15565,N_15143,N_15092);
nand U15566 (N_15566,N_15205,N_15084);
xor U15567 (N_15567,N_15116,N_15339);
nor U15568 (N_15568,N_15153,N_15253);
nor U15569 (N_15569,N_15008,N_15493);
nor U15570 (N_15570,N_15376,N_15334);
nor U15571 (N_15571,N_15410,N_15001);
and U15572 (N_15572,N_15260,N_15329);
xnor U15573 (N_15573,N_15022,N_15380);
and U15574 (N_15574,N_15227,N_15291);
or U15575 (N_15575,N_15048,N_15241);
and U15576 (N_15576,N_15247,N_15046);
and U15577 (N_15577,N_15286,N_15161);
nor U15578 (N_15578,N_15348,N_15290);
xnor U15579 (N_15579,N_15485,N_15117);
nand U15580 (N_15580,N_15128,N_15321);
or U15581 (N_15581,N_15221,N_15389);
or U15582 (N_15582,N_15377,N_15139);
and U15583 (N_15583,N_15054,N_15497);
nand U15584 (N_15584,N_15439,N_15003);
or U15585 (N_15585,N_15250,N_15432);
and U15586 (N_15586,N_15038,N_15297);
or U15587 (N_15587,N_15229,N_15358);
nand U15588 (N_15588,N_15460,N_15366);
and U15589 (N_15589,N_15479,N_15004);
and U15590 (N_15590,N_15378,N_15036);
or U15591 (N_15591,N_15170,N_15072);
nor U15592 (N_15592,N_15238,N_15413);
nor U15593 (N_15593,N_15150,N_15397);
or U15594 (N_15594,N_15327,N_15295);
and U15595 (N_15595,N_15492,N_15308);
and U15596 (N_15596,N_15387,N_15447);
and U15597 (N_15597,N_15299,N_15053);
nand U15598 (N_15598,N_15213,N_15264);
and U15599 (N_15599,N_15401,N_15203);
xor U15600 (N_15600,N_15049,N_15412);
or U15601 (N_15601,N_15296,N_15486);
and U15602 (N_15602,N_15201,N_15174);
or U15603 (N_15603,N_15341,N_15407);
xnor U15604 (N_15604,N_15433,N_15399);
nor U15605 (N_15605,N_15400,N_15373);
nor U15606 (N_15606,N_15305,N_15097);
nor U15607 (N_15607,N_15069,N_15431);
nor U15608 (N_15608,N_15325,N_15142);
or U15609 (N_15609,N_15448,N_15240);
nor U15610 (N_15610,N_15102,N_15498);
xor U15611 (N_15611,N_15235,N_15051);
nand U15612 (N_15612,N_15178,N_15123);
xnor U15613 (N_15613,N_15180,N_15204);
nand U15614 (N_15614,N_15211,N_15067);
nor U15615 (N_15615,N_15457,N_15364);
or U15616 (N_15616,N_15353,N_15246);
nand U15617 (N_15617,N_15473,N_15270);
nor U15618 (N_15618,N_15074,N_15017);
and U15619 (N_15619,N_15061,N_15114);
or U15620 (N_15620,N_15214,N_15289);
nor U15621 (N_15621,N_15464,N_15073);
xor U15622 (N_15622,N_15175,N_15019);
and U15623 (N_15623,N_15121,N_15406);
or U15624 (N_15624,N_15025,N_15352);
nand U15625 (N_15625,N_15179,N_15230);
xnor U15626 (N_15626,N_15255,N_15391);
nand U15627 (N_15627,N_15058,N_15474);
nand U15628 (N_15628,N_15481,N_15082);
nor U15629 (N_15629,N_15089,N_15202);
and U15630 (N_15630,N_15030,N_15335);
and U15631 (N_15631,N_15232,N_15372);
and U15632 (N_15632,N_15332,N_15351);
nor U15633 (N_15633,N_15454,N_15426);
nor U15634 (N_15634,N_15016,N_15422);
or U15635 (N_15635,N_15430,N_15415);
and U15636 (N_15636,N_15060,N_15317);
nor U15637 (N_15637,N_15489,N_15483);
nand U15638 (N_15638,N_15184,N_15110);
and U15639 (N_15639,N_15000,N_15040);
or U15640 (N_15640,N_15133,N_15242);
xnor U15641 (N_15641,N_15311,N_15438);
and U15642 (N_15642,N_15210,N_15243);
or U15643 (N_15643,N_15233,N_15193);
and U15644 (N_15644,N_15023,N_15068);
nand U15645 (N_15645,N_15026,N_15126);
nand U15646 (N_15646,N_15113,N_15013);
and U15647 (N_15647,N_15402,N_15322);
nor U15648 (N_15648,N_15267,N_15275);
nand U15649 (N_15649,N_15395,N_15252);
and U15650 (N_15650,N_15091,N_15472);
or U15651 (N_15651,N_15125,N_15345);
nand U15652 (N_15652,N_15338,N_15343);
or U15653 (N_15653,N_15288,N_15476);
or U15654 (N_15654,N_15181,N_15336);
xor U15655 (N_15655,N_15171,N_15166);
nor U15656 (N_15656,N_15134,N_15182);
nor U15657 (N_15657,N_15313,N_15408);
nor U15658 (N_15658,N_15458,N_15187);
xor U15659 (N_15659,N_15041,N_15132);
nand U15660 (N_15660,N_15367,N_15268);
and U15661 (N_15661,N_15434,N_15006);
and U15662 (N_15662,N_15440,N_15027);
nor U15663 (N_15663,N_15362,N_15212);
and U15664 (N_15664,N_15207,N_15369);
or U15665 (N_15665,N_15354,N_15251);
and U15666 (N_15666,N_15011,N_15108);
or U15667 (N_15667,N_15271,N_15292);
and U15668 (N_15668,N_15446,N_15480);
or U15669 (N_15669,N_15018,N_15122);
and U15670 (N_15670,N_15276,N_15371);
nand U15671 (N_15671,N_15257,N_15478);
and U15672 (N_15672,N_15231,N_15009);
xor U15673 (N_15673,N_15007,N_15109);
nor U15674 (N_15674,N_15236,N_15405);
nor U15675 (N_15675,N_15306,N_15206);
nor U15676 (N_15676,N_15167,N_15470);
nor U15677 (N_15677,N_15265,N_15024);
or U15678 (N_15678,N_15381,N_15070);
nand U15679 (N_15679,N_15244,N_15012);
xnor U15680 (N_15680,N_15451,N_15032);
or U15681 (N_15681,N_15188,N_15183);
xor U15682 (N_15682,N_15031,N_15063);
nand U15683 (N_15683,N_15239,N_15468);
or U15684 (N_15684,N_15044,N_15280);
xor U15685 (N_15685,N_15190,N_15021);
xnor U15686 (N_15686,N_15416,N_15100);
nand U15687 (N_15687,N_15326,N_15262);
xor U15688 (N_15688,N_15087,N_15390);
xnor U15689 (N_15689,N_15284,N_15034);
nand U15690 (N_15690,N_15269,N_15328);
nor U15691 (N_15691,N_15226,N_15196);
nand U15692 (N_15692,N_15169,N_15301);
and U15693 (N_15693,N_15043,N_15340);
and U15694 (N_15694,N_15300,N_15050);
or U15695 (N_15695,N_15140,N_15392);
nand U15696 (N_15696,N_15466,N_15020);
and U15697 (N_15697,N_15456,N_15076);
and U15698 (N_15698,N_15488,N_15467);
nand U15699 (N_15699,N_15098,N_15194);
and U15700 (N_15700,N_15349,N_15429);
nor U15701 (N_15701,N_15278,N_15281);
xor U15702 (N_15702,N_15079,N_15465);
nand U15703 (N_15703,N_15147,N_15081);
nor U15704 (N_15704,N_15158,N_15360);
nand U15705 (N_15705,N_15375,N_15185);
nor U15706 (N_15706,N_15361,N_15418);
nand U15707 (N_15707,N_15263,N_15309);
and U15708 (N_15708,N_15225,N_15208);
nand U15709 (N_15709,N_15112,N_15090);
and U15710 (N_15710,N_15148,N_15445);
nor U15711 (N_15711,N_15085,N_15127);
xnor U15712 (N_15712,N_15383,N_15437);
and U15713 (N_15713,N_15316,N_15192);
and U15714 (N_15714,N_15154,N_15010);
or U15715 (N_15715,N_15427,N_15293);
xor U15716 (N_15716,N_15151,N_15279);
nor U15717 (N_15717,N_15144,N_15283);
nor U15718 (N_15718,N_15428,N_15137);
nand U15719 (N_15719,N_15274,N_15162);
xor U15720 (N_15720,N_15368,N_15499);
nand U15721 (N_15721,N_15197,N_15105);
nand U15722 (N_15722,N_15057,N_15419);
nand U15723 (N_15723,N_15173,N_15104);
nor U15724 (N_15724,N_15398,N_15042);
and U15725 (N_15725,N_15442,N_15459);
or U15726 (N_15726,N_15047,N_15455);
or U15727 (N_15727,N_15223,N_15028);
nand U15728 (N_15728,N_15347,N_15107);
nand U15729 (N_15729,N_15494,N_15319);
nand U15730 (N_15730,N_15318,N_15312);
or U15731 (N_15731,N_15215,N_15409);
nand U15732 (N_15732,N_15396,N_15382);
xor U15733 (N_15733,N_15002,N_15403);
nor U15734 (N_15734,N_15330,N_15272);
and U15735 (N_15735,N_15350,N_15388);
nor U15736 (N_15736,N_15146,N_15315);
nand U15737 (N_15737,N_15145,N_15393);
nor U15738 (N_15738,N_15228,N_15198);
xor U15739 (N_15739,N_15222,N_15379);
nand U15740 (N_15740,N_15172,N_15075);
and U15741 (N_15741,N_15394,N_15249);
and U15742 (N_15742,N_15259,N_15256);
nor U15743 (N_15743,N_15078,N_15055);
nand U15744 (N_15744,N_15333,N_15056);
or U15745 (N_15745,N_15424,N_15266);
nor U15746 (N_15746,N_15093,N_15155);
nor U15747 (N_15747,N_15217,N_15149);
xnor U15748 (N_15748,N_15165,N_15164);
nand U15749 (N_15749,N_15487,N_15129);
nand U15750 (N_15750,N_15022,N_15148);
or U15751 (N_15751,N_15247,N_15018);
or U15752 (N_15752,N_15432,N_15219);
nor U15753 (N_15753,N_15399,N_15347);
xnor U15754 (N_15754,N_15003,N_15410);
or U15755 (N_15755,N_15341,N_15165);
nand U15756 (N_15756,N_15295,N_15367);
or U15757 (N_15757,N_15091,N_15408);
nor U15758 (N_15758,N_15157,N_15444);
or U15759 (N_15759,N_15100,N_15087);
or U15760 (N_15760,N_15208,N_15150);
nand U15761 (N_15761,N_15181,N_15409);
and U15762 (N_15762,N_15401,N_15207);
nand U15763 (N_15763,N_15039,N_15262);
xor U15764 (N_15764,N_15348,N_15306);
or U15765 (N_15765,N_15008,N_15298);
and U15766 (N_15766,N_15495,N_15463);
xor U15767 (N_15767,N_15162,N_15273);
and U15768 (N_15768,N_15034,N_15347);
or U15769 (N_15769,N_15095,N_15268);
nor U15770 (N_15770,N_15471,N_15101);
nor U15771 (N_15771,N_15375,N_15346);
nor U15772 (N_15772,N_15198,N_15442);
nand U15773 (N_15773,N_15480,N_15139);
nor U15774 (N_15774,N_15411,N_15233);
xnor U15775 (N_15775,N_15104,N_15330);
or U15776 (N_15776,N_15082,N_15085);
or U15777 (N_15777,N_15096,N_15026);
xor U15778 (N_15778,N_15437,N_15029);
nand U15779 (N_15779,N_15013,N_15158);
or U15780 (N_15780,N_15171,N_15043);
nand U15781 (N_15781,N_15127,N_15170);
or U15782 (N_15782,N_15312,N_15334);
xnor U15783 (N_15783,N_15082,N_15420);
or U15784 (N_15784,N_15217,N_15260);
xnor U15785 (N_15785,N_15405,N_15094);
nor U15786 (N_15786,N_15201,N_15418);
or U15787 (N_15787,N_15474,N_15317);
nor U15788 (N_15788,N_15024,N_15288);
and U15789 (N_15789,N_15005,N_15022);
or U15790 (N_15790,N_15461,N_15388);
or U15791 (N_15791,N_15010,N_15485);
xnor U15792 (N_15792,N_15430,N_15141);
nor U15793 (N_15793,N_15033,N_15067);
nor U15794 (N_15794,N_15244,N_15475);
or U15795 (N_15795,N_15032,N_15008);
and U15796 (N_15796,N_15319,N_15315);
nand U15797 (N_15797,N_15292,N_15041);
and U15798 (N_15798,N_15172,N_15066);
nand U15799 (N_15799,N_15384,N_15468);
or U15800 (N_15800,N_15012,N_15019);
xnor U15801 (N_15801,N_15204,N_15189);
nand U15802 (N_15802,N_15190,N_15460);
xnor U15803 (N_15803,N_15456,N_15101);
nand U15804 (N_15804,N_15085,N_15462);
and U15805 (N_15805,N_15250,N_15247);
nand U15806 (N_15806,N_15156,N_15431);
xor U15807 (N_15807,N_15466,N_15468);
or U15808 (N_15808,N_15203,N_15177);
and U15809 (N_15809,N_15321,N_15242);
and U15810 (N_15810,N_15073,N_15091);
and U15811 (N_15811,N_15300,N_15052);
or U15812 (N_15812,N_15138,N_15007);
or U15813 (N_15813,N_15391,N_15201);
and U15814 (N_15814,N_15331,N_15123);
nand U15815 (N_15815,N_15116,N_15346);
and U15816 (N_15816,N_15419,N_15472);
xnor U15817 (N_15817,N_15279,N_15109);
or U15818 (N_15818,N_15313,N_15118);
xnor U15819 (N_15819,N_15096,N_15376);
xnor U15820 (N_15820,N_15276,N_15060);
or U15821 (N_15821,N_15251,N_15107);
and U15822 (N_15822,N_15376,N_15358);
and U15823 (N_15823,N_15045,N_15406);
xor U15824 (N_15824,N_15179,N_15245);
and U15825 (N_15825,N_15261,N_15395);
or U15826 (N_15826,N_15080,N_15272);
or U15827 (N_15827,N_15439,N_15456);
nor U15828 (N_15828,N_15053,N_15280);
or U15829 (N_15829,N_15118,N_15190);
nor U15830 (N_15830,N_15372,N_15200);
and U15831 (N_15831,N_15075,N_15380);
and U15832 (N_15832,N_15488,N_15339);
nor U15833 (N_15833,N_15232,N_15150);
nor U15834 (N_15834,N_15182,N_15421);
nor U15835 (N_15835,N_15099,N_15032);
or U15836 (N_15836,N_15157,N_15246);
nor U15837 (N_15837,N_15234,N_15080);
and U15838 (N_15838,N_15391,N_15316);
nand U15839 (N_15839,N_15409,N_15427);
nor U15840 (N_15840,N_15114,N_15356);
xnor U15841 (N_15841,N_15102,N_15195);
xor U15842 (N_15842,N_15173,N_15310);
nand U15843 (N_15843,N_15150,N_15406);
xor U15844 (N_15844,N_15396,N_15322);
or U15845 (N_15845,N_15416,N_15370);
xnor U15846 (N_15846,N_15382,N_15347);
nand U15847 (N_15847,N_15276,N_15301);
nand U15848 (N_15848,N_15152,N_15413);
nor U15849 (N_15849,N_15024,N_15204);
xnor U15850 (N_15850,N_15083,N_15342);
and U15851 (N_15851,N_15316,N_15134);
or U15852 (N_15852,N_15467,N_15081);
nand U15853 (N_15853,N_15222,N_15489);
and U15854 (N_15854,N_15286,N_15073);
nor U15855 (N_15855,N_15470,N_15035);
or U15856 (N_15856,N_15043,N_15001);
or U15857 (N_15857,N_15001,N_15096);
xnor U15858 (N_15858,N_15190,N_15255);
nand U15859 (N_15859,N_15052,N_15202);
or U15860 (N_15860,N_15166,N_15259);
nor U15861 (N_15861,N_15497,N_15485);
and U15862 (N_15862,N_15484,N_15231);
and U15863 (N_15863,N_15241,N_15023);
or U15864 (N_15864,N_15144,N_15376);
or U15865 (N_15865,N_15277,N_15249);
and U15866 (N_15866,N_15017,N_15317);
xnor U15867 (N_15867,N_15143,N_15275);
nor U15868 (N_15868,N_15236,N_15354);
nand U15869 (N_15869,N_15172,N_15092);
nand U15870 (N_15870,N_15095,N_15238);
nand U15871 (N_15871,N_15206,N_15133);
xor U15872 (N_15872,N_15209,N_15439);
xnor U15873 (N_15873,N_15252,N_15172);
nand U15874 (N_15874,N_15208,N_15157);
and U15875 (N_15875,N_15070,N_15373);
nor U15876 (N_15876,N_15079,N_15366);
nand U15877 (N_15877,N_15330,N_15321);
or U15878 (N_15878,N_15058,N_15046);
nand U15879 (N_15879,N_15357,N_15255);
xnor U15880 (N_15880,N_15374,N_15170);
or U15881 (N_15881,N_15268,N_15136);
nor U15882 (N_15882,N_15133,N_15450);
nand U15883 (N_15883,N_15067,N_15408);
nand U15884 (N_15884,N_15147,N_15095);
xor U15885 (N_15885,N_15087,N_15080);
xor U15886 (N_15886,N_15135,N_15319);
or U15887 (N_15887,N_15119,N_15082);
nor U15888 (N_15888,N_15037,N_15155);
nand U15889 (N_15889,N_15003,N_15462);
xor U15890 (N_15890,N_15163,N_15337);
nand U15891 (N_15891,N_15090,N_15468);
and U15892 (N_15892,N_15161,N_15282);
and U15893 (N_15893,N_15014,N_15299);
nand U15894 (N_15894,N_15030,N_15139);
nor U15895 (N_15895,N_15437,N_15059);
or U15896 (N_15896,N_15399,N_15045);
xnor U15897 (N_15897,N_15449,N_15372);
or U15898 (N_15898,N_15046,N_15073);
nand U15899 (N_15899,N_15467,N_15245);
nand U15900 (N_15900,N_15263,N_15120);
nor U15901 (N_15901,N_15013,N_15128);
and U15902 (N_15902,N_15390,N_15315);
and U15903 (N_15903,N_15109,N_15198);
and U15904 (N_15904,N_15421,N_15146);
or U15905 (N_15905,N_15185,N_15386);
xnor U15906 (N_15906,N_15393,N_15367);
nor U15907 (N_15907,N_15354,N_15279);
nor U15908 (N_15908,N_15443,N_15322);
nor U15909 (N_15909,N_15195,N_15281);
or U15910 (N_15910,N_15165,N_15337);
nor U15911 (N_15911,N_15050,N_15469);
and U15912 (N_15912,N_15339,N_15348);
nor U15913 (N_15913,N_15116,N_15034);
nor U15914 (N_15914,N_15464,N_15345);
nor U15915 (N_15915,N_15206,N_15100);
xnor U15916 (N_15916,N_15416,N_15192);
or U15917 (N_15917,N_15432,N_15136);
and U15918 (N_15918,N_15108,N_15442);
xnor U15919 (N_15919,N_15427,N_15189);
xor U15920 (N_15920,N_15479,N_15014);
and U15921 (N_15921,N_15096,N_15127);
nor U15922 (N_15922,N_15194,N_15483);
nand U15923 (N_15923,N_15498,N_15424);
nand U15924 (N_15924,N_15241,N_15081);
or U15925 (N_15925,N_15174,N_15145);
and U15926 (N_15926,N_15228,N_15021);
or U15927 (N_15927,N_15484,N_15265);
nand U15928 (N_15928,N_15272,N_15122);
or U15929 (N_15929,N_15376,N_15351);
or U15930 (N_15930,N_15385,N_15483);
xor U15931 (N_15931,N_15433,N_15042);
and U15932 (N_15932,N_15255,N_15250);
nor U15933 (N_15933,N_15121,N_15485);
xor U15934 (N_15934,N_15077,N_15143);
and U15935 (N_15935,N_15032,N_15125);
and U15936 (N_15936,N_15296,N_15401);
or U15937 (N_15937,N_15248,N_15366);
nor U15938 (N_15938,N_15427,N_15239);
nor U15939 (N_15939,N_15333,N_15109);
nor U15940 (N_15940,N_15282,N_15370);
or U15941 (N_15941,N_15075,N_15308);
and U15942 (N_15942,N_15268,N_15294);
or U15943 (N_15943,N_15371,N_15177);
xnor U15944 (N_15944,N_15062,N_15098);
and U15945 (N_15945,N_15090,N_15154);
and U15946 (N_15946,N_15300,N_15372);
xnor U15947 (N_15947,N_15078,N_15218);
and U15948 (N_15948,N_15466,N_15158);
xnor U15949 (N_15949,N_15145,N_15182);
or U15950 (N_15950,N_15413,N_15411);
and U15951 (N_15951,N_15098,N_15433);
nand U15952 (N_15952,N_15390,N_15305);
nand U15953 (N_15953,N_15396,N_15076);
nand U15954 (N_15954,N_15060,N_15412);
nand U15955 (N_15955,N_15460,N_15417);
xnor U15956 (N_15956,N_15484,N_15499);
xor U15957 (N_15957,N_15035,N_15409);
nor U15958 (N_15958,N_15327,N_15358);
nor U15959 (N_15959,N_15205,N_15282);
and U15960 (N_15960,N_15411,N_15357);
xor U15961 (N_15961,N_15037,N_15492);
nand U15962 (N_15962,N_15229,N_15036);
xnor U15963 (N_15963,N_15314,N_15373);
and U15964 (N_15964,N_15020,N_15063);
nand U15965 (N_15965,N_15046,N_15308);
nand U15966 (N_15966,N_15275,N_15146);
or U15967 (N_15967,N_15345,N_15170);
or U15968 (N_15968,N_15068,N_15416);
and U15969 (N_15969,N_15354,N_15162);
and U15970 (N_15970,N_15374,N_15299);
or U15971 (N_15971,N_15304,N_15244);
and U15972 (N_15972,N_15469,N_15452);
or U15973 (N_15973,N_15345,N_15457);
and U15974 (N_15974,N_15355,N_15493);
nor U15975 (N_15975,N_15463,N_15191);
nor U15976 (N_15976,N_15204,N_15241);
or U15977 (N_15977,N_15455,N_15273);
xor U15978 (N_15978,N_15285,N_15137);
xor U15979 (N_15979,N_15388,N_15028);
nand U15980 (N_15980,N_15052,N_15064);
nand U15981 (N_15981,N_15051,N_15310);
or U15982 (N_15982,N_15220,N_15061);
and U15983 (N_15983,N_15013,N_15306);
xor U15984 (N_15984,N_15223,N_15116);
nor U15985 (N_15985,N_15409,N_15317);
or U15986 (N_15986,N_15137,N_15205);
and U15987 (N_15987,N_15101,N_15213);
or U15988 (N_15988,N_15254,N_15488);
xor U15989 (N_15989,N_15250,N_15467);
and U15990 (N_15990,N_15491,N_15016);
or U15991 (N_15991,N_15118,N_15155);
nor U15992 (N_15992,N_15052,N_15289);
nor U15993 (N_15993,N_15296,N_15069);
or U15994 (N_15994,N_15122,N_15248);
and U15995 (N_15995,N_15256,N_15455);
nand U15996 (N_15996,N_15155,N_15302);
xor U15997 (N_15997,N_15184,N_15168);
nor U15998 (N_15998,N_15480,N_15070);
nor U15999 (N_15999,N_15132,N_15255);
nor U16000 (N_16000,N_15511,N_15903);
or U16001 (N_16001,N_15921,N_15916);
or U16002 (N_16002,N_15934,N_15678);
xnor U16003 (N_16003,N_15800,N_15614);
nor U16004 (N_16004,N_15835,N_15600);
and U16005 (N_16005,N_15851,N_15913);
or U16006 (N_16006,N_15679,N_15905);
nor U16007 (N_16007,N_15624,N_15620);
and U16008 (N_16008,N_15636,N_15820);
nor U16009 (N_16009,N_15541,N_15500);
nor U16010 (N_16010,N_15822,N_15946);
nor U16011 (N_16011,N_15900,N_15713);
or U16012 (N_16012,N_15551,N_15648);
xor U16013 (N_16013,N_15881,N_15766);
and U16014 (N_16014,N_15911,N_15988);
nor U16015 (N_16015,N_15544,N_15659);
nor U16016 (N_16016,N_15663,N_15944);
and U16017 (N_16017,N_15828,N_15676);
or U16018 (N_16018,N_15969,N_15780);
xor U16019 (N_16019,N_15645,N_15744);
nand U16020 (N_16020,N_15644,N_15816);
and U16021 (N_16021,N_15973,N_15897);
or U16022 (N_16022,N_15700,N_15737);
and U16023 (N_16023,N_15601,N_15703);
nand U16024 (N_16024,N_15824,N_15777);
or U16025 (N_16025,N_15653,N_15637);
nor U16026 (N_16026,N_15596,N_15697);
nor U16027 (N_16027,N_15962,N_15891);
and U16028 (N_16028,N_15517,N_15751);
nor U16029 (N_16029,N_15638,N_15559);
xor U16030 (N_16030,N_15603,N_15955);
xnor U16031 (N_16031,N_15981,N_15927);
and U16032 (N_16032,N_15890,N_15506);
nand U16033 (N_16033,N_15712,N_15733);
nor U16034 (N_16034,N_15692,N_15536);
nand U16035 (N_16035,N_15887,N_15761);
and U16036 (N_16036,N_15862,N_15707);
nor U16037 (N_16037,N_15910,N_15831);
or U16038 (N_16038,N_15554,N_15612);
or U16039 (N_16039,N_15677,N_15635);
nor U16040 (N_16040,N_15959,N_15529);
or U16041 (N_16041,N_15542,N_15995);
nor U16042 (N_16042,N_15634,N_15804);
nand U16043 (N_16043,N_15985,N_15740);
and U16044 (N_16044,N_15513,N_15920);
nor U16045 (N_16045,N_15523,N_15772);
nor U16046 (N_16046,N_15923,N_15791);
nor U16047 (N_16047,N_15509,N_15912);
nand U16048 (N_16048,N_15618,N_15527);
xnor U16049 (N_16049,N_15884,N_15814);
or U16050 (N_16050,N_15746,N_15615);
xor U16051 (N_16051,N_15844,N_15811);
and U16052 (N_16052,N_15882,N_15664);
nand U16053 (N_16053,N_15798,N_15970);
nand U16054 (N_16054,N_15555,N_15901);
or U16055 (N_16055,N_15584,N_15602);
nor U16056 (N_16056,N_15854,N_15594);
nand U16057 (N_16057,N_15963,N_15670);
and U16058 (N_16058,N_15764,N_15702);
or U16059 (N_16059,N_15731,N_15688);
nor U16060 (N_16060,N_15585,N_15694);
or U16061 (N_16061,N_15753,N_15704);
nand U16062 (N_16062,N_15756,N_15986);
nor U16063 (N_16063,N_15619,N_15657);
xnor U16064 (N_16064,N_15793,N_15718);
nand U16065 (N_16065,N_15558,N_15721);
nand U16066 (N_16066,N_15609,N_15629);
or U16067 (N_16067,N_15691,N_15507);
nor U16068 (N_16068,N_15987,N_15743);
and U16069 (N_16069,N_15829,N_15656);
and U16070 (N_16070,N_15690,N_15747);
or U16071 (N_16071,N_15840,N_15550);
xor U16072 (N_16072,N_15931,N_15752);
nor U16073 (N_16073,N_15611,N_15906);
or U16074 (N_16074,N_15525,N_15658);
and U16075 (N_16075,N_15505,N_15871);
nor U16076 (N_16076,N_15849,N_15661);
nand U16077 (N_16077,N_15982,N_15592);
xnor U16078 (N_16078,N_15873,N_15984);
or U16079 (N_16079,N_15874,N_15787);
and U16080 (N_16080,N_15514,N_15760);
nor U16081 (N_16081,N_15683,N_15860);
xnor U16082 (N_16082,N_15604,N_15672);
nand U16083 (N_16083,N_15586,N_15528);
or U16084 (N_16084,N_15671,N_15735);
and U16085 (N_16085,N_15714,N_15922);
or U16086 (N_16086,N_15641,N_15813);
or U16087 (N_16087,N_15686,N_15533);
xnor U16088 (N_16088,N_15781,N_15974);
xnor U16089 (N_16089,N_15966,N_15834);
or U16090 (N_16090,N_15655,N_15877);
and U16091 (N_16091,N_15545,N_15680);
or U16092 (N_16092,N_15958,N_15940);
nand U16093 (N_16093,N_15622,N_15745);
and U16094 (N_16094,N_15832,N_15732);
nand U16095 (N_16095,N_15979,N_15626);
nor U16096 (N_16096,N_15767,N_15783);
or U16097 (N_16097,N_15510,N_15786);
and U16098 (N_16098,N_15796,N_15976);
nand U16099 (N_16099,N_15765,N_15968);
and U16100 (N_16100,N_15728,N_15886);
or U16101 (N_16101,N_15843,N_15599);
nand U16102 (N_16102,N_15883,N_15810);
nand U16103 (N_16103,N_15625,N_15817);
or U16104 (N_16104,N_15908,N_15865);
or U16105 (N_16105,N_15924,N_15939);
nor U16106 (N_16106,N_15956,N_15583);
and U16107 (N_16107,N_15830,N_15571);
xnor U16108 (N_16108,N_15972,N_15711);
nand U16109 (N_16109,N_15848,N_15633);
and U16110 (N_16110,N_15964,N_15701);
nand U16111 (N_16111,N_15763,N_15898);
nand U16112 (N_16112,N_15647,N_15685);
and U16113 (N_16113,N_15806,N_15738);
or U16114 (N_16114,N_15917,N_15557);
or U16115 (N_16115,N_15994,N_15943);
or U16116 (N_16116,N_15674,N_15868);
or U16117 (N_16117,N_15942,N_15705);
nand U16118 (N_16118,N_15710,N_15642);
and U16119 (N_16119,N_15520,N_15784);
xnor U16120 (N_16120,N_15965,N_15621);
nor U16121 (N_16121,N_15856,N_15792);
xnor U16122 (N_16122,N_15858,N_15899);
and U16123 (N_16123,N_15548,N_15823);
xnor U16124 (N_16124,N_15613,N_15902);
nand U16125 (N_16125,N_15805,N_15947);
and U16126 (N_16126,N_15651,N_15715);
nand U16127 (N_16127,N_15773,N_15932);
nor U16128 (N_16128,N_15825,N_15503);
nor U16129 (N_16129,N_15538,N_15930);
nand U16130 (N_16130,N_15859,N_15826);
and U16131 (N_16131,N_15867,N_15579);
xor U16132 (N_16132,N_15549,N_15998);
nand U16133 (N_16133,N_15543,N_15996);
nand U16134 (N_16134,N_15853,N_15526);
or U16135 (N_16135,N_15606,N_15821);
xnor U16136 (N_16136,N_15808,N_15778);
nor U16137 (N_16137,N_15807,N_15667);
xor U16138 (N_16138,N_15630,N_15669);
nor U16139 (N_16139,N_15833,N_15954);
and U16140 (N_16140,N_15650,N_15597);
and U16141 (N_16141,N_15782,N_15696);
xor U16142 (N_16142,N_15546,N_15501);
xnor U16143 (N_16143,N_15504,N_15730);
or U16144 (N_16144,N_15951,N_15852);
and U16145 (N_16145,N_15582,N_15904);
or U16146 (N_16146,N_15580,N_15578);
and U16147 (N_16147,N_15990,N_15864);
nor U16148 (N_16148,N_15631,N_15770);
and U16149 (N_16149,N_15693,N_15553);
or U16150 (N_16150,N_15723,N_15960);
and U16151 (N_16151,N_15741,N_15566);
xnor U16152 (N_16152,N_15768,N_15572);
and U16153 (N_16153,N_15872,N_15515);
xnor U16154 (N_16154,N_15983,N_15587);
or U16155 (N_16155,N_15878,N_15521);
xor U16156 (N_16156,N_15660,N_15518);
nand U16157 (N_16157,N_15623,N_15819);
nand U16158 (N_16158,N_15950,N_15531);
xor U16159 (N_16159,N_15563,N_15775);
nor U16160 (N_16160,N_15547,N_15845);
or U16161 (N_16161,N_15590,N_15598);
and U16162 (N_16162,N_15552,N_15725);
or U16163 (N_16163,N_15861,N_15855);
nor U16164 (N_16164,N_15759,N_15846);
xnor U16165 (N_16165,N_15789,N_15573);
nor U16166 (N_16166,N_15564,N_15698);
nor U16167 (N_16167,N_15895,N_15726);
or U16168 (N_16168,N_15668,N_15708);
xor U16169 (N_16169,N_15742,N_15896);
nand U16170 (N_16170,N_15560,N_15790);
nor U16171 (N_16171,N_15556,N_15941);
and U16172 (N_16172,N_15575,N_15681);
xor U16173 (N_16173,N_15616,N_15999);
nand U16174 (N_16174,N_15617,N_15762);
nand U16175 (N_16175,N_15729,N_15802);
nand U16176 (N_16176,N_15610,N_15978);
and U16177 (N_16177,N_15794,N_15971);
xnor U16178 (N_16178,N_15757,N_15919);
xor U16179 (N_16179,N_15516,N_15842);
xor U16180 (N_16180,N_15839,N_15928);
and U16181 (N_16181,N_15608,N_15640);
or U16182 (N_16182,N_15841,N_15749);
nor U16183 (N_16183,N_15926,N_15524);
and U16184 (N_16184,N_15706,N_15837);
nor U16185 (N_16185,N_15776,N_15565);
or U16186 (N_16186,N_15540,N_15534);
nor U16187 (N_16187,N_15665,N_15720);
and U16188 (N_16188,N_15695,N_15576);
xnor U16189 (N_16189,N_15888,N_15722);
and U16190 (N_16190,N_15997,N_15727);
nor U16191 (N_16191,N_15605,N_15577);
xor U16192 (N_16192,N_15748,N_15980);
or U16193 (N_16193,N_15799,N_15628);
nor U16194 (N_16194,N_15673,N_15535);
nor U16195 (N_16195,N_15893,N_15532);
nor U16196 (N_16196,N_15863,N_15795);
or U16197 (N_16197,N_15581,N_15769);
and U16198 (N_16198,N_15975,N_15836);
or U16199 (N_16199,N_15632,N_15682);
xnor U16200 (N_16200,N_15591,N_15918);
or U16201 (N_16201,N_15639,N_15914);
nand U16202 (N_16202,N_15937,N_15774);
xnor U16203 (N_16203,N_15953,N_15909);
and U16204 (N_16204,N_15870,N_15539);
nor U16205 (N_16205,N_15522,N_15797);
nor U16206 (N_16206,N_15687,N_15929);
xnor U16207 (N_16207,N_15643,N_15689);
xnor U16208 (N_16208,N_15967,N_15562);
and U16209 (N_16209,N_15945,N_15717);
or U16210 (N_16210,N_15818,N_15991);
or U16211 (N_16211,N_15827,N_15627);
xor U16212 (N_16212,N_15815,N_15993);
nor U16213 (N_16213,N_15754,N_15935);
or U16214 (N_16214,N_15734,N_15662);
and U16215 (N_16215,N_15809,N_15838);
nand U16216 (N_16216,N_15699,N_15812);
or U16217 (N_16217,N_15880,N_15709);
nand U16218 (N_16218,N_15875,N_15936);
nand U16219 (N_16219,N_15654,N_15850);
nor U16220 (N_16220,N_15779,N_15652);
and U16221 (N_16221,N_15739,N_15588);
xor U16222 (N_16222,N_15607,N_15907);
nand U16223 (N_16223,N_15961,N_15892);
nor U16224 (N_16224,N_15561,N_15675);
and U16225 (N_16225,N_15957,N_15803);
and U16226 (N_16226,N_15889,N_15876);
xor U16227 (N_16227,N_15537,N_15570);
and U16228 (N_16228,N_15646,N_15530);
or U16229 (N_16229,N_15938,N_15866);
xor U16230 (N_16230,N_15574,N_15649);
or U16231 (N_16231,N_15847,N_15569);
and U16232 (N_16232,N_15894,N_15593);
xor U16233 (N_16233,N_15724,N_15589);
or U16234 (N_16234,N_15519,N_15885);
nor U16235 (N_16235,N_15952,N_15508);
nor U16236 (N_16236,N_15788,N_15568);
and U16237 (N_16237,N_15755,N_15977);
xnor U16238 (N_16238,N_15869,N_15925);
xnor U16239 (N_16239,N_15989,N_15801);
or U16240 (N_16240,N_15567,N_15915);
xnor U16241 (N_16241,N_15758,N_15992);
and U16242 (N_16242,N_15771,N_15785);
xor U16243 (N_16243,N_15736,N_15750);
or U16244 (N_16244,N_15716,N_15719);
or U16245 (N_16245,N_15684,N_15857);
xnor U16246 (N_16246,N_15502,N_15666);
or U16247 (N_16247,N_15933,N_15512);
nand U16248 (N_16248,N_15595,N_15949);
or U16249 (N_16249,N_15948,N_15879);
or U16250 (N_16250,N_15926,N_15958);
nand U16251 (N_16251,N_15916,N_15986);
nand U16252 (N_16252,N_15546,N_15548);
nor U16253 (N_16253,N_15670,N_15836);
and U16254 (N_16254,N_15979,N_15658);
or U16255 (N_16255,N_15888,N_15640);
xor U16256 (N_16256,N_15600,N_15846);
nor U16257 (N_16257,N_15721,N_15929);
nor U16258 (N_16258,N_15674,N_15783);
xor U16259 (N_16259,N_15832,N_15646);
and U16260 (N_16260,N_15795,N_15781);
and U16261 (N_16261,N_15959,N_15810);
xnor U16262 (N_16262,N_15628,N_15553);
nand U16263 (N_16263,N_15756,N_15793);
nor U16264 (N_16264,N_15993,N_15880);
nor U16265 (N_16265,N_15875,N_15909);
nand U16266 (N_16266,N_15999,N_15846);
xnor U16267 (N_16267,N_15504,N_15714);
and U16268 (N_16268,N_15812,N_15948);
xnor U16269 (N_16269,N_15740,N_15590);
nor U16270 (N_16270,N_15872,N_15669);
xnor U16271 (N_16271,N_15588,N_15551);
or U16272 (N_16272,N_15967,N_15570);
or U16273 (N_16273,N_15655,N_15592);
nand U16274 (N_16274,N_15929,N_15823);
nor U16275 (N_16275,N_15660,N_15763);
xnor U16276 (N_16276,N_15577,N_15908);
nor U16277 (N_16277,N_15901,N_15702);
nand U16278 (N_16278,N_15770,N_15873);
nand U16279 (N_16279,N_15785,N_15835);
or U16280 (N_16280,N_15795,N_15791);
or U16281 (N_16281,N_15702,N_15913);
nor U16282 (N_16282,N_15732,N_15512);
xnor U16283 (N_16283,N_15892,N_15934);
nand U16284 (N_16284,N_15709,N_15737);
or U16285 (N_16285,N_15797,N_15669);
or U16286 (N_16286,N_15942,N_15621);
nor U16287 (N_16287,N_15601,N_15575);
nand U16288 (N_16288,N_15675,N_15788);
xnor U16289 (N_16289,N_15862,N_15980);
or U16290 (N_16290,N_15881,N_15911);
and U16291 (N_16291,N_15602,N_15596);
nor U16292 (N_16292,N_15978,N_15526);
or U16293 (N_16293,N_15861,N_15943);
or U16294 (N_16294,N_15909,N_15726);
and U16295 (N_16295,N_15850,N_15798);
xnor U16296 (N_16296,N_15735,N_15557);
xor U16297 (N_16297,N_15875,N_15910);
xnor U16298 (N_16298,N_15521,N_15520);
nor U16299 (N_16299,N_15899,N_15748);
and U16300 (N_16300,N_15770,N_15502);
xnor U16301 (N_16301,N_15915,N_15947);
nand U16302 (N_16302,N_15648,N_15645);
nand U16303 (N_16303,N_15574,N_15648);
nand U16304 (N_16304,N_15577,N_15937);
and U16305 (N_16305,N_15836,N_15633);
nor U16306 (N_16306,N_15779,N_15841);
xnor U16307 (N_16307,N_15589,N_15939);
and U16308 (N_16308,N_15532,N_15686);
nand U16309 (N_16309,N_15576,N_15799);
nor U16310 (N_16310,N_15970,N_15816);
or U16311 (N_16311,N_15839,N_15863);
xnor U16312 (N_16312,N_15872,N_15512);
and U16313 (N_16313,N_15780,N_15836);
xnor U16314 (N_16314,N_15759,N_15942);
and U16315 (N_16315,N_15770,N_15938);
or U16316 (N_16316,N_15757,N_15548);
nand U16317 (N_16317,N_15675,N_15713);
nand U16318 (N_16318,N_15602,N_15744);
nor U16319 (N_16319,N_15792,N_15957);
xor U16320 (N_16320,N_15772,N_15702);
and U16321 (N_16321,N_15779,N_15972);
xor U16322 (N_16322,N_15821,N_15647);
nor U16323 (N_16323,N_15956,N_15747);
and U16324 (N_16324,N_15690,N_15639);
nand U16325 (N_16325,N_15668,N_15532);
nand U16326 (N_16326,N_15761,N_15672);
nand U16327 (N_16327,N_15677,N_15824);
or U16328 (N_16328,N_15997,N_15500);
or U16329 (N_16329,N_15565,N_15646);
and U16330 (N_16330,N_15825,N_15561);
and U16331 (N_16331,N_15584,N_15714);
or U16332 (N_16332,N_15735,N_15509);
nand U16333 (N_16333,N_15665,N_15588);
and U16334 (N_16334,N_15973,N_15746);
nand U16335 (N_16335,N_15511,N_15887);
nand U16336 (N_16336,N_15606,N_15954);
or U16337 (N_16337,N_15593,N_15818);
nor U16338 (N_16338,N_15911,N_15877);
xnor U16339 (N_16339,N_15872,N_15724);
nand U16340 (N_16340,N_15750,N_15731);
xor U16341 (N_16341,N_15926,N_15677);
nor U16342 (N_16342,N_15610,N_15751);
or U16343 (N_16343,N_15980,N_15510);
xnor U16344 (N_16344,N_15591,N_15864);
nand U16345 (N_16345,N_15740,N_15998);
nand U16346 (N_16346,N_15615,N_15728);
or U16347 (N_16347,N_15860,N_15717);
or U16348 (N_16348,N_15944,N_15550);
or U16349 (N_16349,N_15993,N_15848);
nor U16350 (N_16350,N_15706,N_15761);
and U16351 (N_16351,N_15648,N_15743);
and U16352 (N_16352,N_15642,N_15625);
nor U16353 (N_16353,N_15557,N_15747);
and U16354 (N_16354,N_15952,N_15861);
and U16355 (N_16355,N_15931,N_15766);
and U16356 (N_16356,N_15882,N_15938);
or U16357 (N_16357,N_15531,N_15714);
nor U16358 (N_16358,N_15973,N_15905);
xor U16359 (N_16359,N_15779,N_15656);
and U16360 (N_16360,N_15927,N_15951);
nand U16361 (N_16361,N_15658,N_15600);
or U16362 (N_16362,N_15980,N_15701);
nand U16363 (N_16363,N_15935,N_15977);
xor U16364 (N_16364,N_15822,N_15940);
or U16365 (N_16365,N_15919,N_15820);
and U16366 (N_16366,N_15597,N_15681);
xnor U16367 (N_16367,N_15591,N_15715);
xor U16368 (N_16368,N_15723,N_15555);
or U16369 (N_16369,N_15801,N_15821);
and U16370 (N_16370,N_15980,N_15909);
and U16371 (N_16371,N_15917,N_15559);
xor U16372 (N_16372,N_15804,N_15781);
and U16373 (N_16373,N_15841,N_15554);
xor U16374 (N_16374,N_15752,N_15919);
or U16375 (N_16375,N_15971,N_15672);
nand U16376 (N_16376,N_15667,N_15936);
and U16377 (N_16377,N_15956,N_15574);
xor U16378 (N_16378,N_15730,N_15953);
and U16379 (N_16379,N_15561,N_15569);
and U16380 (N_16380,N_15619,N_15630);
nand U16381 (N_16381,N_15522,N_15684);
or U16382 (N_16382,N_15620,N_15530);
nand U16383 (N_16383,N_15681,N_15505);
nand U16384 (N_16384,N_15521,N_15703);
or U16385 (N_16385,N_15946,N_15987);
xnor U16386 (N_16386,N_15648,N_15884);
xor U16387 (N_16387,N_15934,N_15563);
and U16388 (N_16388,N_15845,N_15780);
and U16389 (N_16389,N_15879,N_15919);
and U16390 (N_16390,N_15877,N_15633);
or U16391 (N_16391,N_15568,N_15696);
or U16392 (N_16392,N_15586,N_15737);
nor U16393 (N_16393,N_15897,N_15906);
xor U16394 (N_16394,N_15993,N_15691);
nor U16395 (N_16395,N_15902,N_15736);
or U16396 (N_16396,N_15506,N_15979);
nand U16397 (N_16397,N_15708,N_15659);
or U16398 (N_16398,N_15865,N_15909);
nand U16399 (N_16399,N_15713,N_15984);
and U16400 (N_16400,N_15646,N_15947);
xor U16401 (N_16401,N_15695,N_15804);
or U16402 (N_16402,N_15814,N_15555);
xnor U16403 (N_16403,N_15944,N_15949);
or U16404 (N_16404,N_15937,N_15804);
nand U16405 (N_16405,N_15549,N_15740);
nand U16406 (N_16406,N_15632,N_15910);
and U16407 (N_16407,N_15592,N_15781);
nand U16408 (N_16408,N_15604,N_15750);
xor U16409 (N_16409,N_15508,N_15672);
nor U16410 (N_16410,N_15733,N_15913);
or U16411 (N_16411,N_15516,N_15851);
and U16412 (N_16412,N_15703,N_15949);
or U16413 (N_16413,N_15545,N_15964);
xnor U16414 (N_16414,N_15930,N_15628);
and U16415 (N_16415,N_15769,N_15946);
xor U16416 (N_16416,N_15695,N_15877);
and U16417 (N_16417,N_15688,N_15714);
nand U16418 (N_16418,N_15526,N_15986);
xor U16419 (N_16419,N_15952,N_15949);
and U16420 (N_16420,N_15856,N_15913);
or U16421 (N_16421,N_15617,N_15769);
nand U16422 (N_16422,N_15609,N_15945);
nand U16423 (N_16423,N_15950,N_15830);
or U16424 (N_16424,N_15543,N_15633);
nand U16425 (N_16425,N_15811,N_15867);
or U16426 (N_16426,N_15958,N_15868);
and U16427 (N_16427,N_15698,N_15822);
xnor U16428 (N_16428,N_15665,N_15602);
and U16429 (N_16429,N_15692,N_15862);
nand U16430 (N_16430,N_15738,N_15688);
or U16431 (N_16431,N_15795,N_15957);
xor U16432 (N_16432,N_15536,N_15937);
nand U16433 (N_16433,N_15960,N_15534);
nor U16434 (N_16434,N_15913,N_15505);
or U16435 (N_16435,N_15999,N_15670);
or U16436 (N_16436,N_15704,N_15998);
xnor U16437 (N_16437,N_15819,N_15502);
xnor U16438 (N_16438,N_15775,N_15635);
xor U16439 (N_16439,N_15609,N_15768);
nand U16440 (N_16440,N_15541,N_15915);
nand U16441 (N_16441,N_15716,N_15852);
and U16442 (N_16442,N_15982,N_15880);
and U16443 (N_16443,N_15814,N_15641);
or U16444 (N_16444,N_15932,N_15661);
xnor U16445 (N_16445,N_15913,N_15912);
and U16446 (N_16446,N_15766,N_15716);
nand U16447 (N_16447,N_15997,N_15889);
nand U16448 (N_16448,N_15870,N_15546);
nand U16449 (N_16449,N_15589,N_15707);
xor U16450 (N_16450,N_15765,N_15912);
nand U16451 (N_16451,N_15915,N_15982);
xor U16452 (N_16452,N_15732,N_15525);
xnor U16453 (N_16453,N_15955,N_15957);
nand U16454 (N_16454,N_15777,N_15551);
nor U16455 (N_16455,N_15904,N_15920);
nand U16456 (N_16456,N_15527,N_15631);
or U16457 (N_16457,N_15673,N_15852);
xor U16458 (N_16458,N_15674,N_15542);
xnor U16459 (N_16459,N_15894,N_15726);
or U16460 (N_16460,N_15917,N_15794);
xor U16461 (N_16461,N_15804,N_15562);
nand U16462 (N_16462,N_15986,N_15712);
xnor U16463 (N_16463,N_15777,N_15922);
nand U16464 (N_16464,N_15510,N_15830);
or U16465 (N_16465,N_15873,N_15875);
xor U16466 (N_16466,N_15592,N_15790);
nand U16467 (N_16467,N_15840,N_15920);
or U16468 (N_16468,N_15532,N_15536);
xor U16469 (N_16469,N_15542,N_15626);
nor U16470 (N_16470,N_15754,N_15679);
nand U16471 (N_16471,N_15888,N_15526);
xor U16472 (N_16472,N_15889,N_15822);
xor U16473 (N_16473,N_15817,N_15642);
nand U16474 (N_16474,N_15535,N_15847);
nor U16475 (N_16475,N_15996,N_15657);
nor U16476 (N_16476,N_15893,N_15594);
nand U16477 (N_16477,N_15724,N_15829);
or U16478 (N_16478,N_15887,N_15818);
nor U16479 (N_16479,N_15876,N_15808);
xor U16480 (N_16480,N_15612,N_15837);
nand U16481 (N_16481,N_15769,N_15523);
and U16482 (N_16482,N_15746,N_15753);
and U16483 (N_16483,N_15745,N_15669);
xor U16484 (N_16484,N_15786,N_15588);
nand U16485 (N_16485,N_15557,N_15963);
nor U16486 (N_16486,N_15858,N_15995);
or U16487 (N_16487,N_15907,N_15905);
nor U16488 (N_16488,N_15800,N_15653);
nand U16489 (N_16489,N_15865,N_15973);
xnor U16490 (N_16490,N_15610,N_15713);
nor U16491 (N_16491,N_15612,N_15725);
xnor U16492 (N_16492,N_15998,N_15547);
or U16493 (N_16493,N_15641,N_15915);
and U16494 (N_16494,N_15666,N_15529);
or U16495 (N_16495,N_15787,N_15756);
or U16496 (N_16496,N_15510,N_15600);
nand U16497 (N_16497,N_15730,N_15831);
nand U16498 (N_16498,N_15982,N_15599);
nand U16499 (N_16499,N_15536,N_15984);
nand U16500 (N_16500,N_16079,N_16449);
nand U16501 (N_16501,N_16160,N_16401);
or U16502 (N_16502,N_16265,N_16280);
and U16503 (N_16503,N_16292,N_16225);
nand U16504 (N_16504,N_16161,N_16402);
or U16505 (N_16505,N_16195,N_16392);
and U16506 (N_16506,N_16335,N_16259);
or U16507 (N_16507,N_16015,N_16497);
xnor U16508 (N_16508,N_16074,N_16427);
nor U16509 (N_16509,N_16221,N_16474);
nand U16510 (N_16510,N_16033,N_16170);
xnor U16511 (N_16511,N_16260,N_16013);
xnor U16512 (N_16512,N_16168,N_16287);
and U16513 (N_16513,N_16360,N_16438);
nand U16514 (N_16514,N_16247,N_16143);
nor U16515 (N_16515,N_16190,N_16254);
nand U16516 (N_16516,N_16064,N_16141);
xnor U16517 (N_16517,N_16044,N_16258);
nor U16518 (N_16518,N_16413,N_16273);
nor U16519 (N_16519,N_16208,N_16131);
or U16520 (N_16520,N_16086,N_16434);
nor U16521 (N_16521,N_16129,N_16005);
xnor U16522 (N_16522,N_16178,N_16341);
or U16523 (N_16523,N_16472,N_16130);
nand U16524 (N_16524,N_16271,N_16450);
xor U16525 (N_16525,N_16187,N_16183);
or U16526 (N_16526,N_16433,N_16473);
nand U16527 (N_16527,N_16317,N_16337);
or U16528 (N_16528,N_16169,N_16461);
nand U16529 (N_16529,N_16344,N_16493);
or U16530 (N_16530,N_16381,N_16027);
nand U16531 (N_16531,N_16037,N_16175);
nor U16532 (N_16532,N_16336,N_16499);
xor U16533 (N_16533,N_16115,N_16091);
and U16534 (N_16534,N_16243,N_16471);
and U16535 (N_16535,N_16025,N_16238);
or U16536 (N_16536,N_16274,N_16426);
nor U16537 (N_16537,N_16105,N_16107);
xnor U16538 (N_16538,N_16111,N_16241);
nand U16539 (N_16539,N_16496,N_16255);
and U16540 (N_16540,N_16199,N_16355);
and U16541 (N_16541,N_16207,N_16191);
xor U16542 (N_16542,N_16149,N_16332);
xnor U16543 (N_16543,N_16443,N_16420);
nor U16544 (N_16544,N_16491,N_16441);
nand U16545 (N_16545,N_16069,N_16051);
xor U16546 (N_16546,N_16366,N_16132);
or U16547 (N_16547,N_16047,N_16018);
and U16548 (N_16548,N_16387,N_16284);
and U16549 (N_16549,N_16327,N_16429);
or U16550 (N_16550,N_16182,N_16222);
nand U16551 (N_16551,N_16290,N_16093);
or U16552 (N_16552,N_16275,N_16193);
nor U16553 (N_16553,N_16395,N_16328);
nor U16554 (N_16554,N_16237,N_16101);
and U16555 (N_16555,N_16088,N_16068);
and U16556 (N_16556,N_16140,N_16468);
and U16557 (N_16557,N_16278,N_16055);
or U16558 (N_16558,N_16298,N_16148);
and U16559 (N_16559,N_16010,N_16176);
nor U16560 (N_16560,N_16418,N_16021);
xor U16561 (N_16561,N_16397,N_16089);
or U16562 (N_16562,N_16244,N_16030);
nor U16563 (N_16563,N_16293,N_16407);
nor U16564 (N_16564,N_16261,N_16017);
nor U16565 (N_16565,N_16447,N_16145);
nor U16566 (N_16566,N_16362,N_16467);
nor U16567 (N_16567,N_16318,N_16403);
xor U16568 (N_16568,N_16453,N_16215);
or U16569 (N_16569,N_16098,N_16390);
nor U16570 (N_16570,N_16321,N_16478);
nor U16571 (N_16571,N_16349,N_16262);
or U16572 (N_16572,N_16286,N_16266);
nand U16573 (N_16573,N_16489,N_16052);
nor U16574 (N_16574,N_16465,N_16230);
nor U16575 (N_16575,N_16248,N_16269);
xnor U16576 (N_16576,N_16113,N_16108);
nor U16577 (N_16577,N_16001,N_16311);
or U16578 (N_16578,N_16134,N_16151);
xor U16579 (N_16579,N_16307,N_16014);
nand U16580 (N_16580,N_16227,N_16322);
and U16581 (N_16581,N_16167,N_16367);
and U16582 (N_16582,N_16296,N_16029);
nor U16583 (N_16583,N_16379,N_16206);
and U16584 (N_16584,N_16186,N_16184);
nor U16585 (N_16585,N_16439,N_16359);
or U16586 (N_16586,N_16109,N_16155);
nor U16587 (N_16587,N_16120,N_16228);
nor U16588 (N_16588,N_16316,N_16100);
nor U16589 (N_16589,N_16357,N_16118);
xnor U16590 (N_16590,N_16097,N_16022);
nor U16591 (N_16591,N_16048,N_16343);
nor U16592 (N_16592,N_16385,N_16209);
or U16593 (N_16593,N_16409,N_16179);
and U16594 (N_16594,N_16194,N_16095);
or U16595 (N_16595,N_16200,N_16437);
and U16596 (N_16596,N_16481,N_16043);
xor U16597 (N_16597,N_16365,N_16263);
xor U16598 (N_16598,N_16484,N_16204);
and U16599 (N_16599,N_16440,N_16272);
nor U16600 (N_16600,N_16459,N_16174);
nor U16601 (N_16601,N_16210,N_16404);
or U16602 (N_16602,N_16007,N_16342);
and U16603 (N_16603,N_16198,N_16116);
or U16604 (N_16604,N_16487,N_16488);
nor U16605 (N_16605,N_16012,N_16067);
nor U16606 (N_16606,N_16085,N_16235);
nor U16607 (N_16607,N_16137,N_16483);
nand U16608 (N_16608,N_16319,N_16038);
nand U16609 (N_16609,N_16162,N_16495);
and U16610 (N_16610,N_16076,N_16405);
xor U16611 (N_16611,N_16345,N_16425);
and U16612 (N_16612,N_16092,N_16233);
nor U16613 (N_16613,N_16053,N_16417);
and U16614 (N_16614,N_16049,N_16371);
nand U16615 (N_16615,N_16370,N_16331);
or U16616 (N_16616,N_16070,N_16351);
nor U16617 (N_16617,N_16135,N_16333);
and U16618 (N_16618,N_16494,N_16415);
or U16619 (N_16619,N_16348,N_16324);
nand U16620 (N_16620,N_16352,N_16096);
and U16621 (N_16621,N_16119,N_16083);
nand U16622 (N_16622,N_16419,N_16020);
nor U16623 (N_16623,N_16011,N_16398);
and U16624 (N_16624,N_16159,N_16006);
xnor U16625 (N_16625,N_16231,N_16136);
or U16626 (N_16626,N_16264,N_16354);
or U16627 (N_16627,N_16364,N_16312);
and U16628 (N_16628,N_16087,N_16173);
or U16629 (N_16629,N_16466,N_16171);
xor U16630 (N_16630,N_16428,N_16277);
or U16631 (N_16631,N_16300,N_16391);
or U16632 (N_16632,N_16464,N_16445);
or U16633 (N_16633,N_16040,N_16330);
nand U16634 (N_16634,N_16229,N_16374);
or U16635 (N_16635,N_16384,N_16080);
nor U16636 (N_16636,N_16283,N_16114);
or U16637 (N_16637,N_16034,N_16172);
nand U16638 (N_16638,N_16024,N_16216);
nor U16639 (N_16639,N_16454,N_16432);
xnor U16640 (N_16640,N_16389,N_16054);
nor U16641 (N_16641,N_16008,N_16480);
nor U16642 (N_16642,N_16347,N_16185);
nor U16643 (N_16643,N_16456,N_16063);
or U16644 (N_16644,N_16455,N_16072);
or U16645 (N_16645,N_16346,N_16490);
nand U16646 (N_16646,N_16061,N_16126);
nand U16647 (N_16647,N_16106,N_16276);
or U16648 (N_16648,N_16205,N_16469);
nor U16649 (N_16649,N_16081,N_16016);
nor U16650 (N_16650,N_16128,N_16152);
and U16651 (N_16651,N_16125,N_16246);
nand U16652 (N_16652,N_16253,N_16138);
nand U16653 (N_16653,N_16133,N_16485);
and U16654 (N_16654,N_16103,N_16285);
nor U16655 (N_16655,N_16094,N_16380);
nor U16656 (N_16656,N_16462,N_16301);
or U16657 (N_16657,N_16394,N_16060);
nor U16658 (N_16658,N_16482,N_16314);
nor U16659 (N_16659,N_16019,N_16435);
nor U16660 (N_16660,N_16041,N_16486);
nor U16661 (N_16661,N_16122,N_16373);
nor U16662 (N_16662,N_16257,N_16112);
or U16663 (N_16663,N_16234,N_16026);
and U16664 (N_16664,N_16309,N_16201);
nor U16665 (N_16665,N_16153,N_16213);
or U16666 (N_16666,N_16315,N_16142);
and U16667 (N_16667,N_16306,N_16256);
or U16668 (N_16668,N_16323,N_16303);
xor U16669 (N_16669,N_16164,N_16180);
and U16670 (N_16670,N_16028,N_16310);
nand U16671 (N_16671,N_16356,N_16075);
or U16672 (N_16672,N_16304,N_16305);
nor U16673 (N_16673,N_16123,N_16150);
or U16674 (N_16674,N_16416,N_16203);
and U16675 (N_16675,N_16197,N_16004);
and U16676 (N_16676,N_16009,N_16031);
xor U16677 (N_16677,N_16412,N_16476);
and U16678 (N_16678,N_16400,N_16430);
nor U16679 (N_16679,N_16460,N_16039);
nor U16680 (N_16680,N_16165,N_16358);
or U16681 (N_16681,N_16457,N_16406);
xnor U16682 (N_16682,N_16299,N_16369);
nand U16683 (N_16683,N_16372,N_16410);
and U16684 (N_16684,N_16268,N_16214);
and U16685 (N_16685,N_16448,N_16224);
or U16686 (N_16686,N_16196,N_16062);
and U16687 (N_16687,N_16289,N_16382);
nor U16688 (N_16688,N_16117,N_16239);
or U16689 (N_16689,N_16036,N_16212);
nor U16690 (N_16690,N_16188,N_16334);
or U16691 (N_16691,N_16361,N_16000);
and U16692 (N_16692,N_16057,N_16383);
and U16693 (N_16693,N_16032,N_16463);
xor U16694 (N_16694,N_16045,N_16078);
nand U16695 (N_16695,N_16393,N_16219);
xnor U16696 (N_16696,N_16326,N_16090);
nand U16697 (N_16697,N_16424,N_16442);
xor U16698 (N_16698,N_16320,N_16077);
and U16699 (N_16699,N_16250,N_16073);
or U16700 (N_16700,N_16408,N_16154);
nand U16701 (N_16701,N_16378,N_16375);
and U16702 (N_16702,N_16281,N_16279);
xnor U16703 (N_16703,N_16340,N_16399);
xor U16704 (N_16704,N_16189,N_16127);
nor U16705 (N_16705,N_16377,N_16308);
nor U16706 (N_16706,N_16302,N_16084);
nand U16707 (N_16707,N_16002,N_16050);
nand U16708 (N_16708,N_16065,N_16339);
xnor U16709 (N_16709,N_16217,N_16414);
and U16710 (N_16710,N_16350,N_16245);
or U16711 (N_16711,N_16270,N_16156);
nand U16712 (N_16712,N_16252,N_16421);
nor U16713 (N_16713,N_16056,N_16313);
nor U16714 (N_16714,N_16329,N_16376);
and U16715 (N_16715,N_16232,N_16035);
nor U16716 (N_16716,N_16436,N_16192);
nor U16717 (N_16717,N_16059,N_16223);
xnor U16718 (N_16718,N_16282,N_16363);
xor U16719 (N_16719,N_16338,N_16422);
and U16720 (N_16720,N_16158,N_16166);
and U16721 (N_16721,N_16470,N_16444);
nor U16722 (N_16722,N_16295,N_16236);
nor U16723 (N_16723,N_16446,N_16368);
or U16724 (N_16724,N_16411,N_16388);
nor U16725 (N_16725,N_16042,N_16297);
nor U16726 (N_16726,N_16181,N_16082);
xnor U16727 (N_16727,N_16251,N_16492);
or U16728 (N_16728,N_16353,N_16211);
nand U16729 (N_16729,N_16202,N_16157);
nand U16730 (N_16730,N_16475,N_16003);
nor U16731 (N_16731,N_16071,N_16226);
and U16732 (N_16732,N_16451,N_16121);
nand U16733 (N_16733,N_16218,N_16294);
nand U16734 (N_16734,N_16249,N_16177);
or U16735 (N_16735,N_16139,N_16110);
nand U16736 (N_16736,N_16104,N_16046);
nand U16737 (N_16737,N_16023,N_16452);
and U16738 (N_16738,N_16146,N_16288);
xnor U16739 (N_16739,N_16431,N_16099);
nor U16740 (N_16740,N_16144,N_16220);
or U16741 (N_16741,N_16325,N_16102);
nand U16742 (N_16742,N_16147,N_16458);
or U16743 (N_16743,N_16423,N_16386);
or U16744 (N_16744,N_16124,N_16163);
xnor U16745 (N_16745,N_16396,N_16240);
nand U16746 (N_16746,N_16477,N_16291);
nor U16747 (N_16747,N_16498,N_16058);
nand U16748 (N_16748,N_16242,N_16066);
xor U16749 (N_16749,N_16267,N_16479);
and U16750 (N_16750,N_16145,N_16423);
xnor U16751 (N_16751,N_16466,N_16470);
nor U16752 (N_16752,N_16197,N_16382);
nand U16753 (N_16753,N_16134,N_16157);
and U16754 (N_16754,N_16300,N_16395);
xor U16755 (N_16755,N_16197,N_16389);
nor U16756 (N_16756,N_16428,N_16154);
nor U16757 (N_16757,N_16356,N_16236);
xnor U16758 (N_16758,N_16017,N_16298);
or U16759 (N_16759,N_16336,N_16449);
nand U16760 (N_16760,N_16489,N_16449);
and U16761 (N_16761,N_16454,N_16281);
xnor U16762 (N_16762,N_16281,N_16387);
nor U16763 (N_16763,N_16170,N_16394);
or U16764 (N_16764,N_16297,N_16205);
nand U16765 (N_16765,N_16384,N_16199);
nor U16766 (N_16766,N_16194,N_16123);
nor U16767 (N_16767,N_16467,N_16041);
nor U16768 (N_16768,N_16169,N_16349);
xor U16769 (N_16769,N_16254,N_16020);
nor U16770 (N_16770,N_16121,N_16335);
or U16771 (N_16771,N_16441,N_16127);
nand U16772 (N_16772,N_16079,N_16109);
nor U16773 (N_16773,N_16487,N_16384);
nor U16774 (N_16774,N_16079,N_16263);
or U16775 (N_16775,N_16079,N_16157);
xor U16776 (N_16776,N_16437,N_16319);
or U16777 (N_16777,N_16057,N_16035);
nand U16778 (N_16778,N_16117,N_16298);
or U16779 (N_16779,N_16075,N_16003);
nor U16780 (N_16780,N_16482,N_16156);
xor U16781 (N_16781,N_16303,N_16428);
or U16782 (N_16782,N_16174,N_16234);
xor U16783 (N_16783,N_16105,N_16005);
xor U16784 (N_16784,N_16443,N_16304);
nor U16785 (N_16785,N_16087,N_16197);
or U16786 (N_16786,N_16105,N_16179);
nand U16787 (N_16787,N_16460,N_16333);
xnor U16788 (N_16788,N_16170,N_16295);
or U16789 (N_16789,N_16430,N_16134);
xor U16790 (N_16790,N_16178,N_16054);
nor U16791 (N_16791,N_16272,N_16067);
nand U16792 (N_16792,N_16044,N_16240);
xnor U16793 (N_16793,N_16028,N_16488);
nor U16794 (N_16794,N_16173,N_16205);
and U16795 (N_16795,N_16378,N_16463);
nor U16796 (N_16796,N_16080,N_16180);
or U16797 (N_16797,N_16199,N_16256);
xor U16798 (N_16798,N_16474,N_16464);
and U16799 (N_16799,N_16050,N_16475);
and U16800 (N_16800,N_16130,N_16070);
or U16801 (N_16801,N_16036,N_16333);
or U16802 (N_16802,N_16096,N_16338);
nor U16803 (N_16803,N_16394,N_16174);
nand U16804 (N_16804,N_16153,N_16421);
xor U16805 (N_16805,N_16119,N_16346);
nand U16806 (N_16806,N_16372,N_16390);
nand U16807 (N_16807,N_16300,N_16438);
nor U16808 (N_16808,N_16203,N_16356);
nand U16809 (N_16809,N_16259,N_16446);
and U16810 (N_16810,N_16117,N_16032);
nand U16811 (N_16811,N_16210,N_16363);
and U16812 (N_16812,N_16142,N_16322);
nor U16813 (N_16813,N_16251,N_16313);
or U16814 (N_16814,N_16204,N_16263);
nand U16815 (N_16815,N_16447,N_16289);
and U16816 (N_16816,N_16313,N_16170);
xnor U16817 (N_16817,N_16319,N_16206);
nor U16818 (N_16818,N_16195,N_16095);
nor U16819 (N_16819,N_16482,N_16347);
and U16820 (N_16820,N_16314,N_16301);
xor U16821 (N_16821,N_16208,N_16364);
and U16822 (N_16822,N_16419,N_16093);
and U16823 (N_16823,N_16006,N_16057);
nand U16824 (N_16824,N_16377,N_16246);
nor U16825 (N_16825,N_16467,N_16488);
xnor U16826 (N_16826,N_16472,N_16078);
or U16827 (N_16827,N_16076,N_16272);
nor U16828 (N_16828,N_16168,N_16030);
and U16829 (N_16829,N_16014,N_16473);
nor U16830 (N_16830,N_16441,N_16293);
nand U16831 (N_16831,N_16308,N_16132);
nor U16832 (N_16832,N_16407,N_16202);
nand U16833 (N_16833,N_16311,N_16303);
xor U16834 (N_16834,N_16464,N_16061);
nand U16835 (N_16835,N_16047,N_16231);
and U16836 (N_16836,N_16049,N_16325);
xor U16837 (N_16837,N_16069,N_16206);
nand U16838 (N_16838,N_16411,N_16272);
and U16839 (N_16839,N_16345,N_16142);
or U16840 (N_16840,N_16479,N_16089);
and U16841 (N_16841,N_16245,N_16394);
xnor U16842 (N_16842,N_16458,N_16421);
xor U16843 (N_16843,N_16473,N_16432);
nor U16844 (N_16844,N_16201,N_16262);
or U16845 (N_16845,N_16365,N_16417);
xnor U16846 (N_16846,N_16488,N_16228);
or U16847 (N_16847,N_16108,N_16130);
and U16848 (N_16848,N_16342,N_16110);
or U16849 (N_16849,N_16045,N_16044);
xor U16850 (N_16850,N_16456,N_16433);
nor U16851 (N_16851,N_16251,N_16257);
nand U16852 (N_16852,N_16105,N_16319);
and U16853 (N_16853,N_16249,N_16127);
xnor U16854 (N_16854,N_16216,N_16259);
and U16855 (N_16855,N_16161,N_16327);
nand U16856 (N_16856,N_16324,N_16223);
and U16857 (N_16857,N_16078,N_16244);
and U16858 (N_16858,N_16132,N_16332);
and U16859 (N_16859,N_16193,N_16224);
or U16860 (N_16860,N_16493,N_16397);
and U16861 (N_16861,N_16418,N_16130);
xnor U16862 (N_16862,N_16283,N_16176);
nand U16863 (N_16863,N_16358,N_16347);
nand U16864 (N_16864,N_16189,N_16427);
nand U16865 (N_16865,N_16364,N_16224);
nand U16866 (N_16866,N_16432,N_16356);
nor U16867 (N_16867,N_16356,N_16273);
and U16868 (N_16868,N_16279,N_16269);
or U16869 (N_16869,N_16066,N_16268);
and U16870 (N_16870,N_16408,N_16264);
nor U16871 (N_16871,N_16160,N_16028);
xnor U16872 (N_16872,N_16102,N_16315);
xor U16873 (N_16873,N_16306,N_16150);
nor U16874 (N_16874,N_16469,N_16182);
xor U16875 (N_16875,N_16212,N_16070);
xor U16876 (N_16876,N_16106,N_16033);
nor U16877 (N_16877,N_16006,N_16126);
xnor U16878 (N_16878,N_16046,N_16370);
nor U16879 (N_16879,N_16365,N_16189);
nand U16880 (N_16880,N_16195,N_16447);
nor U16881 (N_16881,N_16059,N_16320);
nand U16882 (N_16882,N_16072,N_16395);
xor U16883 (N_16883,N_16269,N_16307);
nand U16884 (N_16884,N_16110,N_16134);
xnor U16885 (N_16885,N_16326,N_16148);
xor U16886 (N_16886,N_16219,N_16067);
and U16887 (N_16887,N_16454,N_16254);
xnor U16888 (N_16888,N_16005,N_16312);
or U16889 (N_16889,N_16457,N_16316);
nand U16890 (N_16890,N_16485,N_16149);
or U16891 (N_16891,N_16383,N_16108);
and U16892 (N_16892,N_16375,N_16332);
nor U16893 (N_16893,N_16024,N_16123);
and U16894 (N_16894,N_16262,N_16411);
xnor U16895 (N_16895,N_16129,N_16382);
and U16896 (N_16896,N_16113,N_16015);
and U16897 (N_16897,N_16460,N_16081);
and U16898 (N_16898,N_16357,N_16106);
nor U16899 (N_16899,N_16006,N_16199);
and U16900 (N_16900,N_16249,N_16331);
nor U16901 (N_16901,N_16126,N_16090);
nand U16902 (N_16902,N_16047,N_16256);
nand U16903 (N_16903,N_16275,N_16024);
and U16904 (N_16904,N_16202,N_16428);
or U16905 (N_16905,N_16239,N_16430);
nand U16906 (N_16906,N_16296,N_16244);
and U16907 (N_16907,N_16049,N_16152);
xor U16908 (N_16908,N_16362,N_16464);
nor U16909 (N_16909,N_16060,N_16037);
nor U16910 (N_16910,N_16215,N_16239);
or U16911 (N_16911,N_16009,N_16455);
or U16912 (N_16912,N_16473,N_16116);
and U16913 (N_16913,N_16093,N_16191);
and U16914 (N_16914,N_16417,N_16124);
or U16915 (N_16915,N_16399,N_16495);
nor U16916 (N_16916,N_16303,N_16294);
or U16917 (N_16917,N_16294,N_16044);
nand U16918 (N_16918,N_16347,N_16490);
or U16919 (N_16919,N_16009,N_16168);
nor U16920 (N_16920,N_16231,N_16206);
nor U16921 (N_16921,N_16268,N_16251);
xor U16922 (N_16922,N_16343,N_16212);
xor U16923 (N_16923,N_16439,N_16210);
nand U16924 (N_16924,N_16313,N_16478);
xnor U16925 (N_16925,N_16207,N_16379);
or U16926 (N_16926,N_16340,N_16131);
or U16927 (N_16927,N_16391,N_16027);
nand U16928 (N_16928,N_16238,N_16146);
xor U16929 (N_16929,N_16123,N_16184);
and U16930 (N_16930,N_16094,N_16333);
nand U16931 (N_16931,N_16013,N_16025);
nor U16932 (N_16932,N_16086,N_16481);
nand U16933 (N_16933,N_16123,N_16237);
or U16934 (N_16934,N_16390,N_16180);
nor U16935 (N_16935,N_16239,N_16012);
xor U16936 (N_16936,N_16426,N_16285);
nor U16937 (N_16937,N_16429,N_16140);
nand U16938 (N_16938,N_16104,N_16294);
nand U16939 (N_16939,N_16131,N_16039);
and U16940 (N_16940,N_16331,N_16106);
nor U16941 (N_16941,N_16152,N_16299);
or U16942 (N_16942,N_16097,N_16237);
xor U16943 (N_16943,N_16333,N_16256);
xor U16944 (N_16944,N_16297,N_16022);
nand U16945 (N_16945,N_16487,N_16263);
nand U16946 (N_16946,N_16283,N_16396);
and U16947 (N_16947,N_16136,N_16226);
nor U16948 (N_16948,N_16186,N_16116);
or U16949 (N_16949,N_16052,N_16442);
or U16950 (N_16950,N_16481,N_16130);
or U16951 (N_16951,N_16212,N_16380);
nor U16952 (N_16952,N_16357,N_16055);
or U16953 (N_16953,N_16381,N_16108);
nand U16954 (N_16954,N_16061,N_16015);
or U16955 (N_16955,N_16050,N_16453);
or U16956 (N_16956,N_16230,N_16378);
nor U16957 (N_16957,N_16203,N_16057);
nand U16958 (N_16958,N_16053,N_16113);
and U16959 (N_16959,N_16233,N_16314);
xor U16960 (N_16960,N_16006,N_16379);
xnor U16961 (N_16961,N_16063,N_16289);
and U16962 (N_16962,N_16301,N_16342);
xnor U16963 (N_16963,N_16249,N_16333);
nand U16964 (N_16964,N_16416,N_16244);
nor U16965 (N_16965,N_16199,N_16069);
and U16966 (N_16966,N_16374,N_16184);
xnor U16967 (N_16967,N_16408,N_16440);
or U16968 (N_16968,N_16323,N_16477);
or U16969 (N_16969,N_16024,N_16329);
nand U16970 (N_16970,N_16243,N_16082);
nand U16971 (N_16971,N_16350,N_16427);
xnor U16972 (N_16972,N_16391,N_16037);
xnor U16973 (N_16973,N_16028,N_16349);
nand U16974 (N_16974,N_16208,N_16400);
and U16975 (N_16975,N_16209,N_16498);
or U16976 (N_16976,N_16041,N_16000);
or U16977 (N_16977,N_16440,N_16316);
xor U16978 (N_16978,N_16034,N_16230);
nand U16979 (N_16979,N_16233,N_16103);
xnor U16980 (N_16980,N_16086,N_16313);
and U16981 (N_16981,N_16429,N_16258);
nor U16982 (N_16982,N_16146,N_16428);
xor U16983 (N_16983,N_16482,N_16473);
xnor U16984 (N_16984,N_16182,N_16142);
and U16985 (N_16985,N_16457,N_16369);
nand U16986 (N_16986,N_16494,N_16350);
nand U16987 (N_16987,N_16290,N_16174);
nand U16988 (N_16988,N_16404,N_16392);
and U16989 (N_16989,N_16469,N_16282);
nand U16990 (N_16990,N_16291,N_16063);
xor U16991 (N_16991,N_16369,N_16492);
nand U16992 (N_16992,N_16114,N_16182);
nand U16993 (N_16993,N_16053,N_16143);
or U16994 (N_16994,N_16120,N_16473);
and U16995 (N_16995,N_16284,N_16160);
xor U16996 (N_16996,N_16012,N_16133);
xnor U16997 (N_16997,N_16154,N_16437);
and U16998 (N_16998,N_16082,N_16131);
or U16999 (N_16999,N_16197,N_16376);
xor U17000 (N_17000,N_16895,N_16859);
nand U17001 (N_17001,N_16936,N_16643);
or U17002 (N_17002,N_16552,N_16650);
nor U17003 (N_17003,N_16724,N_16710);
or U17004 (N_17004,N_16907,N_16788);
or U17005 (N_17005,N_16686,N_16893);
xnor U17006 (N_17006,N_16598,N_16974);
nor U17007 (N_17007,N_16933,N_16753);
and U17008 (N_17008,N_16688,N_16916);
nor U17009 (N_17009,N_16756,N_16655);
xor U17010 (N_17010,N_16969,N_16563);
nor U17011 (N_17011,N_16813,N_16910);
nand U17012 (N_17012,N_16755,N_16508);
or U17013 (N_17013,N_16944,N_16727);
nor U17014 (N_17014,N_16808,N_16978);
and U17015 (N_17015,N_16578,N_16677);
xnor U17016 (N_17016,N_16558,N_16805);
or U17017 (N_17017,N_16719,N_16676);
nor U17018 (N_17018,N_16664,N_16751);
xnor U17019 (N_17019,N_16990,N_16546);
nand U17020 (N_17020,N_16564,N_16766);
nor U17021 (N_17021,N_16775,N_16601);
xnor U17022 (N_17022,N_16663,N_16966);
nand U17023 (N_17023,N_16887,N_16784);
and U17024 (N_17024,N_16603,N_16848);
and U17025 (N_17025,N_16674,N_16732);
nand U17026 (N_17026,N_16994,N_16604);
or U17027 (N_17027,N_16747,N_16891);
nand U17028 (N_17028,N_16696,N_16524);
and U17029 (N_17029,N_16595,N_16768);
nor U17030 (N_17030,N_16807,N_16960);
or U17031 (N_17031,N_16884,N_16901);
or U17032 (N_17032,N_16894,N_16925);
and U17033 (N_17033,N_16685,N_16689);
or U17034 (N_17034,N_16928,N_16659);
nand U17035 (N_17035,N_16568,N_16919);
nor U17036 (N_17036,N_16512,N_16608);
and U17037 (N_17037,N_16758,N_16804);
nand U17038 (N_17038,N_16959,N_16577);
xor U17039 (N_17039,N_16941,N_16507);
xor U17040 (N_17040,N_16557,N_16708);
nor U17041 (N_17041,N_16729,N_16678);
nor U17042 (N_17042,N_16583,N_16647);
or U17043 (N_17043,N_16717,N_16556);
nand U17044 (N_17044,N_16544,N_16826);
nor U17045 (N_17045,N_16971,N_16581);
and U17046 (N_17046,N_16737,N_16913);
nor U17047 (N_17047,N_16930,N_16923);
nor U17048 (N_17048,N_16818,N_16856);
or U17049 (N_17049,N_16954,N_16612);
nand U17050 (N_17050,N_16860,N_16855);
or U17051 (N_17051,N_16515,N_16638);
or U17052 (N_17052,N_16709,N_16740);
and U17053 (N_17053,N_16824,N_16942);
and U17054 (N_17054,N_16926,N_16730);
and U17055 (N_17055,N_16857,N_16833);
xnor U17056 (N_17056,N_16949,N_16772);
or U17057 (N_17057,N_16531,N_16550);
and U17058 (N_17058,N_16782,N_16800);
and U17059 (N_17059,N_16796,N_16774);
nand U17060 (N_17060,N_16523,N_16757);
nand U17061 (N_17061,N_16665,N_16870);
and U17062 (N_17062,N_16844,N_16554);
nor U17063 (N_17063,N_16513,N_16864);
nor U17064 (N_17064,N_16537,N_16828);
xor U17065 (N_17065,N_16921,N_16605);
nor U17066 (N_17066,N_16549,N_16632);
nand U17067 (N_17067,N_16534,N_16705);
and U17068 (N_17068,N_16720,N_16946);
or U17069 (N_17069,N_16816,N_16871);
nor U17070 (N_17070,N_16885,N_16883);
nand U17071 (N_17071,N_16505,N_16561);
xnor U17072 (N_17072,N_16511,N_16514);
nor U17073 (N_17073,N_16504,N_16914);
nor U17074 (N_17074,N_16763,N_16517);
or U17075 (N_17075,N_16792,N_16892);
or U17076 (N_17076,N_16559,N_16692);
nor U17077 (N_17077,N_16915,N_16952);
nor U17078 (N_17078,N_16723,N_16634);
or U17079 (N_17079,N_16739,N_16527);
nand U17080 (N_17080,N_16849,N_16526);
xor U17081 (N_17081,N_16831,N_16794);
xnor U17082 (N_17082,N_16721,N_16789);
nand U17083 (N_17083,N_16519,N_16759);
or U17084 (N_17084,N_16798,N_16786);
and U17085 (N_17085,N_16738,N_16728);
nor U17086 (N_17086,N_16834,N_16840);
nor U17087 (N_17087,N_16842,N_16636);
nor U17088 (N_17088,N_16745,N_16991);
nand U17089 (N_17089,N_16722,N_16889);
and U17090 (N_17090,N_16779,N_16585);
xnor U17091 (N_17091,N_16836,N_16879);
or U17092 (N_17092,N_16701,N_16725);
and U17093 (N_17093,N_16547,N_16579);
xnor U17094 (N_17094,N_16839,N_16847);
xor U17095 (N_17095,N_16961,N_16752);
xnor U17096 (N_17096,N_16771,N_16982);
nor U17097 (N_17097,N_16580,N_16811);
nor U17098 (N_17098,N_16851,N_16918);
nand U17099 (N_17099,N_16897,N_16555);
xor U17100 (N_17100,N_16814,N_16642);
xor U17101 (N_17101,N_16702,N_16861);
xnor U17102 (N_17102,N_16645,N_16648);
and U17103 (N_17103,N_16661,N_16633);
nor U17104 (N_17104,N_16778,N_16781);
and U17105 (N_17105,N_16687,N_16509);
nand U17106 (N_17106,N_16637,N_16525);
nand U17107 (N_17107,N_16518,N_16905);
nand U17108 (N_17108,N_16596,N_16968);
xor U17109 (N_17109,N_16592,N_16572);
nor U17110 (N_17110,N_16651,N_16510);
nand U17111 (N_17111,N_16715,N_16931);
and U17112 (N_17112,N_16667,N_16690);
or U17113 (N_17113,N_16875,N_16629);
or U17114 (N_17114,N_16657,N_16570);
nand U17115 (N_17115,N_16573,N_16750);
or U17116 (N_17116,N_16618,N_16821);
xnor U17117 (N_17117,N_16769,N_16791);
or U17118 (N_17118,N_16909,N_16520);
nor U17119 (N_17119,N_16736,N_16924);
xnor U17120 (N_17120,N_16770,N_16869);
xnor U17121 (N_17121,N_16972,N_16516);
nor U17122 (N_17122,N_16530,N_16830);
nor U17123 (N_17123,N_16929,N_16673);
nor U17124 (N_17124,N_16854,N_16850);
or U17125 (N_17125,N_16669,N_16627);
xnor U17126 (N_17126,N_16992,N_16899);
and U17127 (N_17127,N_16876,N_16761);
nand U17128 (N_17128,N_16743,N_16939);
and U17129 (N_17129,N_16541,N_16917);
xor U17130 (N_17130,N_16660,N_16963);
and U17131 (N_17131,N_16584,N_16588);
and U17132 (N_17132,N_16841,N_16858);
xor U17133 (N_17133,N_16896,N_16666);
and U17134 (N_17134,N_16704,N_16746);
xor U17135 (N_17135,N_16668,N_16565);
or U17136 (N_17136,N_16987,N_16589);
xor U17137 (N_17137,N_16560,N_16908);
and U17138 (N_17138,N_16873,N_16631);
nor U17139 (N_17139,N_16812,N_16881);
or U17140 (N_17140,N_16548,N_16874);
nand U17141 (N_17141,N_16865,N_16853);
nor U17142 (N_17142,N_16962,N_16543);
nand U17143 (N_17143,N_16695,N_16846);
or U17144 (N_17144,N_16607,N_16571);
and U17145 (N_17145,N_16538,N_16681);
nand U17146 (N_17146,N_16569,N_16947);
nand U17147 (N_17147,N_16979,N_16935);
nor U17148 (N_17148,N_16641,N_16981);
or U17149 (N_17149,N_16780,N_16773);
or U17150 (N_17150,N_16802,N_16996);
xor U17151 (N_17151,N_16953,N_16640);
xor U17152 (N_17152,N_16888,N_16906);
nand U17153 (N_17153,N_16820,N_16653);
and U17154 (N_17154,N_16619,N_16613);
nor U17155 (N_17155,N_16733,N_16711);
or U17156 (N_17156,N_16767,N_16716);
xor U17157 (N_17157,N_16670,N_16652);
xnor U17158 (N_17158,N_16799,N_16591);
xnor U17159 (N_17159,N_16691,N_16989);
xor U17160 (N_17160,N_16958,N_16997);
xor U17161 (N_17161,N_16683,N_16940);
or U17162 (N_17162,N_16600,N_16658);
or U17163 (N_17163,N_16809,N_16706);
xnor U17164 (N_17164,N_16934,N_16882);
xnor U17165 (N_17165,N_16500,N_16718);
xnor U17166 (N_17166,N_16587,N_16562);
or U17167 (N_17167,N_16662,N_16622);
xnor U17168 (N_17168,N_16693,N_16922);
nor U17169 (N_17169,N_16748,N_16582);
nand U17170 (N_17170,N_16983,N_16726);
nor U17171 (N_17171,N_16503,N_16599);
xor U17172 (N_17172,N_16542,N_16810);
nor U17173 (N_17173,N_16575,N_16528);
nand U17174 (N_17174,N_16819,N_16602);
nor U17175 (N_17175,N_16694,N_16988);
or U17176 (N_17176,N_16529,N_16630);
nand U17177 (N_17177,N_16617,N_16540);
nor U17178 (N_17178,N_16644,N_16938);
nand U17179 (N_17179,N_16815,N_16976);
xor U17180 (N_17180,N_16998,N_16521);
xnor U17181 (N_17181,N_16535,N_16593);
and U17182 (N_17182,N_16679,N_16795);
and U17183 (N_17183,N_16606,N_16539);
or U17184 (N_17184,N_16522,N_16867);
xor U17185 (N_17185,N_16903,N_16964);
nand U17186 (N_17186,N_16700,N_16806);
xor U17187 (N_17187,N_16698,N_16880);
xor U17188 (N_17188,N_16999,N_16623);
or U17189 (N_17189,N_16551,N_16912);
or U17190 (N_17190,N_16793,N_16862);
or U17191 (N_17191,N_16672,N_16506);
xnor U17192 (N_17192,N_16586,N_16948);
and U17193 (N_17193,N_16590,N_16735);
nor U17194 (N_17194,N_16945,N_16615);
and U17195 (N_17195,N_16843,N_16731);
and U17196 (N_17196,N_16980,N_16754);
or U17197 (N_17197,N_16984,N_16832);
xor U17198 (N_17198,N_16911,N_16951);
xor U17199 (N_17199,N_16975,N_16712);
nand U17200 (N_17200,N_16898,N_16823);
xnor U17201 (N_17201,N_16625,N_16713);
or U17202 (N_17202,N_16878,N_16868);
nand U17203 (N_17203,N_16621,N_16682);
and U17204 (N_17204,N_16801,N_16533);
nand U17205 (N_17205,N_16734,N_16852);
xnor U17206 (N_17206,N_16785,N_16872);
xor U17207 (N_17207,N_16610,N_16699);
nor U17208 (N_17208,N_16635,N_16822);
nor U17209 (N_17209,N_16703,N_16797);
or U17210 (N_17210,N_16646,N_16576);
nand U17211 (N_17211,N_16943,N_16765);
and U17212 (N_17212,N_16609,N_16762);
xor U17213 (N_17213,N_16827,N_16900);
nor U17214 (N_17214,N_16967,N_16567);
nand U17215 (N_17215,N_16532,N_16863);
and U17216 (N_17216,N_16680,N_16626);
nor U17217 (N_17217,N_16714,N_16744);
or U17218 (N_17218,N_16993,N_16838);
and U17219 (N_17219,N_16611,N_16937);
xnor U17220 (N_17220,N_16671,N_16639);
and U17221 (N_17221,N_16920,N_16985);
and U17222 (N_17222,N_16742,N_16986);
nor U17223 (N_17223,N_16835,N_16656);
and U17224 (N_17224,N_16536,N_16825);
nor U17225 (N_17225,N_16886,N_16955);
and U17226 (N_17226,N_16553,N_16877);
nand U17227 (N_17227,N_16957,N_16829);
or U17228 (N_17228,N_16904,N_16866);
nand U17229 (N_17229,N_16890,N_16817);
xnor U17230 (N_17230,N_16614,N_16950);
nand U17231 (N_17231,N_16749,N_16616);
xor U17232 (N_17232,N_16654,N_16502);
nand U17233 (N_17233,N_16675,N_16684);
nand U17234 (N_17234,N_16927,N_16597);
nand U17235 (N_17235,N_16837,N_16956);
nand U17236 (N_17236,N_16777,N_16566);
nor U17237 (N_17237,N_16741,N_16760);
nor U17238 (N_17238,N_16620,N_16977);
nand U17239 (N_17239,N_16932,N_16628);
or U17240 (N_17240,N_16545,N_16783);
nor U17241 (N_17241,N_16776,N_16707);
nand U17242 (N_17242,N_16790,N_16649);
nand U17243 (N_17243,N_16574,N_16803);
and U17244 (N_17244,N_16624,N_16965);
and U17245 (N_17245,N_16902,N_16697);
nand U17246 (N_17246,N_16845,N_16764);
or U17247 (N_17247,N_16970,N_16973);
and U17248 (N_17248,N_16594,N_16995);
nor U17249 (N_17249,N_16787,N_16501);
nor U17250 (N_17250,N_16879,N_16895);
and U17251 (N_17251,N_16604,N_16911);
xor U17252 (N_17252,N_16979,N_16998);
nor U17253 (N_17253,N_16933,N_16939);
nor U17254 (N_17254,N_16851,N_16999);
and U17255 (N_17255,N_16973,N_16590);
and U17256 (N_17256,N_16773,N_16633);
nand U17257 (N_17257,N_16521,N_16776);
xnor U17258 (N_17258,N_16856,N_16774);
nand U17259 (N_17259,N_16524,N_16722);
nor U17260 (N_17260,N_16805,N_16997);
xnor U17261 (N_17261,N_16936,N_16529);
xor U17262 (N_17262,N_16960,N_16718);
nor U17263 (N_17263,N_16740,N_16970);
nor U17264 (N_17264,N_16732,N_16563);
xnor U17265 (N_17265,N_16528,N_16814);
nand U17266 (N_17266,N_16933,N_16573);
and U17267 (N_17267,N_16639,N_16939);
xnor U17268 (N_17268,N_16503,N_16948);
or U17269 (N_17269,N_16793,N_16715);
nor U17270 (N_17270,N_16772,N_16807);
nor U17271 (N_17271,N_16570,N_16942);
nor U17272 (N_17272,N_16963,N_16627);
or U17273 (N_17273,N_16677,N_16591);
or U17274 (N_17274,N_16994,N_16575);
nor U17275 (N_17275,N_16982,N_16745);
nor U17276 (N_17276,N_16687,N_16640);
or U17277 (N_17277,N_16577,N_16894);
or U17278 (N_17278,N_16774,N_16726);
nand U17279 (N_17279,N_16669,N_16989);
or U17280 (N_17280,N_16615,N_16575);
and U17281 (N_17281,N_16712,N_16536);
or U17282 (N_17282,N_16685,N_16676);
xor U17283 (N_17283,N_16744,N_16549);
nor U17284 (N_17284,N_16694,N_16927);
nand U17285 (N_17285,N_16581,N_16596);
or U17286 (N_17286,N_16603,N_16771);
nor U17287 (N_17287,N_16968,N_16821);
and U17288 (N_17288,N_16989,N_16747);
nand U17289 (N_17289,N_16832,N_16888);
nor U17290 (N_17290,N_16611,N_16796);
xor U17291 (N_17291,N_16783,N_16822);
nand U17292 (N_17292,N_16842,N_16769);
nor U17293 (N_17293,N_16584,N_16626);
xor U17294 (N_17294,N_16660,N_16970);
xor U17295 (N_17295,N_16941,N_16572);
nor U17296 (N_17296,N_16690,N_16665);
nor U17297 (N_17297,N_16535,N_16788);
and U17298 (N_17298,N_16827,N_16815);
or U17299 (N_17299,N_16982,N_16570);
xnor U17300 (N_17300,N_16804,N_16566);
or U17301 (N_17301,N_16722,N_16806);
or U17302 (N_17302,N_16801,N_16774);
and U17303 (N_17303,N_16620,N_16607);
nor U17304 (N_17304,N_16845,N_16879);
xnor U17305 (N_17305,N_16770,N_16713);
nor U17306 (N_17306,N_16842,N_16980);
xnor U17307 (N_17307,N_16523,N_16916);
or U17308 (N_17308,N_16962,N_16607);
or U17309 (N_17309,N_16766,N_16610);
nand U17310 (N_17310,N_16802,N_16649);
nand U17311 (N_17311,N_16790,N_16885);
nor U17312 (N_17312,N_16695,N_16738);
and U17313 (N_17313,N_16794,N_16511);
and U17314 (N_17314,N_16905,N_16759);
and U17315 (N_17315,N_16641,N_16819);
nor U17316 (N_17316,N_16820,N_16948);
or U17317 (N_17317,N_16939,N_16991);
nor U17318 (N_17318,N_16503,N_16777);
xnor U17319 (N_17319,N_16537,N_16582);
xnor U17320 (N_17320,N_16538,N_16583);
nand U17321 (N_17321,N_16878,N_16986);
nor U17322 (N_17322,N_16690,N_16911);
or U17323 (N_17323,N_16968,N_16925);
xor U17324 (N_17324,N_16576,N_16687);
nor U17325 (N_17325,N_16852,N_16517);
nand U17326 (N_17326,N_16863,N_16653);
xnor U17327 (N_17327,N_16903,N_16578);
nor U17328 (N_17328,N_16972,N_16695);
and U17329 (N_17329,N_16605,N_16927);
and U17330 (N_17330,N_16950,N_16794);
nand U17331 (N_17331,N_16552,N_16793);
xor U17332 (N_17332,N_16929,N_16674);
or U17333 (N_17333,N_16958,N_16939);
or U17334 (N_17334,N_16984,N_16634);
nor U17335 (N_17335,N_16571,N_16991);
xnor U17336 (N_17336,N_16688,N_16543);
nand U17337 (N_17337,N_16587,N_16758);
xor U17338 (N_17338,N_16533,N_16851);
nor U17339 (N_17339,N_16585,N_16500);
nor U17340 (N_17340,N_16705,N_16883);
nor U17341 (N_17341,N_16804,N_16626);
and U17342 (N_17342,N_16967,N_16733);
nand U17343 (N_17343,N_16980,N_16984);
and U17344 (N_17344,N_16945,N_16713);
xnor U17345 (N_17345,N_16916,N_16985);
or U17346 (N_17346,N_16624,N_16926);
xnor U17347 (N_17347,N_16825,N_16767);
nor U17348 (N_17348,N_16875,N_16772);
or U17349 (N_17349,N_16725,N_16735);
nand U17350 (N_17350,N_16512,N_16865);
nand U17351 (N_17351,N_16681,N_16905);
nand U17352 (N_17352,N_16723,N_16782);
or U17353 (N_17353,N_16945,N_16607);
and U17354 (N_17354,N_16658,N_16602);
xor U17355 (N_17355,N_16587,N_16873);
and U17356 (N_17356,N_16831,N_16631);
nor U17357 (N_17357,N_16815,N_16673);
and U17358 (N_17358,N_16905,N_16840);
xor U17359 (N_17359,N_16591,N_16574);
and U17360 (N_17360,N_16998,N_16657);
xor U17361 (N_17361,N_16759,N_16904);
nor U17362 (N_17362,N_16539,N_16942);
nand U17363 (N_17363,N_16987,N_16934);
xnor U17364 (N_17364,N_16627,N_16847);
or U17365 (N_17365,N_16540,N_16564);
nand U17366 (N_17366,N_16788,N_16507);
xor U17367 (N_17367,N_16633,N_16687);
nor U17368 (N_17368,N_16915,N_16638);
or U17369 (N_17369,N_16631,N_16621);
or U17370 (N_17370,N_16711,N_16630);
or U17371 (N_17371,N_16946,N_16973);
nor U17372 (N_17372,N_16690,N_16822);
nor U17373 (N_17373,N_16827,N_16516);
xnor U17374 (N_17374,N_16762,N_16865);
nor U17375 (N_17375,N_16700,N_16821);
nand U17376 (N_17376,N_16734,N_16503);
and U17377 (N_17377,N_16927,N_16846);
or U17378 (N_17378,N_16785,N_16926);
or U17379 (N_17379,N_16788,N_16970);
nand U17380 (N_17380,N_16528,N_16993);
or U17381 (N_17381,N_16703,N_16550);
or U17382 (N_17382,N_16594,N_16672);
nor U17383 (N_17383,N_16742,N_16825);
nor U17384 (N_17384,N_16961,N_16911);
nor U17385 (N_17385,N_16678,N_16810);
xnor U17386 (N_17386,N_16560,N_16862);
nor U17387 (N_17387,N_16511,N_16541);
or U17388 (N_17388,N_16923,N_16786);
nor U17389 (N_17389,N_16933,N_16659);
nand U17390 (N_17390,N_16647,N_16640);
and U17391 (N_17391,N_16791,N_16656);
or U17392 (N_17392,N_16539,N_16616);
nor U17393 (N_17393,N_16975,N_16869);
or U17394 (N_17394,N_16700,N_16839);
xor U17395 (N_17395,N_16589,N_16956);
nand U17396 (N_17396,N_16562,N_16863);
nand U17397 (N_17397,N_16552,N_16586);
xor U17398 (N_17398,N_16895,N_16725);
or U17399 (N_17399,N_16601,N_16638);
xor U17400 (N_17400,N_16840,N_16545);
nor U17401 (N_17401,N_16571,N_16567);
xor U17402 (N_17402,N_16797,N_16867);
xor U17403 (N_17403,N_16828,N_16660);
nand U17404 (N_17404,N_16534,N_16942);
and U17405 (N_17405,N_16515,N_16524);
and U17406 (N_17406,N_16560,N_16722);
or U17407 (N_17407,N_16524,N_16666);
nand U17408 (N_17408,N_16512,N_16599);
and U17409 (N_17409,N_16515,N_16559);
or U17410 (N_17410,N_16961,N_16516);
xnor U17411 (N_17411,N_16895,N_16952);
nor U17412 (N_17412,N_16563,N_16946);
nor U17413 (N_17413,N_16987,N_16971);
xnor U17414 (N_17414,N_16727,N_16604);
xor U17415 (N_17415,N_16592,N_16761);
nand U17416 (N_17416,N_16956,N_16916);
nand U17417 (N_17417,N_16903,N_16879);
nand U17418 (N_17418,N_16553,N_16665);
nand U17419 (N_17419,N_16506,N_16774);
and U17420 (N_17420,N_16861,N_16792);
xnor U17421 (N_17421,N_16736,N_16515);
and U17422 (N_17422,N_16628,N_16550);
and U17423 (N_17423,N_16789,N_16745);
nand U17424 (N_17424,N_16732,N_16768);
or U17425 (N_17425,N_16625,N_16874);
and U17426 (N_17426,N_16855,N_16695);
xor U17427 (N_17427,N_16729,N_16607);
or U17428 (N_17428,N_16548,N_16651);
nand U17429 (N_17429,N_16813,N_16998);
or U17430 (N_17430,N_16817,N_16888);
nand U17431 (N_17431,N_16627,N_16619);
nand U17432 (N_17432,N_16661,N_16897);
or U17433 (N_17433,N_16966,N_16772);
nand U17434 (N_17434,N_16542,N_16928);
or U17435 (N_17435,N_16676,N_16671);
nor U17436 (N_17436,N_16520,N_16711);
xnor U17437 (N_17437,N_16626,N_16758);
and U17438 (N_17438,N_16559,N_16765);
and U17439 (N_17439,N_16845,N_16563);
or U17440 (N_17440,N_16918,N_16512);
or U17441 (N_17441,N_16922,N_16750);
nand U17442 (N_17442,N_16563,N_16882);
nor U17443 (N_17443,N_16867,N_16619);
or U17444 (N_17444,N_16547,N_16787);
nor U17445 (N_17445,N_16722,N_16878);
nor U17446 (N_17446,N_16809,N_16791);
nand U17447 (N_17447,N_16814,N_16806);
and U17448 (N_17448,N_16774,N_16532);
xor U17449 (N_17449,N_16892,N_16775);
nand U17450 (N_17450,N_16660,N_16727);
or U17451 (N_17451,N_16702,N_16835);
or U17452 (N_17452,N_16818,N_16730);
nor U17453 (N_17453,N_16944,N_16956);
nand U17454 (N_17454,N_16649,N_16526);
nor U17455 (N_17455,N_16566,N_16567);
nand U17456 (N_17456,N_16911,N_16580);
nor U17457 (N_17457,N_16735,N_16771);
xor U17458 (N_17458,N_16647,N_16802);
nand U17459 (N_17459,N_16567,N_16803);
nand U17460 (N_17460,N_16712,N_16503);
and U17461 (N_17461,N_16511,N_16834);
xnor U17462 (N_17462,N_16643,N_16642);
nor U17463 (N_17463,N_16971,N_16815);
and U17464 (N_17464,N_16845,N_16605);
nor U17465 (N_17465,N_16847,N_16858);
nand U17466 (N_17466,N_16557,N_16727);
or U17467 (N_17467,N_16736,N_16501);
nor U17468 (N_17468,N_16711,N_16894);
or U17469 (N_17469,N_16827,N_16546);
nand U17470 (N_17470,N_16704,N_16549);
and U17471 (N_17471,N_16769,N_16705);
nand U17472 (N_17472,N_16550,N_16781);
nor U17473 (N_17473,N_16707,N_16964);
nor U17474 (N_17474,N_16955,N_16743);
nor U17475 (N_17475,N_16714,N_16713);
and U17476 (N_17476,N_16945,N_16865);
or U17477 (N_17477,N_16699,N_16626);
or U17478 (N_17478,N_16803,N_16762);
xnor U17479 (N_17479,N_16782,N_16765);
nand U17480 (N_17480,N_16581,N_16818);
nand U17481 (N_17481,N_16607,N_16613);
or U17482 (N_17482,N_16568,N_16590);
xor U17483 (N_17483,N_16815,N_16993);
nand U17484 (N_17484,N_16654,N_16977);
xor U17485 (N_17485,N_16886,N_16508);
nor U17486 (N_17486,N_16723,N_16599);
nand U17487 (N_17487,N_16620,N_16549);
xor U17488 (N_17488,N_16543,N_16867);
nor U17489 (N_17489,N_16623,N_16956);
and U17490 (N_17490,N_16700,N_16719);
xor U17491 (N_17491,N_16779,N_16956);
xnor U17492 (N_17492,N_16652,N_16982);
xor U17493 (N_17493,N_16886,N_16733);
and U17494 (N_17494,N_16887,N_16611);
or U17495 (N_17495,N_16734,N_16641);
and U17496 (N_17496,N_16522,N_16702);
or U17497 (N_17497,N_16785,N_16656);
xor U17498 (N_17498,N_16516,N_16923);
nand U17499 (N_17499,N_16559,N_16716);
or U17500 (N_17500,N_17007,N_17439);
nand U17501 (N_17501,N_17183,N_17464);
nor U17502 (N_17502,N_17392,N_17247);
and U17503 (N_17503,N_17368,N_17362);
and U17504 (N_17504,N_17115,N_17395);
or U17505 (N_17505,N_17109,N_17371);
or U17506 (N_17506,N_17287,N_17129);
xor U17507 (N_17507,N_17022,N_17231);
nor U17508 (N_17508,N_17164,N_17270);
and U17509 (N_17509,N_17015,N_17035);
nand U17510 (N_17510,N_17289,N_17044);
nand U17511 (N_17511,N_17469,N_17322);
nand U17512 (N_17512,N_17112,N_17188);
nor U17513 (N_17513,N_17204,N_17203);
and U17514 (N_17514,N_17011,N_17190);
nor U17515 (N_17515,N_17485,N_17092);
and U17516 (N_17516,N_17209,N_17060);
nor U17517 (N_17517,N_17151,N_17423);
or U17518 (N_17518,N_17000,N_17202);
xor U17519 (N_17519,N_17279,N_17215);
nand U17520 (N_17520,N_17297,N_17354);
nand U17521 (N_17521,N_17402,N_17144);
or U17522 (N_17522,N_17388,N_17126);
nand U17523 (N_17523,N_17298,N_17207);
or U17524 (N_17524,N_17430,N_17259);
nor U17525 (N_17525,N_17266,N_17226);
nor U17526 (N_17526,N_17271,N_17108);
nor U17527 (N_17527,N_17017,N_17383);
nand U17528 (N_17528,N_17038,N_17021);
nor U17529 (N_17529,N_17356,N_17361);
nor U17530 (N_17530,N_17101,N_17481);
or U17531 (N_17531,N_17462,N_17104);
nor U17532 (N_17532,N_17331,N_17032);
nor U17533 (N_17533,N_17219,N_17014);
and U17534 (N_17534,N_17292,N_17347);
xnor U17535 (N_17535,N_17024,N_17065);
xnor U17536 (N_17536,N_17382,N_17278);
nand U17537 (N_17537,N_17489,N_17212);
or U17538 (N_17538,N_17053,N_17290);
xor U17539 (N_17539,N_17414,N_17317);
xnor U17540 (N_17540,N_17078,N_17432);
nand U17541 (N_17541,N_17338,N_17477);
nand U17542 (N_17542,N_17249,N_17142);
xor U17543 (N_17543,N_17156,N_17170);
or U17544 (N_17544,N_17380,N_17458);
and U17545 (N_17545,N_17146,N_17118);
or U17546 (N_17546,N_17025,N_17174);
and U17547 (N_17547,N_17265,N_17048);
or U17548 (N_17548,N_17302,N_17498);
xnor U17549 (N_17549,N_17268,N_17140);
nand U17550 (N_17550,N_17093,N_17213);
xor U17551 (N_17551,N_17475,N_17312);
xor U17552 (N_17552,N_17028,N_17367);
nor U17553 (N_17553,N_17348,N_17301);
nor U17554 (N_17554,N_17026,N_17411);
and U17555 (N_17555,N_17443,N_17206);
and U17556 (N_17556,N_17358,N_17150);
xor U17557 (N_17557,N_17124,N_17161);
nand U17558 (N_17558,N_17111,N_17133);
xor U17559 (N_17559,N_17341,N_17186);
nor U17560 (N_17560,N_17318,N_17479);
nand U17561 (N_17561,N_17130,N_17088);
xnor U17562 (N_17562,N_17470,N_17377);
xor U17563 (N_17563,N_17343,N_17474);
nand U17564 (N_17564,N_17490,N_17172);
xor U17565 (N_17565,N_17145,N_17393);
xnor U17566 (N_17566,N_17154,N_17454);
and U17567 (N_17567,N_17366,N_17099);
nor U17568 (N_17568,N_17461,N_17050);
or U17569 (N_17569,N_17373,N_17094);
nand U17570 (N_17570,N_17448,N_17196);
and U17571 (N_17571,N_17210,N_17019);
or U17572 (N_17572,N_17004,N_17193);
nand U17573 (N_17573,N_17275,N_17173);
xor U17574 (N_17574,N_17002,N_17023);
and U17575 (N_17575,N_17072,N_17391);
and U17576 (N_17576,N_17419,N_17030);
nor U17577 (N_17577,N_17143,N_17401);
or U17578 (N_17578,N_17057,N_17089);
and U17579 (N_17579,N_17321,N_17463);
or U17580 (N_17580,N_17037,N_17216);
or U17581 (N_17581,N_17169,N_17310);
or U17582 (N_17582,N_17267,N_17255);
or U17583 (N_17583,N_17230,N_17390);
and U17584 (N_17584,N_17486,N_17201);
nor U17585 (N_17585,N_17457,N_17328);
or U17586 (N_17586,N_17106,N_17309);
nand U17587 (N_17587,N_17323,N_17184);
nor U17588 (N_17588,N_17372,N_17234);
and U17589 (N_17589,N_17339,N_17125);
xnor U17590 (N_17590,N_17334,N_17293);
nor U17591 (N_17591,N_17082,N_17436);
or U17592 (N_17592,N_17191,N_17229);
or U17593 (N_17593,N_17333,N_17018);
nand U17594 (N_17594,N_17337,N_17425);
xnor U17595 (N_17595,N_17283,N_17049);
and U17596 (N_17596,N_17484,N_17379);
nor U17597 (N_17597,N_17246,N_17314);
or U17598 (N_17598,N_17488,N_17324);
nor U17599 (N_17599,N_17285,N_17385);
xnor U17600 (N_17600,N_17428,N_17256);
nand U17601 (N_17601,N_17059,N_17222);
nand U17602 (N_17602,N_17098,N_17420);
and U17603 (N_17603,N_17137,N_17149);
and U17604 (N_17604,N_17211,N_17325);
nor U17605 (N_17605,N_17272,N_17467);
xor U17606 (N_17606,N_17413,N_17459);
or U17607 (N_17607,N_17307,N_17465);
nor U17608 (N_17608,N_17426,N_17157);
or U17609 (N_17609,N_17499,N_17166);
or U17610 (N_17610,N_17442,N_17009);
xor U17611 (N_17611,N_17386,N_17406);
xnor U17612 (N_17612,N_17340,N_17178);
or U17613 (N_17613,N_17330,N_17336);
or U17614 (N_17614,N_17446,N_17300);
or U17615 (N_17615,N_17412,N_17497);
xor U17616 (N_17616,N_17223,N_17158);
xnor U17617 (N_17617,N_17295,N_17478);
nor U17618 (N_17618,N_17319,N_17352);
or U17619 (N_17619,N_17244,N_17122);
nand U17620 (N_17620,N_17036,N_17280);
and U17621 (N_17621,N_17253,N_17236);
and U17622 (N_17622,N_17311,N_17117);
or U17623 (N_17623,N_17068,N_17076);
nor U17624 (N_17624,N_17052,N_17153);
nor U17625 (N_17625,N_17085,N_17116);
or U17626 (N_17626,N_17080,N_17214);
xnor U17627 (N_17627,N_17006,N_17029);
and U17628 (N_17628,N_17062,N_17198);
xor U17629 (N_17629,N_17276,N_17357);
xnor U17630 (N_17630,N_17274,N_17148);
or U17631 (N_17631,N_17364,N_17043);
and U17632 (N_17632,N_17254,N_17303);
xor U17633 (N_17633,N_17107,N_17180);
or U17634 (N_17634,N_17189,N_17139);
and U17635 (N_17635,N_17453,N_17041);
xor U17636 (N_17636,N_17422,N_17431);
nand U17637 (N_17637,N_17286,N_17273);
and U17638 (N_17638,N_17480,N_17389);
or U17639 (N_17639,N_17194,N_17110);
nor U17640 (N_17640,N_17387,N_17447);
or U17641 (N_17641,N_17013,N_17429);
or U17642 (N_17642,N_17232,N_17208);
nand U17643 (N_17643,N_17167,N_17012);
nor U17644 (N_17644,N_17260,N_17353);
nor U17645 (N_17645,N_17128,N_17086);
xor U17646 (N_17646,N_17033,N_17056);
nor U17647 (N_17647,N_17248,N_17200);
or U17648 (N_17648,N_17218,N_17123);
xor U17649 (N_17649,N_17359,N_17163);
nand U17650 (N_17650,N_17398,N_17070);
and U17651 (N_17651,N_17308,N_17455);
nor U17652 (N_17652,N_17205,N_17228);
xnor U17653 (N_17653,N_17327,N_17363);
and U17654 (N_17654,N_17020,N_17042);
nand U17655 (N_17655,N_17472,N_17039);
nor U17656 (N_17656,N_17421,N_17135);
xor U17657 (N_17657,N_17103,N_17066);
and U17658 (N_17658,N_17171,N_17179);
and U17659 (N_17659,N_17090,N_17493);
nand U17660 (N_17660,N_17119,N_17055);
nand U17661 (N_17661,N_17160,N_17242);
xor U17662 (N_17662,N_17081,N_17181);
and U17663 (N_17663,N_17240,N_17299);
and U17664 (N_17664,N_17258,N_17010);
nor U17665 (N_17665,N_17394,N_17045);
nor U17666 (N_17666,N_17460,N_17054);
or U17667 (N_17667,N_17378,N_17305);
nor U17668 (N_17668,N_17400,N_17073);
and U17669 (N_17669,N_17491,N_17440);
nor U17670 (N_17670,N_17277,N_17496);
nand U17671 (N_17671,N_17438,N_17031);
or U17672 (N_17672,N_17427,N_17077);
nor U17673 (N_17673,N_17239,N_17482);
nor U17674 (N_17674,N_17165,N_17349);
and U17675 (N_17675,N_17224,N_17071);
nor U17676 (N_17676,N_17264,N_17445);
or U17677 (N_17677,N_17435,N_17177);
nand U17678 (N_17678,N_17233,N_17087);
or U17679 (N_17679,N_17155,N_17404);
and U17680 (N_17680,N_17063,N_17396);
nand U17681 (N_17681,N_17441,N_17105);
or U17682 (N_17682,N_17005,N_17175);
and U17683 (N_17683,N_17083,N_17345);
nand U17684 (N_17684,N_17064,N_17369);
nor U17685 (N_17685,N_17221,N_17091);
xor U17686 (N_17686,N_17433,N_17217);
or U17687 (N_17687,N_17408,N_17350);
or U17688 (N_17688,N_17261,N_17192);
or U17689 (N_17689,N_17437,N_17100);
nor U17690 (N_17690,N_17138,N_17113);
nor U17691 (N_17691,N_17027,N_17252);
nor U17692 (N_17692,N_17132,N_17147);
and U17693 (N_17693,N_17399,N_17306);
or U17694 (N_17694,N_17034,N_17296);
or U17695 (N_17695,N_17152,N_17416);
nand U17696 (N_17696,N_17096,N_17243);
or U17697 (N_17697,N_17058,N_17238);
and U17698 (N_17698,N_17409,N_17225);
xor U17699 (N_17699,N_17251,N_17374);
xor U17700 (N_17700,N_17492,N_17182);
or U17701 (N_17701,N_17079,N_17001);
nor U17702 (N_17702,N_17235,N_17284);
nand U17703 (N_17703,N_17227,N_17282);
nand U17704 (N_17704,N_17075,N_17185);
and U17705 (N_17705,N_17136,N_17141);
and U17706 (N_17706,N_17351,N_17120);
xnor U17707 (N_17707,N_17294,N_17487);
nand U17708 (N_17708,N_17262,N_17449);
nand U17709 (N_17709,N_17127,N_17121);
nand U17710 (N_17710,N_17046,N_17410);
or U17711 (N_17711,N_17291,N_17199);
or U17712 (N_17712,N_17370,N_17250);
nand U17713 (N_17713,N_17397,N_17407);
and U17714 (N_17714,N_17061,N_17102);
xnor U17715 (N_17715,N_17245,N_17365);
xnor U17716 (N_17716,N_17269,N_17040);
and U17717 (N_17717,N_17220,N_17051);
nand U17718 (N_17718,N_17003,N_17281);
and U17719 (N_17719,N_17424,N_17417);
or U17720 (N_17720,N_17195,N_17326);
nand U17721 (N_17721,N_17008,N_17335);
or U17722 (N_17722,N_17468,N_17329);
nor U17723 (N_17723,N_17315,N_17263);
nand U17724 (N_17724,N_17187,N_17176);
and U17725 (N_17725,N_17476,N_17434);
or U17726 (N_17726,N_17466,N_17483);
and U17727 (N_17727,N_17320,N_17168);
nand U17728 (N_17728,N_17355,N_17452);
nand U17729 (N_17729,N_17444,N_17313);
and U17730 (N_17730,N_17342,N_17403);
xor U17731 (N_17731,N_17381,N_17346);
or U17732 (N_17732,N_17494,N_17405);
xor U17733 (N_17733,N_17237,N_17074);
xor U17734 (N_17734,N_17495,N_17197);
nand U17735 (N_17735,N_17332,N_17450);
xnor U17736 (N_17736,N_17344,N_17418);
xor U17737 (N_17737,N_17376,N_17288);
nand U17738 (N_17738,N_17159,N_17375);
xnor U17739 (N_17739,N_17384,N_17097);
or U17740 (N_17740,N_17257,N_17456);
and U17741 (N_17741,N_17162,N_17304);
nor U17742 (N_17742,N_17095,N_17415);
xnor U17743 (N_17743,N_17316,N_17131);
nor U17744 (N_17744,N_17016,N_17451);
or U17745 (N_17745,N_17067,N_17047);
nor U17746 (N_17746,N_17134,N_17114);
nand U17747 (N_17747,N_17360,N_17084);
or U17748 (N_17748,N_17069,N_17473);
and U17749 (N_17749,N_17241,N_17471);
and U17750 (N_17750,N_17273,N_17108);
nor U17751 (N_17751,N_17465,N_17005);
xor U17752 (N_17752,N_17130,N_17432);
and U17753 (N_17753,N_17358,N_17386);
nand U17754 (N_17754,N_17386,N_17253);
nor U17755 (N_17755,N_17384,N_17006);
xnor U17756 (N_17756,N_17401,N_17307);
xnor U17757 (N_17757,N_17392,N_17480);
nand U17758 (N_17758,N_17378,N_17370);
xnor U17759 (N_17759,N_17135,N_17221);
and U17760 (N_17760,N_17006,N_17108);
nand U17761 (N_17761,N_17176,N_17052);
nor U17762 (N_17762,N_17395,N_17218);
nor U17763 (N_17763,N_17421,N_17399);
xnor U17764 (N_17764,N_17332,N_17146);
xnor U17765 (N_17765,N_17245,N_17016);
nand U17766 (N_17766,N_17084,N_17307);
nand U17767 (N_17767,N_17456,N_17436);
xnor U17768 (N_17768,N_17095,N_17067);
or U17769 (N_17769,N_17331,N_17047);
nor U17770 (N_17770,N_17454,N_17177);
xnor U17771 (N_17771,N_17065,N_17224);
and U17772 (N_17772,N_17171,N_17486);
nand U17773 (N_17773,N_17135,N_17271);
nor U17774 (N_17774,N_17198,N_17113);
nand U17775 (N_17775,N_17416,N_17196);
and U17776 (N_17776,N_17347,N_17323);
or U17777 (N_17777,N_17178,N_17418);
nand U17778 (N_17778,N_17092,N_17270);
nor U17779 (N_17779,N_17233,N_17120);
nor U17780 (N_17780,N_17417,N_17163);
xor U17781 (N_17781,N_17359,N_17125);
xnor U17782 (N_17782,N_17140,N_17131);
or U17783 (N_17783,N_17300,N_17487);
or U17784 (N_17784,N_17400,N_17101);
or U17785 (N_17785,N_17206,N_17438);
nand U17786 (N_17786,N_17147,N_17078);
nand U17787 (N_17787,N_17198,N_17057);
and U17788 (N_17788,N_17257,N_17334);
nor U17789 (N_17789,N_17060,N_17219);
nor U17790 (N_17790,N_17318,N_17271);
nor U17791 (N_17791,N_17220,N_17156);
nor U17792 (N_17792,N_17063,N_17308);
xnor U17793 (N_17793,N_17238,N_17128);
xor U17794 (N_17794,N_17342,N_17375);
xor U17795 (N_17795,N_17495,N_17159);
and U17796 (N_17796,N_17009,N_17127);
xor U17797 (N_17797,N_17399,N_17250);
nor U17798 (N_17798,N_17027,N_17403);
nand U17799 (N_17799,N_17397,N_17472);
nand U17800 (N_17800,N_17377,N_17220);
or U17801 (N_17801,N_17265,N_17151);
or U17802 (N_17802,N_17282,N_17073);
xnor U17803 (N_17803,N_17234,N_17474);
xnor U17804 (N_17804,N_17177,N_17038);
or U17805 (N_17805,N_17003,N_17131);
and U17806 (N_17806,N_17173,N_17494);
and U17807 (N_17807,N_17344,N_17044);
or U17808 (N_17808,N_17332,N_17031);
and U17809 (N_17809,N_17393,N_17146);
and U17810 (N_17810,N_17338,N_17143);
and U17811 (N_17811,N_17315,N_17074);
xor U17812 (N_17812,N_17442,N_17334);
and U17813 (N_17813,N_17433,N_17484);
nand U17814 (N_17814,N_17240,N_17028);
and U17815 (N_17815,N_17008,N_17423);
or U17816 (N_17816,N_17217,N_17031);
xor U17817 (N_17817,N_17316,N_17060);
nand U17818 (N_17818,N_17373,N_17277);
nor U17819 (N_17819,N_17468,N_17038);
nand U17820 (N_17820,N_17485,N_17052);
and U17821 (N_17821,N_17381,N_17011);
nor U17822 (N_17822,N_17332,N_17085);
nand U17823 (N_17823,N_17198,N_17454);
nor U17824 (N_17824,N_17100,N_17258);
nor U17825 (N_17825,N_17182,N_17272);
xor U17826 (N_17826,N_17247,N_17049);
or U17827 (N_17827,N_17139,N_17354);
and U17828 (N_17828,N_17347,N_17490);
nor U17829 (N_17829,N_17036,N_17158);
nor U17830 (N_17830,N_17286,N_17497);
or U17831 (N_17831,N_17160,N_17007);
nor U17832 (N_17832,N_17393,N_17258);
xnor U17833 (N_17833,N_17153,N_17443);
xor U17834 (N_17834,N_17168,N_17275);
nand U17835 (N_17835,N_17475,N_17163);
and U17836 (N_17836,N_17367,N_17035);
nor U17837 (N_17837,N_17252,N_17041);
nand U17838 (N_17838,N_17304,N_17003);
nor U17839 (N_17839,N_17186,N_17148);
xor U17840 (N_17840,N_17240,N_17144);
or U17841 (N_17841,N_17466,N_17173);
nand U17842 (N_17842,N_17145,N_17469);
nor U17843 (N_17843,N_17344,N_17458);
xnor U17844 (N_17844,N_17318,N_17127);
xor U17845 (N_17845,N_17331,N_17275);
nand U17846 (N_17846,N_17216,N_17010);
nand U17847 (N_17847,N_17004,N_17046);
nand U17848 (N_17848,N_17211,N_17446);
nand U17849 (N_17849,N_17108,N_17426);
or U17850 (N_17850,N_17443,N_17004);
and U17851 (N_17851,N_17302,N_17214);
nand U17852 (N_17852,N_17484,N_17409);
or U17853 (N_17853,N_17432,N_17047);
nand U17854 (N_17854,N_17415,N_17016);
nor U17855 (N_17855,N_17140,N_17397);
nand U17856 (N_17856,N_17168,N_17019);
and U17857 (N_17857,N_17313,N_17110);
xnor U17858 (N_17858,N_17275,N_17192);
nand U17859 (N_17859,N_17184,N_17473);
nand U17860 (N_17860,N_17482,N_17433);
and U17861 (N_17861,N_17062,N_17393);
and U17862 (N_17862,N_17020,N_17169);
nand U17863 (N_17863,N_17411,N_17328);
and U17864 (N_17864,N_17078,N_17061);
and U17865 (N_17865,N_17336,N_17127);
nand U17866 (N_17866,N_17437,N_17436);
and U17867 (N_17867,N_17114,N_17083);
and U17868 (N_17868,N_17312,N_17151);
xnor U17869 (N_17869,N_17322,N_17004);
nor U17870 (N_17870,N_17376,N_17403);
or U17871 (N_17871,N_17123,N_17263);
and U17872 (N_17872,N_17245,N_17203);
xor U17873 (N_17873,N_17387,N_17265);
nand U17874 (N_17874,N_17218,N_17246);
or U17875 (N_17875,N_17141,N_17228);
and U17876 (N_17876,N_17077,N_17230);
or U17877 (N_17877,N_17043,N_17203);
xor U17878 (N_17878,N_17425,N_17044);
nand U17879 (N_17879,N_17236,N_17121);
or U17880 (N_17880,N_17348,N_17479);
xor U17881 (N_17881,N_17396,N_17410);
xnor U17882 (N_17882,N_17455,N_17468);
and U17883 (N_17883,N_17169,N_17367);
nor U17884 (N_17884,N_17447,N_17464);
or U17885 (N_17885,N_17337,N_17122);
nand U17886 (N_17886,N_17483,N_17173);
and U17887 (N_17887,N_17105,N_17303);
and U17888 (N_17888,N_17290,N_17275);
nor U17889 (N_17889,N_17331,N_17163);
xor U17890 (N_17890,N_17194,N_17322);
and U17891 (N_17891,N_17332,N_17206);
xnor U17892 (N_17892,N_17091,N_17171);
and U17893 (N_17893,N_17336,N_17308);
nor U17894 (N_17894,N_17001,N_17227);
and U17895 (N_17895,N_17488,N_17382);
nand U17896 (N_17896,N_17458,N_17435);
nand U17897 (N_17897,N_17434,N_17234);
and U17898 (N_17898,N_17101,N_17388);
nand U17899 (N_17899,N_17333,N_17476);
xnor U17900 (N_17900,N_17336,N_17019);
or U17901 (N_17901,N_17189,N_17095);
nand U17902 (N_17902,N_17207,N_17436);
xor U17903 (N_17903,N_17041,N_17155);
and U17904 (N_17904,N_17470,N_17068);
nand U17905 (N_17905,N_17140,N_17433);
or U17906 (N_17906,N_17056,N_17173);
or U17907 (N_17907,N_17278,N_17283);
nand U17908 (N_17908,N_17496,N_17490);
nor U17909 (N_17909,N_17373,N_17405);
or U17910 (N_17910,N_17490,N_17061);
nand U17911 (N_17911,N_17380,N_17412);
nand U17912 (N_17912,N_17264,N_17381);
or U17913 (N_17913,N_17155,N_17495);
nand U17914 (N_17914,N_17478,N_17489);
or U17915 (N_17915,N_17229,N_17378);
and U17916 (N_17916,N_17046,N_17471);
and U17917 (N_17917,N_17173,N_17329);
nand U17918 (N_17918,N_17363,N_17328);
xnor U17919 (N_17919,N_17386,N_17202);
nand U17920 (N_17920,N_17497,N_17396);
xor U17921 (N_17921,N_17293,N_17269);
and U17922 (N_17922,N_17276,N_17306);
and U17923 (N_17923,N_17158,N_17375);
nand U17924 (N_17924,N_17094,N_17483);
xor U17925 (N_17925,N_17029,N_17454);
nand U17926 (N_17926,N_17260,N_17372);
nand U17927 (N_17927,N_17254,N_17181);
xor U17928 (N_17928,N_17384,N_17320);
xnor U17929 (N_17929,N_17067,N_17023);
and U17930 (N_17930,N_17351,N_17216);
and U17931 (N_17931,N_17461,N_17049);
nand U17932 (N_17932,N_17245,N_17085);
nor U17933 (N_17933,N_17052,N_17210);
nand U17934 (N_17934,N_17052,N_17457);
or U17935 (N_17935,N_17137,N_17232);
and U17936 (N_17936,N_17379,N_17463);
nor U17937 (N_17937,N_17055,N_17113);
nand U17938 (N_17938,N_17172,N_17457);
xor U17939 (N_17939,N_17188,N_17307);
nor U17940 (N_17940,N_17462,N_17420);
or U17941 (N_17941,N_17015,N_17406);
nand U17942 (N_17942,N_17369,N_17258);
and U17943 (N_17943,N_17194,N_17125);
nor U17944 (N_17944,N_17408,N_17188);
xor U17945 (N_17945,N_17276,N_17210);
nand U17946 (N_17946,N_17399,N_17205);
and U17947 (N_17947,N_17055,N_17034);
nand U17948 (N_17948,N_17429,N_17034);
nor U17949 (N_17949,N_17112,N_17255);
and U17950 (N_17950,N_17320,N_17306);
and U17951 (N_17951,N_17318,N_17315);
nand U17952 (N_17952,N_17084,N_17349);
and U17953 (N_17953,N_17477,N_17418);
and U17954 (N_17954,N_17388,N_17395);
nand U17955 (N_17955,N_17408,N_17177);
xor U17956 (N_17956,N_17040,N_17076);
nor U17957 (N_17957,N_17143,N_17013);
nand U17958 (N_17958,N_17104,N_17401);
nor U17959 (N_17959,N_17142,N_17091);
and U17960 (N_17960,N_17438,N_17445);
nand U17961 (N_17961,N_17283,N_17111);
or U17962 (N_17962,N_17154,N_17319);
xnor U17963 (N_17963,N_17335,N_17281);
nor U17964 (N_17964,N_17263,N_17023);
xor U17965 (N_17965,N_17204,N_17407);
xnor U17966 (N_17966,N_17132,N_17042);
xnor U17967 (N_17967,N_17455,N_17369);
xor U17968 (N_17968,N_17148,N_17023);
nor U17969 (N_17969,N_17061,N_17443);
nor U17970 (N_17970,N_17012,N_17255);
or U17971 (N_17971,N_17444,N_17388);
xor U17972 (N_17972,N_17303,N_17251);
or U17973 (N_17973,N_17271,N_17103);
xor U17974 (N_17974,N_17294,N_17467);
or U17975 (N_17975,N_17081,N_17084);
nor U17976 (N_17976,N_17401,N_17013);
nor U17977 (N_17977,N_17325,N_17179);
and U17978 (N_17978,N_17120,N_17392);
xor U17979 (N_17979,N_17308,N_17372);
and U17980 (N_17980,N_17328,N_17312);
xnor U17981 (N_17981,N_17386,N_17283);
nand U17982 (N_17982,N_17327,N_17235);
and U17983 (N_17983,N_17275,N_17439);
or U17984 (N_17984,N_17313,N_17226);
nor U17985 (N_17985,N_17248,N_17196);
or U17986 (N_17986,N_17427,N_17358);
and U17987 (N_17987,N_17358,N_17115);
and U17988 (N_17988,N_17205,N_17030);
and U17989 (N_17989,N_17190,N_17391);
nand U17990 (N_17990,N_17247,N_17072);
and U17991 (N_17991,N_17029,N_17188);
or U17992 (N_17992,N_17480,N_17004);
or U17993 (N_17993,N_17338,N_17497);
nor U17994 (N_17994,N_17246,N_17041);
or U17995 (N_17995,N_17332,N_17472);
and U17996 (N_17996,N_17197,N_17133);
xor U17997 (N_17997,N_17183,N_17375);
xnor U17998 (N_17998,N_17380,N_17173);
nor U17999 (N_17999,N_17262,N_17136);
or U18000 (N_18000,N_17966,N_17612);
and U18001 (N_18001,N_17733,N_17639);
or U18002 (N_18002,N_17556,N_17978);
nand U18003 (N_18003,N_17632,N_17601);
or U18004 (N_18004,N_17805,N_17864);
and U18005 (N_18005,N_17546,N_17767);
nand U18006 (N_18006,N_17960,N_17976);
nor U18007 (N_18007,N_17653,N_17509);
or U18008 (N_18008,N_17929,N_17902);
or U18009 (N_18009,N_17814,N_17687);
nand U18010 (N_18010,N_17967,N_17825);
nor U18011 (N_18011,N_17849,N_17598);
and U18012 (N_18012,N_17840,N_17554);
and U18013 (N_18013,N_17842,N_17587);
nor U18014 (N_18014,N_17510,N_17874);
or U18015 (N_18015,N_17924,N_17547);
xnor U18016 (N_18016,N_17827,N_17775);
nor U18017 (N_18017,N_17685,N_17530);
nand U18018 (N_18018,N_17717,N_17736);
nor U18019 (N_18019,N_17906,N_17590);
or U18020 (N_18020,N_17517,N_17972);
xor U18021 (N_18021,N_17720,N_17742);
nor U18022 (N_18022,N_17732,N_17529);
xor U18023 (N_18023,N_17769,N_17996);
and U18024 (N_18024,N_17748,N_17868);
nor U18025 (N_18025,N_17950,N_17689);
xor U18026 (N_18026,N_17974,N_17946);
xnor U18027 (N_18027,N_17543,N_17971);
nor U18028 (N_18028,N_17558,N_17887);
nand U18029 (N_18029,N_17765,N_17995);
nor U18030 (N_18030,N_17502,N_17956);
nand U18031 (N_18031,N_17658,N_17931);
nor U18032 (N_18032,N_17968,N_17566);
or U18033 (N_18033,N_17700,N_17757);
and U18034 (N_18034,N_17561,N_17584);
nor U18035 (N_18035,N_17774,N_17883);
xor U18036 (N_18036,N_17731,N_17707);
and U18037 (N_18037,N_17730,N_17711);
or U18038 (N_18038,N_17522,N_17672);
nor U18039 (N_18039,N_17988,N_17993);
xor U18040 (N_18040,N_17633,N_17740);
or U18041 (N_18041,N_17698,N_17831);
xor U18042 (N_18042,N_17679,N_17872);
nand U18043 (N_18043,N_17702,N_17713);
xnor U18044 (N_18044,N_17613,N_17766);
or U18045 (N_18045,N_17819,N_17808);
nand U18046 (N_18046,N_17750,N_17693);
or U18047 (N_18047,N_17991,N_17662);
or U18048 (N_18048,N_17563,N_17620);
nor U18049 (N_18049,N_17667,N_17777);
and U18050 (N_18050,N_17668,N_17745);
or U18051 (N_18051,N_17705,N_17594);
and U18052 (N_18052,N_17673,N_17512);
or U18053 (N_18053,N_17837,N_17596);
or U18054 (N_18054,N_17920,N_17696);
and U18055 (N_18055,N_17643,N_17803);
xnor U18056 (N_18056,N_17895,N_17782);
and U18057 (N_18057,N_17884,N_17790);
xor U18058 (N_18058,N_17744,N_17869);
nand U18059 (N_18059,N_17627,N_17604);
nand U18060 (N_18060,N_17888,N_17801);
xor U18061 (N_18061,N_17918,N_17875);
nand U18062 (N_18062,N_17629,N_17877);
or U18063 (N_18063,N_17710,N_17800);
nor U18064 (N_18064,N_17553,N_17861);
xor U18065 (N_18065,N_17990,N_17893);
nor U18066 (N_18066,N_17822,N_17795);
nor U18067 (N_18067,N_17749,N_17504);
and U18068 (N_18068,N_17751,N_17835);
nor U18069 (N_18069,N_17674,N_17501);
nor U18070 (N_18070,N_17885,N_17951);
and U18071 (N_18071,N_17536,N_17614);
xnor U18072 (N_18072,N_17778,N_17694);
nand U18073 (N_18073,N_17826,N_17818);
or U18074 (N_18074,N_17834,N_17845);
xnor U18075 (N_18075,N_17855,N_17592);
or U18076 (N_18076,N_17706,N_17508);
nor U18077 (N_18077,N_17666,N_17903);
or U18078 (N_18078,N_17626,N_17630);
and U18079 (N_18079,N_17937,N_17534);
xor U18080 (N_18080,N_17779,N_17727);
nor U18081 (N_18081,N_17984,N_17813);
or U18082 (N_18082,N_17880,N_17661);
nor U18083 (N_18083,N_17898,N_17608);
nand U18084 (N_18084,N_17934,N_17911);
xor U18085 (N_18085,N_17870,N_17645);
xor U18086 (N_18086,N_17891,N_17642);
xor U18087 (N_18087,N_17505,N_17725);
nand U18088 (N_18088,N_17539,N_17853);
and U18089 (N_18089,N_17680,N_17616);
and U18090 (N_18090,N_17586,N_17654);
and U18091 (N_18091,N_17958,N_17682);
or U18092 (N_18092,N_17677,N_17992);
and U18093 (N_18093,N_17724,N_17722);
and U18094 (N_18094,N_17938,N_17901);
nand U18095 (N_18095,N_17862,N_17595);
nor U18096 (N_18096,N_17635,N_17761);
or U18097 (N_18097,N_17921,N_17823);
or U18098 (N_18098,N_17860,N_17985);
nand U18099 (N_18099,N_17816,N_17737);
xnor U18100 (N_18100,N_17876,N_17847);
xor U18101 (N_18101,N_17686,N_17802);
nor U18102 (N_18102,N_17909,N_17760);
nand U18103 (N_18103,N_17764,N_17809);
nor U18104 (N_18104,N_17575,N_17610);
nand U18105 (N_18105,N_17570,N_17507);
or U18106 (N_18106,N_17537,N_17832);
and U18107 (N_18107,N_17549,N_17548);
or U18108 (N_18108,N_17759,N_17973);
xnor U18109 (N_18109,N_17591,N_17515);
nand U18110 (N_18110,N_17640,N_17589);
and U18111 (N_18111,N_17784,N_17599);
and U18112 (N_18112,N_17828,N_17754);
or U18113 (N_18113,N_17681,N_17573);
or U18114 (N_18114,N_17544,N_17848);
or U18115 (N_18115,N_17657,N_17899);
and U18116 (N_18116,N_17799,N_17542);
xor U18117 (N_18117,N_17856,N_17572);
nand U18118 (N_18118,N_17969,N_17678);
nand U18119 (N_18119,N_17794,N_17602);
and U18120 (N_18120,N_17622,N_17583);
and U18121 (N_18121,N_17904,N_17793);
nor U18122 (N_18122,N_17588,N_17569);
nand U18123 (N_18123,N_17838,N_17792);
nand U18124 (N_18124,N_17982,N_17511);
nor U18125 (N_18125,N_17965,N_17611);
or U18126 (N_18126,N_17551,N_17735);
and U18127 (N_18127,N_17810,N_17701);
nand U18128 (N_18128,N_17987,N_17528);
xnor U18129 (N_18129,N_17843,N_17562);
nand U18130 (N_18130,N_17624,N_17663);
and U18131 (N_18131,N_17646,N_17647);
and U18132 (N_18132,N_17697,N_17664);
or U18133 (N_18133,N_17912,N_17747);
and U18134 (N_18134,N_17723,N_17896);
xnor U18135 (N_18135,N_17936,N_17928);
nand U18136 (N_18136,N_17684,N_17550);
xnor U18137 (N_18137,N_17821,N_17582);
xor U18138 (N_18138,N_17752,N_17671);
xnor U18139 (N_18139,N_17941,N_17879);
and U18140 (N_18140,N_17715,N_17649);
nand U18141 (N_18141,N_17783,N_17948);
xnor U18142 (N_18142,N_17836,N_17797);
nand U18143 (N_18143,N_17866,N_17979);
and U18144 (N_18144,N_17669,N_17631);
nor U18145 (N_18145,N_17520,N_17621);
nor U18146 (N_18146,N_17789,N_17786);
nand U18147 (N_18147,N_17726,N_17863);
xor U18148 (N_18148,N_17516,N_17655);
nand U18149 (N_18149,N_17756,N_17665);
nor U18150 (N_18150,N_17567,N_17578);
and U18151 (N_18151,N_17980,N_17581);
nand U18152 (N_18152,N_17540,N_17670);
nor U18153 (N_18153,N_17758,N_17961);
and U18154 (N_18154,N_17704,N_17683);
xor U18155 (N_18155,N_17850,N_17609);
and U18156 (N_18156,N_17557,N_17699);
and U18157 (N_18157,N_17606,N_17709);
and U18158 (N_18158,N_17975,N_17503);
or U18159 (N_18159,N_17989,N_17852);
nand U18160 (N_18160,N_17952,N_17933);
xor U18161 (N_18161,N_17882,N_17617);
or U18162 (N_18162,N_17953,N_17734);
and U18163 (N_18163,N_17518,N_17648);
nor U18164 (N_18164,N_17533,N_17957);
xnor U18165 (N_18165,N_17935,N_17807);
nand U18166 (N_18166,N_17812,N_17641);
and U18167 (N_18167,N_17771,N_17675);
nor U18168 (N_18168,N_17762,N_17708);
xnor U18169 (N_18169,N_17506,N_17743);
nor U18170 (N_18170,N_17787,N_17527);
nand U18171 (N_18171,N_17538,N_17983);
and U18172 (N_18172,N_17927,N_17897);
and U18173 (N_18173,N_17636,N_17603);
nand U18174 (N_18174,N_17628,N_17576);
or U18175 (N_18175,N_17500,N_17728);
and U18176 (N_18176,N_17889,N_17867);
nand U18177 (N_18177,N_17521,N_17788);
or U18178 (N_18178,N_17577,N_17650);
nor U18179 (N_18179,N_17986,N_17955);
xor U18180 (N_18180,N_17833,N_17525);
or U18181 (N_18181,N_17524,N_17605);
and U18182 (N_18182,N_17922,N_17691);
nor U18183 (N_18183,N_17585,N_17970);
nand U18184 (N_18184,N_17894,N_17829);
or U18185 (N_18185,N_17712,N_17555);
nand U18186 (N_18186,N_17820,N_17651);
nand U18187 (N_18187,N_17824,N_17768);
and U18188 (N_18188,N_17804,N_17580);
nor U18189 (N_18189,N_17579,N_17781);
nand U18190 (N_18190,N_17519,N_17905);
nor U18191 (N_18191,N_17890,N_17716);
nand U18192 (N_18192,N_17858,N_17859);
or U18193 (N_18193,N_17571,N_17660);
xor U18194 (N_18194,N_17981,N_17703);
nor U18195 (N_18195,N_17977,N_17531);
or U18196 (N_18196,N_17552,N_17692);
nor U18197 (N_18197,N_17634,N_17846);
or U18198 (N_18198,N_17773,N_17690);
or U18199 (N_18199,N_17830,N_17913);
xor U18200 (N_18200,N_17564,N_17695);
and U18201 (N_18201,N_17526,N_17560);
and U18202 (N_18202,N_17910,N_17718);
xor U18203 (N_18203,N_17676,N_17900);
xor U18204 (N_18204,N_17593,N_17939);
or U18205 (N_18205,N_17776,N_17963);
or U18206 (N_18206,N_17932,N_17780);
nor U18207 (N_18207,N_17513,N_17959);
and U18208 (N_18208,N_17944,N_17607);
nor U18209 (N_18209,N_17619,N_17659);
or U18210 (N_18210,N_17656,N_17817);
nor U18211 (N_18211,N_17839,N_17719);
xor U18212 (N_18212,N_17844,N_17615);
nor U18213 (N_18213,N_17772,N_17878);
xor U18214 (N_18214,N_17623,N_17541);
nor U18215 (N_18215,N_17994,N_17997);
nand U18216 (N_18216,N_17791,N_17926);
nor U18217 (N_18217,N_17942,N_17798);
nand U18218 (N_18218,N_17597,N_17916);
and U18219 (N_18219,N_17871,N_17600);
xnor U18220 (N_18220,N_17714,N_17741);
nor U18221 (N_18221,N_17943,N_17892);
xnor U18222 (N_18222,N_17947,N_17999);
xor U18223 (N_18223,N_17907,N_17865);
or U18224 (N_18224,N_17914,N_17873);
xor U18225 (N_18225,N_17915,N_17739);
xnor U18226 (N_18226,N_17755,N_17886);
and U18227 (N_18227,N_17746,N_17753);
nor U18228 (N_18228,N_17919,N_17688);
xor U18229 (N_18229,N_17908,N_17523);
and U18230 (N_18230,N_17559,N_17565);
xnor U18231 (N_18231,N_17729,N_17763);
xnor U18232 (N_18232,N_17954,N_17940);
nor U18233 (N_18233,N_17881,N_17535);
xor U18234 (N_18234,N_17738,N_17917);
and U18235 (N_18235,N_17841,N_17574);
and U18236 (N_18236,N_17532,N_17625);
nand U18237 (N_18237,N_17964,N_17806);
xnor U18238 (N_18238,N_17998,N_17638);
and U18239 (N_18239,N_17545,N_17637);
xor U18240 (N_18240,N_17854,N_17568);
and U18241 (N_18241,N_17945,N_17925);
or U18242 (N_18242,N_17514,N_17770);
and U18243 (N_18243,N_17811,N_17815);
or U18244 (N_18244,N_17857,N_17785);
nand U18245 (N_18245,N_17949,N_17618);
nor U18246 (N_18246,N_17930,N_17962);
xor U18247 (N_18247,N_17721,N_17851);
and U18248 (N_18248,N_17796,N_17923);
nand U18249 (N_18249,N_17652,N_17644);
nor U18250 (N_18250,N_17809,N_17836);
xnor U18251 (N_18251,N_17505,N_17904);
and U18252 (N_18252,N_17925,N_17740);
or U18253 (N_18253,N_17798,N_17773);
nand U18254 (N_18254,N_17917,N_17977);
or U18255 (N_18255,N_17790,N_17561);
nor U18256 (N_18256,N_17922,N_17644);
nand U18257 (N_18257,N_17866,N_17795);
xor U18258 (N_18258,N_17646,N_17529);
and U18259 (N_18259,N_17865,N_17963);
nand U18260 (N_18260,N_17981,N_17701);
or U18261 (N_18261,N_17650,N_17647);
or U18262 (N_18262,N_17521,N_17796);
nor U18263 (N_18263,N_17836,N_17667);
and U18264 (N_18264,N_17951,N_17809);
or U18265 (N_18265,N_17717,N_17748);
and U18266 (N_18266,N_17569,N_17814);
and U18267 (N_18267,N_17960,N_17533);
or U18268 (N_18268,N_17787,N_17669);
xor U18269 (N_18269,N_17646,N_17771);
or U18270 (N_18270,N_17644,N_17703);
nand U18271 (N_18271,N_17629,N_17541);
xor U18272 (N_18272,N_17554,N_17921);
and U18273 (N_18273,N_17815,N_17887);
xor U18274 (N_18274,N_17704,N_17809);
nor U18275 (N_18275,N_17701,N_17595);
or U18276 (N_18276,N_17891,N_17797);
and U18277 (N_18277,N_17982,N_17650);
or U18278 (N_18278,N_17945,N_17703);
nor U18279 (N_18279,N_17982,N_17556);
or U18280 (N_18280,N_17555,N_17612);
xor U18281 (N_18281,N_17684,N_17725);
nand U18282 (N_18282,N_17793,N_17918);
nor U18283 (N_18283,N_17723,N_17583);
or U18284 (N_18284,N_17562,N_17910);
or U18285 (N_18285,N_17668,N_17808);
and U18286 (N_18286,N_17805,N_17612);
nand U18287 (N_18287,N_17842,N_17678);
nand U18288 (N_18288,N_17855,N_17739);
xnor U18289 (N_18289,N_17645,N_17975);
xnor U18290 (N_18290,N_17987,N_17711);
or U18291 (N_18291,N_17729,N_17616);
xnor U18292 (N_18292,N_17748,N_17631);
xor U18293 (N_18293,N_17627,N_17811);
nand U18294 (N_18294,N_17557,N_17801);
and U18295 (N_18295,N_17530,N_17600);
and U18296 (N_18296,N_17702,N_17764);
nand U18297 (N_18297,N_17988,N_17789);
and U18298 (N_18298,N_17757,N_17848);
and U18299 (N_18299,N_17579,N_17703);
or U18300 (N_18300,N_17871,N_17619);
xnor U18301 (N_18301,N_17666,N_17597);
nand U18302 (N_18302,N_17939,N_17879);
nand U18303 (N_18303,N_17508,N_17902);
or U18304 (N_18304,N_17677,N_17869);
or U18305 (N_18305,N_17976,N_17798);
xnor U18306 (N_18306,N_17980,N_17618);
xor U18307 (N_18307,N_17815,N_17950);
nand U18308 (N_18308,N_17928,N_17817);
nand U18309 (N_18309,N_17770,N_17638);
and U18310 (N_18310,N_17521,N_17969);
and U18311 (N_18311,N_17567,N_17651);
or U18312 (N_18312,N_17856,N_17823);
nor U18313 (N_18313,N_17976,N_17965);
xnor U18314 (N_18314,N_17836,N_17581);
or U18315 (N_18315,N_17501,N_17556);
and U18316 (N_18316,N_17956,N_17854);
nor U18317 (N_18317,N_17740,N_17526);
or U18318 (N_18318,N_17521,N_17810);
xnor U18319 (N_18319,N_17595,N_17597);
nand U18320 (N_18320,N_17670,N_17662);
xnor U18321 (N_18321,N_17520,N_17609);
and U18322 (N_18322,N_17703,N_17728);
nand U18323 (N_18323,N_17786,N_17741);
nor U18324 (N_18324,N_17910,N_17657);
nand U18325 (N_18325,N_17755,N_17943);
xnor U18326 (N_18326,N_17673,N_17598);
or U18327 (N_18327,N_17633,N_17629);
or U18328 (N_18328,N_17903,N_17668);
and U18329 (N_18329,N_17523,N_17800);
nand U18330 (N_18330,N_17504,N_17703);
or U18331 (N_18331,N_17881,N_17864);
nand U18332 (N_18332,N_17916,N_17906);
nand U18333 (N_18333,N_17647,N_17758);
and U18334 (N_18334,N_17983,N_17736);
nor U18335 (N_18335,N_17629,N_17765);
nor U18336 (N_18336,N_17569,N_17942);
nor U18337 (N_18337,N_17786,N_17994);
nand U18338 (N_18338,N_17929,N_17595);
xor U18339 (N_18339,N_17821,N_17827);
nor U18340 (N_18340,N_17534,N_17912);
nor U18341 (N_18341,N_17582,N_17847);
xor U18342 (N_18342,N_17936,N_17714);
xor U18343 (N_18343,N_17667,N_17587);
or U18344 (N_18344,N_17946,N_17735);
nor U18345 (N_18345,N_17674,N_17506);
nand U18346 (N_18346,N_17534,N_17948);
or U18347 (N_18347,N_17947,N_17797);
and U18348 (N_18348,N_17657,N_17642);
nand U18349 (N_18349,N_17651,N_17726);
and U18350 (N_18350,N_17720,N_17708);
and U18351 (N_18351,N_17632,N_17587);
nor U18352 (N_18352,N_17606,N_17902);
xor U18353 (N_18353,N_17888,N_17602);
nor U18354 (N_18354,N_17817,N_17861);
and U18355 (N_18355,N_17584,N_17810);
or U18356 (N_18356,N_17563,N_17725);
xnor U18357 (N_18357,N_17647,N_17885);
nand U18358 (N_18358,N_17595,N_17980);
nand U18359 (N_18359,N_17648,N_17900);
and U18360 (N_18360,N_17732,N_17769);
or U18361 (N_18361,N_17699,N_17502);
and U18362 (N_18362,N_17908,N_17610);
xnor U18363 (N_18363,N_17566,N_17870);
or U18364 (N_18364,N_17996,N_17663);
and U18365 (N_18365,N_17769,N_17552);
and U18366 (N_18366,N_17958,N_17867);
or U18367 (N_18367,N_17595,N_17802);
and U18368 (N_18368,N_17717,N_17540);
nand U18369 (N_18369,N_17801,N_17645);
or U18370 (N_18370,N_17706,N_17532);
and U18371 (N_18371,N_17637,N_17910);
nor U18372 (N_18372,N_17796,N_17501);
xor U18373 (N_18373,N_17677,N_17731);
xnor U18374 (N_18374,N_17764,N_17590);
nand U18375 (N_18375,N_17706,N_17885);
xor U18376 (N_18376,N_17827,N_17974);
and U18377 (N_18377,N_17660,N_17646);
nor U18378 (N_18378,N_17786,N_17973);
nand U18379 (N_18379,N_17723,N_17647);
xor U18380 (N_18380,N_17639,N_17774);
nand U18381 (N_18381,N_17978,N_17960);
nand U18382 (N_18382,N_17906,N_17731);
nand U18383 (N_18383,N_17564,N_17525);
or U18384 (N_18384,N_17658,N_17616);
or U18385 (N_18385,N_17530,N_17981);
and U18386 (N_18386,N_17548,N_17993);
xnor U18387 (N_18387,N_17594,N_17532);
or U18388 (N_18388,N_17741,N_17522);
xnor U18389 (N_18389,N_17751,N_17631);
nand U18390 (N_18390,N_17781,N_17670);
or U18391 (N_18391,N_17656,N_17852);
nand U18392 (N_18392,N_17818,N_17586);
nand U18393 (N_18393,N_17854,N_17629);
or U18394 (N_18394,N_17873,N_17743);
and U18395 (N_18395,N_17674,N_17967);
nor U18396 (N_18396,N_17999,N_17589);
or U18397 (N_18397,N_17525,N_17874);
nor U18398 (N_18398,N_17798,N_17591);
xor U18399 (N_18399,N_17649,N_17691);
xor U18400 (N_18400,N_17587,N_17871);
nor U18401 (N_18401,N_17962,N_17892);
nand U18402 (N_18402,N_17782,N_17980);
xnor U18403 (N_18403,N_17810,N_17631);
or U18404 (N_18404,N_17511,N_17665);
nand U18405 (N_18405,N_17717,N_17902);
xnor U18406 (N_18406,N_17584,N_17588);
and U18407 (N_18407,N_17654,N_17863);
and U18408 (N_18408,N_17541,N_17720);
or U18409 (N_18409,N_17630,N_17820);
and U18410 (N_18410,N_17552,N_17932);
nor U18411 (N_18411,N_17768,N_17558);
xnor U18412 (N_18412,N_17693,N_17955);
or U18413 (N_18413,N_17809,N_17612);
or U18414 (N_18414,N_17766,N_17770);
nor U18415 (N_18415,N_17910,N_17706);
and U18416 (N_18416,N_17756,N_17956);
or U18417 (N_18417,N_17744,N_17639);
nor U18418 (N_18418,N_17850,N_17733);
or U18419 (N_18419,N_17674,N_17561);
nor U18420 (N_18420,N_17978,N_17782);
or U18421 (N_18421,N_17548,N_17838);
xnor U18422 (N_18422,N_17995,N_17662);
and U18423 (N_18423,N_17565,N_17502);
and U18424 (N_18424,N_17756,N_17684);
and U18425 (N_18425,N_17628,N_17654);
and U18426 (N_18426,N_17991,N_17769);
nor U18427 (N_18427,N_17768,N_17779);
nand U18428 (N_18428,N_17713,N_17763);
and U18429 (N_18429,N_17769,N_17975);
nor U18430 (N_18430,N_17669,N_17749);
nand U18431 (N_18431,N_17840,N_17563);
and U18432 (N_18432,N_17860,N_17688);
nor U18433 (N_18433,N_17610,N_17561);
nand U18434 (N_18434,N_17671,N_17707);
or U18435 (N_18435,N_17609,N_17848);
or U18436 (N_18436,N_17853,N_17541);
nor U18437 (N_18437,N_17893,N_17859);
nand U18438 (N_18438,N_17776,N_17667);
and U18439 (N_18439,N_17921,N_17895);
or U18440 (N_18440,N_17903,N_17907);
nor U18441 (N_18441,N_17973,N_17572);
nor U18442 (N_18442,N_17536,N_17613);
or U18443 (N_18443,N_17816,N_17752);
xor U18444 (N_18444,N_17501,N_17707);
nand U18445 (N_18445,N_17662,N_17926);
or U18446 (N_18446,N_17635,N_17956);
nor U18447 (N_18447,N_17992,N_17629);
xnor U18448 (N_18448,N_17771,N_17812);
nor U18449 (N_18449,N_17940,N_17930);
xor U18450 (N_18450,N_17913,N_17540);
xor U18451 (N_18451,N_17906,N_17681);
xnor U18452 (N_18452,N_17799,N_17895);
xnor U18453 (N_18453,N_17715,N_17605);
nand U18454 (N_18454,N_17684,N_17976);
and U18455 (N_18455,N_17658,N_17601);
nand U18456 (N_18456,N_17831,N_17815);
xor U18457 (N_18457,N_17947,N_17940);
xnor U18458 (N_18458,N_17902,N_17937);
xor U18459 (N_18459,N_17651,N_17725);
or U18460 (N_18460,N_17810,N_17956);
nand U18461 (N_18461,N_17702,N_17604);
nand U18462 (N_18462,N_17819,N_17992);
xor U18463 (N_18463,N_17603,N_17661);
or U18464 (N_18464,N_17995,N_17642);
or U18465 (N_18465,N_17825,N_17717);
nor U18466 (N_18466,N_17855,N_17690);
nand U18467 (N_18467,N_17863,N_17759);
and U18468 (N_18468,N_17623,N_17558);
or U18469 (N_18469,N_17942,N_17970);
xor U18470 (N_18470,N_17877,N_17549);
xnor U18471 (N_18471,N_17551,N_17917);
and U18472 (N_18472,N_17558,N_17795);
nand U18473 (N_18473,N_17661,N_17591);
nor U18474 (N_18474,N_17843,N_17730);
nor U18475 (N_18475,N_17970,N_17761);
nand U18476 (N_18476,N_17769,N_17921);
xor U18477 (N_18477,N_17619,N_17988);
or U18478 (N_18478,N_17710,N_17911);
or U18479 (N_18479,N_17590,N_17619);
nor U18480 (N_18480,N_17828,N_17709);
nand U18481 (N_18481,N_17539,N_17921);
or U18482 (N_18482,N_17706,N_17972);
nor U18483 (N_18483,N_17829,N_17811);
or U18484 (N_18484,N_17580,N_17905);
or U18485 (N_18485,N_17909,N_17749);
or U18486 (N_18486,N_17587,N_17907);
nor U18487 (N_18487,N_17851,N_17564);
nor U18488 (N_18488,N_17593,N_17582);
and U18489 (N_18489,N_17949,N_17639);
xnor U18490 (N_18490,N_17589,N_17685);
nand U18491 (N_18491,N_17863,N_17810);
or U18492 (N_18492,N_17727,N_17545);
nor U18493 (N_18493,N_17784,N_17520);
nor U18494 (N_18494,N_17963,N_17686);
and U18495 (N_18495,N_17675,N_17656);
or U18496 (N_18496,N_17945,N_17989);
xor U18497 (N_18497,N_17830,N_17566);
and U18498 (N_18498,N_17729,N_17507);
xnor U18499 (N_18499,N_17887,N_17568);
xor U18500 (N_18500,N_18414,N_18235);
nand U18501 (N_18501,N_18335,N_18229);
xnor U18502 (N_18502,N_18195,N_18069);
and U18503 (N_18503,N_18003,N_18178);
xor U18504 (N_18504,N_18361,N_18005);
nand U18505 (N_18505,N_18445,N_18308);
nand U18506 (N_18506,N_18127,N_18274);
nor U18507 (N_18507,N_18175,N_18112);
nor U18508 (N_18508,N_18253,N_18122);
and U18509 (N_18509,N_18219,N_18214);
or U18510 (N_18510,N_18225,N_18306);
or U18511 (N_18511,N_18464,N_18425);
xor U18512 (N_18512,N_18139,N_18140);
xnor U18513 (N_18513,N_18465,N_18418);
xnor U18514 (N_18514,N_18037,N_18338);
xor U18515 (N_18515,N_18288,N_18357);
or U18516 (N_18516,N_18083,N_18384);
nand U18517 (N_18517,N_18018,N_18364);
or U18518 (N_18518,N_18411,N_18055);
or U18519 (N_18519,N_18146,N_18359);
or U18520 (N_18520,N_18071,N_18371);
nand U18521 (N_18521,N_18290,N_18313);
nand U18522 (N_18522,N_18365,N_18156);
or U18523 (N_18523,N_18260,N_18232);
or U18524 (N_18524,N_18120,N_18377);
or U18525 (N_18525,N_18047,N_18258);
nor U18526 (N_18526,N_18309,N_18215);
or U18527 (N_18527,N_18142,N_18378);
xnor U18528 (N_18528,N_18278,N_18349);
nand U18529 (N_18529,N_18273,N_18135);
xnor U18530 (N_18530,N_18486,N_18149);
and U18531 (N_18531,N_18315,N_18342);
or U18532 (N_18532,N_18136,N_18102);
xor U18533 (N_18533,N_18459,N_18341);
nor U18534 (N_18534,N_18011,N_18054);
nand U18535 (N_18535,N_18360,N_18036);
nor U18536 (N_18536,N_18247,N_18297);
or U18537 (N_18537,N_18492,N_18105);
or U18538 (N_18538,N_18075,N_18048);
or U18539 (N_18539,N_18035,N_18222);
nand U18540 (N_18540,N_18299,N_18166);
xor U18541 (N_18541,N_18420,N_18057);
nand U18542 (N_18542,N_18201,N_18022);
and U18543 (N_18543,N_18433,N_18443);
and U18544 (N_18544,N_18391,N_18343);
xnor U18545 (N_18545,N_18482,N_18434);
and U18546 (N_18546,N_18440,N_18495);
nand U18547 (N_18547,N_18056,N_18436);
xor U18548 (N_18548,N_18027,N_18279);
and U18549 (N_18549,N_18295,N_18330);
nor U18550 (N_18550,N_18028,N_18402);
or U18551 (N_18551,N_18078,N_18064);
nor U18552 (N_18552,N_18204,N_18403);
nand U18553 (N_18553,N_18059,N_18467);
or U18554 (N_18554,N_18192,N_18052);
nand U18555 (N_18555,N_18183,N_18014);
nor U18556 (N_18556,N_18179,N_18234);
nor U18557 (N_18557,N_18173,N_18487);
or U18558 (N_18558,N_18145,N_18199);
nor U18559 (N_18559,N_18489,N_18220);
and U18560 (N_18560,N_18478,N_18224);
and U18561 (N_18561,N_18162,N_18472);
nand U18562 (N_18562,N_18031,N_18358);
xnor U18563 (N_18563,N_18292,N_18494);
and U18564 (N_18564,N_18038,N_18163);
or U18565 (N_18565,N_18413,N_18227);
and U18566 (N_18566,N_18421,N_18042);
or U18567 (N_18567,N_18339,N_18311);
xnor U18568 (N_18568,N_18405,N_18032);
or U18569 (N_18569,N_18165,N_18280);
nor U18570 (N_18570,N_18293,N_18491);
or U18571 (N_18571,N_18319,N_18101);
nand U18572 (N_18572,N_18020,N_18068);
nand U18573 (N_18573,N_18372,N_18438);
or U18574 (N_18574,N_18417,N_18114);
nor U18575 (N_18575,N_18354,N_18089);
nand U18576 (N_18576,N_18488,N_18058);
nor U18577 (N_18577,N_18161,N_18226);
xnor U18578 (N_18578,N_18062,N_18450);
xor U18579 (N_18579,N_18133,N_18460);
nor U18580 (N_18580,N_18348,N_18016);
or U18581 (N_18581,N_18250,N_18040);
or U18582 (N_18582,N_18332,N_18408);
or U18583 (N_18583,N_18240,N_18189);
xnor U18584 (N_18584,N_18277,N_18079);
xor U18585 (N_18585,N_18174,N_18256);
and U18586 (N_18586,N_18119,N_18108);
xor U18587 (N_18587,N_18115,N_18254);
nor U18588 (N_18588,N_18001,N_18369);
nand U18589 (N_18589,N_18375,N_18347);
and U18590 (N_18590,N_18368,N_18281);
nand U18591 (N_18591,N_18380,N_18024);
nor U18592 (N_18592,N_18305,N_18289);
or U18593 (N_18593,N_18437,N_18210);
nor U18594 (N_18594,N_18211,N_18117);
and U18595 (N_18595,N_18107,N_18287);
or U18596 (N_18596,N_18294,N_18353);
and U18597 (N_18597,N_18045,N_18216);
nor U18598 (N_18598,N_18186,N_18025);
xor U18599 (N_18599,N_18009,N_18376);
xor U18600 (N_18600,N_18041,N_18346);
xor U18601 (N_18601,N_18096,N_18033);
or U18602 (N_18602,N_18252,N_18385);
nand U18603 (N_18603,N_18030,N_18147);
xor U18604 (N_18604,N_18328,N_18185);
nor U18605 (N_18605,N_18208,N_18312);
and U18606 (N_18606,N_18099,N_18132);
and U18607 (N_18607,N_18326,N_18406);
or U18608 (N_18608,N_18259,N_18271);
nand U18609 (N_18609,N_18412,N_18134);
xnor U18610 (N_18610,N_18017,N_18023);
nor U18611 (N_18611,N_18100,N_18498);
nand U18612 (N_18612,N_18461,N_18409);
or U18613 (N_18613,N_18113,N_18327);
xnor U18614 (N_18614,N_18243,N_18217);
nor U18615 (N_18615,N_18331,N_18382);
and U18616 (N_18616,N_18424,N_18270);
nor U18617 (N_18617,N_18285,N_18388);
or U18618 (N_18618,N_18070,N_18233);
nor U18619 (N_18619,N_18496,N_18065);
and U18620 (N_18620,N_18272,N_18334);
xor U18621 (N_18621,N_18473,N_18021);
nor U18622 (N_18622,N_18060,N_18157);
nand U18623 (N_18623,N_18203,N_18286);
and U18624 (N_18624,N_18144,N_18169);
nor U18625 (N_18625,N_18188,N_18053);
nor U18626 (N_18626,N_18483,N_18439);
and U18627 (N_18627,N_18302,N_18230);
and U18628 (N_18628,N_18257,N_18152);
and U18629 (N_18629,N_18310,N_18410);
nor U18630 (N_18630,N_18168,N_18263);
nand U18631 (N_18631,N_18194,N_18291);
nand U18632 (N_18632,N_18352,N_18479);
xor U18633 (N_18633,N_18092,N_18477);
and U18634 (N_18634,N_18441,N_18088);
nand U18635 (N_18635,N_18457,N_18296);
xor U18636 (N_18636,N_18324,N_18301);
nor U18637 (N_18637,N_18284,N_18317);
and U18638 (N_18638,N_18351,N_18451);
nor U18639 (N_18639,N_18264,N_18176);
and U18640 (N_18640,N_18363,N_18164);
nand U18641 (N_18641,N_18074,N_18399);
xor U18642 (N_18642,N_18000,N_18137);
and U18643 (N_18643,N_18367,N_18172);
xor U18644 (N_18644,N_18141,N_18190);
nor U18645 (N_18645,N_18344,N_18435);
xnor U18646 (N_18646,N_18430,N_18322);
nand U18647 (N_18647,N_18431,N_18298);
or U18648 (N_18648,N_18043,N_18276);
nand U18649 (N_18649,N_18044,N_18387);
and U18650 (N_18650,N_18381,N_18323);
nor U18651 (N_18651,N_18126,N_18366);
or U18652 (N_18652,N_18318,N_18106);
nor U18653 (N_18653,N_18239,N_18193);
or U18654 (N_18654,N_18091,N_18255);
or U18655 (N_18655,N_18104,N_18066);
and U18656 (N_18656,N_18497,N_18238);
and U18657 (N_18657,N_18350,N_18268);
and U18658 (N_18658,N_18029,N_18452);
and U18659 (N_18659,N_18307,N_18373);
or U18660 (N_18660,N_18202,N_18007);
or U18661 (N_18661,N_18182,N_18470);
or U18662 (N_18662,N_18072,N_18077);
nor U18663 (N_18663,N_18475,N_18448);
and U18664 (N_18664,N_18063,N_18223);
or U18665 (N_18665,N_18356,N_18400);
and U18666 (N_18666,N_18158,N_18415);
nand U18667 (N_18667,N_18170,N_18244);
xor U18668 (N_18668,N_18428,N_18006);
and U18669 (N_18669,N_18490,N_18076);
xnor U18670 (N_18670,N_18389,N_18370);
or U18671 (N_18671,N_18466,N_18087);
nand U18672 (N_18672,N_18447,N_18051);
and U18673 (N_18673,N_18432,N_18004);
xnor U18674 (N_18674,N_18167,N_18187);
or U18675 (N_18675,N_18393,N_18148);
nand U18676 (N_18676,N_18196,N_18444);
and U18677 (N_18677,N_18468,N_18419);
and U18678 (N_18678,N_18129,N_18143);
nand U18679 (N_18679,N_18050,N_18159);
nor U18680 (N_18680,N_18153,N_18394);
and U18681 (N_18681,N_18345,N_18265);
nor U18682 (N_18682,N_18218,N_18008);
xnor U18683 (N_18683,N_18177,N_18124);
nor U18684 (N_18684,N_18304,N_18454);
and U18685 (N_18685,N_18160,N_18205);
and U18686 (N_18686,N_18484,N_18336);
xor U18687 (N_18687,N_18407,N_18397);
or U18688 (N_18688,N_18383,N_18171);
and U18689 (N_18689,N_18480,N_18325);
nor U18690 (N_18690,N_18002,N_18155);
nand U18691 (N_18691,N_18207,N_18321);
nand U18692 (N_18692,N_18362,N_18191);
or U18693 (N_18693,N_18493,N_18426);
nor U18694 (N_18694,N_18098,N_18095);
nand U18695 (N_18695,N_18118,N_18404);
nor U18696 (N_18696,N_18320,N_18455);
or U18697 (N_18697,N_18248,N_18019);
nand U18698 (N_18698,N_18228,N_18453);
and U18699 (N_18699,N_18423,N_18231);
and U18700 (N_18700,N_18474,N_18427);
xor U18701 (N_18701,N_18390,N_18396);
and U18702 (N_18702,N_18446,N_18481);
nor U18703 (N_18703,N_18046,N_18249);
nand U18704 (N_18704,N_18109,N_18151);
or U18705 (N_18705,N_18471,N_18476);
xor U18706 (N_18706,N_18355,N_18180);
nor U18707 (N_18707,N_18084,N_18469);
nand U18708 (N_18708,N_18499,N_18485);
xor U18709 (N_18709,N_18121,N_18337);
and U18710 (N_18710,N_18333,N_18340);
nor U18711 (N_18711,N_18422,N_18283);
nor U18712 (N_18712,N_18429,N_18067);
or U18713 (N_18713,N_18209,N_18246);
or U18714 (N_18714,N_18081,N_18269);
nor U18715 (N_18715,N_18090,N_18379);
xor U18716 (N_18716,N_18010,N_18110);
nor U18717 (N_18717,N_18316,N_18462);
and U18718 (N_18718,N_18442,N_18015);
nand U18719 (N_18719,N_18449,N_18131);
nand U18720 (N_18720,N_18103,N_18237);
and U18721 (N_18721,N_18374,N_18049);
nor U18722 (N_18722,N_18080,N_18012);
nand U18723 (N_18723,N_18275,N_18150);
nor U18724 (N_18724,N_18086,N_18034);
and U18725 (N_18725,N_18073,N_18456);
xnor U18726 (N_18726,N_18221,N_18463);
xor U18727 (N_18727,N_18300,N_18097);
and U18728 (N_18728,N_18266,N_18116);
nand U18729 (N_18729,N_18094,N_18154);
xor U18730 (N_18730,N_18181,N_18262);
nor U18731 (N_18731,N_18245,N_18213);
and U18732 (N_18732,N_18200,N_18184);
nor U18733 (N_18733,N_18314,N_18267);
or U18734 (N_18734,N_18398,N_18401);
and U18735 (N_18735,N_18130,N_18082);
and U18736 (N_18736,N_18303,N_18395);
xor U18737 (N_18737,N_18386,N_18212);
and U18738 (N_18738,N_18242,N_18261);
and U18739 (N_18739,N_18458,N_18093);
xnor U18740 (N_18740,N_18125,N_18282);
or U18741 (N_18741,N_18392,N_18061);
or U18742 (N_18742,N_18111,N_18416);
xnor U18743 (N_18743,N_18085,N_18329);
nor U18744 (N_18744,N_18013,N_18138);
and U18745 (N_18745,N_18236,N_18123);
nor U18746 (N_18746,N_18198,N_18197);
and U18747 (N_18747,N_18128,N_18026);
nor U18748 (N_18748,N_18206,N_18241);
nor U18749 (N_18749,N_18039,N_18251);
xor U18750 (N_18750,N_18085,N_18497);
or U18751 (N_18751,N_18442,N_18453);
nand U18752 (N_18752,N_18391,N_18258);
and U18753 (N_18753,N_18117,N_18027);
nand U18754 (N_18754,N_18456,N_18070);
nand U18755 (N_18755,N_18161,N_18267);
or U18756 (N_18756,N_18367,N_18349);
nand U18757 (N_18757,N_18328,N_18301);
xnor U18758 (N_18758,N_18379,N_18035);
nor U18759 (N_18759,N_18329,N_18203);
and U18760 (N_18760,N_18411,N_18230);
xor U18761 (N_18761,N_18092,N_18292);
and U18762 (N_18762,N_18092,N_18418);
nor U18763 (N_18763,N_18014,N_18319);
xnor U18764 (N_18764,N_18253,N_18383);
or U18765 (N_18765,N_18286,N_18298);
and U18766 (N_18766,N_18035,N_18368);
and U18767 (N_18767,N_18261,N_18220);
nor U18768 (N_18768,N_18452,N_18210);
xnor U18769 (N_18769,N_18099,N_18001);
nor U18770 (N_18770,N_18016,N_18244);
or U18771 (N_18771,N_18102,N_18209);
nor U18772 (N_18772,N_18314,N_18264);
nor U18773 (N_18773,N_18091,N_18371);
and U18774 (N_18774,N_18355,N_18219);
and U18775 (N_18775,N_18057,N_18222);
xnor U18776 (N_18776,N_18475,N_18034);
nor U18777 (N_18777,N_18188,N_18111);
nor U18778 (N_18778,N_18285,N_18027);
xor U18779 (N_18779,N_18049,N_18478);
nand U18780 (N_18780,N_18409,N_18426);
xor U18781 (N_18781,N_18348,N_18394);
nor U18782 (N_18782,N_18151,N_18365);
nor U18783 (N_18783,N_18346,N_18480);
and U18784 (N_18784,N_18391,N_18463);
xnor U18785 (N_18785,N_18265,N_18166);
nand U18786 (N_18786,N_18384,N_18239);
or U18787 (N_18787,N_18132,N_18300);
nand U18788 (N_18788,N_18262,N_18303);
or U18789 (N_18789,N_18184,N_18437);
and U18790 (N_18790,N_18465,N_18307);
or U18791 (N_18791,N_18188,N_18395);
and U18792 (N_18792,N_18346,N_18195);
nand U18793 (N_18793,N_18437,N_18151);
or U18794 (N_18794,N_18423,N_18003);
and U18795 (N_18795,N_18426,N_18367);
nor U18796 (N_18796,N_18495,N_18130);
and U18797 (N_18797,N_18250,N_18360);
nand U18798 (N_18798,N_18268,N_18126);
nor U18799 (N_18799,N_18324,N_18071);
nand U18800 (N_18800,N_18442,N_18367);
nor U18801 (N_18801,N_18220,N_18181);
xor U18802 (N_18802,N_18142,N_18060);
and U18803 (N_18803,N_18440,N_18196);
nor U18804 (N_18804,N_18378,N_18038);
nor U18805 (N_18805,N_18400,N_18100);
nor U18806 (N_18806,N_18180,N_18224);
nand U18807 (N_18807,N_18107,N_18024);
or U18808 (N_18808,N_18021,N_18468);
xor U18809 (N_18809,N_18040,N_18225);
nor U18810 (N_18810,N_18411,N_18287);
and U18811 (N_18811,N_18144,N_18337);
xnor U18812 (N_18812,N_18319,N_18424);
and U18813 (N_18813,N_18148,N_18135);
nand U18814 (N_18814,N_18300,N_18108);
nand U18815 (N_18815,N_18005,N_18150);
nand U18816 (N_18816,N_18103,N_18404);
nor U18817 (N_18817,N_18035,N_18109);
nand U18818 (N_18818,N_18376,N_18219);
nand U18819 (N_18819,N_18377,N_18335);
nor U18820 (N_18820,N_18038,N_18030);
nor U18821 (N_18821,N_18260,N_18011);
nor U18822 (N_18822,N_18243,N_18004);
or U18823 (N_18823,N_18013,N_18185);
nand U18824 (N_18824,N_18275,N_18009);
and U18825 (N_18825,N_18363,N_18175);
or U18826 (N_18826,N_18367,N_18049);
nor U18827 (N_18827,N_18326,N_18380);
and U18828 (N_18828,N_18152,N_18357);
nand U18829 (N_18829,N_18139,N_18369);
xor U18830 (N_18830,N_18104,N_18272);
xor U18831 (N_18831,N_18360,N_18302);
nand U18832 (N_18832,N_18102,N_18442);
nor U18833 (N_18833,N_18052,N_18312);
and U18834 (N_18834,N_18183,N_18227);
and U18835 (N_18835,N_18147,N_18057);
nor U18836 (N_18836,N_18094,N_18463);
or U18837 (N_18837,N_18295,N_18227);
nand U18838 (N_18838,N_18344,N_18097);
or U18839 (N_18839,N_18371,N_18147);
or U18840 (N_18840,N_18324,N_18098);
nor U18841 (N_18841,N_18428,N_18049);
nor U18842 (N_18842,N_18025,N_18365);
nand U18843 (N_18843,N_18325,N_18463);
nor U18844 (N_18844,N_18132,N_18380);
xor U18845 (N_18845,N_18088,N_18179);
xnor U18846 (N_18846,N_18364,N_18406);
xor U18847 (N_18847,N_18467,N_18447);
or U18848 (N_18848,N_18199,N_18091);
or U18849 (N_18849,N_18052,N_18000);
or U18850 (N_18850,N_18058,N_18144);
nor U18851 (N_18851,N_18075,N_18333);
nor U18852 (N_18852,N_18469,N_18138);
nor U18853 (N_18853,N_18099,N_18426);
xor U18854 (N_18854,N_18192,N_18428);
xor U18855 (N_18855,N_18162,N_18319);
nor U18856 (N_18856,N_18188,N_18416);
and U18857 (N_18857,N_18462,N_18214);
and U18858 (N_18858,N_18423,N_18083);
xnor U18859 (N_18859,N_18460,N_18065);
nor U18860 (N_18860,N_18488,N_18170);
or U18861 (N_18861,N_18355,N_18485);
and U18862 (N_18862,N_18376,N_18106);
nand U18863 (N_18863,N_18219,N_18383);
and U18864 (N_18864,N_18092,N_18391);
xnor U18865 (N_18865,N_18350,N_18155);
and U18866 (N_18866,N_18396,N_18085);
or U18867 (N_18867,N_18156,N_18205);
nand U18868 (N_18868,N_18449,N_18263);
nor U18869 (N_18869,N_18415,N_18397);
nor U18870 (N_18870,N_18037,N_18422);
xor U18871 (N_18871,N_18332,N_18086);
nand U18872 (N_18872,N_18135,N_18270);
and U18873 (N_18873,N_18122,N_18076);
xor U18874 (N_18874,N_18065,N_18008);
or U18875 (N_18875,N_18027,N_18197);
or U18876 (N_18876,N_18206,N_18057);
nand U18877 (N_18877,N_18221,N_18472);
nor U18878 (N_18878,N_18478,N_18172);
or U18879 (N_18879,N_18186,N_18187);
xnor U18880 (N_18880,N_18422,N_18005);
nor U18881 (N_18881,N_18173,N_18284);
and U18882 (N_18882,N_18493,N_18194);
and U18883 (N_18883,N_18288,N_18222);
and U18884 (N_18884,N_18267,N_18367);
xnor U18885 (N_18885,N_18184,N_18047);
nand U18886 (N_18886,N_18184,N_18315);
nor U18887 (N_18887,N_18323,N_18443);
or U18888 (N_18888,N_18276,N_18089);
nor U18889 (N_18889,N_18054,N_18398);
or U18890 (N_18890,N_18129,N_18220);
xor U18891 (N_18891,N_18089,N_18487);
and U18892 (N_18892,N_18249,N_18168);
nand U18893 (N_18893,N_18002,N_18063);
nor U18894 (N_18894,N_18145,N_18365);
nor U18895 (N_18895,N_18326,N_18236);
nor U18896 (N_18896,N_18158,N_18070);
or U18897 (N_18897,N_18244,N_18302);
nor U18898 (N_18898,N_18443,N_18037);
xnor U18899 (N_18899,N_18255,N_18166);
xor U18900 (N_18900,N_18257,N_18177);
nand U18901 (N_18901,N_18028,N_18295);
and U18902 (N_18902,N_18035,N_18210);
and U18903 (N_18903,N_18289,N_18388);
xnor U18904 (N_18904,N_18151,N_18025);
or U18905 (N_18905,N_18206,N_18306);
nor U18906 (N_18906,N_18438,N_18381);
nand U18907 (N_18907,N_18239,N_18131);
or U18908 (N_18908,N_18476,N_18301);
nand U18909 (N_18909,N_18017,N_18323);
nor U18910 (N_18910,N_18331,N_18299);
nor U18911 (N_18911,N_18125,N_18451);
or U18912 (N_18912,N_18482,N_18017);
and U18913 (N_18913,N_18310,N_18377);
nand U18914 (N_18914,N_18372,N_18016);
and U18915 (N_18915,N_18461,N_18326);
nor U18916 (N_18916,N_18417,N_18392);
nor U18917 (N_18917,N_18483,N_18094);
nor U18918 (N_18918,N_18189,N_18306);
and U18919 (N_18919,N_18141,N_18133);
or U18920 (N_18920,N_18232,N_18218);
nor U18921 (N_18921,N_18434,N_18419);
nor U18922 (N_18922,N_18385,N_18220);
xnor U18923 (N_18923,N_18285,N_18083);
or U18924 (N_18924,N_18142,N_18413);
and U18925 (N_18925,N_18485,N_18030);
xor U18926 (N_18926,N_18266,N_18327);
and U18927 (N_18927,N_18033,N_18293);
or U18928 (N_18928,N_18004,N_18008);
xnor U18929 (N_18929,N_18091,N_18015);
or U18930 (N_18930,N_18060,N_18253);
xor U18931 (N_18931,N_18205,N_18494);
or U18932 (N_18932,N_18272,N_18013);
xor U18933 (N_18933,N_18455,N_18220);
nand U18934 (N_18934,N_18057,N_18279);
and U18935 (N_18935,N_18089,N_18065);
and U18936 (N_18936,N_18409,N_18051);
nand U18937 (N_18937,N_18182,N_18008);
nand U18938 (N_18938,N_18009,N_18184);
or U18939 (N_18939,N_18484,N_18445);
or U18940 (N_18940,N_18261,N_18167);
or U18941 (N_18941,N_18049,N_18479);
and U18942 (N_18942,N_18209,N_18164);
or U18943 (N_18943,N_18461,N_18119);
or U18944 (N_18944,N_18266,N_18333);
nand U18945 (N_18945,N_18386,N_18205);
and U18946 (N_18946,N_18099,N_18104);
or U18947 (N_18947,N_18003,N_18105);
nor U18948 (N_18948,N_18270,N_18066);
nand U18949 (N_18949,N_18221,N_18246);
xor U18950 (N_18950,N_18370,N_18459);
nand U18951 (N_18951,N_18228,N_18002);
nor U18952 (N_18952,N_18414,N_18156);
and U18953 (N_18953,N_18343,N_18255);
or U18954 (N_18954,N_18311,N_18142);
or U18955 (N_18955,N_18469,N_18181);
nor U18956 (N_18956,N_18467,N_18472);
or U18957 (N_18957,N_18286,N_18288);
or U18958 (N_18958,N_18413,N_18314);
nor U18959 (N_18959,N_18174,N_18354);
or U18960 (N_18960,N_18497,N_18455);
nand U18961 (N_18961,N_18197,N_18459);
nor U18962 (N_18962,N_18125,N_18244);
or U18963 (N_18963,N_18189,N_18376);
xnor U18964 (N_18964,N_18078,N_18079);
nand U18965 (N_18965,N_18116,N_18104);
and U18966 (N_18966,N_18058,N_18149);
or U18967 (N_18967,N_18236,N_18477);
nor U18968 (N_18968,N_18045,N_18317);
xor U18969 (N_18969,N_18182,N_18446);
nor U18970 (N_18970,N_18190,N_18367);
nor U18971 (N_18971,N_18483,N_18049);
nor U18972 (N_18972,N_18173,N_18163);
nand U18973 (N_18973,N_18216,N_18499);
xor U18974 (N_18974,N_18435,N_18145);
or U18975 (N_18975,N_18465,N_18147);
or U18976 (N_18976,N_18466,N_18038);
or U18977 (N_18977,N_18328,N_18252);
nor U18978 (N_18978,N_18044,N_18034);
nand U18979 (N_18979,N_18148,N_18259);
nor U18980 (N_18980,N_18247,N_18125);
xnor U18981 (N_18981,N_18455,N_18143);
xor U18982 (N_18982,N_18002,N_18146);
and U18983 (N_18983,N_18110,N_18462);
nand U18984 (N_18984,N_18333,N_18407);
nor U18985 (N_18985,N_18342,N_18220);
nor U18986 (N_18986,N_18165,N_18163);
nor U18987 (N_18987,N_18084,N_18448);
nor U18988 (N_18988,N_18043,N_18201);
or U18989 (N_18989,N_18002,N_18287);
xnor U18990 (N_18990,N_18126,N_18127);
nand U18991 (N_18991,N_18210,N_18465);
nand U18992 (N_18992,N_18187,N_18345);
or U18993 (N_18993,N_18419,N_18377);
or U18994 (N_18994,N_18071,N_18245);
nand U18995 (N_18995,N_18394,N_18068);
nor U18996 (N_18996,N_18118,N_18293);
nand U18997 (N_18997,N_18020,N_18099);
and U18998 (N_18998,N_18473,N_18208);
and U18999 (N_18999,N_18425,N_18125);
nor U19000 (N_19000,N_18983,N_18703);
and U19001 (N_19001,N_18578,N_18612);
or U19002 (N_19002,N_18812,N_18710);
nor U19003 (N_19003,N_18616,N_18760);
xnor U19004 (N_19004,N_18668,N_18518);
and U19005 (N_19005,N_18842,N_18776);
xnor U19006 (N_19006,N_18650,N_18550);
and U19007 (N_19007,N_18818,N_18528);
xnor U19008 (N_19008,N_18510,N_18836);
and U19009 (N_19009,N_18920,N_18608);
and U19010 (N_19010,N_18553,N_18505);
or U19011 (N_19011,N_18744,N_18924);
nor U19012 (N_19012,N_18774,N_18551);
nor U19013 (N_19013,N_18831,N_18893);
xnor U19014 (N_19014,N_18979,N_18565);
nor U19015 (N_19015,N_18596,N_18954);
nand U19016 (N_19016,N_18537,N_18527);
xnor U19017 (N_19017,N_18991,N_18795);
xor U19018 (N_19018,N_18908,N_18732);
or U19019 (N_19019,N_18641,N_18764);
xnor U19020 (N_19020,N_18789,N_18839);
nand U19021 (N_19021,N_18891,N_18773);
and U19022 (N_19022,N_18688,N_18988);
nor U19023 (N_19023,N_18873,N_18556);
nor U19024 (N_19024,N_18782,N_18532);
xnor U19025 (N_19025,N_18677,N_18853);
xor U19026 (N_19026,N_18880,N_18855);
or U19027 (N_19027,N_18775,N_18605);
xnor U19028 (N_19028,N_18548,N_18731);
and U19029 (N_19029,N_18944,N_18826);
or U19030 (N_19030,N_18741,N_18506);
and U19031 (N_19031,N_18805,N_18856);
or U19032 (N_19032,N_18808,N_18657);
nand U19033 (N_19033,N_18685,N_18561);
nand U19034 (N_19034,N_18566,N_18523);
or U19035 (N_19035,N_18723,N_18588);
nor U19036 (N_19036,N_18549,N_18928);
xor U19037 (N_19037,N_18841,N_18868);
nor U19038 (N_19038,N_18984,N_18654);
or U19039 (N_19039,N_18835,N_18909);
nand U19040 (N_19040,N_18907,N_18937);
nor U19041 (N_19041,N_18697,N_18675);
and U19042 (N_19042,N_18680,N_18739);
nor U19043 (N_19043,N_18575,N_18681);
and U19044 (N_19044,N_18734,N_18579);
nand U19045 (N_19045,N_18899,N_18889);
xor U19046 (N_19046,N_18699,N_18923);
and U19047 (N_19047,N_18693,N_18646);
and U19048 (N_19048,N_18500,N_18756);
or U19049 (N_19049,N_18562,N_18571);
or U19050 (N_19050,N_18981,N_18746);
and U19051 (N_19051,N_18629,N_18765);
xor U19052 (N_19052,N_18648,N_18897);
and U19053 (N_19053,N_18757,N_18918);
xnor U19054 (N_19054,N_18963,N_18622);
or U19055 (N_19055,N_18664,N_18535);
nor U19056 (N_19056,N_18867,N_18798);
nor U19057 (N_19057,N_18936,N_18813);
nor U19058 (N_19058,N_18541,N_18787);
nand U19059 (N_19059,N_18905,N_18584);
xnor U19060 (N_19060,N_18559,N_18686);
nand U19061 (N_19061,N_18982,N_18726);
nor U19062 (N_19062,N_18625,N_18717);
xor U19063 (N_19063,N_18806,N_18793);
xor U19064 (N_19064,N_18547,N_18817);
and U19065 (N_19065,N_18887,N_18783);
xnor U19066 (N_19066,N_18862,N_18607);
or U19067 (N_19067,N_18956,N_18847);
nand U19068 (N_19068,N_18930,N_18993);
nand U19069 (N_19069,N_18828,N_18581);
or U19070 (N_19070,N_18632,N_18845);
and U19071 (N_19071,N_18784,N_18910);
and U19072 (N_19072,N_18800,N_18786);
xnor U19073 (N_19073,N_18833,N_18788);
or U19074 (N_19074,N_18978,N_18933);
xnor U19075 (N_19075,N_18673,N_18921);
nor U19076 (N_19076,N_18507,N_18850);
xnor U19077 (N_19077,N_18859,N_18737);
or U19078 (N_19078,N_18687,N_18906);
and U19079 (N_19079,N_18959,N_18848);
and U19080 (N_19080,N_18614,N_18879);
nand U19081 (N_19081,N_18558,N_18631);
xor U19082 (N_19082,N_18722,N_18729);
xnor U19083 (N_19083,N_18792,N_18672);
nand U19084 (N_19084,N_18969,N_18881);
xor U19085 (N_19085,N_18640,N_18740);
or U19086 (N_19086,N_18875,N_18663);
nor U19087 (N_19087,N_18590,N_18595);
and U19088 (N_19088,N_18896,N_18763);
nand U19089 (N_19089,N_18560,N_18957);
nand U19090 (N_19090,N_18621,N_18583);
and U19091 (N_19091,N_18951,N_18700);
nand U19092 (N_19092,N_18692,N_18635);
or U19093 (N_19093,N_18997,N_18724);
nor U19094 (N_19094,N_18846,N_18803);
and U19095 (N_19095,N_18942,N_18623);
and U19096 (N_19096,N_18519,N_18934);
nor U19097 (N_19097,N_18514,N_18759);
xor U19098 (N_19098,N_18667,N_18938);
nor U19099 (N_19099,N_18671,N_18914);
or U19100 (N_19100,N_18515,N_18998);
and U19101 (N_19101,N_18865,N_18554);
nor U19102 (N_19102,N_18661,N_18586);
nand U19103 (N_19103,N_18878,N_18655);
or U19104 (N_19104,N_18642,N_18718);
or U19105 (N_19105,N_18508,N_18949);
and U19106 (N_19106,N_18652,N_18968);
and U19107 (N_19107,N_18609,N_18526);
or U19108 (N_19108,N_18684,N_18822);
xnor U19109 (N_19109,N_18513,N_18585);
and U19110 (N_19110,N_18945,N_18733);
or U19111 (N_19111,N_18962,N_18987);
nand U19112 (N_19112,N_18976,N_18602);
xor U19113 (N_19113,N_18639,N_18854);
and U19114 (N_19114,N_18864,N_18534);
xnor U19115 (N_19115,N_18662,N_18857);
nand U19116 (N_19116,N_18720,N_18502);
nand U19117 (N_19117,N_18870,N_18791);
nand U19118 (N_19118,N_18704,N_18886);
nand U19119 (N_19119,N_18778,N_18863);
or U19120 (N_19120,N_18913,N_18858);
and U19121 (N_19121,N_18917,N_18589);
or U19122 (N_19122,N_18814,N_18545);
xor U19123 (N_19123,N_18838,N_18751);
nand U19124 (N_19124,N_18748,N_18725);
nand U19125 (N_19125,N_18592,N_18999);
and U19126 (N_19126,N_18972,N_18844);
xnor U19127 (N_19127,N_18772,N_18630);
nand U19128 (N_19128,N_18970,N_18929);
nand U19129 (N_19129,N_18883,N_18882);
and U19130 (N_19130,N_18816,N_18678);
or U19131 (N_19131,N_18660,N_18900);
xor U19132 (N_19132,N_18604,N_18536);
or U19133 (N_19133,N_18790,N_18811);
nor U19134 (N_19134,N_18679,N_18591);
and U19135 (N_19135,N_18567,N_18620);
or U19136 (N_19136,N_18649,N_18797);
nand U19137 (N_19137,N_18644,N_18990);
xor U19138 (N_19138,N_18659,N_18960);
xnor U19139 (N_19139,N_18745,N_18587);
xor U19140 (N_19140,N_18669,N_18851);
xor U19141 (N_19141,N_18898,N_18511);
nand U19142 (N_19142,N_18919,N_18958);
or U19143 (N_19143,N_18721,N_18613);
xnor U19144 (N_19144,N_18766,N_18830);
nor U19145 (N_19145,N_18840,N_18645);
and U19146 (N_19146,N_18555,N_18994);
and U19147 (N_19147,N_18824,N_18533);
or U19148 (N_19148,N_18606,N_18577);
xor U19149 (N_19149,N_18735,N_18837);
and U19150 (N_19150,N_18569,N_18593);
xnor U19151 (N_19151,N_18785,N_18985);
nor U19152 (N_19152,N_18801,N_18767);
nand U19153 (N_19153,N_18869,N_18911);
and U19154 (N_19154,N_18706,N_18574);
nand U19155 (N_19155,N_18651,N_18769);
or U19156 (N_19156,N_18807,N_18568);
nor U19157 (N_19157,N_18627,N_18696);
xnor U19158 (N_19158,N_18834,N_18618);
nand U19159 (N_19159,N_18599,N_18825);
and U19160 (N_19160,N_18600,N_18827);
and U19161 (N_19161,N_18674,N_18582);
nand U19162 (N_19162,N_18711,N_18705);
nand U19163 (N_19163,N_18973,N_18638);
or U19164 (N_19164,N_18516,N_18974);
and U19165 (N_19165,N_18815,N_18939);
nor U19166 (N_19166,N_18762,N_18503);
xor U19167 (N_19167,N_18819,N_18755);
nor U19168 (N_19168,N_18989,N_18915);
and U19169 (N_19169,N_18779,N_18892);
or U19170 (N_19170,N_18967,N_18563);
and U19171 (N_19171,N_18714,N_18610);
nor U19172 (N_19172,N_18643,N_18542);
or U19173 (N_19173,N_18932,N_18922);
or U19174 (N_19174,N_18829,N_18874);
nor U19175 (N_19175,N_18916,N_18964);
and U19176 (N_19176,N_18529,N_18953);
and U19177 (N_19177,N_18890,N_18580);
xor U19178 (N_19178,N_18927,N_18736);
nand U19179 (N_19179,N_18658,N_18955);
xor U19180 (N_19180,N_18540,N_18777);
nor U19181 (N_19181,N_18634,N_18738);
or U19182 (N_19182,N_18977,N_18780);
and U19183 (N_19183,N_18617,N_18823);
or U19184 (N_19184,N_18971,N_18520);
or U19185 (N_19185,N_18950,N_18771);
and U19186 (N_19186,N_18702,N_18799);
nand U19187 (N_19187,N_18647,N_18931);
nor U19188 (N_19188,N_18624,N_18576);
xnor U19189 (N_19189,N_18947,N_18986);
nand U19190 (N_19190,N_18758,N_18866);
nor U19191 (N_19191,N_18728,N_18689);
and U19192 (N_19192,N_18531,N_18902);
xnor U19193 (N_19193,N_18885,N_18603);
nand U19194 (N_19194,N_18996,N_18727);
xor U19195 (N_19195,N_18636,N_18543);
nand U19196 (N_19196,N_18925,N_18716);
nand U19197 (N_19197,N_18901,N_18849);
or U19198 (N_19198,N_18653,N_18894);
and U19199 (N_19199,N_18539,N_18572);
nand U19200 (N_19200,N_18517,N_18564);
nand U19201 (N_19201,N_18712,N_18665);
nand U19202 (N_19202,N_18750,N_18530);
nor U19203 (N_19203,N_18707,N_18743);
nand U19204 (N_19204,N_18952,N_18601);
and U19205 (N_19205,N_18912,N_18552);
xnor U19206 (N_19206,N_18796,N_18980);
nor U19207 (N_19207,N_18820,N_18941);
nand U19208 (N_19208,N_18666,N_18754);
xnor U19209 (N_19209,N_18903,N_18676);
xnor U19210 (N_19210,N_18943,N_18656);
nor U19211 (N_19211,N_18695,N_18573);
nand U19212 (N_19212,N_18877,N_18749);
xnor U19213 (N_19213,N_18521,N_18753);
xnor U19214 (N_19214,N_18872,N_18809);
or U19215 (N_19215,N_18935,N_18690);
xnor U19216 (N_19216,N_18966,N_18948);
and U19217 (N_19217,N_18946,N_18509);
and U19218 (N_19218,N_18633,N_18628);
xnor U19219 (N_19219,N_18904,N_18843);
xor U19220 (N_19220,N_18557,N_18670);
xnor U19221 (N_19221,N_18691,N_18730);
nor U19222 (N_19222,N_18876,N_18683);
and U19223 (N_19223,N_18810,N_18995);
and U19224 (N_19224,N_18611,N_18715);
xor U19225 (N_19225,N_18512,N_18501);
nand U19226 (N_19226,N_18709,N_18852);
and U19227 (N_19227,N_18992,N_18522);
and U19228 (N_19228,N_18719,N_18940);
xnor U19229 (N_19229,N_18965,N_18708);
or U19230 (N_19230,N_18975,N_18701);
nor U19231 (N_19231,N_18747,N_18832);
nand U19232 (N_19232,N_18761,N_18861);
nor U19233 (N_19233,N_18926,N_18694);
and U19234 (N_19234,N_18713,N_18544);
xnor U19235 (N_19235,N_18504,N_18619);
xnor U19236 (N_19236,N_18615,N_18637);
nand U19237 (N_19237,N_18794,N_18525);
and U19238 (N_19238,N_18961,N_18802);
or U19239 (N_19239,N_18538,N_18871);
nor U19240 (N_19240,N_18594,N_18570);
or U19241 (N_19241,N_18888,N_18781);
nand U19242 (N_19242,N_18626,N_18682);
nand U19243 (N_19243,N_18598,N_18597);
nor U19244 (N_19244,N_18821,N_18770);
nand U19245 (N_19245,N_18860,N_18698);
nor U19246 (N_19246,N_18546,N_18768);
nand U19247 (N_19247,N_18524,N_18752);
or U19248 (N_19248,N_18895,N_18804);
nand U19249 (N_19249,N_18884,N_18742);
and U19250 (N_19250,N_18858,N_18693);
nand U19251 (N_19251,N_18615,N_18508);
xnor U19252 (N_19252,N_18793,N_18625);
or U19253 (N_19253,N_18551,N_18513);
nand U19254 (N_19254,N_18613,N_18617);
and U19255 (N_19255,N_18847,N_18551);
and U19256 (N_19256,N_18548,N_18961);
nand U19257 (N_19257,N_18625,N_18901);
xor U19258 (N_19258,N_18526,N_18798);
and U19259 (N_19259,N_18661,N_18599);
xor U19260 (N_19260,N_18994,N_18629);
and U19261 (N_19261,N_18625,N_18528);
nor U19262 (N_19262,N_18575,N_18915);
nor U19263 (N_19263,N_18525,N_18817);
xor U19264 (N_19264,N_18596,N_18908);
nor U19265 (N_19265,N_18692,N_18590);
nor U19266 (N_19266,N_18759,N_18734);
xor U19267 (N_19267,N_18949,N_18718);
xnor U19268 (N_19268,N_18998,N_18590);
nand U19269 (N_19269,N_18516,N_18522);
xor U19270 (N_19270,N_18603,N_18771);
xor U19271 (N_19271,N_18897,N_18962);
xnor U19272 (N_19272,N_18527,N_18868);
or U19273 (N_19273,N_18685,N_18934);
and U19274 (N_19274,N_18713,N_18902);
xnor U19275 (N_19275,N_18505,N_18609);
nor U19276 (N_19276,N_18744,N_18507);
nor U19277 (N_19277,N_18575,N_18998);
or U19278 (N_19278,N_18816,N_18962);
nor U19279 (N_19279,N_18687,N_18815);
nor U19280 (N_19280,N_18874,N_18588);
nand U19281 (N_19281,N_18513,N_18715);
nor U19282 (N_19282,N_18741,N_18663);
or U19283 (N_19283,N_18632,N_18655);
nor U19284 (N_19284,N_18544,N_18667);
nand U19285 (N_19285,N_18704,N_18651);
xor U19286 (N_19286,N_18953,N_18769);
nor U19287 (N_19287,N_18677,N_18781);
xor U19288 (N_19288,N_18975,N_18519);
nand U19289 (N_19289,N_18556,N_18772);
and U19290 (N_19290,N_18640,N_18979);
nand U19291 (N_19291,N_18803,N_18754);
or U19292 (N_19292,N_18584,N_18558);
or U19293 (N_19293,N_18879,N_18968);
xnor U19294 (N_19294,N_18584,N_18709);
and U19295 (N_19295,N_18547,N_18611);
nor U19296 (N_19296,N_18996,N_18748);
nor U19297 (N_19297,N_18755,N_18672);
nor U19298 (N_19298,N_18654,N_18674);
xor U19299 (N_19299,N_18731,N_18782);
xor U19300 (N_19300,N_18748,N_18626);
nor U19301 (N_19301,N_18820,N_18932);
nand U19302 (N_19302,N_18589,N_18755);
nand U19303 (N_19303,N_18966,N_18961);
nor U19304 (N_19304,N_18742,N_18711);
xnor U19305 (N_19305,N_18754,N_18692);
and U19306 (N_19306,N_18685,N_18889);
nor U19307 (N_19307,N_18647,N_18511);
and U19308 (N_19308,N_18605,N_18663);
or U19309 (N_19309,N_18580,N_18528);
or U19310 (N_19310,N_18656,N_18850);
or U19311 (N_19311,N_18704,N_18935);
and U19312 (N_19312,N_18807,N_18943);
or U19313 (N_19313,N_18639,N_18878);
nor U19314 (N_19314,N_18771,N_18876);
and U19315 (N_19315,N_18764,N_18848);
or U19316 (N_19316,N_18840,N_18584);
nor U19317 (N_19317,N_18694,N_18655);
nor U19318 (N_19318,N_18608,N_18756);
nor U19319 (N_19319,N_18640,N_18879);
xnor U19320 (N_19320,N_18647,N_18830);
or U19321 (N_19321,N_18661,N_18639);
xnor U19322 (N_19322,N_18706,N_18980);
xor U19323 (N_19323,N_18628,N_18967);
or U19324 (N_19324,N_18731,N_18644);
nor U19325 (N_19325,N_18648,N_18700);
xnor U19326 (N_19326,N_18732,N_18803);
xnor U19327 (N_19327,N_18901,N_18833);
and U19328 (N_19328,N_18510,N_18844);
and U19329 (N_19329,N_18742,N_18689);
or U19330 (N_19330,N_18862,N_18824);
and U19331 (N_19331,N_18981,N_18730);
nor U19332 (N_19332,N_18862,N_18852);
xor U19333 (N_19333,N_18985,N_18578);
nand U19334 (N_19334,N_18600,N_18901);
or U19335 (N_19335,N_18533,N_18905);
nor U19336 (N_19336,N_18568,N_18569);
or U19337 (N_19337,N_18851,N_18931);
nand U19338 (N_19338,N_18721,N_18534);
and U19339 (N_19339,N_18963,N_18835);
nor U19340 (N_19340,N_18754,N_18914);
nor U19341 (N_19341,N_18518,N_18938);
xnor U19342 (N_19342,N_18676,N_18809);
xor U19343 (N_19343,N_18532,N_18737);
nand U19344 (N_19344,N_18518,N_18587);
or U19345 (N_19345,N_18637,N_18594);
nor U19346 (N_19346,N_18899,N_18937);
nor U19347 (N_19347,N_18756,N_18819);
nor U19348 (N_19348,N_18657,N_18773);
nand U19349 (N_19349,N_18946,N_18876);
nand U19350 (N_19350,N_18944,N_18671);
nand U19351 (N_19351,N_18907,N_18579);
or U19352 (N_19352,N_18842,N_18672);
nand U19353 (N_19353,N_18905,N_18648);
xor U19354 (N_19354,N_18728,N_18618);
nand U19355 (N_19355,N_18796,N_18849);
xnor U19356 (N_19356,N_18540,N_18805);
and U19357 (N_19357,N_18863,N_18835);
and U19358 (N_19358,N_18965,N_18613);
and U19359 (N_19359,N_18827,N_18914);
and U19360 (N_19360,N_18898,N_18632);
nor U19361 (N_19361,N_18858,N_18613);
nand U19362 (N_19362,N_18588,N_18653);
or U19363 (N_19363,N_18885,N_18569);
and U19364 (N_19364,N_18536,N_18637);
or U19365 (N_19365,N_18769,N_18975);
or U19366 (N_19366,N_18792,N_18848);
or U19367 (N_19367,N_18538,N_18790);
and U19368 (N_19368,N_18843,N_18621);
and U19369 (N_19369,N_18525,N_18544);
nor U19370 (N_19370,N_18837,N_18631);
and U19371 (N_19371,N_18872,N_18650);
or U19372 (N_19372,N_18832,N_18625);
nand U19373 (N_19373,N_18647,N_18705);
nor U19374 (N_19374,N_18545,N_18572);
nor U19375 (N_19375,N_18812,N_18804);
and U19376 (N_19376,N_18791,N_18695);
xnor U19377 (N_19377,N_18567,N_18804);
or U19378 (N_19378,N_18738,N_18984);
or U19379 (N_19379,N_18694,N_18525);
and U19380 (N_19380,N_18640,N_18933);
and U19381 (N_19381,N_18812,N_18614);
nand U19382 (N_19382,N_18538,N_18710);
or U19383 (N_19383,N_18666,N_18642);
and U19384 (N_19384,N_18946,N_18877);
or U19385 (N_19385,N_18619,N_18875);
and U19386 (N_19386,N_18964,N_18696);
nand U19387 (N_19387,N_18983,N_18773);
and U19388 (N_19388,N_18605,N_18818);
and U19389 (N_19389,N_18743,N_18511);
xnor U19390 (N_19390,N_18703,N_18625);
or U19391 (N_19391,N_18720,N_18976);
nor U19392 (N_19392,N_18833,N_18622);
nand U19393 (N_19393,N_18790,N_18700);
or U19394 (N_19394,N_18755,N_18901);
or U19395 (N_19395,N_18589,N_18579);
and U19396 (N_19396,N_18860,N_18929);
nor U19397 (N_19397,N_18777,N_18738);
and U19398 (N_19398,N_18660,N_18707);
nor U19399 (N_19399,N_18680,N_18556);
nor U19400 (N_19400,N_18939,N_18908);
or U19401 (N_19401,N_18894,N_18884);
and U19402 (N_19402,N_18519,N_18681);
or U19403 (N_19403,N_18665,N_18701);
nand U19404 (N_19404,N_18953,N_18723);
nor U19405 (N_19405,N_18995,N_18586);
or U19406 (N_19406,N_18772,N_18568);
and U19407 (N_19407,N_18647,N_18699);
nor U19408 (N_19408,N_18539,N_18589);
nand U19409 (N_19409,N_18695,N_18651);
and U19410 (N_19410,N_18856,N_18955);
nand U19411 (N_19411,N_18830,N_18750);
nor U19412 (N_19412,N_18914,N_18631);
nor U19413 (N_19413,N_18628,N_18744);
xnor U19414 (N_19414,N_18751,N_18852);
nor U19415 (N_19415,N_18747,N_18791);
or U19416 (N_19416,N_18504,N_18572);
xnor U19417 (N_19417,N_18617,N_18600);
nand U19418 (N_19418,N_18953,N_18993);
xnor U19419 (N_19419,N_18849,N_18801);
and U19420 (N_19420,N_18504,N_18579);
nor U19421 (N_19421,N_18786,N_18815);
nor U19422 (N_19422,N_18503,N_18734);
and U19423 (N_19423,N_18617,N_18949);
nor U19424 (N_19424,N_18698,N_18657);
xnor U19425 (N_19425,N_18922,N_18698);
nor U19426 (N_19426,N_18658,N_18684);
nand U19427 (N_19427,N_18741,N_18563);
xnor U19428 (N_19428,N_18531,N_18545);
nand U19429 (N_19429,N_18730,N_18605);
nand U19430 (N_19430,N_18523,N_18872);
nor U19431 (N_19431,N_18985,N_18833);
xor U19432 (N_19432,N_18589,N_18892);
nor U19433 (N_19433,N_18625,N_18676);
and U19434 (N_19434,N_18710,N_18865);
xnor U19435 (N_19435,N_18900,N_18714);
nand U19436 (N_19436,N_18629,N_18696);
nand U19437 (N_19437,N_18584,N_18950);
or U19438 (N_19438,N_18546,N_18796);
nand U19439 (N_19439,N_18852,N_18985);
and U19440 (N_19440,N_18563,N_18963);
nand U19441 (N_19441,N_18528,N_18967);
nand U19442 (N_19442,N_18852,N_18551);
and U19443 (N_19443,N_18875,N_18605);
xnor U19444 (N_19444,N_18895,N_18714);
nor U19445 (N_19445,N_18520,N_18725);
nand U19446 (N_19446,N_18752,N_18511);
or U19447 (N_19447,N_18564,N_18682);
nor U19448 (N_19448,N_18640,N_18617);
nor U19449 (N_19449,N_18910,N_18632);
or U19450 (N_19450,N_18514,N_18636);
nand U19451 (N_19451,N_18607,N_18915);
xor U19452 (N_19452,N_18525,N_18735);
nor U19453 (N_19453,N_18895,N_18869);
xnor U19454 (N_19454,N_18709,N_18712);
and U19455 (N_19455,N_18672,N_18573);
nor U19456 (N_19456,N_18586,N_18999);
xnor U19457 (N_19457,N_18739,N_18913);
nor U19458 (N_19458,N_18842,N_18513);
nand U19459 (N_19459,N_18811,N_18740);
xnor U19460 (N_19460,N_18892,N_18588);
nor U19461 (N_19461,N_18524,N_18991);
xnor U19462 (N_19462,N_18770,N_18689);
or U19463 (N_19463,N_18657,N_18812);
and U19464 (N_19464,N_18508,N_18663);
or U19465 (N_19465,N_18885,N_18531);
nand U19466 (N_19466,N_18811,N_18879);
or U19467 (N_19467,N_18583,N_18994);
nand U19468 (N_19468,N_18848,N_18993);
nor U19469 (N_19469,N_18980,N_18734);
nand U19470 (N_19470,N_18701,N_18951);
or U19471 (N_19471,N_18897,N_18890);
or U19472 (N_19472,N_18616,N_18712);
xnor U19473 (N_19473,N_18760,N_18643);
and U19474 (N_19474,N_18919,N_18942);
or U19475 (N_19475,N_18670,N_18993);
or U19476 (N_19476,N_18566,N_18873);
nor U19477 (N_19477,N_18684,N_18772);
and U19478 (N_19478,N_18668,N_18545);
nor U19479 (N_19479,N_18541,N_18771);
and U19480 (N_19480,N_18623,N_18990);
nor U19481 (N_19481,N_18902,N_18911);
nor U19482 (N_19482,N_18963,N_18644);
nand U19483 (N_19483,N_18870,N_18705);
and U19484 (N_19484,N_18843,N_18722);
nor U19485 (N_19485,N_18781,N_18836);
xor U19486 (N_19486,N_18711,N_18807);
nor U19487 (N_19487,N_18867,N_18743);
nand U19488 (N_19488,N_18900,N_18636);
and U19489 (N_19489,N_18906,N_18600);
nor U19490 (N_19490,N_18517,N_18979);
or U19491 (N_19491,N_18885,N_18735);
nand U19492 (N_19492,N_18599,N_18783);
nand U19493 (N_19493,N_18969,N_18897);
nor U19494 (N_19494,N_18653,N_18699);
or U19495 (N_19495,N_18987,N_18929);
nand U19496 (N_19496,N_18642,N_18796);
and U19497 (N_19497,N_18616,N_18955);
and U19498 (N_19498,N_18535,N_18906);
and U19499 (N_19499,N_18805,N_18701);
or U19500 (N_19500,N_19251,N_19385);
nor U19501 (N_19501,N_19407,N_19244);
nand U19502 (N_19502,N_19393,N_19491);
and U19503 (N_19503,N_19367,N_19169);
xor U19504 (N_19504,N_19143,N_19261);
and U19505 (N_19505,N_19135,N_19262);
nand U19506 (N_19506,N_19125,N_19126);
or U19507 (N_19507,N_19032,N_19316);
xor U19508 (N_19508,N_19395,N_19119);
and U19509 (N_19509,N_19483,N_19268);
xor U19510 (N_19510,N_19083,N_19120);
nor U19511 (N_19511,N_19109,N_19495);
nand U19512 (N_19512,N_19200,N_19285);
nor U19513 (N_19513,N_19248,N_19409);
and U19514 (N_19514,N_19026,N_19089);
nor U19515 (N_19515,N_19353,N_19490);
xor U19516 (N_19516,N_19423,N_19192);
nor U19517 (N_19517,N_19401,N_19412);
nor U19518 (N_19518,N_19343,N_19272);
or U19519 (N_19519,N_19184,N_19332);
nand U19520 (N_19520,N_19070,N_19374);
nand U19521 (N_19521,N_19445,N_19267);
nand U19522 (N_19522,N_19221,N_19336);
nor U19523 (N_19523,N_19290,N_19339);
or U19524 (N_19524,N_19060,N_19094);
nand U19525 (N_19525,N_19075,N_19213);
xnor U19526 (N_19526,N_19039,N_19322);
or U19527 (N_19527,N_19313,N_19054);
and U19528 (N_19528,N_19325,N_19159);
xor U19529 (N_19529,N_19074,N_19266);
nand U19530 (N_19530,N_19277,N_19252);
or U19531 (N_19531,N_19052,N_19034);
xnor U19532 (N_19532,N_19150,N_19116);
nor U19533 (N_19533,N_19370,N_19319);
nand U19534 (N_19534,N_19173,N_19376);
nand U19535 (N_19535,N_19097,N_19382);
or U19536 (N_19536,N_19420,N_19241);
nor U19537 (N_19537,N_19431,N_19455);
nand U19538 (N_19538,N_19471,N_19334);
xnor U19539 (N_19539,N_19003,N_19225);
nor U19540 (N_19540,N_19410,N_19389);
and U19541 (N_19541,N_19162,N_19098);
nor U19542 (N_19542,N_19207,N_19247);
or U19543 (N_19543,N_19442,N_19182);
and U19544 (N_19544,N_19007,N_19388);
nand U19545 (N_19545,N_19246,N_19362);
nand U19546 (N_19546,N_19363,N_19286);
nor U19547 (N_19547,N_19292,N_19335);
nor U19548 (N_19548,N_19327,N_19373);
xnor U19549 (N_19549,N_19440,N_19172);
nand U19550 (N_19550,N_19441,N_19149);
nand U19551 (N_19551,N_19309,N_19137);
or U19552 (N_19552,N_19183,N_19411);
nand U19553 (N_19553,N_19085,N_19274);
xor U19554 (N_19554,N_19293,N_19091);
nor U19555 (N_19555,N_19042,N_19078);
and U19556 (N_19556,N_19458,N_19379);
or U19557 (N_19557,N_19047,N_19381);
xor U19558 (N_19558,N_19044,N_19051);
or U19559 (N_19559,N_19392,N_19289);
and U19560 (N_19560,N_19228,N_19038);
nor U19561 (N_19561,N_19255,N_19354);
xor U19562 (N_19562,N_19204,N_19396);
nand U19563 (N_19563,N_19421,N_19488);
nand U19564 (N_19564,N_19282,N_19259);
and U19565 (N_19565,N_19180,N_19002);
nand U19566 (N_19566,N_19498,N_19114);
or U19567 (N_19567,N_19365,N_19337);
or U19568 (N_19568,N_19364,N_19361);
xnor U19569 (N_19569,N_19022,N_19186);
and U19570 (N_19570,N_19185,N_19131);
xnor U19571 (N_19571,N_19233,N_19095);
nand U19572 (N_19572,N_19256,N_19099);
xnor U19573 (N_19573,N_19071,N_19346);
nand U19574 (N_19574,N_19000,N_19090);
nand U19575 (N_19575,N_19459,N_19171);
nand U19576 (N_19576,N_19064,N_19310);
xnor U19577 (N_19577,N_19201,N_19303);
and U19578 (N_19578,N_19275,N_19477);
nor U19579 (N_19579,N_19073,N_19250);
or U19580 (N_19580,N_19174,N_19219);
and U19581 (N_19581,N_19470,N_19300);
and U19582 (N_19582,N_19062,N_19128);
nor U19583 (N_19583,N_19462,N_19359);
or U19584 (N_19584,N_19140,N_19072);
xnor U19585 (N_19585,N_19168,N_19108);
xnor U19586 (N_19586,N_19156,N_19017);
or U19587 (N_19587,N_19058,N_19028);
or U19588 (N_19588,N_19155,N_19176);
or U19589 (N_19589,N_19190,N_19066);
xnor U19590 (N_19590,N_19245,N_19306);
xor U19591 (N_19591,N_19350,N_19144);
xor U19592 (N_19592,N_19428,N_19311);
or U19593 (N_19593,N_19271,N_19341);
and U19594 (N_19594,N_19175,N_19307);
and U19595 (N_19595,N_19209,N_19068);
or U19596 (N_19596,N_19480,N_19013);
and U19597 (N_19597,N_19076,N_19067);
xnor U19598 (N_19598,N_19460,N_19181);
xnor U19599 (N_19599,N_19467,N_19427);
nand U19600 (N_19600,N_19351,N_19419);
or U19601 (N_19601,N_19036,N_19400);
or U19602 (N_19602,N_19340,N_19096);
nand U19603 (N_19603,N_19375,N_19088);
nor U19604 (N_19604,N_19291,N_19435);
or U19605 (N_19605,N_19029,N_19283);
or U19606 (N_19606,N_19104,N_19386);
and U19607 (N_19607,N_19280,N_19199);
xnor U19608 (N_19608,N_19037,N_19284);
or U19609 (N_19609,N_19197,N_19105);
and U19610 (N_19610,N_19206,N_19012);
nand U19611 (N_19611,N_19254,N_19122);
nor U19612 (N_19612,N_19321,N_19496);
xor U19613 (N_19613,N_19258,N_19178);
nor U19614 (N_19614,N_19242,N_19317);
or U19615 (N_19615,N_19232,N_19004);
or U19616 (N_19616,N_19234,N_19314);
nand U19617 (N_19617,N_19148,N_19408);
nand U19618 (N_19618,N_19499,N_19205);
and U19619 (N_19619,N_19451,N_19299);
nor U19620 (N_19620,N_19492,N_19121);
nand U19621 (N_19621,N_19448,N_19265);
xor U19622 (N_19622,N_19124,N_19236);
or U19623 (N_19623,N_19239,N_19253);
nand U19624 (N_19624,N_19461,N_19115);
nor U19625 (N_19625,N_19323,N_19330);
nand U19626 (N_19626,N_19019,N_19413);
xnor U19627 (N_19627,N_19151,N_19117);
nor U19628 (N_19628,N_19005,N_19422);
nand U19629 (N_19629,N_19191,N_19216);
and U19630 (N_19630,N_19018,N_19161);
and U19631 (N_19631,N_19304,N_19160);
and U19632 (N_19632,N_19482,N_19298);
or U19633 (N_19633,N_19223,N_19033);
xor U19634 (N_19634,N_19348,N_19404);
or U19635 (N_19635,N_19100,N_19092);
nand U19636 (N_19636,N_19009,N_19086);
nor U19637 (N_19637,N_19424,N_19065);
nand U19638 (N_19638,N_19043,N_19390);
and U19639 (N_19639,N_19011,N_19473);
nor U19640 (N_19640,N_19456,N_19152);
nor U19641 (N_19641,N_19006,N_19249);
nand U19642 (N_19642,N_19497,N_19080);
and U19643 (N_19643,N_19194,N_19118);
xnor U19644 (N_19644,N_19287,N_19464);
or U19645 (N_19645,N_19438,N_19481);
and U19646 (N_19646,N_19103,N_19203);
xor U19647 (N_19647,N_19113,N_19046);
and U19648 (N_19648,N_19057,N_19315);
nor U19649 (N_19649,N_19479,N_19305);
and U19650 (N_19650,N_19188,N_19264);
nor U19651 (N_19651,N_19406,N_19243);
or U19652 (N_19652,N_19324,N_19031);
nand U19653 (N_19653,N_19202,N_19278);
or U19654 (N_19654,N_19157,N_19165);
or U19655 (N_19655,N_19050,N_19452);
or U19656 (N_19656,N_19449,N_19329);
and U19657 (N_19657,N_19147,N_19312);
or U19658 (N_19658,N_19237,N_19081);
and U19659 (N_19659,N_19153,N_19399);
and U19660 (N_19660,N_19023,N_19465);
and U19661 (N_19661,N_19260,N_19432);
nand U19662 (N_19662,N_19338,N_19053);
xnor U19663 (N_19663,N_19403,N_19416);
nor U19664 (N_19664,N_19391,N_19195);
and U19665 (N_19665,N_19133,N_19356);
xnor U19666 (N_19666,N_19257,N_19487);
nand U19667 (N_19667,N_19270,N_19357);
nor U19668 (N_19668,N_19418,N_19468);
nor U19669 (N_19669,N_19166,N_19426);
nor U19670 (N_19670,N_19218,N_19170);
or U19671 (N_19671,N_19387,N_19102);
nor U19672 (N_19672,N_19358,N_19222);
or U19673 (N_19673,N_19443,N_19189);
and U19674 (N_19674,N_19417,N_19110);
and U19675 (N_19675,N_19444,N_19301);
xnor U19676 (N_19676,N_19484,N_19235);
or U19677 (N_19677,N_19154,N_19130);
or U19678 (N_19678,N_19297,N_19035);
xnor U19679 (N_19679,N_19106,N_19308);
xnor U19680 (N_19680,N_19405,N_19048);
and U19681 (N_19681,N_19326,N_19024);
nor U19682 (N_19682,N_19331,N_19238);
or U19683 (N_19683,N_19472,N_19215);
nand U19684 (N_19684,N_19025,N_19129);
xnor U19685 (N_19685,N_19021,N_19476);
or U19686 (N_19686,N_19041,N_19141);
nand U19687 (N_19687,N_19055,N_19457);
xor U19688 (N_19688,N_19352,N_19177);
and U19689 (N_19689,N_19123,N_19415);
xnor U19690 (N_19690,N_19230,N_19059);
xnor U19691 (N_19691,N_19107,N_19224);
nor U19692 (N_19692,N_19402,N_19061);
or U19693 (N_19693,N_19077,N_19378);
or U19694 (N_19694,N_19069,N_19474);
nand U19695 (N_19695,N_19210,N_19231);
xor U19696 (N_19696,N_19214,N_19030);
xor U19697 (N_19697,N_19138,N_19229);
nor U19698 (N_19698,N_19295,N_19447);
and U19699 (N_19699,N_19016,N_19145);
xor U19700 (N_19700,N_19478,N_19079);
xor U19701 (N_19701,N_19276,N_19014);
and U19702 (N_19702,N_19369,N_19333);
and U19703 (N_19703,N_19198,N_19084);
or U19704 (N_19704,N_19063,N_19093);
and U19705 (N_19705,N_19087,N_19494);
nor U19706 (N_19706,N_19429,N_19439);
or U19707 (N_19707,N_19227,N_19040);
or U19708 (N_19708,N_19240,N_19273);
nor U19709 (N_19709,N_19027,N_19134);
nand U19710 (N_19710,N_19366,N_19434);
nor U19711 (N_19711,N_19394,N_19454);
nor U19712 (N_19712,N_19463,N_19008);
xor U19713 (N_19713,N_19049,N_19453);
and U19714 (N_19714,N_19020,N_19486);
nand U19715 (N_19715,N_19111,N_19001);
nor U19716 (N_19716,N_19318,N_19187);
and U19717 (N_19717,N_19475,N_19045);
and U19718 (N_19718,N_19485,N_19212);
nor U19719 (N_19719,N_19056,N_19146);
nand U19720 (N_19720,N_19398,N_19211);
nor U19721 (N_19721,N_19437,N_19281);
nor U19722 (N_19722,N_19344,N_19158);
nand U19723 (N_19723,N_19446,N_19371);
or U19724 (N_19724,N_19163,N_19164);
or U19725 (N_19725,N_19279,N_19179);
or U19726 (N_19726,N_19112,N_19302);
xnor U19727 (N_19727,N_19368,N_19493);
and U19728 (N_19728,N_19372,N_19489);
xnor U19729 (N_19729,N_19217,N_19433);
or U19730 (N_19730,N_19015,N_19127);
nand U19731 (N_19731,N_19132,N_19136);
and U19732 (N_19732,N_19196,N_19377);
nand U19733 (N_19733,N_19355,N_19430);
nand U19734 (N_19734,N_19263,N_19101);
nor U19735 (N_19735,N_19397,N_19167);
and U19736 (N_19736,N_19328,N_19220);
nand U19737 (N_19737,N_19414,N_19347);
xor U19738 (N_19738,N_19082,N_19269);
and U19739 (N_19739,N_19320,N_19466);
xor U19740 (N_19740,N_19383,N_19139);
xor U19741 (N_19741,N_19384,N_19349);
nor U19742 (N_19742,N_19436,N_19226);
or U19743 (N_19743,N_19469,N_19380);
xor U19744 (N_19744,N_19296,N_19193);
nand U19745 (N_19745,N_19360,N_19342);
xor U19746 (N_19746,N_19142,N_19425);
or U19747 (N_19747,N_19010,N_19345);
or U19748 (N_19748,N_19450,N_19294);
nand U19749 (N_19749,N_19288,N_19208);
and U19750 (N_19750,N_19204,N_19493);
xnor U19751 (N_19751,N_19102,N_19377);
or U19752 (N_19752,N_19149,N_19097);
xnor U19753 (N_19753,N_19370,N_19260);
xnor U19754 (N_19754,N_19223,N_19284);
and U19755 (N_19755,N_19467,N_19091);
or U19756 (N_19756,N_19384,N_19156);
nor U19757 (N_19757,N_19361,N_19434);
nand U19758 (N_19758,N_19017,N_19476);
or U19759 (N_19759,N_19404,N_19205);
or U19760 (N_19760,N_19359,N_19436);
or U19761 (N_19761,N_19244,N_19198);
xnor U19762 (N_19762,N_19477,N_19102);
nand U19763 (N_19763,N_19361,N_19471);
xor U19764 (N_19764,N_19033,N_19465);
nand U19765 (N_19765,N_19273,N_19258);
xor U19766 (N_19766,N_19257,N_19279);
or U19767 (N_19767,N_19102,N_19098);
xor U19768 (N_19768,N_19082,N_19482);
nor U19769 (N_19769,N_19120,N_19162);
nor U19770 (N_19770,N_19417,N_19264);
and U19771 (N_19771,N_19443,N_19181);
nor U19772 (N_19772,N_19149,N_19400);
nand U19773 (N_19773,N_19407,N_19239);
and U19774 (N_19774,N_19272,N_19333);
xor U19775 (N_19775,N_19033,N_19350);
or U19776 (N_19776,N_19097,N_19011);
nand U19777 (N_19777,N_19453,N_19289);
xor U19778 (N_19778,N_19365,N_19297);
nor U19779 (N_19779,N_19240,N_19175);
nand U19780 (N_19780,N_19201,N_19254);
xor U19781 (N_19781,N_19149,N_19044);
nor U19782 (N_19782,N_19084,N_19416);
and U19783 (N_19783,N_19269,N_19442);
nor U19784 (N_19784,N_19067,N_19031);
and U19785 (N_19785,N_19043,N_19317);
or U19786 (N_19786,N_19013,N_19344);
nand U19787 (N_19787,N_19230,N_19003);
or U19788 (N_19788,N_19131,N_19049);
and U19789 (N_19789,N_19304,N_19189);
nand U19790 (N_19790,N_19404,N_19322);
nand U19791 (N_19791,N_19450,N_19002);
xor U19792 (N_19792,N_19469,N_19313);
or U19793 (N_19793,N_19017,N_19135);
or U19794 (N_19794,N_19207,N_19064);
and U19795 (N_19795,N_19426,N_19327);
nand U19796 (N_19796,N_19252,N_19342);
and U19797 (N_19797,N_19358,N_19302);
nor U19798 (N_19798,N_19096,N_19469);
xnor U19799 (N_19799,N_19080,N_19293);
nor U19800 (N_19800,N_19263,N_19230);
or U19801 (N_19801,N_19171,N_19140);
nor U19802 (N_19802,N_19034,N_19012);
and U19803 (N_19803,N_19379,N_19273);
or U19804 (N_19804,N_19415,N_19354);
nor U19805 (N_19805,N_19053,N_19128);
nand U19806 (N_19806,N_19473,N_19055);
xor U19807 (N_19807,N_19404,N_19136);
xnor U19808 (N_19808,N_19401,N_19131);
xnor U19809 (N_19809,N_19199,N_19256);
xor U19810 (N_19810,N_19143,N_19010);
xor U19811 (N_19811,N_19385,N_19359);
nand U19812 (N_19812,N_19386,N_19207);
nand U19813 (N_19813,N_19107,N_19278);
and U19814 (N_19814,N_19481,N_19487);
nor U19815 (N_19815,N_19154,N_19102);
and U19816 (N_19816,N_19463,N_19450);
xnor U19817 (N_19817,N_19478,N_19499);
xnor U19818 (N_19818,N_19389,N_19468);
nor U19819 (N_19819,N_19393,N_19486);
xor U19820 (N_19820,N_19183,N_19335);
and U19821 (N_19821,N_19358,N_19351);
or U19822 (N_19822,N_19218,N_19090);
and U19823 (N_19823,N_19429,N_19321);
nand U19824 (N_19824,N_19407,N_19066);
xnor U19825 (N_19825,N_19446,N_19135);
and U19826 (N_19826,N_19485,N_19108);
nand U19827 (N_19827,N_19306,N_19392);
nor U19828 (N_19828,N_19386,N_19391);
and U19829 (N_19829,N_19308,N_19306);
nand U19830 (N_19830,N_19250,N_19378);
nand U19831 (N_19831,N_19042,N_19276);
nand U19832 (N_19832,N_19151,N_19171);
nand U19833 (N_19833,N_19093,N_19251);
or U19834 (N_19834,N_19071,N_19497);
nor U19835 (N_19835,N_19212,N_19414);
and U19836 (N_19836,N_19231,N_19303);
and U19837 (N_19837,N_19404,N_19098);
or U19838 (N_19838,N_19462,N_19026);
nand U19839 (N_19839,N_19439,N_19155);
nand U19840 (N_19840,N_19006,N_19314);
nand U19841 (N_19841,N_19312,N_19471);
xor U19842 (N_19842,N_19170,N_19015);
and U19843 (N_19843,N_19412,N_19150);
nor U19844 (N_19844,N_19290,N_19393);
xnor U19845 (N_19845,N_19184,N_19491);
nor U19846 (N_19846,N_19114,N_19087);
nor U19847 (N_19847,N_19237,N_19408);
xnor U19848 (N_19848,N_19297,N_19468);
nand U19849 (N_19849,N_19276,N_19401);
nor U19850 (N_19850,N_19206,N_19315);
or U19851 (N_19851,N_19207,N_19146);
or U19852 (N_19852,N_19098,N_19402);
and U19853 (N_19853,N_19200,N_19017);
nor U19854 (N_19854,N_19473,N_19433);
or U19855 (N_19855,N_19154,N_19354);
xor U19856 (N_19856,N_19200,N_19140);
and U19857 (N_19857,N_19174,N_19069);
and U19858 (N_19858,N_19446,N_19056);
nor U19859 (N_19859,N_19057,N_19372);
and U19860 (N_19860,N_19414,N_19329);
nand U19861 (N_19861,N_19027,N_19156);
xor U19862 (N_19862,N_19305,N_19142);
nand U19863 (N_19863,N_19422,N_19414);
and U19864 (N_19864,N_19191,N_19136);
and U19865 (N_19865,N_19360,N_19206);
nor U19866 (N_19866,N_19281,N_19004);
and U19867 (N_19867,N_19408,N_19139);
and U19868 (N_19868,N_19423,N_19420);
xnor U19869 (N_19869,N_19032,N_19449);
and U19870 (N_19870,N_19257,N_19080);
nand U19871 (N_19871,N_19231,N_19011);
and U19872 (N_19872,N_19310,N_19176);
xnor U19873 (N_19873,N_19482,N_19047);
nor U19874 (N_19874,N_19458,N_19331);
nor U19875 (N_19875,N_19398,N_19338);
xnor U19876 (N_19876,N_19006,N_19254);
and U19877 (N_19877,N_19059,N_19093);
and U19878 (N_19878,N_19097,N_19304);
nand U19879 (N_19879,N_19169,N_19207);
nand U19880 (N_19880,N_19460,N_19441);
xor U19881 (N_19881,N_19292,N_19485);
xor U19882 (N_19882,N_19010,N_19445);
nand U19883 (N_19883,N_19280,N_19279);
or U19884 (N_19884,N_19017,N_19130);
or U19885 (N_19885,N_19457,N_19307);
and U19886 (N_19886,N_19043,N_19487);
nor U19887 (N_19887,N_19126,N_19448);
xnor U19888 (N_19888,N_19262,N_19108);
nor U19889 (N_19889,N_19231,N_19152);
or U19890 (N_19890,N_19234,N_19340);
xnor U19891 (N_19891,N_19222,N_19469);
nand U19892 (N_19892,N_19351,N_19340);
nor U19893 (N_19893,N_19022,N_19496);
nand U19894 (N_19894,N_19498,N_19226);
xnor U19895 (N_19895,N_19040,N_19402);
nand U19896 (N_19896,N_19284,N_19464);
nand U19897 (N_19897,N_19477,N_19071);
or U19898 (N_19898,N_19290,N_19338);
or U19899 (N_19899,N_19288,N_19242);
nor U19900 (N_19900,N_19419,N_19284);
xor U19901 (N_19901,N_19078,N_19447);
nor U19902 (N_19902,N_19320,N_19281);
and U19903 (N_19903,N_19165,N_19095);
nor U19904 (N_19904,N_19114,N_19365);
xor U19905 (N_19905,N_19164,N_19170);
nand U19906 (N_19906,N_19492,N_19325);
nor U19907 (N_19907,N_19126,N_19341);
nand U19908 (N_19908,N_19253,N_19414);
and U19909 (N_19909,N_19013,N_19120);
nand U19910 (N_19910,N_19398,N_19004);
xnor U19911 (N_19911,N_19429,N_19157);
and U19912 (N_19912,N_19170,N_19385);
or U19913 (N_19913,N_19489,N_19186);
or U19914 (N_19914,N_19345,N_19198);
nor U19915 (N_19915,N_19222,N_19062);
or U19916 (N_19916,N_19279,N_19050);
xnor U19917 (N_19917,N_19345,N_19172);
or U19918 (N_19918,N_19304,N_19397);
or U19919 (N_19919,N_19195,N_19011);
or U19920 (N_19920,N_19196,N_19192);
and U19921 (N_19921,N_19385,N_19059);
nand U19922 (N_19922,N_19365,N_19256);
xor U19923 (N_19923,N_19392,N_19105);
nand U19924 (N_19924,N_19176,N_19246);
nor U19925 (N_19925,N_19482,N_19290);
or U19926 (N_19926,N_19275,N_19254);
or U19927 (N_19927,N_19251,N_19114);
and U19928 (N_19928,N_19386,N_19282);
or U19929 (N_19929,N_19417,N_19412);
nand U19930 (N_19930,N_19499,N_19103);
xor U19931 (N_19931,N_19268,N_19383);
and U19932 (N_19932,N_19383,N_19154);
or U19933 (N_19933,N_19287,N_19030);
nand U19934 (N_19934,N_19088,N_19220);
or U19935 (N_19935,N_19040,N_19006);
and U19936 (N_19936,N_19357,N_19323);
and U19937 (N_19937,N_19233,N_19081);
and U19938 (N_19938,N_19159,N_19431);
nand U19939 (N_19939,N_19452,N_19321);
and U19940 (N_19940,N_19366,N_19491);
nor U19941 (N_19941,N_19046,N_19464);
and U19942 (N_19942,N_19393,N_19418);
nor U19943 (N_19943,N_19467,N_19487);
and U19944 (N_19944,N_19181,N_19033);
or U19945 (N_19945,N_19394,N_19039);
xor U19946 (N_19946,N_19384,N_19057);
and U19947 (N_19947,N_19442,N_19126);
and U19948 (N_19948,N_19234,N_19217);
and U19949 (N_19949,N_19337,N_19353);
nor U19950 (N_19950,N_19243,N_19239);
and U19951 (N_19951,N_19289,N_19317);
or U19952 (N_19952,N_19226,N_19301);
nand U19953 (N_19953,N_19152,N_19304);
nor U19954 (N_19954,N_19178,N_19112);
nand U19955 (N_19955,N_19449,N_19203);
xnor U19956 (N_19956,N_19285,N_19019);
or U19957 (N_19957,N_19358,N_19117);
or U19958 (N_19958,N_19275,N_19140);
and U19959 (N_19959,N_19222,N_19151);
and U19960 (N_19960,N_19180,N_19243);
nor U19961 (N_19961,N_19093,N_19315);
and U19962 (N_19962,N_19428,N_19149);
nand U19963 (N_19963,N_19249,N_19158);
xnor U19964 (N_19964,N_19449,N_19282);
nand U19965 (N_19965,N_19283,N_19097);
nand U19966 (N_19966,N_19090,N_19072);
and U19967 (N_19967,N_19032,N_19003);
nand U19968 (N_19968,N_19402,N_19250);
xor U19969 (N_19969,N_19337,N_19057);
nand U19970 (N_19970,N_19241,N_19457);
nand U19971 (N_19971,N_19386,N_19449);
nand U19972 (N_19972,N_19351,N_19399);
or U19973 (N_19973,N_19146,N_19151);
nand U19974 (N_19974,N_19336,N_19172);
or U19975 (N_19975,N_19299,N_19290);
nand U19976 (N_19976,N_19258,N_19444);
or U19977 (N_19977,N_19402,N_19107);
and U19978 (N_19978,N_19010,N_19326);
nand U19979 (N_19979,N_19433,N_19108);
or U19980 (N_19980,N_19470,N_19252);
nor U19981 (N_19981,N_19319,N_19132);
xor U19982 (N_19982,N_19128,N_19459);
nand U19983 (N_19983,N_19349,N_19194);
nor U19984 (N_19984,N_19013,N_19465);
nand U19985 (N_19985,N_19277,N_19357);
xor U19986 (N_19986,N_19019,N_19303);
and U19987 (N_19987,N_19432,N_19497);
nand U19988 (N_19988,N_19095,N_19423);
nor U19989 (N_19989,N_19321,N_19431);
or U19990 (N_19990,N_19186,N_19359);
xnor U19991 (N_19991,N_19217,N_19252);
or U19992 (N_19992,N_19457,N_19169);
nor U19993 (N_19993,N_19195,N_19271);
and U19994 (N_19994,N_19163,N_19068);
nor U19995 (N_19995,N_19226,N_19018);
xor U19996 (N_19996,N_19036,N_19186);
nand U19997 (N_19997,N_19025,N_19012);
or U19998 (N_19998,N_19342,N_19044);
nor U19999 (N_19999,N_19352,N_19086);
or U20000 (N_20000,N_19589,N_19528);
or U20001 (N_20001,N_19646,N_19556);
nand U20002 (N_20002,N_19779,N_19650);
nand U20003 (N_20003,N_19816,N_19967);
nand U20004 (N_20004,N_19615,N_19711);
or U20005 (N_20005,N_19707,N_19503);
nand U20006 (N_20006,N_19795,N_19899);
nand U20007 (N_20007,N_19643,N_19935);
nor U20008 (N_20008,N_19818,N_19680);
xnor U20009 (N_20009,N_19530,N_19738);
and U20010 (N_20010,N_19681,N_19790);
nand U20011 (N_20011,N_19671,N_19732);
and U20012 (N_20012,N_19662,N_19888);
and U20013 (N_20013,N_19989,N_19629);
nand U20014 (N_20014,N_19870,N_19939);
xnor U20015 (N_20015,N_19983,N_19927);
nor U20016 (N_20016,N_19801,N_19729);
xnor U20017 (N_20017,N_19630,N_19976);
nor U20018 (N_20018,N_19830,N_19676);
nand U20019 (N_20019,N_19514,N_19552);
nand U20020 (N_20020,N_19708,N_19743);
and U20021 (N_20021,N_19561,N_19992);
nand U20022 (N_20022,N_19597,N_19858);
nor U20023 (N_20023,N_19600,N_19672);
and U20024 (N_20024,N_19544,N_19808);
and U20025 (N_20025,N_19928,N_19756);
and U20026 (N_20026,N_19962,N_19762);
xor U20027 (N_20027,N_19796,N_19724);
and U20028 (N_20028,N_19894,N_19938);
nand U20029 (N_20029,N_19917,N_19698);
or U20030 (N_20030,N_19730,N_19506);
nand U20031 (N_20031,N_19523,N_19726);
or U20032 (N_20032,N_19820,N_19909);
nand U20033 (N_20033,N_19720,N_19865);
xor U20034 (N_20034,N_19896,N_19925);
and U20035 (N_20035,N_19573,N_19777);
nor U20036 (N_20036,N_19673,N_19863);
xnor U20037 (N_20037,N_19789,N_19933);
nand U20038 (N_20038,N_19731,N_19803);
nor U20039 (N_20039,N_19821,N_19970);
or U20040 (N_20040,N_19778,N_19594);
xnor U20041 (N_20041,N_19761,N_19860);
or U20042 (N_20042,N_19807,N_19524);
nor U20043 (N_20043,N_19554,N_19620);
xnor U20044 (N_20044,N_19575,N_19760);
nand U20045 (N_20045,N_19607,N_19840);
nand U20046 (N_20046,N_19640,N_19563);
and U20047 (N_20047,N_19621,N_19576);
and U20048 (N_20048,N_19966,N_19519);
xnor U20049 (N_20049,N_19531,N_19715);
or U20050 (N_20050,N_19583,N_19608);
nand U20051 (N_20051,N_19587,N_19771);
or U20052 (N_20052,N_19866,N_19787);
nor U20053 (N_20053,N_19581,N_19892);
and U20054 (N_20054,N_19659,N_19986);
xnor U20055 (N_20055,N_19669,N_19915);
nor U20056 (N_20056,N_19695,N_19572);
and U20057 (N_20057,N_19522,N_19831);
xor U20058 (N_20058,N_19977,N_19601);
or U20059 (N_20059,N_19668,N_19532);
or U20060 (N_20060,N_19757,N_19670);
xnor U20061 (N_20061,N_19826,N_19565);
nand U20062 (N_20062,N_19947,N_19623);
xnor U20063 (N_20063,N_19798,N_19759);
xor U20064 (N_20064,N_19658,N_19929);
nand U20065 (N_20065,N_19926,N_19855);
nand U20066 (N_20066,N_19805,N_19919);
and U20067 (N_20067,N_19702,N_19815);
nor U20068 (N_20068,N_19609,N_19722);
xnor U20069 (N_20069,N_19585,N_19534);
and U20070 (N_20070,N_19752,N_19686);
xnor U20071 (N_20071,N_19675,N_19543);
nand U20072 (N_20072,N_19800,N_19644);
nand U20073 (N_20073,N_19758,N_19536);
nor U20074 (N_20074,N_19958,N_19905);
and U20075 (N_20075,N_19748,N_19509);
nor U20076 (N_20076,N_19952,N_19690);
nand U20077 (N_20077,N_19613,N_19973);
or U20078 (N_20078,N_19736,N_19584);
or U20079 (N_20079,N_19737,N_19740);
xor U20080 (N_20080,N_19603,N_19525);
nor U20081 (N_20081,N_19734,N_19971);
or U20082 (N_20082,N_19775,N_19501);
xnor U20083 (N_20083,N_19988,N_19604);
nor U20084 (N_20084,N_19990,N_19867);
nor U20085 (N_20085,N_19555,N_19537);
or U20086 (N_20086,N_19793,N_19912);
nand U20087 (N_20087,N_19904,N_19961);
and U20088 (N_20088,N_19836,N_19750);
and U20089 (N_20089,N_19873,N_19857);
and U20090 (N_20090,N_19746,N_19540);
or U20091 (N_20091,N_19813,N_19879);
or U20092 (N_20092,N_19588,N_19774);
nand U20093 (N_20093,N_19817,N_19665);
nand U20094 (N_20094,N_19957,N_19595);
nor U20095 (N_20095,N_19824,N_19767);
nand U20096 (N_20096,N_19586,N_19780);
and U20097 (N_20097,N_19984,N_19578);
or U20098 (N_20098,N_19797,N_19869);
xnor U20099 (N_20099,N_19985,N_19785);
nor U20100 (N_20100,N_19768,N_19900);
or U20101 (N_20101,N_19764,N_19922);
xnor U20102 (N_20102,N_19940,N_19545);
nor U20103 (N_20103,N_19846,N_19642);
nand U20104 (N_20104,N_19688,N_19747);
and U20105 (N_20105,N_19721,N_19877);
and U20106 (N_20106,N_19645,N_19546);
nand U20107 (N_20107,N_19685,N_19507);
or U20108 (N_20108,N_19728,N_19599);
and U20109 (N_20109,N_19932,N_19923);
or U20110 (N_20110,N_19641,N_19814);
and U20111 (N_20111,N_19626,N_19784);
and U20112 (N_20112,N_19705,N_19710);
nor U20113 (N_20113,N_19974,N_19968);
xnor U20114 (N_20114,N_19852,N_19513);
nand U20115 (N_20115,N_19849,N_19677);
and U20116 (N_20116,N_19618,N_19663);
nor U20117 (N_20117,N_19749,N_19625);
nand U20118 (N_20118,N_19516,N_19825);
nor U20119 (N_20119,N_19794,N_19822);
or U20120 (N_20120,N_19723,N_19874);
nor U20121 (N_20121,N_19713,N_19882);
or U20122 (N_20122,N_19717,N_19689);
nor U20123 (N_20123,N_19885,N_19944);
xor U20124 (N_20124,N_19934,N_19907);
xor U20125 (N_20125,N_19611,N_19886);
nor U20126 (N_20126,N_19636,N_19898);
nor U20127 (N_20127,N_19500,N_19521);
xor U20128 (N_20128,N_19835,N_19624);
nand U20129 (N_20129,N_19804,N_19580);
or U20130 (N_20130,N_19602,N_19833);
or U20131 (N_20131,N_19678,N_19960);
and U20132 (N_20132,N_19511,N_19828);
nor U20133 (N_20133,N_19911,N_19535);
and U20134 (N_20134,N_19570,N_19941);
and U20135 (N_20135,N_19868,N_19776);
and U20136 (N_20136,N_19745,N_19725);
or U20137 (N_20137,N_19943,N_19810);
and U20138 (N_20138,N_19978,N_19802);
and U20139 (N_20139,N_19884,N_19742);
and U20140 (N_20140,N_19812,N_19963);
and U20141 (N_20141,N_19766,N_19861);
nand U20142 (N_20142,N_19949,N_19549);
and U20143 (N_20143,N_19679,N_19508);
and U20144 (N_20144,N_19781,N_19667);
and U20145 (N_20145,N_19755,N_19652);
and U20146 (N_20146,N_19605,N_19741);
and U20147 (N_20147,N_19548,N_19969);
and U20148 (N_20148,N_19862,N_19916);
nand U20149 (N_20149,N_19674,N_19553);
nor U20150 (N_20150,N_19753,N_19950);
xnor U20151 (N_20151,N_19859,N_19591);
or U20152 (N_20152,N_19700,N_19851);
and U20153 (N_20153,N_19829,N_19633);
nor U20154 (N_20154,N_19965,N_19533);
or U20155 (N_20155,N_19878,N_19655);
nor U20156 (N_20156,N_19617,N_19881);
or U20157 (N_20157,N_19632,N_19701);
and U20158 (N_20158,N_19982,N_19538);
and U20159 (N_20159,N_19612,N_19619);
xor U20160 (N_20160,N_19704,N_19693);
and U20161 (N_20161,N_19913,N_19844);
or U20162 (N_20162,N_19582,N_19683);
and U20163 (N_20163,N_19541,N_19845);
xnor U20164 (N_20164,N_19997,N_19930);
xor U20165 (N_20165,N_19651,N_19864);
or U20166 (N_20166,N_19590,N_19527);
nor U20167 (N_20167,N_19991,N_19579);
nor U20168 (N_20168,N_19765,N_19666);
xnor U20169 (N_20169,N_19614,N_19703);
or U20170 (N_20170,N_19931,N_19903);
nand U20171 (N_20171,N_19754,N_19788);
or U20172 (N_20172,N_19924,N_19980);
and U20173 (N_20173,N_19890,N_19637);
and U20174 (N_20174,N_19512,N_19566);
nand U20175 (N_20175,N_19843,N_19712);
or U20176 (N_20176,N_19769,N_19786);
xnor U20177 (N_20177,N_19850,N_19918);
or U20178 (N_20178,N_19975,N_19735);
or U20179 (N_20179,N_19834,N_19593);
and U20180 (N_20180,N_19598,N_19964);
and U20181 (N_20181,N_19838,N_19706);
and U20182 (N_20182,N_19887,N_19856);
or U20183 (N_20183,N_19709,N_19751);
and U20184 (N_20184,N_19647,N_19891);
or U20185 (N_20185,N_19889,N_19773);
or U20186 (N_20186,N_19987,N_19772);
nor U20187 (N_20187,N_19648,N_19517);
nand U20188 (N_20188,N_19687,N_19719);
or U20189 (N_20189,N_19520,N_19994);
nor U20190 (N_20190,N_19691,N_19639);
xnor U20191 (N_20191,N_19592,N_19782);
xor U20192 (N_20192,N_19848,N_19638);
nand U20193 (N_20193,N_19562,N_19956);
nor U20194 (N_20194,N_19569,N_19656);
or U20195 (N_20195,N_19577,N_19610);
or U20196 (N_20196,N_19694,N_19551);
and U20197 (N_20197,N_19951,N_19875);
xor U20198 (N_20198,N_19895,N_19606);
nor U20199 (N_20199,N_19634,N_19854);
and U20200 (N_20200,N_19953,N_19998);
nor U20201 (N_20201,N_19839,N_19799);
nor U20202 (N_20202,N_19574,N_19557);
xor U20203 (N_20203,N_19559,N_19937);
nor U20204 (N_20204,N_19893,N_19832);
nor U20205 (N_20205,N_19946,N_19628);
nand U20206 (N_20206,N_19567,N_19616);
nand U20207 (N_20207,N_19502,N_19999);
xor U20208 (N_20208,N_19550,N_19727);
and U20209 (N_20209,N_19819,N_19979);
or U20210 (N_20210,N_19806,N_19910);
nand U20211 (N_20211,N_19547,N_19504);
nor U20212 (N_20212,N_19542,N_19635);
or U20213 (N_20213,N_19718,N_19841);
nand U20214 (N_20214,N_19995,N_19906);
nor U20215 (N_20215,N_19770,N_19955);
xnor U20216 (N_20216,N_19847,N_19733);
nor U20217 (N_20217,N_19872,N_19954);
or U20218 (N_20218,N_19791,N_19653);
nor U20219 (N_20219,N_19526,N_19972);
or U20220 (N_20220,N_19661,N_19897);
xnor U20221 (N_20221,N_19827,N_19853);
or U20222 (N_20222,N_19518,N_19837);
nand U20223 (N_20223,N_19654,N_19871);
nand U20224 (N_20224,N_19739,N_19842);
and U20225 (N_20225,N_19993,N_19792);
and U20226 (N_20226,N_19914,N_19696);
xnor U20227 (N_20227,N_19783,N_19811);
and U20228 (N_20228,N_19515,N_19959);
nor U20229 (N_20229,N_19908,N_19631);
xnor U20230 (N_20230,N_19981,N_19823);
and U20231 (N_20231,N_19716,N_19948);
xnor U20232 (N_20232,N_19560,N_19763);
xnor U20233 (N_20233,N_19664,N_19505);
or U20234 (N_20234,N_19684,N_19558);
nor U20235 (N_20235,N_19996,N_19649);
xor U20236 (N_20236,N_19902,N_19880);
or U20237 (N_20237,N_19660,N_19809);
nand U20238 (N_20238,N_19622,N_19627);
or U20239 (N_20239,N_19921,N_19699);
nor U20240 (N_20240,N_19682,N_19744);
nor U20241 (N_20241,N_19596,N_19564);
nor U20242 (N_20242,N_19571,N_19920);
nor U20243 (N_20243,N_19539,N_19657);
nand U20244 (N_20244,N_19942,N_19692);
or U20245 (N_20245,N_19510,N_19697);
nand U20246 (N_20246,N_19901,N_19568);
nor U20247 (N_20247,N_19529,N_19945);
nand U20248 (N_20248,N_19714,N_19936);
or U20249 (N_20249,N_19876,N_19883);
xor U20250 (N_20250,N_19568,N_19966);
nand U20251 (N_20251,N_19747,N_19671);
nor U20252 (N_20252,N_19676,N_19620);
or U20253 (N_20253,N_19645,N_19960);
nand U20254 (N_20254,N_19939,N_19840);
nand U20255 (N_20255,N_19696,N_19817);
or U20256 (N_20256,N_19556,N_19871);
nor U20257 (N_20257,N_19577,N_19608);
nand U20258 (N_20258,N_19961,N_19988);
or U20259 (N_20259,N_19639,N_19961);
or U20260 (N_20260,N_19927,N_19970);
xnor U20261 (N_20261,N_19720,N_19832);
and U20262 (N_20262,N_19905,N_19770);
nor U20263 (N_20263,N_19920,N_19872);
xnor U20264 (N_20264,N_19716,N_19651);
or U20265 (N_20265,N_19560,N_19984);
and U20266 (N_20266,N_19521,N_19796);
xnor U20267 (N_20267,N_19894,N_19779);
and U20268 (N_20268,N_19887,N_19828);
nand U20269 (N_20269,N_19836,N_19920);
xor U20270 (N_20270,N_19791,N_19890);
and U20271 (N_20271,N_19532,N_19885);
nand U20272 (N_20272,N_19913,N_19617);
xor U20273 (N_20273,N_19890,N_19754);
or U20274 (N_20274,N_19735,N_19873);
xor U20275 (N_20275,N_19799,N_19615);
or U20276 (N_20276,N_19619,N_19679);
nand U20277 (N_20277,N_19698,N_19923);
nor U20278 (N_20278,N_19869,N_19995);
nand U20279 (N_20279,N_19736,N_19970);
nor U20280 (N_20280,N_19862,N_19588);
or U20281 (N_20281,N_19852,N_19770);
nand U20282 (N_20282,N_19937,N_19976);
nand U20283 (N_20283,N_19755,N_19572);
and U20284 (N_20284,N_19808,N_19691);
and U20285 (N_20285,N_19954,N_19598);
xor U20286 (N_20286,N_19666,N_19994);
or U20287 (N_20287,N_19746,N_19524);
nor U20288 (N_20288,N_19943,N_19582);
nor U20289 (N_20289,N_19756,N_19975);
nor U20290 (N_20290,N_19586,N_19577);
xnor U20291 (N_20291,N_19785,N_19942);
and U20292 (N_20292,N_19794,N_19696);
nand U20293 (N_20293,N_19517,N_19815);
or U20294 (N_20294,N_19504,N_19754);
and U20295 (N_20295,N_19906,N_19700);
nor U20296 (N_20296,N_19952,N_19757);
and U20297 (N_20297,N_19866,N_19594);
nor U20298 (N_20298,N_19938,N_19577);
or U20299 (N_20299,N_19803,N_19954);
xor U20300 (N_20300,N_19818,N_19589);
and U20301 (N_20301,N_19861,N_19813);
and U20302 (N_20302,N_19538,N_19570);
nand U20303 (N_20303,N_19829,N_19557);
nor U20304 (N_20304,N_19613,N_19974);
and U20305 (N_20305,N_19699,N_19746);
nand U20306 (N_20306,N_19748,N_19757);
and U20307 (N_20307,N_19633,N_19528);
nand U20308 (N_20308,N_19568,N_19828);
and U20309 (N_20309,N_19687,N_19981);
and U20310 (N_20310,N_19676,N_19942);
nor U20311 (N_20311,N_19876,N_19821);
or U20312 (N_20312,N_19638,N_19681);
nand U20313 (N_20313,N_19932,N_19546);
or U20314 (N_20314,N_19606,N_19555);
and U20315 (N_20315,N_19705,N_19713);
xor U20316 (N_20316,N_19793,N_19980);
or U20317 (N_20317,N_19571,N_19583);
or U20318 (N_20318,N_19902,N_19576);
nor U20319 (N_20319,N_19672,N_19875);
or U20320 (N_20320,N_19979,N_19895);
xnor U20321 (N_20321,N_19934,N_19936);
nor U20322 (N_20322,N_19829,N_19698);
nand U20323 (N_20323,N_19553,N_19817);
nor U20324 (N_20324,N_19632,N_19872);
xnor U20325 (N_20325,N_19747,N_19692);
nor U20326 (N_20326,N_19782,N_19725);
and U20327 (N_20327,N_19924,N_19725);
or U20328 (N_20328,N_19858,N_19706);
nand U20329 (N_20329,N_19713,N_19579);
nor U20330 (N_20330,N_19823,N_19561);
nor U20331 (N_20331,N_19530,N_19795);
and U20332 (N_20332,N_19838,N_19870);
xor U20333 (N_20333,N_19789,N_19585);
and U20334 (N_20334,N_19815,N_19832);
and U20335 (N_20335,N_19734,N_19942);
or U20336 (N_20336,N_19704,N_19780);
xnor U20337 (N_20337,N_19753,N_19640);
and U20338 (N_20338,N_19523,N_19567);
or U20339 (N_20339,N_19710,N_19838);
and U20340 (N_20340,N_19905,N_19581);
nor U20341 (N_20341,N_19783,N_19571);
and U20342 (N_20342,N_19932,N_19837);
xnor U20343 (N_20343,N_19757,N_19974);
nand U20344 (N_20344,N_19724,N_19937);
nand U20345 (N_20345,N_19875,N_19562);
nand U20346 (N_20346,N_19692,N_19886);
nor U20347 (N_20347,N_19865,N_19665);
xor U20348 (N_20348,N_19751,N_19752);
and U20349 (N_20349,N_19754,N_19640);
and U20350 (N_20350,N_19801,N_19912);
nand U20351 (N_20351,N_19879,N_19981);
and U20352 (N_20352,N_19940,N_19927);
xor U20353 (N_20353,N_19710,N_19756);
nor U20354 (N_20354,N_19632,N_19821);
and U20355 (N_20355,N_19504,N_19635);
or U20356 (N_20356,N_19888,N_19533);
xor U20357 (N_20357,N_19660,N_19805);
nor U20358 (N_20358,N_19997,N_19531);
nor U20359 (N_20359,N_19619,N_19794);
nand U20360 (N_20360,N_19783,N_19865);
nor U20361 (N_20361,N_19705,N_19656);
or U20362 (N_20362,N_19702,N_19715);
nor U20363 (N_20363,N_19708,N_19675);
xor U20364 (N_20364,N_19946,N_19764);
nor U20365 (N_20365,N_19522,N_19608);
and U20366 (N_20366,N_19953,N_19964);
and U20367 (N_20367,N_19573,N_19871);
or U20368 (N_20368,N_19771,N_19821);
or U20369 (N_20369,N_19701,N_19694);
nor U20370 (N_20370,N_19634,N_19514);
or U20371 (N_20371,N_19801,N_19861);
xor U20372 (N_20372,N_19680,N_19971);
or U20373 (N_20373,N_19961,N_19835);
xnor U20374 (N_20374,N_19758,N_19520);
and U20375 (N_20375,N_19883,N_19878);
nand U20376 (N_20376,N_19767,N_19980);
nor U20377 (N_20377,N_19826,N_19913);
and U20378 (N_20378,N_19702,N_19958);
nor U20379 (N_20379,N_19571,N_19938);
nor U20380 (N_20380,N_19978,N_19839);
nor U20381 (N_20381,N_19575,N_19828);
nand U20382 (N_20382,N_19559,N_19638);
or U20383 (N_20383,N_19866,N_19592);
nor U20384 (N_20384,N_19633,N_19593);
xor U20385 (N_20385,N_19722,N_19595);
nor U20386 (N_20386,N_19740,N_19754);
xnor U20387 (N_20387,N_19568,N_19732);
xor U20388 (N_20388,N_19547,N_19946);
xnor U20389 (N_20389,N_19713,N_19592);
nand U20390 (N_20390,N_19759,N_19775);
nand U20391 (N_20391,N_19986,N_19501);
nand U20392 (N_20392,N_19606,N_19620);
nor U20393 (N_20393,N_19810,N_19898);
nor U20394 (N_20394,N_19857,N_19604);
and U20395 (N_20395,N_19655,N_19912);
nor U20396 (N_20396,N_19603,N_19748);
or U20397 (N_20397,N_19553,N_19753);
nand U20398 (N_20398,N_19762,N_19846);
or U20399 (N_20399,N_19931,N_19842);
nand U20400 (N_20400,N_19898,N_19579);
xor U20401 (N_20401,N_19929,N_19580);
or U20402 (N_20402,N_19921,N_19865);
and U20403 (N_20403,N_19689,N_19798);
and U20404 (N_20404,N_19665,N_19813);
and U20405 (N_20405,N_19978,N_19588);
or U20406 (N_20406,N_19610,N_19700);
nand U20407 (N_20407,N_19921,N_19873);
nand U20408 (N_20408,N_19724,N_19744);
or U20409 (N_20409,N_19892,N_19502);
and U20410 (N_20410,N_19899,N_19837);
nand U20411 (N_20411,N_19520,N_19912);
xor U20412 (N_20412,N_19942,N_19788);
nand U20413 (N_20413,N_19912,N_19800);
nand U20414 (N_20414,N_19649,N_19794);
nor U20415 (N_20415,N_19878,N_19608);
nand U20416 (N_20416,N_19765,N_19536);
xor U20417 (N_20417,N_19951,N_19735);
nand U20418 (N_20418,N_19994,N_19933);
and U20419 (N_20419,N_19953,N_19922);
xor U20420 (N_20420,N_19806,N_19829);
xor U20421 (N_20421,N_19524,N_19550);
nand U20422 (N_20422,N_19797,N_19615);
and U20423 (N_20423,N_19871,N_19555);
nand U20424 (N_20424,N_19504,N_19748);
or U20425 (N_20425,N_19915,N_19710);
and U20426 (N_20426,N_19936,N_19908);
or U20427 (N_20427,N_19723,N_19846);
nor U20428 (N_20428,N_19804,N_19617);
xor U20429 (N_20429,N_19857,N_19913);
or U20430 (N_20430,N_19626,N_19663);
or U20431 (N_20431,N_19771,N_19972);
nand U20432 (N_20432,N_19570,N_19556);
nor U20433 (N_20433,N_19720,N_19601);
nor U20434 (N_20434,N_19735,N_19656);
nand U20435 (N_20435,N_19793,N_19820);
and U20436 (N_20436,N_19617,N_19759);
nand U20437 (N_20437,N_19783,N_19747);
nor U20438 (N_20438,N_19559,N_19545);
or U20439 (N_20439,N_19836,N_19527);
or U20440 (N_20440,N_19712,N_19514);
and U20441 (N_20441,N_19653,N_19871);
and U20442 (N_20442,N_19721,N_19527);
and U20443 (N_20443,N_19679,N_19894);
or U20444 (N_20444,N_19837,N_19641);
or U20445 (N_20445,N_19848,N_19832);
nand U20446 (N_20446,N_19549,N_19955);
and U20447 (N_20447,N_19713,N_19703);
nor U20448 (N_20448,N_19737,N_19808);
xor U20449 (N_20449,N_19511,N_19964);
nand U20450 (N_20450,N_19588,N_19842);
nor U20451 (N_20451,N_19645,N_19751);
or U20452 (N_20452,N_19708,N_19600);
or U20453 (N_20453,N_19589,N_19839);
or U20454 (N_20454,N_19958,N_19945);
xor U20455 (N_20455,N_19946,N_19732);
nand U20456 (N_20456,N_19710,N_19638);
xor U20457 (N_20457,N_19539,N_19999);
or U20458 (N_20458,N_19512,N_19519);
and U20459 (N_20459,N_19971,N_19621);
or U20460 (N_20460,N_19573,N_19825);
nor U20461 (N_20461,N_19981,N_19862);
nor U20462 (N_20462,N_19842,N_19854);
or U20463 (N_20463,N_19875,N_19698);
nand U20464 (N_20464,N_19963,N_19583);
nand U20465 (N_20465,N_19600,N_19868);
or U20466 (N_20466,N_19818,N_19986);
or U20467 (N_20467,N_19833,N_19909);
nor U20468 (N_20468,N_19601,N_19595);
xor U20469 (N_20469,N_19774,N_19690);
or U20470 (N_20470,N_19526,N_19957);
nand U20471 (N_20471,N_19647,N_19610);
or U20472 (N_20472,N_19704,N_19903);
nand U20473 (N_20473,N_19963,N_19956);
xor U20474 (N_20474,N_19835,N_19719);
nand U20475 (N_20475,N_19537,N_19849);
nor U20476 (N_20476,N_19601,N_19617);
and U20477 (N_20477,N_19881,N_19583);
xnor U20478 (N_20478,N_19812,N_19557);
nor U20479 (N_20479,N_19704,N_19817);
xnor U20480 (N_20480,N_19729,N_19513);
nand U20481 (N_20481,N_19776,N_19618);
xor U20482 (N_20482,N_19949,N_19976);
xnor U20483 (N_20483,N_19834,N_19865);
nand U20484 (N_20484,N_19522,N_19715);
or U20485 (N_20485,N_19752,N_19532);
nor U20486 (N_20486,N_19744,N_19780);
and U20487 (N_20487,N_19872,N_19533);
and U20488 (N_20488,N_19698,N_19993);
and U20489 (N_20489,N_19501,N_19949);
and U20490 (N_20490,N_19927,N_19883);
or U20491 (N_20491,N_19585,N_19677);
xor U20492 (N_20492,N_19535,N_19799);
nor U20493 (N_20493,N_19542,N_19773);
nor U20494 (N_20494,N_19520,N_19939);
nand U20495 (N_20495,N_19981,N_19751);
and U20496 (N_20496,N_19543,N_19879);
or U20497 (N_20497,N_19500,N_19997);
nor U20498 (N_20498,N_19512,N_19995);
nor U20499 (N_20499,N_19564,N_19685);
xnor U20500 (N_20500,N_20077,N_20176);
or U20501 (N_20501,N_20262,N_20268);
nand U20502 (N_20502,N_20399,N_20273);
or U20503 (N_20503,N_20103,N_20412);
or U20504 (N_20504,N_20290,N_20130);
or U20505 (N_20505,N_20180,N_20123);
xnor U20506 (N_20506,N_20096,N_20187);
xor U20507 (N_20507,N_20026,N_20174);
nand U20508 (N_20508,N_20189,N_20163);
nand U20509 (N_20509,N_20377,N_20051);
or U20510 (N_20510,N_20479,N_20379);
or U20511 (N_20511,N_20141,N_20284);
and U20512 (N_20512,N_20069,N_20138);
nor U20513 (N_20513,N_20373,N_20211);
and U20514 (N_20514,N_20229,N_20129);
nand U20515 (N_20515,N_20046,N_20318);
or U20516 (N_20516,N_20116,N_20212);
nor U20517 (N_20517,N_20342,N_20220);
nand U20518 (N_20518,N_20246,N_20252);
nor U20519 (N_20519,N_20192,N_20428);
xnor U20520 (N_20520,N_20283,N_20094);
nor U20521 (N_20521,N_20242,N_20425);
nor U20522 (N_20522,N_20397,N_20119);
xnor U20523 (N_20523,N_20167,N_20148);
nor U20524 (N_20524,N_20477,N_20156);
xnor U20525 (N_20525,N_20074,N_20169);
xor U20526 (N_20526,N_20300,N_20054);
nor U20527 (N_20527,N_20408,N_20392);
and U20528 (N_20528,N_20272,N_20150);
xnor U20529 (N_20529,N_20128,N_20291);
and U20530 (N_20530,N_20228,N_20437);
or U20531 (N_20531,N_20249,N_20430);
or U20532 (N_20532,N_20222,N_20137);
nand U20533 (N_20533,N_20048,N_20055);
nand U20534 (N_20534,N_20151,N_20115);
nand U20535 (N_20535,N_20172,N_20010);
xor U20536 (N_20536,N_20380,N_20294);
nand U20537 (N_20537,N_20213,N_20226);
and U20538 (N_20538,N_20101,N_20064);
nand U20539 (N_20539,N_20001,N_20317);
nor U20540 (N_20540,N_20121,N_20155);
xor U20541 (N_20541,N_20359,N_20429);
or U20542 (N_20542,N_20022,N_20417);
xor U20543 (N_20543,N_20039,N_20241);
nor U20544 (N_20544,N_20025,N_20339);
nand U20545 (N_20545,N_20144,N_20409);
xor U20546 (N_20546,N_20480,N_20234);
nor U20547 (N_20547,N_20427,N_20364);
or U20548 (N_20548,N_20251,N_20303);
or U20549 (N_20549,N_20170,N_20072);
nor U20550 (N_20550,N_20413,N_20095);
xnor U20551 (N_20551,N_20470,N_20104);
or U20552 (N_20552,N_20011,N_20227);
and U20553 (N_20553,N_20200,N_20035);
nor U20554 (N_20554,N_20476,N_20231);
and U20555 (N_20555,N_20062,N_20085);
xnor U20556 (N_20556,N_20154,N_20166);
and U20557 (N_20557,N_20441,N_20183);
nand U20558 (N_20558,N_20327,N_20240);
nor U20559 (N_20559,N_20366,N_20335);
or U20560 (N_20560,N_20206,N_20045);
nand U20561 (N_20561,N_20391,N_20132);
and U20562 (N_20562,N_20471,N_20450);
nand U20563 (N_20563,N_20308,N_20447);
nand U20564 (N_20564,N_20275,N_20322);
xor U20565 (N_20565,N_20415,N_20345);
nand U20566 (N_20566,N_20149,N_20021);
nor U20567 (N_20567,N_20147,N_20081);
xnor U20568 (N_20568,N_20245,N_20473);
xnor U20569 (N_20569,N_20032,N_20000);
nor U20570 (N_20570,N_20495,N_20168);
or U20571 (N_20571,N_20203,N_20173);
xnor U20572 (N_20572,N_20467,N_20018);
nor U20573 (N_20573,N_20434,N_20400);
nor U20574 (N_20574,N_20067,N_20185);
nand U20575 (N_20575,N_20086,N_20188);
or U20576 (N_20576,N_20351,N_20233);
nand U20577 (N_20577,N_20182,N_20131);
xor U20578 (N_20578,N_20316,N_20134);
nor U20579 (N_20579,N_20389,N_20133);
nor U20580 (N_20580,N_20029,N_20099);
xor U20581 (N_20581,N_20264,N_20463);
nand U20582 (N_20582,N_20209,N_20293);
nor U20583 (N_20583,N_20207,N_20255);
and U20584 (N_20584,N_20199,N_20286);
nor U20585 (N_20585,N_20088,N_20406);
nor U20586 (N_20586,N_20248,N_20421);
nor U20587 (N_20587,N_20423,N_20157);
and U20588 (N_20588,N_20334,N_20091);
nor U20589 (N_20589,N_20337,N_20443);
nor U20590 (N_20590,N_20260,N_20020);
or U20591 (N_20591,N_20354,N_20432);
xnor U20592 (N_20592,N_20060,N_20033);
nor U20593 (N_20593,N_20279,N_20028);
xnor U20594 (N_20594,N_20374,N_20385);
or U20595 (N_20595,N_20365,N_20336);
nand U20596 (N_20596,N_20224,N_20216);
nand U20597 (N_20597,N_20023,N_20093);
nor U20598 (N_20598,N_20363,N_20490);
or U20599 (N_20599,N_20098,N_20120);
xnor U20600 (N_20600,N_20475,N_20258);
and U20601 (N_20601,N_20263,N_20092);
or U20602 (N_20602,N_20247,N_20462);
nand U20603 (N_20603,N_20261,N_20356);
and U20604 (N_20604,N_20311,N_20304);
or U20605 (N_20605,N_20269,N_20482);
xor U20606 (N_20606,N_20461,N_20041);
or U20607 (N_20607,N_20497,N_20422);
or U20608 (N_20608,N_20012,N_20280);
nand U20609 (N_20609,N_20487,N_20418);
and U20610 (N_20610,N_20070,N_20175);
and U20611 (N_20611,N_20464,N_20139);
nor U20612 (N_20612,N_20319,N_20158);
or U20613 (N_20613,N_20488,N_20436);
nor U20614 (N_20614,N_20469,N_20333);
and U20615 (N_20615,N_20369,N_20315);
nor U20616 (N_20616,N_20438,N_20014);
nor U20617 (N_20617,N_20071,N_20402);
nor U20618 (N_20618,N_20448,N_20005);
or U20619 (N_20619,N_20061,N_20003);
or U20620 (N_20620,N_20358,N_20007);
xnor U20621 (N_20621,N_20375,N_20455);
and U20622 (N_20622,N_20355,N_20494);
nand U20623 (N_20623,N_20118,N_20050);
nand U20624 (N_20624,N_20320,N_20282);
nor U20625 (N_20625,N_20449,N_20426);
and U20626 (N_20626,N_20352,N_20357);
or U20627 (N_20627,N_20368,N_20287);
and U20628 (N_20628,N_20186,N_20177);
or U20629 (N_20629,N_20405,N_20338);
nor U20630 (N_20630,N_20223,N_20178);
or U20631 (N_20631,N_20326,N_20127);
nand U20632 (N_20632,N_20410,N_20306);
or U20633 (N_20633,N_20034,N_20420);
xnor U20634 (N_20634,N_20198,N_20340);
and U20635 (N_20635,N_20274,N_20344);
or U20636 (N_20636,N_20056,N_20190);
nand U20637 (N_20637,N_20217,N_20110);
or U20638 (N_20638,N_20411,N_20004);
and U20639 (N_20639,N_20431,N_20196);
or U20640 (N_20640,N_20075,N_20367);
or U20641 (N_20641,N_20250,N_20277);
nor U20642 (N_20642,N_20499,N_20452);
xor U20643 (N_20643,N_20194,N_20458);
and U20644 (N_20644,N_20205,N_20016);
nor U20645 (N_20645,N_20243,N_20270);
nor U20646 (N_20646,N_20135,N_20312);
xor U20647 (N_20647,N_20387,N_20396);
xnor U20648 (N_20648,N_20299,N_20083);
or U20649 (N_20649,N_20219,N_20384);
or U20650 (N_20650,N_20446,N_20257);
nor U20651 (N_20651,N_20314,N_20065);
nor U20652 (N_20652,N_20237,N_20297);
or U20653 (N_20653,N_20002,N_20047);
and U20654 (N_20654,N_20136,N_20407);
and U20655 (N_20655,N_20161,N_20030);
and U20656 (N_20656,N_20378,N_20038);
or U20657 (N_20657,N_20109,N_20042);
or U20658 (N_20658,N_20301,N_20281);
and U20659 (N_20659,N_20078,N_20302);
nor U20660 (N_20660,N_20341,N_20232);
nand U20661 (N_20661,N_20453,N_20040);
nand U20662 (N_20662,N_20459,N_20013);
and U20663 (N_20663,N_20063,N_20419);
nor U20664 (N_20664,N_20360,N_20201);
or U20665 (N_20665,N_20361,N_20372);
and U20666 (N_20666,N_20371,N_20235);
xor U20667 (N_20667,N_20124,N_20031);
nor U20668 (N_20668,N_20433,N_20254);
or U20669 (N_20669,N_20179,N_20090);
or U20670 (N_20670,N_20238,N_20265);
nor U20671 (N_20671,N_20017,N_20498);
xor U20672 (N_20672,N_20171,N_20230);
or U20673 (N_20673,N_20310,N_20496);
nor U20674 (N_20674,N_20285,N_20324);
or U20675 (N_20675,N_20159,N_20383);
nand U20676 (N_20676,N_20424,N_20152);
and U20677 (N_20677,N_20457,N_20142);
xor U20678 (N_20678,N_20451,N_20444);
or U20679 (N_20679,N_20259,N_20370);
or U20680 (N_20680,N_20298,N_20215);
and U20681 (N_20681,N_20197,N_20466);
nor U20682 (N_20682,N_20276,N_20309);
xor U20683 (N_20683,N_20126,N_20395);
nor U20684 (N_20684,N_20489,N_20008);
xnor U20685 (N_20685,N_20478,N_20165);
or U20686 (N_20686,N_20140,N_20037);
or U20687 (N_20687,N_20468,N_20330);
nand U20688 (N_20688,N_20493,N_20208);
and U20689 (N_20689,N_20331,N_20465);
and U20690 (N_20690,N_20350,N_20388);
xor U20691 (N_20691,N_20210,N_20289);
or U20692 (N_20692,N_20105,N_20348);
and U20693 (N_20693,N_20439,N_20347);
xnor U20694 (N_20694,N_20068,N_20454);
nor U20695 (N_20695,N_20256,N_20332);
xnor U20696 (N_20696,N_20492,N_20145);
nor U20697 (N_20697,N_20416,N_20146);
and U20698 (N_20698,N_20195,N_20343);
or U20699 (N_20699,N_20346,N_20398);
xnor U20700 (N_20700,N_20024,N_20321);
nor U20701 (N_20701,N_20288,N_20403);
and U20702 (N_20702,N_20009,N_20376);
and U20703 (N_20703,N_20043,N_20362);
nor U20704 (N_20704,N_20049,N_20394);
or U20705 (N_20705,N_20112,N_20381);
and U20706 (N_20706,N_20329,N_20082);
or U20707 (N_20707,N_20036,N_20106);
nor U20708 (N_20708,N_20221,N_20204);
xnor U20709 (N_20709,N_20382,N_20271);
and U20710 (N_20710,N_20076,N_20485);
xor U20711 (N_20711,N_20295,N_20044);
and U20712 (N_20712,N_20117,N_20100);
or U20713 (N_20713,N_20218,N_20202);
nor U20714 (N_20714,N_20267,N_20184);
nor U20715 (N_20715,N_20027,N_20253);
xnor U20716 (N_20716,N_20080,N_20239);
nand U20717 (N_20717,N_20481,N_20486);
nand U20718 (N_20718,N_20108,N_20390);
nand U20719 (N_20719,N_20328,N_20225);
or U20720 (N_20720,N_20052,N_20353);
nor U20721 (N_20721,N_20474,N_20305);
and U20722 (N_20722,N_20440,N_20181);
nand U20723 (N_20723,N_20404,N_20435);
nand U20724 (N_20724,N_20006,N_20244);
nor U20725 (N_20725,N_20483,N_20278);
nor U20726 (N_20726,N_20059,N_20162);
xor U20727 (N_20727,N_20114,N_20015);
xor U20728 (N_20728,N_20193,N_20191);
nor U20729 (N_20729,N_20313,N_20160);
xnor U20730 (N_20730,N_20053,N_20484);
nor U20731 (N_20731,N_20019,N_20266);
nor U20732 (N_20732,N_20442,N_20107);
or U20733 (N_20733,N_20472,N_20491);
xor U20734 (N_20734,N_20097,N_20386);
nand U20735 (N_20735,N_20102,N_20307);
nor U20736 (N_20736,N_20084,N_20393);
nand U20737 (N_20737,N_20236,N_20087);
or U20738 (N_20738,N_20292,N_20057);
or U20739 (N_20739,N_20153,N_20089);
and U20740 (N_20740,N_20456,N_20073);
nand U20741 (N_20741,N_20460,N_20414);
and U20742 (N_20742,N_20349,N_20058);
nor U20743 (N_20743,N_20445,N_20066);
xor U20744 (N_20744,N_20111,N_20125);
and U20745 (N_20745,N_20164,N_20325);
nand U20746 (N_20746,N_20113,N_20079);
nor U20747 (N_20747,N_20323,N_20296);
and U20748 (N_20748,N_20401,N_20122);
xnor U20749 (N_20749,N_20214,N_20143);
or U20750 (N_20750,N_20105,N_20427);
and U20751 (N_20751,N_20080,N_20493);
or U20752 (N_20752,N_20443,N_20126);
nand U20753 (N_20753,N_20100,N_20238);
xor U20754 (N_20754,N_20469,N_20061);
nor U20755 (N_20755,N_20443,N_20380);
or U20756 (N_20756,N_20266,N_20219);
and U20757 (N_20757,N_20160,N_20217);
xnor U20758 (N_20758,N_20471,N_20219);
and U20759 (N_20759,N_20189,N_20214);
nor U20760 (N_20760,N_20189,N_20278);
xnor U20761 (N_20761,N_20384,N_20011);
nor U20762 (N_20762,N_20492,N_20204);
or U20763 (N_20763,N_20369,N_20417);
xnor U20764 (N_20764,N_20216,N_20424);
xnor U20765 (N_20765,N_20098,N_20312);
nand U20766 (N_20766,N_20458,N_20219);
nand U20767 (N_20767,N_20098,N_20248);
and U20768 (N_20768,N_20292,N_20209);
and U20769 (N_20769,N_20161,N_20162);
nor U20770 (N_20770,N_20202,N_20027);
nor U20771 (N_20771,N_20304,N_20379);
nor U20772 (N_20772,N_20392,N_20436);
or U20773 (N_20773,N_20477,N_20006);
xnor U20774 (N_20774,N_20309,N_20399);
nor U20775 (N_20775,N_20340,N_20310);
xor U20776 (N_20776,N_20358,N_20479);
and U20777 (N_20777,N_20393,N_20193);
xor U20778 (N_20778,N_20108,N_20142);
nand U20779 (N_20779,N_20081,N_20365);
nor U20780 (N_20780,N_20286,N_20249);
nor U20781 (N_20781,N_20033,N_20045);
or U20782 (N_20782,N_20102,N_20339);
and U20783 (N_20783,N_20094,N_20446);
and U20784 (N_20784,N_20050,N_20103);
xor U20785 (N_20785,N_20180,N_20182);
nor U20786 (N_20786,N_20163,N_20181);
xnor U20787 (N_20787,N_20361,N_20299);
xnor U20788 (N_20788,N_20410,N_20492);
xnor U20789 (N_20789,N_20388,N_20340);
nand U20790 (N_20790,N_20395,N_20483);
nand U20791 (N_20791,N_20272,N_20153);
and U20792 (N_20792,N_20457,N_20270);
nor U20793 (N_20793,N_20224,N_20295);
or U20794 (N_20794,N_20286,N_20207);
xnor U20795 (N_20795,N_20151,N_20316);
and U20796 (N_20796,N_20474,N_20214);
nand U20797 (N_20797,N_20160,N_20203);
nor U20798 (N_20798,N_20044,N_20299);
nand U20799 (N_20799,N_20051,N_20040);
and U20800 (N_20800,N_20497,N_20384);
nand U20801 (N_20801,N_20224,N_20075);
or U20802 (N_20802,N_20305,N_20329);
or U20803 (N_20803,N_20361,N_20069);
nand U20804 (N_20804,N_20267,N_20120);
or U20805 (N_20805,N_20352,N_20134);
nand U20806 (N_20806,N_20032,N_20075);
nor U20807 (N_20807,N_20063,N_20422);
nand U20808 (N_20808,N_20265,N_20125);
nor U20809 (N_20809,N_20286,N_20430);
xnor U20810 (N_20810,N_20301,N_20002);
and U20811 (N_20811,N_20158,N_20162);
and U20812 (N_20812,N_20418,N_20485);
nand U20813 (N_20813,N_20212,N_20457);
and U20814 (N_20814,N_20202,N_20050);
or U20815 (N_20815,N_20241,N_20042);
and U20816 (N_20816,N_20233,N_20190);
or U20817 (N_20817,N_20326,N_20342);
nor U20818 (N_20818,N_20202,N_20320);
xnor U20819 (N_20819,N_20052,N_20013);
nand U20820 (N_20820,N_20156,N_20231);
nor U20821 (N_20821,N_20326,N_20035);
xnor U20822 (N_20822,N_20053,N_20379);
or U20823 (N_20823,N_20318,N_20425);
xnor U20824 (N_20824,N_20248,N_20396);
and U20825 (N_20825,N_20277,N_20398);
and U20826 (N_20826,N_20030,N_20271);
and U20827 (N_20827,N_20270,N_20067);
nor U20828 (N_20828,N_20206,N_20384);
nand U20829 (N_20829,N_20105,N_20093);
or U20830 (N_20830,N_20307,N_20133);
or U20831 (N_20831,N_20344,N_20119);
xnor U20832 (N_20832,N_20327,N_20059);
and U20833 (N_20833,N_20285,N_20343);
or U20834 (N_20834,N_20257,N_20036);
xnor U20835 (N_20835,N_20306,N_20439);
or U20836 (N_20836,N_20239,N_20253);
or U20837 (N_20837,N_20278,N_20057);
xor U20838 (N_20838,N_20051,N_20444);
nor U20839 (N_20839,N_20426,N_20173);
or U20840 (N_20840,N_20383,N_20234);
nor U20841 (N_20841,N_20253,N_20481);
nand U20842 (N_20842,N_20210,N_20124);
nand U20843 (N_20843,N_20382,N_20199);
or U20844 (N_20844,N_20362,N_20086);
and U20845 (N_20845,N_20404,N_20473);
or U20846 (N_20846,N_20274,N_20120);
nand U20847 (N_20847,N_20272,N_20217);
nand U20848 (N_20848,N_20454,N_20456);
nor U20849 (N_20849,N_20016,N_20209);
and U20850 (N_20850,N_20415,N_20201);
nor U20851 (N_20851,N_20237,N_20348);
nand U20852 (N_20852,N_20077,N_20079);
and U20853 (N_20853,N_20067,N_20266);
nand U20854 (N_20854,N_20382,N_20166);
or U20855 (N_20855,N_20264,N_20289);
or U20856 (N_20856,N_20255,N_20304);
nand U20857 (N_20857,N_20368,N_20124);
xnor U20858 (N_20858,N_20157,N_20458);
and U20859 (N_20859,N_20220,N_20226);
nor U20860 (N_20860,N_20092,N_20446);
or U20861 (N_20861,N_20304,N_20404);
xnor U20862 (N_20862,N_20143,N_20320);
xnor U20863 (N_20863,N_20107,N_20333);
and U20864 (N_20864,N_20073,N_20120);
xor U20865 (N_20865,N_20157,N_20411);
nand U20866 (N_20866,N_20442,N_20056);
and U20867 (N_20867,N_20437,N_20053);
nand U20868 (N_20868,N_20335,N_20351);
or U20869 (N_20869,N_20217,N_20093);
nand U20870 (N_20870,N_20362,N_20058);
nor U20871 (N_20871,N_20020,N_20068);
or U20872 (N_20872,N_20345,N_20150);
nor U20873 (N_20873,N_20047,N_20499);
nand U20874 (N_20874,N_20280,N_20080);
xnor U20875 (N_20875,N_20469,N_20435);
and U20876 (N_20876,N_20412,N_20470);
and U20877 (N_20877,N_20316,N_20382);
and U20878 (N_20878,N_20476,N_20337);
nor U20879 (N_20879,N_20209,N_20017);
or U20880 (N_20880,N_20124,N_20299);
xor U20881 (N_20881,N_20011,N_20041);
nor U20882 (N_20882,N_20454,N_20092);
xor U20883 (N_20883,N_20302,N_20104);
nor U20884 (N_20884,N_20418,N_20384);
nor U20885 (N_20885,N_20319,N_20475);
nand U20886 (N_20886,N_20486,N_20033);
and U20887 (N_20887,N_20078,N_20160);
or U20888 (N_20888,N_20312,N_20119);
xnor U20889 (N_20889,N_20317,N_20048);
xor U20890 (N_20890,N_20375,N_20079);
and U20891 (N_20891,N_20484,N_20493);
or U20892 (N_20892,N_20079,N_20388);
and U20893 (N_20893,N_20373,N_20124);
xor U20894 (N_20894,N_20369,N_20017);
and U20895 (N_20895,N_20368,N_20191);
nand U20896 (N_20896,N_20428,N_20431);
nor U20897 (N_20897,N_20318,N_20485);
or U20898 (N_20898,N_20307,N_20078);
nand U20899 (N_20899,N_20088,N_20157);
nand U20900 (N_20900,N_20045,N_20180);
xor U20901 (N_20901,N_20450,N_20493);
nor U20902 (N_20902,N_20474,N_20134);
xor U20903 (N_20903,N_20306,N_20277);
nor U20904 (N_20904,N_20363,N_20144);
and U20905 (N_20905,N_20388,N_20433);
and U20906 (N_20906,N_20154,N_20151);
nor U20907 (N_20907,N_20111,N_20273);
nand U20908 (N_20908,N_20481,N_20032);
nand U20909 (N_20909,N_20413,N_20112);
or U20910 (N_20910,N_20478,N_20226);
or U20911 (N_20911,N_20188,N_20322);
or U20912 (N_20912,N_20094,N_20317);
nand U20913 (N_20913,N_20159,N_20034);
xnor U20914 (N_20914,N_20489,N_20042);
or U20915 (N_20915,N_20088,N_20387);
xor U20916 (N_20916,N_20463,N_20065);
nor U20917 (N_20917,N_20353,N_20073);
xor U20918 (N_20918,N_20029,N_20103);
nand U20919 (N_20919,N_20476,N_20091);
nor U20920 (N_20920,N_20335,N_20287);
nor U20921 (N_20921,N_20042,N_20046);
or U20922 (N_20922,N_20423,N_20237);
xor U20923 (N_20923,N_20387,N_20005);
or U20924 (N_20924,N_20015,N_20480);
or U20925 (N_20925,N_20303,N_20465);
nor U20926 (N_20926,N_20159,N_20180);
or U20927 (N_20927,N_20398,N_20143);
and U20928 (N_20928,N_20491,N_20259);
xor U20929 (N_20929,N_20128,N_20217);
or U20930 (N_20930,N_20089,N_20302);
nand U20931 (N_20931,N_20083,N_20062);
nand U20932 (N_20932,N_20189,N_20394);
nor U20933 (N_20933,N_20273,N_20427);
nor U20934 (N_20934,N_20073,N_20266);
xnor U20935 (N_20935,N_20438,N_20202);
xnor U20936 (N_20936,N_20390,N_20418);
or U20937 (N_20937,N_20361,N_20283);
nand U20938 (N_20938,N_20168,N_20088);
xor U20939 (N_20939,N_20032,N_20127);
and U20940 (N_20940,N_20214,N_20097);
or U20941 (N_20941,N_20146,N_20411);
and U20942 (N_20942,N_20129,N_20459);
nand U20943 (N_20943,N_20459,N_20348);
xor U20944 (N_20944,N_20082,N_20066);
nand U20945 (N_20945,N_20015,N_20016);
xor U20946 (N_20946,N_20080,N_20351);
nor U20947 (N_20947,N_20287,N_20406);
xnor U20948 (N_20948,N_20076,N_20373);
nand U20949 (N_20949,N_20273,N_20434);
xor U20950 (N_20950,N_20276,N_20057);
nand U20951 (N_20951,N_20068,N_20084);
and U20952 (N_20952,N_20430,N_20171);
nor U20953 (N_20953,N_20409,N_20213);
or U20954 (N_20954,N_20454,N_20180);
xor U20955 (N_20955,N_20227,N_20000);
or U20956 (N_20956,N_20487,N_20370);
and U20957 (N_20957,N_20327,N_20155);
nor U20958 (N_20958,N_20021,N_20461);
xor U20959 (N_20959,N_20389,N_20373);
and U20960 (N_20960,N_20017,N_20458);
or U20961 (N_20961,N_20057,N_20064);
nor U20962 (N_20962,N_20391,N_20336);
nor U20963 (N_20963,N_20232,N_20056);
xor U20964 (N_20964,N_20383,N_20434);
xor U20965 (N_20965,N_20279,N_20154);
and U20966 (N_20966,N_20175,N_20291);
nand U20967 (N_20967,N_20131,N_20373);
xnor U20968 (N_20968,N_20483,N_20021);
or U20969 (N_20969,N_20417,N_20228);
and U20970 (N_20970,N_20140,N_20299);
nand U20971 (N_20971,N_20471,N_20160);
nor U20972 (N_20972,N_20269,N_20271);
xor U20973 (N_20973,N_20375,N_20430);
nor U20974 (N_20974,N_20338,N_20171);
nand U20975 (N_20975,N_20350,N_20136);
nor U20976 (N_20976,N_20455,N_20313);
nand U20977 (N_20977,N_20313,N_20411);
and U20978 (N_20978,N_20353,N_20261);
xnor U20979 (N_20979,N_20183,N_20498);
nor U20980 (N_20980,N_20183,N_20060);
or U20981 (N_20981,N_20458,N_20299);
nor U20982 (N_20982,N_20120,N_20042);
or U20983 (N_20983,N_20184,N_20023);
or U20984 (N_20984,N_20102,N_20219);
xor U20985 (N_20985,N_20122,N_20011);
nor U20986 (N_20986,N_20086,N_20396);
nand U20987 (N_20987,N_20479,N_20292);
nor U20988 (N_20988,N_20379,N_20130);
nor U20989 (N_20989,N_20051,N_20302);
xor U20990 (N_20990,N_20096,N_20381);
xor U20991 (N_20991,N_20058,N_20475);
nand U20992 (N_20992,N_20352,N_20448);
nor U20993 (N_20993,N_20215,N_20297);
nor U20994 (N_20994,N_20359,N_20352);
nor U20995 (N_20995,N_20354,N_20006);
xor U20996 (N_20996,N_20010,N_20044);
nor U20997 (N_20997,N_20062,N_20004);
and U20998 (N_20998,N_20371,N_20296);
nand U20999 (N_20999,N_20261,N_20336);
or U21000 (N_21000,N_20984,N_20720);
nor U21001 (N_21001,N_20834,N_20937);
nand U21002 (N_21002,N_20796,N_20963);
or U21003 (N_21003,N_20759,N_20610);
nor U21004 (N_21004,N_20560,N_20953);
nor U21005 (N_21005,N_20525,N_20865);
or U21006 (N_21006,N_20848,N_20593);
nor U21007 (N_21007,N_20800,N_20678);
xor U21008 (N_21008,N_20816,N_20840);
and U21009 (N_21009,N_20779,N_20641);
nor U21010 (N_21010,N_20620,N_20773);
or U21011 (N_21011,N_20512,N_20889);
xor U21012 (N_21012,N_20944,N_20867);
nor U21013 (N_21013,N_20942,N_20938);
nand U21014 (N_21014,N_20813,N_20544);
nor U21015 (N_21015,N_20915,N_20957);
or U21016 (N_21016,N_20814,N_20740);
xnor U21017 (N_21017,N_20661,N_20973);
nand U21018 (N_21018,N_20896,N_20507);
and U21019 (N_21019,N_20885,N_20844);
nand U21020 (N_21020,N_20968,N_20851);
nor U21021 (N_21021,N_20836,N_20835);
and U21022 (N_21022,N_20529,N_20586);
xnor U21023 (N_21023,N_20989,N_20786);
xor U21024 (N_21024,N_20781,N_20683);
or U21025 (N_21025,N_20501,N_20563);
and U21026 (N_21026,N_20760,N_20613);
or U21027 (N_21027,N_20907,N_20695);
xor U21028 (N_21028,N_20662,N_20684);
or U21029 (N_21029,N_20673,N_20991);
or U21030 (N_21030,N_20746,N_20862);
xor U21031 (N_21031,N_20802,N_20723);
xnor U21032 (N_21032,N_20932,N_20928);
nor U21033 (N_21033,N_20546,N_20743);
xor U21034 (N_21034,N_20993,N_20561);
nor U21035 (N_21035,N_20667,N_20839);
nor U21036 (N_21036,N_20705,N_20841);
and U21037 (N_21037,N_20628,N_20599);
nand U21038 (N_21038,N_20863,N_20821);
nand U21039 (N_21039,N_20846,N_20579);
xor U21040 (N_21040,N_20888,N_20564);
or U21041 (N_21041,N_20543,N_20549);
and U21042 (N_21042,N_20726,N_20995);
nor U21043 (N_21043,N_20539,N_20556);
or U21044 (N_21044,N_20765,N_20569);
or U21045 (N_21045,N_20734,N_20985);
or U21046 (N_21046,N_20858,N_20671);
xnor U21047 (N_21047,N_20633,N_20807);
xnor U21048 (N_21048,N_20890,N_20905);
and U21049 (N_21049,N_20595,N_20847);
nor U21050 (N_21050,N_20693,N_20606);
and U21051 (N_21051,N_20589,N_20541);
and U21052 (N_21052,N_20535,N_20715);
xnor U21053 (N_21053,N_20506,N_20689);
xnor U21054 (N_21054,N_20598,N_20670);
and U21055 (N_21055,N_20675,N_20604);
or U21056 (N_21056,N_20513,N_20892);
nor U21057 (N_21057,N_20755,N_20536);
or U21058 (N_21058,N_20645,N_20592);
and U21059 (N_21059,N_20990,N_20769);
and U21060 (N_21060,N_20766,N_20660);
xor U21061 (N_21061,N_20524,N_20774);
nor U21062 (N_21062,N_20902,N_20698);
xnor U21063 (N_21063,N_20971,N_20584);
nand U21064 (N_21064,N_20980,N_20624);
nor U21065 (N_21065,N_20502,N_20988);
nor U21066 (N_21066,N_20917,N_20653);
nor U21067 (N_21067,N_20987,N_20580);
or U21068 (N_21068,N_20934,N_20571);
nand U21069 (N_21069,N_20871,N_20866);
and U21070 (N_21070,N_20679,N_20597);
xnor U21071 (N_21071,N_20655,N_20951);
or U21072 (N_21072,N_20916,N_20767);
xor U21073 (N_21073,N_20758,N_20808);
nor U21074 (N_21074,N_20964,N_20837);
nand U21075 (N_21075,N_20665,N_20982);
xor U21076 (N_21076,N_20614,N_20946);
xnor U21077 (N_21077,N_20656,N_20643);
and U21078 (N_21078,N_20815,N_20911);
and U21079 (N_21079,N_20729,N_20674);
and U21080 (N_21080,N_20966,N_20873);
xnor U21081 (N_21081,N_20623,N_20828);
or U21082 (N_21082,N_20714,N_20898);
nand U21083 (N_21083,N_20687,N_20859);
nor U21084 (N_21084,N_20882,N_20702);
xnor U21085 (N_21085,N_20831,N_20538);
and U21086 (N_21086,N_20733,N_20799);
nor U21087 (N_21087,N_20562,N_20872);
or U21088 (N_21088,N_20742,N_20797);
nand U21089 (N_21089,N_20621,N_20752);
xor U21090 (N_21090,N_20912,N_20756);
nor U21091 (N_21091,N_20757,N_20850);
nor U21092 (N_21092,N_20568,N_20778);
or U21093 (N_21093,N_20857,N_20792);
and U21094 (N_21094,N_20876,N_20974);
and U21095 (N_21095,N_20651,N_20978);
xor U21096 (N_21096,N_20554,N_20777);
or U21097 (N_21097,N_20860,N_20735);
and U21098 (N_21098,N_20567,N_20939);
or U21099 (N_21099,N_20886,N_20631);
nand U21100 (N_21100,N_20578,N_20545);
xor U21101 (N_21101,N_20776,N_20878);
xor U21102 (N_21102,N_20530,N_20639);
nand U21103 (N_21103,N_20790,N_20534);
or U21104 (N_21104,N_20772,N_20764);
or U21105 (N_21105,N_20607,N_20899);
xnor U21106 (N_21106,N_20503,N_20869);
nor U21107 (N_21107,N_20969,N_20587);
nand U21108 (N_21108,N_20558,N_20708);
and U21109 (N_21109,N_20956,N_20926);
xnor U21110 (N_21110,N_20591,N_20677);
nor U21111 (N_21111,N_20547,N_20787);
nor U21112 (N_21112,N_20832,N_20699);
nor U21113 (N_21113,N_20718,N_20706);
nand U21114 (N_21114,N_20703,N_20798);
or U21115 (N_21115,N_20642,N_20897);
nor U21116 (N_21116,N_20945,N_20812);
and U21117 (N_21117,N_20793,N_20527);
nor U21118 (N_21118,N_20504,N_20602);
nor U21119 (N_21119,N_20717,N_20618);
xnor U21120 (N_21120,N_20895,N_20998);
or U21121 (N_21121,N_20914,N_20842);
nor U21122 (N_21122,N_20811,N_20780);
xnor U21123 (N_21123,N_20685,N_20694);
xnor U21124 (N_21124,N_20819,N_20979);
or U21125 (N_21125,N_20919,N_20972);
nor U21126 (N_21126,N_20716,N_20731);
or U21127 (N_21127,N_20853,N_20994);
nor U21128 (N_21128,N_20958,N_20596);
and U21129 (N_21129,N_20965,N_20906);
xor U21130 (N_21130,N_20627,N_20881);
and U21131 (N_21131,N_20738,N_20970);
xnor U21132 (N_21132,N_20644,N_20728);
nand U21133 (N_21133,N_20801,N_20654);
xor U21134 (N_21134,N_20789,N_20500);
nor U21135 (N_21135,N_20913,N_20657);
xnor U21136 (N_21136,N_20936,N_20721);
nand U21137 (N_21137,N_20747,N_20508);
nand U21138 (N_21138,N_20894,N_20634);
and U21139 (N_21139,N_20625,N_20852);
nor U21140 (N_21140,N_20696,N_20712);
and U21141 (N_21141,N_20555,N_20730);
nor U21142 (N_21142,N_20635,N_20553);
and U21143 (N_21143,N_20523,N_20537);
xnor U21144 (N_21144,N_20891,N_20818);
xor U21145 (N_21145,N_20750,N_20929);
nor U21146 (N_21146,N_20952,N_20823);
and U21147 (N_21147,N_20532,N_20600);
and U21148 (N_21148,N_20880,N_20804);
and U21149 (N_21149,N_20672,N_20719);
nand U21150 (N_21150,N_20548,N_20868);
xnor U21151 (N_21151,N_20576,N_20638);
or U21152 (N_21152,N_20650,N_20954);
nor U21153 (N_21153,N_20725,N_20825);
nand U21154 (N_21154,N_20557,N_20877);
and U21155 (N_21155,N_20551,N_20583);
nor U21156 (N_21156,N_20515,N_20961);
or U21157 (N_21157,N_20820,N_20609);
xor U21158 (N_21158,N_20676,N_20710);
nor U21159 (N_21159,N_20552,N_20783);
nor U21160 (N_21160,N_20603,N_20887);
nand U21161 (N_21161,N_20658,N_20707);
nand U21162 (N_21162,N_20540,N_20574);
nor U21163 (N_21163,N_20533,N_20771);
and U21164 (N_21164,N_20615,N_20668);
or U21165 (N_21165,N_20565,N_20724);
nor U21166 (N_21166,N_20741,N_20893);
or U21167 (N_21167,N_20577,N_20843);
nand U21168 (N_21168,N_20690,N_20788);
or U21169 (N_21169,N_20748,N_20550);
nand U21170 (N_21170,N_20856,N_20739);
nand U21171 (N_21171,N_20521,N_20999);
nor U21172 (N_21172,N_20997,N_20646);
nand U21173 (N_21173,N_20900,N_20763);
and U21174 (N_21174,N_20669,N_20727);
xnor U21175 (N_21175,N_20903,N_20824);
nand U21176 (N_21176,N_20795,N_20516);
and U21177 (N_21177,N_20930,N_20977);
nand U21178 (N_21178,N_20622,N_20955);
xnor U21179 (N_21179,N_20617,N_20870);
and U21180 (N_21180,N_20570,N_20700);
nand U21181 (N_21181,N_20509,N_20948);
xnor U21182 (N_21182,N_20585,N_20967);
and U21183 (N_21183,N_20829,N_20879);
nor U21184 (N_21184,N_20518,N_20809);
nor U21185 (N_21185,N_20682,N_20761);
nand U21186 (N_21186,N_20616,N_20680);
nand U21187 (N_21187,N_20573,N_20861);
xnor U21188 (N_21188,N_20590,N_20983);
nand U21189 (N_21189,N_20572,N_20612);
nand U21190 (N_21190,N_20782,N_20663);
nand U21191 (N_21191,N_20925,N_20962);
and U21192 (N_21192,N_20753,N_20827);
nand U21193 (N_21193,N_20745,N_20519);
and U21194 (N_21194,N_20806,N_20935);
xor U21195 (N_21195,N_20950,N_20611);
or U21196 (N_21196,N_20659,N_20691);
nand U21197 (N_21197,N_20947,N_20652);
or U21198 (N_21198,N_20921,N_20751);
or U21199 (N_21199,N_20686,N_20855);
and U21200 (N_21200,N_20522,N_20531);
nand U21201 (N_21201,N_20601,N_20854);
nor U21202 (N_21202,N_20864,N_20826);
and U21203 (N_21203,N_20732,N_20838);
nand U21204 (N_21204,N_20701,N_20908);
xnor U21205 (N_21205,N_20647,N_20830);
or U21206 (N_21206,N_20940,N_20975);
nand U21207 (N_21207,N_20528,N_20636);
or U21208 (N_21208,N_20666,N_20649);
or U21209 (N_21209,N_20931,N_20664);
xor U21210 (N_21210,N_20514,N_20817);
xnor U21211 (N_21211,N_20632,N_20630);
and U21212 (N_21212,N_20608,N_20909);
nand U21213 (N_21213,N_20960,N_20736);
and U21214 (N_21214,N_20637,N_20805);
nand U21215 (N_21215,N_20505,N_20692);
xnor U21216 (N_21216,N_20594,N_20629);
nor U21217 (N_21217,N_20688,N_20833);
or U21218 (N_21218,N_20922,N_20784);
nor U21219 (N_21219,N_20575,N_20711);
xnor U21220 (N_21220,N_20981,N_20775);
and U21221 (N_21221,N_20910,N_20883);
and U21222 (N_21222,N_20697,N_20648);
or U21223 (N_21223,N_20992,N_20822);
and U21224 (N_21224,N_20996,N_20875);
nor U21225 (N_21225,N_20794,N_20874);
xnor U21226 (N_21226,N_20754,N_20520);
and U21227 (N_21227,N_20927,N_20722);
xnor U21228 (N_21228,N_20884,N_20933);
nor U21229 (N_21229,N_20959,N_20619);
xnor U21230 (N_21230,N_20681,N_20713);
and U21231 (N_21231,N_20749,N_20920);
or U21232 (N_21232,N_20923,N_20949);
xor U21233 (N_21233,N_20640,N_20904);
nor U21234 (N_21234,N_20976,N_20768);
nand U21235 (N_21235,N_20542,N_20810);
or U21236 (N_21236,N_20924,N_20918);
and U21237 (N_21237,N_20588,N_20791);
or U21238 (N_21238,N_20803,N_20901);
nor U21239 (N_21239,N_20709,N_20845);
and U21240 (N_21240,N_20704,N_20737);
nand U21241 (N_21241,N_20566,N_20785);
or U21242 (N_21242,N_20582,N_20511);
xor U21243 (N_21243,N_20762,N_20744);
nand U21244 (N_21244,N_20849,N_20770);
xor U21245 (N_21245,N_20510,N_20626);
xnor U21246 (N_21246,N_20559,N_20526);
nand U21247 (N_21247,N_20943,N_20581);
and U21248 (N_21248,N_20941,N_20605);
nand U21249 (N_21249,N_20986,N_20517);
xor U21250 (N_21250,N_20973,N_20605);
or U21251 (N_21251,N_20516,N_20596);
xnor U21252 (N_21252,N_20756,N_20652);
or U21253 (N_21253,N_20500,N_20661);
xor U21254 (N_21254,N_20866,N_20674);
and U21255 (N_21255,N_20667,N_20736);
nor U21256 (N_21256,N_20693,N_20508);
and U21257 (N_21257,N_20519,N_20984);
xnor U21258 (N_21258,N_20605,N_20771);
nor U21259 (N_21259,N_20762,N_20842);
and U21260 (N_21260,N_20521,N_20908);
xnor U21261 (N_21261,N_20841,N_20554);
nand U21262 (N_21262,N_20696,N_20785);
and U21263 (N_21263,N_20621,N_20802);
xnor U21264 (N_21264,N_20896,N_20940);
nand U21265 (N_21265,N_20632,N_20968);
xor U21266 (N_21266,N_20849,N_20631);
and U21267 (N_21267,N_20941,N_20889);
xnor U21268 (N_21268,N_20613,N_20912);
xnor U21269 (N_21269,N_20581,N_20738);
nor U21270 (N_21270,N_20802,N_20862);
nand U21271 (N_21271,N_20875,N_20723);
or U21272 (N_21272,N_20890,N_20622);
nor U21273 (N_21273,N_20663,N_20847);
nor U21274 (N_21274,N_20549,N_20848);
or U21275 (N_21275,N_20558,N_20655);
and U21276 (N_21276,N_20939,N_20748);
or U21277 (N_21277,N_20873,N_20596);
and U21278 (N_21278,N_20639,N_20763);
nand U21279 (N_21279,N_20665,N_20669);
nor U21280 (N_21280,N_20608,N_20866);
nor U21281 (N_21281,N_20930,N_20881);
and U21282 (N_21282,N_20634,N_20829);
nand U21283 (N_21283,N_20543,N_20614);
or U21284 (N_21284,N_20698,N_20908);
or U21285 (N_21285,N_20921,N_20576);
and U21286 (N_21286,N_20814,N_20793);
xor U21287 (N_21287,N_20538,N_20640);
nand U21288 (N_21288,N_20803,N_20511);
nand U21289 (N_21289,N_20624,N_20671);
xor U21290 (N_21290,N_20723,N_20848);
or U21291 (N_21291,N_20571,N_20989);
and U21292 (N_21292,N_20796,N_20731);
xnor U21293 (N_21293,N_20815,N_20977);
or U21294 (N_21294,N_20525,N_20983);
nor U21295 (N_21295,N_20520,N_20837);
nand U21296 (N_21296,N_20908,N_20660);
xor U21297 (N_21297,N_20882,N_20829);
or U21298 (N_21298,N_20766,N_20518);
and U21299 (N_21299,N_20629,N_20687);
or U21300 (N_21300,N_20921,N_20897);
nor U21301 (N_21301,N_20693,N_20809);
nor U21302 (N_21302,N_20690,N_20937);
or U21303 (N_21303,N_20726,N_20840);
or U21304 (N_21304,N_20558,N_20600);
and U21305 (N_21305,N_20809,N_20850);
nor U21306 (N_21306,N_20879,N_20831);
nand U21307 (N_21307,N_20764,N_20946);
or U21308 (N_21308,N_20810,N_20879);
or U21309 (N_21309,N_20907,N_20518);
or U21310 (N_21310,N_20508,N_20986);
and U21311 (N_21311,N_20672,N_20527);
xor U21312 (N_21312,N_20744,N_20960);
and U21313 (N_21313,N_20836,N_20772);
nor U21314 (N_21314,N_20594,N_20515);
xnor U21315 (N_21315,N_20657,N_20964);
and U21316 (N_21316,N_20900,N_20797);
nand U21317 (N_21317,N_20779,N_20766);
or U21318 (N_21318,N_20802,N_20899);
xnor U21319 (N_21319,N_20645,N_20671);
xnor U21320 (N_21320,N_20551,N_20733);
xor U21321 (N_21321,N_20878,N_20672);
nor U21322 (N_21322,N_20525,N_20871);
nand U21323 (N_21323,N_20847,N_20709);
nor U21324 (N_21324,N_20935,N_20690);
or U21325 (N_21325,N_20721,N_20649);
or U21326 (N_21326,N_20633,N_20560);
xor U21327 (N_21327,N_20707,N_20995);
xor U21328 (N_21328,N_20648,N_20808);
nor U21329 (N_21329,N_20645,N_20908);
and U21330 (N_21330,N_20979,N_20680);
and U21331 (N_21331,N_20558,N_20837);
xor U21332 (N_21332,N_20729,N_20896);
nor U21333 (N_21333,N_20847,N_20650);
or U21334 (N_21334,N_20619,N_20627);
xor U21335 (N_21335,N_20631,N_20594);
or U21336 (N_21336,N_20904,N_20623);
or U21337 (N_21337,N_20965,N_20866);
and U21338 (N_21338,N_20542,N_20820);
xnor U21339 (N_21339,N_20929,N_20777);
and U21340 (N_21340,N_20510,N_20516);
and U21341 (N_21341,N_20534,N_20900);
nor U21342 (N_21342,N_20565,N_20532);
nor U21343 (N_21343,N_20753,N_20781);
or U21344 (N_21344,N_20959,N_20943);
nor U21345 (N_21345,N_20549,N_20599);
nand U21346 (N_21346,N_20760,N_20784);
nand U21347 (N_21347,N_20554,N_20636);
nor U21348 (N_21348,N_20673,N_20835);
nand U21349 (N_21349,N_20962,N_20941);
nand U21350 (N_21350,N_20718,N_20582);
xor U21351 (N_21351,N_20861,N_20511);
xor U21352 (N_21352,N_20643,N_20869);
xnor U21353 (N_21353,N_20510,N_20976);
or U21354 (N_21354,N_20704,N_20925);
nand U21355 (N_21355,N_20756,N_20741);
nor U21356 (N_21356,N_20587,N_20895);
nand U21357 (N_21357,N_20922,N_20905);
nand U21358 (N_21358,N_20625,N_20646);
or U21359 (N_21359,N_20811,N_20799);
nand U21360 (N_21360,N_20559,N_20606);
xnor U21361 (N_21361,N_20567,N_20989);
xnor U21362 (N_21362,N_20566,N_20810);
nand U21363 (N_21363,N_20973,N_20640);
nand U21364 (N_21364,N_20504,N_20546);
xor U21365 (N_21365,N_20934,N_20728);
or U21366 (N_21366,N_20746,N_20967);
nand U21367 (N_21367,N_20980,N_20930);
xor U21368 (N_21368,N_20631,N_20791);
nor U21369 (N_21369,N_20951,N_20760);
nor U21370 (N_21370,N_20695,N_20733);
nand U21371 (N_21371,N_20670,N_20699);
nor U21372 (N_21372,N_20510,N_20881);
or U21373 (N_21373,N_20537,N_20528);
nor U21374 (N_21374,N_20607,N_20615);
and U21375 (N_21375,N_20587,N_20576);
xnor U21376 (N_21376,N_20564,N_20851);
xor U21377 (N_21377,N_20933,N_20557);
or U21378 (N_21378,N_20585,N_20534);
xnor U21379 (N_21379,N_20638,N_20921);
or U21380 (N_21380,N_20849,N_20782);
and U21381 (N_21381,N_20644,N_20755);
nor U21382 (N_21382,N_20982,N_20729);
or U21383 (N_21383,N_20796,N_20851);
or U21384 (N_21384,N_20555,N_20823);
nor U21385 (N_21385,N_20997,N_20896);
xor U21386 (N_21386,N_20885,N_20905);
or U21387 (N_21387,N_20856,N_20722);
nor U21388 (N_21388,N_20633,N_20973);
and U21389 (N_21389,N_20589,N_20774);
nor U21390 (N_21390,N_20751,N_20845);
or U21391 (N_21391,N_20684,N_20933);
nor U21392 (N_21392,N_20904,N_20867);
nand U21393 (N_21393,N_20622,N_20917);
xnor U21394 (N_21394,N_20500,N_20833);
and U21395 (N_21395,N_20739,N_20773);
nor U21396 (N_21396,N_20941,N_20788);
nor U21397 (N_21397,N_20723,N_20957);
nor U21398 (N_21398,N_20510,N_20686);
nand U21399 (N_21399,N_20722,N_20600);
nand U21400 (N_21400,N_20768,N_20812);
nand U21401 (N_21401,N_20961,N_20868);
and U21402 (N_21402,N_20772,N_20563);
and U21403 (N_21403,N_20919,N_20948);
nor U21404 (N_21404,N_20745,N_20661);
or U21405 (N_21405,N_20544,N_20739);
xnor U21406 (N_21406,N_20836,N_20695);
nor U21407 (N_21407,N_20554,N_20585);
nand U21408 (N_21408,N_20775,N_20644);
nor U21409 (N_21409,N_20758,N_20589);
xnor U21410 (N_21410,N_20992,N_20915);
or U21411 (N_21411,N_20594,N_20778);
nor U21412 (N_21412,N_20983,N_20899);
xor U21413 (N_21413,N_20509,N_20801);
and U21414 (N_21414,N_20791,N_20556);
or U21415 (N_21415,N_20655,N_20989);
and U21416 (N_21416,N_20609,N_20730);
nand U21417 (N_21417,N_20626,N_20787);
xor U21418 (N_21418,N_20983,N_20663);
and U21419 (N_21419,N_20501,N_20922);
nor U21420 (N_21420,N_20547,N_20832);
nand U21421 (N_21421,N_20784,N_20947);
nor U21422 (N_21422,N_20892,N_20518);
nor U21423 (N_21423,N_20644,N_20590);
xnor U21424 (N_21424,N_20851,N_20809);
nand U21425 (N_21425,N_20859,N_20531);
or U21426 (N_21426,N_20910,N_20833);
or U21427 (N_21427,N_20753,N_20680);
or U21428 (N_21428,N_20970,N_20898);
xor U21429 (N_21429,N_20861,N_20994);
nand U21430 (N_21430,N_20764,N_20628);
and U21431 (N_21431,N_20892,N_20568);
nand U21432 (N_21432,N_20504,N_20974);
or U21433 (N_21433,N_20632,N_20871);
and U21434 (N_21434,N_20712,N_20719);
or U21435 (N_21435,N_20578,N_20539);
xnor U21436 (N_21436,N_20717,N_20867);
and U21437 (N_21437,N_20540,N_20954);
and U21438 (N_21438,N_20839,N_20683);
nand U21439 (N_21439,N_20720,N_20830);
xnor U21440 (N_21440,N_20682,N_20566);
xnor U21441 (N_21441,N_20969,N_20555);
nor U21442 (N_21442,N_20784,N_20842);
nor U21443 (N_21443,N_20565,N_20778);
nand U21444 (N_21444,N_20565,N_20999);
nand U21445 (N_21445,N_20765,N_20971);
xnor U21446 (N_21446,N_20963,N_20530);
nand U21447 (N_21447,N_20610,N_20920);
nor U21448 (N_21448,N_20693,N_20585);
or U21449 (N_21449,N_20749,N_20592);
and U21450 (N_21450,N_20537,N_20572);
xor U21451 (N_21451,N_20731,N_20795);
xor U21452 (N_21452,N_20968,N_20975);
nand U21453 (N_21453,N_20751,N_20877);
or U21454 (N_21454,N_20783,N_20838);
nand U21455 (N_21455,N_20629,N_20765);
xnor U21456 (N_21456,N_20822,N_20643);
and U21457 (N_21457,N_20828,N_20621);
nand U21458 (N_21458,N_20960,N_20578);
nand U21459 (N_21459,N_20505,N_20874);
xnor U21460 (N_21460,N_20700,N_20580);
nor U21461 (N_21461,N_20557,N_20999);
or U21462 (N_21462,N_20938,N_20863);
or U21463 (N_21463,N_20569,N_20576);
nor U21464 (N_21464,N_20924,N_20693);
or U21465 (N_21465,N_20706,N_20589);
xnor U21466 (N_21466,N_20615,N_20989);
nor U21467 (N_21467,N_20995,N_20538);
nor U21468 (N_21468,N_20595,N_20919);
and U21469 (N_21469,N_20527,N_20947);
xor U21470 (N_21470,N_20845,N_20589);
xor U21471 (N_21471,N_20804,N_20596);
and U21472 (N_21472,N_20506,N_20954);
and U21473 (N_21473,N_20555,N_20619);
nand U21474 (N_21474,N_20940,N_20966);
xnor U21475 (N_21475,N_20729,N_20857);
or U21476 (N_21476,N_20658,N_20746);
or U21477 (N_21477,N_20975,N_20805);
xnor U21478 (N_21478,N_20998,N_20778);
nand U21479 (N_21479,N_20982,N_20642);
nand U21480 (N_21480,N_20570,N_20521);
nor U21481 (N_21481,N_20854,N_20584);
nor U21482 (N_21482,N_20693,N_20900);
nand U21483 (N_21483,N_20668,N_20808);
nor U21484 (N_21484,N_20663,N_20855);
or U21485 (N_21485,N_20978,N_20739);
nor U21486 (N_21486,N_20638,N_20816);
nor U21487 (N_21487,N_20989,N_20930);
or U21488 (N_21488,N_20761,N_20818);
nor U21489 (N_21489,N_20786,N_20519);
xor U21490 (N_21490,N_20784,N_20568);
xor U21491 (N_21491,N_20600,N_20959);
and U21492 (N_21492,N_20895,N_20855);
nand U21493 (N_21493,N_20764,N_20553);
xnor U21494 (N_21494,N_20647,N_20995);
or U21495 (N_21495,N_20863,N_20700);
and U21496 (N_21496,N_20550,N_20852);
or U21497 (N_21497,N_20603,N_20914);
and U21498 (N_21498,N_20595,N_20835);
nor U21499 (N_21499,N_20702,N_20896);
xnor U21500 (N_21500,N_21152,N_21159);
and U21501 (N_21501,N_21435,N_21222);
xnor U21502 (N_21502,N_21119,N_21232);
nand U21503 (N_21503,N_21493,N_21038);
nand U21504 (N_21504,N_21291,N_21490);
xor U21505 (N_21505,N_21123,N_21132);
nor U21506 (N_21506,N_21498,N_21207);
and U21507 (N_21507,N_21323,N_21486);
xor U21508 (N_21508,N_21220,N_21299);
nand U21509 (N_21509,N_21289,N_21464);
xor U21510 (N_21510,N_21225,N_21111);
nor U21511 (N_21511,N_21445,N_21063);
nor U21512 (N_21512,N_21437,N_21474);
and U21513 (N_21513,N_21124,N_21240);
xor U21514 (N_21514,N_21480,N_21359);
and U21515 (N_21515,N_21326,N_21004);
xor U21516 (N_21516,N_21272,N_21044);
xnor U21517 (N_21517,N_21042,N_21354);
nor U21518 (N_21518,N_21250,N_21165);
nor U21519 (N_21519,N_21430,N_21116);
nor U21520 (N_21520,N_21341,N_21355);
or U21521 (N_21521,N_21115,N_21134);
nor U21522 (N_21522,N_21372,N_21174);
nor U21523 (N_21523,N_21153,N_21495);
or U21524 (N_21524,N_21452,N_21127);
or U21525 (N_21525,N_21425,N_21060);
and U21526 (N_21526,N_21315,N_21343);
nand U21527 (N_21527,N_21394,N_21158);
xnor U21528 (N_21528,N_21109,N_21345);
nor U21529 (N_21529,N_21252,N_21410);
or U21530 (N_21530,N_21338,N_21460);
nor U21531 (N_21531,N_21030,N_21236);
and U21532 (N_21532,N_21344,N_21039);
or U21533 (N_21533,N_21096,N_21121);
nand U21534 (N_21534,N_21277,N_21125);
or U21535 (N_21535,N_21010,N_21237);
xor U21536 (N_21536,N_21456,N_21247);
xnor U21537 (N_21537,N_21248,N_21189);
nand U21538 (N_21538,N_21377,N_21018);
nor U21539 (N_21539,N_21251,N_21228);
nand U21540 (N_21540,N_21477,N_21012);
xor U21541 (N_21541,N_21069,N_21316);
nor U21542 (N_21542,N_21328,N_21348);
xor U21543 (N_21543,N_21330,N_21293);
xnor U21544 (N_21544,N_21395,N_21214);
nor U21545 (N_21545,N_21317,N_21133);
or U21546 (N_21546,N_21131,N_21478);
or U21547 (N_21547,N_21310,N_21161);
or U21548 (N_21548,N_21409,N_21156);
xnor U21549 (N_21549,N_21282,N_21298);
or U21550 (N_21550,N_21249,N_21319);
and U21551 (N_21551,N_21450,N_21365);
and U21552 (N_21552,N_21385,N_21446);
or U21553 (N_21553,N_21184,N_21302);
nand U21554 (N_21554,N_21485,N_21349);
xor U21555 (N_21555,N_21138,N_21175);
nand U21556 (N_21556,N_21095,N_21431);
or U21557 (N_21557,N_21001,N_21101);
xor U21558 (N_21558,N_21139,N_21283);
nand U21559 (N_21559,N_21339,N_21126);
or U21560 (N_21560,N_21242,N_21389);
nand U21561 (N_21561,N_21122,N_21466);
xnor U21562 (N_21562,N_21255,N_21254);
or U21563 (N_21563,N_21489,N_21337);
and U21564 (N_21564,N_21306,N_21419);
xnor U21565 (N_21565,N_21029,N_21241);
and U21566 (N_21566,N_21180,N_21288);
or U21567 (N_21567,N_21427,N_21086);
nor U21568 (N_21568,N_21443,N_21128);
and U21569 (N_21569,N_21032,N_21370);
and U21570 (N_21570,N_21108,N_21142);
xnor U21571 (N_21571,N_21265,N_21083);
or U21572 (N_21572,N_21366,N_21084);
nor U21573 (N_21573,N_21280,N_21428);
or U21574 (N_21574,N_21401,N_21157);
nand U21575 (N_21575,N_21393,N_21423);
xor U21576 (N_21576,N_21488,N_21217);
or U21577 (N_21577,N_21226,N_21424);
and U21578 (N_21578,N_21433,N_21364);
and U21579 (N_21579,N_21303,N_21335);
nor U21580 (N_21580,N_21403,N_21301);
nor U21581 (N_21581,N_21259,N_21376);
or U21582 (N_21582,N_21104,N_21453);
and U21583 (N_21583,N_21448,N_21218);
or U21584 (N_21584,N_21494,N_21094);
nand U21585 (N_21585,N_21099,N_21285);
nand U21586 (N_21586,N_21369,N_21047);
nor U21587 (N_21587,N_21244,N_21422);
and U21588 (N_21588,N_21455,N_21268);
and U21589 (N_21589,N_21002,N_21262);
nor U21590 (N_21590,N_21374,N_21173);
nor U21591 (N_21591,N_21320,N_21404);
and U21592 (N_21592,N_21151,N_21442);
and U21593 (N_21593,N_21436,N_21253);
nor U21594 (N_21594,N_21210,N_21353);
xor U21595 (N_21595,N_21150,N_21076);
or U21596 (N_21596,N_21266,N_21072);
xor U21597 (N_21597,N_21487,N_21234);
nor U21598 (N_21598,N_21304,N_21264);
xnor U21599 (N_21599,N_21491,N_21311);
nand U21600 (N_21600,N_21073,N_21162);
xor U21601 (N_21601,N_21013,N_21065);
nor U21602 (N_21602,N_21031,N_21213);
nand U21603 (N_21603,N_21022,N_21235);
xnor U21604 (N_21604,N_21273,N_21190);
or U21605 (N_21605,N_21281,N_21429);
and U21606 (N_21606,N_21467,N_21172);
and U21607 (N_21607,N_21106,N_21198);
nand U21608 (N_21608,N_21271,N_21239);
nor U21609 (N_21609,N_21463,N_21003);
nor U21610 (N_21610,N_21492,N_21066);
nor U21611 (N_21611,N_21392,N_21461);
nor U21612 (N_21612,N_21459,N_21102);
nand U21613 (N_21613,N_21384,N_21155);
nor U21614 (N_21614,N_21118,N_21347);
or U21615 (N_21615,N_21140,N_21078);
and U21616 (N_21616,N_21089,N_21054);
and U21617 (N_21617,N_21308,N_21256);
xnor U21618 (N_21618,N_21465,N_21216);
nor U21619 (N_21619,N_21048,N_21414);
nand U21620 (N_21620,N_21499,N_21143);
and U21621 (N_21621,N_21219,N_21110);
and U21622 (N_21622,N_21411,N_21027);
and U21623 (N_21623,N_21211,N_21011);
nor U21624 (N_21624,N_21041,N_21399);
nand U21625 (N_21625,N_21398,N_21071);
and U21626 (N_21626,N_21396,N_21373);
or U21627 (N_21627,N_21274,N_21188);
nor U21628 (N_21628,N_21313,N_21473);
nand U21629 (N_21629,N_21238,N_21176);
nor U21630 (N_21630,N_21482,N_21449);
nand U21631 (N_21631,N_21019,N_21154);
and U21632 (N_21632,N_21357,N_21201);
and U21633 (N_21633,N_21245,N_21382);
nand U21634 (N_21634,N_21405,N_21196);
nor U21635 (N_21635,N_21352,N_21481);
and U21636 (N_21636,N_21020,N_21203);
nand U21637 (N_21637,N_21215,N_21426);
nor U21638 (N_21638,N_21340,N_21168);
nor U21639 (N_21639,N_21278,N_21120);
xnor U21640 (N_21640,N_21160,N_21136);
or U21641 (N_21641,N_21324,N_21199);
and U21642 (N_21642,N_21105,N_21223);
xnor U21643 (N_21643,N_21185,N_21141);
xor U21644 (N_21644,N_21439,N_21447);
and U21645 (N_21645,N_21387,N_21418);
xor U21646 (N_21646,N_21087,N_21053);
or U21647 (N_21647,N_21043,N_21358);
nand U21648 (N_21648,N_21227,N_21021);
or U21649 (N_21649,N_21451,N_21112);
and U21650 (N_21650,N_21193,N_21014);
and U21651 (N_21651,N_21181,N_21009);
nor U21652 (N_21652,N_21375,N_21017);
nor U21653 (N_21653,N_21434,N_21100);
nor U21654 (N_21654,N_21284,N_21050);
nor U21655 (N_21655,N_21381,N_21200);
nor U21656 (N_21656,N_21476,N_21224);
nand U21657 (N_21657,N_21144,N_21148);
and U21658 (N_21658,N_21261,N_21233);
or U21659 (N_21659,N_21279,N_21346);
and U21660 (N_21660,N_21379,N_21270);
nor U21661 (N_21661,N_21321,N_21191);
xnor U21662 (N_21662,N_21186,N_21458);
xor U21663 (N_21663,N_21035,N_21230);
nand U21664 (N_21664,N_21361,N_21322);
or U21665 (N_21665,N_21182,N_21081);
nand U21666 (N_21666,N_21204,N_21077);
nand U21667 (N_21667,N_21107,N_21469);
and U21668 (N_21668,N_21415,N_21468);
xnor U21669 (N_21669,N_21046,N_21049);
nand U21670 (N_21670,N_21070,N_21334);
xor U21671 (N_21671,N_21416,N_21179);
xor U21672 (N_21672,N_21388,N_21195);
or U21673 (N_21673,N_21413,N_21212);
nand U21674 (N_21674,N_21064,N_21292);
xor U21675 (N_21675,N_21332,N_21454);
nand U21676 (N_21676,N_21402,N_21231);
xor U21677 (N_21677,N_21058,N_21462);
nand U21678 (N_21678,N_21300,N_21438);
or U21679 (N_21679,N_21333,N_21135);
xnor U21680 (N_21680,N_21386,N_21483);
or U21681 (N_21681,N_21351,N_21342);
xnor U21682 (N_21682,N_21074,N_21325);
xnor U21683 (N_21683,N_21113,N_21258);
or U21684 (N_21684,N_21097,N_21192);
nor U21685 (N_21685,N_21444,N_21380);
or U21686 (N_21686,N_21079,N_21432);
xor U21687 (N_21687,N_21475,N_21205);
nand U21688 (N_21688,N_21057,N_21229);
nor U21689 (N_21689,N_21059,N_21383);
nand U21690 (N_21690,N_21406,N_21075);
nand U21691 (N_21691,N_21037,N_21412);
xnor U21692 (N_21692,N_21336,N_21296);
or U21693 (N_21693,N_21117,N_21260);
nor U21694 (N_21694,N_21114,N_21331);
xnor U21695 (N_21695,N_21000,N_21497);
or U21696 (N_21696,N_21082,N_21052);
or U21697 (N_21697,N_21098,N_21178);
or U21698 (N_21698,N_21085,N_21441);
xnor U21699 (N_21699,N_21091,N_21257);
nand U21700 (N_21700,N_21350,N_21036);
nand U21701 (N_21701,N_21088,N_21170);
or U21702 (N_21702,N_21479,N_21294);
nor U21703 (N_21703,N_21202,N_21149);
nand U21704 (N_21704,N_21163,N_21305);
or U21705 (N_21705,N_21314,N_21329);
nor U21706 (N_21706,N_21484,N_21177);
or U21707 (N_21707,N_21457,N_21062);
or U21708 (N_21708,N_21033,N_21055);
nand U21709 (N_21709,N_21056,N_21297);
nor U21710 (N_21710,N_21471,N_21040);
nor U21711 (N_21711,N_21061,N_21206);
or U21712 (N_21712,N_21397,N_21015);
nand U21713 (N_21713,N_21051,N_21420);
or U21714 (N_21714,N_21130,N_21145);
xnor U21715 (N_21715,N_21440,N_21187);
and U21716 (N_21716,N_21068,N_21093);
xor U21717 (N_21717,N_21290,N_21008);
and U21718 (N_21718,N_21286,N_21208);
and U21719 (N_21719,N_21391,N_21194);
nor U21720 (N_21720,N_21363,N_21221);
or U21721 (N_21721,N_21243,N_21023);
nand U21722 (N_21722,N_21287,N_21390);
xor U21723 (N_21723,N_21103,N_21312);
and U21724 (N_21724,N_21360,N_21025);
or U21725 (N_21725,N_21309,N_21371);
or U21726 (N_21726,N_21378,N_21092);
nor U21727 (N_21727,N_21356,N_21275);
nand U21728 (N_21728,N_21407,N_21263);
xnor U21729 (N_21729,N_21080,N_21026);
nand U21730 (N_21730,N_21267,N_21318);
nor U21731 (N_21731,N_21024,N_21327);
nand U21732 (N_21732,N_21400,N_21146);
nor U21733 (N_21733,N_21367,N_21183);
nand U21734 (N_21734,N_21269,N_21408);
xor U21735 (N_21735,N_21005,N_21028);
and U21736 (N_21736,N_21417,N_21067);
nand U21737 (N_21737,N_21496,N_21137);
xnor U21738 (N_21738,N_21421,N_21016);
xnor U21739 (N_21739,N_21006,N_21169);
nor U21740 (N_21740,N_21246,N_21147);
or U21741 (N_21741,N_21007,N_21209);
nand U21742 (N_21742,N_21362,N_21276);
or U21743 (N_21743,N_21307,N_21166);
nor U21744 (N_21744,N_21164,N_21197);
nand U21745 (N_21745,N_21129,N_21368);
and U21746 (N_21746,N_21045,N_21034);
or U21747 (N_21747,N_21171,N_21470);
nand U21748 (N_21748,N_21472,N_21090);
xnor U21749 (N_21749,N_21295,N_21167);
nand U21750 (N_21750,N_21127,N_21249);
nor U21751 (N_21751,N_21052,N_21340);
or U21752 (N_21752,N_21375,N_21335);
xnor U21753 (N_21753,N_21351,N_21153);
nor U21754 (N_21754,N_21156,N_21493);
or U21755 (N_21755,N_21188,N_21343);
or U21756 (N_21756,N_21058,N_21416);
xor U21757 (N_21757,N_21258,N_21240);
nand U21758 (N_21758,N_21134,N_21236);
nor U21759 (N_21759,N_21266,N_21107);
xnor U21760 (N_21760,N_21157,N_21301);
and U21761 (N_21761,N_21364,N_21074);
nor U21762 (N_21762,N_21292,N_21300);
nand U21763 (N_21763,N_21035,N_21253);
nand U21764 (N_21764,N_21028,N_21068);
xnor U21765 (N_21765,N_21449,N_21409);
nand U21766 (N_21766,N_21372,N_21203);
nor U21767 (N_21767,N_21307,N_21291);
and U21768 (N_21768,N_21430,N_21300);
nand U21769 (N_21769,N_21358,N_21397);
and U21770 (N_21770,N_21087,N_21403);
nor U21771 (N_21771,N_21286,N_21284);
nand U21772 (N_21772,N_21267,N_21246);
nand U21773 (N_21773,N_21330,N_21201);
or U21774 (N_21774,N_21360,N_21039);
and U21775 (N_21775,N_21009,N_21164);
nor U21776 (N_21776,N_21085,N_21173);
nand U21777 (N_21777,N_21052,N_21408);
nor U21778 (N_21778,N_21429,N_21182);
nand U21779 (N_21779,N_21132,N_21158);
nand U21780 (N_21780,N_21020,N_21183);
xnor U21781 (N_21781,N_21251,N_21070);
nand U21782 (N_21782,N_21222,N_21454);
nand U21783 (N_21783,N_21120,N_21425);
nand U21784 (N_21784,N_21225,N_21114);
and U21785 (N_21785,N_21378,N_21279);
nor U21786 (N_21786,N_21304,N_21409);
xnor U21787 (N_21787,N_21496,N_21138);
xor U21788 (N_21788,N_21028,N_21294);
nand U21789 (N_21789,N_21310,N_21482);
nor U21790 (N_21790,N_21265,N_21484);
nand U21791 (N_21791,N_21250,N_21020);
xor U21792 (N_21792,N_21138,N_21120);
or U21793 (N_21793,N_21497,N_21389);
nor U21794 (N_21794,N_21412,N_21432);
xor U21795 (N_21795,N_21093,N_21250);
nor U21796 (N_21796,N_21473,N_21143);
xor U21797 (N_21797,N_21039,N_21042);
xnor U21798 (N_21798,N_21315,N_21301);
nand U21799 (N_21799,N_21045,N_21449);
and U21800 (N_21800,N_21102,N_21487);
xnor U21801 (N_21801,N_21372,N_21014);
and U21802 (N_21802,N_21428,N_21222);
or U21803 (N_21803,N_21279,N_21216);
nor U21804 (N_21804,N_21222,N_21402);
nand U21805 (N_21805,N_21256,N_21361);
and U21806 (N_21806,N_21399,N_21214);
xnor U21807 (N_21807,N_21460,N_21008);
and U21808 (N_21808,N_21410,N_21460);
and U21809 (N_21809,N_21022,N_21095);
and U21810 (N_21810,N_21428,N_21176);
nand U21811 (N_21811,N_21449,N_21218);
and U21812 (N_21812,N_21003,N_21254);
nor U21813 (N_21813,N_21128,N_21244);
or U21814 (N_21814,N_21431,N_21233);
nor U21815 (N_21815,N_21033,N_21227);
xor U21816 (N_21816,N_21225,N_21493);
or U21817 (N_21817,N_21482,N_21113);
nor U21818 (N_21818,N_21230,N_21288);
or U21819 (N_21819,N_21128,N_21103);
or U21820 (N_21820,N_21022,N_21227);
or U21821 (N_21821,N_21450,N_21318);
nand U21822 (N_21822,N_21477,N_21375);
or U21823 (N_21823,N_21413,N_21283);
or U21824 (N_21824,N_21349,N_21208);
xnor U21825 (N_21825,N_21254,N_21091);
xnor U21826 (N_21826,N_21045,N_21073);
xor U21827 (N_21827,N_21207,N_21041);
and U21828 (N_21828,N_21277,N_21138);
or U21829 (N_21829,N_21018,N_21402);
xnor U21830 (N_21830,N_21320,N_21093);
xor U21831 (N_21831,N_21135,N_21202);
or U21832 (N_21832,N_21427,N_21305);
or U21833 (N_21833,N_21078,N_21361);
nor U21834 (N_21834,N_21104,N_21137);
or U21835 (N_21835,N_21062,N_21450);
nand U21836 (N_21836,N_21130,N_21254);
nand U21837 (N_21837,N_21187,N_21131);
and U21838 (N_21838,N_21310,N_21106);
nand U21839 (N_21839,N_21426,N_21296);
xor U21840 (N_21840,N_21114,N_21385);
and U21841 (N_21841,N_21435,N_21476);
or U21842 (N_21842,N_21256,N_21094);
and U21843 (N_21843,N_21460,N_21092);
nand U21844 (N_21844,N_21487,N_21326);
or U21845 (N_21845,N_21490,N_21043);
nor U21846 (N_21846,N_21065,N_21003);
nand U21847 (N_21847,N_21119,N_21158);
and U21848 (N_21848,N_21291,N_21462);
nand U21849 (N_21849,N_21257,N_21302);
or U21850 (N_21850,N_21286,N_21212);
nor U21851 (N_21851,N_21317,N_21156);
and U21852 (N_21852,N_21263,N_21044);
nand U21853 (N_21853,N_21344,N_21399);
or U21854 (N_21854,N_21307,N_21188);
nor U21855 (N_21855,N_21281,N_21117);
nand U21856 (N_21856,N_21465,N_21235);
nand U21857 (N_21857,N_21292,N_21391);
and U21858 (N_21858,N_21190,N_21426);
nor U21859 (N_21859,N_21347,N_21191);
nor U21860 (N_21860,N_21383,N_21082);
or U21861 (N_21861,N_21390,N_21005);
nor U21862 (N_21862,N_21370,N_21149);
xnor U21863 (N_21863,N_21315,N_21264);
or U21864 (N_21864,N_21003,N_21030);
or U21865 (N_21865,N_21349,N_21109);
and U21866 (N_21866,N_21486,N_21303);
nor U21867 (N_21867,N_21257,N_21244);
nand U21868 (N_21868,N_21043,N_21434);
nand U21869 (N_21869,N_21043,N_21040);
nor U21870 (N_21870,N_21416,N_21066);
nand U21871 (N_21871,N_21303,N_21065);
xnor U21872 (N_21872,N_21421,N_21204);
and U21873 (N_21873,N_21479,N_21145);
nor U21874 (N_21874,N_21252,N_21481);
and U21875 (N_21875,N_21469,N_21060);
nand U21876 (N_21876,N_21098,N_21038);
nor U21877 (N_21877,N_21123,N_21174);
or U21878 (N_21878,N_21210,N_21138);
or U21879 (N_21879,N_21471,N_21433);
nand U21880 (N_21880,N_21033,N_21237);
xnor U21881 (N_21881,N_21351,N_21007);
nand U21882 (N_21882,N_21200,N_21078);
xnor U21883 (N_21883,N_21046,N_21164);
nor U21884 (N_21884,N_21009,N_21326);
nor U21885 (N_21885,N_21336,N_21265);
or U21886 (N_21886,N_21428,N_21023);
nor U21887 (N_21887,N_21429,N_21311);
and U21888 (N_21888,N_21412,N_21294);
or U21889 (N_21889,N_21187,N_21447);
and U21890 (N_21890,N_21487,N_21394);
xnor U21891 (N_21891,N_21214,N_21235);
nand U21892 (N_21892,N_21173,N_21118);
nand U21893 (N_21893,N_21062,N_21311);
and U21894 (N_21894,N_21330,N_21254);
and U21895 (N_21895,N_21367,N_21214);
and U21896 (N_21896,N_21317,N_21053);
xnor U21897 (N_21897,N_21098,N_21165);
nor U21898 (N_21898,N_21245,N_21173);
nor U21899 (N_21899,N_21446,N_21433);
nand U21900 (N_21900,N_21310,N_21238);
nor U21901 (N_21901,N_21109,N_21128);
and U21902 (N_21902,N_21246,N_21151);
or U21903 (N_21903,N_21184,N_21035);
xnor U21904 (N_21904,N_21489,N_21178);
nor U21905 (N_21905,N_21470,N_21358);
nor U21906 (N_21906,N_21472,N_21054);
or U21907 (N_21907,N_21492,N_21167);
xnor U21908 (N_21908,N_21095,N_21422);
xor U21909 (N_21909,N_21305,N_21162);
nand U21910 (N_21910,N_21473,N_21141);
xnor U21911 (N_21911,N_21145,N_21270);
xnor U21912 (N_21912,N_21251,N_21282);
xor U21913 (N_21913,N_21014,N_21218);
nor U21914 (N_21914,N_21383,N_21212);
or U21915 (N_21915,N_21399,N_21180);
nand U21916 (N_21916,N_21260,N_21469);
or U21917 (N_21917,N_21426,N_21455);
nand U21918 (N_21918,N_21294,N_21325);
nor U21919 (N_21919,N_21455,N_21077);
nor U21920 (N_21920,N_21448,N_21205);
and U21921 (N_21921,N_21112,N_21394);
or U21922 (N_21922,N_21051,N_21060);
nand U21923 (N_21923,N_21213,N_21473);
nand U21924 (N_21924,N_21300,N_21073);
and U21925 (N_21925,N_21078,N_21137);
nor U21926 (N_21926,N_21012,N_21085);
nand U21927 (N_21927,N_21255,N_21178);
nand U21928 (N_21928,N_21269,N_21011);
nand U21929 (N_21929,N_21156,N_21191);
xor U21930 (N_21930,N_21321,N_21025);
or U21931 (N_21931,N_21201,N_21244);
and U21932 (N_21932,N_21202,N_21335);
nand U21933 (N_21933,N_21342,N_21002);
or U21934 (N_21934,N_21078,N_21356);
or U21935 (N_21935,N_21410,N_21312);
nand U21936 (N_21936,N_21176,N_21046);
xor U21937 (N_21937,N_21031,N_21186);
xnor U21938 (N_21938,N_21277,N_21059);
and U21939 (N_21939,N_21303,N_21184);
or U21940 (N_21940,N_21112,N_21440);
or U21941 (N_21941,N_21318,N_21245);
or U21942 (N_21942,N_21227,N_21395);
xor U21943 (N_21943,N_21095,N_21427);
or U21944 (N_21944,N_21156,N_21478);
nor U21945 (N_21945,N_21273,N_21102);
or U21946 (N_21946,N_21273,N_21236);
and U21947 (N_21947,N_21487,N_21465);
nor U21948 (N_21948,N_21336,N_21285);
nor U21949 (N_21949,N_21319,N_21416);
or U21950 (N_21950,N_21304,N_21158);
nor U21951 (N_21951,N_21133,N_21181);
nor U21952 (N_21952,N_21290,N_21302);
xor U21953 (N_21953,N_21433,N_21063);
and U21954 (N_21954,N_21047,N_21070);
xor U21955 (N_21955,N_21192,N_21431);
and U21956 (N_21956,N_21435,N_21347);
nand U21957 (N_21957,N_21364,N_21272);
or U21958 (N_21958,N_21197,N_21453);
or U21959 (N_21959,N_21442,N_21311);
and U21960 (N_21960,N_21446,N_21274);
and U21961 (N_21961,N_21129,N_21275);
and U21962 (N_21962,N_21441,N_21231);
and U21963 (N_21963,N_21071,N_21157);
or U21964 (N_21964,N_21149,N_21197);
nor U21965 (N_21965,N_21005,N_21119);
nand U21966 (N_21966,N_21408,N_21092);
and U21967 (N_21967,N_21442,N_21126);
nand U21968 (N_21968,N_21419,N_21368);
and U21969 (N_21969,N_21387,N_21300);
nor U21970 (N_21970,N_21235,N_21053);
or U21971 (N_21971,N_21189,N_21453);
and U21972 (N_21972,N_21107,N_21447);
nand U21973 (N_21973,N_21369,N_21176);
and U21974 (N_21974,N_21106,N_21184);
or U21975 (N_21975,N_21301,N_21046);
or U21976 (N_21976,N_21261,N_21322);
or U21977 (N_21977,N_21497,N_21177);
nor U21978 (N_21978,N_21142,N_21442);
xnor U21979 (N_21979,N_21074,N_21298);
or U21980 (N_21980,N_21146,N_21038);
nand U21981 (N_21981,N_21186,N_21268);
or U21982 (N_21982,N_21203,N_21370);
xnor U21983 (N_21983,N_21378,N_21306);
nor U21984 (N_21984,N_21498,N_21232);
nand U21985 (N_21985,N_21270,N_21415);
or U21986 (N_21986,N_21217,N_21357);
and U21987 (N_21987,N_21135,N_21496);
xor U21988 (N_21988,N_21322,N_21173);
and U21989 (N_21989,N_21390,N_21341);
nor U21990 (N_21990,N_21345,N_21427);
nand U21991 (N_21991,N_21447,N_21463);
or U21992 (N_21992,N_21494,N_21373);
nor U21993 (N_21993,N_21293,N_21022);
and U21994 (N_21994,N_21434,N_21168);
nor U21995 (N_21995,N_21282,N_21019);
nand U21996 (N_21996,N_21132,N_21118);
nand U21997 (N_21997,N_21009,N_21093);
nor U21998 (N_21998,N_21469,N_21274);
xor U21999 (N_21999,N_21056,N_21073);
nand U22000 (N_22000,N_21695,N_21988);
nor U22001 (N_22001,N_21781,N_21849);
and U22002 (N_22002,N_21985,N_21569);
xnor U22003 (N_22003,N_21671,N_21623);
nand U22004 (N_22004,N_21593,N_21798);
and U22005 (N_22005,N_21770,N_21823);
nand U22006 (N_22006,N_21601,N_21506);
xor U22007 (N_22007,N_21940,N_21504);
and U22008 (N_22008,N_21537,N_21804);
xor U22009 (N_22009,N_21766,N_21813);
and U22010 (N_22010,N_21732,N_21711);
nand U22011 (N_22011,N_21657,N_21820);
nand U22012 (N_22012,N_21777,N_21689);
and U22013 (N_22013,N_21598,N_21803);
nor U22014 (N_22014,N_21915,N_21752);
nor U22015 (N_22015,N_21586,N_21546);
xor U22016 (N_22016,N_21670,N_21654);
xor U22017 (N_22017,N_21525,N_21522);
and U22018 (N_22018,N_21523,N_21895);
and U22019 (N_22019,N_21821,N_21790);
nand U22020 (N_22020,N_21636,N_21749);
nor U22021 (N_22021,N_21617,N_21706);
xor U22022 (N_22022,N_21656,N_21958);
and U22023 (N_22023,N_21762,N_21782);
and U22024 (N_22024,N_21805,N_21633);
nand U22025 (N_22025,N_21614,N_21784);
or U22026 (N_22026,N_21727,N_21579);
xor U22027 (N_22027,N_21584,N_21621);
or U22028 (N_22028,N_21610,N_21761);
and U22029 (N_22029,N_21744,N_21792);
nor U22030 (N_22030,N_21622,N_21592);
nor U22031 (N_22031,N_21738,N_21899);
nand U22032 (N_22032,N_21952,N_21716);
or U22033 (N_22033,N_21560,N_21853);
nand U22034 (N_22034,N_21948,N_21669);
and U22035 (N_22035,N_21957,N_21649);
or U22036 (N_22036,N_21624,N_21583);
or U22037 (N_22037,N_21517,N_21839);
nand U22038 (N_22038,N_21759,N_21933);
xnor U22039 (N_22039,N_21665,N_21998);
nand U22040 (N_22040,N_21966,N_21942);
or U22041 (N_22041,N_21551,N_21800);
nand U22042 (N_22042,N_21964,N_21765);
nor U22043 (N_22043,N_21846,N_21529);
and U22044 (N_22044,N_21702,N_21926);
or U22045 (N_22045,N_21904,N_21642);
and U22046 (N_22046,N_21746,N_21745);
xnor U22047 (N_22047,N_21993,N_21709);
nor U22048 (N_22048,N_21989,N_21534);
nor U22049 (N_22049,N_21808,N_21870);
or U22050 (N_22050,N_21995,N_21854);
and U22051 (N_22051,N_21986,N_21514);
nand U22052 (N_22052,N_21660,N_21780);
and U22053 (N_22053,N_21673,N_21550);
and U22054 (N_22054,N_21917,N_21962);
or U22055 (N_22055,N_21838,N_21647);
and U22056 (N_22056,N_21675,N_21729);
nand U22057 (N_22057,N_21739,N_21691);
xnor U22058 (N_22058,N_21783,N_21640);
and U22059 (N_22059,N_21789,N_21811);
nand U22060 (N_22060,N_21965,N_21564);
or U22061 (N_22061,N_21878,N_21518);
nand U22062 (N_22062,N_21877,N_21824);
nor U22063 (N_22063,N_21737,N_21947);
nor U22064 (N_22064,N_21543,N_21644);
nor U22065 (N_22065,N_21686,N_21682);
and U22066 (N_22066,N_21949,N_21704);
nand U22067 (N_22067,N_21502,N_21629);
nand U22068 (N_22068,N_21628,N_21845);
xnor U22069 (N_22069,N_21547,N_21630);
nor U22070 (N_22070,N_21907,N_21521);
nor U22071 (N_22071,N_21725,N_21999);
xor U22072 (N_22072,N_21871,N_21501);
nor U22073 (N_22073,N_21581,N_21977);
xnor U22074 (N_22074,N_21715,N_21832);
nand U22075 (N_22075,N_21724,N_21826);
and U22076 (N_22076,N_21690,N_21748);
nand U22077 (N_22077,N_21578,N_21863);
or U22078 (N_22078,N_21978,N_21574);
xor U22079 (N_22079,N_21902,N_21776);
nor U22080 (N_22080,N_21678,N_21666);
or U22081 (N_22081,N_21646,N_21822);
and U22082 (N_22082,N_21509,N_21857);
nand U22083 (N_22083,N_21896,N_21513);
nand U22084 (N_22084,N_21720,N_21515);
xor U22085 (N_22085,N_21953,N_21990);
or U22086 (N_22086,N_21651,N_21612);
nor U22087 (N_22087,N_21662,N_21874);
and U22088 (N_22088,N_21655,N_21963);
xor U22089 (N_22089,N_21873,N_21950);
and U22090 (N_22090,N_21908,N_21728);
or U22091 (N_22091,N_21680,N_21510);
xor U22092 (N_22092,N_21936,N_21843);
xnor U22093 (N_22093,N_21618,N_21722);
and U22094 (N_22094,N_21733,N_21721);
and U22095 (N_22095,N_21856,N_21809);
xor U22096 (N_22096,N_21836,N_21885);
xnor U22097 (N_22097,N_21992,N_21815);
xnor U22098 (N_22098,N_21603,N_21833);
nand U22099 (N_22099,N_21847,N_21771);
nand U22100 (N_22100,N_21890,N_21553);
or U22101 (N_22101,N_21810,N_21788);
and U22102 (N_22102,N_21735,N_21664);
xor U22103 (N_22103,N_21542,N_21883);
or U22104 (N_22104,N_21982,N_21605);
and U22105 (N_22105,N_21596,N_21956);
nand U22106 (N_22106,N_21507,N_21648);
nor U22107 (N_22107,N_21533,N_21613);
and U22108 (N_22108,N_21774,N_21814);
and U22109 (N_22109,N_21677,N_21723);
xor U22110 (N_22110,N_21793,N_21703);
and U22111 (N_22111,N_21595,N_21884);
and U22112 (N_22112,N_21615,N_21632);
nand U22113 (N_22113,N_21787,N_21922);
or U22114 (N_22114,N_21585,N_21609);
xor U22115 (N_22115,N_21693,N_21566);
or U22116 (N_22116,N_21924,N_21858);
and U22117 (N_22117,N_21627,N_21840);
xnor U22118 (N_22118,N_21747,N_21960);
or U22119 (N_22119,N_21927,N_21616);
and U22120 (N_22120,N_21519,N_21736);
nand U22121 (N_22121,N_21987,N_21663);
xor U22122 (N_22122,N_21503,N_21939);
and U22123 (N_22123,N_21828,N_21945);
or U22124 (N_22124,N_21714,N_21921);
nor U22125 (N_22125,N_21684,N_21549);
nand U22126 (N_22126,N_21882,N_21734);
and U22127 (N_22127,N_21799,N_21687);
or U22128 (N_22128,N_21892,N_21937);
nand U22129 (N_22129,N_21568,N_21559);
nand U22130 (N_22130,N_21713,N_21743);
nand U22131 (N_22131,N_21775,N_21555);
nand U22132 (N_22132,N_21968,N_21554);
and U22133 (N_22133,N_21575,N_21756);
nor U22134 (N_22134,N_21842,N_21637);
nor U22135 (N_22135,N_21768,N_21697);
and U22136 (N_22136,N_21891,N_21900);
xor U22137 (N_22137,N_21699,N_21829);
nor U22138 (N_22138,N_21918,N_21505);
nand U22139 (N_22139,N_21512,N_21719);
or U22140 (N_22140,N_21970,N_21641);
nor U22141 (N_22141,N_21912,N_21692);
and U22142 (N_22142,N_21818,N_21797);
nand U22143 (N_22143,N_21879,N_21886);
nor U22144 (N_22144,N_21528,N_21577);
nand U22145 (N_22145,N_21668,N_21919);
and U22146 (N_22146,N_21876,N_21527);
and U22147 (N_22147,N_21909,N_21597);
xor U22148 (N_22148,N_21520,N_21758);
and U22149 (N_22149,N_21973,N_21866);
xnor U22150 (N_22150,N_21760,N_21994);
nand U22151 (N_22151,N_21700,N_21645);
or U22152 (N_22152,N_21548,N_21631);
or U22153 (N_22153,N_21931,N_21906);
nand U22154 (N_22154,N_21905,N_21976);
xnor U22155 (N_22155,N_21802,N_21865);
nand U22156 (N_22156,N_21591,N_21961);
nand U22157 (N_22157,N_21897,N_21565);
nand U22158 (N_22158,N_21812,N_21932);
nand U22159 (N_22159,N_21619,N_21740);
or U22160 (N_22160,N_21951,N_21830);
and U22161 (N_22161,N_21996,N_21844);
xnor U22162 (N_22162,N_21557,N_21508);
nor U22163 (N_22163,N_21903,N_21753);
nand U22164 (N_22164,N_21571,N_21785);
or U22165 (N_22165,N_21626,N_21667);
nand U22166 (N_22166,N_21587,N_21757);
and U22167 (N_22167,N_21779,N_21954);
and U22168 (N_22168,N_21545,N_21570);
xnor U22169 (N_22169,N_21855,N_21552);
or U22170 (N_22170,N_21825,N_21750);
nor U22171 (N_22171,N_21755,N_21572);
and U22172 (N_22172,N_21698,N_21972);
nand U22173 (N_22173,N_21606,N_21974);
nor U22174 (N_22174,N_21531,N_21764);
nor U22175 (N_22175,N_21635,N_21935);
or U22176 (N_22176,N_21590,N_21535);
nand U22177 (N_22177,N_21837,N_21920);
xnor U22178 (N_22178,N_21582,N_21981);
nand U22179 (N_22179,N_21794,N_21530);
and U22180 (N_22180,N_21742,N_21659);
nor U22181 (N_22181,N_21741,N_21850);
xnor U22182 (N_22182,N_21696,N_21643);
or U22183 (N_22183,N_21588,N_21806);
and U22184 (N_22184,N_21538,N_21589);
or U22185 (N_22185,N_21511,N_21661);
nand U22186 (N_22186,N_21639,N_21763);
or U22187 (N_22187,N_21868,N_21707);
xnor U22188 (N_22188,N_21681,N_21889);
or U22189 (N_22189,N_21791,N_21807);
and U22190 (N_22190,N_21929,N_21767);
or U22191 (N_22191,N_21971,N_21819);
and U22192 (N_22192,N_21928,N_21604);
nand U22193 (N_22193,N_21984,N_21708);
or U22194 (N_22194,N_21731,N_21526);
or U22195 (N_22195,N_21558,N_21524);
nor U22196 (N_22196,N_21946,N_21712);
nor U22197 (N_22197,N_21573,N_21969);
nor U22198 (N_22198,N_21967,N_21869);
or U22199 (N_22199,N_21540,N_21816);
or U22200 (N_22200,N_21923,N_21500);
or U22201 (N_22201,N_21608,N_21852);
xnor U22202 (N_22202,N_21625,N_21599);
nand U22203 (N_22203,N_21683,N_21914);
nand U22204 (N_22204,N_21893,N_21860);
nor U22205 (N_22205,N_21834,N_21718);
or U22206 (N_22206,N_21562,N_21817);
xor U22207 (N_22207,N_21979,N_21862);
xor U22208 (N_22208,N_21769,N_21916);
and U22209 (N_22209,N_21676,N_21930);
and U22210 (N_22210,N_21938,N_21717);
nand U22211 (N_22211,N_21851,N_21679);
xnor U22212 (N_22212,N_21576,N_21959);
or U22213 (N_22213,N_21901,N_21941);
xor U22214 (N_22214,N_21594,N_21872);
and U22215 (N_22215,N_21638,N_21796);
nand U22216 (N_22216,N_21913,N_21772);
nor U22217 (N_22217,N_21795,N_21516);
and U22218 (N_22218,N_21848,N_21867);
nand U22219 (N_22219,N_21880,N_21685);
nand U22220 (N_22220,N_21875,N_21556);
or U22221 (N_22221,N_21634,N_21943);
or U22222 (N_22222,N_21539,N_21580);
or U22223 (N_22223,N_21688,N_21786);
and U22224 (N_22224,N_21652,N_21653);
nor U22225 (N_22225,N_21827,N_21600);
nor U22226 (N_22226,N_21754,N_21650);
or U22227 (N_22227,N_21567,N_21726);
xnor U22228 (N_22228,N_21925,N_21898);
and U22229 (N_22229,N_21955,N_21536);
xnor U22230 (N_22230,N_21563,N_21983);
nand U22231 (N_22231,N_21710,N_21602);
nor U22232 (N_22232,N_21674,N_21801);
nor U22233 (N_22233,N_21730,N_21861);
xnor U22234 (N_22234,N_21773,N_21541);
or U22235 (N_22235,N_21841,N_21532);
nand U22236 (N_22236,N_21975,N_21859);
xnor U22237 (N_22237,N_21997,N_21751);
nor U22238 (N_22238,N_21607,N_21881);
xor U22239 (N_22239,N_21705,N_21778);
and U22240 (N_22240,N_21911,N_21701);
and U22241 (N_22241,N_21888,N_21991);
nand U22242 (N_22242,N_21658,N_21672);
xnor U22243 (N_22243,N_21561,N_21611);
xnor U22244 (N_22244,N_21894,N_21694);
xnor U22245 (N_22245,N_21934,N_21544);
and U22246 (N_22246,N_21864,N_21944);
or U22247 (N_22247,N_21831,N_21910);
nand U22248 (N_22248,N_21980,N_21835);
xor U22249 (N_22249,N_21887,N_21620);
xnor U22250 (N_22250,N_21925,N_21965);
or U22251 (N_22251,N_21620,N_21762);
and U22252 (N_22252,N_21606,N_21873);
xnor U22253 (N_22253,N_21768,N_21856);
xnor U22254 (N_22254,N_21672,N_21846);
nand U22255 (N_22255,N_21889,N_21897);
nand U22256 (N_22256,N_21654,N_21855);
nand U22257 (N_22257,N_21834,N_21926);
and U22258 (N_22258,N_21594,N_21849);
or U22259 (N_22259,N_21751,N_21594);
or U22260 (N_22260,N_21806,N_21934);
xnor U22261 (N_22261,N_21789,N_21899);
or U22262 (N_22262,N_21692,N_21817);
nor U22263 (N_22263,N_21687,N_21541);
and U22264 (N_22264,N_21909,N_21768);
xor U22265 (N_22265,N_21672,N_21579);
and U22266 (N_22266,N_21534,N_21558);
and U22267 (N_22267,N_21830,N_21761);
or U22268 (N_22268,N_21540,N_21544);
xor U22269 (N_22269,N_21539,N_21572);
or U22270 (N_22270,N_21834,N_21602);
or U22271 (N_22271,N_21683,N_21515);
and U22272 (N_22272,N_21997,N_21597);
nor U22273 (N_22273,N_21970,N_21818);
and U22274 (N_22274,N_21577,N_21876);
nor U22275 (N_22275,N_21680,N_21792);
or U22276 (N_22276,N_21692,N_21766);
nor U22277 (N_22277,N_21608,N_21804);
and U22278 (N_22278,N_21615,N_21988);
and U22279 (N_22279,N_21682,N_21835);
or U22280 (N_22280,N_21689,N_21766);
nand U22281 (N_22281,N_21563,N_21935);
or U22282 (N_22282,N_21581,N_21551);
xnor U22283 (N_22283,N_21582,N_21605);
and U22284 (N_22284,N_21938,N_21611);
nand U22285 (N_22285,N_21931,N_21972);
xor U22286 (N_22286,N_21752,N_21542);
and U22287 (N_22287,N_21892,N_21641);
or U22288 (N_22288,N_21920,N_21555);
nor U22289 (N_22289,N_21780,N_21544);
nor U22290 (N_22290,N_21826,N_21838);
xnor U22291 (N_22291,N_21787,N_21503);
nor U22292 (N_22292,N_21761,N_21645);
nor U22293 (N_22293,N_21607,N_21800);
and U22294 (N_22294,N_21961,N_21656);
nand U22295 (N_22295,N_21965,N_21985);
and U22296 (N_22296,N_21920,N_21790);
or U22297 (N_22297,N_21772,N_21699);
or U22298 (N_22298,N_21983,N_21808);
and U22299 (N_22299,N_21907,N_21930);
or U22300 (N_22300,N_21794,N_21954);
and U22301 (N_22301,N_21574,N_21955);
and U22302 (N_22302,N_21896,N_21835);
nand U22303 (N_22303,N_21844,N_21997);
nand U22304 (N_22304,N_21863,N_21541);
nand U22305 (N_22305,N_21945,N_21925);
and U22306 (N_22306,N_21947,N_21912);
xnor U22307 (N_22307,N_21976,N_21930);
or U22308 (N_22308,N_21971,N_21607);
nor U22309 (N_22309,N_21626,N_21923);
or U22310 (N_22310,N_21845,N_21709);
nor U22311 (N_22311,N_21549,N_21595);
nor U22312 (N_22312,N_21626,N_21508);
or U22313 (N_22313,N_21769,N_21931);
and U22314 (N_22314,N_21780,N_21549);
and U22315 (N_22315,N_21529,N_21843);
xor U22316 (N_22316,N_21748,N_21819);
xor U22317 (N_22317,N_21958,N_21861);
nor U22318 (N_22318,N_21943,N_21710);
xor U22319 (N_22319,N_21866,N_21711);
nor U22320 (N_22320,N_21841,N_21966);
nand U22321 (N_22321,N_21676,N_21899);
nor U22322 (N_22322,N_21659,N_21665);
or U22323 (N_22323,N_21922,N_21708);
nor U22324 (N_22324,N_21672,N_21799);
or U22325 (N_22325,N_21512,N_21861);
and U22326 (N_22326,N_21526,N_21707);
nor U22327 (N_22327,N_21523,N_21524);
xor U22328 (N_22328,N_21914,N_21974);
or U22329 (N_22329,N_21959,N_21659);
nand U22330 (N_22330,N_21822,N_21526);
and U22331 (N_22331,N_21948,N_21563);
or U22332 (N_22332,N_21679,N_21546);
nand U22333 (N_22333,N_21641,N_21781);
or U22334 (N_22334,N_21568,N_21511);
or U22335 (N_22335,N_21989,N_21668);
xnor U22336 (N_22336,N_21898,N_21614);
and U22337 (N_22337,N_21901,N_21790);
xor U22338 (N_22338,N_21953,N_21858);
and U22339 (N_22339,N_21769,N_21514);
nor U22340 (N_22340,N_21966,N_21602);
xnor U22341 (N_22341,N_21896,N_21629);
nand U22342 (N_22342,N_21530,N_21556);
nand U22343 (N_22343,N_21544,N_21898);
xnor U22344 (N_22344,N_21915,N_21631);
and U22345 (N_22345,N_21766,N_21841);
nand U22346 (N_22346,N_21943,N_21898);
xnor U22347 (N_22347,N_21879,N_21977);
and U22348 (N_22348,N_21921,N_21609);
nand U22349 (N_22349,N_21642,N_21596);
nor U22350 (N_22350,N_21871,N_21602);
nor U22351 (N_22351,N_21620,N_21963);
and U22352 (N_22352,N_21503,N_21538);
nor U22353 (N_22353,N_21968,N_21945);
nand U22354 (N_22354,N_21600,N_21960);
and U22355 (N_22355,N_21645,N_21832);
xor U22356 (N_22356,N_21777,N_21669);
and U22357 (N_22357,N_21966,N_21712);
nand U22358 (N_22358,N_21986,N_21974);
or U22359 (N_22359,N_21522,N_21932);
nand U22360 (N_22360,N_21557,N_21747);
nand U22361 (N_22361,N_21992,N_21825);
nor U22362 (N_22362,N_21623,N_21591);
nand U22363 (N_22363,N_21856,N_21512);
or U22364 (N_22364,N_21621,N_21727);
or U22365 (N_22365,N_21567,N_21885);
and U22366 (N_22366,N_21659,N_21608);
or U22367 (N_22367,N_21751,N_21526);
nand U22368 (N_22368,N_21904,N_21659);
or U22369 (N_22369,N_21656,N_21614);
and U22370 (N_22370,N_21772,N_21620);
or U22371 (N_22371,N_21776,N_21985);
and U22372 (N_22372,N_21965,N_21665);
xnor U22373 (N_22373,N_21845,N_21924);
xnor U22374 (N_22374,N_21659,N_21973);
or U22375 (N_22375,N_21563,N_21882);
and U22376 (N_22376,N_21752,N_21600);
or U22377 (N_22377,N_21516,N_21804);
xnor U22378 (N_22378,N_21725,N_21791);
or U22379 (N_22379,N_21639,N_21942);
xor U22380 (N_22380,N_21648,N_21517);
nor U22381 (N_22381,N_21609,N_21865);
or U22382 (N_22382,N_21542,N_21531);
and U22383 (N_22383,N_21632,N_21777);
and U22384 (N_22384,N_21863,N_21889);
or U22385 (N_22385,N_21615,N_21993);
or U22386 (N_22386,N_21514,N_21972);
nor U22387 (N_22387,N_21545,N_21791);
nand U22388 (N_22388,N_21935,N_21968);
nand U22389 (N_22389,N_21700,N_21788);
xnor U22390 (N_22390,N_21874,N_21648);
nand U22391 (N_22391,N_21998,N_21882);
nor U22392 (N_22392,N_21627,N_21853);
nand U22393 (N_22393,N_21745,N_21828);
nand U22394 (N_22394,N_21530,N_21843);
xnor U22395 (N_22395,N_21980,N_21633);
or U22396 (N_22396,N_21709,N_21870);
and U22397 (N_22397,N_21883,N_21734);
and U22398 (N_22398,N_21596,N_21566);
nand U22399 (N_22399,N_21587,N_21554);
and U22400 (N_22400,N_21994,N_21627);
and U22401 (N_22401,N_21823,N_21556);
xnor U22402 (N_22402,N_21847,N_21831);
nand U22403 (N_22403,N_21818,N_21744);
nand U22404 (N_22404,N_21850,N_21878);
nor U22405 (N_22405,N_21776,N_21735);
and U22406 (N_22406,N_21917,N_21756);
xnor U22407 (N_22407,N_21716,N_21718);
or U22408 (N_22408,N_21547,N_21758);
nor U22409 (N_22409,N_21762,N_21763);
nor U22410 (N_22410,N_21560,N_21861);
or U22411 (N_22411,N_21651,N_21676);
nor U22412 (N_22412,N_21636,N_21919);
and U22413 (N_22413,N_21682,N_21977);
xnor U22414 (N_22414,N_21719,N_21758);
xnor U22415 (N_22415,N_21995,N_21568);
nor U22416 (N_22416,N_21984,N_21729);
nor U22417 (N_22417,N_21856,N_21752);
or U22418 (N_22418,N_21716,N_21648);
nand U22419 (N_22419,N_21841,N_21937);
and U22420 (N_22420,N_21779,N_21823);
or U22421 (N_22421,N_21986,N_21683);
nand U22422 (N_22422,N_21771,N_21750);
and U22423 (N_22423,N_21955,N_21618);
xnor U22424 (N_22424,N_21661,N_21773);
nor U22425 (N_22425,N_21814,N_21858);
xnor U22426 (N_22426,N_21554,N_21867);
xor U22427 (N_22427,N_21728,N_21565);
or U22428 (N_22428,N_21707,N_21823);
and U22429 (N_22429,N_21877,N_21810);
xnor U22430 (N_22430,N_21970,N_21861);
and U22431 (N_22431,N_21876,N_21657);
xor U22432 (N_22432,N_21664,N_21686);
xnor U22433 (N_22433,N_21868,N_21653);
or U22434 (N_22434,N_21928,N_21508);
and U22435 (N_22435,N_21836,N_21638);
nand U22436 (N_22436,N_21565,N_21572);
xnor U22437 (N_22437,N_21792,N_21583);
or U22438 (N_22438,N_21990,N_21879);
or U22439 (N_22439,N_21608,N_21817);
and U22440 (N_22440,N_21833,N_21898);
xnor U22441 (N_22441,N_21825,N_21983);
and U22442 (N_22442,N_21644,N_21906);
and U22443 (N_22443,N_21870,N_21695);
and U22444 (N_22444,N_21869,N_21848);
xor U22445 (N_22445,N_21934,N_21760);
nand U22446 (N_22446,N_21568,N_21809);
nor U22447 (N_22447,N_21762,N_21839);
and U22448 (N_22448,N_21504,N_21977);
and U22449 (N_22449,N_21870,N_21755);
or U22450 (N_22450,N_21728,N_21588);
or U22451 (N_22451,N_21893,N_21561);
and U22452 (N_22452,N_21644,N_21658);
nand U22453 (N_22453,N_21638,N_21938);
or U22454 (N_22454,N_21588,N_21505);
nor U22455 (N_22455,N_21585,N_21816);
xor U22456 (N_22456,N_21648,N_21533);
nand U22457 (N_22457,N_21944,N_21838);
or U22458 (N_22458,N_21649,N_21513);
and U22459 (N_22459,N_21782,N_21895);
nand U22460 (N_22460,N_21721,N_21977);
or U22461 (N_22461,N_21994,N_21706);
xnor U22462 (N_22462,N_21692,N_21937);
xnor U22463 (N_22463,N_21635,N_21692);
nor U22464 (N_22464,N_21794,N_21652);
nand U22465 (N_22465,N_21923,N_21538);
nor U22466 (N_22466,N_21899,N_21584);
and U22467 (N_22467,N_21689,N_21956);
nor U22468 (N_22468,N_21660,N_21827);
and U22469 (N_22469,N_21617,N_21831);
or U22470 (N_22470,N_21887,N_21789);
xor U22471 (N_22471,N_21616,N_21653);
xor U22472 (N_22472,N_21975,N_21651);
and U22473 (N_22473,N_21915,N_21728);
or U22474 (N_22474,N_21847,N_21613);
nand U22475 (N_22475,N_21846,N_21891);
or U22476 (N_22476,N_21621,N_21768);
nor U22477 (N_22477,N_21996,N_21973);
xor U22478 (N_22478,N_21966,N_21555);
nand U22479 (N_22479,N_21716,N_21789);
and U22480 (N_22480,N_21766,N_21973);
nor U22481 (N_22481,N_21776,N_21502);
nor U22482 (N_22482,N_21890,N_21621);
xor U22483 (N_22483,N_21893,N_21965);
xnor U22484 (N_22484,N_21651,N_21866);
or U22485 (N_22485,N_21923,N_21975);
xnor U22486 (N_22486,N_21848,N_21636);
or U22487 (N_22487,N_21518,N_21891);
or U22488 (N_22488,N_21880,N_21527);
and U22489 (N_22489,N_21561,N_21600);
or U22490 (N_22490,N_21753,N_21500);
xor U22491 (N_22491,N_21548,N_21756);
and U22492 (N_22492,N_21744,N_21905);
nor U22493 (N_22493,N_21578,N_21598);
xnor U22494 (N_22494,N_21703,N_21713);
nand U22495 (N_22495,N_21860,N_21857);
and U22496 (N_22496,N_21745,N_21749);
nand U22497 (N_22497,N_21729,N_21607);
nand U22498 (N_22498,N_21752,N_21812);
xnor U22499 (N_22499,N_21584,N_21998);
or U22500 (N_22500,N_22096,N_22356);
xor U22501 (N_22501,N_22146,N_22056);
nand U22502 (N_22502,N_22270,N_22063);
nand U22503 (N_22503,N_22497,N_22495);
nand U22504 (N_22504,N_22088,N_22354);
nand U22505 (N_22505,N_22084,N_22126);
nor U22506 (N_22506,N_22165,N_22049);
xnor U22507 (N_22507,N_22141,N_22311);
xor U22508 (N_22508,N_22180,N_22136);
nand U22509 (N_22509,N_22100,N_22099);
and U22510 (N_22510,N_22064,N_22125);
nand U22511 (N_22511,N_22259,N_22382);
nand U22512 (N_22512,N_22059,N_22480);
nor U22513 (N_22513,N_22021,N_22150);
xnor U22514 (N_22514,N_22291,N_22144);
xor U22515 (N_22515,N_22229,N_22271);
and U22516 (N_22516,N_22122,N_22415);
nand U22517 (N_22517,N_22357,N_22364);
nand U22518 (N_22518,N_22347,N_22097);
xor U22519 (N_22519,N_22460,N_22381);
nand U22520 (N_22520,N_22411,N_22393);
xnor U22521 (N_22521,N_22250,N_22292);
and U22522 (N_22522,N_22067,N_22029);
nor U22523 (N_22523,N_22009,N_22237);
and U22524 (N_22524,N_22030,N_22418);
or U22525 (N_22525,N_22329,N_22394);
nand U22526 (N_22526,N_22476,N_22251);
or U22527 (N_22527,N_22330,N_22413);
nor U22528 (N_22528,N_22328,N_22098);
nor U22529 (N_22529,N_22026,N_22496);
or U22530 (N_22530,N_22261,N_22082);
and U22531 (N_22531,N_22465,N_22403);
and U22532 (N_22532,N_22396,N_22438);
or U22533 (N_22533,N_22445,N_22074);
and U22534 (N_22534,N_22198,N_22078);
nor U22535 (N_22535,N_22266,N_22265);
nand U22536 (N_22536,N_22231,N_22414);
xnor U22537 (N_22537,N_22194,N_22042);
or U22538 (N_22538,N_22478,N_22297);
nor U22539 (N_22539,N_22316,N_22255);
nand U22540 (N_22540,N_22373,N_22363);
or U22541 (N_22541,N_22213,N_22308);
nor U22542 (N_22542,N_22185,N_22424);
nor U22543 (N_22543,N_22060,N_22370);
or U22544 (N_22544,N_22202,N_22473);
nand U22545 (N_22545,N_22066,N_22075);
nor U22546 (N_22546,N_22129,N_22466);
xor U22547 (N_22547,N_22353,N_22483);
and U22548 (N_22548,N_22436,N_22086);
nand U22549 (N_22549,N_22107,N_22239);
nand U22550 (N_22550,N_22040,N_22208);
nand U22551 (N_22551,N_22215,N_22004);
nor U22552 (N_22552,N_22349,N_22222);
or U22553 (N_22553,N_22022,N_22240);
nand U22554 (N_22554,N_22285,N_22178);
xor U22555 (N_22555,N_22020,N_22391);
nand U22556 (N_22556,N_22196,N_22235);
and U22557 (N_22557,N_22390,N_22015);
and U22558 (N_22558,N_22206,N_22337);
and U22559 (N_22559,N_22041,N_22310);
and U22560 (N_22560,N_22207,N_22453);
and U22561 (N_22561,N_22065,N_22048);
nand U22562 (N_22562,N_22233,N_22128);
and U22563 (N_22563,N_22260,N_22116);
and U22564 (N_22564,N_22085,N_22427);
nand U22565 (N_22565,N_22429,N_22119);
nand U22566 (N_22566,N_22158,N_22102);
nand U22567 (N_22567,N_22105,N_22169);
nor U22568 (N_22568,N_22450,N_22053);
nand U22569 (N_22569,N_22317,N_22159);
and U22570 (N_22570,N_22012,N_22286);
or U22571 (N_22571,N_22149,N_22431);
and U22572 (N_22572,N_22033,N_22225);
nand U22573 (N_22573,N_22117,N_22127);
nand U22574 (N_22574,N_22220,N_22470);
and U22575 (N_22575,N_22204,N_22135);
or U22576 (N_22576,N_22183,N_22481);
xor U22577 (N_22577,N_22156,N_22341);
nand U22578 (N_22578,N_22134,N_22050);
nand U22579 (N_22579,N_22314,N_22210);
or U22580 (N_22580,N_22428,N_22492);
nor U22581 (N_22581,N_22167,N_22008);
nor U22582 (N_22582,N_22484,N_22195);
nand U22583 (N_22583,N_22463,N_22248);
xnor U22584 (N_22584,N_22147,N_22121);
nor U22585 (N_22585,N_22023,N_22386);
nand U22586 (N_22586,N_22367,N_22284);
or U22587 (N_22587,N_22342,N_22326);
nor U22588 (N_22588,N_22024,N_22344);
xor U22589 (N_22589,N_22080,N_22234);
or U22590 (N_22590,N_22334,N_22268);
nand U22591 (N_22591,N_22449,N_22209);
xnor U22592 (N_22592,N_22377,N_22166);
nand U22593 (N_22593,N_22368,N_22264);
and U22594 (N_22594,N_22380,N_22432);
xor U22595 (N_22595,N_22152,N_22407);
nand U22596 (N_22596,N_22306,N_22331);
nand U22597 (N_22597,N_22142,N_22174);
nand U22598 (N_22598,N_22361,N_22193);
xor U22599 (N_22599,N_22187,N_22474);
or U22600 (N_22600,N_22175,N_22333);
and U22601 (N_22601,N_22348,N_22355);
nor U22602 (N_22602,N_22387,N_22143);
nand U22603 (N_22603,N_22186,N_22280);
nand U22604 (N_22604,N_22461,N_22154);
xor U22605 (N_22605,N_22254,N_22253);
nand U22606 (N_22606,N_22374,N_22434);
nor U22607 (N_22607,N_22499,N_22351);
and U22608 (N_22608,N_22138,N_22114);
nand U22609 (N_22609,N_22283,N_22435);
and U22610 (N_22610,N_22392,N_22113);
nor U22611 (N_22611,N_22315,N_22412);
xnor U22612 (N_22612,N_22335,N_22038);
and U22613 (N_22613,N_22170,N_22140);
nor U22614 (N_22614,N_22350,N_22153);
nand U22615 (N_22615,N_22115,N_22420);
xnor U22616 (N_22616,N_22073,N_22013);
xnor U22617 (N_22617,N_22464,N_22104);
nand U22618 (N_22618,N_22490,N_22440);
nand U22619 (N_22619,N_22031,N_22275);
and U22620 (N_22620,N_22019,N_22472);
or U22621 (N_22621,N_22010,N_22459);
nand U22622 (N_22622,N_22289,N_22062);
and U22623 (N_22623,N_22035,N_22443);
or U22624 (N_22624,N_22441,N_22406);
nand U22625 (N_22625,N_22421,N_22455);
nor U22626 (N_22626,N_22044,N_22452);
nand U22627 (N_22627,N_22448,N_22477);
xnor U22628 (N_22628,N_22475,N_22027);
and U22629 (N_22629,N_22242,N_22307);
nand U22630 (N_22630,N_22257,N_22224);
and U22631 (N_22631,N_22091,N_22395);
and U22632 (N_22632,N_22148,N_22426);
xnor U22633 (N_22633,N_22485,N_22365);
nor U22634 (N_22634,N_22372,N_22312);
nand U22635 (N_22635,N_22467,N_22243);
or U22636 (N_22636,N_22043,N_22081);
and U22637 (N_22637,N_22155,N_22245);
nor U22638 (N_22638,N_22469,N_22095);
or U22639 (N_22639,N_22087,N_22305);
nor U22640 (N_22640,N_22252,N_22423);
nor U22641 (N_22641,N_22028,N_22422);
or U22642 (N_22642,N_22045,N_22444);
or U22643 (N_22643,N_22325,N_22277);
or U22644 (N_22644,N_22319,N_22036);
xor U22645 (N_22645,N_22236,N_22226);
nor U22646 (N_22646,N_22338,N_22302);
nor U22647 (N_22647,N_22131,N_22139);
nand U22648 (N_22648,N_22456,N_22404);
and U22649 (N_22649,N_22323,N_22112);
nand U22650 (N_22650,N_22006,N_22182);
or U22651 (N_22651,N_22130,N_22072);
or U22652 (N_22652,N_22288,N_22416);
xor U22653 (N_22653,N_22433,N_22190);
nor U22654 (N_22654,N_22232,N_22488);
nand U22655 (N_22655,N_22332,N_22055);
and U22656 (N_22656,N_22238,N_22408);
nor U22657 (N_22657,N_22007,N_22336);
xor U22658 (N_22658,N_22161,N_22047);
nor U22659 (N_22659,N_22057,N_22447);
xor U22660 (N_22660,N_22272,N_22296);
nor U22661 (N_22661,N_22299,N_22103);
nand U22662 (N_22662,N_22458,N_22442);
and U22663 (N_22663,N_22039,N_22227);
and U22664 (N_22664,N_22199,N_22071);
or U22665 (N_22665,N_22179,N_22076);
nor U22666 (N_22666,N_22181,N_22221);
or U22667 (N_22667,N_22137,N_22362);
nand U22668 (N_22668,N_22203,N_22340);
nand U22669 (N_22669,N_22352,N_22157);
nand U22670 (N_22670,N_22046,N_22228);
and U22671 (N_22671,N_22177,N_22313);
nor U22672 (N_22672,N_22322,N_22309);
nand U22673 (N_22673,N_22462,N_22069);
or U22674 (N_22674,N_22223,N_22294);
xnor U22675 (N_22675,N_22375,N_22293);
and U22676 (N_22676,N_22070,N_22437);
or U22677 (N_22677,N_22320,N_22172);
xnor U22678 (N_22678,N_22052,N_22399);
xnor U22679 (N_22679,N_22267,N_22176);
nand U22680 (N_22680,N_22359,N_22120);
nand U22681 (N_22681,N_22300,N_22054);
and U22682 (N_22682,N_22324,N_22118);
nor U22683 (N_22683,N_22110,N_22491);
and U22684 (N_22684,N_22454,N_22287);
xnor U22685 (N_22685,N_22249,N_22191);
xnor U22686 (N_22686,N_22197,N_22439);
nor U22687 (N_22687,N_22327,N_22171);
nor U22688 (N_22688,N_22446,N_22345);
xnor U22689 (N_22689,N_22487,N_22417);
and U22690 (N_22690,N_22014,N_22000);
xor U22691 (N_22691,N_22303,N_22132);
nor U22692 (N_22692,N_22108,N_22145);
nand U22693 (N_22693,N_22419,N_22089);
or U22694 (N_22694,N_22258,N_22219);
and U22695 (N_22695,N_22003,N_22212);
xnor U22696 (N_22696,N_22384,N_22304);
or U22697 (N_22697,N_22184,N_22111);
or U22698 (N_22698,N_22301,N_22124);
or U22699 (N_22699,N_22263,N_22083);
xnor U22700 (N_22700,N_22205,N_22216);
and U22701 (N_22701,N_22401,N_22378);
and U22702 (N_22702,N_22376,N_22274);
nor U22703 (N_22703,N_22358,N_22058);
nor U22704 (N_22704,N_22298,N_22168);
and U22705 (N_22705,N_22388,N_22090);
and U22706 (N_22706,N_22489,N_22200);
and U22707 (N_22707,N_22032,N_22151);
and U22708 (N_22708,N_22281,N_22479);
and U22709 (N_22709,N_22188,N_22468);
xor U22710 (N_22710,N_22189,N_22068);
and U22711 (N_22711,N_22402,N_22494);
xor U22712 (N_22712,N_22400,N_22318);
nor U22713 (N_22713,N_22276,N_22405);
or U22714 (N_22714,N_22369,N_22160);
nand U22715 (N_22715,N_22430,N_22011);
nand U22716 (N_22716,N_22262,N_22339);
nand U22717 (N_22717,N_22493,N_22034);
and U22718 (N_22718,N_22360,N_22343);
or U22719 (N_22719,N_22290,N_22230);
or U22720 (N_22720,N_22133,N_22092);
nand U22721 (N_22721,N_22366,N_22295);
and U22722 (N_22722,N_22214,N_22016);
xor U22723 (N_22723,N_22244,N_22192);
nor U22724 (N_22724,N_22397,N_22101);
or U22725 (N_22725,N_22018,N_22163);
and U22726 (N_22726,N_22173,N_22486);
nor U22727 (N_22727,N_22425,N_22218);
and U22728 (N_22728,N_22246,N_22079);
or U22729 (N_22729,N_22093,N_22077);
and U22730 (N_22730,N_22002,N_22321);
xnor U22731 (N_22731,N_22371,N_22471);
nand U22732 (N_22732,N_22025,N_22217);
nor U22733 (N_22733,N_22379,N_22037);
xnor U22734 (N_22734,N_22498,N_22162);
nand U22735 (N_22735,N_22109,N_22451);
nor U22736 (N_22736,N_22106,N_22201);
and U22737 (N_22737,N_22385,N_22389);
and U22738 (N_22738,N_22051,N_22383);
xnor U22739 (N_22739,N_22269,N_22278);
or U22740 (N_22740,N_22005,N_22211);
xor U22741 (N_22741,N_22241,N_22123);
and U22742 (N_22742,N_22482,N_22398);
xnor U22743 (N_22743,N_22279,N_22282);
xor U22744 (N_22744,N_22017,N_22346);
and U22745 (N_22745,N_22256,N_22001);
xor U22746 (N_22746,N_22164,N_22457);
nand U22747 (N_22747,N_22409,N_22061);
nor U22748 (N_22748,N_22410,N_22094);
or U22749 (N_22749,N_22273,N_22247);
nand U22750 (N_22750,N_22030,N_22439);
and U22751 (N_22751,N_22000,N_22403);
nand U22752 (N_22752,N_22088,N_22438);
and U22753 (N_22753,N_22229,N_22134);
nor U22754 (N_22754,N_22039,N_22437);
and U22755 (N_22755,N_22090,N_22394);
xnor U22756 (N_22756,N_22201,N_22152);
nor U22757 (N_22757,N_22000,N_22497);
and U22758 (N_22758,N_22347,N_22110);
nor U22759 (N_22759,N_22347,N_22451);
nor U22760 (N_22760,N_22460,N_22114);
or U22761 (N_22761,N_22204,N_22006);
or U22762 (N_22762,N_22006,N_22209);
nand U22763 (N_22763,N_22492,N_22176);
or U22764 (N_22764,N_22419,N_22204);
nand U22765 (N_22765,N_22084,N_22286);
or U22766 (N_22766,N_22126,N_22210);
nor U22767 (N_22767,N_22183,N_22029);
xor U22768 (N_22768,N_22062,N_22158);
xnor U22769 (N_22769,N_22290,N_22393);
xnor U22770 (N_22770,N_22358,N_22265);
nand U22771 (N_22771,N_22465,N_22095);
nand U22772 (N_22772,N_22277,N_22452);
nand U22773 (N_22773,N_22481,N_22417);
or U22774 (N_22774,N_22428,N_22459);
nand U22775 (N_22775,N_22368,N_22366);
or U22776 (N_22776,N_22376,N_22125);
or U22777 (N_22777,N_22134,N_22022);
xor U22778 (N_22778,N_22028,N_22215);
nand U22779 (N_22779,N_22428,N_22226);
nor U22780 (N_22780,N_22429,N_22363);
or U22781 (N_22781,N_22273,N_22459);
or U22782 (N_22782,N_22066,N_22496);
and U22783 (N_22783,N_22156,N_22275);
nand U22784 (N_22784,N_22090,N_22044);
and U22785 (N_22785,N_22453,N_22421);
and U22786 (N_22786,N_22216,N_22184);
nor U22787 (N_22787,N_22185,N_22414);
nand U22788 (N_22788,N_22355,N_22255);
nor U22789 (N_22789,N_22298,N_22085);
nor U22790 (N_22790,N_22026,N_22250);
nor U22791 (N_22791,N_22388,N_22239);
nor U22792 (N_22792,N_22215,N_22121);
xor U22793 (N_22793,N_22220,N_22419);
nor U22794 (N_22794,N_22135,N_22280);
xor U22795 (N_22795,N_22431,N_22397);
xor U22796 (N_22796,N_22296,N_22165);
nand U22797 (N_22797,N_22416,N_22044);
nand U22798 (N_22798,N_22482,N_22337);
xnor U22799 (N_22799,N_22446,N_22013);
nand U22800 (N_22800,N_22302,N_22347);
and U22801 (N_22801,N_22322,N_22301);
xor U22802 (N_22802,N_22199,N_22472);
xor U22803 (N_22803,N_22270,N_22206);
or U22804 (N_22804,N_22375,N_22328);
nor U22805 (N_22805,N_22250,N_22321);
nor U22806 (N_22806,N_22359,N_22205);
nor U22807 (N_22807,N_22125,N_22036);
and U22808 (N_22808,N_22017,N_22149);
or U22809 (N_22809,N_22252,N_22167);
or U22810 (N_22810,N_22441,N_22064);
and U22811 (N_22811,N_22068,N_22082);
or U22812 (N_22812,N_22116,N_22395);
xor U22813 (N_22813,N_22243,N_22050);
xnor U22814 (N_22814,N_22231,N_22198);
xor U22815 (N_22815,N_22049,N_22296);
xor U22816 (N_22816,N_22021,N_22300);
and U22817 (N_22817,N_22198,N_22491);
or U22818 (N_22818,N_22002,N_22433);
xor U22819 (N_22819,N_22209,N_22186);
xor U22820 (N_22820,N_22492,N_22172);
or U22821 (N_22821,N_22445,N_22167);
xor U22822 (N_22822,N_22084,N_22274);
nor U22823 (N_22823,N_22467,N_22305);
and U22824 (N_22824,N_22383,N_22057);
nand U22825 (N_22825,N_22372,N_22499);
or U22826 (N_22826,N_22067,N_22091);
or U22827 (N_22827,N_22408,N_22036);
nand U22828 (N_22828,N_22419,N_22277);
or U22829 (N_22829,N_22233,N_22461);
and U22830 (N_22830,N_22340,N_22040);
and U22831 (N_22831,N_22143,N_22054);
nor U22832 (N_22832,N_22280,N_22252);
or U22833 (N_22833,N_22066,N_22215);
and U22834 (N_22834,N_22456,N_22449);
or U22835 (N_22835,N_22322,N_22085);
xnor U22836 (N_22836,N_22373,N_22272);
or U22837 (N_22837,N_22154,N_22243);
and U22838 (N_22838,N_22124,N_22390);
xnor U22839 (N_22839,N_22494,N_22217);
or U22840 (N_22840,N_22065,N_22470);
and U22841 (N_22841,N_22139,N_22196);
nor U22842 (N_22842,N_22325,N_22258);
nor U22843 (N_22843,N_22090,N_22103);
or U22844 (N_22844,N_22213,N_22445);
and U22845 (N_22845,N_22137,N_22363);
nor U22846 (N_22846,N_22248,N_22417);
or U22847 (N_22847,N_22418,N_22034);
nor U22848 (N_22848,N_22265,N_22016);
or U22849 (N_22849,N_22472,N_22028);
xnor U22850 (N_22850,N_22169,N_22153);
or U22851 (N_22851,N_22232,N_22043);
xor U22852 (N_22852,N_22103,N_22316);
nor U22853 (N_22853,N_22271,N_22004);
nand U22854 (N_22854,N_22357,N_22368);
and U22855 (N_22855,N_22436,N_22279);
nand U22856 (N_22856,N_22157,N_22109);
and U22857 (N_22857,N_22190,N_22116);
and U22858 (N_22858,N_22078,N_22352);
or U22859 (N_22859,N_22259,N_22453);
nand U22860 (N_22860,N_22420,N_22397);
and U22861 (N_22861,N_22333,N_22248);
nand U22862 (N_22862,N_22364,N_22206);
and U22863 (N_22863,N_22097,N_22015);
and U22864 (N_22864,N_22474,N_22326);
xor U22865 (N_22865,N_22496,N_22304);
nor U22866 (N_22866,N_22107,N_22236);
and U22867 (N_22867,N_22145,N_22387);
xor U22868 (N_22868,N_22141,N_22472);
or U22869 (N_22869,N_22256,N_22092);
nor U22870 (N_22870,N_22395,N_22261);
and U22871 (N_22871,N_22384,N_22281);
or U22872 (N_22872,N_22468,N_22373);
nor U22873 (N_22873,N_22411,N_22007);
nor U22874 (N_22874,N_22019,N_22351);
nand U22875 (N_22875,N_22030,N_22492);
or U22876 (N_22876,N_22268,N_22031);
and U22877 (N_22877,N_22392,N_22344);
nand U22878 (N_22878,N_22219,N_22429);
nor U22879 (N_22879,N_22321,N_22373);
and U22880 (N_22880,N_22160,N_22447);
xor U22881 (N_22881,N_22189,N_22207);
and U22882 (N_22882,N_22351,N_22099);
and U22883 (N_22883,N_22033,N_22120);
xnor U22884 (N_22884,N_22225,N_22069);
nor U22885 (N_22885,N_22175,N_22015);
xor U22886 (N_22886,N_22315,N_22337);
xor U22887 (N_22887,N_22033,N_22091);
nor U22888 (N_22888,N_22466,N_22369);
and U22889 (N_22889,N_22328,N_22110);
or U22890 (N_22890,N_22121,N_22176);
xnor U22891 (N_22891,N_22108,N_22363);
and U22892 (N_22892,N_22424,N_22158);
and U22893 (N_22893,N_22201,N_22354);
nor U22894 (N_22894,N_22137,N_22123);
xor U22895 (N_22895,N_22092,N_22114);
nor U22896 (N_22896,N_22206,N_22015);
nand U22897 (N_22897,N_22491,N_22220);
nand U22898 (N_22898,N_22309,N_22397);
or U22899 (N_22899,N_22112,N_22119);
xor U22900 (N_22900,N_22049,N_22109);
or U22901 (N_22901,N_22132,N_22187);
and U22902 (N_22902,N_22300,N_22362);
and U22903 (N_22903,N_22180,N_22020);
nor U22904 (N_22904,N_22187,N_22096);
and U22905 (N_22905,N_22130,N_22451);
xor U22906 (N_22906,N_22191,N_22131);
or U22907 (N_22907,N_22074,N_22498);
or U22908 (N_22908,N_22246,N_22204);
nand U22909 (N_22909,N_22061,N_22135);
or U22910 (N_22910,N_22350,N_22414);
xor U22911 (N_22911,N_22064,N_22412);
nand U22912 (N_22912,N_22226,N_22487);
or U22913 (N_22913,N_22127,N_22368);
or U22914 (N_22914,N_22337,N_22049);
xor U22915 (N_22915,N_22388,N_22029);
or U22916 (N_22916,N_22411,N_22208);
and U22917 (N_22917,N_22152,N_22031);
and U22918 (N_22918,N_22256,N_22011);
and U22919 (N_22919,N_22011,N_22253);
and U22920 (N_22920,N_22232,N_22076);
nand U22921 (N_22921,N_22108,N_22027);
xor U22922 (N_22922,N_22338,N_22255);
xor U22923 (N_22923,N_22298,N_22090);
nand U22924 (N_22924,N_22200,N_22047);
nand U22925 (N_22925,N_22377,N_22455);
nor U22926 (N_22926,N_22314,N_22369);
nor U22927 (N_22927,N_22108,N_22349);
nand U22928 (N_22928,N_22149,N_22081);
or U22929 (N_22929,N_22013,N_22118);
xnor U22930 (N_22930,N_22369,N_22230);
xor U22931 (N_22931,N_22463,N_22130);
nor U22932 (N_22932,N_22210,N_22159);
or U22933 (N_22933,N_22106,N_22333);
nor U22934 (N_22934,N_22423,N_22221);
xnor U22935 (N_22935,N_22089,N_22370);
nand U22936 (N_22936,N_22474,N_22050);
and U22937 (N_22937,N_22279,N_22216);
or U22938 (N_22938,N_22385,N_22338);
xnor U22939 (N_22939,N_22468,N_22222);
nand U22940 (N_22940,N_22253,N_22027);
nand U22941 (N_22941,N_22398,N_22455);
nand U22942 (N_22942,N_22400,N_22070);
or U22943 (N_22943,N_22444,N_22038);
and U22944 (N_22944,N_22110,N_22162);
and U22945 (N_22945,N_22370,N_22479);
nand U22946 (N_22946,N_22309,N_22142);
nor U22947 (N_22947,N_22025,N_22365);
or U22948 (N_22948,N_22153,N_22320);
nand U22949 (N_22949,N_22128,N_22261);
nand U22950 (N_22950,N_22368,N_22090);
nor U22951 (N_22951,N_22190,N_22128);
nor U22952 (N_22952,N_22279,N_22074);
or U22953 (N_22953,N_22133,N_22060);
and U22954 (N_22954,N_22223,N_22277);
xnor U22955 (N_22955,N_22345,N_22142);
and U22956 (N_22956,N_22085,N_22024);
or U22957 (N_22957,N_22006,N_22300);
and U22958 (N_22958,N_22133,N_22285);
nand U22959 (N_22959,N_22094,N_22164);
nand U22960 (N_22960,N_22355,N_22120);
nand U22961 (N_22961,N_22068,N_22130);
and U22962 (N_22962,N_22000,N_22009);
and U22963 (N_22963,N_22477,N_22238);
nand U22964 (N_22964,N_22345,N_22430);
or U22965 (N_22965,N_22460,N_22088);
and U22966 (N_22966,N_22112,N_22236);
or U22967 (N_22967,N_22433,N_22135);
nor U22968 (N_22968,N_22275,N_22048);
and U22969 (N_22969,N_22285,N_22316);
or U22970 (N_22970,N_22164,N_22261);
nor U22971 (N_22971,N_22275,N_22089);
nand U22972 (N_22972,N_22097,N_22276);
and U22973 (N_22973,N_22449,N_22229);
and U22974 (N_22974,N_22076,N_22339);
nand U22975 (N_22975,N_22324,N_22276);
nand U22976 (N_22976,N_22143,N_22135);
xnor U22977 (N_22977,N_22051,N_22067);
nor U22978 (N_22978,N_22370,N_22406);
nand U22979 (N_22979,N_22306,N_22239);
and U22980 (N_22980,N_22119,N_22055);
xnor U22981 (N_22981,N_22147,N_22206);
and U22982 (N_22982,N_22249,N_22035);
xor U22983 (N_22983,N_22234,N_22415);
or U22984 (N_22984,N_22462,N_22206);
or U22985 (N_22985,N_22098,N_22486);
nand U22986 (N_22986,N_22127,N_22018);
nand U22987 (N_22987,N_22459,N_22097);
nand U22988 (N_22988,N_22116,N_22358);
nand U22989 (N_22989,N_22496,N_22489);
or U22990 (N_22990,N_22262,N_22216);
xnor U22991 (N_22991,N_22053,N_22007);
nand U22992 (N_22992,N_22007,N_22175);
and U22993 (N_22993,N_22142,N_22324);
and U22994 (N_22994,N_22061,N_22164);
and U22995 (N_22995,N_22397,N_22035);
nor U22996 (N_22996,N_22315,N_22217);
nor U22997 (N_22997,N_22349,N_22354);
nand U22998 (N_22998,N_22424,N_22242);
nor U22999 (N_22999,N_22490,N_22413);
or U23000 (N_23000,N_22886,N_22949);
nand U23001 (N_23001,N_22858,N_22507);
nand U23002 (N_23002,N_22546,N_22624);
and U23003 (N_23003,N_22954,N_22899);
and U23004 (N_23004,N_22629,N_22598);
xor U23005 (N_23005,N_22861,N_22508);
or U23006 (N_23006,N_22797,N_22838);
or U23007 (N_23007,N_22513,N_22511);
and U23008 (N_23008,N_22958,N_22935);
nand U23009 (N_23009,N_22557,N_22763);
nor U23010 (N_23010,N_22810,N_22556);
nor U23011 (N_23011,N_22924,N_22616);
xnor U23012 (N_23012,N_22590,N_22667);
xnor U23013 (N_23013,N_22552,N_22715);
nor U23014 (N_23014,N_22887,N_22894);
and U23015 (N_23015,N_22669,N_22560);
or U23016 (N_23016,N_22712,N_22683);
and U23017 (N_23017,N_22702,N_22581);
nand U23018 (N_23018,N_22966,N_22561);
nor U23019 (N_23019,N_22722,N_22842);
xnor U23020 (N_23020,N_22915,N_22802);
nor U23021 (N_23021,N_22892,N_22536);
nand U23022 (N_23022,N_22694,N_22990);
and U23023 (N_23023,N_22964,N_22878);
nor U23024 (N_23024,N_22545,N_22597);
and U23025 (N_23025,N_22647,N_22870);
and U23026 (N_23026,N_22944,N_22791);
and U23027 (N_23027,N_22516,N_22961);
xnor U23028 (N_23028,N_22829,N_22816);
nand U23029 (N_23029,N_22679,N_22739);
xnor U23030 (N_23030,N_22857,N_22535);
and U23031 (N_23031,N_22913,N_22898);
nor U23032 (N_23032,N_22927,N_22877);
and U23033 (N_23033,N_22879,N_22550);
or U23034 (N_23034,N_22754,N_22606);
and U23035 (N_23035,N_22941,N_22919);
xnor U23036 (N_23036,N_22868,N_22986);
or U23037 (N_23037,N_22741,N_22809);
nand U23038 (N_23038,N_22817,N_22759);
nor U23039 (N_23039,N_22777,N_22768);
and U23040 (N_23040,N_22957,N_22732);
nand U23041 (N_23041,N_22785,N_22834);
and U23042 (N_23042,N_22852,N_22855);
or U23043 (N_23043,N_22635,N_22648);
nand U23044 (N_23044,N_22562,N_22605);
xor U23045 (N_23045,N_22970,N_22976);
nand U23046 (N_23046,N_22888,N_22673);
nor U23047 (N_23047,N_22575,N_22713);
nand U23048 (N_23048,N_22529,N_22850);
and U23049 (N_23049,N_22674,N_22916);
nand U23050 (N_23050,N_22541,N_22952);
or U23051 (N_23051,N_22528,N_22599);
or U23052 (N_23052,N_22746,N_22974);
xnor U23053 (N_23053,N_22853,N_22818);
xor U23054 (N_23054,N_22982,N_22634);
nand U23055 (N_23055,N_22671,N_22984);
nand U23056 (N_23056,N_22865,N_22538);
nand U23057 (N_23057,N_22824,N_22663);
nand U23058 (N_23058,N_22717,N_22757);
nand U23059 (N_23059,N_22764,N_22665);
nor U23060 (N_23060,N_22609,N_22973);
or U23061 (N_23061,N_22839,N_22940);
nand U23062 (N_23062,N_22503,N_22678);
nor U23063 (N_23063,N_22658,N_22577);
or U23064 (N_23064,N_22636,N_22504);
or U23065 (N_23065,N_22705,N_22758);
nand U23066 (N_23066,N_22896,N_22825);
nand U23067 (N_23067,N_22854,N_22977);
xor U23068 (N_23068,N_22847,N_22744);
or U23069 (N_23069,N_22554,N_22718);
nand U23070 (N_23070,N_22716,N_22583);
and U23071 (N_23071,N_22874,N_22639);
or U23072 (N_23072,N_22745,N_22889);
xor U23073 (N_23073,N_22905,N_22698);
xnor U23074 (N_23074,N_22843,N_22523);
nor U23075 (N_23075,N_22837,N_22537);
nor U23076 (N_23076,N_22936,N_22773);
nand U23077 (N_23077,N_22823,N_22519);
or U23078 (N_23078,N_22790,N_22965);
and U23079 (N_23079,N_22567,N_22531);
and U23080 (N_23080,N_22867,N_22738);
xor U23081 (N_23081,N_22814,N_22807);
xor U23082 (N_23082,N_22607,N_22524);
xnor U23083 (N_23083,N_22788,N_22871);
nor U23084 (N_23084,N_22506,N_22626);
or U23085 (N_23085,N_22939,N_22926);
or U23086 (N_23086,N_22580,N_22640);
nor U23087 (N_23087,N_22544,N_22950);
nand U23088 (N_23088,N_22897,N_22903);
xor U23089 (N_23089,N_22666,N_22633);
and U23090 (N_23090,N_22846,N_22645);
nand U23091 (N_23091,N_22863,N_22512);
and U23092 (N_23092,N_22796,N_22589);
or U23093 (N_23093,N_22830,N_22841);
nor U23094 (N_23094,N_22762,N_22547);
and U23095 (N_23095,N_22951,N_22564);
and U23096 (N_23096,N_22617,N_22572);
nor U23097 (N_23097,N_22960,N_22831);
nor U23098 (N_23098,N_22812,N_22735);
and U23099 (N_23099,N_22991,N_22859);
xor U23100 (N_23100,N_22743,N_22568);
xnor U23101 (N_23101,N_22882,N_22637);
or U23102 (N_23102,N_22734,N_22925);
xor U23103 (N_23103,N_22780,N_22769);
nand U23104 (N_23104,N_22928,N_22776);
nor U23105 (N_23105,N_22680,N_22723);
xnor U23106 (N_23106,N_22891,N_22684);
nand U23107 (N_23107,N_22736,N_22917);
nand U23108 (N_23108,N_22630,N_22670);
or U23109 (N_23109,N_22800,N_22584);
xnor U23110 (N_23110,N_22849,N_22500);
xnor U23111 (N_23111,N_22947,N_22709);
nor U23112 (N_23112,N_22992,N_22693);
and U23113 (N_23113,N_22932,N_22860);
or U23114 (N_23114,N_22752,N_22921);
or U23115 (N_23115,N_22959,N_22573);
or U23116 (N_23116,N_22594,N_22934);
nand U23117 (N_23117,N_22920,N_22748);
xor U23118 (N_23118,N_22851,N_22972);
or U23119 (N_23119,N_22969,N_22714);
and U23120 (N_23120,N_22908,N_22621);
nor U23121 (N_23121,N_22760,N_22782);
or U23122 (N_23122,N_22672,N_22601);
or U23123 (N_23123,N_22771,N_22893);
xnor U23124 (N_23124,N_22586,N_22938);
or U23125 (N_23125,N_22755,N_22795);
nor U23126 (N_23126,N_22505,N_22644);
xnor U23127 (N_23127,N_22625,N_22578);
or U23128 (N_23128,N_22930,N_22798);
nand U23129 (N_23129,N_22815,N_22955);
and U23130 (N_23130,N_22750,N_22675);
xor U23131 (N_23131,N_22772,N_22585);
nor U23132 (N_23132,N_22997,N_22983);
and U23133 (N_23133,N_22996,N_22661);
nor U23134 (N_23134,N_22727,N_22613);
nor U23135 (N_23135,N_22682,N_22933);
nand U23136 (N_23136,N_22646,N_22792);
nand U23137 (N_23137,N_22539,N_22828);
nand U23138 (N_23138,N_22628,N_22726);
and U23139 (N_23139,N_22518,N_22642);
or U23140 (N_23140,N_22612,N_22706);
and U23141 (N_23141,N_22962,N_22604);
nand U23142 (N_23142,N_22655,N_22710);
xor U23143 (N_23143,N_22533,N_22866);
or U23144 (N_23144,N_22803,N_22724);
and U23145 (N_23145,N_22627,N_22520);
or U23146 (N_23146,N_22840,N_22565);
and U23147 (N_23147,N_22942,N_22728);
nand U23148 (N_23148,N_22632,N_22844);
nor U23149 (N_23149,N_22593,N_22526);
nand U23150 (N_23150,N_22603,N_22509);
nor U23151 (N_23151,N_22775,N_22967);
and U23152 (N_23152,N_22731,N_22631);
or U23153 (N_23153,N_22953,N_22689);
nand U23154 (N_23154,N_22579,N_22956);
xor U23155 (N_23155,N_22912,N_22923);
and U23156 (N_23156,N_22532,N_22806);
or U23157 (N_23157,N_22574,N_22668);
xor U23158 (N_23158,N_22995,N_22551);
nand U23159 (N_23159,N_22740,N_22558);
or U23160 (N_23160,N_22622,N_22793);
nand U23161 (N_23161,N_22600,N_22826);
and U23162 (N_23162,N_22765,N_22988);
nor U23163 (N_23163,N_22766,N_22761);
and U23164 (N_23164,N_22774,N_22697);
nor U23165 (N_23165,N_22542,N_22742);
nor U23166 (N_23166,N_22566,N_22804);
or U23167 (N_23167,N_22695,N_22999);
or U23168 (N_23168,N_22729,N_22522);
nor U23169 (N_23169,N_22638,N_22548);
or U23170 (N_23170,N_22571,N_22690);
or U23171 (N_23171,N_22657,N_22989);
and U23172 (N_23172,N_22770,N_22827);
and U23173 (N_23173,N_22981,N_22994);
and U23174 (N_23174,N_22813,N_22980);
nand U23175 (N_23175,N_22836,N_22608);
nor U23176 (N_23176,N_22582,N_22975);
or U23177 (N_23177,N_22602,N_22685);
and U23178 (N_23178,N_22811,N_22654);
or U23179 (N_23179,N_22681,N_22971);
nand U23180 (N_23180,N_22721,N_22929);
or U23181 (N_23181,N_22786,N_22649);
or U23182 (N_23182,N_22730,N_22998);
and U23183 (N_23183,N_22659,N_22563);
and U23184 (N_23184,N_22595,N_22869);
and U23185 (N_23185,N_22623,N_22819);
nand U23186 (N_23186,N_22676,N_22821);
and U23187 (N_23187,N_22502,N_22704);
xnor U23188 (N_23188,N_22787,N_22707);
xnor U23189 (N_23189,N_22615,N_22906);
or U23190 (N_23190,N_22688,N_22720);
nand U23191 (N_23191,N_22711,N_22549);
nand U23192 (N_23192,N_22737,N_22588);
and U23193 (N_23193,N_22660,N_22687);
xor U23194 (N_23194,N_22948,N_22559);
and U23195 (N_23195,N_22651,N_22914);
nor U23196 (N_23196,N_22778,N_22864);
and U23197 (N_23197,N_22979,N_22845);
or U23198 (N_23198,N_22569,N_22833);
or U23199 (N_23199,N_22614,N_22880);
xnor U23200 (N_23200,N_22692,N_22756);
nor U23201 (N_23201,N_22643,N_22805);
nor U23202 (N_23202,N_22515,N_22993);
xor U23203 (N_23203,N_22719,N_22872);
xor U23204 (N_23204,N_22619,N_22873);
and U23205 (N_23205,N_22696,N_22904);
and U23206 (N_23206,N_22677,N_22596);
nand U23207 (N_23207,N_22911,N_22856);
or U23208 (N_23208,N_22592,N_22701);
and U23209 (N_23209,N_22781,N_22664);
nand U23210 (N_23210,N_22789,N_22540);
nor U23211 (N_23211,N_22517,N_22591);
xnor U23212 (N_23212,N_22653,N_22820);
or U23213 (N_23213,N_22945,N_22652);
and U23214 (N_23214,N_22747,N_22901);
nand U23215 (N_23215,N_22753,N_22987);
xnor U23216 (N_23216,N_22799,N_22832);
or U23217 (N_23217,N_22978,N_22862);
nor U23218 (N_23218,N_22922,N_22783);
and U23219 (N_23219,N_22848,N_22876);
and U23220 (N_23220,N_22553,N_22686);
and U23221 (N_23221,N_22570,N_22902);
xnor U23222 (N_23222,N_22725,N_22767);
xor U23223 (N_23223,N_22521,N_22703);
nand U23224 (N_23224,N_22885,N_22963);
and U23225 (N_23225,N_22907,N_22931);
nand U23226 (N_23226,N_22937,N_22527);
or U23227 (N_23227,N_22784,N_22910);
and U23228 (N_23228,N_22918,N_22801);
or U23229 (N_23229,N_22620,N_22749);
xnor U23230 (N_23230,N_22883,N_22691);
or U23231 (N_23231,N_22700,N_22530);
or U23232 (N_23232,N_22656,N_22881);
and U23233 (N_23233,N_22543,N_22699);
nor U23234 (N_23234,N_22618,N_22946);
and U23235 (N_23235,N_22835,N_22794);
xor U23236 (N_23236,N_22895,N_22968);
and U23237 (N_23237,N_22751,N_22890);
nor U23238 (N_23238,N_22525,N_22650);
nor U23239 (N_23239,N_22985,N_22779);
nor U23240 (N_23240,N_22501,N_22808);
nand U23241 (N_23241,N_22610,N_22534);
and U23242 (N_23242,N_22884,N_22641);
and U23243 (N_23243,N_22875,N_22708);
nor U23244 (N_23244,N_22909,N_22822);
and U23245 (N_23245,N_22555,N_22587);
xor U23246 (N_23246,N_22900,N_22662);
and U23247 (N_23247,N_22611,N_22733);
nand U23248 (N_23248,N_22576,N_22510);
nor U23249 (N_23249,N_22943,N_22514);
nand U23250 (N_23250,N_22901,N_22859);
xor U23251 (N_23251,N_22986,N_22783);
or U23252 (N_23252,N_22956,N_22752);
nor U23253 (N_23253,N_22606,N_22716);
or U23254 (N_23254,N_22880,N_22969);
nor U23255 (N_23255,N_22848,N_22758);
or U23256 (N_23256,N_22986,N_22899);
or U23257 (N_23257,N_22970,N_22614);
xnor U23258 (N_23258,N_22901,N_22742);
xor U23259 (N_23259,N_22738,N_22636);
and U23260 (N_23260,N_22756,N_22838);
nand U23261 (N_23261,N_22726,N_22673);
nand U23262 (N_23262,N_22939,N_22795);
xor U23263 (N_23263,N_22738,N_22832);
xor U23264 (N_23264,N_22914,N_22869);
and U23265 (N_23265,N_22636,N_22529);
nand U23266 (N_23266,N_22842,N_22847);
nand U23267 (N_23267,N_22874,N_22652);
and U23268 (N_23268,N_22756,N_22574);
or U23269 (N_23269,N_22856,N_22757);
or U23270 (N_23270,N_22661,N_22908);
xor U23271 (N_23271,N_22793,N_22688);
nor U23272 (N_23272,N_22593,N_22650);
and U23273 (N_23273,N_22968,N_22911);
xnor U23274 (N_23274,N_22535,N_22672);
or U23275 (N_23275,N_22893,N_22649);
xor U23276 (N_23276,N_22747,N_22956);
nand U23277 (N_23277,N_22761,N_22527);
and U23278 (N_23278,N_22656,N_22977);
nand U23279 (N_23279,N_22512,N_22810);
nand U23280 (N_23280,N_22598,N_22848);
and U23281 (N_23281,N_22535,N_22778);
xor U23282 (N_23282,N_22864,N_22577);
nand U23283 (N_23283,N_22877,N_22939);
and U23284 (N_23284,N_22795,N_22814);
or U23285 (N_23285,N_22933,N_22628);
nand U23286 (N_23286,N_22533,N_22892);
xnor U23287 (N_23287,N_22905,N_22739);
or U23288 (N_23288,N_22852,N_22869);
xor U23289 (N_23289,N_22810,N_22816);
or U23290 (N_23290,N_22853,N_22993);
nor U23291 (N_23291,N_22812,N_22894);
nor U23292 (N_23292,N_22556,N_22614);
nand U23293 (N_23293,N_22755,N_22598);
xor U23294 (N_23294,N_22950,N_22879);
xnor U23295 (N_23295,N_22617,N_22521);
or U23296 (N_23296,N_22766,N_22840);
or U23297 (N_23297,N_22995,N_22795);
and U23298 (N_23298,N_22613,N_22771);
nand U23299 (N_23299,N_22694,N_22599);
xor U23300 (N_23300,N_22715,N_22889);
nand U23301 (N_23301,N_22635,N_22586);
and U23302 (N_23302,N_22946,N_22763);
and U23303 (N_23303,N_22932,N_22833);
and U23304 (N_23304,N_22732,N_22889);
nand U23305 (N_23305,N_22852,N_22577);
xnor U23306 (N_23306,N_22555,N_22734);
or U23307 (N_23307,N_22902,N_22939);
or U23308 (N_23308,N_22923,N_22765);
or U23309 (N_23309,N_22800,N_22783);
or U23310 (N_23310,N_22500,N_22802);
xor U23311 (N_23311,N_22822,N_22830);
nor U23312 (N_23312,N_22588,N_22764);
nand U23313 (N_23313,N_22559,N_22711);
xnor U23314 (N_23314,N_22825,N_22519);
and U23315 (N_23315,N_22957,N_22777);
xnor U23316 (N_23316,N_22812,N_22989);
xor U23317 (N_23317,N_22727,N_22570);
or U23318 (N_23318,N_22766,N_22880);
xnor U23319 (N_23319,N_22682,N_22582);
nand U23320 (N_23320,N_22764,N_22614);
and U23321 (N_23321,N_22551,N_22945);
nand U23322 (N_23322,N_22570,N_22559);
and U23323 (N_23323,N_22773,N_22657);
or U23324 (N_23324,N_22941,N_22969);
nand U23325 (N_23325,N_22593,N_22569);
nor U23326 (N_23326,N_22868,N_22682);
nand U23327 (N_23327,N_22932,N_22592);
or U23328 (N_23328,N_22632,N_22896);
or U23329 (N_23329,N_22921,N_22555);
nand U23330 (N_23330,N_22972,N_22913);
or U23331 (N_23331,N_22629,N_22697);
or U23332 (N_23332,N_22653,N_22841);
nand U23333 (N_23333,N_22607,N_22549);
or U23334 (N_23334,N_22667,N_22542);
nor U23335 (N_23335,N_22868,N_22689);
or U23336 (N_23336,N_22564,N_22846);
xor U23337 (N_23337,N_22959,N_22514);
or U23338 (N_23338,N_22877,N_22745);
or U23339 (N_23339,N_22690,N_22867);
or U23340 (N_23340,N_22902,N_22630);
and U23341 (N_23341,N_22597,N_22737);
nor U23342 (N_23342,N_22814,N_22976);
xnor U23343 (N_23343,N_22942,N_22703);
nand U23344 (N_23344,N_22913,N_22878);
nand U23345 (N_23345,N_22706,N_22841);
xnor U23346 (N_23346,N_22809,N_22799);
nor U23347 (N_23347,N_22903,N_22917);
xnor U23348 (N_23348,N_22843,N_22528);
and U23349 (N_23349,N_22576,N_22650);
or U23350 (N_23350,N_22597,N_22618);
nor U23351 (N_23351,N_22638,N_22880);
or U23352 (N_23352,N_22891,N_22955);
xor U23353 (N_23353,N_22571,N_22848);
or U23354 (N_23354,N_22730,N_22825);
xor U23355 (N_23355,N_22930,N_22696);
xor U23356 (N_23356,N_22694,N_22535);
or U23357 (N_23357,N_22503,N_22962);
nor U23358 (N_23358,N_22902,N_22643);
nand U23359 (N_23359,N_22644,N_22775);
or U23360 (N_23360,N_22558,N_22576);
xor U23361 (N_23361,N_22863,N_22605);
nand U23362 (N_23362,N_22512,N_22708);
and U23363 (N_23363,N_22606,N_22640);
nor U23364 (N_23364,N_22889,N_22969);
or U23365 (N_23365,N_22863,N_22515);
nor U23366 (N_23366,N_22710,N_22521);
nor U23367 (N_23367,N_22916,N_22842);
nand U23368 (N_23368,N_22558,N_22662);
and U23369 (N_23369,N_22743,N_22536);
nand U23370 (N_23370,N_22521,N_22942);
nor U23371 (N_23371,N_22750,N_22850);
nor U23372 (N_23372,N_22600,N_22501);
or U23373 (N_23373,N_22694,N_22886);
or U23374 (N_23374,N_22853,N_22755);
nand U23375 (N_23375,N_22513,N_22606);
nor U23376 (N_23376,N_22542,N_22987);
and U23377 (N_23377,N_22504,N_22775);
nand U23378 (N_23378,N_22941,N_22713);
nand U23379 (N_23379,N_22806,N_22588);
or U23380 (N_23380,N_22646,N_22703);
or U23381 (N_23381,N_22529,N_22989);
nand U23382 (N_23382,N_22858,N_22998);
nand U23383 (N_23383,N_22946,N_22770);
nand U23384 (N_23384,N_22842,N_22779);
or U23385 (N_23385,N_22739,N_22762);
xnor U23386 (N_23386,N_22664,N_22636);
xnor U23387 (N_23387,N_22512,N_22632);
or U23388 (N_23388,N_22699,N_22565);
and U23389 (N_23389,N_22972,N_22523);
and U23390 (N_23390,N_22644,N_22649);
nand U23391 (N_23391,N_22973,N_22884);
nand U23392 (N_23392,N_22723,N_22625);
nor U23393 (N_23393,N_22618,N_22548);
and U23394 (N_23394,N_22775,N_22734);
nand U23395 (N_23395,N_22584,N_22658);
nand U23396 (N_23396,N_22517,N_22526);
nor U23397 (N_23397,N_22978,N_22747);
and U23398 (N_23398,N_22546,N_22951);
and U23399 (N_23399,N_22838,N_22517);
xnor U23400 (N_23400,N_22835,N_22786);
nand U23401 (N_23401,N_22526,N_22790);
nor U23402 (N_23402,N_22634,N_22523);
nor U23403 (N_23403,N_22836,N_22936);
and U23404 (N_23404,N_22743,N_22821);
nand U23405 (N_23405,N_22957,N_22545);
or U23406 (N_23406,N_22507,N_22969);
and U23407 (N_23407,N_22894,N_22822);
and U23408 (N_23408,N_22592,N_22778);
nand U23409 (N_23409,N_22816,N_22744);
nor U23410 (N_23410,N_22842,N_22561);
nor U23411 (N_23411,N_22612,N_22649);
nand U23412 (N_23412,N_22886,N_22875);
or U23413 (N_23413,N_22685,N_22847);
or U23414 (N_23414,N_22637,N_22853);
nor U23415 (N_23415,N_22831,N_22881);
and U23416 (N_23416,N_22879,N_22938);
and U23417 (N_23417,N_22814,N_22615);
xnor U23418 (N_23418,N_22829,N_22847);
and U23419 (N_23419,N_22729,N_22577);
or U23420 (N_23420,N_22555,N_22690);
and U23421 (N_23421,N_22978,N_22718);
and U23422 (N_23422,N_22705,N_22685);
nor U23423 (N_23423,N_22886,N_22904);
nand U23424 (N_23424,N_22549,N_22763);
xnor U23425 (N_23425,N_22855,N_22672);
or U23426 (N_23426,N_22700,N_22721);
or U23427 (N_23427,N_22712,N_22531);
nand U23428 (N_23428,N_22528,N_22892);
and U23429 (N_23429,N_22898,N_22835);
nor U23430 (N_23430,N_22705,N_22597);
and U23431 (N_23431,N_22731,N_22809);
and U23432 (N_23432,N_22938,N_22612);
or U23433 (N_23433,N_22991,N_22772);
or U23434 (N_23434,N_22995,N_22558);
xnor U23435 (N_23435,N_22785,N_22819);
xor U23436 (N_23436,N_22703,N_22611);
or U23437 (N_23437,N_22627,N_22712);
xor U23438 (N_23438,N_22730,N_22970);
nand U23439 (N_23439,N_22987,N_22609);
xnor U23440 (N_23440,N_22887,N_22518);
xnor U23441 (N_23441,N_22897,N_22514);
xor U23442 (N_23442,N_22798,N_22741);
nand U23443 (N_23443,N_22924,N_22512);
and U23444 (N_23444,N_22952,N_22880);
and U23445 (N_23445,N_22949,N_22506);
and U23446 (N_23446,N_22857,N_22628);
nor U23447 (N_23447,N_22752,N_22606);
and U23448 (N_23448,N_22738,N_22768);
xnor U23449 (N_23449,N_22735,N_22916);
or U23450 (N_23450,N_22524,N_22714);
nand U23451 (N_23451,N_22668,N_22866);
or U23452 (N_23452,N_22568,N_22946);
xor U23453 (N_23453,N_22633,N_22675);
xor U23454 (N_23454,N_22716,N_22997);
nor U23455 (N_23455,N_22516,N_22601);
xor U23456 (N_23456,N_22636,N_22717);
xnor U23457 (N_23457,N_22847,N_22667);
nor U23458 (N_23458,N_22983,N_22665);
nand U23459 (N_23459,N_22756,N_22622);
or U23460 (N_23460,N_22828,N_22731);
xor U23461 (N_23461,N_22820,N_22505);
nor U23462 (N_23462,N_22712,N_22976);
and U23463 (N_23463,N_22719,N_22603);
nor U23464 (N_23464,N_22919,N_22584);
nand U23465 (N_23465,N_22759,N_22652);
nor U23466 (N_23466,N_22505,N_22850);
nand U23467 (N_23467,N_22765,N_22504);
nand U23468 (N_23468,N_22896,N_22570);
or U23469 (N_23469,N_22709,N_22650);
or U23470 (N_23470,N_22505,N_22975);
and U23471 (N_23471,N_22672,N_22702);
nor U23472 (N_23472,N_22785,N_22590);
nand U23473 (N_23473,N_22581,N_22984);
xnor U23474 (N_23474,N_22834,N_22526);
and U23475 (N_23475,N_22916,N_22660);
or U23476 (N_23476,N_22623,N_22961);
nand U23477 (N_23477,N_22569,N_22609);
nand U23478 (N_23478,N_22983,N_22633);
and U23479 (N_23479,N_22692,N_22614);
xor U23480 (N_23480,N_22724,N_22940);
nor U23481 (N_23481,N_22636,N_22570);
or U23482 (N_23482,N_22690,N_22951);
xnor U23483 (N_23483,N_22538,N_22713);
or U23484 (N_23484,N_22592,N_22697);
xnor U23485 (N_23485,N_22622,N_22539);
nand U23486 (N_23486,N_22861,N_22968);
xnor U23487 (N_23487,N_22683,N_22729);
or U23488 (N_23488,N_22853,N_22884);
nand U23489 (N_23489,N_22875,N_22997);
nor U23490 (N_23490,N_22784,N_22740);
and U23491 (N_23491,N_22668,N_22893);
nand U23492 (N_23492,N_22627,N_22573);
nor U23493 (N_23493,N_22807,N_22872);
or U23494 (N_23494,N_22948,N_22968);
nand U23495 (N_23495,N_22985,N_22552);
nand U23496 (N_23496,N_22657,N_22973);
and U23497 (N_23497,N_22549,N_22856);
nand U23498 (N_23498,N_22922,N_22973);
nand U23499 (N_23499,N_22923,N_22638);
nand U23500 (N_23500,N_23092,N_23341);
nand U23501 (N_23501,N_23093,N_23120);
nor U23502 (N_23502,N_23305,N_23184);
xor U23503 (N_23503,N_23339,N_23363);
nand U23504 (N_23504,N_23169,N_23483);
nor U23505 (N_23505,N_23048,N_23259);
nor U23506 (N_23506,N_23155,N_23386);
or U23507 (N_23507,N_23116,N_23369);
and U23508 (N_23508,N_23438,N_23097);
nor U23509 (N_23509,N_23394,N_23233);
nor U23510 (N_23510,N_23274,N_23337);
nand U23511 (N_23511,N_23181,N_23350);
xor U23512 (N_23512,N_23353,N_23293);
xnor U23513 (N_23513,N_23243,N_23471);
or U23514 (N_23514,N_23435,N_23406);
and U23515 (N_23515,N_23290,N_23066);
or U23516 (N_23516,N_23164,N_23316);
and U23517 (N_23517,N_23407,N_23022);
or U23518 (N_23518,N_23037,N_23188);
nor U23519 (N_23519,N_23235,N_23421);
nor U23520 (N_23520,N_23220,N_23298);
nor U23521 (N_23521,N_23027,N_23346);
nor U23522 (N_23522,N_23050,N_23349);
nor U23523 (N_23523,N_23128,N_23067);
and U23524 (N_23524,N_23045,N_23225);
xnor U23525 (N_23525,N_23217,N_23267);
and U23526 (N_23526,N_23417,N_23391);
nor U23527 (N_23527,N_23256,N_23289);
xnor U23528 (N_23528,N_23481,N_23042);
nand U23529 (N_23529,N_23371,N_23152);
xnor U23530 (N_23530,N_23165,N_23306);
or U23531 (N_23531,N_23159,N_23204);
xnor U23532 (N_23532,N_23013,N_23123);
or U23533 (N_23533,N_23433,N_23260);
nor U23534 (N_23534,N_23294,N_23231);
nor U23535 (N_23535,N_23439,N_23213);
nand U23536 (N_23536,N_23318,N_23102);
xor U23537 (N_23537,N_23121,N_23109);
xnor U23538 (N_23538,N_23016,N_23166);
and U23539 (N_23539,N_23324,N_23460);
or U23540 (N_23540,N_23319,N_23499);
and U23541 (N_23541,N_23073,N_23367);
nand U23542 (N_23542,N_23436,N_23244);
nand U23543 (N_23543,N_23418,N_23282);
nand U23544 (N_23544,N_23283,N_23090);
nor U23545 (N_23545,N_23464,N_23182);
nand U23546 (N_23546,N_23124,N_23332);
nand U23547 (N_23547,N_23126,N_23461);
nand U23548 (N_23548,N_23312,N_23281);
xor U23549 (N_23549,N_23467,N_23342);
and U23550 (N_23550,N_23211,N_23393);
nand U23551 (N_23551,N_23226,N_23030);
nor U23552 (N_23552,N_23029,N_23251);
xor U23553 (N_23553,N_23390,N_23223);
nor U23554 (N_23554,N_23362,N_23154);
nand U23555 (N_23555,N_23198,N_23424);
or U23556 (N_23556,N_23262,N_23366);
xnor U23557 (N_23557,N_23161,N_23385);
nor U23558 (N_23558,N_23403,N_23422);
xnor U23559 (N_23559,N_23352,N_23458);
xnor U23560 (N_23560,N_23317,N_23043);
or U23561 (N_23561,N_23426,N_23295);
xor U23562 (N_23562,N_23086,N_23208);
and U23563 (N_23563,N_23047,N_23334);
xor U23564 (N_23564,N_23484,N_23054);
nor U23565 (N_23565,N_23005,N_23375);
or U23566 (N_23566,N_23399,N_23117);
xor U23567 (N_23567,N_23264,N_23404);
nand U23568 (N_23568,N_23162,N_23330);
or U23569 (N_23569,N_23216,N_23437);
nor U23570 (N_23570,N_23008,N_23268);
and U23571 (N_23571,N_23376,N_23398);
xnor U23572 (N_23572,N_23493,N_23201);
or U23573 (N_23573,N_23234,N_23325);
and U23574 (N_23574,N_23333,N_23221);
and U23575 (N_23575,N_23487,N_23019);
nand U23576 (N_23576,N_23345,N_23203);
nor U23577 (N_23577,N_23272,N_23122);
and U23578 (N_23578,N_23100,N_23062);
nand U23579 (N_23579,N_23405,N_23329);
or U23580 (N_23580,N_23380,N_23140);
or U23581 (N_23581,N_23442,N_23018);
nand U23582 (N_23582,N_23300,N_23015);
xor U23583 (N_23583,N_23359,N_23137);
xnor U23584 (N_23584,N_23205,N_23292);
nand U23585 (N_23585,N_23130,N_23070);
nand U23586 (N_23586,N_23082,N_23365);
or U23587 (N_23587,N_23006,N_23309);
nor U23588 (N_23588,N_23237,N_23409);
nor U23589 (N_23589,N_23149,N_23096);
nand U23590 (N_23590,N_23263,N_23046);
and U23591 (N_23591,N_23313,N_23476);
or U23592 (N_23592,N_23469,N_23069);
nand U23593 (N_23593,N_23322,N_23443);
nor U23594 (N_23594,N_23197,N_23423);
xor U23595 (N_23595,N_23445,N_23456);
and U23596 (N_23596,N_23170,N_23158);
and U23597 (N_23597,N_23032,N_23191);
nand U23598 (N_23598,N_23173,N_23147);
nand U23599 (N_23599,N_23248,N_23083);
nand U23600 (N_23600,N_23089,N_23194);
nand U23601 (N_23601,N_23389,N_23299);
xnor U23602 (N_23602,N_23372,N_23098);
nand U23603 (N_23603,N_23133,N_23064);
or U23604 (N_23604,N_23114,N_23450);
xor U23605 (N_23605,N_23434,N_23344);
nor U23606 (N_23606,N_23466,N_23210);
or U23607 (N_23607,N_23072,N_23373);
nand U23608 (N_23608,N_23358,N_23141);
or U23609 (N_23609,N_23270,N_23463);
xnor U23610 (N_23610,N_23459,N_23415);
xnor U23611 (N_23611,N_23266,N_23011);
and U23612 (N_23612,N_23224,N_23475);
xnor U23613 (N_23613,N_23303,N_23049);
or U23614 (N_23614,N_23279,N_23058);
xnor U23615 (N_23615,N_23364,N_23232);
nor U23616 (N_23616,N_23340,N_23452);
nand U23617 (N_23617,N_23347,N_23085);
or U23618 (N_23618,N_23026,N_23419);
or U23619 (N_23619,N_23125,N_23496);
nand U23620 (N_23620,N_23250,N_23039);
nor U23621 (N_23621,N_23257,N_23180);
nor U23622 (N_23622,N_23377,N_23106);
and U23623 (N_23623,N_23304,N_23271);
xnor U23624 (N_23624,N_23041,N_23408);
and U23625 (N_23625,N_23132,N_23025);
or U23626 (N_23626,N_23061,N_23453);
or U23627 (N_23627,N_23374,N_23455);
nand U23628 (N_23628,N_23253,N_23056);
nand U23629 (N_23629,N_23079,N_23143);
and U23630 (N_23630,N_23420,N_23490);
and U23631 (N_23631,N_23228,N_23360);
or U23632 (N_23632,N_23078,N_23477);
nor U23633 (N_23633,N_23355,N_23491);
and U23634 (N_23634,N_23021,N_23044);
or U23635 (N_23635,N_23071,N_23474);
or U23636 (N_23636,N_23077,N_23327);
or U23637 (N_23637,N_23395,N_23115);
and U23638 (N_23638,N_23150,N_23183);
or U23639 (N_23639,N_23003,N_23053);
nand U23640 (N_23640,N_23447,N_23470);
xor U23641 (N_23641,N_23473,N_23351);
xnor U23642 (N_23642,N_23315,N_23052);
xor U23643 (N_23643,N_23088,N_23275);
and U23644 (N_23644,N_23160,N_23209);
xnor U23645 (N_23645,N_23023,N_23427);
and U23646 (N_23646,N_23328,N_23010);
and U23647 (N_23647,N_23105,N_23218);
and U23648 (N_23648,N_23207,N_23055);
or U23649 (N_23649,N_23127,N_23167);
nand U23650 (N_23650,N_23129,N_23196);
nor U23651 (N_23651,N_23172,N_23229);
or U23652 (N_23652,N_23091,N_23472);
nor U23653 (N_23653,N_23119,N_23179);
nor U23654 (N_23654,N_23157,N_23462);
or U23655 (N_23655,N_23242,N_23186);
and U23656 (N_23656,N_23269,N_23382);
xnor U23657 (N_23657,N_23252,N_23156);
or U23658 (N_23658,N_23397,N_23428);
or U23659 (N_23659,N_23036,N_23265);
nor U23660 (N_23660,N_23135,N_23241);
or U23661 (N_23661,N_23038,N_23277);
nor U23662 (N_23662,N_23497,N_23148);
nand U23663 (N_23663,N_23297,N_23336);
nor U23664 (N_23664,N_23195,N_23024);
xnor U23665 (N_23665,N_23110,N_23076);
and U23666 (N_23666,N_23441,N_23498);
nand U23667 (N_23667,N_23368,N_23480);
xnor U23668 (N_23668,N_23227,N_23206);
and U23669 (N_23669,N_23273,N_23307);
nor U23670 (N_23670,N_23370,N_23323);
nand U23671 (N_23671,N_23284,N_23222);
xnor U23672 (N_23672,N_23311,N_23278);
or U23673 (N_23673,N_23214,N_23060);
xor U23674 (N_23674,N_23051,N_23449);
xor U23675 (N_23675,N_23087,N_23356);
xor U23676 (N_23676,N_23200,N_23014);
nor U23677 (N_23677,N_23033,N_23020);
or U23678 (N_23678,N_23301,N_23296);
xor U23679 (N_23679,N_23163,N_23326);
nand U23680 (N_23680,N_23444,N_23193);
and U23681 (N_23681,N_23446,N_23063);
or U23682 (N_23682,N_23348,N_23361);
or U23683 (N_23683,N_23331,N_23431);
and U23684 (N_23684,N_23488,N_23136);
nand U23685 (N_23685,N_23247,N_23002);
or U23686 (N_23686,N_23392,N_23168);
xor U23687 (N_23687,N_23486,N_23396);
nand U23688 (N_23688,N_23202,N_23138);
nand U23689 (N_23689,N_23413,N_23457);
nand U23690 (N_23690,N_23065,N_23075);
nor U23691 (N_23691,N_23101,N_23287);
nor U23692 (N_23692,N_23034,N_23192);
or U23693 (N_23693,N_23320,N_23171);
and U23694 (N_23694,N_23308,N_23255);
nand U23695 (N_23695,N_23286,N_23478);
nand U23696 (N_23696,N_23144,N_23174);
or U23697 (N_23697,N_23357,N_23492);
xor U23698 (N_23698,N_23040,N_23412);
xnor U23699 (N_23699,N_23314,N_23432);
or U23700 (N_23700,N_23245,N_23430);
xor U23701 (N_23701,N_23494,N_23001);
and U23702 (N_23702,N_23112,N_23177);
or U23703 (N_23703,N_23468,N_23215);
nor U23704 (N_23704,N_23068,N_23131);
xnor U23705 (N_23705,N_23178,N_23007);
nor U23706 (N_23706,N_23104,N_23401);
or U23707 (N_23707,N_23000,N_23004);
or U23708 (N_23708,N_23176,N_23354);
nor U23709 (N_23709,N_23118,N_23099);
xnor U23710 (N_23710,N_23291,N_23411);
nor U23711 (N_23711,N_23288,N_23276);
and U23712 (N_23712,N_23387,N_23175);
xnor U23713 (N_23713,N_23012,N_23239);
or U23714 (N_23714,N_23310,N_23081);
nor U23715 (N_23715,N_23335,N_23416);
xor U23716 (N_23716,N_23134,N_23254);
nor U23717 (N_23717,N_23199,N_23028);
or U23718 (N_23718,N_23190,N_23343);
nor U23719 (N_23719,N_23440,N_23465);
nor U23720 (N_23720,N_23240,N_23084);
nor U23721 (N_23721,N_23410,N_23142);
nand U23722 (N_23722,N_23151,N_23429);
or U23723 (N_23723,N_23454,N_23080);
xnor U23724 (N_23724,N_23094,N_23400);
or U23725 (N_23725,N_23383,N_23189);
nor U23726 (N_23726,N_23035,N_23017);
and U23727 (N_23727,N_23479,N_23185);
and U23728 (N_23728,N_23074,N_23495);
and U23729 (N_23729,N_23031,N_23414);
xor U23730 (N_23730,N_23285,N_23057);
nor U23731 (N_23731,N_23146,N_23482);
nor U23732 (N_23732,N_23139,N_23381);
and U23733 (N_23733,N_23230,N_23448);
nor U23734 (N_23734,N_23489,N_23451);
nor U23735 (N_23735,N_23485,N_23402);
nand U23736 (N_23736,N_23111,N_23321);
and U23737 (N_23737,N_23425,N_23238);
nand U23738 (N_23738,N_23219,N_23388);
xnor U23739 (N_23739,N_23103,N_23107);
nor U23740 (N_23740,N_23187,N_23261);
and U23741 (N_23741,N_23258,N_23236);
nand U23742 (N_23742,N_23095,N_23379);
or U23743 (N_23743,N_23108,N_23378);
nor U23744 (N_23744,N_23249,N_23280);
xor U23745 (N_23745,N_23302,N_23059);
nor U23746 (N_23746,N_23009,N_23246);
and U23747 (N_23747,N_23384,N_23145);
nand U23748 (N_23748,N_23338,N_23212);
xnor U23749 (N_23749,N_23153,N_23113);
nand U23750 (N_23750,N_23305,N_23399);
nor U23751 (N_23751,N_23130,N_23354);
nand U23752 (N_23752,N_23057,N_23386);
nand U23753 (N_23753,N_23353,N_23363);
nor U23754 (N_23754,N_23437,N_23245);
or U23755 (N_23755,N_23485,N_23084);
or U23756 (N_23756,N_23049,N_23455);
or U23757 (N_23757,N_23332,N_23168);
and U23758 (N_23758,N_23010,N_23371);
or U23759 (N_23759,N_23433,N_23347);
xnor U23760 (N_23760,N_23314,N_23460);
nand U23761 (N_23761,N_23227,N_23380);
nand U23762 (N_23762,N_23410,N_23431);
nor U23763 (N_23763,N_23122,N_23407);
xnor U23764 (N_23764,N_23105,N_23426);
and U23765 (N_23765,N_23297,N_23010);
nor U23766 (N_23766,N_23083,N_23469);
nor U23767 (N_23767,N_23419,N_23334);
and U23768 (N_23768,N_23280,N_23107);
or U23769 (N_23769,N_23352,N_23070);
and U23770 (N_23770,N_23044,N_23271);
and U23771 (N_23771,N_23006,N_23353);
nand U23772 (N_23772,N_23117,N_23196);
nor U23773 (N_23773,N_23382,N_23437);
nand U23774 (N_23774,N_23229,N_23145);
or U23775 (N_23775,N_23233,N_23173);
nor U23776 (N_23776,N_23086,N_23142);
xor U23777 (N_23777,N_23075,N_23098);
and U23778 (N_23778,N_23267,N_23365);
xor U23779 (N_23779,N_23391,N_23101);
and U23780 (N_23780,N_23263,N_23019);
and U23781 (N_23781,N_23083,N_23029);
and U23782 (N_23782,N_23253,N_23193);
and U23783 (N_23783,N_23276,N_23261);
nor U23784 (N_23784,N_23063,N_23388);
nand U23785 (N_23785,N_23316,N_23428);
nor U23786 (N_23786,N_23094,N_23078);
and U23787 (N_23787,N_23000,N_23047);
nand U23788 (N_23788,N_23267,N_23492);
and U23789 (N_23789,N_23233,N_23097);
or U23790 (N_23790,N_23480,N_23089);
nand U23791 (N_23791,N_23189,N_23093);
nor U23792 (N_23792,N_23384,N_23124);
nand U23793 (N_23793,N_23071,N_23229);
or U23794 (N_23794,N_23365,N_23428);
xnor U23795 (N_23795,N_23438,N_23161);
nand U23796 (N_23796,N_23184,N_23277);
nand U23797 (N_23797,N_23221,N_23157);
and U23798 (N_23798,N_23227,N_23162);
nand U23799 (N_23799,N_23499,N_23467);
nand U23800 (N_23800,N_23394,N_23097);
nand U23801 (N_23801,N_23255,N_23281);
or U23802 (N_23802,N_23368,N_23357);
and U23803 (N_23803,N_23165,N_23053);
and U23804 (N_23804,N_23058,N_23398);
and U23805 (N_23805,N_23456,N_23237);
or U23806 (N_23806,N_23494,N_23474);
or U23807 (N_23807,N_23321,N_23427);
or U23808 (N_23808,N_23305,N_23010);
nor U23809 (N_23809,N_23056,N_23355);
xnor U23810 (N_23810,N_23448,N_23107);
xnor U23811 (N_23811,N_23004,N_23489);
and U23812 (N_23812,N_23270,N_23014);
or U23813 (N_23813,N_23129,N_23051);
nand U23814 (N_23814,N_23134,N_23277);
or U23815 (N_23815,N_23447,N_23287);
or U23816 (N_23816,N_23411,N_23345);
xor U23817 (N_23817,N_23468,N_23251);
and U23818 (N_23818,N_23317,N_23404);
nor U23819 (N_23819,N_23095,N_23014);
xnor U23820 (N_23820,N_23479,N_23443);
and U23821 (N_23821,N_23049,N_23317);
xnor U23822 (N_23822,N_23182,N_23308);
nor U23823 (N_23823,N_23309,N_23076);
and U23824 (N_23824,N_23494,N_23308);
or U23825 (N_23825,N_23143,N_23124);
xor U23826 (N_23826,N_23384,N_23033);
or U23827 (N_23827,N_23344,N_23011);
nand U23828 (N_23828,N_23309,N_23469);
xnor U23829 (N_23829,N_23444,N_23152);
nor U23830 (N_23830,N_23273,N_23434);
nand U23831 (N_23831,N_23481,N_23119);
xor U23832 (N_23832,N_23092,N_23215);
nand U23833 (N_23833,N_23032,N_23277);
nand U23834 (N_23834,N_23239,N_23211);
and U23835 (N_23835,N_23004,N_23360);
and U23836 (N_23836,N_23453,N_23414);
and U23837 (N_23837,N_23100,N_23007);
nand U23838 (N_23838,N_23401,N_23433);
xnor U23839 (N_23839,N_23177,N_23169);
xor U23840 (N_23840,N_23056,N_23292);
xor U23841 (N_23841,N_23048,N_23088);
or U23842 (N_23842,N_23373,N_23095);
or U23843 (N_23843,N_23485,N_23124);
xnor U23844 (N_23844,N_23273,N_23496);
nor U23845 (N_23845,N_23003,N_23071);
nor U23846 (N_23846,N_23491,N_23184);
nor U23847 (N_23847,N_23322,N_23497);
or U23848 (N_23848,N_23262,N_23455);
nor U23849 (N_23849,N_23256,N_23407);
nand U23850 (N_23850,N_23252,N_23270);
and U23851 (N_23851,N_23255,N_23161);
nor U23852 (N_23852,N_23137,N_23265);
nor U23853 (N_23853,N_23448,N_23085);
nor U23854 (N_23854,N_23248,N_23489);
xor U23855 (N_23855,N_23306,N_23200);
or U23856 (N_23856,N_23318,N_23443);
nand U23857 (N_23857,N_23358,N_23021);
xor U23858 (N_23858,N_23239,N_23434);
nand U23859 (N_23859,N_23043,N_23045);
xor U23860 (N_23860,N_23306,N_23291);
or U23861 (N_23861,N_23019,N_23343);
nand U23862 (N_23862,N_23059,N_23136);
and U23863 (N_23863,N_23345,N_23158);
xor U23864 (N_23864,N_23476,N_23053);
xor U23865 (N_23865,N_23141,N_23025);
nor U23866 (N_23866,N_23401,N_23031);
xnor U23867 (N_23867,N_23488,N_23228);
nand U23868 (N_23868,N_23125,N_23356);
xnor U23869 (N_23869,N_23064,N_23179);
or U23870 (N_23870,N_23399,N_23128);
or U23871 (N_23871,N_23162,N_23013);
and U23872 (N_23872,N_23020,N_23058);
xor U23873 (N_23873,N_23037,N_23176);
or U23874 (N_23874,N_23045,N_23133);
xor U23875 (N_23875,N_23117,N_23404);
nor U23876 (N_23876,N_23366,N_23070);
and U23877 (N_23877,N_23026,N_23258);
or U23878 (N_23878,N_23366,N_23104);
or U23879 (N_23879,N_23416,N_23465);
xnor U23880 (N_23880,N_23433,N_23369);
nand U23881 (N_23881,N_23390,N_23013);
nand U23882 (N_23882,N_23433,N_23133);
nand U23883 (N_23883,N_23005,N_23083);
and U23884 (N_23884,N_23253,N_23144);
xnor U23885 (N_23885,N_23156,N_23250);
xnor U23886 (N_23886,N_23378,N_23194);
xnor U23887 (N_23887,N_23167,N_23095);
and U23888 (N_23888,N_23359,N_23386);
or U23889 (N_23889,N_23463,N_23400);
and U23890 (N_23890,N_23106,N_23392);
xor U23891 (N_23891,N_23025,N_23314);
nor U23892 (N_23892,N_23331,N_23379);
or U23893 (N_23893,N_23361,N_23383);
and U23894 (N_23894,N_23275,N_23031);
or U23895 (N_23895,N_23229,N_23311);
xnor U23896 (N_23896,N_23238,N_23406);
and U23897 (N_23897,N_23249,N_23408);
nor U23898 (N_23898,N_23224,N_23228);
nor U23899 (N_23899,N_23016,N_23374);
xnor U23900 (N_23900,N_23250,N_23368);
xor U23901 (N_23901,N_23481,N_23160);
or U23902 (N_23902,N_23197,N_23223);
and U23903 (N_23903,N_23404,N_23471);
nand U23904 (N_23904,N_23233,N_23481);
xor U23905 (N_23905,N_23396,N_23459);
nor U23906 (N_23906,N_23242,N_23475);
xnor U23907 (N_23907,N_23439,N_23222);
or U23908 (N_23908,N_23107,N_23128);
or U23909 (N_23909,N_23179,N_23112);
nor U23910 (N_23910,N_23470,N_23255);
nor U23911 (N_23911,N_23274,N_23328);
or U23912 (N_23912,N_23097,N_23413);
xor U23913 (N_23913,N_23282,N_23251);
xnor U23914 (N_23914,N_23235,N_23188);
or U23915 (N_23915,N_23373,N_23478);
or U23916 (N_23916,N_23306,N_23133);
nor U23917 (N_23917,N_23075,N_23050);
and U23918 (N_23918,N_23204,N_23373);
and U23919 (N_23919,N_23384,N_23263);
and U23920 (N_23920,N_23142,N_23302);
and U23921 (N_23921,N_23331,N_23257);
and U23922 (N_23922,N_23329,N_23340);
nor U23923 (N_23923,N_23115,N_23370);
nand U23924 (N_23924,N_23064,N_23182);
and U23925 (N_23925,N_23105,N_23008);
nand U23926 (N_23926,N_23354,N_23351);
xnor U23927 (N_23927,N_23478,N_23088);
xor U23928 (N_23928,N_23152,N_23005);
and U23929 (N_23929,N_23416,N_23486);
and U23930 (N_23930,N_23064,N_23091);
nand U23931 (N_23931,N_23475,N_23315);
nand U23932 (N_23932,N_23199,N_23202);
and U23933 (N_23933,N_23054,N_23036);
nand U23934 (N_23934,N_23358,N_23400);
xor U23935 (N_23935,N_23483,N_23017);
nor U23936 (N_23936,N_23167,N_23499);
and U23937 (N_23937,N_23177,N_23037);
xnor U23938 (N_23938,N_23200,N_23296);
or U23939 (N_23939,N_23147,N_23264);
and U23940 (N_23940,N_23323,N_23347);
and U23941 (N_23941,N_23313,N_23483);
and U23942 (N_23942,N_23266,N_23213);
nor U23943 (N_23943,N_23322,N_23164);
or U23944 (N_23944,N_23350,N_23117);
nor U23945 (N_23945,N_23285,N_23329);
nor U23946 (N_23946,N_23405,N_23496);
xor U23947 (N_23947,N_23347,N_23212);
or U23948 (N_23948,N_23372,N_23355);
xor U23949 (N_23949,N_23185,N_23092);
nand U23950 (N_23950,N_23455,N_23229);
or U23951 (N_23951,N_23152,N_23140);
nor U23952 (N_23952,N_23279,N_23481);
or U23953 (N_23953,N_23463,N_23405);
and U23954 (N_23954,N_23418,N_23169);
xor U23955 (N_23955,N_23152,N_23393);
or U23956 (N_23956,N_23342,N_23293);
xnor U23957 (N_23957,N_23315,N_23219);
xnor U23958 (N_23958,N_23211,N_23314);
xor U23959 (N_23959,N_23267,N_23382);
nor U23960 (N_23960,N_23103,N_23499);
and U23961 (N_23961,N_23140,N_23184);
or U23962 (N_23962,N_23126,N_23011);
nand U23963 (N_23963,N_23298,N_23055);
or U23964 (N_23964,N_23337,N_23459);
and U23965 (N_23965,N_23494,N_23038);
and U23966 (N_23966,N_23315,N_23135);
or U23967 (N_23967,N_23408,N_23338);
nand U23968 (N_23968,N_23153,N_23071);
nand U23969 (N_23969,N_23213,N_23468);
nand U23970 (N_23970,N_23263,N_23325);
nor U23971 (N_23971,N_23072,N_23032);
and U23972 (N_23972,N_23313,N_23208);
and U23973 (N_23973,N_23368,N_23397);
or U23974 (N_23974,N_23263,N_23153);
xnor U23975 (N_23975,N_23033,N_23244);
or U23976 (N_23976,N_23195,N_23267);
or U23977 (N_23977,N_23328,N_23038);
and U23978 (N_23978,N_23434,N_23120);
and U23979 (N_23979,N_23027,N_23466);
nor U23980 (N_23980,N_23391,N_23157);
or U23981 (N_23981,N_23167,N_23091);
xor U23982 (N_23982,N_23199,N_23298);
and U23983 (N_23983,N_23042,N_23119);
xnor U23984 (N_23984,N_23482,N_23266);
and U23985 (N_23985,N_23148,N_23327);
and U23986 (N_23986,N_23483,N_23317);
and U23987 (N_23987,N_23393,N_23125);
nand U23988 (N_23988,N_23055,N_23282);
nand U23989 (N_23989,N_23342,N_23358);
or U23990 (N_23990,N_23047,N_23159);
nor U23991 (N_23991,N_23136,N_23288);
xor U23992 (N_23992,N_23327,N_23060);
nor U23993 (N_23993,N_23113,N_23480);
nor U23994 (N_23994,N_23436,N_23418);
xor U23995 (N_23995,N_23401,N_23170);
xnor U23996 (N_23996,N_23424,N_23230);
nor U23997 (N_23997,N_23248,N_23444);
or U23998 (N_23998,N_23177,N_23294);
and U23999 (N_23999,N_23184,N_23444);
nor U24000 (N_24000,N_23669,N_23577);
and U24001 (N_24001,N_23798,N_23737);
or U24002 (N_24002,N_23827,N_23627);
xor U24003 (N_24003,N_23881,N_23565);
xnor U24004 (N_24004,N_23712,N_23569);
nand U24005 (N_24005,N_23987,N_23804);
nand U24006 (N_24006,N_23525,N_23620);
xor U24007 (N_24007,N_23631,N_23920);
and U24008 (N_24008,N_23666,N_23986);
nand U24009 (N_24009,N_23951,N_23801);
and U24010 (N_24010,N_23658,N_23865);
nand U24011 (N_24011,N_23518,N_23610);
nand U24012 (N_24012,N_23958,N_23901);
nor U24013 (N_24013,N_23813,N_23953);
nand U24014 (N_24014,N_23899,N_23926);
xor U24015 (N_24015,N_23571,N_23811);
nor U24016 (N_24016,N_23786,N_23819);
nand U24017 (N_24017,N_23719,N_23547);
nand U24018 (N_24018,N_23529,N_23661);
or U24019 (N_24019,N_23607,N_23623);
xor U24020 (N_24020,N_23932,N_23918);
or U24021 (N_24021,N_23853,N_23982);
or U24022 (N_24022,N_23612,N_23676);
and U24023 (N_24023,N_23989,N_23649);
nand U24024 (N_24024,N_23678,N_23578);
nand U24025 (N_24025,N_23904,N_23534);
nand U24026 (N_24026,N_23749,N_23916);
and U24027 (N_24027,N_23628,N_23775);
or U24028 (N_24028,N_23929,N_23652);
and U24029 (N_24029,N_23934,N_23815);
or U24030 (N_24030,N_23734,N_23871);
nand U24031 (N_24031,N_23657,N_23966);
nor U24032 (N_24032,N_23803,N_23875);
nor U24033 (N_24033,N_23823,N_23973);
and U24034 (N_24034,N_23992,N_23595);
nand U24035 (N_24035,N_23878,N_23683);
and U24036 (N_24036,N_23614,N_23931);
or U24037 (N_24037,N_23852,N_23639);
nor U24038 (N_24038,N_23945,N_23507);
nand U24039 (N_24039,N_23670,N_23651);
nand U24040 (N_24040,N_23630,N_23706);
xor U24041 (N_24041,N_23511,N_23758);
nor U24042 (N_24042,N_23519,N_23751);
and U24043 (N_24043,N_23622,N_23778);
xor U24044 (N_24044,N_23842,N_23655);
nand U24045 (N_24045,N_23910,N_23856);
xnor U24046 (N_24046,N_23956,N_23922);
and U24047 (N_24047,N_23543,N_23641);
nor U24048 (N_24048,N_23545,N_23959);
and U24049 (N_24049,N_23830,N_23917);
and U24050 (N_24050,N_23691,N_23807);
or U24051 (N_24051,N_23558,N_23667);
or U24052 (N_24052,N_23869,N_23996);
and U24053 (N_24053,N_23841,N_23562);
or U24054 (N_24054,N_23732,N_23970);
nor U24055 (N_24055,N_23660,N_23701);
nand U24056 (N_24056,N_23747,N_23559);
nor U24057 (N_24057,N_23937,N_23760);
and U24058 (N_24058,N_23733,N_23849);
and U24059 (N_24059,N_23840,N_23898);
or U24060 (N_24060,N_23717,N_23727);
nand U24061 (N_24061,N_23697,N_23724);
xnor U24062 (N_24062,N_23995,N_23596);
nand U24063 (N_24063,N_23629,N_23817);
or U24064 (N_24064,N_23527,N_23556);
or U24065 (N_24065,N_23768,N_23574);
xor U24066 (N_24066,N_23709,N_23785);
or U24067 (N_24067,N_23924,N_23650);
and U24068 (N_24068,N_23990,N_23592);
xor U24069 (N_24069,N_23573,N_23954);
or U24070 (N_24070,N_23557,N_23776);
and U24071 (N_24071,N_23928,N_23561);
or U24072 (N_24072,N_23647,N_23590);
xnor U24073 (N_24073,N_23673,N_23598);
xor U24074 (N_24074,N_23605,N_23796);
nor U24075 (N_24075,N_23696,N_23908);
xnor U24076 (N_24076,N_23707,N_23718);
nor U24077 (N_24077,N_23984,N_23548);
or U24078 (N_24078,N_23566,N_23792);
nor U24079 (N_24079,N_23551,N_23584);
or U24080 (N_24080,N_23862,N_23603);
nand U24081 (N_24081,N_23633,N_23714);
nor U24082 (N_24082,N_23788,N_23765);
and U24083 (N_24083,N_23762,N_23872);
nor U24084 (N_24084,N_23618,N_23761);
xnor U24085 (N_24085,N_23824,N_23756);
nand U24086 (N_24086,N_23589,N_23675);
nand U24087 (N_24087,N_23742,N_23748);
nand U24088 (N_24088,N_23820,N_23812);
xnor U24089 (N_24089,N_23593,N_23799);
xnor U24090 (N_24090,N_23602,N_23914);
or U24091 (N_24091,N_23940,N_23905);
nand U24092 (N_24092,N_23983,N_23594);
nand U24093 (N_24093,N_23695,N_23539);
or U24094 (N_24094,N_23848,N_23857);
nand U24095 (N_24095,N_23831,N_23930);
nand U24096 (N_24096,N_23975,N_23874);
and U24097 (N_24097,N_23524,N_23542);
nand U24098 (N_24098,N_23846,N_23659);
nor U24099 (N_24099,N_23893,N_23763);
and U24100 (N_24100,N_23700,N_23526);
and U24101 (N_24101,N_23743,N_23685);
nand U24102 (N_24102,N_23645,N_23535);
nand U24103 (N_24103,N_23994,N_23988);
and U24104 (N_24104,N_23604,N_23611);
nand U24105 (N_24105,N_23814,N_23516);
or U24106 (N_24106,N_23662,N_23962);
and U24107 (N_24107,N_23721,N_23503);
nor U24108 (N_24108,N_23774,N_23771);
nand U24109 (N_24109,N_23508,N_23588);
nand U24110 (N_24110,N_23949,N_23591);
or U24111 (N_24111,N_23541,N_23780);
or U24112 (N_24112,N_23671,N_23863);
or U24113 (N_24113,N_23619,N_23836);
nand U24114 (N_24114,N_23713,N_23907);
and U24115 (N_24115,N_23606,N_23501);
or U24116 (N_24116,N_23883,N_23575);
nor U24117 (N_24117,N_23843,N_23876);
or U24118 (N_24118,N_23802,N_23895);
xor U24119 (N_24119,N_23553,N_23923);
and U24120 (N_24120,N_23927,N_23613);
nand U24121 (N_24121,N_23818,N_23838);
nand U24122 (N_24122,N_23504,N_23757);
nor U24123 (N_24123,N_23935,N_23894);
nand U24124 (N_24124,N_23555,N_23560);
or U24125 (N_24125,N_23939,N_23759);
or U24126 (N_24126,N_23933,N_23528);
nand U24127 (N_24127,N_23769,N_23624);
nor U24128 (N_24128,N_23514,N_23773);
and U24129 (N_24129,N_23617,N_23506);
or U24130 (N_24130,N_23710,N_23942);
and U24131 (N_24131,N_23581,N_23726);
or U24132 (N_24132,N_23510,N_23826);
nor U24133 (N_24133,N_23728,N_23882);
nand U24134 (N_24134,N_23672,N_23698);
nand U24135 (N_24135,N_23580,N_23690);
nor U24136 (N_24136,N_23616,N_23750);
and U24137 (N_24137,N_23889,N_23896);
nand U24138 (N_24138,N_23832,N_23708);
xnor U24139 (N_24139,N_23808,N_23646);
and U24140 (N_24140,N_23974,N_23921);
nor U24141 (N_24141,N_23563,N_23500);
nor U24142 (N_24142,N_23654,N_23746);
or U24143 (N_24143,N_23638,N_23828);
xnor U24144 (N_24144,N_23781,N_23550);
and U24145 (N_24145,N_23834,N_23621);
nor U24146 (N_24146,N_23900,N_23991);
or U24147 (N_24147,N_23665,N_23586);
nor U24148 (N_24148,N_23999,N_23925);
nor U24149 (N_24149,N_23854,N_23972);
xnor U24150 (N_24150,N_23740,N_23998);
xnor U24151 (N_24151,N_23797,N_23608);
and U24152 (N_24152,N_23944,N_23520);
nor U24153 (N_24153,N_23829,N_23766);
or U24154 (N_24154,N_23736,N_23770);
and U24155 (N_24155,N_23686,N_23694);
nand U24156 (N_24156,N_23681,N_23936);
nand U24157 (N_24157,N_23833,N_23976);
or U24158 (N_24158,N_23699,N_23967);
and U24159 (N_24159,N_23585,N_23582);
nor U24160 (N_24160,N_23980,N_23816);
and U24161 (N_24161,N_23656,N_23509);
xor U24162 (N_24162,N_23689,N_23806);
nor U24163 (N_24163,N_23674,N_23892);
and U24164 (N_24164,N_23601,N_23725);
and U24165 (N_24165,N_23947,N_23502);
and U24166 (N_24166,N_23955,N_23512);
nor U24167 (N_24167,N_23861,N_23679);
nand U24168 (N_24168,N_23653,N_23789);
or U24169 (N_24169,N_23723,N_23552);
xnor U24170 (N_24170,N_23523,N_23570);
and U24171 (N_24171,N_23777,N_23731);
and U24172 (N_24172,N_23704,N_23533);
nor U24173 (N_24173,N_23784,N_23885);
nand U24174 (N_24174,N_23549,N_23783);
xor U24175 (N_24175,N_23821,N_23682);
xnor U24176 (N_24176,N_23730,N_23779);
nand U24177 (N_24177,N_23576,N_23978);
and U24178 (N_24178,N_23741,N_23615);
nand U24179 (N_24179,N_23868,N_23755);
nand U24180 (N_24180,N_23715,N_23851);
nand U24181 (N_24181,N_23782,N_23952);
and U24182 (N_24182,N_23993,N_23625);
and U24183 (N_24183,N_23567,N_23963);
xnor U24184 (N_24184,N_23720,N_23795);
xor U24185 (N_24185,N_23716,N_23521);
and U24186 (N_24186,N_23845,N_23583);
or U24187 (N_24187,N_23635,N_23703);
and U24188 (N_24188,N_23879,N_23791);
or U24189 (N_24189,N_23810,N_23711);
xnor U24190 (N_24190,N_23738,N_23825);
nor U24191 (N_24191,N_23637,N_23568);
nor U24192 (N_24192,N_23764,N_23702);
and U24193 (N_24193,N_23544,N_23950);
xnor U24194 (N_24194,N_23870,N_23964);
nor U24195 (N_24195,N_23961,N_23572);
and U24196 (N_24196,N_23536,N_23981);
or U24197 (N_24197,N_23729,N_23579);
xor U24198 (N_24198,N_23599,N_23767);
or U24199 (N_24199,N_23897,N_23902);
nor U24200 (N_24200,N_23587,N_23844);
xor U24201 (N_24201,N_23839,N_23909);
and U24202 (N_24202,N_23919,N_23546);
xnor U24203 (N_24203,N_23906,N_23858);
xnor U24204 (N_24204,N_23877,N_23943);
nor U24205 (N_24205,N_23886,N_23739);
or U24206 (N_24206,N_23687,N_23705);
xor U24207 (N_24207,N_23693,N_23971);
nand U24208 (N_24208,N_23684,N_23867);
nor U24209 (N_24209,N_23754,N_23985);
and U24210 (N_24210,N_23977,N_23517);
nand U24211 (N_24211,N_23847,N_23644);
nor U24212 (N_24212,N_23793,N_23745);
and U24213 (N_24213,N_23634,N_23888);
xor U24214 (N_24214,N_23790,N_23880);
xor U24215 (N_24215,N_23941,N_23532);
nor U24216 (N_24216,N_23538,N_23969);
xnor U24217 (N_24217,N_23968,N_23513);
nor U24218 (N_24218,N_23636,N_23668);
or U24219 (N_24219,N_23866,N_23864);
nor U24220 (N_24220,N_23855,N_23794);
or U24221 (N_24221,N_23787,N_23859);
nor U24222 (N_24222,N_23688,N_23822);
or U24223 (N_24223,N_23522,N_23531);
nand U24224 (N_24224,N_23997,N_23890);
nand U24225 (N_24225,N_23640,N_23692);
nand U24226 (N_24226,N_23643,N_23609);
xnor U24227 (N_24227,N_23505,N_23744);
nand U24228 (N_24228,N_23772,N_23753);
nor U24229 (N_24229,N_23597,N_23915);
and U24230 (N_24230,N_23884,N_23663);
xnor U24231 (N_24231,N_23554,N_23946);
nand U24232 (N_24232,N_23515,N_23887);
xnor U24233 (N_24233,N_23537,N_23735);
xnor U24234 (N_24234,N_23664,N_23648);
xnor U24235 (N_24235,N_23600,N_23809);
xor U24236 (N_24236,N_23800,N_23873);
nand U24237 (N_24237,N_23913,N_23957);
xnor U24238 (N_24238,N_23626,N_23677);
nand U24239 (N_24239,N_23850,N_23530);
or U24240 (N_24240,N_23632,N_23979);
and U24241 (N_24241,N_23835,N_23805);
nand U24242 (N_24242,N_23564,N_23948);
or U24243 (N_24243,N_23911,N_23860);
or U24244 (N_24244,N_23965,N_23837);
nand U24245 (N_24245,N_23680,N_23642);
xnor U24246 (N_24246,N_23722,N_23938);
and U24247 (N_24247,N_23903,N_23891);
nor U24248 (N_24248,N_23912,N_23540);
nand U24249 (N_24249,N_23752,N_23960);
nor U24250 (N_24250,N_23823,N_23699);
nand U24251 (N_24251,N_23872,N_23907);
xor U24252 (N_24252,N_23701,N_23898);
nand U24253 (N_24253,N_23862,N_23912);
or U24254 (N_24254,N_23750,N_23589);
nor U24255 (N_24255,N_23627,N_23565);
and U24256 (N_24256,N_23824,N_23594);
nor U24257 (N_24257,N_23866,N_23718);
nor U24258 (N_24258,N_23828,N_23504);
nand U24259 (N_24259,N_23886,N_23575);
nand U24260 (N_24260,N_23959,N_23553);
nor U24261 (N_24261,N_23658,N_23767);
nor U24262 (N_24262,N_23826,N_23935);
nand U24263 (N_24263,N_23665,N_23843);
nand U24264 (N_24264,N_23801,N_23880);
xnor U24265 (N_24265,N_23754,N_23967);
nand U24266 (N_24266,N_23653,N_23693);
or U24267 (N_24267,N_23847,N_23813);
nor U24268 (N_24268,N_23869,N_23615);
or U24269 (N_24269,N_23706,N_23574);
and U24270 (N_24270,N_23964,N_23685);
and U24271 (N_24271,N_23950,N_23563);
nand U24272 (N_24272,N_23928,N_23959);
and U24273 (N_24273,N_23902,N_23673);
or U24274 (N_24274,N_23626,N_23785);
nand U24275 (N_24275,N_23789,N_23956);
and U24276 (N_24276,N_23749,N_23543);
nor U24277 (N_24277,N_23710,N_23653);
or U24278 (N_24278,N_23673,N_23746);
and U24279 (N_24279,N_23930,N_23978);
nand U24280 (N_24280,N_23829,N_23817);
nor U24281 (N_24281,N_23996,N_23509);
xnor U24282 (N_24282,N_23546,N_23836);
or U24283 (N_24283,N_23969,N_23942);
and U24284 (N_24284,N_23995,N_23775);
or U24285 (N_24285,N_23905,N_23972);
xnor U24286 (N_24286,N_23939,N_23757);
nor U24287 (N_24287,N_23594,N_23734);
and U24288 (N_24288,N_23912,N_23559);
or U24289 (N_24289,N_23593,N_23827);
or U24290 (N_24290,N_23847,N_23536);
and U24291 (N_24291,N_23929,N_23671);
and U24292 (N_24292,N_23673,N_23864);
or U24293 (N_24293,N_23727,N_23678);
or U24294 (N_24294,N_23678,N_23700);
and U24295 (N_24295,N_23641,N_23691);
and U24296 (N_24296,N_23791,N_23971);
or U24297 (N_24297,N_23792,N_23876);
and U24298 (N_24298,N_23833,N_23929);
xnor U24299 (N_24299,N_23766,N_23941);
nor U24300 (N_24300,N_23799,N_23785);
and U24301 (N_24301,N_23875,N_23621);
nand U24302 (N_24302,N_23691,N_23661);
nand U24303 (N_24303,N_23665,N_23707);
nand U24304 (N_24304,N_23646,N_23771);
xor U24305 (N_24305,N_23705,N_23775);
xor U24306 (N_24306,N_23534,N_23814);
or U24307 (N_24307,N_23725,N_23539);
and U24308 (N_24308,N_23722,N_23808);
and U24309 (N_24309,N_23648,N_23850);
xnor U24310 (N_24310,N_23990,N_23826);
nand U24311 (N_24311,N_23688,N_23607);
xor U24312 (N_24312,N_23635,N_23869);
nand U24313 (N_24313,N_23522,N_23963);
nand U24314 (N_24314,N_23584,N_23661);
nor U24315 (N_24315,N_23876,N_23911);
nor U24316 (N_24316,N_23638,N_23586);
or U24317 (N_24317,N_23567,N_23826);
nand U24318 (N_24318,N_23607,N_23518);
nand U24319 (N_24319,N_23532,N_23772);
nand U24320 (N_24320,N_23663,N_23622);
or U24321 (N_24321,N_23502,N_23553);
or U24322 (N_24322,N_23901,N_23962);
xnor U24323 (N_24323,N_23836,N_23755);
and U24324 (N_24324,N_23707,N_23616);
nor U24325 (N_24325,N_23874,N_23928);
nor U24326 (N_24326,N_23982,N_23566);
xor U24327 (N_24327,N_23898,N_23827);
nand U24328 (N_24328,N_23601,N_23717);
or U24329 (N_24329,N_23938,N_23640);
nor U24330 (N_24330,N_23853,N_23640);
and U24331 (N_24331,N_23548,N_23736);
xnor U24332 (N_24332,N_23743,N_23880);
nor U24333 (N_24333,N_23763,N_23889);
or U24334 (N_24334,N_23646,N_23911);
nand U24335 (N_24335,N_23728,N_23779);
or U24336 (N_24336,N_23878,N_23612);
nor U24337 (N_24337,N_23668,N_23557);
or U24338 (N_24338,N_23893,N_23690);
and U24339 (N_24339,N_23972,N_23561);
or U24340 (N_24340,N_23726,N_23712);
xnor U24341 (N_24341,N_23626,N_23515);
nand U24342 (N_24342,N_23723,N_23836);
or U24343 (N_24343,N_23861,N_23848);
nand U24344 (N_24344,N_23863,N_23521);
nor U24345 (N_24345,N_23929,N_23961);
xor U24346 (N_24346,N_23882,N_23953);
xor U24347 (N_24347,N_23918,N_23557);
nor U24348 (N_24348,N_23553,N_23963);
xnor U24349 (N_24349,N_23850,N_23920);
nand U24350 (N_24350,N_23652,N_23970);
nor U24351 (N_24351,N_23970,N_23767);
xor U24352 (N_24352,N_23574,N_23751);
or U24353 (N_24353,N_23904,N_23829);
xnor U24354 (N_24354,N_23776,N_23817);
nor U24355 (N_24355,N_23949,N_23907);
and U24356 (N_24356,N_23982,N_23757);
and U24357 (N_24357,N_23718,N_23809);
xor U24358 (N_24358,N_23645,N_23784);
nor U24359 (N_24359,N_23759,N_23796);
or U24360 (N_24360,N_23880,N_23609);
nor U24361 (N_24361,N_23857,N_23995);
nor U24362 (N_24362,N_23838,N_23548);
nor U24363 (N_24363,N_23512,N_23850);
and U24364 (N_24364,N_23519,N_23667);
and U24365 (N_24365,N_23699,N_23719);
nand U24366 (N_24366,N_23704,N_23800);
or U24367 (N_24367,N_23796,N_23692);
xor U24368 (N_24368,N_23648,N_23919);
xnor U24369 (N_24369,N_23708,N_23777);
nand U24370 (N_24370,N_23991,N_23845);
xor U24371 (N_24371,N_23761,N_23646);
nand U24372 (N_24372,N_23886,N_23967);
and U24373 (N_24373,N_23602,N_23562);
and U24374 (N_24374,N_23848,N_23956);
or U24375 (N_24375,N_23524,N_23689);
xnor U24376 (N_24376,N_23639,N_23648);
or U24377 (N_24377,N_23977,N_23803);
or U24378 (N_24378,N_23725,N_23802);
xor U24379 (N_24379,N_23848,N_23654);
xnor U24380 (N_24380,N_23893,N_23744);
nand U24381 (N_24381,N_23619,N_23818);
nand U24382 (N_24382,N_23948,N_23656);
and U24383 (N_24383,N_23615,N_23535);
nand U24384 (N_24384,N_23836,N_23926);
xor U24385 (N_24385,N_23715,N_23506);
xnor U24386 (N_24386,N_23934,N_23643);
and U24387 (N_24387,N_23640,N_23638);
xnor U24388 (N_24388,N_23791,N_23974);
xnor U24389 (N_24389,N_23546,N_23932);
nor U24390 (N_24390,N_23675,N_23822);
nor U24391 (N_24391,N_23889,N_23571);
nor U24392 (N_24392,N_23597,N_23503);
and U24393 (N_24393,N_23504,N_23650);
nand U24394 (N_24394,N_23746,N_23572);
xnor U24395 (N_24395,N_23993,N_23735);
nor U24396 (N_24396,N_23940,N_23956);
nand U24397 (N_24397,N_23873,N_23516);
or U24398 (N_24398,N_23722,N_23614);
nor U24399 (N_24399,N_23843,N_23902);
or U24400 (N_24400,N_23986,N_23863);
nand U24401 (N_24401,N_23741,N_23632);
and U24402 (N_24402,N_23763,N_23810);
nor U24403 (N_24403,N_23837,N_23815);
nor U24404 (N_24404,N_23779,N_23816);
nand U24405 (N_24405,N_23528,N_23789);
and U24406 (N_24406,N_23658,N_23727);
xnor U24407 (N_24407,N_23883,N_23628);
nor U24408 (N_24408,N_23686,N_23769);
and U24409 (N_24409,N_23562,N_23611);
nor U24410 (N_24410,N_23928,N_23696);
xnor U24411 (N_24411,N_23932,N_23617);
or U24412 (N_24412,N_23602,N_23829);
xnor U24413 (N_24413,N_23910,N_23531);
xor U24414 (N_24414,N_23863,N_23902);
xnor U24415 (N_24415,N_23686,N_23679);
nand U24416 (N_24416,N_23864,N_23745);
nor U24417 (N_24417,N_23582,N_23751);
and U24418 (N_24418,N_23861,N_23871);
nand U24419 (N_24419,N_23896,N_23694);
or U24420 (N_24420,N_23911,N_23750);
xnor U24421 (N_24421,N_23633,N_23700);
nor U24422 (N_24422,N_23664,N_23547);
and U24423 (N_24423,N_23836,N_23779);
and U24424 (N_24424,N_23587,N_23665);
xor U24425 (N_24425,N_23594,N_23939);
nor U24426 (N_24426,N_23545,N_23739);
nand U24427 (N_24427,N_23680,N_23688);
nand U24428 (N_24428,N_23955,N_23844);
xor U24429 (N_24429,N_23527,N_23549);
nor U24430 (N_24430,N_23730,N_23925);
nor U24431 (N_24431,N_23888,N_23971);
xnor U24432 (N_24432,N_23920,N_23971);
nor U24433 (N_24433,N_23861,N_23799);
xnor U24434 (N_24434,N_23524,N_23859);
xnor U24435 (N_24435,N_23506,N_23830);
and U24436 (N_24436,N_23653,N_23668);
or U24437 (N_24437,N_23869,N_23752);
or U24438 (N_24438,N_23628,N_23946);
or U24439 (N_24439,N_23681,N_23872);
or U24440 (N_24440,N_23753,N_23766);
and U24441 (N_24441,N_23721,N_23875);
and U24442 (N_24442,N_23686,N_23677);
or U24443 (N_24443,N_23858,N_23709);
nor U24444 (N_24444,N_23812,N_23659);
xor U24445 (N_24445,N_23980,N_23953);
and U24446 (N_24446,N_23804,N_23610);
xor U24447 (N_24447,N_23938,N_23650);
or U24448 (N_24448,N_23628,N_23751);
or U24449 (N_24449,N_23802,N_23869);
xor U24450 (N_24450,N_23709,N_23983);
nand U24451 (N_24451,N_23788,N_23722);
and U24452 (N_24452,N_23623,N_23675);
or U24453 (N_24453,N_23937,N_23649);
or U24454 (N_24454,N_23681,N_23604);
and U24455 (N_24455,N_23874,N_23544);
xnor U24456 (N_24456,N_23742,N_23801);
nor U24457 (N_24457,N_23922,N_23834);
or U24458 (N_24458,N_23603,N_23850);
and U24459 (N_24459,N_23924,N_23767);
or U24460 (N_24460,N_23610,N_23663);
and U24461 (N_24461,N_23788,N_23753);
xor U24462 (N_24462,N_23771,N_23638);
and U24463 (N_24463,N_23910,N_23646);
nor U24464 (N_24464,N_23997,N_23598);
or U24465 (N_24465,N_23857,N_23647);
nand U24466 (N_24466,N_23624,N_23858);
or U24467 (N_24467,N_23912,N_23696);
and U24468 (N_24468,N_23710,N_23533);
and U24469 (N_24469,N_23926,N_23974);
nand U24470 (N_24470,N_23580,N_23669);
nand U24471 (N_24471,N_23680,N_23902);
or U24472 (N_24472,N_23564,N_23646);
xor U24473 (N_24473,N_23717,N_23567);
or U24474 (N_24474,N_23943,N_23922);
or U24475 (N_24475,N_23502,N_23514);
and U24476 (N_24476,N_23970,N_23670);
nor U24477 (N_24477,N_23923,N_23574);
and U24478 (N_24478,N_23803,N_23510);
xor U24479 (N_24479,N_23990,N_23613);
nor U24480 (N_24480,N_23804,N_23855);
or U24481 (N_24481,N_23657,N_23877);
nand U24482 (N_24482,N_23705,N_23972);
xor U24483 (N_24483,N_23685,N_23602);
or U24484 (N_24484,N_23864,N_23651);
nand U24485 (N_24485,N_23992,N_23851);
nand U24486 (N_24486,N_23907,N_23542);
nand U24487 (N_24487,N_23807,N_23778);
nand U24488 (N_24488,N_23991,N_23735);
xor U24489 (N_24489,N_23932,N_23718);
nand U24490 (N_24490,N_23602,N_23982);
nor U24491 (N_24491,N_23554,N_23778);
or U24492 (N_24492,N_23980,N_23732);
and U24493 (N_24493,N_23625,N_23609);
nand U24494 (N_24494,N_23666,N_23894);
nand U24495 (N_24495,N_23509,N_23901);
and U24496 (N_24496,N_23990,N_23844);
or U24497 (N_24497,N_23689,N_23596);
or U24498 (N_24498,N_23847,N_23799);
or U24499 (N_24499,N_23648,N_23551);
nor U24500 (N_24500,N_24072,N_24463);
nand U24501 (N_24501,N_24049,N_24414);
nor U24502 (N_24502,N_24351,N_24079);
xnor U24503 (N_24503,N_24139,N_24194);
or U24504 (N_24504,N_24377,N_24460);
or U24505 (N_24505,N_24179,N_24020);
xnor U24506 (N_24506,N_24435,N_24078);
nor U24507 (N_24507,N_24278,N_24158);
xor U24508 (N_24508,N_24333,N_24131);
nand U24509 (N_24509,N_24420,N_24439);
and U24510 (N_24510,N_24417,N_24015);
or U24511 (N_24511,N_24418,N_24412);
xnor U24512 (N_24512,N_24248,N_24014);
nand U24513 (N_24513,N_24497,N_24487);
nand U24514 (N_24514,N_24474,N_24483);
xnor U24515 (N_24515,N_24432,N_24383);
or U24516 (N_24516,N_24394,N_24130);
nand U24517 (N_24517,N_24403,N_24301);
nor U24518 (N_24518,N_24096,N_24082);
or U24519 (N_24519,N_24000,N_24461);
xnor U24520 (N_24520,N_24124,N_24093);
and U24521 (N_24521,N_24498,N_24028);
and U24522 (N_24522,N_24293,N_24166);
nor U24523 (N_24523,N_24043,N_24246);
and U24524 (N_24524,N_24327,N_24175);
nor U24525 (N_24525,N_24284,N_24368);
nor U24526 (N_24526,N_24198,N_24308);
and U24527 (N_24527,N_24407,N_24355);
xnor U24528 (N_24528,N_24336,N_24121);
or U24529 (N_24529,N_24322,N_24290);
and U24530 (N_24530,N_24408,N_24136);
nor U24531 (N_24531,N_24359,N_24360);
nor U24532 (N_24532,N_24405,N_24018);
nand U24533 (N_24533,N_24100,N_24098);
xor U24534 (N_24534,N_24392,N_24171);
or U24535 (N_24535,N_24332,N_24236);
nand U24536 (N_24536,N_24346,N_24490);
nor U24537 (N_24537,N_24245,N_24052);
nor U24538 (N_24538,N_24253,N_24307);
xor U24539 (N_24539,N_24187,N_24061);
nand U24540 (N_24540,N_24310,N_24339);
or U24541 (N_24541,N_24492,N_24457);
nor U24542 (N_24542,N_24302,N_24433);
nor U24543 (N_24543,N_24311,N_24444);
nand U24544 (N_24544,N_24160,N_24410);
nor U24545 (N_24545,N_24397,N_24094);
and U24546 (N_24546,N_24331,N_24443);
nand U24547 (N_24547,N_24060,N_24334);
or U24548 (N_24548,N_24050,N_24450);
nor U24549 (N_24549,N_24451,N_24319);
nand U24550 (N_24550,N_24045,N_24476);
xnor U24551 (N_24551,N_24010,N_24204);
nor U24552 (N_24552,N_24207,N_24036);
nor U24553 (N_24553,N_24001,N_24055);
or U24554 (N_24554,N_24480,N_24004);
nand U24555 (N_24555,N_24174,N_24201);
xnor U24556 (N_24556,N_24012,N_24257);
and U24557 (N_24557,N_24149,N_24065);
nand U24558 (N_24558,N_24240,N_24344);
xnor U24559 (N_24559,N_24230,N_24064);
and U24560 (N_24560,N_24318,N_24205);
nand U24561 (N_24561,N_24372,N_24070);
xnor U24562 (N_24562,N_24384,N_24350);
or U24563 (N_24563,N_24140,N_24277);
and U24564 (N_24564,N_24153,N_24002);
and U24565 (N_24565,N_24467,N_24164);
nor U24566 (N_24566,N_24315,N_24430);
and U24567 (N_24567,N_24196,N_24127);
or U24568 (N_24568,N_24202,N_24109);
nor U24569 (N_24569,N_24465,N_24197);
nor U24570 (N_24570,N_24438,N_24495);
xor U24571 (N_24571,N_24494,N_24025);
nand U24572 (N_24572,N_24155,N_24269);
xor U24573 (N_24573,N_24266,N_24343);
or U24574 (N_24574,N_24297,N_24191);
nor U24575 (N_24575,N_24390,N_24272);
nand U24576 (N_24576,N_24401,N_24382);
nand U24577 (N_24577,N_24395,N_24080);
or U24578 (N_24578,N_24108,N_24141);
or U24579 (N_24579,N_24271,N_24056);
nand U24580 (N_24580,N_24200,N_24068);
or U24581 (N_24581,N_24275,N_24157);
and U24582 (N_24582,N_24227,N_24054);
or U24583 (N_24583,N_24466,N_24499);
or U24584 (N_24584,N_24447,N_24422);
or U24585 (N_24585,N_24254,N_24427);
and U24586 (N_24586,N_24256,N_24274);
and U24587 (N_24587,N_24220,N_24459);
and U24588 (N_24588,N_24326,N_24073);
nor U24589 (N_24589,N_24102,N_24416);
nand U24590 (N_24590,N_24247,N_24135);
or U24591 (N_24591,N_24446,N_24469);
nor U24592 (N_24592,N_24085,N_24345);
and U24593 (N_24593,N_24388,N_24371);
or U24594 (N_24594,N_24437,N_24151);
xor U24595 (N_24595,N_24250,N_24262);
or U24596 (N_24596,N_24128,N_24314);
and U24597 (N_24597,N_24285,N_24445);
and U24598 (N_24598,N_24379,N_24429);
nor U24599 (N_24599,N_24142,N_24152);
nor U24600 (N_24600,N_24040,N_24137);
xor U24601 (N_24601,N_24188,N_24145);
or U24602 (N_24602,N_24431,N_24007);
and U24603 (N_24603,N_24481,N_24243);
nor U24604 (N_24604,N_24421,N_24234);
or U24605 (N_24605,N_24129,N_24478);
xnor U24606 (N_24606,N_24287,N_24477);
or U24607 (N_24607,N_24364,N_24428);
nor U24608 (N_24608,N_24365,N_24434);
xnor U24609 (N_24609,N_24242,N_24156);
xnor U24610 (N_24610,N_24270,N_24110);
or U24611 (N_24611,N_24300,N_24017);
and U24612 (N_24612,N_24252,N_24066);
or U24613 (N_24613,N_24386,N_24338);
xnor U24614 (N_24614,N_24340,N_24177);
and U24615 (N_24615,N_24126,N_24409);
and U24616 (N_24616,N_24472,N_24186);
and U24617 (N_24617,N_24212,N_24095);
and U24618 (N_24618,N_24154,N_24406);
xor U24619 (N_24619,N_24321,N_24159);
xor U24620 (N_24620,N_24423,N_24111);
xor U24621 (N_24621,N_24105,N_24122);
or U24622 (N_24622,N_24024,N_24357);
nor U24623 (N_24623,N_24404,N_24218);
xnor U24624 (N_24624,N_24237,N_24486);
or U24625 (N_24625,N_24295,N_24051);
or U24626 (N_24626,N_24172,N_24226);
or U24627 (N_24627,N_24133,N_24279);
nand U24628 (N_24628,N_24458,N_24120);
nand U24629 (N_24629,N_24288,N_24150);
nor U24630 (N_24630,N_24009,N_24273);
or U24631 (N_24631,N_24325,N_24146);
or U24632 (N_24632,N_24342,N_24268);
xor U24633 (N_24633,N_24162,N_24281);
nor U24634 (N_24634,N_24053,N_24489);
and U24635 (N_24635,N_24209,N_24354);
nor U24636 (N_24636,N_24454,N_24267);
xor U24637 (N_24637,N_24448,N_24473);
nand U24638 (N_24638,N_24213,N_24464);
or U24639 (N_24639,N_24228,N_24440);
or U24640 (N_24640,N_24086,N_24038);
or U24641 (N_24641,N_24391,N_24083);
or U24642 (N_24642,N_24488,N_24258);
and U24643 (N_24643,N_24195,N_24022);
and U24644 (N_24644,N_24192,N_24398);
xnor U24645 (N_24645,N_24385,N_24496);
or U24646 (N_24646,N_24077,N_24358);
nor U24647 (N_24647,N_24033,N_24415);
or U24648 (N_24648,N_24493,N_24181);
or U24649 (N_24649,N_24452,N_24099);
nand U24650 (N_24650,N_24259,N_24317);
xnor U24651 (N_24651,N_24104,N_24027);
and U24652 (N_24652,N_24482,N_24441);
or U24653 (N_24653,N_24306,N_24475);
nand U24654 (N_24654,N_24165,N_24147);
nor U24655 (N_24655,N_24449,N_24217);
nor U24656 (N_24656,N_24214,N_24182);
or U24657 (N_24657,N_24030,N_24167);
nand U24658 (N_24658,N_24037,N_24117);
nor U24659 (N_24659,N_24400,N_24341);
nor U24660 (N_24660,N_24393,N_24369);
xor U24661 (N_24661,N_24471,N_24411);
xor U24662 (N_24662,N_24330,N_24442);
nand U24663 (N_24663,N_24426,N_24378);
nand U24664 (N_24664,N_24251,N_24413);
xnor U24665 (N_24665,N_24006,N_24348);
and U24666 (N_24666,N_24041,N_24313);
or U24667 (N_24667,N_24233,N_24203);
xnor U24668 (N_24668,N_24185,N_24180);
nand U24669 (N_24669,N_24143,N_24235);
xnor U24670 (N_24670,N_24046,N_24003);
nand U24671 (N_24671,N_24436,N_24032);
nand U24672 (N_24672,N_24402,N_24106);
xor U24673 (N_24673,N_24485,N_24299);
xnor U24674 (N_24674,N_24380,N_24320);
nand U24675 (N_24675,N_24184,N_24294);
nor U24676 (N_24676,N_24462,N_24329);
nor U24677 (N_24677,N_24224,N_24208);
or U24678 (N_24678,N_24044,N_24238);
and U24679 (N_24679,N_24169,N_24309);
nor U24680 (N_24680,N_24366,N_24016);
or U24681 (N_24681,N_24249,N_24352);
nor U24682 (N_24682,N_24005,N_24215);
nor U24683 (N_24683,N_24168,N_24261);
xnor U24684 (N_24684,N_24035,N_24076);
nor U24685 (N_24685,N_24363,N_24374);
or U24686 (N_24686,N_24479,N_24019);
or U24687 (N_24687,N_24264,N_24190);
nand U24688 (N_24688,N_24029,N_24138);
and U24689 (N_24689,N_24026,N_24023);
or U24690 (N_24690,N_24123,N_24069);
and U24691 (N_24691,N_24260,N_24335);
nor U24692 (N_24692,N_24081,N_24101);
xnor U24693 (N_24693,N_24225,N_24087);
nor U24694 (N_24694,N_24148,N_24088);
and U24695 (N_24695,N_24296,N_24067);
nand U24696 (N_24696,N_24232,N_24362);
xor U24697 (N_24697,N_24206,N_24376);
nor U24698 (N_24698,N_24013,N_24211);
xnor U24699 (N_24699,N_24375,N_24134);
or U24700 (N_24700,N_24298,N_24176);
nor U24701 (N_24701,N_24021,N_24303);
xnor U24702 (N_24702,N_24103,N_24161);
nand U24703 (N_24703,N_24039,N_24324);
nor U24704 (N_24704,N_24216,N_24241);
nor U24705 (N_24705,N_24107,N_24484);
and U24706 (N_24706,N_24048,N_24042);
xor U24707 (N_24707,N_24316,N_24470);
xor U24708 (N_24708,N_24280,N_24491);
xor U24709 (N_24709,N_24170,N_24084);
nand U24710 (N_24710,N_24089,N_24199);
xor U24711 (N_24711,N_24456,N_24381);
nand U24712 (N_24712,N_24074,N_24373);
nor U24713 (N_24713,N_24163,N_24276);
or U24714 (N_24714,N_24291,N_24387);
and U24715 (N_24715,N_24370,N_24091);
nor U24716 (N_24716,N_24057,N_24292);
nor U24717 (N_24717,N_24283,N_24144);
xor U24718 (N_24718,N_24210,N_24305);
nor U24719 (N_24719,N_24071,N_24356);
and U24720 (N_24720,N_24125,N_24113);
xor U24721 (N_24721,N_24058,N_24047);
xnor U24722 (N_24722,N_24114,N_24062);
or U24723 (N_24723,N_24323,N_24222);
and U24724 (N_24724,N_24034,N_24116);
or U24725 (N_24725,N_24178,N_24353);
and U24726 (N_24726,N_24223,N_24229);
and U24727 (N_24727,N_24092,N_24173);
nand U24728 (N_24728,N_24367,N_24221);
nor U24729 (N_24729,N_24265,N_24008);
xor U24730 (N_24730,N_24361,N_24063);
xor U24731 (N_24731,N_24419,N_24347);
and U24732 (N_24732,N_24011,N_24263);
and U24733 (N_24733,N_24219,N_24090);
xnor U24734 (N_24734,N_24118,N_24031);
and U24735 (N_24735,N_24468,N_24425);
xor U24736 (N_24736,N_24289,N_24244);
or U24737 (N_24737,N_24112,N_24183);
and U24738 (N_24738,N_24286,N_24193);
and U24739 (N_24739,N_24115,N_24255);
nand U24740 (N_24740,N_24075,N_24328);
and U24741 (N_24741,N_24304,N_24231);
xor U24742 (N_24742,N_24453,N_24337);
and U24743 (N_24743,N_24424,N_24455);
and U24744 (N_24744,N_24312,N_24389);
or U24745 (N_24745,N_24282,N_24097);
xnor U24746 (N_24746,N_24239,N_24396);
nor U24747 (N_24747,N_24119,N_24132);
xor U24748 (N_24748,N_24349,N_24189);
or U24749 (N_24749,N_24059,N_24399);
nor U24750 (N_24750,N_24177,N_24136);
nand U24751 (N_24751,N_24407,N_24475);
or U24752 (N_24752,N_24338,N_24221);
or U24753 (N_24753,N_24224,N_24018);
xor U24754 (N_24754,N_24065,N_24200);
xnor U24755 (N_24755,N_24219,N_24451);
nand U24756 (N_24756,N_24198,N_24116);
xnor U24757 (N_24757,N_24031,N_24089);
xnor U24758 (N_24758,N_24371,N_24304);
nor U24759 (N_24759,N_24284,N_24347);
nor U24760 (N_24760,N_24063,N_24053);
and U24761 (N_24761,N_24300,N_24262);
or U24762 (N_24762,N_24080,N_24201);
or U24763 (N_24763,N_24240,N_24066);
and U24764 (N_24764,N_24439,N_24402);
and U24765 (N_24765,N_24195,N_24339);
or U24766 (N_24766,N_24236,N_24333);
xnor U24767 (N_24767,N_24051,N_24005);
nand U24768 (N_24768,N_24326,N_24353);
xor U24769 (N_24769,N_24219,N_24313);
xnor U24770 (N_24770,N_24263,N_24369);
nand U24771 (N_24771,N_24236,N_24213);
and U24772 (N_24772,N_24472,N_24382);
or U24773 (N_24773,N_24026,N_24140);
xnor U24774 (N_24774,N_24310,N_24379);
nand U24775 (N_24775,N_24055,N_24464);
xor U24776 (N_24776,N_24293,N_24236);
and U24777 (N_24777,N_24381,N_24072);
xor U24778 (N_24778,N_24449,N_24209);
or U24779 (N_24779,N_24404,N_24018);
nand U24780 (N_24780,N_24414,N_24383);
nor U24781 (N_24781,N_24040,N_24060);
nand U24782 (N_24782,N_24087,N_24164);
xnor U24783 (N_24783,N_24013,N_24303);
xor U24784 (N_24784,N_24134,N_24212);
xnor U24785 (N_24785,N_24191,N_24256);
and U24786 (N_24786,N_24382,N_24351);
xor U24787 (N_24787,N_24403,N_24420);
nand U24788 (N_24788,N_24077,N_24009);
or U24789 (N_24789,N_24063,N_24061);
and U24790 (N_24790,N_24462,N_24471);
or U24791 (N_24791,N_24424,N_24030);
xnor U24792 (N_24792,N_24172,N_24298);
or U24793 (N_24793,N_24370,N_24224);
nand U24794 (N_24794,N_24451,N_24081);
and U24795 (N_24795,N_24446,N_24411);
xor U24796 (N_24796,N_24086,N_24462);
xor U24797 (N_24797,N_24412,N_24241);
xnor U24798 (N_24798,N_24009,N_24005);
nand U24799 (N_24799,N_24123,N_24015);
or U24800 (N_24800,N_24270,N_24155);
or U24801 (N_24801,N_24496,N_24052);
and U24802 (N_24802,N_24055,N_24150);
xor U24803 (N_24803,N_24455,N_24287);
nor U24804 (N_24804,N_24016,N_24047);
xor U24805 (N_24805,N_24234,N_24208);
and U24806 (N_24806,N_24314,N_24494);
and U24807 (N_24807,N_24115,N_24352);
nor U24808 (N_24808,N_24477,N_24359);
and U24809 (N_24809,N_24294,N_24085);
and U24810 (N_24810,N_24464,N_24141);
xnor U24811 (N_24811,N_24206,N_24378);
and U24812 (N_24812,N_24288,N_24052);
or U24813 (N_24813,N_24055,N_24019);
and U24814 (N_24814,N_24153,N_24330);
nand U24815 (N_24815,N_24396,N_24074);
and U24816 (N_24816,N_24310,N_24153);
xor U24817 (N_24817,N_24070,N_24043);
and U24818 (N_24818,N_24110,N_24100);
nor U24819 (N_24819,N_24049,N_24100);
xor U24820 (N_24820,N_24254,N_24326);
xor U24821 (N_24821,N_24124,N_24003);
and U24822 (N_24822,N_24475,N_24404);
or U24823 (N_24823,N_24068,N_24180);
and U24824 (N_24824,N_24089,N_24069);
nand U24825 (N_24825,N_24357,N_24281);
and U24826 (N_24826,N_24196,N_24404);
and U24827 (N_24827,N_24354,N_24147);
nand U24828 (N_24828,N_24151,N_24470);
nor U24829 (N_24829,N_24235,N_24037);
nor U24830 (N_24830,N_24257,N_24135);
or U24831 (N_24831,N_24128,N_24470);
nand U24832 (N_24832,N_24303,N_24380);
xnor U24833 (N_24833,N_24167,N_24332);
nor U24834 (N_24834,N_24432,N_24227);
nor U24835 (N_24835,N_24071,N_24242);
or U24836 (N_24836,N_24195,N_24018);
xor U24837 (N_24837,N_24297,N_24295);
nand U24838 (N_24838,N_24418,N_24196);
nand U24839 (N_24839,N_24326,N_24485);
nor U24840 (N_24840,N_24068,N_24306);
and U24841 (N_24841,N_24078,N_24309);
xor U24842 (N_24842,N_24256,N_24025);
xor U24843 (N_24843,N_24461,N_24438);
xor U24844 (N_24844,N_24319,N_24078);
nand U24845 (N_24845,N_24106,N_24343);
and U24846 (N_24846,N_24459,N_24128);
nor U24847 (N_24847,N_24430,N_24353);
or U24848 (N_24848,N_24231,N_24068);
and U24849 (N_24849,N_24497,N_24237);
or U24850 (N_24850,N_24462,N_24483);
nand U24851 (N_24851,N_24262,N_24269);
nand U24852 (N_24852,N_24132,N_24479);
xor U24853 (N_24853,N_24187,N_24422);
nand U24854 (N_24854,N_24186,N_24121);
and U24855 (N_24855,N_24408,N_24122);
and U24856 (N_24856,N_24061,N_24431);
or U24857 (N_24857,N_24299,N_24076);
nor U24858 (N_24858,N_24050,N_24192);
nor U24859 (N_24859,N_24040,N_24329);
nor U24860 (N_24860,N_24386,N_24053);
nor U24861 (N_24861,N_24268,N_24332);
nand U24862 (N_24862,N_24031,N_24104);
or U24863 (N_24863,N_24292,N_24173);
nor U24864 (N_24864,N_24091,N_24068);
xor U24865 (N_24865,N_24410,N_24322);
nor U24866 (N_24866,N_24110,N_24304);
and U24867 (N_24867,N_24074,N_24427);
nand U24868 (N_24868,N_24178,N_24186);
nor U24869 (N_24869,N_24415,N_24431);
nand U24870 (N_24870,N_24121,N_24041);
xnor U24871 (N_24871,N_24209,N_24466);
or U24872 (N_24872,N_24153,N_24151);
nor U24873 (N_24873,N_24167,N_24161);
xor U24874 (N_24874,N_24485,N_24161);
nor U24875 (N_24875,N_24279,N_24268);
xor U24876 (N_24876,N_24480,N_24140);
nand U24877 (N_24877,N_24397,N_24387);
xnor U24878 (N_24878,N_24007,N_24028);
xnor U24879 (N_24879,N_24105,N_24414);
or U24880 (N_24880,N_24339,N_24009);
nor U24881 (N_24881,N_24207,N_24026);
and U24882 (N_24882,N_24316,N_24100);
nand U24883 (N_24883,N_24377,N_24254);
xnor U24884 (N_24884,N_24273,N_24350);
or U24885 (N_24885,N_24004,N_24362);
xor U24886 (N_24886,N_24288,N_24015);
xor U24887 (N_24887,N_24449,N_24359);
and U24888 (N_24888,N_24217,N_24255);
nor U24889 (N_24889,N_24497,N_24470);
or U24890 (N_24890,N_24225,N_24146);
nand U24891 (N_24891,N_24191,N_24022);
nand U24892 (N_24892,N_24144,N_24042);
nand U24893 (N_24893,N_24123,N_24447);
xor U24894 (N_24894,N_24194,N_24307);
and U24895 (N_24895,N_24277,N_24278);
xnor U24896 (N_24896,N_24397,N_24251);
nor U24897 (N_24897,N_24327,N_24370);
nor U24898 (N_24898,N_24484,N_24011);
xnor U24899 (N_24899,N_24272,N_24471);
nand U24900 (N_24900,N_24133,N_24219);
xnor U24901 (N_24901,N_24466,N_24372);
or U24902 (N_24902,N_24253,N_24471);
nor U24903 (N_24903,N_24316,N_24302);
nand U24904 (N_24904,N_24105,N_24220);
or U24905 (N_24905,N_24111,N_24305);
and U24906 (N_24906,N_24293,N_24123);
or U24907 (N_24907,N_24064,N_24182);
or U24908 (N_24908,N_24435,N_24219);
or U24909 (N_24909,N_24062,N_24255);
xnor U24910 (N_24910,N_24054,N_24044);
and U24911 (N_24911,N_24210,N_24102);
nor U24912 (N_24912,N_24325,N_24009);
nand U24913 (N_24913,N_24210,N_24010);
nand U24914 (N_24914,N_24190,N_24235);
xor U24915 (N_24915,N_24402,N_24320);
xnor U24916 (N_24916,N_24169,N_24471);
and U24917 (N_24917,N_24485,N_24061);
xnor U24918 (N_24918,N_24207,N_24315);
xor U24919 (N_24919,N_24074,N_24459);
and U24920 (N_24920,N_24350,N_24168);
nor U24921 (N_24921,N_24462,N_24475);
xnor U24922 (N_24922,N_24002,N_24346);
nor U24923 (N_24923,N_24156,N_24073);
and U24924 (N_24924,N_24364,N_24072);
and U24925 (N_24925,N_24108,N_24164);
and U24926 (N_24926,N_24044,N_24030);
and U24927 (N_24927,N_24458,N_24125);
xor U24928 (N_24928,N_24494,N_24208);
nor U24929 (N_24929,N_24190,N_24387);
nand U24930 (N_24930,N_24461,N_24166);
xnor U24931 (N_24931,N_24010,N_24482);
nand U24932 (N_24932,N_24012,N_24431);
and U24933 (N_24933,N_24364,N_24006);
xor U24934 (N_24934,N_24061,N_24181);
nand U24935 (N_24935,N_24398,N_24147);
nand U24936 (N_24936,N_24187,N_24498);
xnor U24937 (N_24937,N_24346,N_24405);
or U24938 (N_24938,N_24188,N_24091);
or U24939 (N_24939,N_24226,N_24115);
and U24940 (N_24940,N_24411,N_24190);
nand U24941 (N_24941,N_24161,N_24296);
or U24942 (N_24942,N_24114,N_24274);
or U24943 (N_24943,N_24077,N_24151);
nor U24944 (N_24944,N_24205,N_24002);
nor U24945 (N_24945,N_24414,N_24204);
nor U24946 (N_24946,N_24220,N_24479);
nand U24947 (N_24947,N_24378,N_24078);
xnor U24948 (N_24948,N_24119,N_24056);
or U24949 (N_24949,N_24243,N_24039);
and U24950 (N_24950,N_24132,N_24415);
nand U24951 (N_24951,N_24371,N_24107);
nand U24952 (N_24952,N_24440,N_24402);
xnor U24953 (N_24953,N_24066,N_24235);
and U24954 (N_24954,N_24087,N_24167);
and U24955 (N_24955,N_24406,N_24448);
nor U24956 (N_24956,N_24347,N_24110);
or U24957 (N_24957,N_24029,N_24404);
nor U24958 (N_24958,N_24377,N_24341);
or U24959 (N_24959,N_24073,N_24008);
nor U24960 (N_24960,N_24394,N_24189);
xnor U24961 (N_24961,N_24334,N_24039);
nor U24962 (N_24962,N_24334,N_24433);
or U24963 (N_24963,N_24498,N_24070);
nor U24964 (N_24964,N_24186,N_24034);
xnor U24965 (N_24965,N_24403,N_24303);
nand U24966 (N_24966,N_24300,N_24487);
xnor U24967 (N_24967,N_24301,N_24380);
or U24968 (N_24968,N_24066,N_24041);
nor U24969 (N_24969,N_24386,N_24020);
nand U24970 (N_24970,N_24464,N_24341);
and U24971 (N_24971,N_24482,N_24300);
or U24972 (N_24972,N_24288,N_24007);
or U24973 (N_24973,N_24092,N_24095);
nor U24974 (N_24974,N_24272,N_24377);
nor U24975 (N_24975,N_24078,N_24060);
or U24976 (N_24976,N_24296,N_24241);
or U24977 (N_24977,N_24162,N_24158);
or U24978 (N_24978,N_24026,N_24200);
or U24979 (N_24979,N_24037,N_24209);
or U24980 (N_24980,N_24207,N_24111);
and U24981 (N_24981,N_24080,N_24413);
or U24982 (N_24982,N_24156,N_24490);
nand U24983 (N_24983,N_24075,N_24476);
and U24984 (N_24984,N_24446,N_24431);
nand U24985 (N_24985,N_24270,N_24096);
xnor U24986 (N_24986,N_24187,N_24497);
xor U24987 (N_24987,N_24066,N_24030);
or U24988 (N_24988,N_24333,N_24136);
and U24989 (N_24989,N_24452,N_24291);
or U24990 (N_24990,N_24147,N_24050);
or U24991 (N_24991,N_24182,N_24013);
nand U24992 (N_24992,N_24136,N_24147);
xor U24993 (N_24993,N_24057,N_24060);
nand U24994 (N_24994,N_24192,N_24405);
xor U24995 (N_24995,N_24020,N_24166);
nand U24996 (N_24996,N_24300,N_24489);
nor U24997 (N_24997,N_24482,N_24097);
nand U24998 (N_24998,N_24437,N_24482);
nor U24999 (N_24999,N_24371,N_24102);
nand U25000 (N_25000,N_24812,N_24641);
nor U25001 (N_25001,N_24598,N_24683);
nor U25002 (N_25002,N_24860,N_24829);
nand U25003 (N_25003,N_24875,N_24822);
and U25004 (N_25004,N_24501,N_24697);
nand U25005 (N_25005,N_24536,N_24743);
and U25006 (N_25006,N_24887,N_24821);
nor U25007 (N_25007,N_24966,N_24892);
and U25008 (N_25008,N_24916,N_24525);
xnor U25009 (N_25009,N_24927,N_24959);
and U25010 (N_25010,N_24638,N_24781);
and U25011 (N_25011,N_24589,N_24500);
xnor U25012 (N_25012,N_24775,N_24531);
or U25013 (N_25013,N_24745,N_24649);
or U25014 (N_25014,N_24643,N_24569);
nor U25015 (N_25015,N_24783,N_24958);
nor U25016 (N_25016,N_24604,N_24869);
nor U25017 (N_25017,N_24599,N_24619);
or U25018 (N_25018,N_24856,N_24996);
or U25019 (N_25019,N_24815,N_24660);
xor U25020 (N_25020,N_24735,N_24900);
and U25021 (N_25021,N_24736,N_24684);
and U25022 (N_25022,N_24512,N_24615);
nand U25023 (N_25023,N_24765,N_24950);
and U25024 (N_25024,N_24894,N_24767);
xor U25025 (N_25025,N_24956,N_24579);
nand U25026 (N_25026,N_24814,N_24907);
nor U25027 (N_25027,N_24594,N_24968);
and U25028 (N_25028,N_24626,N_24942);
nand U25029 (N_25029,N_24929,N_24678);
or U25030 (N_25030,N_24964,N_24548);
xor U25031 (N_25031,N_24769,N_24510);
and U25032 (N_25032,N_24945,N_24778);
and U25033 (N_25033,N_24762,N_24692);
nand U25034 (N_25034,N_24562,N_24857);
or U25035 (N_25035,N_24858,N_24596);
or U25036 (N_25036,N_24534,N_24515);
or U25037 (N_25037,N_24664,N_24581);
nand U25038 (N_25038,N_24859,N_24748);
or U25039 (N_25039,N_24839,N_24811);
or U25040 (N_25040,N_24987,N_24928);
nor U25041 (N_25041,N_24819,N_24528);
and U25042 (N_25042,N_24570,N_24939);
nor U25043 (N_25043,N_24618,N_24696);
nor U25044 (N_25044,N_24808,N_24623);
nor U25045 (N_25045,N_24560,N_24522);
and U25046 (N_25046,N_24742,N_24687);
nor U25047 (N_25047,N_24930,N_24764);
xor U25048 (N_25048,N_24637,N_24844);
nand U25049 (N_25049,N_24868,N_24592);
nand U25050 (N_25050,N_24771,N_24688);
or U25051 (N_25051,N_24917,N_24634);
nand U25052 (N_25052,N_24941,N_24518);
xor U25053 (N_25053,N_24524,N_24753);
nor U25054 (N_25054,N_24972,N_24609);
and U25055 (N_25055,N_24636,N_24555);
or U25056 (N_25056,N_24951,N_24792);
or U25057 (N_25057,N_24997,N_24572);
or U25058 (N_25058,N_24804,N_24985);
or U25059 (N_25059,N_24582,N_24905);
or U25060 (N_25060,N_24866,N_24788);
nand U25061 (N_25061,N_24969,N_24595);
xnor U25062 (N_25062,N_24602,N_24651);
xnor U25063 (N_25063,N_24610,N_24622);
xor U25064 (N_25064,N_24706,N_24890);
xor U25065 (N_25065,N_24909,N_24756);
nor U25066 (N_25066,N_24681,N_24874);
nor U25067 (N_25067,N_24818,N_24865);
nand U25068 (N_25068,N_24708,N_24529);
nor U25069 (N_25069,N_24768,N_24564);
nand U25070 (N_25070,N_24850,N_24910);
or U25071 (N_25071,N_24834,N_24639);
xnor U25072 (N_25072,N_24655,N_24558);
and U25073 (N_25073,N_24652,N_24733);
nand U25074 (N_25074,N_24543,N_24675);
nor U25075 (N_25075,N_24521,N_24547);
xnor U25076 (N_25076,N_24978,N_24566);
nor U25077 (N_25077,N_24898,N_24502);
and U25078 (N_25078,N_24971,N_24871);
xnor U25079 (N_25079,N_24787,N_24730);
xnor U25080 (N_25080,N_24666,N_24741);
and U25081 (N_25081,N_24617,N_24902);
and U25082 (N_25082,N_24995,N_24896);
and U25083 (N_25083,N_24705,N_24879);
or U25084 (N_25084,N_24731,N_24703);
or U25085 (N_25085,N_24751,N_24809);
or U25086 (N_25086,N_24982,N_24785);
xnor U25087 (N_25087,N_24813,N_24593);
and U25088 (N_25088,N_24573,N_24800);
and U25089 (N_25089,N_24870,N_24925);
or U25090 (N_25090,N_24944,N_24663);
or U25091 (N_25091,N_24554,N_24761);
xnor U25092 (N_25092,N_24852,N_24728);
and U25093 (N_25093,N_24517,N_24758);
xor U25094 (N_25094,N_24551,N_24539);
nor U25095 (N_25095,N_24933,N_24556);
xnor U25096 (N_25096,N_24993,N_24565);
nand U25097 (N_25097,N_24689,N_24999);
or U25098 (N_25098,N_24961,N_24931);
nand U25099 (N_25099,N_24983,N_24732);
or U25100 (N_25100,N_24750,N_24509);
xnor U25101 (N_25101,N_24754,N_24801);
or U25102 (N_25102,N_24632,N_24782);
or U25103 (N_25103,N_24737,N_24840);
and U25104 (N_25104,N_24977,N_24780);
xnor U25105 (N_25105,N_24938,N_24571);
nand U25106 (N_25106,N_24913,N_24523);
and U25107 (N_25107,N_24826,N_24552);
and U25108 (N_25108,N_24845,N_24906);
and U25109 (N_25109,N_24885,N_24881);
and U25110 (N_25110,N_24716,N_24876);
nor U25111 (N_25111,N_24511,N_24612);
or U25112 (N_25112,N_24645,N_24616);
or U25113 (N_25113,N_24714,N_24717);
and U25114 (N_25114,N_24676,N_24825);
nand U25115 (N_25115,N_24590,N_24605);
or U25116 (N_25116,N_24685,N_24691);
xnor U25117 (N_25117,N_24624,N_24702);
nor U25118 (N_25118,N_24585,N_24766);
and U25119 (N_25119,N_24770,N_24855);
or U25120 (N_25120,N_24802,N_24607);
nor U25121 (N_25121,N_24970,N_24994);
nor U25122 (N_25122,N_24646,N_24658);
nor U25123 (N_25123,N_24583,N_24704);
xnor U25124 (N_25124,N_24591,N_24823);
and U25125 (N_25125,N_24668,N_24790);
nand U25126 (N_25126,N_24799,N_24990);
and U25127 (N_25127,N_24654,N_24673);
and U25128 (N_25128,N_24810,N_24575);
or U25129 (N_25129,N_24786,N_24606);
or U25130 (N_25130,N_24656,N_24901);
nor U25131 (N_25131,N_24965,N_24806);
and U25132 (N_25132,N_24798,N_24672);
nor U25133 (N_25133,N_24949,N_24984);
nand U25134 (N_25134,N_24757,N_24979);
xor U25135 (N_25135,N_24973,N_24976);
and U25136 (N_25136,N_24659,N_24710);
nand U25137 (N_25137,N_24904,N_24937);
xnor U25138 (N_25138,N_24698,N_24580);
nor U25139 (N_25139,N_24967,N_24888);
nor U25140 (N_25140,N_24739,N_24635);
nand U25141 (N_25141,N_24914,N_24613);
xnor U25142 (N_25142,N_24740,N_24724);
or U25143 (N_25143,N_24648,N_24520);
nand U25144 (N_25144,N_24797,N_24722);
or U25145 (N_25145,N_24989,N_24838);
nand U25146 (N_25146,N_24789,N_24526);
nor U25147 (N_25147,N_24516,N_24549);
nand U25148 (N_25148,N_24709,N_24541);
nor U25149 (N_25149,N_24600,N_24746);
and U25150 (N_25150,N_24694,N_24577);
or U25151 (N_25151,N_24827,N_24795);
and U25152 (N_25152,N_24794,N_24807);
and U25153 (N_25153,N_24640,N_24992);
xnor U25154 (N_25154,N_24584,N_24707);
nor U25155 (N_25155,N_24729,N_24559);
nand U25156 (N_25156,N_24974,N_24621);
and U25157 (N_25157,N_24701,N_24832);
or U25158 (N_25158,N_24837,N_24550);
or U25159 (N_25159,N_24774,N_24922);
or U25160 (N_25160,N_24817,N_24715);
xnor U25161 (N_25161,N_24830,N_24537);
and U25162 (N_25162,N_24680,N_24920);
nor U25163 (N_25163,N_24535,N_24843);
and U25164 (N_25164,N_24503,N_24805);
nand U25165 (N_25165,N_24791,N_24986);
and U25166 (N_25166,N_24587,N_24773);
nor U25167 (N_25167,N_24532,N_24718);
nand U25168 (N_25168,N_24713,N_24744);
or U25169 (N_25169,N_24657,N_24760);
xnor U25170 (N_25170,N_24711,N_24644);
xor U25171 (N_25171,N_24877,N_24864);
nand U25172 (N_25172,N_24527,N_24953);
nand U25173 (N_25173,N_24538,N_24820);
or U25174 (N_25174,N_24936,N_24545);
and U25175 (N_25175,N_24533,N_24915);
nor U25176 (N_25176,N_24625,N_24608);
or U25177 (N_25177,N_24614,N_24514);
xnor U25178 (N_25178,N_24851,N_24847);
and U25179 (N_25179,N_24833,N_24508);
nor U25180 (N_25180,N_24763,N_24627);
and U25181 (N_25181,N_24667,N_24588);
nand U25182 (N_25182,N_24661,N_24828);
xnor U25183 (N_25183,N_24947,N_24563);
nand U25184 (N_25184,N_24557,N_24699);
or U25185 (N_25185,N_24862,N_24723);
nand U25186 (N_25186,N_24700,N_24803);
nor U25187 (N_25187,N_24934,N_24674);
or U25188 (N_25188,N_24923,N_24880);
nor U25189 (N_25189,N_24686,N_24854);
and U25190 (N_25190,N_24630,N_24752);
and U25191 (N_25191,N_24872,N_24882);
nand U25192 (N_25192,N_24749,N_24816);
nand U25193 (N_25193,N_24878,N_24578);
nand U25194 (N_25194,N_24561,N_24677);
nand U25195 (N_25195,N_24633,N_24662);
or U25196 (N_25196,N_24946,N_24886);
nand U25197 (N_25197,N_24988,N_24712);
xor U25198 (N_25198,N_24506,N_24670);
and U25199 (N_25199,N_24779,N_24665);
or U25200 (N_25200,N_24835,N_24542);
and U25201 (N_25201,N_24883,N_24597);
xnor U25202 (N_25202,N_24647,N_24908);
nor U25203 (N_25203,N_24981,N_24793);
xnor U25204 (N_25204,N_24586,N_24921);
nand U25205 (N_25205,N_24897,N_24975);
or U25206 (N_25206,N_24926,N_24553);
nor U25207 (N_25207,N_24867,N_24980);
or U25208 (N_25208,N_24544,N_24629);
nand U25209 (N_25209,N_24690,N_24954);
nand U25210 (N_25210,N_24738,N_24960);
nand U25211 (N_25211,N_24861,N_24924);
or U25212 (N_25212,N_24603,N_24891);
or U25213 (N_25213,N_24889,N_24650);
or U25214 (N_25214,N_24903,N_24601);
nor U25215 (N_25215,N_24940,N_24734);
or U25216 (N_25216,N_24873,N_24935);
nand U25217 (N_25217,N_24679,N_24695);
and U25218 (N_25218,N_24726,N_24759);
xnor U25219 (N_25219,N_24911,N_24620);
and U25220 (N_25220,N_24611,N_24568);
nand U25221 (N_25221,N_24507,N_24671);
nand U25222 (N_25222,N_24574,N_24963);
nor U25223 (N_25223,N_24631,N_24943);
or U25224 (N_25224,N_24895,N_24504);
and U25225 (N_25225,N_24899,N_24853);
nor U25226 (N_25226,N_24777,N_24719);
nor U25227 (N_25227,N_24540,N_24955);
nor U25228 (N_25228,N_24720,N_24932);
or U25229 (N_25229,N_24912,N_24628);
nor U25230 (N_25230,N_24884,N_24919);
and U25231 (N_25231,N_24519,N_24863);
nand U25232 (N_25232,N_24948,N_24842);
and U25233 (N_25233,N_24836,N_24776);
and U25234 (N_25234,N_24831,N_24505);
and U25235 (N_25235,N_24841,N_24772);
nor U25236 (N_25236,N_24784,N_24824);
nand U25237 (N_25237,N_24957,N_24669);
nand U25238 (N_25238,N_24796,N_24747);
xor U25239 (N_25239,N_24962,N_24530);
and U25240 (N_25240,N_24998,N_24721);
xor U25241 (N_25241,N_24513,N_24952);
xnor U25242 (N_25242,N_24693,N_24682);
nand U25243 (N_25243,N_24653,N_24918);
nor U25244 (N_25244,N_24755,N_24567);
nor U25245 (N_25245,N_24849,N_24848);
xor U25246 (N_25246,N_24893,N_24725);
nor U25247 (N_25247,N_24642,N_24846);
nor U25248 (N_25248,N_24727,N_24576);
nor U25249 (N_25249,N_24546,N_24991);
nor U25250 (N_25250,N_24829,N_24657);
or U25251 (N_25251,N_24719,N_24611);
nand U25252 (N_25252,N_24548,N_24937);
and U25253 (N_25253,N_24638,N_24872);
and U25254 (N_25254,N_24832,N_24613);
nor U25255 (N_25255,N_24641,N_24507);
or U25256 (N_25256,N_24594,N_24566);
and U25257 (N_25257,N_24816,N_24551);
nand U25258 (N_25258,N_24849,N_24993);
or U25259 (N_25259,N_24745,N_24603);
nor U25260 (N_25260,N_24738,N_24732);
or U25261 (N_25261,N_24774,N_24959);
nor U25262 (N_25262,N_24816,N_24612);
and U25263 (N_25263,N_24622,N_24765);
or U25264 (N_25264,N_24712,N_24520);
nand U25265 (N_25265,N_24712,N_24524);
xor U25266 (N_25266,N_24677,N_24753);
and U25267 (N_25267,N_24882,N_24630);
nor U25268 (N_25268,N_24731,N_24503);
xor U25269 (N_25269,N_24614,N_24763);
xor U25270 (N_25270,N_24847,N_24967);
nor U25271 (N_25271,N_24682,N_24916);
xnor U25272 (N_25272,N_24800,N_24878);
and U25273 (N_25273,N_24569,N_24707);
nand U25274 (N_25274,N_24981,N_24530);
or U25275 (N_25275,N_24971,N_24911);
nand U25276 (N_25276,N_24971,N_24524);
xnor U25277 (N_25277,N_24861,N_24671);
or U25278 (N_25278,N_24886,N_24987);
nand U25279 (N_25279,N_24683,N_24621);
nand U25280 (N_25280,N_24787,N_24968);
xor U25281 (N_25281,N_24838,N_24576);
xnor U25282 (N_25282,N_24522,N_24975);
and U25283 (N_25283,N_24561,N_24922);
and U25284 (N_25284,N_24584,N_24537);
nand U25285 (N_25285,N_24576,N_24530);
or U25286 (N_25286,N_24594,N_24698);
or U25287 (N_25287,N_24725,N_24898);
nor U25288 (N_25288,N_24818,N_24814);
nor U25289 (N_25289,N_24572,N_24594);
xor U25290 (N_25290,N_24663,N_24986);
nand U25291 (N_25291,N_24753,N_24532);
nand U25292 (N_25292,N_24767,N_24739);
xnor U25293 (N_25293,N_24784,N_24926);
and U25294 (N_25294,N_24879,N_24912);
or U25295 (N_25295,N_24511,N_24679);
or U25296 (N_25296,N_24955,N_24905);
nand U25297 (N_25297,N_24739,N_24869);
nor U25298 (N_25298,N_24986,N_24587);
or U25299 (N_25299,N_24524,N_24997);
nor U25300 (N_25300,N_24576,N_24941);
nand U25301 (N_25301,N_24639,N_24667);
xnor U25302 (N_25302,N_24547,N_24605);
or U25303 (N_25303,N_24681,N_24940);
and U25304 (N_25304,N_24844,N_24749);
xor U25305 (N_25305,N_24833,N_24884);
or U25306 (N_25306,N_24815,N_24650);
or U25307 (N_25307,N_24816,N_24779);
xor U25308 (N_25308,N_24689,N_24902);
or U25309 (N_25309,N_24987,N_24639);
and U25310 (N_25310,N_24541,N_24846);
nor U25311 (N_25311,N_24881,N_24737);
or U25312 (N_25312,N_24551,N_24906);
nor U25313 (N_25313,N_24574,N_24568);
nand U25314 (N_25314,N_24806,N_24837);
nor U25315 (N_25315,N_24769,N_24533);
nor U25316 (N_25316,N_24656,N_24841);
nor U25317 (N_25317,N_24720,N_24500);
nor U25318 (N_25318,N_24853,N_24964);
nand U25319 (N_25319,N_24878,N_24560);
nand U25320 (N_25320,N_24993,N_24620);
xor U25321 (N_25321,N_24673,N_24915);
xnor U25322 (N_25322,N_24685,N_24861);
and U25323 (N_25323,N_24957,N_24758);
nand U25324 (N_25324,N_24579,N_24797);
or U25325 (N_25325,N_24609,N_24952);
nand U25326 (N_25326,N_24688,N_24719);
nor U25327 (N_25327,N_24646,N_24576);
nor U25328 (N_25328,N_24579,N_24504);
and U25329 (N_25329,N_24800,N_24520);
nor U25330 (N_25330,N_24840,N_24825);
or U25331 (N_25331,N_24595,N_24684);
xor U25332 (N_25332,N_24783,N_24613);
or U25333 (N_25333,N_24801,N_24572);
nand U25334 (N_25334,N_24883,N_24592);
nand U25335 (N_25335,N_24679,N_24950);
and U25336 (N_25336,N_24714,N_24637);
xor U25337 (N_25337,N_24538,N_24877);
or U25338 (N_25338,N_24659,N_24768);
nand U25339 (N_25339,N_24950,N_24609);
xnor U25340 (N_25340,N_24989,N_24988);
nor U25341 (N_25341,N_24895,N_24869);
nand U25342 (N_25342,N_24544,N_24983);
xnor U25343 (N_25343,N_24852,N_24945);
nand U25344 (N_25344,N_24985,N_24590);
nor U25345 (N_25345,N_24596,N_24944);
and U25346 (N_25346,N_24928,N_24884);
or U25347 (N_25347,N_24508,N_24888);
nor U25348 (N_25348,N_24998,N_24629);
nor U25349 (N_25349,N_24966,N_24574);
or U25350 (N_25350,N_24965,N_24845);
xnor U25351 (N_25351,N_24797,N_24810);
xnor U25352 (N_25352,N_24599,N_24709);
nand U25353 (N_25353,N_24501,N_24559);
nand U25354 (N_25354,N_24725,N_24677);
or U25355 (N_25355,N_24950,N_24756);
nand U25356 (N_25356,N_24515,N_24875);
xor U25357 (N_25357,N_24535,N_24624);
xor U25358 (N_25358,N_24584,N_24950);
xor U25359 (N_25359,N_24731,N_24800);
xor U25360 (N_25360,N_24762,N_24825);
and U25361 (N_25361,N_24552,N_24777);
or U25362 (N_25362,N_24682,N_24906);
nand U25363 (N_25363,N_24550,N_24584);
xnor U25364 (N_25364,N_24642,N_24982);
or U25365 (N_25365,N_24997,N_24797);
xor U25366 (N_25366,N_24960,N_24668);
and U25367 (N_25367,N_24813,N_24917);
nor U25368 (N_25368,N_24717,N_24547);
nor U25369 (N_25369,N_24683,N_24876);
nand U25370 (N_25370,N_24576,N_24820);
or U25371 (N_25371,N_24841,N_24644);
and U25372 (N_25372,N_24738,N_24935);
nand U25373 (N_25373,N_24704,N_24501);
or U25374 (N_25374,N_24514,N_24697);
or U25375 (N_25375,N_24556,N_24970);
or U25376 (N_25376,N_24993,N_24554);
and U25377 (N_25377,N_24681,N_24933);
nor U25378 (N_25378,N_24888,N_24992);
or U25379 (N_25379,N_24757,N_24701);
nor U25380 (N_25380,N_24625,N_24996);
nand U25381 (N_25381,N_24513,N_24814);
and U25382 (N_25382,N_24552,N_24811);
and U25383 (N_25383,N_24704,N_24932);
and U25384 (N_25384,N_24745,N_24965);
or U25385 (N_25385,N_24811,N_24881);
xnor U25386 (N_25386,N_24525,N_24794);
xor U25387 (N_25387,N_24591,N_24624);
xor U25388 (N_25388,N_24919,N_24535);
xnor U25389 (N_25389,N_24793,N_24610);
xnor U25390 (N_25390,N_24698,N_24770);
xnor U25391 (N_25391,N_24666,N_24718);
and U25392 (N_25392,N_24513,N_24580);
or U25393 (N_25393,N_24668,N_24957);
or U25394 (N_25394,N_24602,N_24703);
nand U25395 (N_25395,N_24945,N_24953);
nand U25396 (N_25396,N_24566,N_24688);
xor U25397 (N_25397,N_24924,N_24853);
and U25398 (N_25398,N_24887,N_24591);
nor U25399 (N_25399,N_24682,N_24579);
nor U25400 (N_25400,N_24709,N_24863);
and U25401 (N_25401,N_24845,N_24759);
nand U25402 (N_25402,N_24757,N_24627);
nor U25403 (N_25403,N_24647,N_24926);
or U25404 (N_25404,N_24552,N_24619);
xor U25405 (N_25405,N_24579,N_24601);
or U25406 (N_25406,N_24680,N_24838);
and U25407 (N_25407,N_24712,N_24586);
or U25408 (N_25408,N_24901,N_24573);
and U25409 (N_25409,N_24551,N_24623);
xor U25410 (N_25410,N_24761,N_24863);
or U25411 (N_25411,N_24899,N_24780);
or U25412 (N_25412,N_24863,N_24744);
or U25413 (N_25413,N_24947,N_24508);
nor U25414 (N_25414,N_24992,N_24504);
and U25415 (N_25415,N_24934,N_24530);
nand U25416 (N_25416,N_24677,N_24668);
and U25417 (N_25417,N_24997,N_24575);
nor U25418 (N_25418,N_24574,N_24546);
xnor U25419 (N_25419,N_24995,N_24716);
nor U25420 (N_25420,N_24663,N_24650);
and U25421 (N_25421,N_24674,N_24949);
and U25422 (N_25422,N_24599,N_24844);
xnor U25423 (N_25423,N_24638,N_24610);
nor U25424 (N_25424,N_24527,N_24929);
xor U25425 (N_25425,N_24903,N_24832);
nand U25426 (N_25426,N_24712,N_24866);
xor U25427 (N_25427,N_24896,N_24512);
and U25428 (N_25428,N_24582,N_24508);
nand U25429 (N_25429,N_24593,N_24788);
and U25430 (N_25430,N_24781,N_24749);
nor U25431 (N_25431,N_24599,N_24522);
or U25432 (N_25432,N_24565,N_24645);
or U25433 (N_25433,N_24558,N_24680);
or U25434 (N_25434,N_24756,N_24777);
or U25435 (N_25435,N_24683,N_24875);
nand U25436 (N_25436,N_24887,N_24943);
nor U25437 (N_25437,N_24772,N_24642);
and U25438 (N_25438,N_24869,N_24953);
nor U25439 (N_25439,N_24635,N_24709);
xor U25440 (N_25440,N_24914,N_24884);
xnor U25441 (N_25441,N_24888,N_24619);
nor U25442 (N_25442,N_24523,N_24785);
and U25443 (N_25443,N_24966,N_24748);
nand U25444 (N_25444,N_24877,N_24539);
xnor U25445 (N_25445,N_24860,N_24887);
xnor U25446 (N_25446,N_24518,N_24869);
xor U25447 (N_25447,N_24936,N_24691);
nand U25448 (N_25448,N_24688,N_24614);
xnor U25449 (N_25449,N_24601,N_24604);
or U25450 (N_25450,N_24999,N_24580);
and U25451 (N_25451,N_24940,N_24866);
and U25452 (N_25452,N_24646,N_24981);
and U25453 (N_25453,N_24983,N_24949);
nand U25454 (N_25454,N_24770,N_24679);
nor U25455 (N_25455,N_24641,N_24867);
and U25456 (N_25456,N_24777,N_24983);
nor U25457 (N_25457,N_24655,N_24822);
and U25458 (N_25458,N_24641,N_24724);
or U25459 (N_25459,N_24540,N_24909);
xor U25460 (N_25460,N_24841,N_24837);
and U25461 (N_25461,N_24886,N_24718);
xor U25462 (N_25462,N_24881,N_24744);
xor U25463 (N_25463,N_24976,N_24649);
and U25464 (N_25464,N_24577,N_24786);
and U25465 (N_25465,N_24917,N_24522);
nor U25466 (N_25466,N_24570,N_24598);
and U25467 (N_25467,N_24638,N_24849);
and U25468 (N_25468,N_24929,N_24914);
nand U25469 (N_25469,N_24662,N_24968);
nor U25470 (N_25470,N_24980,N_24914);
or U25471 (N_25471,N_24779,N_24661);
or U25472 (N_25472,N_24791,N_24928);
nor U25473 (N_25473,N_24879,N_24528);
xnor U25474 (N_25474,N_24855,N_24932);
nor U25475 (N_25475,N_24902,N_24527);
nor U25476 (N_25476,N_24599,N_24542);
nor U25477 (N_25477,N_24647,N_24679);
nor U25478 (N_25478,N_24788,N_24764);
nor U25479 (N_25479,N_24955,N_24978);
nor U25480 (N_25480,N_24944,N_24812);
or U25481 (N_25481,N_24770,N_24867);
xnor U25482 (N_25482,N_24924,N_24505);
xnor U25483 (N_25483,N_24831,N_24541);
nand U25484 (N_25484,N_24774,N_24506);
and U25485 (N_25485,N_24643,N_24693);
nand U25486 (N_25486,N_24856,N_24850);
xor U25487 (N_25487,N_24604,N_24536);
or U25488 (N_25488,N_24634,N_24772);
nor U25489 (N_25489,N_24753,N_24709);
and U25490 (N_25490,N_24595,N_24761);
xor U25491 (N_25491,N_24794,N_24971);
and U25492 (N_25492,N_24655,N_24594);
nand U25493 (N_25493,N_24782,N_24539);
xor U25494 (N_25494,N_24713,N_24894);
and U25495 (N_25495,N_24618,N_24633);
nand U25496 (N_25496,N_24599,N_24560);
nand U25497 (N_25497,N_24964,N_24635);
xnor U25498 (N_25498,N_24605,N_24828);
nor U25499 (N_25499,N_24741,N_24960);
and U25500 (N_25500,N_25015,N_25306);
xor U25501 (N_25501,N_25158,N_25161);
and U25502 (N_25502,N_25346,N_25344);
nand U25503 (N_25503,N_25123,N_25408);
and U25504 (N_25504,N_25477,N_25374);
nand U25505 (N_25505,N_25108,N_25294);
nor U25506 (N_25506,N_25203,N_25319);
nor U25507 (N_25507,N_25117,N_25036);
and U25508 (N_25508,N_25233,N_25153);
nand U25509 (N_25509,N_25449,N_25366);
xor U25510 (N_25510,N_25225,N_25019);
nand U25511 (N_25511,N_25375,N_25240);
xor U25512 (N_25512,N_25467,N_25013);
xor U25513 (N_25513,N_25051,N_25212);
xor U25514 (N_25514,N_25341,N_25269);
nor U25515 (N_25515,N_25328,N_25050);
xor U25516 (N_25516,N_25043,N_25323);
xor U25517 (N_25517,N_25059,N_25263);
nand U25518 (N_25518,N_25247,N_25245);
and U25519 (N_25519,N_25211,N_25446);
and U25520 (N_25520,N_25264,N_25114);
and U25521 (N_25521,N_25499,N_25170);
or U25522 (N_25522,N_25016,N_25018);
or U25523 (N_25523,N_25388,N_25064);
or U25524 (N_25524,N_25073,N_25389);
xor U25525 (N_25525,N_25033,N_25260);
or U25526 (N_25526,N_25397,N_25066);
nand U25527 (N_25527,N_25201,N_25402);
or U25528 (N_25528,N_25001,N_25125);
and U25529 (N_25529,N_25332,N_25287);
nand U25530 (N_25530,N_25035,N_25055);
and U25531 (N_25531,N_25415,N_25062);
xnor U25532 (N_25532,N_25364,N_25229);
nor U25533 (N_25533,N_25483,N_25451);
nor U25534 (N_25534,N_25098,N_25411);
nand U25535 (N_25535,N_25352,N_25045);
and U25536 (N_25536,N_25488,N_25285);
xnor U25537 (N_25537,N_25453,N_25381);
xor U25538 (N_25538,N_25259,N_25307);
xnor U25539 (N_25539,N_25143,N_25171);
nor U25540 (N_25540,N_25335,N_25262);
or U25541 (N_25541,N_25168,N_25443);
and U25542 (N_25542,N_25003,N_25111);
nand U25543 (N_25543,N_25008,N_25276);
and U25544 (N_25544,N_25215,N_25314);
or U25545 (N_25545,N_25497,N_25138);
and U25546 (N_25546,N_25012,N_25102);
or U25547 (N_25547,N_25345,N_25355);
xnor U25548 (N_25548,N_25057,N_25023);
nand U25549 (N_25549,N_25393,N_25156);
nor U25550 (N_25550,N_25297,N_25442);
nor U25551 (N_25551,N_25096,N_25172);
xnor U25552 (N_25552,N_25126,N_25046);
and U25553 (N_25553,N_25009,N_25014);
nand U25554 (N_25554,N_25079,N_25427);
or U25555 (N_25555,N_25083,N_25282);
nand U25556 (N_25556,N_25007,N_25325);
xor U25557 (N_25557,N_25218,N_25406);
nor U25558 (N_25558,N_25481,N_25095);
xor U25559 (N_25559,N_25464,N_25296);
and U25560 (N_25560,N_25498,N_25140);
nor U25561 (N_25561,N_25040,N_25400);
xnor U25562 (N_25562,N_25152,N_25162);
or U25563 (N_25563,N_25091,N_25025);
nor U25564 (N_25564,N_25405,N_25222);
or U25565 (N_25565,N_25317,N_25458);
or U25566 (N_25566,N_25454,N_25354);
and U25567 (N_25567,N_25430,N_25227);
nor U25568 (N_25568,N_25032,N_25437);
and U25569 (N_25569,N_25137,N_25093);
nand U25570 (N_25570,N_25363,N_25078);
xor U25571 (N_25571,N_25334,N_25353);
or U25572 (N_25572,N_25268,N_25253);
nand U25573 (N_25573,N_25432,N_25252);
or U25574 (N_25574,N_25122,N_25301);
xnor U25575 (N_25575,N_25452,N_25204);
or U25576 (N_25576,N_25136,N_25447);
xor U25577 (N_25577,N_25228,N_25338);
nor U25578 (N_25578,N_25473,N_25283);
and U25579 (N_25579,N_25286,N_25305);
nor U25580 (N_25580,N_25470,N_25132);
nand U25581 (N_25581,N_25075,N_25416);
and U25582 (N_25582,N_25250,N_25261);
or U25583 (N_25583,N_25094,N_25365);
nor U25584 (N_25584,N_25026,N_25217);
xnor U25585 (N_25585,N_25315,N_25490);
xnor U25586 (N_25586,N_25150,N_25254);
or U25587 (N_25587,N_25292,N_25060);
xnor U25588 (N_25588,N_25326,N_25068);
nand U25589 (N_25589,N_25462,N_25348);
nand U25590 (N_25590,N_25076,N_25424);
nor U25591 (N_25591,N_25238,N_25209);
nand U25592 (N_25592,N_25378,N_25082);
nor U25593 (N_25593,N_25255,N_25048);
or U25594 (N_25594,N_25173,N_25113);
and U25595 (N_25595,N_25220,N_25187);
and U25596 (N_25596,N_25193,N_25119);
xnor U25597 (N_25597,N_25109,N_25127);
nand U25598 (N_25598,N_25189,N_25004);
and U25599 (N_25599,N_25207,N_25495);
and U25600 (N_25600,N_25165,N_25100);
nor U25601 (N_25601,N_25199,N_25104);
nand U25602 (N_25602,N_25084,N_25038);
nand U25603 (N_25603,N_25476,N_25129);
xor U25604 (N_25604,N_25281,N_25020);
nor U25605 (N_25605,N_25154,N_25049);
or U25606 (N_25606,N_25249,N_25373);
xor U25607 (N_25607,N_25435,N_25052);
or U25608 (N_25608,N_25144,N_25185);
nand U25609 (N_25609,N_25417,N_25460);
nor U25610 (N_25610,N_25372,N_25112);
nor U25611 (N_25611,N_25368,N_25257);
or U25612 (N_25612,N_25320,N_25438);
xnor U25613 (N_25613,N_25280,N_25339);
nor U25614 (N_25614,N_25478,N_25029);
xnor U25615 (N_25615,N_25466,N_25469);
nand U25616 (N_25616,N_25224,N_25058);
and U25617 (N_25617,N_25006,N_25321);
and U25618 (N_25618,N_25436,N_25433);
nand U25619 (N_25619,N_25146,N_25174);
or U25620 (N_25620,N_25471,N_25316);
xor U25621 (N_25621,N_25128,N_25196);
nand U25622 (N_25622,N_25237,N_25367);
nor U25623 (N_25623,N_25457,N_25248);
nand U25624 (N_25624,N_25230,N_25336);
and U25625 (N_25625,N_25182,N_25309);
nor U25626 (N_25626,N_25439,N_25147);
nand U25627 (N_25627,N_25166,N_25181);
nand U25628 (N_25628,N_25271,N_25420);
and U25629 (N_25629,N_25157,N_25485);
or U25630 (N_25630,N_25422,N_25226);
or U25631 (N_25631,N_25206,N_25221);
and U25632 (N_25632,N_25465,N_25002);
nand U25633 (N_25633,N_25492,N_25392);
nor U25634 (N_25634,N_25074,N_25067);
xnor U25635 (N_25635,N_25005,N_25099);
nand U25636 (N_25636,N_25071,N_25198);
nor U25637 (N_25637,N_25085,N_25480);
nand U25638 (N_25638,N_25407,N_25340);
or U25639 (N_25639,N_25258,N_25299);
xnor U25640 (N_25640,N_25028,N_25149);
nand U25641 (N_25641,N_25333,N_25183);
xnor U25642 (N_25642,N_25298,N_25398);
nor U25643 (N_25643,N_25246,N_25370);
xnor U25644 (N_25644,N_25011,N_25440);
or U25645 (N_25645,N_25429,N_25421);
nand U25646 (N_25646,N_25080,N_25118);
or U25647 (N_25647,N_25061,N_25063);
nor U25648 (N_25648,N_25379,N_25413);
nand U25649 (N_25649,N_25210,N_25054);
and U25650 (N_25650,N_25376,N_25279);
and U25651 (N_25651,N_25031,N_25192);
nand U25652 (N_25652,N_25350,N_25295);
xor U25653 (N_25653,N_25461,N_25359);
nor U25654 (N_25654,N_25382,N_25491);
nor U25655 (N_25655,N_25409,N_25428);
nand U25656 (N_25656,N_25347,N_25337);
and U25657 (N_25657,N_25414,N_25135);
or U25658 (N_25658,N_25419,N_25131);
nand U25659 (N_25659,N_25234,N_25169);
and U25660 (N_25660,N_25110,N_25101);
nand U25661 (N_25661,N_25474,N_25343);
or U25662 (N_25662,N_25342,N_25361);
and U25663 (N_25663,N_25133,N_25444);
or U25664 (N_25664,N_25239,N_25441);
nand U25665 (N_25665,N_25105,N_25041);
and U25666 (N_25666,N_25194,N_25106);
xor U25667 (N_25667,N_25190,N_25115);
and U25668 (N_25668,N_25303,N_25214);
xor U25669 (N_25669,N_25403,N_25308);
and U25670 (N_25670,N_25431,N_25177);
or U25671 (N_25671,N_25145,N_25394);
nand U25672 (N_25672,N_25232,N_25459);
nor U25673 (N_25673,N_25089,N_25056);
or U25674 (N_25674,N_25356,N_25331);
xnor U25675 (N_25675,N_25244,N_25163);
nor U25676 (N_25676,N_25155,N_25081);
and U25677 (N_25677,N_25304,N_25358);
xnor U25678 (N_25678,N_25487,N_25385);
or U25679 (N_25679,N_25065,N_25475);
and U25680 (N_25680,N_25030,N_25103);
and U25681 (N_25681,N_25266,N_25386);
xor U25682 (N_25682,N_25369,N_25213);
nor U25683 (N_25683,N_25494,N_25357);
nor U25684 (N_25684,N_25377,N_25235);
nor U25685 (N_25685,N_25223,N_25330);
xor U25686 (N_25686,N_25399,N_25371);
nor U25687 (N_25687,N_25418,N_25124);
or U25688 (N_25688,N_25463,N_25097);
nor U25689 (N_25689,N_25380,N_25191);
xnor U25690 (N_25690,N_25396,N_25349);
or U25691 (N_25691,N_25037,N_25291);
and U25692 (N_25692,N_25242,N_25017);
nor U25693 (N_25693,N_25412,N_25121);
xnor U25694 (N_25694,N_25278,N_25022);
xor U25695 (N_25695,N_25077,N_25139);
and U25696 (N_25696,N_25236,N_25404);
xnor U25697 (N_25697,N_25024,N_25395);
nand U25698 (N_25698,N_25456,N_25322);
nor U25699 (N_25699,N_25410,N_25274);
or U25700 (N_25700,N_25448,N_25290);
xor U25701 (N_25701,N_25116,N_25482);
or U25702 (N_25702,N_25455,N_25092);
nor U25703 (N_25703,N_25087,N_25327);
nor U25704 (N_25704,N_25180,N_25265);
or U25705 (N_25705,N_25472,N_25318);
and U25706 (N_25706,N_25272,N_25130);
nand U25707 (N_25707,N_25300,N_25426);
and U25708 (N_25708,N_25179,N_25273);
or U25709 (N_25709,N_25205,N_25069);
nor U25710 (N_25710,N_25047,N_25313);
and U25711 (N_25711,N_25027,N_25362);
nand U25712 (N_25712,N_25202,N_25312);
or U25713 (N_25713,N_25151,N_25390);
nor U25714 (N_25714,N_25445,N_25310);
nand U25715 (N_25715,N_25486,N_25425);
and U25716 (N_25716,N_25142,N_25219);
nand U25717 (N_25717,N_25496,N_25284);
nor U25718 (N_25718,N_25120,N_25423);
or U25719 (N_25719,N_25468,N_25383);
nand U25720 (N_25720,N_25450,N_25256);
and U25721 (N_25721,N_25243,N_25197);
nand U25722 (N_25722,N_25010,N_25107);
nand U25723 (N_25723,N_25302,N_25000);
or U25724 (N_25724,N_25360,N_25148);
and U25725 (N_25725,N_25216,N_25042);
or U25726 (N_25726,N_25270,N_25391);
nand U25727 (N_25727,N_25484,N_25267);
nor U25728 (N_25728,N_25141,N_25134);
xnor U25729 (N_25729,N_25208,N_25176);
and U25730 (N_25730,N_25479,N_25384);
and U25731 (N_25731,N_25053,N_25175);
nand U25732 (N_25732,N_25289,N_25288);
nor U25733 (N_25733,N_25088,N_25186);
nand U25734 (N_25734,N_25329,N_25241);
nand U25735 (N_25735,N_25401,N_25188);
nand U25736 (N_25736,N_25070,N_25231);
or U25737 (N_25737,N_25277,N_25184);
nand U25738 (N_25738,N_25293,N_25090);
xor U25739 (N_25739,N_25164,N_25044);
or U25740 (N_25740,N_25178,N_25086);
xnor U25741 (N_25741,N_25021,N_25160);
and U25742 (N_25742,N_25200,N_25251);
and U25743 (N_25743,N_25034,N_25489);
and U25744 (N_25744,N_25039,N_25072);
xnor U25745 (N_25745,N_25159,N_25311);
and U25746 (N_25746,N_25434,N_25324);
and U25747 (N_25747,N_25493,N_25387);
nand U25748 (N_25748,N_25167,N_25195);
nor U25749 (N_25749,N_25351,N_25275);
or U25750 (N_25750,N_25419,N_25262);
or U25751 (N_25751,N_25371,N_25147);
nand U25752 (N_25752,N_25277,N_25031);
nor U25753 (N_25753,N_25258,N_25149);
or U25754 (N_25754,N_25013,N_25413);
and U25755 (N_25755,N_25038,N_25114);
nor U25756 (N_25756,N_25351,N_25350);
nand U25757 (N_25757,N_25315,N_25375);
or U25758 (N_25758,N_25294,N_25379);
nor U25759 (N_25759,N_25423,N_25435);
and U25760 (N_25760,N_25049,N_25214);
nor U25761 (N_25761,N_25287,N_25297);
and U25762 (N_25762,N_25075,N_25405);
or U25763 (N_25763,N_25165,N_25253);
xnor U25764 (N_25764,N_25313,N_25390);
or U25765 (N_25765,N_25249,N_25453);
xor U25766 (N_25766,N_25173,N_25469);
nand U25767 (N_25767,N_25386,N_25264);
and U25768 (N_25768,N_25435,N_25021);
nand U25769 (N_25769,N_25014,N_25415);
or U25770 (N_25770,N_25192,N_25045);
xnor U25771 (N_25771,N_25017,N_25311);
nor U25772 (N_25772,N_25472,N_25207);
nand U25773 (N_25773,N_25409,N_25438);
nand U25774 (N_25774,N_25357,N_25263);
nand U25775 (N_25775,N_25210,N_25298);
or U25776 (N_25776,N_25204,N_25146);
nor U25777 (N_25777,N_25083,N_25047);
nand U25778 (N_25778,N_25328,N_25213);
nand U25779 (N_25779,N_25275,N_25496);
and U25780 (N_25780,N_25497,N_25105);
or U25781 (N_25781,N_25320,N_25474);
xnor U25782 (N_25782,N_25403,N_25495);
or U25783 (N_25783,N_25278,N_25230);
xor U25784 (N_25784,N_25318,N_25422);
or U25785 (N_25785,N_25068,N_25205);
nor U25786 (N_25786,N_25327,N_25259);
xor U25787 (N_25787,N_25329,N_25204);
and U25788 (N_25788,N_25195,N_25069);
and U25789 (N_25789,N_25488,N_25423);
nand U25790 (N_25790,N_25443,N_25097);
nand U25791 (N_25791,N_25433,N_25014);
nand U25792 (N_25792,N_25089,N_25153);
nor U25793 (N_25793,N_25028,N_25208);
nor U25794 (N_25794,N_25031,N_25005);
or U25795 (N_25795,N_25071,N_25347);
xnor U25796 (N_25796,N_25235,N_25093);
or U25797 (N_25797,N_25376,N_25375);
nand U25798 (N_25798,N_25450,N_25461);
and U25799 (N_25799,N_25249,N_25244);
nand U25800 (N_25800,N_25274,N_25220);
nand U25801 (N_25801,N_25067,N_25395);
nand U25802 (N_25802,N_25124,N_25122);
nor U25803 (N_25803,N_25123,N_25211);
or U25804 (N_25804,N_25334,N_25146);
nand U25805 (N_25805,N_25178,N_25212);
xor U25806 (N_25806,N_25472,N_25111);
nand U25807 (N_25807,N_25041,N_25446);
xnor U25808 (N_25808,N_25399,N_25406);
and U25809 (N_25809,N_25270,N_25198);
and U25810 (N_25810,N_25013,N_25043);
nand U25811 (N_25811,N_25468,N_25425);
and U25812 (N_25812,N_25407,N_25193);
nor U25813 (N_25813,N_25326,N_25315);
nor U25814 (N_25814,N_25109,N_25089);
or U25815 (N_25815,N_25089,N_25247);
xor U25816 (N_25816,N_25266,N_25434);
nor U25817 (N_25817,N_25360,N_25369);
nand U25818 (N_25818,N_25069,N_25225);
nand U25819 (N_25819,N_25384,N_25297);
or U25820 (N_25820,N_25417,N_25259);
nand U25821 (N_25821,N_25203,N_25259);
nor U25822 (N_25822,N_25208,N_25348);
nand U25823 (N_25823,N_25077,N_25101);
nor U25824 (N_25824,N_25001,N_25020);
or U25825 (N_25825,N_25220,N_25231);
nor U25826 (N_25826,N_25340,N_25355);
nor U25827 (N_25827,N_25242,N_25432);
nand U25828 (N_25828,N_25280,N_25160);
and U25829 (N_25829,N_25166,N_25211);
or U25830 (N_25830,N_25034,N_25294);
nand U25831 (N_25831,N_25098,N_25025);
xor U25832 (N_25832,N_25448,N_25327);
xnor U25833 (N_25833,N_25177,N_25375);
nand U25834 (N_25834,N_25296,N_25465);
nand U25835 (N_25835,N_25209,N_25401);
xor U25836 (N_25836,N_25493,N_25104);
or U25837 (N_25837,N_25150,N_25380);
nand U25838 (N_25838,N_25426,N_25291);
nor U25839 (N_25839,N_25121,N_25352);
or U25840 (N_25840,N_25391,N_25042);
and U25841 (N_25841,N_25279,N_25460);
and U25842 (N_25842,N_25491,N_25002);
or U25843 (N_25843,N_25269,N_25442);
and U25844 (N_25844,N_25097,N_25163);
nand U25845 (N_25845,N_25217,N_25246);
nor U25846 (N_25846,N_25177,N_25369);
nor U25847 (N_25847,N_25024,N_25052);
or U25848 (N_25848,N_25119,N_25414);
nor U25849 (N_25849,N_25214,N_25435);
and U25850 (N_25850,N_25308,N_25172);
and U25851 (N_25851,N_25059,N_25104);
and U25852 (N_25852,N_25332,N_25187);
xor U25853 (N_25853,N_25411,N_25229);
or U25854 (N_25854,N_25084,N_25220);
nand U25855 (N_25855,N_25168,N_25170);
and U25856 (N_25856,N_25428,N_25025);
or U25857 (N_25857,N_25380,N_25458);
nor U25858 (N_25858,N_25068,N_25057);
nand U25859 (N_25859,N_25401,N_25189);
xnor U25860 (N_25860,N_25492,N_25047);
and U25861 (N_25861,N_25494,N_25065);
or U25862 (N_25862,N_25420,N_25184);
and U25863 (N_25863,N_25122,N_25252);
nor U25864 (N_25864,N_25210,N_25322);
xor U25865 (N_25865,N_25058,N_25321);
nor U25866 (N_25866,N_25230,N_25307);
or U25867 (N_25867,N_25468,N_25074);
nor U25868 (N_25868,N_25255,N_25107);
and U25869 (N_25869,N_25435,N_25260);
or U25870 (N_25870,N_25121,N_25197);
nor U25871 (N_25871,N_25194,N_25108);
xnor U25872 (N_25872,N_25219,N_25497);
xnor U25873 (N_25873,N_25067,N_25444);
nand U25874 (N_25874,N_25111,N_25362);
and U25875 (N_25875,N_25488,N_25038);
and U25876 (N_25876,N_25432,N_25121);
nor U25877 (N_25877,N_25378,N_25003);
nand U25878 (N_25878,N_25378,N_25097);
nor U25879 (N_25879,N_25068,N_25053);
xor U25880 (N_25880,N_25072,N_25128);
nand U25881 (N_25881,N_25375,N_25100);
nor U25882 (N_25882,N_25228,N_25357);
nor U25883 (N_25883,N_25212,N_25343);
and U25884 (N_25884,N_25447,N_25064);
xor U25885 (N_25885,N_25109,N_25162);
or U25886 (N_25886,N_25091,N_25456);
nand U25887 (N_25887,N_25383,N_25267);
and U25888 (N_25888,N_25369,N_25388);
and U25889 (N_25889,N_25447,N_25173);
and U25890 (N_25890,N_25109,N_25153);
or U25891 (N_25891,N_25275,N_25000);
xor U25892 (N_25892,N_25044,N_25079);
xnor U25893 (N_25893,N_25321,N_25220);
or U25894 (N_25894,N_25243,N_25080);
and U25895 (N_25895,N_25046,N_25130);
or U25896 (N_25896,N_25002,N_25382);
or U25897 (N_25897,N_25302,N_25102);
or U25898 (N_25898,N_25144,N_25490);
nor U25899 (N_25899,N_25132,N_25134);
nor U25900 (N_25900,N_25032,N_25043);
and U25901 (N_25901,N_25015,N_25214);
nand U25902 (N_25902,N_25428,N_25251);
and U25903 (N_25903,N_25365,N_25481);
or U25904 (N_25904,N_25005,N_25294);
xnor U25905 (N_25905,N_25341,N_25477);
or U25906 (N_25906,N_25466,N_25360);
and U25907 (N_25907,N_25357,N_25045);
nor U25908 (N_25908,N_25416,N_25234);
xnor U25909 (N_25909,N_25134,N_25234);
or U25910 (N_25910,N_25225,N_25423);
nor U25911 (N_25911,N_25487,N_25164);
xor U25912 (N_25912,N_25490,N_25477);
and U25913 (N_25913,N_25088,N_25048);
or U25914 (N_25914,N_25334,N_25167);
xor U25915 (N_25915,N_25380,N_25122);
or U25916 (N_25916,N_25149,N_25332);
nand U25917 (N_25917,N_25157,N_25371);
xnor U25918 (N_25918,N_25192,N_25059);
and U25919 (N_25919,N_25329,N_25149);
nand U25920 (N_25920,N_25196,N_25376);
or U25921 (N_25921,N_25458,N_25475);
nor U25922 (N_25922,N_25391,N_25182);
nor U25923 (N_25923,N_25198,N_25486);
and U25924 (N_25924,N_25493,N_25107);
and U25925 (N_25925,N_25072,N_25473);
nor U25926 (N_25926,N_25464,N_25057);
or U25927 (N_25927,N_25221,N_25462);
and U25928 (N_25928,N_25339,N_25354);
or U25929 (N_25929,N_25091,N_25328);
or U25930 (N_25930,N_25027,N_25072);
and U25931 (N_25931,N_25491,N_25333);
nand U25932 (N_25932,N_25424,N_25447);
nor U25933 (N_25933,N_25008,N_25497);
and U25934 (N_25934,N_25175,N_25178);
or U25935 (N_25935,N_25154,N_25341);
xnor U25936 (N_25936,N_25079,N_25018);
or U25937 (N_25937,N_25035,N_25373);
nor U25938 (N_25938,N_25249,N_25348);
nand U25939 (N_25939,N_25026,N_25238);
and U25940 (N_25940,N_25115,N_25311);
xnor U25941 (N_25941,N_25396,N_25017);
nor U25942 (N_25942,N_25137,N_25267);
nor U25943 (N_25943,N_25045,N_25482);
nand U25944 (N_25944,N_25016,N_25214);
and U25945 (N_25945,N_25462,N_25293);
nor U25946 (N_25946,N_25328,N_25063);
or U25947 (N_25947,N_25417,N_25072);
nor U25948 (N_25948,N_25260,N_25092);
and U25949 (N_25949,N_25383,N_25495);
and U25950 (N_25950,N_25187,N_25130);
xnor U25951 (N_25951,N_25077,N_25078);
nand U25952 (N_25952,N_25311,N_25474);
and U25953 (N_25953,N_25407,N_25439);
nand U25954 (N_25954,N_25119,N_25164);
nor U25955 (N_25955,N_25463,N_25261);
nand U25956 (N_25956,N_25237,N_25217);
nor U25957 (N_25957,N_25487,N_25071);
nor U25958 (N_25958,N_25153,N_25450);
or U25959 (N_25959,N_25290,N_25084);
nand U25960 (N_25960,N_25221,N_25029);
and U25961 (N_25961,N_25024,N_25361);
xnor U25962 (N_25962,N_25202,N_25484);
xor U25963 (N_25963,N_25199,N_25375);
nand U25964 (N_25964,N_25469,N_25081);
xor U25965 (N_25965,N_25183,N_25342);
nand U25966 (N_25966,N_25146,N_25068);
nor U25967 (N_25967,N_25353,N_25039);
nand U25968 (N_25968,N_25436,N_25468);
and U25969 (N_25969,N_25215,N_25072);
or U25970 (N_25970,N_25467,N_25254);
nor U25971 (N_25971,N_25095,N_25366);
nand U25972 (N_25972,N_25263,N_25336);
xor U25973 (N_25973,N_25025,N_25389);
xnor U25974 (N_25974,N_25006,N_25482);
and U25975 (N_25975,N_25235,N_25168);
and U25976 (N_25976,N_25256,N_25208);
nor U25977 (N_25977,N_25172,N_25451);
nand U25978 (N_25978,N_25066,N_25373);
xor U25979 (N_25979,N_25002,N_25370);
xor U25980 (N_25980,N_25316,N_25160);
or U25981 (N_25981,N_25173,N_25295);
xnor U25982 (N_25982,N_25432,N_25233);
xor U25983 (N_25983,N_25166,N_25321);
xnor U25984 (N_25984,N_25422,N_25170);
nand U25985 (N_25985,N_25408,N_25170);
and U25986 (N_25986,N_25204,N_25211);
xnor U25987 (N_25987,N_25492,N_25251);
xnor U25988 (N_25988,N_25257,N_25355);
xnor U25989 (N_25989,N_25359,N_25463);
nor U25990 (N_25990,N_25321,N_25046);
nand U25991 (N_25991,N_25180,N_25475);
nor U25992 (N_25992,N_25102,N_25075);
nand U25993 (N_25993,N_25188,N_25144);
nor U25994 (N_25994,N_25415,N_25446);
or U25995 (N_25995,N_25129,N_25380);
nand U25996 (N_25996,N_25058,N_25249);
nor U25997 (N_25997,N_25401,N_25400);
and U25998 (N_25998,N_25444,N_25330);
nand U25999 (N_25999,N_25286,N_25280);
nor U26000 (N_26000,N_25796,N_25668);
xor U26001 (N_26001,N_25861,N_25697);
or U26002 (N_26002,N_25510,N_25850);
or U26003 (N_26003,N_25883,N_25684);
nand U26004 (N_26004,N_25725,N_25920);
nor U26005 (N_26005,N_25691,N_25640);
nor U26006 (N_26006,N_25626,N_25613);
xor U26007 (N_26007,N_25873,N_25599);
nor U26008 (N_26008,N_25543,N_25516);
or U26009 (N_26009,N_25635,N_25502);
and U26010 (N_26010,N_25885,N_25577);
xnor U26011 (N_26011,N_25738,N_25655);
nor U26012 (N_26012,N_25528,N_25734);
and U26013 (N_26013,N_25880,N_25786);
or U26014 (N_26014,N_25568,N_25952);
and U26015 (N_26015,N_25532,N_25824);
or U26016 (N_26016,N_25763,N_25932);
nor U26017 (N_26017,N_25926,N_25911);
and U26018 (N_26018,N_25772,N_25614);
and U26019 (N_26019,N_25870,N_25714);
nand U26020 (N_26020,N_25848,N_25740);
and U26021 (N_26021,N_25788,N_25957);
or U26022 (N_26022,N_25852,N_25969);
nor U26023 (N_26023,N_25758,N_25630);
xor U26024 (N_26024,N_25891,N_25807);
nor U26025 (N_26025,N_25994,N_25660);
and U26026 (N_26026,N_25784,N_25524);
and U26027 (N_26027,N_25562,N_25556);
nand U26028 (N_26028,N_25803,N_25898);
nand U26029 (N_26029,N_25579,N_25742);
and U26030 (N_26030,N_25683,N_25962);
xnor U26031 (N_26031,N_25949,N_25942);
nand U26032 (N_26032,N_25592,N_25720);
xnor U26033 (N_26033,N_25708,N_25521);
xnor U26034 (N_26034,N_25959,N_25970);
or U26035 (N_26035,N_25673,N_25547);
xor U26036 (N_26036,N_25927,N_25564);
xor U26037 (N_26037,N_25661,N_25888);
nor U26038 (N_26038,N_25982,N_25875);
nand U26039 (N_26039,N_25641,N_25857);
xor U26040 (N_26040,N_25677,N_25919);
and U26041 (N_26041,N_25585,N_25810);
and U26042 (N_26042,N_25775,N_25862);
xor U26043 (N_26043,N_25569,N_25854);
nand U26044 (N_26044,N_25645,N_25787);
nor U26045 (N_26045,N_25523,N_25715);
nor U26046 (N_26046,N_25505,N_25809);
nor U26047 (N_26047,N_25755,N_25575);
xor U26048 (N_26048,N_25780,N_25933);
nor U26049 (N_26049,N_25754,N_25559);
or U26050 (N_26050,N_25602,N_25611);
and U26051 (N_26051,N_25806,N_25904);
or U26052 (N_26052,N_25582,N_25943);
or U26053 (N_26053,N_25539,N_25800);
xor U26054 (N_26054,N_25596,N_25607);
nand U26055 (N_26055,N_25874,N_25936);
xor U26056 (N_26056,N_25790,N_25998);
and U26057 (N_26057,N_25934,N_25726);
nand U26058 (N_26058,N_25815,N_25624);
nand U26059 (N_26059,N_25767,N_25843);
xor U26060 (N_26060,N_25839,N_25828);
or U26061 (N_26061,N_25567,N_25925);
nor U26062 (N_26062,N_25931,N_25856);
and U26063 (N_26063,N_25517,N_25744);
and U26064 (N_26064,N_25937,N_25902);
xor U26065 (N_26065,N_25694,N_25745);
nand U26066 (N_26066,N_25858,N_25693);
or U26067 (N_26067,N_25968,N_25612);
and U26068 (N_26068,N_25713,N_25853);
xor U26069 (N_26069,N_25500,N_25648);
or U26070 (N_26070,N_25636,N_25945);
or U26071 (N_26071,N_25699,N_25639);
nor U26072 (N_26072,N_25979,N_25651);
xnor U26073 (N_26073,N_25739,N_25899);
nand U26074 (N_26074,N_25650,N_25872);
and U26075 (N_26075,N_25987,N_25804);
or U26076 (N_26076,N_25871,N_25706);
or U26077 (N_26077,N_25997,N_25519);
nor U26078 (N_26078,N_25618,N_25663);
xor U26079 (N_26079,N_25985,N_25869);
and U26080 (N_26080,N_25604,N_25896);
xor U26081 (N_26081,N_25702,N_25769);
nor U26082 (N_26082,N_25783,N_25541);
xnor U26083 (N_26083,N_25595,N_25574);
and U26084 (N_26084,N_25545,N_25721);
or U26085 (N_26085,N_25583,N_25646);
and U26086 (N_26086,N_25566,N_25924);
nor U26087 (N_26087,N_25948,N_25637);
and U26088 (N_26088,N_25940,N_25867);
nand U26089 (N_26089,N_25703,N_25616);
and U26090 (N_26090,N_25548,N_25736);
and U26091 (N_26091,N_25598,N_25581);
or U26092 (N_26092,N_25704,N_25594);
or U26093 (N_26093,N_25676,N_25723);
nand U26094 (N_26094,N_25608,N_25717);
and U26095 (N_26095,N_25895,N_25832);
nor U26096 (N_26096,N_25812,N_25707);
nor U26097 (N_26097,N_25845,N_25833);
xnor U26098 (N_26098,N_25972,N_25733);
or U26099 (N_26099,N_25914,N_25652);
xnor U26100 (N_26100,N_25819,N_25620);
or U26101 (N_26101,N_25849,N_25747);
nand U26102 (N_26102,N_25609,N_25729);
nand U26103 (N_26103,N_25622,N_25792);
or U26104 (N_26104,N_25601,N_25811);
and U26105 (N_26105,N_25752,N_25976);
or U26106 (N_26106,N_25743,N_25808);
or U26107 (N_26107,N_25981,N_25724);
and U26108 (N_26108,N_25915,N_25587);
and U26109 (N_26109,N_25992,N_25791);
or U26110 (N_26110,N_25737,N_25546);
nand U26111 (N_26111,N_25928,N_25503);
or U26112 (N_26112,N_25825,N_25634);
and U26113 (N_26113,N_25750,N_25712);
and U26114 (N_26114,N_25913,N_25536);
nor U26115 (N_26115,N_25906,N_25728);
xor U26116 (N_26116,N_25844,N_25664);
and U26117 (N_26117,N_25561,N_25756);
nor U26118 (N_26118,N_25776,N_25963);
and U26119 (N_26119,N_25671,N_25782);
xnor U26120 (N_26120,N_25638,N_25847);
or U26121 (N_26121,N_25589,N_25966);
nor U26122 (N_26122,N_25781,N_25610);
nand U26123 (N_26123,N_25978,N_25946);
nor U26124 (N_26124,N_25591,N_25537);
and U26125 (N_26125,N_25542,N_25670);
xor U26126 (N_26126,N_25774,N_25525);
or U26127 (N_26127,N_25793,N_25678);
nand U26128 (N_26128,N_25580,N_25615);
or U26129 (N_26129,N_25603,N_25657);
or U26130 (N_26130,N_25965,N_25533);
nor U26131 (N_26131,N_25908,N_25597);
or U26132 (N_26132,N_25778,N_25798);
xor U26133 (N_26133,N_25578,N_25696);
or U26134 (N_26134,N_25964,N_25893);
xor U26135 (N_26135,N_25897,N_25901);
and U26136 (N_26136,N_25674,N_25649);
nor U26137 (N_26137,N_25560,N_25989);
or U26138 (N_26138,N_25866,N_25518);
nand U26139 (N_26139,N_25584,N_25695);
or U26140 (N_26140,N_25923,N_25529);
xnor U26141 (N_26141,N_25573,N_25823);
xor U26142 (N_26142,N_25760,N_25669);
nand U26143 (N_26143,N_25748,N_25540);
nand U26144 (N_26144,N_25753,N_25513);
and U26145 (N_26145,N_25735,N_25509);
nor U26146 (N_26146,N_25859,N_25868);
or U26147 (N_26147,N_25586,N_25889);
and U26148 (N_26148,N_25813,N_25685);
xnor U26149 (N_26149,N_25700,N_25836);
nand U26150 (N_26150,N_25659,N_25617);
nand U26151 (N_26151,N_25797,N_25826);
and U26152 (N_26152,N_25538,N_25958);
nor U26153 (N_26153,N_25731,N_25680);
xnor U26154 (N_26154,N_25551,N_25527);
and U26155 (N_26155,N_25930,N_25802);
or U26156 (N_26156,N_25894,N_25656);
xor U26157 (N_26157,N_25912,N_25710);
xor U26158 (N_26158,N_25785,N_25922);
or U26159 (N_26159,N_25711,N_25950);
nand U26160 (N_26160,N_25688,N_25623);
nand U26161 (N_26161,N_25765,N_25746);
and U26162 (N_26162,N_25590,N_25555);
nand U26163 (N_26163,N_25929,N_25522);
nand U26164 (N_26164,N_25689,N_25827);
and U26165 (N_26165,N_25644,N_25675);
and U26166 (N_26166,N_25829,N_25916);
nand U26167 (N_26167,N_25764,N_25954);
nor U26168 (N_26168,N_25619,N_25531);
xnor U26169 (N_26169,N_25986,N_25990);
xor U26170 (N_26170,N_25658,N_25917);
and U26171 (N_26171,N_25682,N_25773);
xnor U26172 (N_26172,N_25838,N_25890);
nand U26173 (N_26173,N_25840,N_25507);
xnor U26174 (N_26174,N_25818,N_25627);
xnor U26175 (N_26175,N_25771,N_25654);
nor U26176 (N_26176,N_25534,N_25860);
or U26177 (N_26177,N_25980,N_25606);
xor U26178 (N_26178,N_25512,N_25805);
and U26179 (N_26179,N_25955,N_25687);
or U26180 (N_26180,N_25837,N_25768);
nor U26181 (N_26181,N_25701,N_25831);
nand U26182 (N_26182,N_25905,N_25563);
or U26183 (N_26183,N_25718,N_25506);
xor U26184 (N_26184,N_25886,N_25977);
and U26185 (N_26185,N_25552,N_25921);
nor U26186 (N_26186,N_25681,N_25667);
nor U26187 (N_26187,N_25647,N_25762);
or U26188 (N_26188,N_25642,N_25572);
nor U26189 (N_26189,N_25892,N_25789);
xnor U26190 (N_26190,N_25621,N_25851);
nand U26191 (N_26191,N_25960,N_25632);
nor U26192 (N_26192,N_25863,N_25878);
nand U26193 (N_26193,N_25511,N_25625);
nor U26194 (N_26194,N_25757,N_25909);
nor U26195 (N_26195,N_25709,N_25884);
or U26196 (N_26196,N_25554,N_25741);
and U26197 (N_26197,N_25864,N_25935);
nand U26198 (N_26198,N_25938,N_25501);
nand U26199 (N_26199,N_25515,N_25846);
xor U26200 (N_26200,N_25971,N_25588);
nand U26201 (N_26201,N_25841,N_25907);
or U26202 (N_26202,N_25759,N_25751);
and U26203 (N_26203,N_25941,N_25983);
nor U26204 (N_26204,N_25643,N_25947);
xnor U26205 (N_26205,N_25953,N_25991);
or U26206 (N_26206,N_25801,N_25749);
nand U26207 (N_26207,N_25903,N_25821);
or U26208 (N_26208,N_25631,N_25999);
and U26209 (N_26209,N_25557,N_25679);
nand U26210 (N_26210,N_25975,N_25817);
or U26211 (N_26211,N_25877,N_25727);
or U26212 (N_26212,N_25918,N_25719);
nand U26213 (N_26213,N_25973,N_25530);
nor U26214 (N_26214,N_25865,N_25910);
nor U26215 (N_26215,N_25600,N_25722);
xnor U26216 (N_26216,N_25956,N_25520);
or U26217 (N_26217,N_25514,N_25732);
and U26218 (N_26218,N_25944,N_25628);
and U26219 (N_26219,N_25558,N_25526);
xnor U26220 (N_26220,N_25672,N_25855);
xnor U26221 (N_26221,N_25508,N_25665);
xnor U26222 (N_26222,N_25504,N_25794);
nand U26223 (N_26223,N_25988,N_25766);
xnor U26224 (N_26224,N_25770,N_25705);
xor U26225 (N_26225,N_25814,N_25996);
or U26226 (N_26226,N_25822,N_25961);
nand U26227 (N_26227,N_25799,N_25692);
or U26228 (N_26228,N_25834,N_25662);
and U26229 (N_26229,N_25974,N_25881);
nand U26230 (N_26230,N_25995,N_25549);
or U26231 (N_26231,N_25993,N_25876);
nand U26232 (N_26232,N_25550,N_25967);
nand U26233 (N_26233,N_25879,N_25777);
xor U26234 (N_26234,N_25653,N_25605);
nor U26235 (N_26235,N_25951,N_25544);
nor U26236 (N_26236,N_25816,N_25795);
nor U26237 (N_26237,N_25633,N_25761);
and U26238 (N_26238,N_25939,N_25629);
nor U26239 (N_26239,N_25698,N_25830);
nor U26240 (N_26240,N_25779,N_25571);
and U26241 (N_26241,N_25565,N_25882);
nand U26242 (N_26242,N_25835,N_25666);
xnor U26243 (N_26243,N_25984,N_25686);
nor U26244 (N_26244,N_25690,N_25820);
nand U26245 (N_26245,N_25576,N_25535);
or U26246 (N_26246,N_25730,N_25716);
xor U26247 (N_26247,N_25570,N_25553);
xor U26248 (N_26248,N_25887,N_25900);
and U26249 (N_26249,N_25593,N_25842);
and U26250 (N_26250,N_25991,N_25589);
xor U26251 (N_26251,N_25530,N_25684);
nor U26252 (N_26252,N_25567,N_25801);
and U26253 (N_26253,N_25574,N_25555);
nand U26254 (N_26254,N_25638,N_25518);
nor U26255 (N_26255,N_25862,N_25940);
nor U26256 (N_26256,N_25574,N_25803);
xnor U26257 (N_26257,N_25552,N_25655);
nand U26258 (N_26258,N_25840,N_25837);
nand U26259 (N_26259,N_25506,N_25894);
or U26260 (N_26260,N_25668,N_25677);
nor U26261 (N_26261,N_25638,N_25852);
or U26262 (N_26262,N_25542,N_25816);
and U26263 (N_26263,N_25680,N_25710);
and U26264 (N_26264,N_25935,N_25572);
and U26265 (N_26265,N_25813,N_25772);
nor U26266 (N_26266,N_25853,N_25721);
nand U26267 (N_26267,N_25995,N_25984);
and U26268 (N_26268,N_25572,N_25612);
and U26269 (N_26269,N_25580,N_25679);
and U26270 (N_26270,N_25944,N_25619);
and U26271 (N_26271,N_25825,N_25900);
and U26272 (N_26272,N_25648,N_25708);
nor U26273 (N_26273,N_25764,N_25623);
nor U26274 (N_26274,N_25963,N_25823);
nand U26275 (N_26275,N_25968,N_25662);
and U26276 (N_26276,N_25874,N_25989);
or U26277 (N_26277,N_25548,N_25927);
nor U26278 (N_26278,N_25985,N_25836);
nor U26279 (N_26279,N_25582,N_25901);
or U26280 (N_26280,N_25508,N_25782);
nor U26281 (N_26281,N_25929,N_25907);
nand U26282 (N_26282,N_25951,N_25676);
or U26283 (N_26283,N_25859,N_25905);
nor U26284 (N_26284,N_25736,N_25923);
and U26285 (N_26285,N_25798,N_25734);
or U26286 (N_26286,N_25942,N_25576);
nor U26287 (N_26287,N_25979,N_25802);
nand U26288 (N_26288,N_25803,N_25698);
and U26289 (N_26289,N_25810,N_25915);
nor U26290 (N_26290,N_25784,N_25981);
nor U26291 (N_26291,N_25786,N_25933);
xor U26292 (N_26292,N_25602,N_25695);
xor U26293 (N_26293,N_25582,N_25854);
or U26294 (N_26294,N_25829,N_25563);
or U26295 (N_26295,N_25895,N_25904);
and U26296 (N_26296,N_25542,N_25676);
or U26297 (N_26297,N_25779,N_25868);
nor U26298 (N_26298,N_25660,N_25813);
nor U26299 (N_26299,N_25646,N_25777);
nor U26300 (N_26300,N_25890,N_25920);
nand U26301 (N_26301,N_25831,N_25959);
and U26302 (N_26302,N_25796,N_25991);
and U26303 (N_26303,N_25931,N_25731);
and U26304 (N_26304,N_25794,N_25508);
nor U26305 (N_26305,N_25550,N_25798);
xor U26306 (N_26306,N_25723,N_25513);
or U26307 (N_26307,N_25859,N_25945);
xor U26308 (N_26308,N_25913,N_25885);
nor U26309 (N_26309,N_25852,N_25529);
nand U26310 (N_26310,N_25665,N_25817);
and U26311 (N_26311,N_25585,N_25921);
nor U26312 (N_26312,N_25574,N_25947);
or U26313 (N_26313,N_25915,N_25672);
xnor U26314 (N_26314,N_25980,N_25712);
or U26315 (N_26315,N_25788,N_25853);
and U26316 (N_26316,N_25520,N_25505);
and U26317 (N_26317,N_25989,N_25963);
nor U26318 (N_26318,N_25634,N_25694);
and U26319 (N_26319,N_25856,N_25995);
or U26320 (N_26320,N_25750,N_25533);
and U26321 (N_26321,N_25813,N_25535);
nor U26322 (N_26322,N_25693,N_25603);
and U26323 (N_26323,N_25737,N_25669);
xor U26324 (N_26324,N_25763,N_25992);
or U26325 (N_26325,N_25702,N_25880);
or U26326 (N_26326,N_25865,N_25955);
nand U26327 (N_26327,N_25614,N_25822);
or U26328 (N_26328,N_25897,N_25597);
xor U26329 (N_26329,N_25605,N_25585);
nand U26330 (N_26330,N_25816,N_25980);
and U26331 (N_26331,N_25922,N_25792);
and U26332 (N_26332,N_25553,N_25828);
nand U26333 (N_26333,N_25950,N_25980);
and U26334 (N_26334,N_25993,N_25806);
or U26335 (N_26335,N_25621,N_25501);
nor U26336 (N_26336,N_25929,N_25565);
xnor U26337 (N_26337,N_25688,N_25555);
nor U26338 (N_26338,N_25841,N_25965);
nor U26339 (N_26339,N_25998,N_25692);
and U26340 (N_26340,N_25980,N_25734);
and U26341 (N_26341,N_25843,N_25934);
and U26342 (N_26342,N_25633,N_25728);
and U26343 (N_26343,N_25846,N_25776);
xor U26344 (N_26344,N_25538,N_25607);
nand U26345 (N_26345,N_25622,N_25603);
and U26346 (N_26346,N_25980,N_25800);
nand U26347 (N_26347,N_25674,N_25758);
xnor U26348 (N_26348,N_25589,N_25555);
or U26349 (N_26349,N_25986,N_25881);
nand U26350 (N_26350,N_25710,N_25744);
nand U26351 (N_26351,N_25665,N_25961);
nor U26352 (N_26352,N_25928,N_25956);
nand U26353 (N_26353,N_25766,N_25874);
nand U26354 (N_26354,N_25960,N_25881);
xor U26355 (N_26355,N_25888,N_25884);
nor U26356 (N_26356,N_25609,N_25560);
nand U26357 (N_26357,N_25700,N_25802);
and U26358 (N_26358,N_25687,N_25967);
or U26359 (N_26359,N_25791,N_25642);
and U26360 (N_26360,N_25968,N_25886);
xor U26361 (N_26361,N_25895,N_25626);
xor U26362 (N_26362,N_25542,N_25685);
xnor U26363 (N_26363,N_25852,N_25839);
or U26364 (N_26364,N_25608,N_25986);
and U26365 (N_26365,N_25835,N_25668);
nand U26366 (N_26366,N_25563,N_25729);
and U26367 (N_26367,N_25980,N_25744);
xor U26368 (N_26368,N_25929,N_25539);
nor U26369 (N_26369,N_25888,N_25969);
nand U26370 (N_26370,N_25556,N_25584);
xnor U26371 (N_26371,N_25838,N_25695);
nor U26372 (N_26372,N_25583,N_25592);
nor U26373 (N_26373,N_25503,N_25883);
nor U26374 (N_26374,N_25989,N_25564);
or U26375 (N_26375,N_25581,N_25603);
xor U26376 (N_26376,N_25684,N_25778);
and U26377 (N_26377,N_25891,N_25604);
or U26378 (N_26378,N_25943,N_25581);
nand U26379 (N_26379,N_25684,N_25732);
and U26380 (N_26380,N_25720,N_25630);
or U26381 (N_26381,N_25682,N_25655);
nor U26382 (N_26382,N_25613,N_25846);
or U26383 (N_26383,N_25893,N_25743);
nand U26384 (N_26384,N_25794,N_25517);
nor U26385 (N_26385,N_25748,N_25792);
nor U26386 (N_26386,N_25924,N_25726);
nor U26387 (N_26387,N_25937,N_25567);
or U26388 (N_26388,N_25702,N_25839);
and U26389 (N_26389,N_25894,N_25518);
or U26390 (N_26390,N_25966,N_25855);
xor U26391 (N_26391,N_25532,N_25696);
or U26392 (N_26392,N_25680,N_25825);
nand U26393 (N_26393,N_25697,N_25998);
nand U26394 (N_26394,N_25617,N_25595);
nand U26395 (N_26395,N_25957,N_25820);
and U26396 (N_26396,N_25564,N_25509);
and U26397 (N_26397,N_25971,N_25556);
and U26398 (N_26398,N_25894,N_25565);
and U26399 (N_26399,N_25951,N_25689);
or U26400 (N_26400,N_25832,N_25680);
and U26401 (N_26401,N_25884,N_25996);
or U26402 (N_26402,N_25875,N_25654);
nor U26403 (N_26403,N_25961,N_25942);
or U26404 (N_26404,N_25514,N_25638);
and U26405 (N_26405,N_25838,N_25617);
xnor U26406 (N_26406,N_25957,N_25930);
or U26407 (N_26407,N_25699,N_25890);
and U26408 (N_26408,N_25699,N_25646);
or U26409 (N_26409,N_25977,N_25773);
xnor U26410 (N_26410,N_25983,N_25931);
nand U26411 (N_26411,N_25537,N_25667);
or U26412 (N_26412,N_25982,N_25992);
or U26413 (N_26413,N_25545,N_25894);
nand U26414 (N_26414,N_25878,N_25637);
and U26415 (N_26415,N_25674,N_25810);
nor U26416 (N_26416,N_25860,N_25571);
nand U26417 (N_26417,N_25551,N_25687);
and U26418 (N_26418,N_25508,N_25699);
nor U26419 (N_26419,N_25765,N_25946);
nand U26420 (N_26420,N_25999,N_25533);
or U26421 (N_26421,N_25934,N_25846);
nor U26422 (N_26422,N_25995,N_25685);
xor U26423 (N_26423,N_25871,N_25569);
xnor U26424 (N_26424,N_25762,N_25639);
nand U26425 (N_26425,N_25755,N_25686);
and U26426 (N_26426,N_25934,N_25704);
xnor U26427 (N_26427,N_25554,N_25860);
or U26428 (N_26428,N_25930,N_25701);
or U26429 (N_26429,N_25568,N_25776);
and U26430 (N_26430,N_25902,N_25867);
xor U26431 (N_26431,N_25963,N_25637);
nand U26432 (N_26432,N_25946,N_25673);
and U26433 (N_26433,N_25522,N_25547);
or U26434 (N_26434,N_25905,N_25815);
nor U26435 (N_26435,N_25858,N_25606);
nor U26436 (N_26436,N_25750,N_25937);
or U26437 (N_26437,N_25660,N_25936);
or U26438 (N_26438,N_25751,N_25788);
xnor U26439 (N_26439,N_25863,N_25992);
nand U26440 (N_26440,N_25984,N_25936);
nor U26441 (N_26441,N_25671,N_25514);
nand U26442 (N_26442,N_25621,N_25753);
xnor U26443 (N_26443,N_25665,N_25504);
nor U26444 (N_26444,N_25896,N_25528);
and U26445 (N_26445,N_25864,N_25972);
xnor U26446 (N_26446,N_25668,N_25563);
or U26447 (N_26447,N_25949,N_25516);
nand U26448 (N_26448,N_25907,N_25972);
or U26449 (N_26449,N_25766,N_25896);
nor U26450 (N_26450,N_25759,N_25546);
nand U26451 (N_26451,N_25902,N_25818);
or U26452 (N_26452,N_25977,N_25873);
xor U26453 (N_26453,N_25677,N_25525);
nand U26454 (N_26454,N_25601,N_25810);
nand U26455 (N_26455,N_25658,N_25557);
xor U26456 (N_26456,N_25766,N_25738);
and U26457 (N_26457,N_25883,N_25944);
nor U26458 (N_26458,N_25650,N_25611);
and U26459 (N_26459,N_25638,N_25646);
nand U26460 (N_26460,N_25981,N_25543);
and U26461 (N_26461,N_25517,N_25941);
or U26462 (N_26462,N_25518,N_25876);
and U26463 (N_26463,N_25990,N_25873);
and U26464 (N_26464,N_25984,N_25650);
nor U26465 (N_26465,N_25690,N_25786);
xnor U26466 (N_26466,N_25857,N_25706);
or U26467 (N_26467,N_25916,N_25632);
or U26468 (N_26468,N_25638,N_25950);
xnor U26469 (N_26469,N_25889,N_25979);
or U26470 (N_26470,N_25612,N_25735);
and U26471 (N_26471,N_25634,N_25878);
xnor U26472 (N_26472,N_25801,N_25785);
nand U26473 (N_26473,N_25990,N_25945);
and U26474 (N_26474,N_25870,N_25847);
and U26475 (N_26475,N_25902,N_25802);
xnor U26476 (N_26476,N_25831,N_25747);
xnor U26477 (N_26477,N_25864,N_25791);
nand U26478 (N_26478,N_25948,N_25885);
xnor U26479 (N_26479,N_25600,N_25575);
nand U26480 (N_26480,N_25750,N_25601);
xnor U26481 (N_26481,N_25570,N_25566);
xnor U26482 (N_26482,N_25877,N_25794);
xor U26483 (N_26483,N_25870,N_25607);
and U26484 (N_26484,N_25583,N_25982);
xnor U26485 (N_26485,N_25919,N_25739);
or U26486 (N_26486,N_25677,N_25928);
and U26487 (N_26487,N_25550,N_25546);
and U26488 (N_26488,N_25647,N_25821);
and U26489 (N_26489,N_25795,N_25535);
and U26490 (N_26490,N_25820,N_25727);
xnor U26491 (N_26491,N_25531,N_25747);
nor U26492 (N_26492,N_25521,N_25910);
or U26493 (N_26493,N_25924,N_25758);
and U26494 (N_26494,N_25783,N_25890);
or U26495 (N_26495,N_25835,N_25538);
or U26496 (N_26496,N_25918,N_25716);
xor U26497 (N_26497,N_25717,N_25742);
xnor U26498 (N_26498,N_25992,N_25550);
nor U26499 (N_26499,N_25608,N_25553);
or U26500 (N_26500,N_26191,N_26382);
and U26501 (N_26501,N_26195,N_26045);
and U26502 (N_26502,N_26440,N_26247);
nor U26503 (N_26503,N_26465,N_26262);
nor U26504 (N_26504,N_26277,N_26105);
and U26505 (N_26505,N_26334,N_26080);
nor U26506 (N_26506,N_26032,N_26222);
nand U26507 (N_26507,N_26321,N_26455);
and U26508 (N_26508,N_26299,N_26364);
or U26509 (N_26509,N_26392,N_26237);
or U26510 (N_26510,N_26259,N_26429);
or U26511 (N_26511,N_26112,N_26064);
or U26512 (N_26512,N_26088,N_26043);
xnor U26513 (N_26513,N_26090,N_26154);
nand U26514 (N_26514,N_26451,N_26342);
nor U26515 (N_26515,N_26493,N_26351);
or U26516 (N_26516,N_26478,N_26256);
xnor U26517 (N_26517,N_26018,N_26404);
nand U26518 (N_26518,N_26196,N_26391);
or U26519 (N_26519,N_26374,N_26115);
nor U26520 (N_26520,N_26483,N_26225);
nand U26521 (N_26521,N_26120,N_26179);
nand U26522 (N_26522,N_26371,N_26425);
xor U26523 (N_26523,N_26092,N_26298);
or U26524 (N_26524,N_26056,N_26280);
nor U26525 (N_26525,N_26472,N_26111);
and U26526 (N_26526,N_26294,N_26014);
or U26527 (N_26527,N_26323,N_26049);
nand U26528 (N_26528,N_26175,N_26012);
nor U26529 (N_26529,N_26213,N_26362);
or U26530 (N_26530,N_26171,N_26481);
nor U26531 (N_26531,N_26135,N_26331);
xnor U26532 (N_26532,N_26082,N_26091);
and U26533 (N_26533,N_26123,N_26424);
xnor U26534 (N_26534,N_26075,N_26365);
or U26535 (N_26535,N_26022,N_26060);
and U26536 (N_26536,N_26416,N_26489);
xnor U26537 (N_26537,N_26488,N_26445);
xnor U26538 (N_26538,N_26305,N_26418);
or U26539 (N_26539,N_26227,N_26132);
and U26540 (N_26540,N_26485,N_26363);
xnor U26541 (N_26541,N_26077,N_26428);
and U26542 (N_26542,N_26186,N_26332);
nand U26543 (N_26543,N_26347,N_26410);
or U26544 (N_26544,N_26017,N_26005);
nand U26545 (N_26545,N_26435,N_26098);
xor U26546 (N_26546,N_26315,N_26184);
nor U26547 (N_26547,N_26333,N_26031);
nand U26548 (N_26548,N_26216,N_26456);
nand U26549 (N_26549,N_26433,N_26140);
nor U26550 (N_26550,N_26272,N_26193);
and U26551 (N_26551,N_26036,N_26176);
nor U26552 (N_26552,N_26393,N_26151);
or U26553 (N_26553,N_26177,N_26172);
and U26554 (N_26554,N_26412,N_26265);
or U26555 (N_26555,N_26198,N_26245);
and U26556 (N_26556,N_26073,N_26377);
xnor U26557 (N_26557,N_26288,N_26419);
nand U26558 (N_26558,N_26449,N_26166);
nor U26559 (N_26559,N_26128,N_26182);
or U26560 (N_26560,N_26352,N_26349);
xnor U26561 (N_26561,N_26441,N_26070);
nand U26562 (N_26562,N_26477,N_26139);
nor U26563 (N_26563,N_26069,N_26313);
or U26564 (N_26564,N_26055,N_26284);
xnor U26565 (N_26565,N_26226,N_26215);
nor U26566 (N_26566,N_26137,N_26345);
xor U26567 (N_26567,N_26348,N_26497);
xor U26568 (N_26568,N_26264,N_26223);
or U26569 (N_26569,N_26181,N_26214);
or U26570 (N_26570,N_26071,N_26311);
nor U26571 (N_26571,N_26430,N_26464);
or U26572 (N_26572,N_26194,N_26443);
or U26573 (N_26573,N_26230,N_26384);
or U26574 (N_26574,N_26189,N_26356);
or U26575 (N_26575,N_26268,N_26087);
nand U26576 (N_26576,N_26174,N_26233);
nor U26577 (N_26577,N_26234,N_26006);
nor U26578 (N_26578,N_26258,N_26355);
nor U26579 (N_26579,N_26178,N_26318);
or U26580 (N_26580,N_26468,N_26496);
nor U26581 (N_26581,N_26307,N_26257);
nor U26582 (N_26582,N_26113,N_26165);
nand U26583 (N_26583,N_26293,N_26336);
xor U26584 (N_26584,N_26415,N_26490);
and U26585 (N_26585,N_26303,N_26471);
nand U26586 (N_26586,N_26252,N_26061);
or U26587 (N_26587,N_26266,N_26357);
and U26588 (N_26588,N_26057,N_26021);
xnor U26589 (N_26589,N_26386,N_26063);
xor U26590 (N_26590,N_26224,N_26188);
and U26591 (N_26591,N_26089,N_26370);
and U26592 (N_26592,N_26450,N_26251);
and U26593 (N_26593,N_26387,N_26281);
nor U26594 (N_26594,N_26327,N_26062);
nand U26595 (N_26595,N_26326,N_26405);
xnor U26596 (N_26596,N_26218,N_26271);
xor U26597 (N_26597,N_26422,N_26246);
xnor U26598 (N_26598,N_26129,N_26187);
nand U26599 (N_26599,N_26495,N_26448);
nand U26600 (N_26600,N_26461,N_26379);
and U26601 (N_26601,N_26125,N_26053);
and U26602 (N_26602,N_26499,N_26316);
xor U26603 (N_26603,N_26396,N_26388);
or U26604 (N_26604,N_26086,N_26236);
nand U26605 (N_26605,N_26058,N_26343);
and U26606 (N_26606,N_26161,N_26498);
nand U26607 (N_26607,N_26205,N_26402);
xnor U26608 (N_26608,N_26152,N_26423);
xor U26609 (N_26609,N_26003,N_26159);
or U26610 (N_26610,N_26400,N_26104);
xnor U26611 (N_26611,N_26397,N_26426);
nand U26612 (N_26612,N_26029,N_26038);
or U26613 (N_26613,N_26147,N_26011);
nor U26614 (N_26614,N_26420,N_26249);
nor U26615 (N_26615,N_26118,N_26395);
nand U26616 (N_26616,N_26050,N_26285);
or U26617 (N_26617,N_26150,N_26354);
or U26618 (N_26618,N_26040,N_26008);
xnor U26619 (N_26619,N_26051,N_26406);
and U26620 (N_26620,N_26106,N_26241);
and U26621 (N_26621,N_26367,N_26009);
nor U26622 (N_26622,N_26119,N_26452);
and U26623 (N_26623,N_26254,N_26399);
and U26624 (N_26624,N_26207,N_26183);
and U26625 (N_26625,N_26099,N_26028);
xnor U26626 (N_26626,N_26155,N_26153);
xnor U26627 (N_26627,N_26231,N_26217);
nor U26628 (N_26628,N_26344,N_26286);
or U26629 (N_26629,N_26476,N_26039);
xor U26630 (N_26630,N_26110,N_26494);
or U26631 (N_26631,N_26016,N_26243);
xor U26632 (N_26632,N_26211,N_26117);
xor U26633 (N_26633,N_26170,N_26442);
nor U26634 (N_26634,N_26295,N_26078);
nand U26635 (N_26635,N_26304,N_26296);
nand U26636 (N_26636,N_26096,N_26221);
nor U26637 (N_26637,N_26001,N_26401);
xnor U26638 (N_26638,N_26491,N_26368);
xor U26639 (N_26639,N_26261,N_26066);
nand U26640 (N_26640,N_26042,N_26000);
or U26641 (N_26641,N_26270,N_26173);
nand U26642 (N_26642,N_26358,N_26143);
and U26643 (N_26643,N_26025,N_26320);
or U26644 (N_26644,N_26127,N_26130);
and U26645 (N_26645,N_26201,N_26157);
nand U26646 (N_26646,N_26287,N_26024);
and U26647 (N_26647,N_26475,N_26065);
or U26648 (N_26648,N_26330,N_26302);
nor U26649 (N_26649,N_26030,N_26116);
xnor U26650 (N_26650,N_26164,N_26375);
and U26651 (N_26651,N_26467,N_26114);
nand U26652 (N_26652,N_26010,N_26454);
and U26653 (N_26653,N_26278,N_26260);
nand U26654 (N_26654,N_26235,N_26479);
nor U26655 (N_26655,N_26160,N_26054);
or U26656 (N_26656,N_26212,N_26250);
xor U26657 (N_26657,N_26228,N_26473);
and U26658 (N_26658,N_26121,N_26200);
xor U26659 (N_26659,N_26308,N_26136);
nor U26660 (N_26660,N_26074,N_26142);
xnor U26661 (N_26661,N_26366,N_26197);
or U26662 (N_26662,N_26353,N_26329);
nor U26663 (N_26663,N_26108,N_26274);
nor U26664 (N_26664,N_26163,N_26289);
nor U26665 (N_26665,N_26421,N_26390);
or U26666 (N_26666,N_26141,N_26403);
xor U26667 (N_26667,N_26457,N_26168);
nor U26668 (N_26668,N_26037,N_26148);
and U26669 (N_26669,N_26310,N_26301);
nand U26670 (N_26670,N_26431,N_26297);
nor U26671 (N_26671,N_26269,N_26378);
nand U26672 (N_26672,N_26324,N_26340);
and U26673 (N_26673,N_26480,N_26026);
and U26674 (N_26674,N_26094,N_26041);
or U26675 (N_26675,N_26263,N_26109);
or U26676 (N_26676,N_26047,N_26462);
xnor U26677 (N_26677,N_26439,N_26275);
or U26678 (N_26678,N_26338,N_26414);
nor U26679 (N_26679,N_26460,N_26020);
or U26680 (N_26680,N_26255,N_26447);
nor U26681 (N_26681,N_26267,N_26328);
or U26682 (N_26682,N_26007,N_26209);
or U26683 (N_26683,N_26232,N_26015);
nor U26684 (N_26684,N_26239,N_26474);
nor U26685 (N_26685,N_26202,N_26314);
and U26686 (N_26686,N_26122,N_26072);
or U26687 (N_26687,N_26048,N_26102);
xor U26688 (N_26688,N_26145,N_26359);
or U26689 (N_26689,N_26282,N_26046);
and U26690 (N_26690,N_26023,N_26002);
nand U26691 (N_26691,N_26124,N_26131);
or U26692 (N_26692,N_26436,N_26156);
nor U26693 (N_26693,N_26079,N_26149);
or U26694 (N_26694,N_26244,N_26229);
nand U26695 (N_26695,N_26167,N_26210);
xnor U26696 (N_26696,N_26335,N_26453);
or U26697 (N_26697,N_26059,N_26219);
xnor U26698 (N_26698,N_26407,N_26291);
nand U26699 (N_26699,N_26097,N_26095);
and U26700 (N_26700,N_26319,N_26417);
xor U26701 (N_26701,N_26437,N_26434);
nor U26702 (N_26702,N_26103,N_26385);
or U26703 (N_26703,N_26411,N_26484);
xor U26704 (N_26704,N_26279,N_26208);
nand U26705 (N_26705,N_26067,N_26276);
nor U26706 (N_26706,N_26180,N_26206);
and U26707 (N_26707,N_26083,N_26346);
nand U26708 (N_26708,N_26459,N_26427);
xor U26709 (N_26709,N_26192,N_26482);
xor U26710 (N_26710,N_26238,N_26413);
nand U26711 (N_26711,N_26027,N_26013);
xor U26712 (N_26712,N_26019,N_26081);
or U26713 (N_26713,N_26133,N_26381);
nand U26714 (N_26714,N_26034,N_26470);
or U26715 (N_26715,N_26350,N_26076);
and U26716 (N_26716,N_26052,N_26273);
nor U26717 (N_26717,N_26486,N_26492);
or U26718 (N_26718,N_26101,N_26389);
or U26719 (N_26719,N_26292,N_26369);
xnor U26720 (N_26720,N_26068,N_26376);
and U26721 (N_26721,N_26085,N_26100);
and U26722 (N_26722,N_26487,N_26373);
and U26723 (N_26723,N_26204,N_26337);
nand U26724 (N_26724,N_26312,N_26169);
nand U26725 (N_26725,N_26199,N_26146);
nor U26726 (N_26726,N_26469,N_26126);
or U26727 (N_26727,N_26162,N_26394);
or U26728 (N_26728,N_26325,N_26300);
or U26729 (N_26729,N_26138,N_26408);
or U26730 (N_26730,N_26383,N_26283);
nand U26731 (N_26731,N_26309,N_26290);
nand U26732 (N_26732,N_26463,N_26360);
nor U26733 (N_26733,N_26398,N_26190);
nor U26734 (N_26734,N_26240,N_26004);
nor U26735 (N_26735,N_26220,N_26084);
nor U26736 (N_26736,N_26253,N_26380);
xnor U26737 (N_26737,N_26322,N_26093);
and U26738 (N_26738,N_26409,N_26432);
or U26739 (N_26739,N_26203,N_26339);
nor U26740 (N_26740,N_26134,N_26044);
or U26741 (N_26741,N_26458,N_26317);
and U26742 (N_26742,N_26035,N_26466);
and U26743 (N_26743,N_26444,N_26438);
or U26744 (N_26744,N_26158,N_26372);
and U26745 (N_26745,N_26341,N_26107);
xnor U26746 (N_26746,N_26248,N_26361);
xor U26747 (N_26747,N_26446,N_26033);
xnor U26748 (N_26748,N_26185,N_26306);
nor U26749 (N_26749,N_26242,N_26144);
nor U26750 (N_26750,N_26490,N_26059);
xnor U26751 (N_26751,N_26021,N_26182);
xor U26752 (N_26752,N_26319,N_26390);
xor U26753 (N_26753,N_26134,N_26321);
nor U26754 (N_26754,N_26495,N_26273);
nor U26755 (N_26755,N_26370,N_26147);
and U26756 (N_26756,N_26020,N_26022);
nor U26757 (N_26757,N_26324,N_26339);
nor U26758 (N_26758,N_26068,N_26378);
and U26759 (N_26759,N_26344,N_26135);
and U26760 (N_26760,N_26380,N_26042);
xor U26761 (N_26761,N_26458,N_26415);
nor U26762 (N_26762,N_26170,N_26341);
xnor U26763 (N_26763,N_26060,N_26115);
or U26764 (N_26764,N_26459,N_26489);
and U26765 (N_26765,N_26125,N_26405);
and U26766 (N_26766,N_26442,N_26035);
nor U26767 (N_26767,N_26407,N_26228);
xnor U26768 (N_26768,N_26486,N_26111);
and U26769 (N_26769,N_26172,N_26406);
xor U26770 (N_26770,N_26460,N_26184);
nor U26771 (N_26771,N_26135,N_26210);
or U26772 (N_26772,N_26163,N_26465);
xor U26773 (N_26773,N_26346,N_26263);
nand U26774 (N_26774,N_26318,N_26284);
and U26775 (N_26775,N_26490,N_26096);
xor U26776 (N_26776,N_26207,N_26273);
or U26777 (N_26777,N_26343,N_26441);
and U26778 (N_26778,N_26489,N_26280);
nand U26779 (N_26779,N_26193,N_26495);
nor U26780 (N_26780,N_26422,N_26001);
or U26781 (N_26781,N_26213,N_26044);
or U26782 (N_26782,N_26284,N_26074);
nor U26783 (N_26783,N_26194,N_26416);
or U26784 (N_26784,N_26229,N_26239);
nand U26785 (N_26785,N_26144,N_26248);
or U26786 (N_26786,N_26492,N_26047);
or U26787 (N_26787,N_26227,N_26117);
nand U26788 (N_26788,N_26240,N_26470);
nand U26789 (N_26789,N_26419,N_26228);
and U26790 (N_26790,N_26415,N_26273);
xnor U26791 (N_26791,N_26166,N_26152);
nand U26792 (N_26792,N_26138,N_26004);
or U26793 (N_26793,N_26208,N_26061);
xnor U26794 (N_26794,N_26467,N_26291);
or U26795 (N_26795,N_26265,N_26304);
xnor U26796 (N_26796,N_26016,N_26219);
nor U26797 (N_26797,N_26474,N_26425);
nor U26798 (N_26798,N_26190,N_26022);
and U26799 (N_26799,N_26192,N_26075);
nand U26800 (N_26800,N_26457,N_26004);
nor U26801 (N_26801,N_26211,N_26218);
xor U26802 (N_26802,N_26187,N_26105);
nand U26803 (N_26803,N_26036,N_26364);
or U26804 (N_26804,N_26395,N_26282);
nand U26805 (N_26805,N_26250,N_26159);
or U26806 (N_26806,N_26139,N_26040);
nor U26807 (N_26807,N_26398,N_26348);
and U26808 (N_26808,N_26296,N_26320);
xnor U26809 (N_26809,N_26215,N_26330);
xor U26810 (N_26810,N_26004,N_26460);
nor U26811 (N_26811,N_26186,N_26088);
xor U26812 (N_26812,N_26209,N_26474);
xnor U26813 (N_26813,N_26027,N_26067);
nand U26814 (N_26814,N_26003,N_26020);
nor U26815 (N_26815,N_26209,N_26388);
nand U26816 (N_26816,N_26278,N_26062);
or U26817 (N_26817,N_26478,N_26467);
nand U26818 (N_26818,N_26109,N_26191);
or U26819 (N_26819,N_26003,N_26332);
nand U26820 (N_26820,N_26305,N_26442);
nor U26821 (N_26821,N_26062,N_26454);
nor U26822 (N_26822,N_26489,N_26396);
nand U26823 (N_26823,N_26353,N_26175);
nand U26824 (N_26824,N_26247,N_26345);
and U26825 (N_26825,N_26075,N_26028);
and U26826 (N_26826,N_26211,N_26068);
and U26827 (N_26827,N_26064,N_26166);
nand U26828 (N_26828,N_26228,N_26157);
and U26829 (N_26829,N_26492,N_26156);
and U26830 (N_26830,N_26086,N_26302);
nor U26831 (N_26831,N_26148,N_26287);
nor U26832 (N_26832,N_26399,N_26264);
and U26833 (N_26833,N_26030,N_26019);
and U26834 (N_26834,N_26145,N_26319);
xor U26835 (N_26835,N_26097,N_26450);
or U26836 (N_26836,N_26418,N_26215);
nand U26837 (N_26837,N_26037,N_26337);
xnor U26838 (N_26838,N_26441,N_26270);
and U26839 (N_26839,N_26463,N_26348);
and U26840 (N_26840,N_26466,N_26425);
and U26841 (N_26841,N_26114,N_26300);
nand U26842 (N_26842,N_26186,N_26215);
nor U26843 (N_26843,N_26121,N_26144);
and U26844 (N_26844,N_26221,N_26276);
nor U26845 (N_26845,N_26277,N_26020);
or U26846 (N_26846,N_26150,N_26312);
or U26847 (N_26847,N_26218,N_26216);
nand U26848 (N_26848,N_26362,N_26186);
nand U26849 (N_26849,N_26263,N_26295);
or U26850 (N_26850,N_26098,N_26336);
nand U26851 (N_26851,N_26277,N_26198);
xnor U26852 (N_26852,N_26248,N_26430);
or U26853 (N_26853,N_26320,N_26099);
and U26854 (N_26854,N_26314,N_26039);
and U26855 (N_26855,N_26150,N_26015);
nand U26856 (N_26856,N_26279,N_26039);
nor U26857 (N_26857,N_26366,N_26342);
and U26858 (N_26858,N_26041,N_26457);
and U26859 (N_26859,N_26074,N_26227);
nor U26860 (N_26860,N_26044,N_26357);
nand U26861 (N_26861,N_26241,N_26476);
nor U26862 (N_26862,N_26019,N_26266);
xor U26863 (N_26863,N_26248,N_26219);
and U26864 (N_26864,N_26345,N_26008);
nor U26865 (N_26865,N_26270,N_26306);
nand U26866 (N_26866,N_26132,N_26386);
nand U26867 (N_26867,N_26413,N_26188);
xor U26868 (N_26868,N_26263,N_26009);
xnor U26869 (N_26869,N_26219,N_26291);
and U26870 (N_26870,N_26108,N_26499);
or U26871 (N_26871,N_26423,N_26421);
nand U26872 (N_26872,N_26138,N_26084);
nand U26873 (N_26873,N_26229,N_26137);
or U26874 (N_26874,N_26201,N_26098);
nand U26875 (N_26875,N_26270,N_26367);
nand U26876 (N_26876,N_26160,N_26083);
nor U26877 (N_26877,N_26422,N_26289);
nor U26878 (N_26878,N_26053,N_26313);
and U26879 (N_26879,N_26335,N_26279);
xnor U26880 (N_26880,N_26119,N_26339);
nand U26881 (N_26881,N_26244,N_26445);
xor U26882 (N_26882,N_26059,N_26310);
and U26883 (N_26883,N_26338,N_26343);
xnor U26884 (N_26884,N_26158,N_26190);
nand U26885 (N_26885,N_26063,N_26161);
nor U26886 (N_26886,N_26454,N_26102);
or U26887 (N_26887,N_26384,N_26460);
nor U26888 (N_26888,N_26187,N_26180);
xor U26889 (N_26889,N_26469,N_26397);
xnor U26890 (N_26890,N_26166,N_26199);
and U26891 (N_26891,N_26234,N_26045);
and U26892 (N_26892,N_26440,N_26201);
and U26893 (N_26893,N_26073,N_26259);
or U26894 (N_26894,N_26257,N_26190);
nand U26895 (N_26895,N_26417,N_26285);
xor U26896 (N_26896,N_26419,N_26174);
nand U26897 (N_26897,N_26366,N_26109);
nor U26898 (N_26898,N_26434,N_26288);
nor U26899 (N_26899,N_26252,N_26163);
nor U26900 (N_26900,N_26068,N_26173);
or U26901 (N_26901,N_26063,N_26110);
nor U26902 (N_26902,N_26134,N_26493);
and U26903 (N_26903,N_26045,N_26103);
or U26904 (N_26904,N_26045,N_26087);
and U26905 (N_26905,N_26046,N_26396);
nand U26906 (N_26906,N_26266,N_26027);
nand U26907 (N_26907,N_26408,N_26101);
xor U26908 (N_26908,N_26453,N_26188);
xnor U26909 (N_26909,N_26233,N_26461);
or U26910 (N_26910,N_26356,N_26408);
and U26911 (N_26911,N_26196,N_26492);
or U26912 (N_26912,N_26099,N_26178);
xor U26913 (N_26913,N_26034,N_26198);
or U26914 (N_26914,N_26380,N_26132);
nor U26915 (N_26915,N_26150,N_26228);
or U26916 (N_26916,N_26236,N_26477);
nand U26917 (N_26917,N_26401,N_26131);
and U26918 (N_26918,N_26472,N_26094);
nand U26919 (N_26919,N_26034,N_26267);
nor U26920 (N_26920,N_26375,N_26448);
nor U26921 (N_26921,N_26045,N_26448);
xnor U26922 (N_26922,N_26364,N_26060);
and U26923 (N_26923,N_26148,N_26167);
nand U26924 (N_26924,N_26384,N_26200);
nand U26925 (N_26925,N_26457,N_26284);
xnor U26926 (N_26926,N_26349,N_26444);
xor U26927 (N_26927,N_26010,N_26108);
or U26928 (N_26928,N_26291,N_26379);
nand U26929 (N_26929,N_26360,N_26426);
nand U26930 (N_26930,N_26011,N_26429);
xnor U26931 (N_26931,N_26194,N_26185);
or U26932 (N_26932,N_26363,N_26061);
nand U26933 (N_26933,N_26386,N_26482);
or U26934 (N_26934,N_26362,N_26266);
nor U26935 (N_26935,N_26417,N_26340);
xnor U26936 (N_26936,N_26008,N_26252);
nand U26937 (N_26937,N_26333,N_26264);
nor U26938 (N_26938,N_26172,N_26007);
and U26939 (N_26939,N_26148,N_26428);
nor U26940 (N_26940,N_26292,N_26360);
and U26941 (N_26941,N_26262,N_26046);
nand U26942 (N_26942,N_26129,N_26240);
nor U26943 (N_26943,N_26299,N_26252);
xor U26944 (N_26944,N_26175,N_26132);
xnor U26945 (N_26945,N_26353,N_26152);
nor U26946 (N_26946,N_26331,N_26316);
or U26947 (N_26947,N_26197,N_26494);
nor U26948 (N_26948,N_26071,N_26477);
or U26949 (N_26949,N_26203,N_26232);
xnor U26950 (N_26950,N_26032,N_26083);
and U26951 (N_26951,N_26389,N_26208);
nor U26952 (N_26952,N_26278,N_26303);
nand U26953 (N_26953,N_26327,N_26407);
nand U26954 (N_26954,N_26201,N_26410);
xor U26955 (N_26955,N_26471,N_26164);
or U26956 (N_26956,N_26308,N_26064);
or U26957 (N_26957,N_26322,N_26174);
or U26958 (N_26958,N_26390,N_26423);
xnor U26959 (N_26959,N_26395,N_26077);
xor U26960 (N_26960,N_26053,N_26069);
or U26961 (N_26961,N_26056,N_26279);
nor U26962 (N_26962,N_26149,N_26021);
or U26963 (N_26963,N_26273,N_26474);
xor U26964 (N_26964,N_26401,N_26099);
and U26965 (N_26965,N_26432,N_26124);
xor U26966 (N_26966,N_26131,N_26062);
nand U26967 (N_26967,N_26020,N_26122);
nor U26968 (N_26968,N_26328,N_26460);
nor U26969 (N_26969,N_26395,N_26032);
nand U26970 (N_26970,N_26350,N_26347);
nand U26971 (N_26971,N_26189,N_26109);
xor U26972 (N_26972,N_26031,N_26451);
and U26973 (N_26973,N_26339,N_26262);
or U26974 (N_26974,N_26226,N_26317);
or U26975 (N_26975,N_26211,N_26268);
and U26976 (N_26976,N_26161,N_26224);
and U26977 (N_26977,N_26478,N_26342);
or U26978 (N_26978,N_26261,N_26056);
or U26979 (N_26979,N_26091,N_26438);
nor U26980 (N_26980,N_26085,N_26089);
and U26981 (N_26981,N_26140,N_26205);
nand U26982 (N_26982,N_26463,N_26099);
or U26983 (N_26983,N_26360,N_26225);
or U26984 (N_26984,N_26468,N_26105);
xor U26985 (N_26985,N_26096,N_26363);
nand U26986 (N_26986,N_26494,N_26453);
xnor U26987 (N_26987,N_26425,N_26020);
and U26988 (N_26988,N_26391,N_26304);
and U26989 (N_26989,N_26007,N_26051);
and U26990 (N_26990,N_26092,N_26381);
nand U26991 (N_26991,N_26182,N_26020);
or U26992 (N_26992,N_26272,N_26016);
xnor U26993 (N_26993,N_26218,N_26490);
or U26994 (N_26994,N_26415,N_26270);
or U26995 (N_26995,N_26234,N_26442);
nor U26996 (N_26996,N_26301,N_26135);
nand U26997 (N_26997,N_26190,N_26420);
and U26998 (N_26998,N_26393,N_26230);
nand U26999 (N_26999,N_26075,N_26298);
or U27000 (N_27000,N_26639,N_26938);
nor U27001 (N_27001,N_26547,N_26595);
nand U27002 (N_27002,N_26799,N_26872);
nor U27003 (N_27003,N_26915,N_26786);
xnor U27004 (N_27004,N_26679,N_26979);
or U27005 (N_27005,N_26768,N_26849);
or U27006 (N_27006,N_26984,N_26845);
and U27007 (N_27007,N_26716,N_26956);
xor U27008 (N_27008,N_26589,N_26794);
nor U27009 (N_27009,N_26905,N_26505);
nor U27010 (N_27010,N_26687,N_26593);
or U27011 (N_27011,N_26896,N_26631);
nand U27012 (N_27012,N_26667,N_26583);
or U27013 (N_27013,N_26753,N_26556);
xor U27014 (N_27014,N_26777,N_26999);
nor U27015 (N_27015,N_26946,N_26611);
or U27016 (N_27016,N_26800,N_26507);
and U27017 (N_27017,N_26994,N_26742);
and U27018 (N_27018,N_26801,N_26871);
xor U27019 (N_27019,N_26617,N_26581);
xor U27020 (N_27020,N_26566,N_26628);
nand U27021 (N_27021,N_26763,N_26750);
or U27022 (N_27022,N_26823,N_26587);
nand U27023 (N_27023,N_26645,N_26541);
nand U27024 (N_27024,N_26525,N_26771);
nand U27025 (N_27025,N_26895,N_26726);
nand U27026 (N_27026,N_26598,N_26546);
nand U27027 (N_27027,N_26944,N_26676);
or U27028 (N_27028,N_26839,N_26736);
nand U27029 (N_27029,N_26898,N_26625);
or U27030 (N_27030,N_26666,N_26773);
nand U27031 (N_27031,N_26616,N_26684);
nand U27032 (N_27032,N_26803,N_26513);
or U27033 (N_27033,N_26521,N_26860);
xor U27034 (N_27034,N_26538,N_26685);
nor U27035 (N_27035,N_26699,N_26635);
and U27036 (N_27036,N_26772,N_26833);
or U27037 (N_27037,N_26958,N_26862);
and U27038 (N_27038,N_26535,N_26897);
nand U27039 (N_27039,N_26952,N_26634);
or U27040 (N_27040,N_26993,N_26848);
nor U27041 (N_27041,N_26718,N_26919);
xnor U27042 (N_27042,N_26602,N_26935);
or U27043 (N_27043,N_26814,N_26881);
or U27044 (N_27044,N_26606,N_26749);
nor U27045 (N_27045,N_26879,N_26551);
nor U27046 (N_27046,N_26618,N_26545);
or U27047 (N_27047,N_26534,N_26868);
or U27048 (N_27048,N_26623,N_26506);
nand U27049 (N_27049,N_26629,N_26561);
xnor U27050 (N_27050,N_26519,N_26990);
nand U27051 (N_27051,N_26955,N_26932);
xor U27052 (N_27052,N_26820,N_26605);
nand U27053 (N_27053,N_26909,N_26832);
and U27054 (N_27054,N_26882,N_26517);
xnor U27055 (N_27055,N_26853,N_26532);
nand U27056 (N_27056,N_26648,N_26758);
nor U27057 (N_27057,N_26592,N_26787);
or U27058 (N_27058,N_26904,N_26811);
or U27059 (N_27059,N_26885,N_26825);
xnor U27060 (N_27060,N_26664,N_26731);
nor U27061 (N_27061,N_26810,N_26789);
and U27062 (N_27062,N_26708,N_26981);
nor U27063 (N_27063,N_26913,N_26917);
nand U27064 (N_27064,N_26797,N_26805);
and U27065 (N_27065,N_26949,N_26908);
nand U27066 (N_27066,N_26527,N_26930);
and U27067 (N_27067,N_26796,N_26948);
nor U27068 (N_27068,N_26921,N_26533);
nor U27069 (N_27069,N_26992,N_26638);
nand U27070 (N_27070,N_26980,N_26696);
nor U27071 (N_27071,N_26876,N_26883);
xor U27072 (N_27072,N_26859,N_26830);
or U27073 (N_27073,N_26945,N_26609);
nor U27074 (N_27074,N_26614,N_26974);
and U27075 (N_27075,N_26580,N_26711);
nor U27076 (N_27076,N_26619,N_26636);
nor U27077 (N_27077,N_26514,N_26512);
or U27078 (N_27078,N_26572,N_26855);
or U27079 (N_27079,N_26858,N_26693);
nand U27080 (N_27080,N_26596,N_26567);
nand U27081 (N_27081,N_26933,N_26929);
nor U27082 (N_27082,N_26864,N_26704);
or U27083 (N_27083,N_26559,N_26548);
nor U27084 (N_27084,N_26809,N_26804);
or U27085 (N_27085,N_26986,N_26542);
nand U27086 (N_27086,N_26892,N_26788);
nor U27087 (N_27087,N_26818,N_26791);
xor U27088 (N_27088,N_26682,N_26727);
and U27089 (N_27089,N_26827,N_26874);
and U27090 (N_27090,N_26660,N_26694);
xor U27091 (N_27091,N_26709,N_26594);
nor U27092 (N_27092,N_26808,N_26508);
nand U27093 (N_27093,N_26515,N_26939);
nor U27094 (N_27094,N_26722,N_26637);
nor U27095 (N_27095,N_26813,N_26601);
or U27096 (N_27096,N_26672,N_26910);
or U27097 (N_27097,N_26558,N_26747);
nor U27098 (N_27098,N_26560,N_26900);
nand U27099 (N_27099,N_26738,N_26537);
or U27100 (N_27100,N_26653,N_26755);
or U27101 (N_27101,N_26931,N_26646);
and U27102 (N_27102,N_26942,N_26779);
nand U27103 (N_27103,N_26972,N_26838);
or U27104 (N_27104,N_26982,N_26651);
xnor U27105 (N_27105,N_26745,N_26522);
xnor U27106 (N_27106,N_26925,N_26783);
xor U27107 (N_27107,N_26654,N_26970);
or U27108 (N_27108,N_26914,N_26621);
nor U27109 (N_27109,N_26509,N_26826);
or U27110 (N_27110,N_26705,N_26698);
and U27111 (N_27111,N_26840,N_26540);
nand U27112 (N_27112,N_26903,N_26652);
nor U27113 (N_27113,N_26670,N_26675);
and U27114 (N_27114,N_26966,N_26843);
xnor U27115 (N_27115,N_26977,N_26700);
or U27116 (N_27116,N_26969,N_26888);
and U27117 (N_27117,N_26819,N_26995);
and U27118 (N_27118,N_26978,N_26630);
nor U27119 (N_27119,N_26543,N_26923);
and U27120 (N_27120,N_26615,N_26782);
xor U27121 (N_27121,N_26574,N_26756);
nor U27122 (N_27122,N_26626,N_26659);
and U27123 (N_27123,N_26907,N_26937);
xor U27124 (N_27124,N_26926,N_26766);
nor U27125 (N_27125,N_26816,N_26835);
and U27126 (N_27126,N_26683,N_26934);
or U27127 (N_27127,N_26585,N_26961);
nand U27128 (N_27128,N_26940,N_26856);
nand U27129 (N_27129,N_26590,N_26841);
nand U27130 (N_27130,N_26671,N_26837);
or U27131 (N_27131,N_26662,N_26578);
nor U27132 (N_27132,N_26656,N_26821);
nor U27133 (N_27133,N_26951,N_26962);
nand U27134 (N_27134,N_26889,N_26953);
xor U27135 (N_27135,N_26761,N_26922);
nor U27136 (N_27136,N_26706,N_26989);
xnor U27137 (N_27137,N_26746,N_26902);
or U27138 (N_27138,N_26744,N_26834);
and U27139 (N_27139,N_26529,N_26996);
or U27140 (N_27140,N_26557,N_26680);
xor U27141 (N_27141,N_26875,N_26957);
xor U27142 (N_27142,N_26918,N_26644);
and U27143 (N_27143,N_26586,N_26523);
or U27144 (N_27144,N_26715,N_26866);
or U27145 (N_27145,N_26959,N_26569);
and U27146 (N_27146,N_26734,N_26752);
and U27147 (N_27147,N_26649,N_26524);
nand U27148 (N_27148,N_26599,N_26516);
nand U27149 (N_27149,N_26751,N_26518);
xnor U27150 (N_27150,N_26668,N_26714);
or U27151 (N_27151,N_26658,N_26555);
xor U27152 (N_27152,N_26579,N_26985);
or U27153 (N_27153,N_26822,N_26719);
nor U27154 (N_27154,N_26988,N_26733);
xor U27155 (N_27155,N_26776,N_26703);
or U27156 (N_27156,N_26576,N_26728);
xor U27157 (N_27157,N_26760,N_26829);
and U27158 (N_27158,N_26790,N_26836);
and U27159 (N_27159,N_26530,N_26661);
nor U27160 (N_27160,N_26943,N_26911);
and U27161 (N_27161,N_26554,N_26947);
nand U27162 (N_27162,N_26565,N_26887);
nor U27163 (N_27163,N_26600,N_26681);
or U27164 (N_27164,N_26612,N_26991);
or U27165 (N_27165,N_26765,N_26591);
nor U27166 (N_27166,N_26552,N_26812);
and U27167 (N_27167,N_26998,N_26573);
nor U27168 (N_27168,N_26880,N_26500);
xnor U27169 (N_27169,N_26689,N_26575);
and U27170 (N_27170,N_26739,N_26778);
and U27171 (N_27171,N_26633,N_26971);
xor U27172 (N_27172,N_26987,N_26536);
nand U27173 (N_27173,N_26713,N_26607);
or U27174 (N_27174,N_26857,N_26824);
and U27175 (N_27175,N_26976,N_26865);
and U27176 (N_27176,N_26632,N_26526);
xnor U27177 (N_27177,N_26608,N_26690);
or U27178 (N_27178,N_26620,N_26544);
xnor U27179 (N_27179,N_26568,N_26807);
and U27180 (N_27180,N_26692,N_26828);
and U27181 (N_27181,N_26793,N_26725);
and U27182 (N_27182,N_26846,N_26964);
nand U27183 (N_27183,N_26870,N_26806);
xor U27184 (N_27184,N_26844,N_26759);
nor U27185 (N_27185,N_26960,N_26784);
nor U27186 (N_27186,N_26973,N_26798);
and U27187 (N_27187,N_26686,N_26924);
nand U27188 (N_27188,N_26894,N_26588);
nand U27189 (N_27189,N_26732,N_26702);
nand U27190 (N_27190,N_26674,N_26622);
nand U27191 (N_27191,N_26564,N_26710);
xor U27192 (N_27192,N_26877,N_26640);
xor U27193 (N_27193,N_26737,N_26701);
and U27194 (N_27194,N_26717,N_26663);
and U27195 (N_27195,N_26669,N_26764);
nor U27196 (N_27196,N_26886,N_26603);
or U27197 (N_27197,N_26582,N_26531);
and U27198 (N_27198,N_26740,N_26539);
xnor U27199 (N_27199,N_26642,N_26743);
xor U27200 (N_27200,N_26968,N_26785);
xor U27201 (N_27201,N_26920,N_26624);
nand U27202 (N_27202,N_26780,N_26950);
nor U27203 (N_27203,N_26965,N_26678);
xor U27204 (N_27204,N_26748,N_26815);
nor U27205 (N_27205,N_26847,N_26975);
nand U27206 (N_27206,N_26503,N_26650);
or U27207 (N_27207,N_26899,N_26712);
xor U27208 (N_27208,N_26842,N_26802);
and U27209 (N_27209,N_26720,N_26673);
nor U27210 (N_27210,N_26584,N_26647);
nand U27211 (N_27211,N_26610,N_26997);
nand U27212 (N_27212,N_26511,N_26549);
or U27213 (N_27213,N_26854,N_26571);
nor U27214 (N_27214,N_26707,N_26502);
nor U27215 (N_27215,N_26657,N_26691);
nor U27216 (N_27216,N_26852,N_26873);
and U27217 (N_27217,N_26963,N_26901);
and U27218 (N_27218,N_26695,N_26643);
or U27219 (N_27219,N_26863,N_26928);
nor U27220 (N_27220,N_26562,N_26604);
or U27221 (N_27221,N_26884,N_26735);
nand U27222 (N_27222,N_26831,N_26641);
or U27223 (N_27223,N_26677,N_26665);
xor U27224 (N_27224,N_26520,N_26553);
nand U27225 (N_27225,N_26954,N_26906);
nor U27226 (N_27226,N_26869,N_26817);
nor U27227 (N_27227,N_26781,N_26501);
and U27228 (N_27228,N_26767,N_26510);
and U27229 (N_27229,N_26570,N_26613);
nor U27230 (N_27230,N_26721,N_26770);
and U27231 (N_27231,N_26577,N_26697);
or U27232 (N_27232,N_26891,N_26850);
xor U27233 (N_27233,N_26878,N_26775);
and U27234 (N_27234,N_26757,N_26550);
nor U27235 (N_27235,N_26741,N_26528);
nand U27236 (N_27236,N_26936,N_26688);
nand U27237 (N_27237,N_26627,N_26867);
and U27238 (N_27238,N_26851,N_26916);
nand U27239 (N_27239,N_26724,N_26861);
xor U27240 (N_27240,N_26504,N_26729);
xnor U27241 (N_27241,N_26730,N_26983);
and U27242 (N_27242,N_26792,N_26795);
nand U27243 (N_27243,N_26754,N_26893);
nor U27244 (N_27244,N_26597,N_26774);
nor U27245 (N_27245,N_26563,N_26927);
or U27246 (N_27246,N_26967,N_26941);
nor U27247 (N_27247,N_26655,N_26723);
xor U27248 (N_27248,N_26912,N_26769);
or U27249 (N_27249,N_26762,N_26890);
nor U27250 (N_27250,N_26544,N_26910);
nand U27251 (N_27251,N_26661,N_26799);
and U27252 (N_27252,N_26951,N_26544);
and U27253 (N_27253,N_26602,N_26810);
nor U27254 (N_27254,N_26764,N_26555);
nor U27255 (N_27255,N_26547,N_26577);
nor U27256 (N_27256,N_26845,N_26733);
xor U27257 (N_27257,N_26592,N_26970);
nor U27258 (N_27258,N_26984,N_26745);
xnor U27259 (N_27259,N_26995,N_26949);
or U27260 (N_27260,N_26529,N_26993);
nor U27261 (N_27261,N_26713,N_26909);
or U27262 (N_27262,N_26886,N_26915);
or U27263 (N_27263,N_26896,N_26628);
xnor U27264 (N_27264,N_26594,N_26597);
and U27265 (N_27265,N_26796,N_26727);
nand U27266 (N_27266,N_26922,N_26738);
nor U27267 (N_27267,N_26610,N_26559);
xnor U27268 (N_27268,N_26617,N_26590);
and U27269 (N_27269,N_26641,N_26967);
nor U27270 (N_27270,N_26973,N_26943);
nor U27271 (N_27271,N_26886,N_26727);
nand U27272 (N_27272,N_26983,N_26950);
nor U27273 (N_27273,N_26731,N_26604);
or U27274 (N_27274,N_26812,N_26965);
or U27275 (N_27275,N_26824,N_26845);
nor U27276 (N_27276,N_26956,N_26666);
nand U27277 (N_27277,N_26781,N_26913);
nor U27278 (N_27278,N_26788,N_26546);
and U27279 (N_27279,N_26967,N_26554);
nand U27280 (N_27280,N_26957,N_26836);
xnor U27281 (N_27281,N_26941,N_26772);
nor U27282 (N_27282,N_26795,N_26713);
nor U27283 (N_27283,N_26636,N_26951);
nand U27284 (N_27284,N_26553,N_26918);
xor U27285 (N_27285,N_26859,N_26750);
nand U27286 (N_27286,N_26937,N_26672);
nor U27287 (N_27287,N_26902,N_26732);
and U27288 (N_27288,N_26791,N_26785);
nand U27289 (N_27289,N_26918,N_26878);
or U27290 (N_27290,N_26873,N_26652);
nand U27291 (N_27291,N_26828,N_26560);
nand U27292 (N_27292,N_26708,N_26531);
or U27293 (N_27293,N_26922,N_26567);
nor U27294 (N_27294,N_26618,N_26557);
or U27295 (N_27295,N_26897,N_26984);
and U27296 (N_27296,N_26743,N_26980);
or U27297 (N_27297,N_26564,N_26864);
nor U27298 (N_27298,N_26968,N_26588);
and U27299 (N_27299,N_26802,N_26962);
nand U27300 (N_27300,N_26974,N_26538);
nand U27301 (N_27301,N_26930,N_26837);
and U27302 (N_27302,N_26757,N_26679);
and U27303 (N_27303,N_26755,N_26569);
or U27304 (N_27304,N_26730,N_26544);
xor U27305 (N_27305,N_26644,N_26910);
nor U27306 (N_27306,N_26863,N_26802);
nand U27307 (N_27307,N_26898,N_26751);
nand U27308 (N_27308,N_26738,N_26801);
nand U27309 (N_27309,N_26571,N_26917);
nand U27310 (N_27310,N_26769,N_26807);
nand U27311 (N_27311,N_26748,N_26751);
nand U27312 (N_27312,N_26588,N_26607);
or U27313 (N_27313,N_26660,N_26689);
or U27314 (N_27314,N_26617,N_26722);
nand U27315 (N_27315,N_26549,N_26838);
nor U27316 (N_27316,N_26697,N_26789);
nand U27317 (N_27317,N_26661,N_26787);
nand U27318 (N_27318,N_26504,N_26717);
or U27319 (N_27319,N_26883,N_26800);
nand U27320 (N_27320,N_26507,N_26819);
nand U27321 (N_27321,N_26896,N_26888);
nand U27322 (N_27322,N_26911,N_26780);
or U27323 (N_27323,N_26797,N_26848);
nor U27324 (N_27324,N_26564,N_26578);
xor U27325 (N_27325,N_26893,N_26765);
and U27326 (N_27326,N_26879,N_26712);
and U27327 (N_27327,N_26755,N_26890);
or U27328 (N_27328,N_26517,N_26690);
nand U27329 (N_27329,N_26598,N_26592);
nor U27330 (N_27330,N_26948,N_26984);
xnor U27331 (N_27331,N_26545,N_26522);
xor U27332 (N_27332,N_26511,N_26695);
and U27333 (N_27333,N_26973,N_26823);
and U27334 (N_27334,N_26687,N_26969);
nand U27335 (N_27335,N_26676,N_26724);
or U27336 (N_27336,N_26694,N_26904);
and U27337 (N_27337,N_26636,N_26747);
and U27338 (N_27338,N_26782,N_26889);
or U27339 (N_27339,N_26953,N_26635);
or U27340 (N_27340,N_26595,N_26605);
or U27341 (N_27341,N_26864,N_26681);
xor U27342 (N_27342,N_26591,N_26707);
or U27343 (N_27343,N_26591,N_26697);
xor U27344 (N_27344,N_26620,N_26727);
nand U27345 (N_27345,N_26925,N_26602);
nor U27346 (N_27346,N_26637,N_26983);
nor U27347 (N_27347,N_26637,N_26941);
xnor U27348 (N_27348,N_26615,N_26797);
nor U27349 (N_27349,N_26837,N_26749);
nor U27350 (N_27350,N_26801,N_26817);
and U27351 (N_27351,N_26867,N_26681);
nand U27352 (N_27352,N_26936,N_26971);
and U27353 (N_27353,N_26941,N_26940);
or U27354 (N_27354,N_26849,N_26798);
nand U27355 (N_27355,N_26981,N_26818);
nor U27356 (N_27356,N_26979,N_26761);
or U27357 (N_27357,N_26761,N_26950);
nand U27358 (N_27358,N_26598,N_26905);
nand U27359 (N_27359,N_26873,N_26965);
nor U27360 (N_27360,N_26992,N_26500);
xor U27361 (N_27361,N_26897,N_26539);
nor U27362 (N_27362,N_26855,N_26838);
or U27363 (N_27363,N_26590,N_26615);
xnor U27364 (N_27364,N_26752,N_26826);
nand U27365 (N_27365,N_26606,N_26623);
xnor U27366 (N_27366,N_26516,N_26659);
nand U27367 (N_27367,N_26953,N_26982);
xor U27368 (N_27368,N_26533,N_26992);
xnor U27369 (N_27369,N_26664,N_26986);
and U27370 (N_27370,N_26901,N_26604);
or U27371 (N_27371,N_26991,N_26516);
nand U27372 (N_27372,N_26507,N_26568);
or U27373 (N_27373,N_26793,N_26937);
nor U27374 (N_27374,N_26864,N_26970);
or U27375 (N_27375,N_26739,N_26562);
or U27376 (N_27376,N_26952,N_26845);
xor U27377 (N_27377,N_26508,N_26851);
xnor U27378 (N_27378,N_26795,N_26977);
xor U27379 (N_27379,N_26790,N_26882);
nand U27380 (N_27380,N_26710,N_26764);
nor U27381 (N_27381,N_26640,N_26847);
xor U27382 (N_27382,N_26811,N_26625);
or U27383 (N_27383,N_26959,N_26533);
nand U27384 (N_27384,N_26975,N_26716);
nor U27385 (N_27385,N_26720,N_26504);
and U27386 (N_27386,N_26659,N_26664);
xor U27387 (N_27387,N_26879,N_26717);
nor U27388 (N_27388,N_26638,N_26760);
or U27389 (N_27389,N_26709,N_26808);
or U27390 (N_27390,N_26813,N_26742);
nor U27391 (N_27391,N_26875,N_26717);
or U27392 (N_27392,N_26882,N_26636);
nand U27393 (N_27393,N_26609,N_26591);
or U27394 (N_27394,N_26766,N_26619);
and U27395 (N_27395,N_26793,N_26524);
nor U27396 (N_27396,N_26872,N_26502);
nand U27397 (N_27397,N_26599,N_26523);
and U27398 (N_27398,N_26944,N_26823);
or U27399 (N_27399,N_26603,N_26928);
nand U27400 (N_27400,N_26732,N_26673);
and U27401 (N_27401,N_26835,N_26849);
xor U27402 (N_27402,N_26999,N_26625);
nand U27403 (N_27403,N_26842,N_26542);
nor U27404 (N_27404,N_26544,N_26698);
nand U27405 (N_27405,N_26585,N_26659);
nand U27406 (N_27406,N_26960,N_26799);
nand U27407 (N_27407,N_26646,N_26633);
xor U27408 (N_27408,N_26803,N_26615);
nor U27409 (N_27409,N_26753,N_26713);
or U27410 (N_27410,N_26972,N_26730);
and U27411 (N_27411,N_26946,N_26730);
and U27412 (N_27412,N_26626,N_26670);
nand U27413 (N_27413,N_26802,N_26688);
nor U27414 (N_27414,N_26591,N_26778);
and U27415 (N_27415,N_26680,N_26590);
xnor U27416 (N_27416,N_26586,N_26629);
or U27417 (N_27417,N_26873,N_26670);
nand U27418 (N_27418,N_26550,N_26914);
nand U27419 (N_27419,N_26578,N_26685);
nor U27420 (N_27420,N_26628,N_26798);
and U27421 (N_27421,N_26936,N_26885);
nand U27422 (N_27422,N_26503,N_26838);
nor U27423 (N_27423,N_26865,N_26906);
and U27424 (N_27424,N_26753,N_26983);
xnor U27425 (N_27425,N_26622,N_26611);
and U27426 (N_27426,N_26962,N_26729);
or U27427 (N_27427,N_26945,N_26933);
nor U27428 (N_27428,N_26990,N_26661);
nor U27429 (N_27429,N_26805,N_26808);
nand U27430 (N_27430,N_26660,N_26960);
and U27431 (N_27431,N_26758,N_26849);
xor U27432 (N_27432,N_26887,N_26652);
or U27433 (N_27433,N_26539,N_26552);
nor U27434 (N_27434,N_26825,N_26644);
xnor U27435 (N_27435,N_26535,N_26793);
xor U27436 (N_27436,N_26696,N_26941);
nor U27437 (N_27437,N_26580,N_26672);
xor U27438 (N_27438,N_26881,N_26952);
nor U27439 (N_27439,N_26572,N_26797);
nor U27440 (N_27440,N_26878,N_26581);
xnor U27441 (N_27441,N_26759,N_26850);
nand U27442 (N_27442,N_26698,N_26617);
xor U27443 (N_27443,N_26859,N_26749);
nand U27444 (N_27444,N_26581,N_26883);
and U27445 (N_27445,N_26638,N_26776);
nor U27446 (N_27446,N_26636,N_26729);
and U27447 (N_27447,N_26776,N_26772);
nand U27448 (N_27448,N_26567,N_26907);
xor U27449 (N_27449,N_26941,N_26869);
or U27450 (N_27450,N_26954,N_26566);
or U27451 (N_27451,N_26956,N_26785);
or U27452 (N_27452,N_26661,N_26591);
nor U27453 (N_27453,N_26721,N_26728);
nor U27454 (N_27454,N_26855,N_26600);
nor U27455 (N_27455,N_26723,N_26764);
nand U27456 (N_27456,N_26704,N_26665);
nor U27457 (N_27457,N_26988,N_26876);
xnor U27458 (N_27458,N_26930,N_26554);
nor U27459 (N_27459,N_26881,N_26669);
xor U27460 (N_27460,N_26708,N_26866);
or U27461 (N_27461,N_26723,N_26641);
nand U27462 (N_27462,N_26707,N_26578);
xor U27463 (N_27463,N_26517,N_26724);
and U27464 (N_27464,N_26867,N_26944);
or U27465 (N_27465,N_26818,N_26597);
nand U27466 (N_27466,N_26510,N_26829);
nor U27467 (N_27467,N_26809,N_26511);
xnor U27468 (N_27468,N_26719,N_26647);
or U27469 (N_27469,N_26973,N_26965);
or U27470 (N_27470,N_26794,N_26553);
nor U27471 (N_27471,N_26826,N_26788);
nor U27472 (N_27472,N_26801,N_26564);
nand U27473 (N_27473,N_26636,N_26924);
nor U27474 (N_27474,N_26511,N_26538);
nand U27475 (N_27475,N_26653,N_26513);
xnor U27476 (N_27476,N_26834,N_26937);
and U27477 (N_27477,N_26885,N_26792);
nor U27478 (N_27478,N_26678,N_26707);
nand U27479 (N_27479,N_26629,N_26829);
and U27480 (N_27480,N_26555,N_26749);
nor U27481 (N_27481,N_26795,N_26872);
xnor U27482 (N_27482,N_26937,N_26566);
nand U27483 (N_27483,N_26551,N_26680);
xnor U27484 (N_27484,N_26849,N_26847);
nand U27485 (N_27485,N_26700,N_26514);
xor U27486 (N_27486,N_26507,N_26523);
nor U27487 (N_27487,N_26546,N_26714);
nor U27488 (N_27488,N_26962,N_26608);
and U27489 (N_27489,N_26850,N_26544);
or U27490 (N_27490,N_26858,N_26919);
nor U27491 (N_27491,N_26811,N_26798);
nand U27492 (N_27492,N_26921,N_26866);
nand U27493 (N_27493,N_26862,N_26691);
or U27494 (N_27494,N_26747,N_26801);
and U27495 (N_27495,N_26909,N_26739);
and U27496 (N_27496,N_26956,N_26829);
nor U27497 (N_27497,N_26963,N_26835);
or U27498 (N_27498,N_26553,N_26910);
nor U27499 (N_27499,N_26997,N_26773);
nand U27500 (N_27500,N_27147,N_27109);
xnor U27501 (N_27501,N_27234,N_27061);
or U27502 (N_27502,N_27418,N_27226);
xnor U27503 (N_27503,N_27427,N_27272);
nor U27504 (N_27504,N_27192,N_27123);
nand U27505 (N_27505,N_27170,N_27454);
xor U27506 (N_27506,N_27166,N_27012);
nand U27507 (N_27507,N_27080,N_27283);
and U27508 (N_27508,N_27139,N_27494);
xnor U27509 (N_27509,N_27342,N_27303);
and U27510 (N_27510,N_27372,N_27230);
or U27511 (N_27511,N_27047,N_27261);
xnor U27512 (N_27512,N_27287,N_27370);
or U27513 (N_27513,N_27135,N_27193);
and U27514 (N_27514,N_27441,N_27207);
xor U27515 (N_27515,N_27020,N_27463);
nand U27516 (N_27516,N_27247,N_27296);
xor U27517 (N_27517,N_27264,N_27255);
nand U27518 (N_27518,N_27155,N_27411);
nor U27519 (N_27519,N_27112,N_27348);
xnor U27520 (N_27520,N_27071,N_27163);
nor U27521 (N_27521,N_27154,N_27110);
nand U27522 (N_27522,N_27239,N_27381);
xnor U27523 (N_27523,N_27251,N_27040);
or U27524 (N_27524,N_27467,N_27334);
nor U27525 (N_27525,N_27305,N_27027);
nor U27526 (N_27526,N_27329,N_27295);
nand U27527 (N_27527,N_27219,N_27006);
and U27528 (N_27528,N_27188,N_27113);
or U27529 (N_27529,N_27439,N_27216);
xnor U27530 (N_27530,N_27438,N_27033);
xnor U27531 (N_27531,N_27351,N_27285);
nand U27532 (N_27532,N_27457,N_27086);
and U27533 (N_27533,N_27298,N_27346);
nand U27534 (N_27534,N_27314,N_27249);
and U27535 (N_27535,N_27489,N_27477);
or U27536 (N_27536,N_27194,N_27294);
and U27537 (N_27537,N_27099,N_27140);
nor U27538 (N_27538,N_27082,N_27420);
nand U27539 (N_27539,N_27374,N_27366);
and U27540 (N_27540,N_27365,N_27018);
or U27541 (N_27541,N_27383,N_27380);
or U27542 (N_27542,N_27256,N_27393);
xnor U27543 (N_27543,N_27078,N_27354);
or U27544 (N_27544,N_27324,N_27440);
or U27545 (N_27545,N_27395,N_27468);
and U27546 (N_27546,N_27036,N_27406);
xor U27547 (N_27547,N_27311,N_27414);
nor U27548 (N_27548,N_27423,N_27446);
nand U27549 (N_27549,N_27300,N_27394);
nand U27550 (N_27550,N_27054,N_27160);
or U27551 (N_27551,N_27369,N_27431);
nand U27552 (N_27552,N_27461,N_27279);
and U27553 (N_27553,N_27382,N_27146);
xor U27554 (N_27554,N_27421,N_27055);
nor U27555 (N_27555,N_27385,N_27217);
nor U27556 (N_27556,N_27443,N_27399);
or U27557 (N_27557,N_27100,N_27465);
and U27558 (N_27558,N_27043,N_27085);
nor U27559 (N_27559,N_27072,N_27453);
or U27560 (N_27560,N_27073,N_27191);
or U27561 (N_27561,N_27321,N_27144);
xor U27562 (N_27562,N_27211,N_27037);
and U27563 (N_27563,N_27108,N_27297);
xor U27564 (N_27564,N_27093,N_27433);
nor U27565 (N_27565,N_27445,N_27464);
or U27566 (N_27566,N_27025,N_27143);
nand U27567 (N_27567,N_27102,N_27499);
and U27568 (N_27568,N_27153,N_27031);
or U27569 (N_27569,N_27125,N_27103);
or U27570 (N_27570,N_27315,N_27128);
and U27571 (N_27571,N_27435,N_27200);
xnor U27572 (N_27572,N_27456,N_27046);
nand U27573 (N_27573,N_27316,N_27208);
or U27574 (N_27574,N_27024,N_27449);
and U27575 (N_27575,N_27032,N_27437);
or U27576 (N_27576,N_27087,N_27097);
or U27577 (N_27577,N_27023,N_27487);
and U27578 (N_27578,N_27238,N_27084);
and U27579 (N_27579,N_27229,N_27044);
or U27580 (N_27580,N_27232,N_27042);
xnor U27581 (N_27581,N_27426,N_27083);
nor U27582 (N_27582,N_27386,N_27246);
and U27583 (N_27583,N_27330,N_27403);
nor U27584 (N_27584,N_27245,N_27258);
and U27585 (N_27585,N_27045,N_27126);
or U27586 (N_27586,N_27002,N_27428);
nand U27587 (N_27587,N_27384,N_27336);
nor U27588 (N_27588,N_27168,N_27145);
nand U27589 (N_27589,N_27471,N_27377);
and U27590 (N_27590,N_27352,N_27114);
xor U27591 (N_27591,N_27187,N_27225);
nor U27592 (N_27592,N_27243,N_27323);
nor U27593 (N_27593,N_27450,N_27360);
and U27594 (N_27594,N_27274,N_27172);
nor U27595 (N_27595,N_27302,N_27095);
and U27596 (N_27596,N_27379,N_27017);
or U27597 (N_27597,N_27290,N_27179);
nor U27598 (N_27598,N_27409,N_27201);
or U27599 (N_27599,N_27176,N_27356);
nor U27600 (N_27600,N_27057,N_27396);
and U27601 (N_27601,N_27028,N_27149);
xor U27602 (N_27602,N_27318,N_27419);
nand U27603 (N_27603,N_27488,N_27292);
nand U27604 (N_27604,N_27313,N_27310);
nor U27605 (N_27605,N_27479,N_27483);
xor U27606 (N_27606,N_27069,N_27304);
nor U27607 (N_27607,N_27412,N_27401);
and U27608 (N_27608,N_27118,N_27052);
nand U27609 (N_27609,N_27391,N_27417);
nor U27610 (N_27610,N_27429,N_27432);
or U27611 (N_27611,N_27184,N_27011);
xor U27612 (N_27612,N_27138,N_27010);
and U27613 (N_27613,N_27280,N_27000);
xnor U27614 (N_27614,N_27130,N_27266);
nor U27615 (N_27615,N_27241,N_27121);
nor U27616 (N_27616,N_27325,N_27152);
nand U27617 (N_27617,N_27485,N_27227);
nor U27618 (N_27618,N_27021,N_27157);
nand U27619 (N_27619,N_27065,N_27268);
or U27620 (N_27620,N_27008,N_27240);
and U27621 (N_27621,N_27462,N_27344);
nor U27622 (N_27622,N_27415,N_27473);
xnor U27623 (N_27623,N_27224,N_27062);
nor U27624 (N_27624,N_27016,N_27094);
nor U27625 (N_27625,N_27452,N_27480);
xnor U27626 (N_27626,N_27349,N_27425);
or U27627 (N_27627,N_27408,N_27066);
nor U27628 (N_27628,N_27376,N_27068);
nand U27629 (N_27629,N_27362,N_27368);
nand U27630 (N_27630,N_27291,N_27159);
or U27631 (N_27631,N_27048,N_27286);
or U27632 (N_27632,N_27288,N_27339);
xor U27633 (N_27633,N_27206,N_27129);
nor U27634 (N_27634,N_27358,N_27004);
xor U27635 (N_27635,N_27252,N_27469);
nand U27636 (N_27636,N_27183,N_27470);
or U27637 (N_27637,N_27038,N_27132);
nand U27638 (N_27638,N_27448,N_27174);
nor U27639 (N_27639,N_27150,N_27478);
nand U27640 (N_27640,N_27177,N_27030);
nor U27641 (N_27641,N_27398,N_27116);
and U27642 (N_27642,N_27375,N_27253);
nand U27643 (N_27643,N_27332,N_27492);
nor U27644 (N_27644,N_27293,N_27106);
or U27645 (N_27645,N_27034,N_27156);
nand U27646 (N_27646,N_27067,N_27273);
nor U27647 (N_27647,N_27436,N_27079);
nor U27648 (N_27648,N_27387,N_27019);
nand U27649 (N_27649,N_27289,N_27322);
and U27650 (N_27650,N_27039,N_27111);
or U27651 (N_27651,N_27064,N_27338);
nor U27652 (N_27652,N_27136,N_27430);
and U27653 (N_27653,N_27141,N_27361);
nand U27654 (N_27654,N_27026,N_27378);
and U27655 (N_27655,N_27312,N_27058);
nand U27656 (N_27656,N_27005,N_27131);
xor U27657 (N_27657,N_27204,N_27257);
xor U27658 (N_27658,N_27231,N_27444);
or U27659 (N_27659,N_27271,N_27001);
and U27660 (N_27660,N_27220,N_27307);
or U27661 (N_27661,N_27096,N_27405);
nand U27662 (N_27662,N_27148,N_27390);
xor U27663 (N_27663,N_27355,N_27049);
and U27664 (N_27664,N_27169,N_27333);
and U27665 (N_27665,N_27015,N_27388);
nand U27666 (N_27666,N_27053,N_27215);
and U27667 (N_27667,N_27422,N_27205);
nor U27668 (N_27668,N_27284,N_27178);
nor U27669 (N_27669,N_27308,N_27331);
xor U27670 (N_27670,N_27014,N_27203);
or U27671 (N_27671,N_27345,N_27434);
or U27672 (N_27672,N_27413,N_27173);
and U27673 (N_27673,N_27495,N_27063);
and U27674 (N_27674,N_27481,N_27490);
nor U27675 (N_27675,N_27107,N_27190);
and U27676 (N_27676,N_27022,N_27282);
nor U27677 (N_27677,N_27142,N_27185);
nand U27678 (N_27678,N_27363,N_27496);
or U27679 (N_27679,N_27357,N_27459);
nand U27680 (N_27680,N_27309,N_27407);
or U27681 (N_27681,N_27041,N_27262);
and U27682 (N_27682,N_27158,N_27035);
nand U27683 (N_27683,N_27392,N_27077);
or U27684 (N_27684,N_27180,N_27353);
nor U27685 (N_27685,N_27250,N_27197);
and U27686 (N_27686,N_27416,N_27088);
and U27687 (N_27687,N_27267,N_27167);
nor U27688 (N_27688,N_27076,N_27491);
xnor U27689 (N_27689,N_27460,N_27402);
or U27690 (N_27690,N_27242,N_27127);
nand U27691 (N_27691,N_27104,N_27451);
or U27692 (N_27692,N_27013,N_27320);
xor U27693 (N_27693,N_27214,N_27081);
or U27694 (N_27694,N_27228,N_27341);
and U27695 (N_27695,N_27455,N_27359);
or U27696 (N_27696,N_27181,N_27458);
and U27697 (N_27697,N_27115,N_27189);
and U27698 (N_27698,N_27447,N_27400);
xor U27699 (N_27699,N_27209,N_27367);
nand U27700 (N_27700,N_27105,N_27003);
nand U27701 (N_27701,N_27474,N_27498);
or U27702 (N_27702,N_27133,N_27404);
and U27703 (N_27703,N_27328,N_27486);
or U27704 (N_27704,N_27410,N_27196);
nand U27705 (N_27705,N_27007,N_27056);
nand U27706 (N_27706,N_27171,N_27212);
xnor U27707 (N_27707,N_27319,N_27497);
and U27708 (N_27708,N_27326,N_27233);
or U27709 (N_27709,N_27424,N_27472);
nand U27710 (N_27710,N_27151,N_27340);
xor U27711 (N_27711,N_27074,N_27335);
nor U27712 (N_27712,N_27124,N_27343);
and U27713 (N_27713,N_27122,N_27260);
and U27714 (N_27714,N_27221,N_27223);
nand U27715 (N_27715,N_27092,N_27198);
nand U27716 (N_27716,N_27210,N_27161);
and U27717 (N_27717,N_27186,N_27244);
or U27718 (N_27718,N_27484,N_27199);
or U27719 (N_27719,N_27029,N_27098);
nand U27720 (N_27720,N_27218,N_27275);
xnor U27721 (N_27721,N_27134,N_27164);
or U27722 (N_27722,N_27350,N_27270);
xor U27723 (N_27723,N_27301,N_27306);
or U27724 (N_27724,N_27337,N_27259);
nand U27725 (N_27725,N_27269,N_27009);
xor U27726 (N_27726,N_27051,N_27070);
nor U27727 (N_27727,N_27397,N_27075);
or U27728 (N_27728,N_27119,N_27120);
nor U27729 (N_27729,N_27182,N_27442);
xnor U27730 (N_27730,N_27248,N_27089);
nor U27731 (N_27731,N_27327,N_27137);
and U27732 (N_27732,N_27165,N_27278);
xor U27733 (N_27733,N_27299,N_27213);
and U27734 (N_27734,N_27101,N_27263);
nor U27735 (N_27735,N_27475,N_27493);
xor U27736 (N_27736,N_27281,N_27050);
and U27737 (N_27737,N_27060,N_27117);
nand U27738 (N_27738,N_27276,N_27090);
nand U27739 (N_27739,N_27222,N_27236);
and U27740 (N_27740,N_27237,N_27175);
or U27741 (N_27741,N_27364,N_27389);
and U27742 (N_27742,N_27277,N_27162);
and U27743 (N_27743,N_27466,N_27235);
nor U27744 (N_27744,N_27482,N_27371);
or U27745 (N_27745,N_27317,N_27091);
or U27746 (N_27746,N_27059,N_27265);
and U27747 (N_27747,N_27347,N_27202);
nor U27748 (N_27748,N_27254,N_27476);
or U27749 (N_27749,N_27373,N_27195);
nand U27750 (N_27750,N_27047,N_27160);
or U27751 (N_27751,N_27179,N_27029);
nand U27752 (N_27752,N_27424,N_27099);
xor U27753 (N_27753,N_27361,N_27493);
nand U27754 (N_27754,N_27287,N_27383);
nor U27755 (N_27755,N_27005,N_27099);
xnor U27756 (N_27756,N_27215,N_27288);
and U27757 (N_27757,N_27294,N_27196);
nor U27758 (N_27758,N_27327,N_27211);
nor U27759 (N_27759,N_27163,N_27332);
nor U27760 (N_27760,N_27343,N_27465);
and U27761 (N_27761,N_27191,N_27441);
or U27762 (N_27762,N_27217,N_27111);
nor U27763 (N_27763,N_27116,N_27043);
xnor U27764 (N_27764,N_27121,N_27467);
and U27765 (N_27765,N_27076,N_27384);
and U27766 (N_27766,N_27212,N_27123);
and U27767 (N_27767,N_27239,N_27244);
nand U27768 (N_27768,N_27315,N_27150);
and U27769 (N_27769,N_27357,N_27319);
or U27770 (N_27770,N_27021,N_27353);
and U27771 (N_27771,N_27483,N_27359);
or U27772 (N_27772,N_27304,N_27038);
xor U27773 (N_27773,N_27328,N_27109);
and U27774 (N_27774,N_27013,N_27111);
nand U27775 (N_27775,N_27343,N_27295);
nand U27776 (N_27776,N_27272,N_27474);
xnor U27777 (N_27777,N_27114,N_27031);
xor U27778 (N_27778,N_27241,N_27250);
and U27779 (N_27779,N_27163,N_27135);
nand U27780 (N_27780,N_27143,N_27392);
xor U27781 (N_27781,N_27147,N_27072);
nand U27782 (N_27782,N_27358,N_27096);
or U27783 (N_27783,N_27487,N_27365);
and U27784 (N_27784,N_27062,N_27496);
or U27785 (N_27785,N_27359,N_27339);
or U27786 (N_27786,N_27459,N_27237);
nor U27787 (N_27787,N_27330,N_27281);
xnor U27788 (N_27788,N_27098,N_27069);
xor U27789 (N_27789,N_27498,N_27382);
nor U27790 (N_27790,N_27457,N_27280);
nand U27791 (N_27791,N_27143,N_27093);
xor U27792 (N_27792,N_27124,N_27070);
xor U27793 (N_27793,N_27248,N_27279);
and U27794 (N_27794,N_27497,N_27453);
xor U27795 (N_27795,N_27390,N_27277);
or U27796 (N_27796,N_27307,N_27209);
or U27797 (N_27797,N_27096,N_27344);
xnor U27798 (N_27798,N_27139,N_27192);
nand U27799 (N_27799,N_27144,N_27111);
nand U27800 (N_27800,N_27217,N_27386);
nand U27801 (N_27801,N_27009,N_27370);
or U27802 (N_27802,N_27382,N_27024);
or U27803 (N_27803,N_27361,N_27459);
or U27804 (N_27804,N_27456,N_27201);
or U27805 (N_27805,N_27016,N_27259);
or U27806 (N_27806,N_27488,N_27106);
or U27807 (N_27807,N_27476,N_27058);
and U27808 (N_27808,N_27080,N_27129);
nor U27809 (N_27809,N_27108,N_27417);
nand U27810 (N_27810,N_27113,N_27436);
nor U27811 (N_27811,N_27332,N_27189);
and U27812 (N_27812,N_27015,N_27330);
and U27813 (N_27813,N_27053,N_27236);
xor U27814 (N_27814,N_27307,N_27265);
nor U27815 (N_27815,N_27000,N_27279);
xnor U27816 (N_27816,N_27045,N_27344);
and U27817 (N_27817,N_27313,N_27234);
nand U27818 (N_27818,N_27252,N_27093);
nor U27819 (N_27819,N_27193,N_27419);
and U27820 (N_27820,N_27081,N_27264);
nor U27821 (N_27821,N_27265,N_27167);
and U27822 (N_27822,N_27171,N_27075);
xor U27823 (N_27823,N_27302,N_27328);
xor U27824 (N_27824,N_27159,N_27149);
nand U27825 (N_27825,N_27162,N_27497);
or U27826 (N_27826,N_27441,N_27105);
nand U27827 (N_27827,N_27376,N_27326);
and U27828 (N_27828,N_27491,N_27230);
nand U27829 (N_27829,N_27203,N_27254);
nand U27830 (N_27830,N_27193,N_27007);
or U27831 (N_27831,N_27402,N_27026);
nor U27832 (N_27832,N_27201,N_27093);
nand U27833 (N_27833,N_27040,N_27169);
nor U27834 (N_27834,N_27387,N_27118);
nor U27835 (N_27835,N_27168,N_27321);
nor U27836 (N_27836,N_27400,N_27292);
and U27837 (N_27837,N_27092,N_27368);
xnor U27838 (N_27838,N_27225,N_27220);
nor U27839 (N_27839,N_27100,N_27197);
nor U27840 (N_27840,N_27030,N_27128);
and U27841 (N_27841,N_27297,N_27471);
and U27842 (N_27842,N_27284,N_27458);
and U27843 (N_27843,N_27117,N_27051);
and U27844 (N_27844,N_27374,N_27341);
or U27845 (N_27845,N_27242,N_27211);
nand U27846 (N_27846,N_27496,N_27462);
xor U27847 (N_27847,N_27299,N_27358);
nor U27848 (N_27848,N_27238,N_27320);
nor U27849 (N_27849,N_27408,N_27379);
nand U27850 (N_27850,N_27457,N_27028);
nor U27851 (N_27851,N_27224,N_27473);
xor U27852 (N_27852,N_27034,N_27070);
nor U27853 (N_27853,N_27192,N_27224);
or U27854 (N_27854,N_27107,N_27123);
nand U27855 (N_27855,N_27234,N_27103);
xor U27856 (N_27856,N_27393,N_27407);
xnor U27857 (N_27857,N_27285,N_27346);
xor U27858 (N_27858,N_27111,N_27327);
and U27859 (N_27859,N_27015,N_27497);
and U27860 (N_27860,N_27382,N_27279);
nand U27861 (N_27861,N_27247,N_27067);
and U27862 (N_27862,N_27488,N_27003);
xor U27863 (N_27863,N_27258,N_27255);
nand U27864 (N_27864,N_27281,N_27403);
and U27865 (N_27865,N_27366,N_27011);
and U27866 (N_27866,N_27292,N_27276);
and U27867 (N_27867,N_27154,N_27406);
nor U27868 (N_27868,N_27420,N_27349);
and U27869 (N_27869,N_27406,N_27120);
nor U27870 (N_27870,N_27157,N_27433);
or U27871 (N_27871,N_27443,N_27178);
or U27872 (N_27872,N_27474,N_27308);
or U27873 (N_27873,N_27361,N_27356);
nand U27874 (N_27874,N_27049,N_27151);
and U27875 (N_27875,N_27140,N_27319);
nand U27876 (N_27876,N_27246,N_27362);
nand U27877 (N_27877,N_27370,N_27044);
nand U27878 (N_27878,N_27172,N_27462);
or U27879 (N_27879,N_27213,N_27254);
or U27880 (N_27880,N_27444,N_27428);
and U27881 (N_27881,N_27311,N_27160);
xnor U27882 (N_27882,N_27443,N_27001);
and U27883 (N_27883,N_27438,N_27186);
or U27884 (N_27884,N_27163,N_27348);
and U27885 (N_27885,N_27490,N_27289);
or U27886 (N_27886,N_27069,N_27064);
or U27887 (N_27887,N_27271,N_27252);
xor U27888 (N_27888,N_27266,N_27034);
nor U27889 (N_27889,N_27100,N_27291);
and U27890 (N_27890,N_27378,N_27039);
and U27891 (N_27891,N_27295,N_27024);
xnor U27892 (N_27892,N_27254,N_27239);
xnor U27893 (N_27893,N_27466,N_27018);
or U27894 (N_27894,N_27038,N_27247);
and U27895 (N_27895,N_27237,N_27391);
xor U27896 (N_27896,N_27477,N_27326);
xor U27897 (N_27897,N_27177,N_27187);
or U27898 (N_27898,N_27150,N_27257);
xnor U27899 (N_27899,N_27191,N_27318);
nor U27900 (N_27900,N_27409,N_27369);
and U27901 (N_27901,N_27135,N_27002);
nor U27902 (N_27902,N_27192,N_27366);
and U27903 (N_27903,N_27311,N_27048);
nor U27904 (N_27904,N_27339,N_27441);
and U27905 (N_27905,N_27181,N_27022);
nand U27906 (N_27906,N_27451,N_27459);
nor U27907 (N_27907,N_27110,N_27106);
nor U27908 (N_27908,N_27371,N_27252);
xnor U27909 (N_27909,N_27144,N_27428);
and U27910 (N_27910,N_27454,N_27432);
or U27911 (N_27911,N_27074,N_27189);
xnor U27912 (N_27912,N_27298,N_27387);
and U27913 (N_27913,N_27383,N_27019);
nor U27914 (N_27914,N_27496,N_27384);
nor U27915 (N_27915,N_27118,N_27217);
and U27916 (N_27916,N_27438,N_27045);
nor U27917 (N_27917,N_27295,N_27455);
nand U27918 (N_27918,N_27452,N_27265);
nor U27919 (N_27919,N_27327,N_27038);
xor U27920 (N_27920,N_27331,N_27419);
or U27921 (N_27921,N_27300,N_27160);
nor U27922 (N_27922,N_27223,N_27075);
nand U27923 (N_27923,N_27383,N_27446);
or U27924 (N_27924,N_27427,N_27320);
nand U27925 (N_27925,N_27331,N_27247);
and U27926 (N_27926,N_27176,N_27063);
xnor U27927 (N_27927,N_27300,N_27046);
or U27928 (N_27928,N_27238,N_27289);
xnor U27929 (N_27929,N_27018,N_27407);
nor U27930 (N_27930,N_27223,N_27176);
xor U27931 (N_27931,N_27036,N_27353);
or U27932 (N_27932,N_27373,N_27323);
or U27933 (N_27933,N_27462,N_27150);
xor U27934 (N_27934,N_27291,N_27270);
nand U27935 (N_27935,N_27383,N_27345);
or U27936 (N_27936,N_27100,N_27174);
or U27937 (N_27937,N_27214,N_27091);
nand U27938 (N_27938,N_27249,N_27033);
and U27939 (N_27939,N_27436,N_27017);
xor U27940 (N_27940,N_27427,N_27106);
and U27941 (N_27941,N_27253,N_27123);
nand U27942 (N_27942,N_27084,N_27426);
or U27943 (N_27943,N_27168,N_27039);
nand U27944 (N_27944,N_27317,N_27270);
or U27945 (N_27945,N_27231,N_27311);
nor U27946 (N_27946,N_27182,N_27185);
xor U27947 (N_27947,N_27019,N_27421);
nor U27948 (N_27948,N_27395,N_27473);
nand U27949 (N_27949,N_27046,N_27281);
nor U27950 (N_27950,N_27095,N_27068);
xnor U27951 (N_27951,N_27039,N_27014);
and U27952 (N_27952,N_27261,N_27118);
nor U27953 (N_27953,N_27328,N_27400);
nand U27954 (N_27954,N_27080,N_27375);
nand U27955 (N_27955,N_27047,N_27331);
nor U27956 (N_27956,N_27069,N_27290);
and U27957 (N_27957,N_27121,N_27100);
nor U27958 (N_27958,N_27235,N_27202);
nand U27959 (N_27959,N_27036,N_27027);
or U27960 (N_27960,N_27406,N_27266);
and U27961 (N_27961,N_27187,N_27104);
nand U27962 (N_27962,N_27437,N_27302);
nor U27963 (N_27963,N_27358,N_27226);
nand U27964 (N_27964,N_27226,N_27144);
xnor U27965 (N_27965,N_27026,N_27009);
or U27966 (N_27966,N_27417,N_27435);
xor U27967 (N_27967,N_27004,N_27311);
xnor U27968 (N_27968,N_27474,N_27353);
or U27969 (N_27969,N_27156,N_27416);
or U27970 (N_27970,N_27108,N_27455);
and U27971 (N_27971,N_27399,N_27182);
and U27972 (N_27972,N_27281,N_27262);
or U27973 (N_27973,N_27463,N_27096);
and U27974 (N_27974,N_27283,N_27220);
or U27975 (N_27975,N_27094,N_27407);
nor U27976 (N_27976,N_27169,N_27209);
nor U27977 (N_27977,N_27453,N_27323);
nor U27978 (N_27978,N_27070,N_27013);
xor U27979 (N_27979,N_27171,N_27175);
or U27980 (N_27980,N_27008,N_27388);
xor U27981 (N_27981,N_27252,N_27437);
xor U27982 (N_27982,N_27304,N_27278);
xnor U27983 (N_27983,N_27211,N_27416);
or U27984 (N_27984,N_27167,N_27062);
xor U27985 (N_27985,N_27433,N_27428);
and U27986 (N_27986,N_27073,N_27358);
nor U27987 (N_27987,N_27018,N_27078);
nor U27988 (N_27988,N_27019,N_27204);
xnor U27989 (N_27989,N_27051,N_27098);
nand U27990 (N_27990,N_27458,N_27300);
nor U27991 (N_27991,N_27275,N_27053);
nor U27992 (N_27992,N_27437,N_27310);
xor U27993 (N_27993,N_27438,N_27419);
nand U27994 (N_27994,N_27175,N_27061);
and U27995 (N_27995,N_27198,N_27483);
or U27996 (N_27996,N_27211,N_27375);
and U27997 (N_27997,N_27403,N_27268);
nor U27998 (N_27998,N_27158,N_27056);
nand U27999 (N_27999,N_27392,N_27498);
or U28000 (N_28000,N_27709,N_27678);
xnor U28001 (N_28001,N_27582,N_27650);
xor U28002 (N_28002,N_27797,N_27707);
nor U28003 (N_28003,N_27549,N_27932);
nor U28004 (N_28004,N_27899,N_27601);
nor U28005 (N_28005,N_27577,N_27662);
nand U28006 (N_28006,N_27552,N_27634);
nand U28007 (N_28007,N_27863,N_27727);
or U28008 (N_28008,N_27668,N_27531);
and U28009 (N_28009,N_27837,N_27908);
xor U28010 (N_28010,N_27706,N_27640);
and U28011 (N_28011,N_27853,N_27567);
xnor U28012 (N_28012,N_27597,N_27902);
nand U28013 (N_28013,N_27819,N_27578);
nor U28014 (N_28014,N_27741,N_27782);
nand U28015 (N_28015,N_27951,N_27547);
xnor U28016 (N_28016,N_27528,N_27967);
nand U28017 (N_28017,N_27935,N_27992);
or U28018 (N_28018,N_27664,N_27912);
nand U28019 (N_28019,N_27649,N_27906);
nor U28020 (N_28020,N_27755,N_27776);
xnor U28021 (N_28021,N_27871,N_27551);
xnor U28022 (N_28022,N_27895,N_27950);
nand U28023 (N_28023,N_27856,N_27620);
xor U28024 (N_28024,N_27897,N_27639);
or U28025 (N_28025,N_27659,N_27811);
xor U28026 (N_28026,N_27826,N_27993);
nand U28027 (N_28027,N_27956,N_27680);
nand U28028 (N_28028,N_27787,N_27999);
or U28029 (N_28029,N_27892,N_27584);
and U28030 (N_28030,N_27847,N_27980);
and U28031 (N_28031,N_27983,N_27687);
nor U28032 (N_28032,N_27541,N_27571);
nor U28033 (N_28033,N_27865,N_27881);
and U28034 (N_28034,N_27548,N_27576);
or U28035 (N_28035,N_27886,N_27593);
nor U28036 (N_28036,N_27922,N_27810);
xnor U28037 (N_28037,N_27596,N_27937);
nand U28038 (N_28038,N_27672,N_27929);
xnor U28039 (N_28039,N_27719,N_27708);
nor U28040 (N_28040,N_27633,N_27798);
xor U28041 (N_28041,N_27774,N_27772);
nor U28042 (N_28042,N_27512,N_27809);
nand U28043 (N_28043,N_27690,N_27845);
and U28044 (N_28044,N_27984,N_27995);
or U28045 (N_28045,N_27813,N_27920);
and U28046 (N_28046,N_27764,N_27927);
nand U28047 (N_28047,N_27978,N_27611);
and U28048 (N_28048,N_27889,N_27830);
and U28049 (N_28049,N_27945,N_27833);
and U28050 (N_28050,N_27900,N_27532);
nor U28051 (N_28051,N_27533,N_27624);
and U28052 (N_28052,N_27511,N_27595);
nor U28053 (N_28053,N_27862,N_27904);
or U28054 (N_28054,N_27786,N_27867);
nor U28055 (N_28055,N_27759,N_27622);
or U28056 (N_28056,N_27580,N_27699);
xor U28057 (N_28057,N_27939,N_27989);
or U28058 (N_28058,N_27665,N_27702);
and U28059 (N_28059,N_27911,N_27733);
and U28060 (N_28060,N_27523,N_27740);
xnor U28061 (N_28061,N_27641,N_27645);
nor U28062 (N_28062,N_27606,N_27613);
and U28063 (N_28063,N_27635,N_27824);
nand U28064 (N_28064,N_27808,N_27944);
or U28065 (N_28065,N_27598,N_27569);
nand U28066 (N_28066,N_27693,N_27679);
or U28067 (N_28067,N_27694,N_27969);
nor U28068 (N_28068,N_27568,N_27636);
nor U28069 (N_28069,N_27973,N_27521);
and U28070 (N_28070,N_27850,N_27591);
or U28071 (N_28071,N_27793,N_27677);
or U28072 (N_28072,N_27643,N_27943);
nand U28073 (N_28073,N_27946,N_27626);
nor U28074 (N_28074,N_27898,N_27891);
and U28075 (N_28075,N_27804,N_27818);
and U28076 (N_28076,N_27996,N_27987);
or U28077 (N_28077,N_27802,N_27617);
and U28078 (N_28078,N_27812,N_27942);
and U28079 (N_28079,N_27689,N_27625);
nor U28080 (N_28080,N_27763,N_27730);
nand U28081 (N_28081,N_27725,N_27988);
nor U28082 (N_28082,N_27926,N_27647);
and U28083 (N_28083,N_27949,N_27785);
or U28084 (N_28084,N_27681,N_27981);
or U28085 (N_28085,N_27803,N_27734);
xor U28086 (N_28086,N_27508,N_27746);
xor U28087 (N_28087,N_27917,N_27752);
nand U28088 (N_28088,N_27692,N_27757);
nand U28089 (N_28089,N_27514,N_27632);
nand U28090 (N_28090,N_27933,N_27843);
nand U28091 (N_28091,N_27691,N_27685);
xor U28092 (N_28092,N_27976,N_27963);
nand U28093 (N_28093,N_27779,N_27873);
and U28094 (N_28094,N_27673,N_27637);
xnor U28095 (N_28095,N_27602,N_27783);
or U28096 (N_28096,N_27924,N_27792);
or U28097 (N_28097,N_27907,N_27657);
and U28098 (N_28098,N_27587,N_27505);
or U28099 (N_28099,N_27948,N_27866);
xnor U28100 (N_28100,N_27775,N_27952);
and U28101 (N_28101,N_27841,N_27758);
xnor U28102 (N_28102,N_27769,N_27807);
and U28103 (N_28103,N_27966,N_27543);
or U28104 (N_28104,N_27638,N_27544);
nand U28105 (N_28105,N_27742,N_27655);
nand U28106 (N_28106,N_27542,N_27799);
nand U28107 (N_28107,N_27723,N_27663);
xor U28108 (N_28108,N_27695,N_27796);
nand U28109 (N_28109,N_27852,N_27923);
nor U28110 (N_28110,N_27817,N_27513);
or U28111 (N_28111,N_27522,N_27502);
and U28112 (N_28112,N_27832,N_27820);
nor U28113 (N_28113,N_27631,N_27936);
xnor U28114 (N_28114,N_27849,N_27930);
or U28115 (N_28115,N_27526,N_27816);
and U28116 (N_28116,N_27844,N_27559);
xor U28117 (N_28117,N_27765,N_27985);
or U28118 (N_28118,N_27729,N_27997);
or U28119 (N_28119,N_27982,N_27861);
nand U28120 (N_28120,N_27656,N_27700);
nand U28121 (N_28121,N_27573,N_27781);
xor U28122 (N_28122,N_27965,N_27768);
and U28123 (N_28123,N_27605,N_27537);
nor U28124 (N_28124,N_27675,N_27676);
xnor U28125 (N_28125,N_27744,N_27516);
nand U28126 (N_28126,N_27991,N_27518);
xor U28127 (N_28127,N_27915,N_27722);
nand U28128 (N_28128,N_27957,N_27860);
xor U28129 (N_28129,N_27747,N_27955);
and U28130 (N_28130,N_27737,N_27885);
nand U28131 (N_28131,N_27652,N_27726);
and U28132 (N_28132,N_27712,N_27884);
nand U28133 (N_28133,N_27750,N_27520);
nor U28134 (N_28134,N_27507,N_27918);
nor U28135 (N_28135,N_27974,N_27960);
and U28136 (N_28136,N_27696,N_27599);
nor U28137 (N_28137,N_27654,N_27877);
nand U28138 (N_28138,N_27749,N_27743);
nor U28139 (N_28139,N_27790,N_27869);
and U28140 (N_28140,N_27686,N_27938);
xor U28141 (N_28141,N_27890,N_27831);
nand U28142 (N_28142,N_27585,N_27773);
xor U28143 (N_28143,N_27684,N_27941);
nor U28144 (N_28144,N_27961,N_27887);
xnor U28145 (N_28145,N_27771,N_27540);
nand U28146 (N_28146,N_27575,N_27754);
nand U28147 (N_28147,N_27829,N_27848);
nand U28148 (N_28148,N_27583,N_27674);
or U28149 (N_28149,N_27834,N_27838);
or U28150 (N_28150,N_27827,N_27697);
and U28151 (N_28151,N_27959,N_27962);
and U28152 (N_28152,N_27555,N_27646);
nor U28153 (N_28153,N_27581,N_27784);
or U28154 (N_28154,N_27565,N_27868);
and U28155 (N_28155,N_27713,N_27500);
nand U28156 (N_28156,N_27735,N_27921);
and U28157 (N_28157,N_27629,N_27710);
and U28158 (N_28158,N_27558,N_27728);
nand U28159 (N_28159,N_27994,N_27736);
nand U28160 (N_28160,N_27627,N_27715);
nand U28161 (N_28161,N_27660,N_27928);
nor U28162 (N_28162,N_27711,N_27964);
or U28163 (N_28163,N_27828,N_27510);
xor U28164 (N_28164,N_27835,N_27971);
nor U28165 (N_28165,N_27671,N_27590);
nand U28166 (N_28166,N_27556,N_27851);
nor U28167 (N_28167,N_27896,N_27751);
xor U28168 (N_28168,N_27954,N_27714);
nor U28169 (N_28169,N_27509,N_27958);
or U28170 (N_28170,N_27731,N_27880);
nand U28171 (N_28171,N_27604,N_27801);
and U28172 (N_28172,N_27854,N_27519);
nand U28173 (N_28173,N_27846,N_27610);
or U28174 (N_28174,N_27986,N_27653);
and U28175 (N_28175,N_27570,N_27839);
nor U28176 (N_28176,N_27574,N_27883);
xor U28177 (N_28177,N_27720,N_27623);
or U28178 (N_28178,N_27872,N_27795);
and U28179 (N_28179,N_27683,N_27882);
and U28180 (N_28180,N_27536,N_27562);
or U28181 (N_28181,N_27608,N_27762);
nor U28182 (N_28182,N_27539,N_27527);
xnor U28183 (N_28183,N_27703,N_27651);
nor U28184 (N_28184,N_27858,N_27893);
nand U28185 (N_28185,N_27588,N_27572);
nor U28186 (N_28186,N_27778,N_27721);
nor U28187 (N_28187,N_27756,N_27910);
and U28188 (N_28188,N_27879,N_27716);
nor U28189 (N_28189,N_27825,N_27990);
nand U28190 (N_28190,N_27717,N_27970);
and U28191 (N_28191,N_27688,N_27524);
nand U28192 (N_28192,N_27972,N_27529);
nor U28193 (N_28193,N_27564,N_27557);
or U28194 (N_28194,N_27934,N_27916);
nor U28195 (N_28195,N_27586,N_27864);
xor U28196 (N_28196,N_27550,N_27615);
nand U28197 (N_28197,N_27770,N_27738);
xnor U28198 (N_28198,N_27621,N_27561);
or U28199 (N_28199,N_27953,N_27682);
nor U28200 (N_28200,N_27822,N_27925);
xor U28201 (N_28201,N_27805,N_27670);
xnor U28202 (N_28202,N_27840,N_27628);
or U28203 (N_28203,N_27517,N_27592);
and U28204 (N_28204,N_27501,N_27913);
and U28205 (N_28205,N_27698,N_27530);
nand U28206 (N_28206,N_27648,N_27780);
nand U28207 (N_28207,N_27594,N_27903);
and U28208 (N_28208,N_27515,N_27732);
xor U28209 (N_28209,N_27503,N_27905);
and U28210 (N_28210,N_27619,N_27876);
and U28211 (N_28211,N_27909,N_27745);
and U28212 (N_28212,N_27975,N_27607);
nor U28213 (N_28213,N_27870,N_27603);
or U28214 (N_28214,N_27800,N_27761);
or U28215 (N_28215,N_27894,N_27998);
nor U28216 (N_28216,N_27614,N_27718);
nor U28217 (N_28217,N_27566,N_27612);
xor U28218 (N_28218,N_27609,N_27525);
and U28219 (N_28219,N_27667,N_27748);
nand U28220 (N_28220,N_27791,N_27875);
or U28221 (N_28221,N_27901,N_27669);
xnor U28222 (N_28222,N_27506,N_27979);
and U28223 (N_28223,N_27724,N_27579);
xor U28224 (N_28224,N_27767,N_27788);
xnor U28225 (N_28225,N_27821,N_27947);
nor U28226 (N_28226,N_27630,N_27968);
or U28227 (N_28227,N_27560,N_27546);
nor U28228 (N_28228,N_27538,N_27794);
nor U28229 (N_28229,N_27642,N_27545);
or U28230 (N_28230,N_27704,N_27842);
nand U28231 (N_28231,N_27589,N_27874);
and U28232 (N_28232,N_27919,N_27777);
or U28233 (N_28233,N_27616,N_27701);
and U28234 (N_28234,N_27814,N_27705);
or U28235 (N_28235,N_27658,N_27644);
xor U28236 (N_28236,N_27766,N_27661);
nor U28237 (N_28237,N_27823,N_27666);
nand U28238 (N_28238,N_27940,N_27815);
xor U28239 (N_28239,N_27504,N_27855);
and U28240 (N_28240,N_27888,N_27931);
or U28241 (N_28241,N_27534,N_27914);
xnor U28242 (N_28242,N_27739,N_27836);
nand U28243 (N_28243,N_27554,N_27563);
xnor U28244 (N_28244,N_27857,N_27553);
and U28245 (N_28245,N_27753,N_27535);
xor U28246 (N_28246,N_27977,N_27789);
nand U28247 (N_28247,N_27618,N_27600);
nand U28248 (N_28248,N_27760,N_27878);
nand U28249 (N_28249,N_27859,N_27806);
or U28250 (N_28250,N_27628,N_27984);
or U28251 (N_28251,N_27500,N_27820);
and U28252 (N_28252,N_27959,N_27609);
xor U28253 (N_28253,N_27610,N_27512);
and U28254 (N_28254,N_27742,N_27716);
and U28255 (N_28255,N_27923,N_27520);
nand U28256 (N_28256,N_27942,N_27768);
xor U28257 (N_28257,N_27637,N_27646);
and U28258 (N_28258,N_27760,N_27647);
xor U28259 (N_28259,N_27885,N_27909);
and U28260 (N_28260,N_27961,N_27526);
nor U28261 (N_28261,N_27959,N_27654);
nand U28262 (N_28262,N_27561,N_27997);
nor U28263 (N_28263,N_27807,N_27665);
nor U28264 (N_28264,N_27598,N_27929);
xnor U28265 (N_28265,N_27797,N_27965);
nor U28266 (N_28266,N_27862,N_27924);
or U28267 (N_28267,N_27723,N_27859);
and U28268 (N_28268,N_27991,N_27554);
and U28269 (N_28269,N_27538,N_27925);
nor U28270 (N_28270,N_27524,N_27801);
xor U28271 (N_28271,N_27609,N_27956);
or U28272 (N_28272,N_27881,N_27522);
and U28273 (N_28273,N_27734,N_27571);
and U28274 (N_28274,N_27580,N_27889);
and U28275 (N_28275,N_27935,N_27625);
xor U28276 (N_28276,N_27888,N_27536);
xor U28277 (N_28277,N_27543,N_27544);
and U28278 (N_28278,N_27609,N_27771);
nand U28279 (N_28279,N_27704,N_27910);
nor U28280 (N_28280,N_27680,N_27691);
or U28281 (N_28281,N_27868,N_27629);
xnor U28282 (N_28282,N_27912,N_27675);
xnor U28283 (N_28283,N_27914,N_27543);
nor U28284 (N_28284,N_27599,N_27559);
nand U28285 (N_28285,N_27994,N_27688);
xnor U28286 (N_28286,N_27637,N_27743);
and U28287 (N_28287,N_27967,N_27988);
xor U28288 (N_28288,N_27849,N_27788);
or U28289 (N_28289,N_27984,N_27675);
xor U28290 (N_28290,N_27577,N_27921);
or U28291 (N_28291,N_27820,N_27671);
or U28292 (N_28292,N_27765,N_27805);
or U28293 (N_28293,N_27625,N_27620);
or U28294 (N_28294,N_27800,N_27707);
and U28295 (N_28295,N_27575,N_27581);
or U28296 (N_28296,N_27962,N_27658);
nand U28297 (N_28297,N_27800,N_27876);
nor U28298 (N_28298,N_27732,N_27559);
nor U28299 (N_28299,N_27936,N_27651);
and U28300 (N_28300,N_27786,N_27620);
nor U28301 (N_28301,N_27892,N_27872);
xnor U28302 (N_28302,N_27739,N_27780);
nand U28303 (N_28303,N_27669,N_27605);
nor U28304 (N_28304,N_27521,N_27718);
nand U28305 (N_28305,N_27580,N_27680);
nor U28306 (N_28306,N_27572,N_27959);
xnor U28307 (N_28307,N_27632,N_27995);
or U28308 (N_28308,N_27750,N_27937);
or U28309 (N_28309,N_27552,N_27538);
nand U28310 (N_28310,N_27775,N_27794);
nor U28311 (N_28311,N_27551,N_27532);
and U28312 (N_28312,N_27787,N_27893);
and U28313 (N_28313,N_27885,N_27984);
nor U28314 (N_28314,N_27593,N_27623);
xor U28315 (N_28315,N_27689,N_27659);
and U28316 (N_28316,N_27822,N_27958);
nor U28317 (N_28317,N_27770,N_27797);
or U28318 (N_28318,N_27554,N_27733);
or U28319 (N_28319,N_27771,N_27935);
nand U28320 (N_28320,N_27700,N_27968);
and U28321 (N_28321,N_27562,N_27853);
xor U28322 (N_28322,N_27604,N_27966);
nor U28323 (N_28323,N_27524,N_27838);
xnor U28324 (N_28324,N_27882,N_27655);
xnor U28325 (N_28325,N_27610,N_27884);
nand U28326 (N_28326,N_27782,N_27922);
nand U28327 (N_28327,N_27646,N_27868);
nand U28328 (N_28328,N_27678,N_27632);
nor U28329 (N_28329,N_27575,N_27626);
xor U28330 (N_28330,N_27815,N_27865);
nor U28331 (N_28331,N_27740,N_27822);
nor U28332 (N_28332,N_27844,N_27912);
or U28333 (N_28333,N_27594,N_27835);
nand U28334 (N_28334,N_27566,N_27623);
nor U28335 (N_28335,N_27520,N_27739);
and U28336 (N_28336,N_27869,N_27508);
or U28337 (N_28337,N_27714,N_27510);
and U28338 (N_28338,N_27860,N_27539);
nor U28339 (N_28339,N_27593,N_27832);
nor U28340 (N_28340,N_27504,N_27740);
xor U28341 (N_28341,N_27750,N_27566);
xnor U28342 (N_28342,N_27907,N_27914);
nor U28343 (N_28343,N_27890,N_27840);
and U28344 (N_28344,N_27567,N_27970);
or U28345 (N_28345,N_27935,N_27592);
and U28346 (N_28346,N_27624,N_27809);
nor U28347 (N_28347,N_27779,N_27617);
nand U28348 (N_28348,N_27732,N_27934);
or U28349 (N_28349,N_27993,N_27779);
nand U28350 (N_28350,N_27915,N_27648);
xor U28351 (N_28351,N_27956,N_27779);
nand U28352 (N_28352,N_27550,N_27999);
xor U28353 (N_28353,N_27553,N_27942);
xor U28354 (N_28354,N_27522,N_27503);
nand U28355 (N_28355,N_27615,N_27706);
and U28356 (N_28356,N_27803,N_27723);
or U28357 (N_28357,N_27540,N_27704);
xor U28358 (N_28358,N_27962,N_27820);
and U28359 (N_28359,N_27855,N_27949);
nor U28360 (N_28360,N_27947,N_27557);
or U28361 (N_28361,N_27617,N_27750);
xnor U28362 (N_28362,N_27864,N_27573);
and U28363 (N_28363,N_27690,N_27594);
or U28364 (N_28364,N_27642,N_27707);
nor U28365 (N_28365,N_27693,N_27866);
and U28366 (N_28366,N_27840,N_27543);
nor U28367 (N_28367,N_27786,N_27543);
xnor U28368 (N_28368,N_27502,N_27715);
and U28369 (N_28369,N_27552,N_27847);
nand U28370 (N_28370,N_27734,N_27601);
xnor U28371 (N_28371,N_27789,N_27791);
and U28372 (N_28372,N_27636,N_27788);
nor U28373 (N_28373,N_27777,N_27619);
and U28374 (N_28374,N_27952,N_27909);
nor U28375 (N_28375,N_27779,N_27758);
or U28376 (N_28376,N_27752,N_27790);
or U28377 (N_28377,N_27647,N_27952);
nor U28378 (N_28378,N_27751,N_27673);
nand U28379 (N_28379,N_27599,N_27821);
nand U28380 (N_28380,N_27682,N_27525);
or U28381 (N_28381,N_27535,N_27582);
and U28382 (N_28382,N_27948,N_27553);
and U28383 (N_28383,N_27630,N_27908);
or U28384 (N_28384,N_27738,N_27843);
xor U28385 (N_28385,N_27741,N_27876);
or U28386 (N_28386,N_27761,N_27516);
xor U28387 (N_28387,N_27886,N_27743);
or U28388 (N_28388,N_27552,N_27504);
or U28389 (N_28389,N_27668,N_27566);
or U28390 (N_28390,N_27528,N_27588);
xor U28391 (N_28391,N_27966,N_27760);
nor U28392 (N_28392,N_27542,N_27764);
nand U28393 (N_28393,N_27846,N_27694);
xor U28394 (N_28394,N_27971,N_27707);
nor U28395 (N_28395,N_27998,N_27772);
or U28396 (N_28396,N_27528,N_27648);
nand U28397 (N_28397,N_27529,N_27689);
or U28398 (N_28398,N_27706,N_27702);
nand U28399 (N_28399,N_27804,N_27751);
and U28400 (N_28400,N_27965,N_27512);
nor U28401 (N_28401,N_27959,N_27954);
nand U28402 (N_28402,N_27904,N_27838);
and U28403 (N_28403,N_27808,N_27711);
nand U28404 (N_28404,N_27500,N_27793);
nor U28405 (N_28405,N_27862,N_27539);
nor U28406 (N_28406,N_27609,N_27546);
xnor U28407 (N_28407,N_27976,N_27577);
xnor U28408 (N_28408,N_27801,N_27536);
nand U28409 (N_28409,N_27669,N_27861);
nor U28410 (N_28410,N_27880,N_27618);
or U28411 (N_28411,N_27842,N_27854);
xnor U28412 (N_28412,N_27875,N_27521);
and U28413 (N_28413,N_27669,N_27931);
xor U28414 (N_28414,N_27791,N_27855);
nor U28415 (N_28415,N_27908,N_27648);
nor U28416 (N_28416,N_27976,N_27959);
and U28417 (N_28417,N_27876,N_27745);
xnor U28418 (N_28418,N_27667,N_27799);
nor U28419 (N_28419,N_27957,N_27638);
xnor U28420 (N_28420,N_27886,N_27827);
nand U28421 (N_28421,N_27624,N_27677);
xor U28422 (N_28422,N_27601,N_27903);
or U28423 (N_28423,N_27769,N_27635);
nor U28424 (N_28424,N_27956,N_27891);
nand U28425 (N_28425,N_27670,N_27639);
nor U28426 (N_28426,N_27834,N_27701);
and U28427 (N_28427,N_27740,N_27881);
nor U28428 (N_28428,N_27703,N_27612);
xnor U28429 (N_28429,N_27519,N_27995);
nand U28430 (N_28430,N_27836,N_27768);
nand U28431 (N_28431,N_27748,N_27664);
and U28432 (N_28432,N_27948,N_27635);
nand U28433 (N_28433,N_27856,N_27869);
or U28434 (N_28434,N_27563,N_27705);
and U28435 (N_28435,N_27686,N_27804);
nor U28436 (N_28436,N_27702,N_27771);
or U28437 (N_28437,N_27519,N_27839);
and U28438 (N_28438,N_27501,N_27705);
xnor U28439 (N_28439,N_27898,N_27924);
nor U28440 (N_28440,N_27748,N_27830);
xor U28441 (N_28441,N_27618,N_27884);
or U28442 (N_28442,N_27977,N_27693);
xor U28443 (N_28443,N_27996,N_27525);
xor U28444 (N_28444,N_27819,N_27858);
nor U28445 (N_28445,N_27979,N_27797);
nor U28446 (N_28446,N_27815,N_27691);
xnor U28447 (N_28447,N_27847,N_27661);
nor U28448 (N_28448,N_27799,N_27980);
or U28449 (N_28449,N_27710,N_27961);
or U28450 (N_28450,N_27836,N_27720);
nand U28451 (N_28451,N_27888,N_27964);
and U28452 (N_28452,N_27707,N_27873);
nor U28453 (N_28453,N_27766,N_27534);
or U28454 (N_28454,N_27624,N_27939);
and U28455 (N_28455,N_27750,N_27995);
xor U28456 (N_28456,N_27745,N_27697);
nand U28457 (N_28457,N_27744,N_27807);
and U28458 (N_28458,N_27894,N_27620);
nand U28459 (N_28459,N_27794,N_27866);
xnor U28460 (N_28460,N_27782,N_27882);
nand U28461 (N_28461,N_27942,N_27830);
and U28462 (N_28462,N_27961,N_27760);
nor U28463 (N_28463,N_27637,N_27676);
and U28464 (N_28464,N_27912,N_27753);
and U28465 (N_28465,N_27564,N_27877);
nor U28466 (N_28466,N_27941,N_27892);
or U28467 (N_28467,N_27954,N_27547);
nor U28468 (N_28468,N_27630,N_27762);
xor U28469 (N_28469,N_27689,N_27873);
nand U28470 (N_28470,N_27901,N_27703);
or U28471 (N_28471,N_27780,N_27886);
and U28472 (N_28472,N_27981,N_27800);
nor U28473 (N_28473,N_27833,N_27508);
and U28474 (N_28474,N_27611,N_27706);
and U28475 (N_28475,N_27557,N_27909);
xnor U28476 (N_28476,N_27857,N_27675);
nor U28477 (N_28477,N_27576,N_27858);
xor U28478 (N_28478,N_27651,N_27989);
xnor U28479 (N_28479,N_27933,N_27502);
or U28480 (N_28480,N_27864,N_27643);
or U28481 (N_28481,N_27826,N_27587);
or U28482 (N_28482,N_27888,N_27968);
nor U28483 (N_28483,N_27943,N_27756);
or U28484 (N_28484,N_27535,N_27854);
xnor U28485 (N_28485,N_27787,N_27586);
nor U28486 (N_28486,N_27717,N_27605);
nand U28487 (N_28487,N_27954,N_27923);
and U28488 (N_28488,N_27991,N_27617);
or U28489 (N_28489,N_27574,N_27847);
xor U28490 (N_28490,N_27852,N_27738);
nand U28491 (N_28491,N_27987,N_27691);
and U28492 (N_28492,N_27970,N_27688);
xnor U28493 (N_28493,N_27571,N_27623);
and U28494 (N_28494,N_27597,N_27839);
or U28495 (N_28495,N_27789,N_27957);
nand U28496 (N_28496,N_27555,N_27504);
nand U28497 (N_28497,N_27694,N_27776);
nand U28498 (N_28498,N_27604,N_27671);
nor U28499 (N_28499,N_27725,N_27782);
nand U28500 (N_28500,N_28048,N_28244);
nand U28501 (N_28501,N_28465,N_28371);
and U28502 (N_28502,N_28387,N_28334);
and U28503 (N_28503,N_28132,N_28006);
xor U28504 (N_28504,N_28112,N_28360);
and U28505 (N_28505,N_28150,N_28097);
nand U28506 (N_28506,N_28369,N_28215);
and U28507 (N_28507,N_28299,N_28038);
nor U28508 (N_28508,N_28264,N_28256);
nor U28509 (N_28509,N_28399,N_28195);
or U28510 (N_28510,N_28217,N_28318);
and U28511 (N_28511,N_28446,N_28303);
xnor U28512 (N_28512,N_28285,N_28449);
or U28513 (N_28513,N_28122,N_28356);
and U28514 (N_28514,N_28070,N_28065);
nor U28515 (N_28515,N_28407,N_28290);
or U28516 (N_28516,N_28379,N_28046);
or U28517 (N_28517,N_28296,N_28293);
xnor U28518 (N_28518,N_28301,N_28436);
xnor U28519 (N_28519,N_28343,N_28140);
or U28520 (N_28520,N_28003,N_28312);
nand U28521 (N_28521,N_28309,N_28052);
nor U28522 (N_28522,N_28317,N_28497);
nor U28523 (N_28523,N_28345,N_28137);
nor U28524 (N_28524,N_28492,N_28222);
nand U28525 (N_28525,N_28372,N_28289);
or U28526 (N_28526,N_28454,N_28035);
and U28527 (N_28527,N_28287,N_28120);
xnor U28528 (N_28528,N_28457,N_28258);
or U28529 (N_28529,N_28431,N_28197);
nand U28530 (N_28530,N_28490,N_28023);
or U28531 (N_28531,N_28445,N_28257);
nor U28532 (N_28532,N_28094,N_28022);
and U28533 (N_28533,N_28152,N_28327);
and U28534 (N_28534,N_28131,N_28057);
nand U28535 (N_28535,N_28267,N_28425);
and U28536 (N_28536,N_28169,N_28037);
or U28537 (N_28537,N_28040,N_28423);
or U28538 (N_28538,N_28242,N_28300);
and U28539 (N_28539,N_28216,N_28391);
and U28540 (N_28540,N_28382,N_28366);
nand U28541 (N_28541,N_28085,N_28098);
nand U28542 (N_28542,N_28471,N_28117);
and U28543 (N_28543,N_28050,N_28253);
nor U28544 (N_28544,N_28495,N_28370);
or U28545 (N_28545,N_28136,N_28283);
and U28546 (N_28546,N_28077,N_28437);
and U28547 (N_28547,N_28376,N_28108);
nand U28548 (N_28548,N_28208,N_28075);
and U28549 (N_28549,N_28099,N_28450);
or U28550 (N_28550,N_28126,N_28173);
and U28551 (N_28551,N_28196,N_28170);
xnor U28552 (N_28552,N_28246,N_28281);
xor U28553 (N_28553,N_28092,N_28335);
nand U28554 (N_28554,N_28073,N_28282);
and U28555 (N_28555,N_28359,N_28165);
or U28556 (N_28556,N_28347,N_28466);
nor U28557 (N_28557,N_28453,N_28314);
and U28558 (N_28558,N_28090,N_28459);
or U28559 (N_28559,N_28342,N_28109);
nor U28560 (N_28560,N_28072,N_28395);
nand U28561 (N_28561,N_28306,N_28275);
nor U28562 (N_28562,N_28115,N_28033);
or U28563 (N_28563,N_28199,N_28451);
or U28564 (N_28564,N_28234,N_28354);
nand U28565 (N_28565,N_28277,N_28361);
xor U28566 (N_28566,N_28381,N_28491);
or U28567 (N_28567,N_28460,N_28262);
or U28568 (N_28568,N_28499,N_28420);
nand U28569 (N_28569,N_28002,N_28426);
and U28570 (N_28570,N_28144,N_28212);
nor U28571 (N_28571,N_28185,N_28326);
nand U28572 (N_28572,N_28175,N_28268);
xnor U28573 (N_28573,N_28427,N_28053);
nor U28574 (N_28574,N_28367,N_28153);
or U28575 (N_28575,N_28396,N_28486);
and U28576 (N_28576,N_28424,N_28051);
or U28577 (N_28577,N_28042,N_28362);
and U28578 (N_28578,N_28406,N_28164);
nand U28579 (N_28579,N_28288,N_28076);
xor U28580 (N_28580,N_28266,N_28435);
xnor U28581 (N_28581,N_28167,N_28284);
nor U28582 (N_28582,N_28104,N_28337);
nand U28583 (N_28583,N_28349,N_28438);
and U28584 (N_28584,N_28422,N_28021);
or U28585 (N_28585,N_28404,N_28027);
or U28586 (N_28586,N_28029,N_28232);
nor U28587 (N_28587,N_28470,N_28194);
nor U28588 (N_28588,N_28355,N_28031);
and U28589 (N_28589,N_28074,N_28239);
nor U28590 (N_28590,N_28125,N_28351);
nand U28591 (N_28591,N_28339,N_28341);
xor U28592 (N_28592,N_28352,N_28340);
nor U28593 (N_28593,N_28313,N_28014);
nand U28594 (N_28594,N_28020,N_28237);
and U28595 (N_28595,N_28363,N_28260);
or U28596 (N_28596,N_28114,N_28214);
and U28597 (N_28597,N_28015,N_28079);
nand U28598 (N_28598,N_28291,N_28478);
nor U28599 (N_28599,N_28064,N_28297);
xnor U28600 (N_28600,N_28101,N_28328);
or U28601 (N_28601,N_28154,N_28276);
nand U28602 (N_28602,N_28250,N_28129);
or U28603 (N_28603,N_28026,N_28148);
xor U28604 (N_28604,N_28230,N_28388);
xnor U28605 (N_28605,N_28025,N_28008);
or U28606 (N_28606,N_28482,N_28383);
or U28607 (N_28607,N_28107,N_28146);
nand U28608 (N_28608,N_28187,N_28028);
or U28609 (N_28609,N_28413,N_28163);
xor U28610 (N_28610,N_28350,N_28274);
xnor U28611 (N_28611,N_28261,N_28385);
nor U28612 (N_28612,N_28389,N_28176);
and U28613 (N_28613,N_28200,N_28496);
xor U28614 (N_28614,N_28224,N_28178);
and U28615 (N_28615,N_28087,N_28294);
and U28616 (N_28616,N_28494,N_28047);
xor U28617 (N_28617,N_28174,N_28304);
and U28618 (N_28618,N_28201,N_28102);
and U28619 (N_28619,N_28130,N_28330);
xor U28620 (N_28620,N_28213,N_28166);
xor U28621 (N_28621,N_28316,N_28365);
or U28622 (N_28622,N_28429,N_28059);
and U28623 (N_28623,N_28123,N_28386);
xor U28624 (N_28624,N_28447,N_28093);
or U28625 (N_28625,N_28182,N_28039);
nor U28626 (N_28626,N_28333,N_28018);
and U28627 (N_28627,N_28373,N_28408);
nand U28628 (N_28628,N_28469,N_28010);
xor U28629 (N_28629,N_28134,N_28004);
xnor U28630 (N_28630,N_28251,N_28172);
nand U28631 (N_28631,N_28433,N_28078);
or U28632 (N_28632,N_28226,N_28168);
xor U28633 (N_28633,N_28045,N_28069);
xnor U28634 (N_28634,N_28011,N_28088);
nand U28635 (N_28635,N_28189,N_28374);
or U28636 (N_28636,N_28398,N_28181);
nand U28637 (N_28637,N_28394,N_28206);
nor U28638 (N_28638,N_28468,N_28302);
nor U28639 (N_28639,N_28411,N_28151);
and U28640 (N_28640,N_28141,N_28060);
xor U28641 (N_28641,N_28205,N_28241);
nor U28642 (N_28642,N_28418,N_28012);
nor U28643 (N_28643,N_28209,N_28332);
nor U28644 (N_28644,N_28311,N_28179);
nor U28645 (N_28645,N_28116,N_28013);
nor U28646 (N_28646,N_28377,N_28259);
nand U28647 (N_28647,N_28248,N_28477);
xor U28648 (N_28648,N_28041,N_28400);
or U28649 (N_28649,N_28443,N_28393);
or U28650 (N_28650,N_28384,N_28127);
xnor U28651 (N_28651,N_28061,N_28448);
nand U28652 (N_28652,N_28485,N_28188);
xor U28653 (N_28653,N_28263,N_28473);
and U28654 (N_28654,N_28358,N_28110);
nor U28655 (N_28655,N_28286,N_28236);
or U28656 (N_28656,N_28410,N_28211);
nand U28657 (N_28657,N_28062,N_28017);
nand U28658 (N_28658,N_28269,N_28489);
xnor U28659 (N_28659,N_28220,N_28005);
nand U28660 (N_28660,N_28001,N_28229);
xor U28661 (N_28661,N_28066,N_28193);
nor U28662 (N_28662,N_28105,N_28055);
nand U28663 (N_28663,N_28180,N_28476);
nand U28664 (N_28664,N_28414,N_28219);
and U28665 (N_28665,N_28428,N_28320);
nand U28666 (N_28666,N_28081,N_28067);
and U28667 (N_28667,N_28484,N_28121);
nand U28668 (N_28668,N_28292,N_28095);
xor U28669 (N_28669,N_28442,N_28083);
nand U28670 (N_28670,N_28156,N_28171);
nand U28671 (N_28671,N_28049,N_28016);
xor U28672 (N_28672,N_28159,N_28397);
or U28673 (N_28673,N_28056,N_28405);
and U28674 (N_28674,N_28135,N_28124);
nand U28675 (N_28675,N_28307,N_28338);
and U28676 (N_28676,N_28128,N_28331);
nor U28677 (N_28677,N_28145,N_28392);
or U28678 (N_28678,N_28207,N_28009);
xnor U28679 (N_28679,N_28249,N_28390);
xor U28680 (N_28680,N_28402,N_28329);
xor U28681 (N_28681,N_28007,N_28325);
or U28682 (N_28682,N_28380,N_28255);
and U28683 (N_28683,N_28203,N_28142);
and U28684 (N_28684,N_28462,N_28401);
nand U28685 (N_28685,N_28498,N_28147);
xor U28686 (N_28686,N_28487,N_28063);
xor U28687 (N_28687,N_28254,N_28158);
nor U28688 (N_28688,N_28440,N_28235);
nor U28689 (N_28689,N_28421,N_28204);
nor U28690 (N_28690,N_28344,N_28278);
and U28691 (N_28691,N_28412,N_28080);
nand U28692 (N_28692,N_28223,N_28228);
and U28693 (N_28693,N_28032,N_28348);
and U28694 (N_28694,N_28475,N_28084);
or U28695 (N_28695,N_28044,N_28240);
xor U28696 (N_28696,N_28430,N_28096);
or U28697 (N_28697,N_28210,N_28310);
xor U28698 (N_28698,N_28456,N_28324);
nor U28699 (N_28699,N_28162,N_28184);
xor U28700 (N_28700,N_28227,N_28265);
and U28701 (N_28701,N_28243,N_28225);
xor U28702 (N_28702,N_28272,N_28054);
xor U28703 (N_28703,N_28036,N_28375);
nor U28704 (N_28704,N_28118,N_28472);
and U28705 (N_28705,N_28247,N_28364);
xnor U28706 (N_28706,N_28091,N_28419);
or U28707 (N_28707,N_28068,N_28202);
or U28708 (N_28708,N_28280,N_28493);
or U28709 (N_28709,N_28415,N_28019);
and U28710 (N_28710,N_28160,N_28319);
nor U28711 (N_28711,N_28461,N_28321);
and U28712 (N_28712,N_28298,N_28191);
xor U28713 (N_28713,N_28416,N_28183);
and U28714 (N_28714,N_28481,N_28024);
nand U28715 (N_28715,N_28353,N_28441);
or U28716 (N_28716,N_28323,N_28138);
xnor U28717 (N_28717,N_28030,N_28043);
nor U28718 (N_28718,N_28058,N_28368);
nand U28719 (N_28719,N_28198,N_28089);
or U28720 (N_28720,N_28157,N_28270);
nor U28721 (N_28721,N_28467,N_28100);
nor U28722 (N_28722,N_28322,N_28161);
and U28723 (N_28723,N_28474,N_28119);
nor U28724 (N_28724,N_28279,N_28452);
xor U28725 (N_28725,N_28315,N_28177);
xnor U28726 (N_28726,N_28455,N_28403);
or U28727 (N_28727,N_28488,N_28133);
nor U28728 (N_28728,N_28218,N_28308);
or U28729 (N_28729,N_28082,N_28221);
xnor U28730 (N_28730,N_28238,N_28463);
nand U28731 (N_28731,N_28439,N_28252);
xnor U28732 (N_28732,N_28458,N_28143);
and U28733 (N_28733,N_28378,N_28417);
and U28734 (N_28734,N_28444,N_28357);
nor U28735 (N_28735,N_28409,N_28305);
xnor U28736 (N_28736,N_28231,N_28479);
or U28737 (N_28737,N_28000,N_28245);
xnor U28738 (N_28738,N_28071,N_28346);
and U28739 (N_28739,N_28271,N_28106);
xnor U28740 (N_28740,N_28464,N_28034);
nor U28741 (N_28741,N_28186,N_28434);
nand U28742 (N_28742,N_28155,N_28190);
and U28743 (N_28743,N_28113,N_28111);
nand U28744 (N_28744,N_28483,N_28295);
and U28745 (N_28745,N_28273,N_28086);
nand U28746 (N_28746,N_28336,N_28432);
or U28747 (N_28747,N_28192,N_28103);
nand U28748 (N_28748,N_28480,N_28149);
or U28749 (N_28749,N_28139,N_28233);
or U28750 (N_28750,N_28228,N_28186);
and U28751 (N_28751,N_28467,N_28082);
xor U28752 (N_28752,N_28192,N_28117);
xnor U28753 (N_28753,N_28005,N_28150);
nor U28754 (N_28754,N_28314,N_28351);
nand U28755 (N_28755,N_28250,N_28004);
nor U28756 (N_28756,N_28264,N_28067);
or U28757 (N_28757,N_28397,N_28170);
nor U28758 (N_28758,N_28492,N_28371);
and U28759 (N_28759,N_28442,N_28348);
or U28760 (N_28760,N_28303,N_28167);
nand U28761 (N_28761,N_28255,N_28186);
or U28762 (N_28762,N_28189,N_28339);
nand U28763 (N_28763,N_28140,N_28346);
nor U28764 (N_28764,N_28285,N_28025);
or U28765 (N_28765,N_28347,N_28022);
and U28766 (N_28766,N_28162,N_28367);
or U28767 (N_28767,N_28306,N_28324);
nor U28768 (N_28768,N_28183,N_28032);
nor U28769 (N_28769,N_28224,N_28435);
or U28770 (N_28770,N_28213,N_28448);
xnor U28771 (N_28771,N_28347,N_28475);
xnor U28772 (N_28772,N_28359,N_28422);
nand U28773 (N_28773,N_28151,N_28023);
nor U28774 (N_28774,N_28339,N_28029);
nor U28775 (N_28775,N_28265,N_28109);
xor U28776 (N_28776,N_28301,N_28387);
and U28777 (N_28777,N_28376,N_28493);
nand U28778 (N_28778,N_28337,N_28261);
nor U28779 (N_28779,N_28317,N_28106);
or U28780 (N_28780,N_28093,N_28211);
xnor U28781 (N_28781,N_28158,N_28199);
nand U28782 (N_28782,N_28148,N_28357);
xnor U28783 (N_28783,N_28431,N_28192);
nand U28784 (N_28784,N_28395,N_28219);
xor U28785 (N_28785,N_28311,N_28233);
nor U28786 (N_28786,N_28190,N_28206);
or U28787 (N_28787,N_28005,N_28191);
or U28788 (N_28788,N_28169,N_28141);
and U28789 (N_28789,N_28061,N_28015);
nand U28790 (N_28790,N_28009,N_28485);
and U28791 (N_28791,N_28196,N_28437);
xor U28792 (N_28792,N_28445,N_28021);
or U28793 (N_28793,N_28440,N_28450);
nand U28794 (N_28794,N_28259,N_28196);
xnor U28795 (N_28795,N_28005,N_28226);
or U28796 (N_28796,N_28351,N_28372);
and U28797 (N_28797,N_28236,N_28360);
nand U28798 (N_28798,N_28251,N_28177);
or U28799 (N_28799,N_28303,N_28043);
xnor U28800 (N_28800,N_28154,N_28091);
nor U28801 (N_28801,N_28348,N_28163);
and U28802 (N_28802,N_28055,N_28384);
nand U28803 (N_28803,N_28105,N_28414);
nor U28804 (N_28804,N_28494,N_28230);
nor U28805 (N_28805,N_28130,N_28273);
or U28806 (N_28806,N_28391,N_28496);
or U28807 (N_28807,N_28102,N_28217);
nor U28808 (N_28808,N_28389,N_28254);
or U28809 (N_28809,N_28203,N_28008);
nand U28810 (N_28810,N_28370,N_28237);
nand U28811 (N_28811,N_28233,N_28044);
or U28812 (N_28812,N_28101,N_28287);
xnor U28813 (N_28813,N_28022,N_28153);
nor U28814 (N_28814,N_28110,N_28053);
nor U28815 (N_28815,N_28136,N_28080);
or U28816 (N_28816,N_28379,N_28414);
nor U28817 (N_28817,N_28194,N_28123);
or U28818 (N_28818,N_28487,N_28453);
and U28819 (N_28819,N_28131,N_28127);
xnor U28820 (N_28820,N_28380,N_28049);
nand U28821 (N_28821,N_28439,N_28408);
or U28822 (N_28822,N_28387,N_28253);
nor U28823 (N_28823,N_28361,N_28341);
xor U28824 (N_28824,N_28132,N_28093);
nand U28825 (N_28825,N_28073,N_28213);
xnor U28826 (N_28826,N_28189,N_28351);
or U28827 (N_28827,N_28054,N_28276);
xnor U28828 (N_28828,N_28288,N_28011);
nand U28829 (N_28829,N_28221,N_28405);
or U28830 (N_28830,N_28031,N_28042);
and U28831 (N_28831,N_28185,N_28216);
nand U28832 (N_28832,N_28223,N_28126);
xor U28833 (N_28833,N_28356,N_28386);
nand U28834 (N_28834,N_28061,N_28317);
or U28835 (N_28835,N_28448,N_28218);
and U28836 (N_28836,N_28351,N_28244);
nand U28837 (N_28837,N_28333,N_28306);
and U28838 (N_28838,N_28426,N_28184);
or U28839 (N_28839,N_28218,N_28489);
and U28840 (N_28840,N_28143,N_28446);
nand U28841 (N_28841,N_28268,N_28313);
or U28842 (N_28842,N_28059,N_28353);
xor U28843 (N_28843,N_28184,N_28322);
nand U28844 (N_28844,N_28151,N_28407);
nor U28845 (N_28845,N_28498,N_28377);
nand U28846 (N_28846,N_28175,N_28020);
xnor U28847 (N_28847,N_28281,N_28088);
nor U28848 (N_28848,N_28443,N_28128);
or U28849 (N_28849,N_28495,N_28275);
nor U28850 (N_28850,N_28049,N_28210);
nor U28851 (N_28851,N_28143,N_28375);
nor U28852 (N_28852,N_28217,N_28299);
xor U28853 (N_28853,N_28154,N_28287);
or U28854 (N_28854,N_28356,N_28347);
nand U28855 (N_28855,N_28148,N_28177);
or U28856 (N_28856,N_28334,N_28146);
xnor U28857 (N_28857,N_28415,N_28002);
and U28858 (N_28858,N_28450,N_28493);
or U28859 (N_28859,N_28498,N_28120);
and U28860 (N_28860,N_28093,N_28021);
and U28861 (N_28861,N_28016,N_28050);
and U28862 (N_28862,N_28186,N_28355);
xor U28863 (N_28863,N_28245,N_28097);
or U28864 (N_28864,N_28459,N_28321);
nor U28865 (N_28865,N_28485,N_28419);
nor U28866 (N_28866,N_28392,N_28288);
xor U28867 (N_28867,N_28476,N_28322);
xor U28868 (N_28868,N_28025,N_28304);
nand U28869 (N_28869,N_28018,N_28288);
xnor U28870 (N_28870,N_28461,N_28170);
xnor U28871 (N_28871,N_28377,N_28338);
nor U28872 (N_28872,N_28138,N_28452);
nand U28873 (N_28873,N_28456,N_28082);
nor U28874 (N_28874,N_28360,N_28221);
or U28875 (N_28875,N_28351,N_28382);
xnor U28876 (N_28876,N_28005,N_28411);
nand U28877 (N_28877,N_28483,N_28325);
and U28878 (N_28878,N_28200,N_28351);
nor U28879 (N_28879,N_28430,N_28388);
nand U28880 (N_28880,N_28138,N_28196);
nand U28881 (N_28881,N_28459,N_28478);
and U28882 (N_28882,N_28427,N_28294);
and U28883 (N_28883,N_28004,N_28317);
nand U28884 (N_28884,N_28244,N_28445);
xor U28885 (N_28885,N_28420,N_28007);
nor U28886 (N_28886,N_28017,N_28403);
nor U28887 (N_28887,N_28467,N_28230);
xnor U28888 (N_28888,N_28216,N_28371);
xnor U28889 (N_28889,N_28376,N_28059);
nor U28890 (N_28890,N_28433,N_28346);
nand U28891 (N_28891,N_28019,N_28390);
nor U28892 (N_28892,N_28247,N_28223);
nand U28893 (N_28893,N_28053,N_28363);
or U28894 (N_28894,N_28432,N_28420);
nor U28895 (N_28895,N_28088,N_28041);
nand U28896 (N_28896,N_28299,N_28197);
and U28897 (N_28897,N_28275,N_28218);
and U28898 (N_28898,N_28369,N_28318);
or U28899 (N_28899,N_28126,N_28467);
and U28900 (N_28900,N_28098,N_28276);
nor U28901 (N_28901,N_28328,N_28002);
xnor U28902 (N_28902,N_28039,N_28223);
nor U28903 (N_28903,N_28178,N_28150);
xnor U28904 (N_28904,N_28102,N_28354);
nor U28905 (N_28905,N_28172,N_28407);
and U28906 (N_28906,N_28442,N_28429);
xnor U28907 (N_28907,N_28196,N_28343);
nand U28908 (N_28908,N_28083,N_28047);
or U28909 (N_28909,N_28441,N_28169);
nor U28910 (N_28910,N_28419,N_28295);
nor U28911 (N_28911,N_28103,N_28100);
or U28912 (N_28912,N_28265,N_28056);
nand U28913 (N_28913,N_28021,N_28141);
and U28914 (N_28914,N_28219,N_28237);
nand U28915 (N_28915,N_28267,N_28470);
xnor U28916 (N_28916,N_28036,N_28116);
nor U28917 (N_28917,N_28358,N_28295);
or U28918 (N_28918,N_28205,N_28444);
nand U28919 (N_28919,N_28014,N_28364);
nor U28920 (N_28920,N_28038,N_28376);
and U28921 (N_28921,N_28241,N_28394);
nor U28922 (N_28922,N_28060,N_28086);
nand U28923 (N_28923,N_28301,N_28484);
nand U28924 (N_28924,N_28112,N_28142);
nor U28925 (N_28925,N_28091,N_28382);
and U28926 (N_28926,N_28421,N_28372);
or U28927 (N_28927,N_28132,N_28431);
and U28928 (N_28928,N_28490,N_28379);
xor U28929 (N_28929,N_28108,N_28113);
or U28930 (N_28930,N_28486,N_28051);
xnor U28931 (N_28931,N_28084,N_28117);
and U28932 (N_28932,N_28296,N_28488);
and U28933 (N_28933,N_28223,N_28497);
nor U28934 (N_28934,N_28172,N_28341);
nor U28935 (N_28935,N_28334,N_28180);
nor U28936 (N_28936,N_28076,N_28240);
or U28937 (N_28937,N_28081,N_28242);
nor U28938 (N_28938,N_28290,N_28348);
nor U28939 (N_28939,N_28201,N_28258);
nand U28940 (N_28940,N_28173,N_28294);
nor U28941 (N_28941,N_28195,N_28055);
nor U28942 (N_28942,N_28260,N_28185);
nand U28943 (N_28943,N_28153,N_28457);
nand U28944 (N_28944,N_28365,N_28148);
or U28945 (N_28945,N_28188,N_28338);
nand U28946 (N_28946,N_28120,N_28185);
or U28947 (N_28947,N_28205,N_28282);
or U28948 (N_28948,N_28265,N_28135);
and U28949 (N_28949,N_28342,N_28214);
nor U28950 (N_28950,N_28375,N_28356);
nor U28951 (N_28951,N_28139,N_28133);
nand U28952 (N_28952,N_28095,N_28012);
nand U28953 (N_28953,N_28300,N_28059);
xor U28954 (N_28954,N_28352,N_28161);
or U28955 (N_28955,N_28431,N_28424);
and U28956 (N_28956,N_28284,N_28399);
xnor U28957 (N_28957,N_28045,N_28363);
xnor U28958 (N_28958,N_28229,N_28297);
or U28959 (N_28959,N_28310,N_28447);
and U28960 (N_28960,N_28225,N_28202);
or U28961 (N_28961,N_28207,N_28020);
xor U28962 (N_28962,N_28237,N_28170);
and U28963 (N_28963,N_28300,N_28423);
or U28964 (N_28964,N_28382,N_28482);
xor U28965 (N_28965,N_28334,N_28227);
and U28966 (N_28966,N_28240,N_28122);
and U28967 (N_28967,N_28196,N_28153);
nor U28968 (N_28968,N_28094,N_28374);
nand U28969 (N_28969,N_28046,N_28123);
xor U28970 (N_28970,N_28020,N_28059);
xnor U28971 (N_28971,N_28250,N_28224);
nor U28972 (N_28972,N_28026,N_28152);
nor U28973 (N_28973,N_28191,N_28303);
xor U28974 (N_28974,N_28202,N_28268);
nand U28975 (N_28975,N_28177,N_28477);
nor U28976 (N_28976,N_28351,N_28234);
nor U28977 (N_28977,N_28369,N_28476);
xnor U28978 (N_28978,N_28410,N_28266);
xnor U28979 (N_28979,N_28224,N_28095);
and U28980 (N_28980,N_28142,N_28123);
nor U28981 (N_28981,N_28355,N_28017);
xor U28982 (N_28982,N_28480,N_28463);
xnor U28983 (N_28983,N_28035,N_28366);
and U28984 (N_28984,N_28053,N_28461);
nor U28985 (N_28985,N_28187,N_28407);
and U28986 (N_28986,N_28037,N_28054);
xor U28987 (N_28987,N_28294,N_28110);
or U28988 (N_28988,N_28391,N_28276);
nor U28989 (N_28989,N_28281,N_28400);
and U28990 (N_28990,N_28282,N_28360);
and U28991 (N_28991,N_28028,N_28180);
and U28992 (N_28992,N_28441,N_28330);
nand U28993 (N_28993,N_28375,N_28323);
and U28994 (N_28994,N_28111,N_28443);
nand U28995 (N_28995,N_28101,N_28116);
nor U28996 (N_28996,N_28475,N_28031);
xnor U28997 (N_28997,N_28430,N_28452);
nand U28998 (N_28998,N_28259,N_28186);
and U28999 (N_28999,N_28320,N_28151);
nor U29000 (N_29000,N_28919,N_28563);
and U29001 (N_29001,N_28577,N_28962);
or U29002 (N_29002,N_28939,N_28782);
xor U29003 (N_29003,N_28602,N_28935);
nand U29004 (N_29004,N_28501,N_28612);
nand U29005 (N_29005,N_28977,N_28908);
nand U29006 (N_29006,N_28837,N_28812);
nand U29007 (N_29007,N_28692,N_28702);
nand U29008 (N_29008,N_28830,N_28661);
nand U29009 (N_29009,N_28701,N_28773);
and U29010 (N_29010,N_28526,N_28504);
or U29011 (N_29011,N_28964,N_28691);
xor U29012 (N_29012,N_28828,N_28776);
nor U29013 (N_29013,N_28804,N_28983);
nand U29014 (N_29014,N_28934,N_28597);
or U29015 (N_29015,N_28646,N_28660);
nand U29016 (N_29016,N_28752,N_28922);
xor U29017 (N_29017,N_28832,N_28751);
nand U29018 (N_29018,N_28936,N_28657);
or U29019 (N_29019,N_28579,N_28860);
and U29020 (N_29020,N_28829,N_28790);
nor U29021 (N_29021,N_28650,N_28547);
xnor U29022 (N_29022,N_28550,N_28627);
xnor U29023 (N_29023,N_28856,N_28861);
and U29024 (N_29024,N_28622,N_28635);
xnor U29025 (N_29025,N_28544,N_28867);
or U29026 (N_29026,N_28823,N_28566);
nor U29027 (N_29027,N_28567,N_28806);
or U29028 (N_29028,N_28619,N_28959);
nand U29029 (N_29029,N_28878,N_28879);
or U29030 (N_29030,N_28899,N_28576);
nand U29031 (N_29031,N_28710,N_28863);
nor U29032 (N_29032,N_28677,N_28531);
xor U29033 (N_29033,N_28881,N_28674);
nor U29034 (N_29034,N_28606,N_28551);
and U29035 (N_29035,N_28523,N_28670);
xor U29036 (N_29036,N_28819,N_28665);
nor U29037 (N_29037,N_28810,N_28872);
nor U29038 (N_29038,N_28673,N_28520);
xor U29039 (N_29039,N_28578,N_28783);
xor U29040 (N_29040,N_28889,N_28689);
or U29041 (N_29041,N_28965,N_28814);
and U29042 (N_29042,N_28958,N_28685);
nor U29043 (N_29043,N_28630,N_28928);
nand U29044 (N_29044,N_28565,N_28847);
nand U29045 (N_29045,N_28900,N_28938);
xnor U29046 (N_29046,N_28641,N_28826);
xor U29047 (N_29047,N_28756,N_28596);
or U29048 (N_29048,N_28754,N_28536);
or U29049 (N_29049,N_28822,N_28880);
nor U29050 (N_29050,N_28791,N_28852);
and U29051 (N_29051,N_28996,N_28690);
and U29052 (N_29052,N_28873,N_28820);
and U29053 (N_29053,N_28686,N_28532);
nand U29054 (N_29054,N_28700,N_28802);
and U29055 (N_29055,N_28877,N_28855);
nor U29056 (N_29056,N_28604,N_28705);
nand U29057 (N_29057,N_28584,N_28594);
or U29058 (N_29058,N_28582,N_28857);
nor U29059 (N_29059,N_28623,N_28628);
xor U29060 (N_29060,N_28666,N_28617);
xnor U29061 (N_29061,N_28683,N_28745);
xnor U29062 (N_29062,N_28981,N_28987);
nor U29063 (N_29063,N_28769,N_28724);
and U29064 (N_29064,N_28771,N_28995);
nand U29065 (N_29065,N_28805,N_28664);
nor U29066 (N_29066,N_28592,N_28795);
nand U29067 (N_29067,N_28868,N_28775);
and U29068 (N_29068,N_28809,N_28985);
nand U29069 (N_29069,N_28718,N_28560);
or U29070 (N_29070,N_28671,N_28957);
and U29071 (N_29071,N_28559,N_28825);
nor U29072 (N_29072,N_28599,N_28748);
nand U29073 (N_29073,N_28510,N_28941);
or U29074 (N_29074,N_28555,N_28815);
or U29075 (N_29075,N_28633,N_28716);
and U29076 (N_29076,N_28763,N_28914);
xor U29077 (N_29077,N_28610,N_28948);
nor U29078 (N_29078,N_28572,N_28731);
or U29079 (N_29079,N_28909,N_28672);
and U29080 (N_29080,N_28961,N_28569);
and U29081 (N_29081,N_28761,N_28758);
or U29082 (N_29082,N_28605,N_28545);
or U29083 (N_29083,N_28695,N_28574);
xor U29084 (N_29084,N_28573,N_28539);
or U29085 (N_29085,N_28858,N_28548);
or U29086 (N_29086,N_28838,N_28854);
xor U29087 (N_29087,N_28946,N_28581);
nor U29088 (N_29088,N_28515,N_28780);
or U29089 (N_29089,N_28750,N_28937);
nor U29090 (N_29090,N_28730,N_28513);
nand U29091 (N_29091,N_28723,N_28557);
xor U29092 (N_29092,N_28912,N_28891);
and U29093 (N_29093,N_28944,N_28918);
and U29094 (N_29094,N_28915,N_28543);
or U29095 (N_29095,N_28570,N_28834);
xnor U29096 (N_29096,N_28765,N_28534);
and U29097 (N_29097,N_28991,N_28926);
nand U29098 (N_29098,N_28675,N_28840);
xnor U29099 (N_29099,N_28580,N_28553);
nand U29100 (N_29100,N_28967,N_28571);
nor U29101 (N_29101,N_28818,N_28933);
nor U29102 (N_29102,N_28801,N_28739);
or U29103 (N_29103,N_28892,N_28652);
xor U29104 (N_29104,N_28629,N_28703);
and U29105 (N_29105,N_28634,N_28921);
and U29106 (N_29106,N_28740,N_28917);
nor U29107 (N_29107,N_28649,N_28757);
nor U29108 (N_29108,N_28653,N_28549);
xnor U29109 (N_29109,N_28713,N_28762);
nor U29110 (N_29110,N_28898,N_28833);
nand U29111 (N_29111,N_28509,N_28800);
and U29112 (N_29112,N_28680,N_28734);
xnor U29113 (N_29113,N_28608,N_28992);
or U29114 (N_29114,N_28799,N_28642);
and U29115 (N_29115,N_28681,N_28621);
nor U29116 (N_29116,N_28506,N_28706);
nand U29117 (N_29117,N_28910,N_28979);
nand U29118 (N_29118,N_28753,N_28853);
xnor U29119 (N_29119,N_28911,N_28647);
nand U29120 (N_29120,N_28907,N_28950);
xnor U29121 (N_29121,N_28960,N_28744);
xor U29122 (N_29122,N_28717,N_28940);
nand U29123 (N_29123,N_28916,N_28888);
nor U29124 (N_29124,N_28742,N_28552);
and U29125 (N_29125,N_28614,N_28698);
or U29126 (N_29126,N_28781,N_28516);
nand U29127 (N_29127,N_28870,N_28732);
or U29128 (N_29128,N_28736,N_28785);
and U29129 (N_29129,N_28986,N_28772);
nand U29130 (N_29130,N_28824,N_28500);
nand U29131 (N_29131,N_28658,N_28639);
xor U29132 (N_29132,N_28601,N_28648);
nor U29133 (N_29133,N_28778,N_28904);
nand U29134 (N_29134,N_28841,N_28827);
xor U29135 (N_29135,N_28529,N_28835);
xor U29136 (N_29136,N_28616,N_28787);
and U29137 (N_29137,N_28583,N_28746);
xnor U29138 (N_29138,N_28722,N_28932);
nor U29139 (N_29139,N_28714,N_28561);
or U29140 (N_29140,N_28659,N_28593);
xnor U29141 (N_29141,N_28786,N_28528);
nand U29142 (N_29142,N_28945,N_28969);
nor U29143 (N_29143,N_28988,N_28953);
nor U29144 (N_29144,N_28848,N_28952);
xor U29145 (N_29145,N_28862,N_28931);
nand U29146 (N_29146,N_28990,N_28808);
and U29147 (N_29147,N_28728,N_28759);
xnor U29148 (N_29148,N_28893,N_28600);
or U29149 (N_29149,N_28951,N_28591);
nand U29150 (N_29150,N_28866,N_28803);
and U29151 (N_29151,N_28788,N_28793);
and U29152 (N_29152,N_28546,N_28792);
nand U29153 (N_29153,N_28954,N_28715);
and U29154 (N_29154,N_28949,N_28844);
nor U29155 (N_29155,N_28760,N_28678);
nand U29156 (N_29156,N_28682,N_28654);
nand U29157 (N_29157,N_28737,N_28625);
nand U29158 (N_29158,N_28874,N_28883);
or U29159 (N_29159,N_28503,N_28514);
nor U29160 (N_29160,N_28568,N_28598);
and U29161 (N_29161,N_28924,N_28846);
nand U29162 (N_29162,N_28684,N_28975);
xnor U29163 (N_29163,N_28517,N_28927);
xnor U29164 (N_29164,N_28699,N_28644);
and U29165 (N_29165,N_28595,N_28632);
or U29166 (N_29166,N_28709,N_28943);
nor U29167 (N_29167,N_28538,N_28743);
nand U29168 (N_29168,N_28807,N_28895);
and U29169 (N_29169,N_28890,N_28735);
or U29170 (N_29170,N_28527,N_28587);
or U29171 (N_29171,N_28925,N_28668);
nand U29172 (N_29172,N_28558,N_28609);
xnor U29173 (N_29173,N_28886,N_28929);
and U29174 (N_29174,N_28956,N_28694);
nor U29175 (N_29175,N_28978,N_28697);
nand U29176 (N_29176,N_28679,N_28966);
and U29177 (N_29177,N_28541,N_28507);
xnor U29178 (N_29178,N_28884,N_28643);
nand U29179 (N_29179,N_28618,N_28817);
nand U29180 (N_29180,N_28947,N_28708);
xnor U29181 (N_29181,N_28511,N_28721);
nor U29182 (N_29182,N_28656,N_28770);
xnor U29183 (N_29183,N_28611,N_28720);
xor U29184 (N_29184,N_28738,N_28796);
and U29185 (N_29185,N_28535,N_28980);
and U29186 (N_29186,N_28859,N_28688);
or U29187 (N_29187,N_28839,N_28725);
nand U29188 (N_29188,N_28747,N_28882);
nand U29189 (N_29189,N_28663,N_28777);
or U29190 (N_29190,N_28850,N_28588);
xnor U29191 (N_29191,N_28849,N_28955);
nand U29192 (N_29192,N_28519,N_28997);
nand U29193 (N_29193,N_28774,N_28667);
nand U29194 (N_29194,N_28971,N_28533);
nand U29195 (N_29195,N_28887,N_28845);
and U29196 (N_29196,N_28537,N_28903);
or U29197 (N_29197,N_28562,N_28590);
nand U29198 (N_29198,N_28631,N_28897);
nand U29199 (N_29199,N_28637,N_28993);
xnor U29200 (N_29200,N_28712,N_28508);
nor U29201 (N_29201,N_28662,N_28586);
or U29202 (N_29202,N_28871,N_28901);
nand U29203 (N_29203,N_28645,N_28896);
xor U29204 (N_29204,N_28972,N_28851);
nand U29205 (N_29205,N_28696,N_28784);
nand U29206 (N_29206,N_28865,N_28726);
and U29207 (N_29207,N_28768,N_28512);
nor U29208 (N_29208,N_28984,N_28755);
xnor U29209 (N_29209,N_28518,N_28963);
nand U29210 (N_29210,N_28651,N_28797);
xnor U29211 (N_29211,N_28970,N_28585);
nand U29212 (N_29212,N_28749,N_28816);
or U29213 (N_29213,N_28974,N_28729);
and U29214 (N_29214,N_28636,N_28811);
and U29215 (N_29215,N_28813,N_28733);
nor U29216 (N_29216,N_28607,N_28556);
or U29217 (N_29217,N_28930,N_28542);
or U29218 (N_29218,N_28779,N_28789);
or U29219 (N_29219,N_28693,N_28913);
nor U29220 (N_29220,N_28505,N_28842);
nand U29221 (N_29221,N_28968,N_28906);
nand U29222 (N_29222,N_28741,N_28766);
nor U29223 (N_29223,N_28836,N_28894);
xor U29224 (N_29224,N_28626,N_28831);
nor U29225 (N_29225,N_28589,N_28976);
and U29226 (N_29226,N_28687,N_28624);
or U29227 (N_29227,N_28994,N_28620);
xor U29228 (N_29228,N_28640,N_28719);
and U29229 (N_29229,N_28821,N_28521);
nand U29230 (N_29230,N_28885,N_28704);
and U29231 (N_29231,N_28942,N_28869);
nor U29232 (N_29232,N_28905,N_28794);
or U29233 (N_29233,N_28676,N_28655);
nor U29234 (N_29234,N_28502,N_28669);
nor U29235 (N_29235,N_28727,N_28999);
nand U29236 (N_29236,N_28989,N_28603);
nor U29237 (N_29237,N_28998,N_28554);
or U29238 (N_29238,N_28613,N_28923);
or U29239 (N_29239,N_28564,N_28876);
nand U29240 (N_29240,N_28575,N_28982);
xnor U29241 (N_29241,N_28638,N_28767);
nand U29242 (N_29242,N_28711,N_28524);
or U29243 (N_29243,N_28707,N_28764);
nor U29244 (N_29244,N_28920,N_28875);
xor U29245 (N_29245,N_28540,N_28530);
and U29246 (N_29246,N_28864,N_28798);
and U29247 (N_29247,N_28525,N_28973);
nor U29248 (N_29248,N_28843,N_28522);
nor U29249 (N_29249,N_28902,N_28615);
and U29250 (N_29250,N_28809,N_28856);
nand U29251 (N_29251,N_28962,N_28805);
nand U29252 (N_29252,N_28821,N_28853);
nor U29253 (N_29253,N_28876,N_28559);
nor U29254 (N_29254,N_28600,N_28566);
or U29255 (N_29255,N_28702,N_28749);
nor U29256 (N_29256,N_28790,N_28945);
or U29257 (N_29257,N_28950,N_28997);
or U29258 (N_29258,N_28517,N_28875);
or U29259 (N_29259,N_28916,N_28992);
and U29260 (N_29260,N_28970,N_28814);
nor U29261 (N_29261,N_28755,N_28718);
xor U29262 (N_29262,N_28752,N_28882);
nor U29263 (N_29263,N_28945,N_28931);
nor U29264 (N_29264,N_28781,N_28627);
xor U29265 (N_29265,N_28862,N_28609);
xnor U29266 (N_29266,N_28527,N_28546);
xnor U29267 (N_29267,N_28533,N_28736);
nand U29268 (N_29268,N_28888,N_28698);
nor U29269 (N_29269,N_28588,N_28787);
nor U29270 (N_29270,N_28983,N_28794);
nand U29271 (N_29271,N_28684,N_28609);
xor U29272 (N_29272,N_28625,N_28551);
nand U29273 (N_29273,N_28951,N_28807);
nor U29274 (N_29274,N_28877,N_28826);
and U29275 (N_29275,N_28587,N_28927);
and U29276 (N_29276,N_28764,N_28712);
and U29277 (N_29277,N_28714,N_28977);
nor U29278 (N_29278,N_28623,N_28674);
nand U29279 (N_29279,N_28871,N_28680);
nand U29280 (N_29280,N_28727,N_28816);
and U29281 (N_29281,N_28513,N_28996);
xnor U29282 (N_29282,N_28620,N_28593);
and U29283 (N_29283,N_28869,N_28719);
or U29284 (N_29284,N_28760,N_28743);
nand U29285 (N_29285,N_28543,N_28678);
nor U29286 (N_29286,N_28879,N_28574);
and U29287 (N_29287,N_28978,N_28673);
nand U29288 (N_29288,N_28649,N_28638);
nor U29289 (N_29289,N_28899,N_28650);
or U29290 (N_29290,N_28622,N_28697);
nor U29291 (N_29291,N_28765,N_28653);
nor U29292 (N_29292,N_28850,N_28683);
xnor U29293 (N_29293,N_28918,N_28755);
xnor U29294 (N_29294,N_28636,N_28973);
or U29295 (N_29295,N_28792,N_28731);
nor U29296 (N_29296,N_28701,N_28767);
nand U29297 (N_29297,N_28612,N_28651);
nand U29298 (N_29298,N_28986,N_28705);
nor U29299 (N_29299,N_28843,N_28678);
nor U29300 (N_29300,N_28580,N_28981);
or U29301 (N_29301,N_28874,N_28766);
nor U29302 (N_29302,N_28933,N_28559);
nor U29303 (N_29303,N_28532,N_28817);
xnor U29304 (N_29304,N_28649,N_28950);
and U29305 (N_29305,N_28978,N_28826);
xor U29306 (N_29306,N_28590,N_28819);
nor U29307 (N_29307,N_28737,N_28728);
and U29308 (N_29308,N_28658,N_28994);
or U29309 (N_29309,N_28563,N_28578);
nor U29310 (N_29310,N_28964,N_28735);
nor U29311 (N_29311,N_28662,N_28675);
nor U29312 (N_29312,N_28822,N_28631);
or U29313 (N_29313,N_28737,N_28572);
and U29314 (N_29314,N_28916,N_28877);
nor U29315 (N_29315,N_28630,N_28809);
xnor U29316 (N_29316,N_28706,N_28913);
nand U29317 (N_29317,N_28607,N_28906);
xor U29318 (N_29318,N_28951,N_28668);
nor U29319 (N_29319,N_28679,N_28816);
nor U29320 (N_29320,N_28805,N_28514);
nand U29321 (N_29321,N_28611,N_28810);
nand U29322 (N_29322,N_28689,N_28542);
or U29323 (N_29323,N_28912,N_28712);
xnor U29324 (N_29324,N_28827,N_28939);
nand U29325 (N_29325,N_28541,N_28636);
xor U29326 (N_29326,N_28722,N_28625);
or U29327 (N_29327,N_28667,N_28936);
xnor U29328 (N_29328,N_28961,N_28970);
nand U29329 (N_29329,N_28690,N_28577);
nand U29330 (N_29330,N_28921,N_28818);
and U29331 (N_29331,N_28689,N_28892);
or U29332 (N_29332,N_28613,N_28904);
or U29333 (N_29333,N_28637,N_28778);
xnor U29334 (N_29334,N_28579,N_28927);
and U29335 (N_29335,N_28842,N_28637);
nand U29336 (N_29336,N_28709,N_28831);
nand U29337 (N_29337,N_28572,N_28591);
or U29338 (N_29338,N_28851,N_28866);
and U29339 (N_29339,N_28652,N_28532);
nand U29340 (N_29340,N_28793,N_28562);
xnor U29341 (N_29341,N_28732,N_28879);
nand U29342 (N_29342,N_28831,N_28896);
xnor U29343 (N_29343,N_28949,N_28582);
or U29344 (N_29344,N_28726,N_28777);
nand U29345 (N_29345,N_28603,N_28578);
xnor U29346 (N_29346,N_28799,N_28981);
nand U29347 (N_29347,N_28772,N_28533);
nor U29348 (N_29348,N_28982,N_28675);
nand U29349 (N_29349,N_28619,N_28850);
nor U29350 (N_29350,N_28843,N_28601);
xnor U29351 (N_29351,N_28524,N_28531);
xor U29352 (N_29352,N_28542,N_28870);
or U29353 (N_29353,N_28626,N_28896);
nand U29354 (N_29354,N_28518,N_28949);
or U29355 (N_29355,N_28710,N_28950);
xor U29356 (N_29356,N_28576,N_28525);
and U29357 (N_29357,N_28699,N_28615);
nor U29358 (N_29358,N_28582,N_28731);
or U29359 (N_29359,N_28750,N_28848);
nor U29360 (N_29360,N_28766,N_28795);
xnor U29361 (N_29361,N_28816,N_28984);
nor U29362 (N_29362,N_28540,N_28753);
nor U29363 (N_29363,N_28530,N_28986);
xor U29364 (N_29364,N_28605,N_28778);
xnor U29365 (N_29365,N_28509,N_28948);
xnor U29366 (N_29366,N_28621,N_28997);
xor U29367 (N_29367,N_28817,N_28928);
xor U29368 (N_29368,N_28891,N_28549);
or U29369 (N_29369,N_28849,N_28665);
xnor U29370 (N_29370,N_28502,N_28531);
xor U29371 (N_29371,N_28731,N_28877);
nor U29372 (N_29372,N_28896,N_28894);
and U29373 (N_29373,N_28750,N_28519);
and U29374 (N_29374,N_28678,N_28579);
nand U29375 (N_29375,N_28777,N_28826);
or U29376 (N_29376,N_28908,N_28843);
nand U29377 (N_29377,N_28973,N_28830);
nand U29378 (N_29378,N_28648,N_28785);
and U29379 (N_29379,N_28835,N_28594);
nand U29380 (N_29380,N_28524,N_28663);
nand U29381 (N_29381,N_28908,N_28633);
nor U29382 (N_29382,N_28958,N_28971);
or U29383 (N_29383,N_28938,N_28905);
nand U29384 (N_29384,N_28873,N_28603);
and U29385 (N_29385,N_28967,N_28932);
or U29386 (N_29386,N_28881,N_28525);
nor U29387 (N_29387,N_28655,N_28557);
and U29388 (N_29388,N_28581,N_28659);
nand U29389 (N_29389,N_28624,N_28656);
and U29390 (N_29390,N_28548,N_28844);
nor U29391 (N_29391,N_28547,N_28995);
nor U29392 (N_29392,N_28706,N_28821);
and U29393 (N_29393,N_28942,N_28976);
nand U29394 (N_29394,N_28930,N_28869);
or U29395 (N_29395,N_28521,N_28875);
or U29396 (N_29396,N_28874,N_28672);
xnor U29397 (N_29397,N_28785,N_28587);
and U29398 (N_29398,N_28590,N_28523);
nor U29399 (N_29399,N_28931,N_28528);
or U29400 (N_29400,N_28895,N_28771);
nand U29401 (N_29401,N_28544,N_28621);
or U29402 (N_29402,N_28577,N_28770);
and U29403 (N_29403,N_28792,N_28990);
nand U29404 (N_29404,N_28845,N_28972);
nor U29405 (N_29405,N_28571,N_28545);
nand U29406 (N_29406,N_28830,N_28665);
nand U29407 (N_29407,N_28737,N_28618);
xor U29408 (N_29408,N_28666,N_28630);
and U29409 (N_29409,N_28988,N_28838);
or U29410 (N_29410,N_28622,N_28704);
or U29411 (N_29411,N_28948,N_28934);
nor U29412 (N_29412,N_28877,N_28729);
nor U29413 (N_29413,N_28736,N_28720);
nor U29414 (N_29414,N_28746,N_28560);
or U29415 (N_29415,N_28798,N_28548);
nor U29416 (N_29416,N_28640,N_28725);
nand U29417 (N_29417,N_28642,N_28789);
or U29418 (N_29418,N_28593,N_28561);
nand U29419 (N_29419,N_28860,N_28656);
or U29420 (N_29420,N_28934,N_28908);
and U29421 (N_29421,N_28579,N_28707);
and U29422 (N_29422,N_28671,N_28940);
or U29423 (N_29423,N_28860,N_28649);
and U29424 (N_29424,N_28823,N_28766);
nor U29425 (N_29425,N_28811,N_28855);
xor U29426 (N_29426,N_28654,N_28626);
xnor U29427 (N_29427,N_28740,N_28779);
nand U29428 (N_29428,N_28985,N_28951);
or U29429 (N_29429,N_28661,N_28925);
or U29430 (N_29430,N_28676,N_28986);
xnor U29431 (N_29431,N_28761,N_28664);
and U29432 (N_29432,N_28654,N_28824);
nand U29433 (N_29433,N_28964,N_28591);
or U29434 (N_29434,N_28849,N_28707);
nand U29435 (N_29435,N_28915,N_28940);
xnor U29436 (N_29436,N_28534,N_28734);
or U29437 (N_29437,N_28679,N_28544);
or U29438 (N_29438,N_28530,N_28919);
nor U29439 (N_29439,N_28911,N_28983);
xor U29440 (N_29440,N_28918,N_28745);
and U29441 (N_29441,N_28919,N_28837);
and U29442 (N_29442,N_28579,N_28590);
or U29443 (N_29443,N_28792,N_28836);
nand U29444 (N_29444,N_28740,N_28777);
or U29445 (N_29445,N_28560,N_28934);
and U29446 (N_29446,N_28895,N_28676);
and U29447 (N_29447,N_28663,N_28884);
nor U29448 (N_29448,N_28765,N_28999);
nor U29449 (N_29449,N_28907,N_28741);
or U29450 (N_29450,N_28692,N_28727);
nand U29451 (N_29451,N_28719,N_28900);
xor U29452 (N_29452,N_28564,N_28825);
nor U29453 (N_29453,N_28849,N_28765);
nor U29454 (N_29454,N_28880,N_28757);
xor U29455 (N_29455,N_28692,N_28967);
or U29456 (N_29456,N_28896,N_28818);
nor U29457 (N_29457,N_28638,N_28737);
nor U29458 (N_29458,N_28759,N_28925);
xnor U29459 (N_29459,N_28573,N_28789);
and U29460 (N_29460,N_28882,N_28875);
nor U29461 (N_29461,N_28681,N_28914);
or U29462 (N_29462,N_28946,N_28550);
nand U29463 (N_29463,N_28564,N_28703);
nand U29464 (N_29464,N_28939,N_28803);
nor U29465 (N_29465,N_28643,N_28645);
or U29466 (N_29466,N_28547,N_28745);
nand U29467 (N_29467,N_28957,N_28985);
nor U29468 (N_29468,N_28765,N_28987);
or U29469 (N_29469,N_28563,N_28903);
and U29470 (N_29470,N_28919,N_28676);
xnor U29471 (N_29471,N_28733,N_28705);
and U29472 (N_29472,N_28858,N_28957);
and U29473 (N_29473,N_28917,N_28559);
xnor U29474 (N_29474,N_28621,N_28683);
nor U29475 (N_29475,N_28724,N_28941);
xor U29476 (N_29476,N_28881,N_28789);
nand U29477 (N_29477,N_28543,N_28557);
or U29478 (N_29478,N_28996,N_28843);
and U29479 (N_29479,N_28931,N_28933);
nor U29480 (N_29480,N_28900,N_28560);
or U29481 (N_29481,N_28545,N_28705);
or U29482 (N_29482,N_28961,N_28924);
nand U29483 (N_29483,N_28849,N_28551);
or U29484 (N_29484,N_28586,N_28806);
xnor U29485 (N_29485,N_28603,N_28703);
and U29486 (N_29486,N_28968,N_28519);
xnor U29487 (N_29487,N_28869,N_28713);
xnor U29488 (N_29488,N_28917,N_28653);
nand U29489 (N_29489,N_28980,N_28799);
or U29490 (N_29490,N_28532,N_28940);
nor U29491 (N_29491,N_28512,N_28678);
or U29492 (N_29492,N_28995,N_28879);
nor U29493 (N_29493,N_28792,N_28671);
xnor U29494 (N_29494,N_28520,N_28630);
nor U29495 (N_29495,N_28946,N_28768);
xnor U29496 (N_29496,N_28592,N_28551);
or U29497 (N_29497,N_28635,N_28842);
nand U29498 (N_29498,N_28731,N_28574);
xnor U29499 (N_29499,N_28948,N_28914);
or U29500 (N_29500,N_29281,N_29486);
or U29501 (N_29501,N_29349,N_29095);
nor U29502 (N_29502,N_29037,N_29490);
nor U29503 (N_29503,N_29260,N_29302);
or U29504 (N_29504,N_29307,N_29033);
and U29505 (N_29505,N_29227,N_29136);
nand U29506 (N_29506,N_29419,N_29259);
nor U29507 (N_29507,N_29323,N_29380);
or U29508 (N_29508,N_29097,N_29296);
and U29509 (N_29509,N_29241,N_29014);
and U29510 (N_29510,N_29476,N_29204);
and U29511 (N_29511,N_29129,N_29447);
and U29512 (N_29512,N_29218,N_29466);
and U29513 (N_29513,N_29000,N_29454);
or U29514 (N_29514,N_29190,N_29305);
or U29515 (N_29515,N_29107,N_29217);
xnor U29516 (N_29516,N_29406,N_29461);
or U29517 (N_29517,N_29038,N_29261);
nor U29518 (N_29518,N_29079,N_29184);
or U29519 (N_29519,N_29155,N_29188);
nor U29520 (N_29520,N_29379,N_29146);
or U29521 (N_29521,N_29298,N_29243);
or U29522 (N_29522,N_29437,N_29424);
xor U29523 (N_29523,N_29220,N_29099);
or U29524 (N_29524,N_29224,N_29057);
nor U29525 (N_29525,N_29264,N_29026);
nand U29526 (N_29526,N_29032,N_29169);
nand U29527 (N_29527,N_29414,N_29101);
nand U29528 (N_29528,N_29374,N_29131);
xnor U29529 (N_29529,N_29276,N_29152);
and U29530 (N_29530,N_29211,N_29321);
nor U29531 (N_29531,N_29130,N_29340);
nand U29532 (N_29532,N_29334,N_29090);
nor U29533 (N_29533,N_29159,N_29103);
nand U29534 (N_29534,N_29157,N_29358);
and U29535 (N_29535,N_29207,N_29128);
and U29536 (N_29536,N_29392,N_29044);
or U29537 (N_29537,N_29285,N_29408);
or U29538 (N_29538,N_29343,N_29435);
and U29539 (N_29539,N_29096,N_29463);
xnor U29540 (N_29540,N_29470,N_29077);
nor U29541 (N_29541,N_29117,N_29040);
xor U29542 (N_29542,N_29402,N_29138);
and U29543 (N_29543,N_29072,N_29456);
and U29544 (N_29544,N_29127,N_29059);
xnor U29545 (N_29545,N_29313,N_29240);
nor U29546 (N_29546,N_29052,N_29479);
or U29547 (N_29547,N_29233,N_29303);
and U29548 (N_29548,N_29208,N_29335);
xnor U29549 (N_29549,N_29404,N_29371);
and U29550 (N_29550,N_29398,N_29194);
or U29551 (N_29551,N_29306,N_29149);
nor U29552 (N_29552,N_29308,N_29082);
nor U29553 (N_29553,N_29247,N_29473);
nor U29554 (N_29554,N_29314,N_29137);
or U29555 (N_29555,N_29439,N_29248);
nand U29556 (N_29556,N_29265,N_29327);
xnor U29557 (N_29557,N_29223,N_29244);
xor U29558 (N_29558,N_29141,N_29168);
and U29559 (N_29559,N_29142,N_29186);
or U29560 (N_29560,N_29332,N_29199);
or U29561 (N_29561,N_29464,N_29198);
nand U29562 (N_29562,N_29140,N_29451);
nand U29563 (N_29563,N_29200,N_29460);
nor U29564 (N_29564,N_29375,N_29106);
or U29565 (N_29565,N_29084,N_29287);
nor U29566 (N_29566,N_29145,N_29295);
or U29567 (N_29567,N_29354,N_29093);
or U29568 (N_29568,N_29029,N_29377);
nor U29569 (N_29569,N_29187,N_29412);
and U29570 (N_29570,N_29267,N_29489);
or U29571 (N_29571,N_29094,N_29177);
nor U29572 (N_29572,N_29448,N_29368);
nand U29573 (N_29573,N_29274,N_29042);
xnor U29574 (N_29574,N_29030,N_29309);
nand U29575 (N_29575,N_29041,N_29023);
nand U29576 (N_29576,N_29280,N_29139);
nor U29577 (N_29577,N_29221,N_29469);
or U29578 (N_29578,N_29191,N_29425);
nor U29579 (N_29579,N_29182,N_29495);
or U29580 (N_29580,N_29318,N_29053);
or U29581 (N_29581,N_29143,N_29273);
or U29582 (N_29582,N_29232,N_29108);
xor U29583 (N_29583,N_29115,N_29331);
nand U29584 (N_29584,N_29234,N_29381);
and U29585 (N_29585,N_29058,N_29284);
xor U29586 (N_29586,N_29409,N_29089);
or U29587 (N_29587,N_29201,N_29269);
nor U29588 (N_29588,N_29275,N_29403);
xor U29589 (N_29589,N_29474,N_29125);
or U29590 (N_29590,N_29337,N_29468);
nor U29591 (N_29591,N_29205,N_29440);
or U29592 (N_29592,N_29283,N_29310);
and U29593 (N_29593,N_29317,N_29166);
nor U29594 (N_29594,N_29135,N_29452);
or U29595 (N_29595,N_29016,N_29076);
xor U29596 (N_29596,N_29299,N_29005);
or U29597 (N_29597,N_29329,N_29423);
and U29598 (N_29598,N_29213,N_29121);
xor U29599 (N_29599,N_29181,N_29228);
and U29600 (N_29600,N_29104,N_29258);
nor U29601 (N_29601,N_29399,N_29055);
and U29602 (N_29602,N_29382,N_29420);
or U29603 (N_29603,N_29214,N_29178);
and U29604 (N_29604,N_29278,N_29304);
and U29605 (N_29605,N_29075,N_29286);
xor U29606 (N_29606,N_29158,N_29475);
xnor U29607 (N_29607,N_29297,N_29415);
xnor U29608 (N_29608,N_29002,N_29396);
nand U29609 (N_29609,N_29039,N_29235);
nand U29610 (N_29610,N_29179,N_29036);
or U29611 (N_29611,N_29357,N_29443);
or U29612 (N_29612,N_29362,N_29065);
xnor U29613 (N_29613,N_29345,N_29197);
nand U29614 (N_29614,N_29373,N_29134);
and U29615 (N_29615,N_29338,N_29458);
nand U29616 (N_29616,N_29395,N_29153);
xnor U29617 (N_29617,N_29092,N_29459);
and U29618 (N_29618,N_29416,N_29301);
xor U29619 (N_29619,N_29432,N_29256);
and U29620 (N_29620,N_29118,N_29352);
nand U29621 (N_29621,N_29100,N_29427);
and U29622 (N_29622,N_29480,N_29497);
or U29623 (N_29623,N_29193,N_29110);
nand U29624 (N_29624,N_29262,N_29066);
or U29625 (N_29625,N_29422,N_29027);
xor U29626 (N_29626,N_29291,N_29342);
nor U29627 (N_29627,N_29124,N_29325);
or U29628 (N_29628,N_29481,N_29315);
or U29629 (N_29629,N_29351,N_29434);
nor U29630 (N_29630,N_29133,N_29102);
or U29631 (N_29631,N_29483,N_29359);
nor U29632 (N_29632,N_29383,N_29418);
xnor U29633 (N_29633,N_29087,N_29226);
or U29634 (N_29634,N_29252,N_29421);
nand U29635 (N_29635,N_29341,N_29477);
or U29636 (N_29636,N_29031,N_29405);
or U29637 (N_29637,N_29161,N_29492);
or U29638 (N_29638,N_29189,N_29018);
nor U29639 (N_29639,N_29230,N_29484);
and U29640 (N_29640,N_29339,N_29071);
or U29641 (N_29641,N_29330,N_29068);
nand U29642 (N_29642,N_29385,N_29455);
and U29643 (N_29643,N_29450,N_29070);
nor U29644 (N_29644,N_29147,N_29263);
xnor U29645 (N_29645,N_29001,N_29022);
and U29646 (N_29646,N_29144,N_29289);
nor U29647 (N_29647,N_29431,N_29063);
and U29648 (N_29648,N_29397,N_29465);
or U29649 (N_29649,N_29328,N_29320);
xor U29650 (N_29650,N_29246,N_29078);
nor U29651 (N_29651,N_29237,N_29245);
xnor U29652 (N_29652,N_29206,N_29113);
or U29653 (N_29653,N_29098,N_29360);
nor U29654 (N_29654,N_29433,N_29255);
or U29655 (N_29655,N_29498,N_29294);
xnor U29656 (N_29656,N_29012,N_29279);
or U29657 (N_29657,N_29156,N_29319);
and U29658 (N_29658,N_29061,N_29024);
nor U29659 (N_29659,N_29438,N_29088);
and U29660 (N_29660,N_29292,N_29457);
nand U29661 (N_29661,N_29196,N_29391);
xnor U29662 (N_29662,N_29364,N_29048);
nand U29663 (N_29663,N_29311,N_29444);
and U29664 (N_29664,N_29407,N_29290);
nor U29665 (N_29665,N_29148,N_29046);
and U29666 (N_29666,N_29499,N_29333);
xnor U29667 (N_29667,N_29192,N_29366);
nand U29668 (N_29668,N_29253,N_29344);
nor U29669 (N_29669,N_29176,N_29154);
or U29670 (N_29670,N_29049,N_29160);
nor U29671 (N_29671,N_29185,N_29047);
nand U29672 (N_29672,N_29293,N_29449);
nand U29673 (N_29673,N_29180,N_29060);
or U29674 (N_29674,N_29170,N_29426);
nand U29675 (N_29675,N_29111,N_29015);
nor U29676 (N_29676,N_29011,N_29347);
nand U29677 (N_29677,N_29355,N_29043);
nand U29678 (N_29678,N_29203,N_29250);
or U29679 (N_29679,N_29493,N_29056);
nor U29680 (N_29680,N_29394,N_29288);
xnor U29681 (N_29681,N_29091,N_29085);
nor U29682 (N_29682,N_29209,N_29120);
and U29683 (N_29683,N_29163,N_29277);
nor U29684 (N_29684,N_29312,N_29123);
xnor U29685 (N_29685,N_29478,N_29080);
xor U29686 (N_29686,N_29105,N_29150);
nor U29687 (N_29687,N_29050,N_29491);
nand U29688 (N_29688,N_29367,N_29035);
nand U29689 (N_29689,N_29257,N_29471);
or U29690 (N_29690,N_29238,N_29054);
nand U29691 (N_29691,N_29013,N_29009);
nor U29692 (N_29692,N_29212,N_29174);
xor U29693 (N_29693,N_29034,N_29282);
nor U29694 (N_29694,N_29175,N_29376);
nand U29695 (N_29695,N_29442,N_29219);
nor U29696 (N_29696,N_29073,N_29485);
and U29697 (N_29697,N_29172,N_29430);
nand U29698 (N_29698,N_29112,N_29010);
nor U29699 (N_29699,N_29370,N_29350);
or U29700 (N_29700,N_29028,N_29114);
nand U29701 (N_29701,N_29271,N_29231);
xor U29702 (N_29702,N_29361,N_29007);
or U29703 (N_29703,N_29401,N_29249);
nor U29704 (N_29704,N_29369,N_29020);
nor U29705 (N_29705,N_29215,N_29126);
or U29706 (N_29706,N_29062,N_29348);
nand U29707 (N_29707,N_29216,N_29356);
nand U29708 (N_29708,N_29006,N_29239);
nor U29709 (N_29709,N_29109,N_29446);
xnor U29710 (N_29710,N_29270,N_29482);
nor U29711 (N_29711,N_29171,N_29004);
xor U29712 (N_29712,N_29428,N_29389);
nand U29713 (N_29713,N_29336,N_29487);
nor U29714 (N_29714,N_29167,N_29324);
or U29715 (N_29715,N_29225,N_29393);
nand U29716 (N_29716,N_29202,N_29019);
xor U29717 (N_29717,N_29086,N_29467);
xnor U29718 (N_29718,N_29064,N_29173);
nand U29719 (N_29719,N_29122,N_29021);
and U29720 (N_29720,N_29045,N_29183);
and U29721 (N_29721,N_29413,N_29496);
nand U29722 (N_29722,N_29008,N_29210);
nand U29723 (N_29723,N_29411,N_29378);
and U29724 (N_29724,N_29363,N_29229);
and U29725 (N_29725,N_29453,N_29195);
xor U29726 (N_29726,N_29488,N_29119);
xor U29727 (N_29727,N_29387,N_29472);
nor U29728 (N_29728,N_29436,N_29417);
xnor U29729 (N_29729,N_29164,N_29372);
and U29730 (N_29730,N_29116,N_29326);
xor U29731 (N_29731,N_29242,N_29390);
or U29732 (N_29732,N_29165,N_29222);
nor U29733 (N_29733,N_29462,N_29272);
or U29734 (N_29734,N_29236,N_29074);
nor U29735 (N_29735,N_29441,N_29445);
or U29736 (N_29736,N_29322,N_29300);
xor U29737 (N_29737,N_29083,N_29025);
nor U29738 (N_29738,N_29268,N_29386);
xnor U29739 (N_29739,N_29132,N_29410);
nand U29740 (N_29740,N_29003,N_29081);
and U29741 (N_29741,N_29400,N_29069);
nand U29742 (N_29742,N_29067,N_29346);
or U29743 (N_29743,N_29254,N_29251);
nand U29744 (N_29744,N_29151,N_29429);
or U29745 (N_29745,N_29388,N_29162);
nand U29746 (N_29746,N_29051,N_29316);
xnor U29747 (N_29747,N_29017,N_29384);
xnor U29748 (N_29748,N_29266,N_29494);
xor U29749 (N_29749,N_29353,N_29365);
or U29750 (N_29750,N_29282,N_29347);
nand U29751 (N_29751,N_29459,N_29001);
nand U29752 (N_29752,N_29472,N_29199);
nand U29753 (N_29753,N_29167,N_29115);
and U29754 (N_29754,N_29078,N_29378);
xnor U29755 (N_29755,N_29223,N_29467);
nand U29756 (N_29756,N_29286,N_29283);
or U29757 (N_29757,N_29426,N_29497);
or U29758 (N_29758,N_29214,N_29423);
nor U29759 (N_29759,N_29413,N_29211);
or U29760 (N_29760,N_29236,N_29362);
and U29761 (N_29761,N_29369,N_29033);
nand U29762 (N_29762,N_29111,N_29216);
and U29763 (N_29763,N_29133,N_29031);
or U29764 (N_29764,N_29032,N_29057);
nor U29765 (N_29765,N_29496,N_29364);
and U29766 (N_29766,N_29072,N_29166);
nand U29767 (N_29767,N_29318,N_29106);
xor U29768 (N_29768,N_29416,N_29421);
or U29769 (N_29769,N_29485,N_29166);
nor U29770 (N_29770,N_29314,N_29148);
nor U29771 (N_29771,N_29094,N_29432);
and U29772 (N_29772,N_29382,N_29464);
nand U29773 (N_29773,N_29349,N_29144);
and U29774 (N_29774,N_29424,N_29400);
and U29775 (N_29775,N_29380,N_29061);
and U29776 (N_29776,N_29099,N_29177);
or U29777 (N_29777,N_29338,N_29224);
nor U29778 (N_29778,N_29417,N_29001);
or U29779 (N_29779,N_29348,N_29434);
nor U29780 (N_29780,N_29422,N_29053);
or U29781 (N_29781,N_29030,N_29217);
or U29782 (N_29782,N_29492,N_29210);
or U29783 (N_29783,N_29216,N_29014);
nor U29784 (N_29784,N_29438,N_29334);
nand U29785 (N_29785,N_29023,N_29311);
and U29786 (N_29786,N_29179,N_29020);
nor U29787 (N_29787,N_29183,N_29109);
and U29788 (N_29788,N_29072,N_29178);
xor U29789 (N_29789,N_29002,N_29307);
or U29790 (N_29790,N_29321,N_29347);
nor U29791 (N_29791,N_29036,N_29213);
or U29792 (N_29792,N_29243,N_29138);
nor U29793 (N_29793,N_29075,N_29018);
and U29794 (N_29794,N_29101,N_29253);
nor U29795 (N_29795,N_29242,N_29148);
nand U29796 (N_29796,N_29318,N_29460);
xor U29797 (N_29797,N_29372,N_29326);
and U29798 (N_29798,N_29282,N_29459);
xnor U29799 (N_29799,N_29207,N_29453);
nand U29800 (N_29800,N_29242,N_29108);
nor U29801 (N_29801,N_29164,N_29028);
or U29802 (N_29802,N_29122,N_29166);
nand U29803 (N_29803,N_29254,N_29011);
nor U29804 (N_29804,N_29151,N_29419);
xor U29805 (N_29805,N_29146,N_29316);
and U29806 (N_29806,N_29203,N_29242);
and U29807 (N_29807,N_29160,N_29434);
nand U29808 (N_29808,N_29383,N_29024);
nand U29809 (N_29809,N_29000,N_29470);
and U29810 (N_29810,N_29471,N_29327);
or U29811 (N_29811,N_29422,N_29067);
or U29812 (N_29812,N_29325,N_29481);
xor U29813 (N_29813,N_29126,N_29179);
nor U29814 (N_29814,N_29185,N_29209);
nor U29815 (N_29815,N_29434,N_29239);
nor U29816 (N_29816,N_29098,N_29058);
nand U29817 (N_29817,N_29427,N_29199);
or U29818 (N_29818,N_29298,N_29494);
and U29819 (N_29819,N_29334,N_29201);
xor U29820 (N_29820,N_29127,N_29181);
nor U29821 (N_29821,N_29343,N_29336);
or U29822 (N_29822,N_29238,N_29325);
and U29823 (N_29823,N_29229,N_29220);
and U29824 (N_29824,N_29219,N_29159);
xor U29825 (N_29825,N_29484,N_29004);
nor U29826 (N_29826,N_29192,N_29094);
and U29827 (N_29827,N_29275,N_29482);
xor U29828 (N_29828,N_29229,N_29366);
nand U29829 (N_29829,N_29261,N_29264);
nand U29830 (N_29830,N_29174,N_29202);
or U29831 (N_29831,N_29296,N_29243);
xor U29832 (N_29832,N_29044,N_29174);
or U29833 (N_29833,N_29476,N_29399);
nand U29834 (N_29834,N_29460,N_29410);
nor U29835 (N_29835,N_29384,N_29391);
nor U29836 (N_29836,N_29463,N_29031);
xor U29837 (N_29837,N_29164,N_29205);
or U29838 (N_29838,N_29322,N_29099);
xnor U29839 (N_29839,N_29140,N_29436);
or U29840 (N_29840,N_29075,N_29200);
nor U29841 (N_29841,N_29274,N_29072);
nand U29842 (N_29842,N_29103,N_29376);
and U29843 (N_29843,N_29120,N_29485);
and U29844 (N_29844,N_29189,N_29354);
xor U29845 (N_29845,N_29158,N_29275);
nor U29846 (N_29846,N_29245,N_29231);
nor U29847 (N_29847,N_29244,N_29207);
nor U29848 (N_29848,N_29378,N_29005);
xor U29849 (N_29849,N_29152,N_29314);
and U29850 (N_29850,N_29081,N_29089);
xnor U29851 (N_29851,N_29307,N_29001);
or U29852 (N_29852,N_29091,N_29397);
nand U29853 (N_29853,N_29014,N_29126);
nor U29854 (N_29854,N_29115,N_29326);
nand U29855 (N_29855,N_29462,N_29498);
and U29856 (N_29856,N_29317,N_29029);
nand U29857 (N_29857,N_29441,N_29053);
xnor U29858 (N_29858,N_29116,N_29265);
and U29859 (N_29859,N_29287,N_29142);
and U29860 (N_29860,N_29195,N_29412);
xor U29861 (N_29861,N_29030,N_29154);
nor U29862 (N_29862,N_29288,N_29174);
nand U29863 (N_29863,N_29289,N_29238);
xnor U29864 (N_29864,N_29345,N_29120);
xor U29865 (N_29865,N_29440,N_29208);
nor U29866 (N_29866,N_29218,N_29246);
and U29867 (N_29867,N_29215,N_29112);
and U29868 (N_29868,N_29281,N_29470);
and U29869 (N_29869,N_29077,N_29118);
nand U29870 (N_29870,N_29467,N_29091);
or U29871 (N_29871,N_29278,N_29249);
nor U29872 (N_29872,N_29160,N_29146);
xor U29873 (N_29873,N_29495,N_29383);
xor U29874 (N_29874,N_29123,N_29489);
and U29875 (N_29875,N_29124,N_29265);
nor U29876 (N_29876,N_29288,N_29002);
xor U29877 (N_29877,N_29102,N_29359);
nor U29878 (N_29878,N_29395,N_29164);
or U29879 (N_29879,N_29377,N_29497);
nand U29880 (N_29880,N_29484,N_29025);
or U29881 (N_29881,N_29126,N_29463);
and U29882 (N_29882,N_29475,N_29001);
nand U29883 (N_29883,N_29066,N_29168);
nor U29884 (N_29884,N_29412,N_29154);
nor U29885 (N_29885,N_29342,N_29078);
nand U29886 (N_29886,N_29421,N_29186);
nor U29887 (N_29887,N_29336,N_29294);
nand U29888 (N_29888,N_29042,N_29196);
nand U29889 (N_29889,N_29328,N_29369);
and U29890 (N_29890,N_29263,N_29156);
nor U29891 (N_29891,N_29158,N_29232);
or U29892 (N_29892,N_29443,N_29311);
nor U29893 (N_29893,N_29145,N_29429);
xnor U29894 (N_29894,N_29043,N_29494);
nand U29895 (N_29895,N_29458,N_29098);
or U29896 (N_29896,N_29484,N_29254);
xnor U29897 (N_29897,N_29334,N_29278);
xor U29898 (N_29898,N_29303,N_29321);
xnor U29899 (N_29899,N_29120,N_29048);
nand U29900 (N_29900,N_29317,N_29400);
xor U29901 (N_29901,N_29097,N_29361);
and U29902 (N_29902,N_29111,N_29466);
nand U29903 (N_29903,N_29269,N_29073);
nand U29904 (N_29904,N_29205,N_29352);
nor U29905 (N_29905,N_29063,N_29026);
xor U29906 (N_29906,N_29148,N_29029);
and U29907 (N_29907,N_29453,N_29051);
or U29908 (N_29908,N_29045,N_29433);
xnor U29909 (N_29909,N_29467,N_29364);
and U29910 (N_29910,N_29111,N_29152);
nand U29911 (N_29911,N_29405,N_29163);
and U29912 (N_29912,N_29313,N_29058);
or U29913 (N_29913,N_29128,N_29482);
nand U29914 (N_29914,N_29051,N_29447);
or U29915 (N_29915,N_29493,N_29482);
xnor U29916 (N_29916,N_29451,N_29251);
nand U29917 (N_29917,N_29262,N_29095);
nor U29918 (N_29918,N_29288,N_29032);
or U29919 (N_29919,N_29049,N_29342);
or U29920 (N_29920,N_29085,N_29128);
or U29921 (N_29921,N_29323,N_29257);
and U29922 (N_29922,N_29274,N_29077);
nor U29923 (N_29923,N_29160,N_29446);
nand U29924 (N_29924,N_29014,N_29155);
nand U29925 (N_29925,N_29420,N_29031);
xnor U29926 (N_29926,N_29061,N_29498);
xnor U29927 (N_29927,N_29073,N_29473);
nor U29928 (N_29928,N_29463,N_29475);
nor U29929 (N_29929,N_29339,N_29489);
or U29930 (N_29930,N_29126,N_29480);
nand U29931 (N_29931,N_29082,N_29140);
and U29932 (N_29932,N_29093,N_29197);
nor U29933 (N_29933,N_29338,N_29388);
nand U29934 (N_29934,N_29448,N_29295);
nand U29935 (N_29935,N_29474,N_29497);
nand U29936 (N_29936,N_29451,N_29003);
nor U29937 (N_29937,N_29162,N_29305);
nor U29938 (N_29938,N_29048,N_29486);
and U29939 (N_29939,N_29391,N_29105);
or U29940 (N_29940,N_29317,N_29190);
or U29941 (N_29941,N_29129,N_29060);
or U29942 (N_29942,N_29287,N_29124);
xnor U29943 (N_29943,N_29474,N_29088);
and U29944 (N_29944,N_29359,N_29028);
and U29945 (N_29945,N_29050,N_29208);
xor U29946 (N_29946,N_29274,N_29132);
xnor U29947 (N_29947,N_29449,N_29361);
nand U29948 (N_29948,N_29427,N_29262);
xor U29949 (N_29949,N_29233,N_29446);
nor U29950 (N_29950,N_29224,N_29436);
nor U29951 (N_29951,N_29045,N_29429);
nand U29952 (N_29952,N_29364,N_29213);
nand U29953 (N_29953,N_29141,N_29425);
and U29954 (N_29954,N_29463,N_29471);
nor U29955 (N_29955,N_29335,N_29072);
and U29956 (N_29956,N_29467,N_29151);
nand U29957 (N_29957,N_29286,N_29064);
nor U29958 (N_29958,N_29487,N_29022);
nand U29959 (N_29959,N_29246,N_29436);
nand U29960 (N_29960,N_29477,N_29438);
xor U29961 (N_29961,N_29185,N_29138);
and U29962 (N_29962,N_29227,N_29412);
xnor U29963 (N_29963,N_29308,N_29330);
and U29964 (N_29964,N_29267,N_29132);
nor U29965 (N_29965,N_29491,N_29403);
nand U29966 (N_29966,N_29297,N_29237);
nand U29967 (N_29967,N_29019,N_29280);
or U29968 (N_29968,N_29217,N_29091);
nor U29969 (N_29969,N_29271,N_29215);
or U29970 (N_29970,N_29383,N_29189);
and U29971 (N_29971,N_29346,N_29070);
nor U29972 (N_29972,N_29167,N_29425);
nor U29973 (N_29973,N_29464,N_29389);
xor U29974 (N_29974,N_29136,N_29316);
xnor U29975 (N_29975,N_29105,N_29134);
xor U29976 (N_29976,N_29330,N_29053);
xnor U29977 (N_29977,N_29082,N_29187);
and U29978 (N_29978,N_29112,N_29003);
or U29979 (N_29979,N_29478,N_29332);
xor U29980 (N_29980,N_29185,N_29487);
or U29981 (N_29981,N_29318,N_29181);
or U29982 (N_29982,N_29142,N_29439);
nand U29983 (N_29983,N_29117,N_29470);
or U29984 (N_29984,N_29043,N_29174);
or U29985 (N_29985,N_29403,N_29037);
or U29986 (N_29986,N_29385,N_29318);
or U29987 (N_29987,N_29088,N_29019);
or U29988 (N_29988,N_29023,N_29037);
or U29989 (N_29989,N_29319,N_29392);
or U29990 (N_29990,N_29225,N_29254);
nor U29991 (N_29991,N_29365,N_29445);
nand U29992 (N_29992,N_29015,N_29156);
xnor U29993 (N_29993,N_29438,N_29451);
xnor U29994 (N_29994,N_29080,N_29150);
nand U29995 (N_29995,N_29355,N_29472);
nand U29996 (N_29996,N_29073,N_29317);
and U29997 (N_29997,N_29497,N_29077);
xnor U29998 (N_29998,N_29427,N_29361);
and U29999 (N_29999,N_29184,N_29050);
nor UO_0 (O_0,N_29673,N_29931);
nor UO_1 (O_1,N_29956,N_29926);
xor UO_2 (O_2,N_29593,N_29776);
and UO_3 (O_3,N_29906,N_29561);
and UO_4 (O_4,N_29840,N_29694);
nor UO_5 (O_5,N_29912,N_29891);
nand UO_6 (O_6,N_29811,N_29702);
nand UO_7 (O_7,N_29869,N_29873);
nand UO_8 (O_8,N_29944,N_29616);
nor UO_9 (O_9,N_29790,N_29831);
and UO_10 (O_10,N_29656,N_29661);
and UO_11 (O_11,N_29630,N_29989);
nor UO_12 (O_12,N_29670,N_29535);
or UO_13 (O_13,N_29826,N_29844);
and UO_14 (O_14,N_29932,N_29584);
or UO_15 (O_15,N_29868,N_29765);
xnor UO_16 (O_16,N_29686,N_29692);
or UO_17 (O_17,N_29958,N_29745);
and UO_18 (O_18,N_29585,N_29981);
and UO_19 (O_19,N_29708,N_29730);
and UO_20 (O_20,N_29591,N_29624);
nand UO_21 (O_21,N_29978,N_29977);
xnor UO_22 (O_22,N_29506,N_29774);
xor UO_23 (O_23,N_29987,N_29798);
nor UO_24 (O_24,N_29700,N_29613);
and UO_25 (O_25,N_29773,N_29666);
nor UO_26 (O_26,N_29922,N_29777);
xnor UO_27 (O_27,N_29703,N_29679);
nand UO_28 (O_28,N_29847,N_29523);
or UO_29 (O_29,N_29598,N_29684);
xor UO_30 (O_30,N_29541,N_29890);
and UO_31 (O_31,N_29893,N_29812);
xnor UO_32 (O_32,N_29783,N_29542);
xnor UO_33 (O_33,N_29964,N_29683);
xnor UO_34 (O_34,N_29736,N_29509);
xnor UO_35 (O_35,N_29642,N_29696);
or UO_36 (O_36,N_29522,N_29784);
or UO_37 (O_37,N_29508,N_29728);
xnor UO_38 (O_38,N_29809,N_29941);
xnor UO_39 (O_39,N_29665,N_29725);
nor UO_40 (O_40,N_29967,N_29654);
and UO_41 (O_41,N_29646,N_29636);
nor UO_42 (O_42,N_29907,N_29594);
and UO_43 (O_43,N_29763,N_29918);
and UO_44 (O_44,N_29878,N_29799);
xor UO_45 (O_45,N_29780,N_29995);
or UO_46 (O_46,N_29603,N_29856);
nand UO_47 (O_47,N_29933,N_29620);
nand UO_48 (O_48,N_29752,N_29996);
nor UO_49 (O_49,N_29807,N_29667);
xnor UO_50 (O_50,N_29657,N_29836);
and UO_51 (O_51,N_29822,N_29959);
nand UO_52 (O_52,N_29921,N_29568);
nand UO_53 (O_53,N_29729,N_29530);
or UO_54 (O_54,N_29991,N_29500);
or UO_55 (O_55,N_29533,N_29724);
nor UO_56 (O_56,N_29575,N_29827);
or UO_57 (O_57,N_29808,N_29501);
nand UO_58 (O_58,N_29574,N_29910);
nor UO_59 (O_59,N_29688,N_29737);
xnor UO_60 (O_60,N_29985,N_29528);
nand UO_61 (O_61,N_29539,N_29767);
or UO_62 (O_62,N_29817,N_29655);
and UO_63 (O_63,N_29502,N_29587);
xor UO_64 (O_64,N_29659,N_29547);
and UO_65 (O_65,N_29888,N_29992);
xnor UO_66 (O_66,N_29953,N_29791);
or UO_67 (O_67,N_29653,N_29747);
and UO_68 (O_68,N_29572,N_29560);
xor UO_69 (O_69,N_29599,N_29607);
nor UO_70 (O_70,N_29813,N_29693);
nand UO_71 (O_71,N_29548,N_29706);
nor UO_72 (O_72,N_29704,N_29723);
nor UO_73 (O_73,N_29875,N_29916);
or UO_74 (O_74,N_29942,N_29870);
or UO_75 (O_75,N_29556,N_29677);
nand UO_76 (O_76,N_29512,N_29757);
and UO_77 (O_77,N_29830,N_29590);
nand UO_78 (O_78,N_29586,N_29862);
and UO_79 (O_79,N_29573,N_29538);
xor UO_80 (O_80,N_29604,N_29866);
nand UO_81 (O_81,N_29674,N_29592);
xnor UO_82 (O_82,N_29897,N_29764);
xnor UO_83 (O_83,N_29838,N_29520);
or UO_84 (O_84,N_29966,N_29562);
and UO_85 (O_85,N_29879,N_29761);
or UO_86 (O_86,N_29505,N_29705);
nor UO_87 (O_87,N_29672,N_29682);
xnor UO_88 (O_88,N_29563,N_29731);
xor UO_89 (O_89,N_29880,N_29720);
nor UO_90 (O_90,N_29732,N_29871);
xor UO_91 (O_91,N_29643,N_29526);
nor UO_92 (O_92,N_29895,N_29837);
nand UO_93 (O_93,N_29972,N_29975);
nor UO_94 (O_94,N_29680,N_29537);
and UO_95 (O_95,N_29639,N_29908);
xor UO_96 (O_96,N_29796,N_29717);
or UO_97 (O_97,N_29637,N_29804);
nand UO_98 (O_98,N_29718,N_29621);
and UO_99 (O_99,N_29510,N_29716);
nand UO_100 (O_100,N_29531,N_29885);
and UO_101 (O_101,N_29845,N_29557);
xnor UO_102 (O_102,N_29821,N_29928);
nand UO_103 (O_103,N_29632,N_29652);
nand UO_104 (O_104,N_29943,N_29853);
and UO_105 (O_105,N_29711,N_29819);
or UO_106 (O_106,N_29823,N_29962);
and UO_107 (O_107,N_29927,N_29748);
and UO_108 (O_108,N_29519,N_29618);
xor UO_109 (O_109,N_29750,N_29608);
nor UO_110 (O_110,N_29581,N_29877);
xor UO_111 (O_111,N_29828,N_29899);
or UO_112 (O_112,N_29920,N_29852);
xnor UO_113 (O_113,N_29833,N_29957);
nand UO_114 (O_114,N_29936,N_29638);
xnor UO_115 (O_115,N_29758,N_29676);
or UO_116 (O_116,N_29825,N_29759);
nor UO_117 (O_117,N_29923,N_29628);
nand UO_118 (O_118,N_29946,N_29954);
or UO_119 (O_119,N_29970,N_29884);
nand UO_120 (O_120,N_29818,N_29785);
xnor UO_121 (O_121,N_29876,N_29851);
nor UO_122 (O_122,N_29629,N_29649);
nand UO_123 (O_123,N_29779,N_29947);
nor UO_124 (O_124,N_29612,N_29881);
nor UO_125 (O_125,N_29754,N_29669);
nor UO_126 (O_126,N_29648,N_29769);
or UO_127 (O_127,N_29787,N_29513);
and UO_128 (O_128,N_29645,N_29606);
nor UO_129 (O_129,N_29915,N_29631);
nand UO_130 (O_130,N_29960,N_29850);
and UO_131 (O_131,N_29635,N_29545);
nand UO_132 (O_132,N_29940,N_29609);
nand UO_133 (O_133,N_29503,N_29719);
and UO_134 (O_134,N_29514,N_29846);
and UO_135 (O_135,N_29794,N_29605);
nand UO_136 (O_136,N_29647,N_29625);
and UO_137 (O_137,N_29734,N_29998);
xor UO_138 (O_138,N_29892,N_29671);
nand UO_139 (O_139,N_29615,N_29715);
and UO_140 (O_140,N_29651,N_29595);
nand UO_141 (O_141,N_29986,N_29546);
or UO_142 (O_142,N_29663,N_29552);
or UO_143 (O_143,N_29622,N_29740);
xnor UO_144 (O_144,N_29951,N_29980);
nand UO_145 (O_145,N_29567,N_29633);
and UO_146 (O_146,N_29577,N_29861);
xor UO_147 (O_147,N_29801,N_29660);
and UO_148 (O_148,N_29532,N_29760);
nor UO_149 (O_149,N_29948,N_29739);
and UO_150 (O_150,N_29699,N_29945);
nand UO_151 (O_151,N_29619,N_29746);
nor UO_152 (O_152,N_29849,N_29865);
nand UO_153 (O_153,N_29925,N_29623);
nand UO_154 (O_154,N_29969,N_29990);
and UO_155 (O_155,N_29889,N_29938);
xnor UO_156 (O_156,N_29858,N_29722);
or UO_157 (O_157,N_29534,N_29733);
nor UO_158 (O_158,N_29540,N_29976);
or UO_159 (O_159,N_29580,N_29668);
xnor UO_160 (O_160,N_29793,N_29903);
and UO_161 (O_161,N_29707,N_29601);
nor UO_162 (O_162,N_29697,N_29775);
xor UO_163 (O_163,N_29582,N_29588);
nor UO_164 (O_164,N_29681,N_29919);
or UO_165 (O_165,N_29579,N_29781);
or UO_166 (O_166,N_29968,N_29507);
nand UO_167 (O_167,N_29641,N_29887);
nor UO_168 (O_168,N_29596,N_29685);
xnor UO_169 (O_169,N_29924,N_29566);
or UO_170 (O_170,N_29600,N_29786);
and UO_171 (O_171,N_29744,N_29952);
or UO_172 (O_172,N_29886,N_29762);
xor UO_173 (O_173,N_29771,N_29741);
nor UO_174 (O_174,N_29905,N_29900);
and UO_175 (O_175,N_29614,N_29626);
nor UO_176 (O_176,N_29743,N_29738);
nor UO_177 (O_177,N_29714,N_29511);
xnor UO_178 (O_178,N_29902,N_29742);
and UO_179 (O_179,N_29555,N_29883);
and UO_180 (O_180,N_29904,N_29549);
nand UO_181 (O_181,N_29982,N_29617);
xor UO_182 (O_182,N_29820,N_29553);
nand UO_183 (O_183,N_29835,N_29955);
nand UO_184 (O_184,N_29517,N_29857);
nand UO_185 (O_185,N_29901,N_29569);
xor UO_186 (O_186,N_29788,N_29735);
nand UO_187 (O_187,N_29710,N_29806);
and UO_188 (O_188,N_29937,N_29814);
nor UO_189 (O_189,N_29690,N_29695);
xnor UO_190 (O_190,N_29749,N_29999);
nor UO_191 (O_191,N_29611,N_29518);
or UO_192 (O_192,N_29678,N_29650);
nor UO_193 (O_193,N_29515,N_29894);
xnor UO_194 (O_194,N_29855,N_29721);
nor UO_195 (O_195,N_29644,N_29839);
nand UO_196 (O_196,N_29691,N_29755);
nand UO_197 (O_197,N_29554,N_29997);
or UO_198 (O_198,N_29766,N_29634);
nand UO_199 (O_199,N_29898,N_29701);
xor UO_200 (O_200,N_29864,N_29524);
xor UO_201 (O_201,N_29832,N_29854);
nor UO_202 (O_202,N_29860,N_29558);
or UO_203 (O_203,N_29504,N_29583);
nor UO_204 (O_204,N_29689,N_29536);
or UO_205 (O_205,N_29842,N_29917);
nand UO_206 (O_206,N_29727,N_29815);
nor UO_207 (O_207,N_29726,N_29973);
nand UO_208 (O_208,N_29963,N_29930);
and UO_209 (O_209,N_29802,N_29929);
or UO_210 (O_210,N_29803,N_29516);
nor UO_211 (O_211,N_29965,N_29602);
nor UO_212 (O_212,N_29529,N_29709);
nand UO_213 (O_213,N_29994,N_29627);
nand UO_214 (O_214,N_29589,N_29565);
nand UO_215 (O_215,N_29770,N_29834);
nor UO_216 (O_216,N_29824,N_29939);
nand UO_217 (O_217,N_29753,N_29578);
or UO_218 (O_218,N_29800,N_29527);
nand UO_219 (O_219,N_29874,N_29640);
and UO_220 (O_220,N_29843,N_29979);
xor UO_221 (O_221,N_29848,N_29950);
xor UO_222 (O_222,N_29984,N_29521);
nor UO_223 (O_223,N_29792,N_29551);
xor UO_224 (O_224,N_29772,N_29756);
xor UO_225 (O_225,N_29934,N_29789);
xnor UO_226 (O_226,N_29914,N_29971);
or UO_227 (O_227,N_29571,N_29778);
or UO_228 (O_228,N_29658,N_29882);
or UO_229 (O_229,N_29859,N_29687);
nand UO_230 (O_230,N_29795,N_29543);
xnor UO_231 (O_231,N_29768,N_29961);
nor UO_232 (O_232,N_29713,N_29782);
xor UO_233 (O_233,N_29576,N_29610);
or UO_234 (O_234,N_29867,N_29829);
or UO_235 (O_235,N_29974,N_29664);
or UO_236 (O_236,N_29751,N_29896);
xor UO_237 (O_237,N_29841,N_29550);
xnor UO_238 (O_238,N_29662,N_29810);
nor UO_239 (O_239,N_29570,N_29913);
xor UO_240 (O_240,N_29816,N_29564);
nor UO_241 (O_241,N_29993,N_29698);
or UO_242 (O_242,N_29805,N_29988);
nand UO_243 (O_243,N_29949,N_29525);
xor UO_244 (O_244,N_29872,N_29863);
nand UO_245 (O_245,N_29909,N_29911);
nand UO_246 (O_246,N_29544,N_29712);
nor UO_247 (O_247,N_29983,N_29597);
or UO_248 (O_248,N_29675,N_29935);
or UO_249 (O_249,N_29559,N_29797);
or UO_250 (O_250,N_29740,N_29863);
or UO_251 (O_251,N_29668,N_29890);
or UO_252 (O_252,N_29656,N_29783);
and UO_253 (O_253,N_29967,N_29954);
nand UO_254 (O_254,N_29716,N_29529);
nand UO_255 (O_255,N_29578,N_29631);
and UO_256 (O_256,N_29954,N_29611);
nor UO_257 (O_257,N_29640,N_29669);
xor UO_258 (O_258,N_29626,N_29565);
nand UO_259 (O_259,N_29599,N_29888);
nand UO_260 (O_260,N_29836,N_29523);
and UO_261 (O_261,N_29931,N_29883);
nor UO_262 (O_262,N_29698,N_29983);
and UO_263 (O_263,N_29861,N_29995);
or UO_264 (O_264,N_29674,N_29596);
or UO_265 (O_265,N_29804,N_29998);
or UO_266 (O_266,N_29870,N_29962);
nand UO_267 (O_267,N_29501,N_29747);
nor UO_268 (O_268,N_29747,N_29647);
xor UO_269 (O_269,N_29859,N_29968);
xnor UO_270 (O_270,N_29999,N_29815);
or UO_271 (O_271,N_29932,N_29806);
or UO_272 (O_272,N_29652,N_29902);
xor UO_273 (O_273,N_29731,N_29508);
or UO_274 (O_274,N_29544,N_29911);
nand UO_275 (O_275,N_29796,N_29967);
nor UO_276 (O_276,N_29937,N_29513);
and UO_277 (O_277,N_29983,N_29911);
and UO_278 (O_278,N_29516,N_29826);
xor UO_279 (O_279,N_29535,N_29521);
and UO_280 (O_280,N_29937,N_29939);
or UO_281 (O_281,N_29997,N_29788);
and UO_282 (O_282,N_29514,N_29877);
and UO_283 (O_283,N_29838,N_29781);
or UO_284 (O_284,N_29893,N_29629);
and UO_285 (O_285,N_29703,N_29544);
nor UO_286 (O_286,N_29919,N_29962);
xor UO_287 (O_287,N_29570,N_29561);
xor UO_288 (O_288,N_29997,N_29510);
nor UO_289 (O_289,N_29763,N_29564);
xor UO_290 (O_290,N_29629,N_29806);
and UO_291 (O_291,N_29516,N_29943);
or UO_292 (O_292,N_29619,N_29689);
and UO_293 (O_293,N_29862,N_29915);
or UO_294 (O_294,N_29789,N_29741);
or UO_295 (O_295,N_29702,N_29758);
nand UO_296 (O_296,N_29967,N_29850);
nor UO_297 (O_297,N_29509,N_29504);
xor UO_298 (O_298,N_29556,N_29951);
nand UO_299 (O_299,N_29884,N_29691);
nor UO_300 (O_300,N_29708,N_29881);
nor UO_301 (O_301,N_29700,N_29562);
xnor UO_302 (O_302,N_29872,N_29674);
and UO_303 (O_303,N_29522,N_29821);
and UO_304 (O_304,N_29986,N_29985);
and UO_305 (O_305,N_29953,N_29979);
nand UO_306 (O_306,N_29948,N_29629);
and UO_307 (O_307,N_29746,N_29867);
or UO_308 (O_308,N_29870,N_29856);
or UO_309 (O_309,N_29764,N_29844);
nand UO_310 (O_310,N_29623,N_29653);
nand UO_311 (O_311,N_29750,N_29956);
and UO_312 (O_312,N_29765,N_29959);
nand UO_313 (O_313,N_29734,N_29777);
nand UO_314 (O_314,N_29936,N_29845);
or UO_315 (O_315,N_29520,N_29924);
nor UO_316 (O_316,N_29766,N_29904);
or UO_317 (O_317,N_29514,N_29699);
or UO_318 (O_318,N_29828,N_29787);
nor UO_319 (O_319,N_29543,N_29662);
and UO_320 (O_320,N_29548,N_29573);
and UO_321 (O_321,N_29772,N_29712);
nand UO_322 (O_322,N_29520,N_29829);
nor UO_323 (O_323,N_29644,N_29922);
and UO_324 (O_324,N_29846,N_29718);
and UO_325 (O_325,N_29844,N_29676);
and UO_326 (O_326,N_29606,N_29888);
and UO_327 (O_327,N_29576,N_29523);
nor UO_328 (O_328,N_29979,N_29868);
xnor UO_329 (O_329,N_29612,N_29676);
and UO_330 (O_330,N_29952,N_29692);
and UO_331 (O_331,N_29796,N_29753);
or UO_332 (O_332,N_29724,N_29502);
xor UO_333 (O_333,N_29658,N_29690);
and UO_334 (O_334,N_29837,N_29812);
xor UO_335 (O_335,N_29966,N_29873);
and UO_336 (O_336,N_29964,N_29707);
and UO_337 (O_337,N_29855,N_29605);
nand UO_338 (O_338,N_29988,N_29580);
or UO_339 (O_339,N_29835,N_29524);
xnor UO_340 (O_340,N_29653,N_29584);
and UO_341 (O_341,N_29926,N_29616);
and UO_342 (O_342,N_29766,N_29706);
nor UO_343 (O_343,N_29852,N_29529);
or UO_344 (O_344,N_29805,N_29964);
and UO_345 (O_345,N_29791,N_29741);
or UO_346 (O_346,N_29934,N_29998);
and UO_347 (O_347,N_29787,N_29532);
nor UO_348 (O_348,N_29822,N_29607);
or UO_349 (O_349,N_29911,N_29826);
nor UO_350 (O_350,N_29927,N_29759);
nand UO_351 (O_351,N_29812,N_29621);
nor UO_352 (O_352,N_29711,N_29677);
nor UO_353 (O_353,N_29562,N_29911);
nand UO_354 (O_354,N_29706,N_29750);
and UO_355 (O_355,N_29838,N_29721);
or UO_356 (O_356,N_29839,N_29853);
nand UO_357 (O_357,N_29966,N_29835);
xor UO_358 (O_358,N_29525,N_29663);
xnor UO_359 (O_359,N_29845,N_29522);
and UO_360 (O_360,N_29849,N_29826);
and UO_361 (O_361,N_29631,N_29548);
and UO_362 (O_362,N_29792,N_29962);
and UO_363 (O_363,N_29655,N_29644);
xor UO_364 (O_364,N_29871,N_29531);
xnor UO_365 (O_365,N_29987,N_29956);
xnor UO_366 (O_366,N_29579,N_29547);
and UO_367 (O_367,N_29651,N_29885);
nand UO_368 (O_368,N_29557,N_29930);
or UO_369 (O_369,N_29970,N_29718);
nand UO_370 (O_370,N_29835,N_29957);
xor UO_371 (O_371,N_29645,N_29524);
xor UO_372 (O_372,N_29649,N_29843);
xor UO_373 (O_373,N_29623,N_29517);
or UO_374 (O_374,N_29808,N_29755);
or UO_375 (O_375,N_29921,N_29606);
and UO_376 (O_376,N_29946,N_29963);
and UO_377 (O_377,N_29933,N_29858);
xor UO_378 (O_378,N_29921,N_29961);
or UO_379 (O_379,N_29724,N_29623);
nor UO_380 (O_380,N_29793,N_29886);
nor UO_381 (O_381,N_29655,N_29764);
xor UO_382 (O_382,N_29855,N_29816);
xnor UO_383 (O_383,N_29893,N_29590);
xnor UO_384 (O_384,N_29579,N_29679);
nor UO_385 (O_385,N_29529,N_29977);
nand UO_386 (O_386,N_29760,N_29757);
nand UO_387 (O_387,N_29800,N_29812);
or UO_388 (O_388,N_29548,N_29595);
and UO_389 (O_389,N_29724,N_29678);
nor UO_390 (O_390,N_29910,N_29552);
or UO_391 (O_391,N_29875,N_29635);
nor UO_392 (O_392,N_29664,N_29533);
nand UO_393 (O_393,N_29678,N_29781);
nand UO_394 (O_394,N_29551,N_29970);
or UO_395 (O_395,N_29612,N_29568);
nor UO_396 (O_396,N_29980,N_29867);
or UO_397 (O_397,N_29810,N_29511);
nor UO_398 (O_398,N_29869,N_29563);
or UO_399 (O_399,N_29711,N_29507);
or UO_400 (O_400,N_29910,N_29505);
nor UO_401 (O_401,N_29897,N_29617);
xnor UO_402 (O_402,N_29959,N_29698);
nand UO_403 (O_403,N_29739,N_29703);
xnor UO_404 (O_404,N_29565,N_29703);
and UO_405 (O_405,N_29509,N_29580);
and UO_406 (O_406,N_29555,N_29737);
nor UO_407 (O_407,N_29873,N_29759);
xnor UO_408 (O_408,N_29614,N_29887);
or UO_409 (O_409,N_29988,N_29841);
nand UO_410 (O_410,N_29819,N_29859);
xnor UO_411 (O_411,N_29790,N_29937);
or UO_412 (O_412,N_29712,N_29956);
and UO_413 (O_413,N_29915,N_29870);
or UO_414 (O_414,N_29734,N_29794);
nand UO_415 (O_415,N_29522,N_29943);
nand UO_416 (O_416,N_29592,N_29854);
nor UO_417 (O_417,N_29870,N_29850);
and UO_418 (O_418,N_29578,N_29621);
xor UO_419 (O_419,N_29709,N_29933);
and UO_420 (O_420,N_29800,N_29760);
nand UO_421 (O_421,N_29815,N_29816);
nor UO_422 (O_422,N_29929,N_29747);
or UO_423 (O_423,N_29732,N_29780);
nor UO_424 (O_424,N_29787,N_29937);
and UO_425 (O_425,N_29769,N_29674);
nor UO_426 (O_426,N_29972,N_29639);
nor UO_427 (O_427,N_29970,N_29579);
xnor UO_428 (O_428,N_29803,N_29558);
and UO_429 (O_429,N_29709,N_29685);
or UO_430 (O_430,N_29698,N_29553);
nand UO_431 (O_431,N_29702,N_29848);
xor UO_432 (O_432,N_29595,N_29918);
xnor UO_433 (O_433,N_29516,N_29766);
nand UO_434 (O_434,N_29613,N_29739);
xor UO_435 (O_435,N_29904,N_29908);
or UO_436 (O_436,N_29724,N_29946);
nand UO_437 (O_437,N_29765,N_29553);
xnor UO_438 (O_438,N_29759,N_29675);
nand UO_439 (O_439,N_29661,N_29588);
or UO_440 (O_440,N_29551,N_29532);
or UO_441 (O_441,N_29991,N_29663);
nand UO_442 (O_442,N_29759,N_29620);
nor UO_443 (O_443,N_29617,N_29950);
nor UO_444 (O_444,N_29843,N_29815);
nor UO_445 (O_445,N_29500,N_29631);
or UO_446 (O_446,N_29702,N_29596);
or UO_447 (O_447,N_29954,N_29821);
nor UO_448 (O_448,N_29915,N_29566);
or UO_449 (O_449,N_29827,N_29970);
xnor UO_450 (O_450,N_29912,N_29905);
and UO_451 (O_451,N_29947,N_29634);
xnor UO_452 (O_452,N_29647,N_29538);
and UO_453 (O_453,N_29788,N_29619);
xnor UO_454 (O_454,N_29960,N_29533);
or UO_455 (O_455,N_29533,N_29919);
and UO_456 (O_456,N_29867,N_29920);
or UO_457 (O_457,N_29694,N_29689);
xnor UO_458 (O_458,N_29860,N_29537);
xnor UO_459 (O_459,N_29675,N_29565);
nor UO_460 (O_460,N_29844,N_29941);
xnor UO_461 (O_461,N_29748,N_29566);
nor UO_462 (O_462,N_29744,N_29529);
or UO_463 (O_463,N_29974,N_29791);
and UO_464 (O_464,N_29817,N_29740);
and UO_465 (O_465,N_29761,N_29914);
nor UO_466 (O_466,N_29646,N_29950);
xor UO_467 (O_467,N_29944,N_29676);
nand UO_468 (O_468,N_29638,N_29618);
and UO_469 (O_469,N_29510,N_29521);
or UO_470 (O_470,N_29842,N_29644);
and UO_471 (O_471,N_29923,N_29685);
or UO_472 (O_472,N_29868,N_29575);
nor UO_473 (O_473,N_29836,N_29978);
nor UO_474 (O_474,N_29965,N_29666);
xor UO_475 (O_475,N_29997,N_29854);
and UO_476 (O_476,N_29699,N_29984);
and UO_477 (O_477,N_29978,N_29872);
nor UO_478 (O_478,N_29982,N_29874);
and UO_479 (O_479,N_29501,N_29932);
xnor UO_480 (O_480,N_29744,N_29523);
or UO_481 (O_481,N_29907,N_29753);
nand UO_482 (O_482,N_29816,N_29635);
nor UO_483 (O_483,N_29867,N_29599);
and UO_484 (O_484,N_29880,N_29943);
and UO_485 (O_485,N_29635,N_29844);
xor UO_486 (O_486,N_29969,N_29515);
and UO_487 (O_487,N_29616,N_29580);
xor UO_488 (O_488,N_29741,N_29576);
or UO_489 (O_489,N_29728,N_29581);
xnor UO_490 (O_490,N_29856,N_29547);
and UO_491 (O_491,N_29597,N_29982);
nor UO_492 (O_492,N_29996,N_29977);
xnor UO_493 (O_493,N_29604,N_29733);
and UO_494 (O_494,N_29925,N_29742);
nor UO_495 (O_495,N_29528,N_29556);
nor UO_496 (O_496,N_29995,N_29840);
and UO_497 (O_497,N_29887,N_29752);
and UO_498 (O_498,N_29833,N_29715);
or UO_499 (O_499,N_29917,N_29665);
nand UO_500 (O_500,N_29747,N_29953);
or UO_501 (O_501,N_29923,N_29900);
xor UO_502 (O_502,N_29973,N_29944);
or UO_503 (O_503,N_29769,N_29659);
and UO_504 (O_504,N_29657,N_29504);
nand UO_505 (O_505,N_29617,N_29664);
and UO_506 (O_506,N_29576,N_29730);
or UO_507 (O_507,N_29624,N_29509);
and UO_508 (O_508,N_29785,N_29681);
nand UO_509 (O_509,N_29937,N_29505);
or UO_510 (O_510,N_29819,N_29700);
nor UO_511 (O_511,N_29714,N_29791);
nand UO_512 (O_512,N_29859,N_29996);
or UO_513 (O_513,N_29675,N_29512);
or UO_514 (O_514,N_29618,N_29930);
and UO_515 (O_515,N_29581,N_29797);
nand UO_516 (O_516,N_29899,N_29547);
xnor UO_517 (O_517,N_29655,N_29964);
nand UO_518 (O_518,N_29555,N_29690);
xnor UO_519 (O_519,N_29832,N_29953);
nand UO_520 (O_520,N_29878,N_29933);
and UO_521 (O_521,N_29872,N_29556);
xnor UO_522 (O_522,N_29708,N_29548);
nor UO_523 (O_523,N_29751,N_29685);
and UO_524 (O_524,N_29652,N_29702);
or UO_525 (O_525,N_29702,N_29565);
and UO_526 (O_526,N_29918,N_29847);
and UO_527 (O_527,N_29821,N_29662);
xnor UO_528 (O_528,N_29610,N_29730);
and UO_529 (O_529,N_29965,N_29516);
xor UO_530 (O_530,N_29665,N_29672);
or UO_531 (O_531,N_29799,N_29598);
xnor UO_532 (O_532,N_29968,N_29594);
nor UO_533 (O_533,N_29963,N_29671);
xnor UO_534 (O_534,N_29956,N_29556);
nor UO_535 (O_535,N_29565,N_29832);
nand UO_536 (O_536,N_29738,N_29684);
nor UO_537 (O_537,N_29824,N_29812);
or UO_538 (O_538,N_29843,N_29917);
nand UO_539 (O_539,N_29528,N_29754);
or UO_540 (O_540,N_29521,N_29590);
xor UO_541 (O_541,N_29619,N_29510);
or UO_542 (O_542,N_29683,N_29781);
nand UO_543 (O_543,N_29994,N_29634);
and UO_544 (O_544,N_29747,N_29585);
nand UO_545 (O_545,N_29718,N_29687);
and UO_546 (O_546,N_29604,N_29616);
or UO_547 (O_547,N_29614,N_29675);
xnor UO_548 (O_548,N_29510,N_29674);
nand UO_549 (O_549,N_29505,N_29889);
and UO_550 (O_550,N_29756,N_29650);
or UO_551 (O_551,N_29682,N_29608);
nand UO_552 (O_552,N_29814,N_29570);
and UO_553 (O_553,N_29879,N_29925);
and UO_554 (O_554,N_29935,N_29853);
nand UO_555 (O_555,N_29834,N_29871);
nor UO_556 (O_556,N_29675,N_29570);
nor UO_557 (O_557,N_29503,N_29963);
xnor UO_558 (O_558,N_29634,N_29622);
nand UO_559 (O_559,N_29626,N_29586);
nand UO_560 (O_560,N_29558,N_29500);
nand UO_561 (O_561,N_29592,N_29961);
nor UO_562 (O_562,N_29621,N_29540);
nor UO_563 (O_563,N_29719,N_29955);
nor UO_564 (O_564,N_29869,N_29971);
or UO_565 (O_565,N_29730,N_29619);
nor UO_566 (O_566,N_29976,N_29697);
or UO_567 (O_567,N_29581,N_29610);
nor UO_568 (O_568,N_29766,N_29612);
nor UO_569 (O_569,N_29765,N_29538);
nor UO_570 (O_570,N_29724,N_29668);
and UO_571 (O_571,N_29766,N_29898);
xnor UO_572 (O_572,N_29826,N_29949);
or UO_573 (O_573,N_29987,N_29669);
nand UO_574 (O_574,N_29713,N_29688);
nor UO_575 (O_575,N_29908,N_29538);
or UO_576 (O_576,N_29704,N_29930);
nand UO_577 (O_577,N_29814,N_29910);
nor UO_578 (O_578,N_29680,N_29504);
or UO_579 (O_579,N_29783,N_29658);
or UO_580 (O_580,N_29575,N_29714);
and UO_581 (O_581,N_29809,N_29945);
xor UO_582 (O_582,N_29952,N_29980);
and UO_583 (O_583,N_29722,N_29734);
nand UO_584 (O_584,N_29783,N_29723);
and UO_585 (O_585,N_29609,N_29991);
or UO_586 (O_586,N_29902,N_29610);
xnor UO_587 (O_587,N_29788,N_29862);
nor UO_588 (O_588,N_29601,N_29544);
nor UO_589 (O_589,N_29746,N_29999);
xnor UO_590 (O_590,N_29925,N_29978);
or UO_591 (O_591,N_29611,N_29570);
nand UO_592 (O_592,N_29672,N_29751);
nor UO_593 (O_593,N_29893,N_29603);
and UO_594 (O_594,N_29622,N_29707);
nand UO_595 (O_595,N_29635,N_29936);
xnor UO_596 (O_596,N_29840,N_29774);
or UO_597 (O_597,N_29722,N_29637);
or UO_598 (O_598,N_29690,N_29881);
nand UO_599 (O_599,N_29526,N_29842);
nand UO_600 (O_600,N_29924,N_29940);
xor UO_601 (O_601,N_29530,N_29656);
nand UO_602 (O_602,N_29640,N_29792);
nor UO_603 (O_603,N_29694,N_29607);
and UO_604 (O_604,N_29662,N_29548);
nand UO_605 (O_605,N_29982,N_29810);
and UO_606 (O_606,N_29835,N_29784);
xor UO_607 (O_607,N_29788,N_29949);
nor UO_608 (O_608,N_29736,N_29553);
nor UO_609 (O_609,N_29922,N_29716);
or UO_610 (O_610,N_29655,N_29839);
nor UO_611 (O_611,N_29771,N_29556);
xnor UO_612 (O_612,N_29986,N_29913);
nand UO_613 (O_613,N_29536,N_29679);
xnor UO_614 (O_614,N_29673,N_29642);
nand UO_615 (O_615,N_29987,N_29522);
xnor UO_616 (O_616,N_29587,N_29707);
or UO_617 (O_617,N_29665,N_29503);
and UO_618 (O_618,N_29614,N_29962);
nand UO_619 (O_619,N_29983,N_29523);
or UO_620 (O_620,N_29684,N_29674);
or UO_621 (O_621,N_29614,N_29863);
nand UO_622 (O_622,N_29613,N_29975);
xor UO_623 (O_623,N_29892,N_29502);
nor UO_624 (O_624,N_29882,N_29585);
xor UO_625 (O_625,N_29560,N_29818);
or UO_626 (O_626,N_29957,N_29885);
xnor UO_627 (O_627,N_29581,N_29722);
nand UO_628 (O_628,N_29562,N_29612);
or UO_629 (O_629,N_29512,N_29771);
xor UO_630 (O_630,N_29816,N_29622);
xnor UO_631 (O_631,N_29983,N_29559);
nand UO_632 (O_632,N_29949,N_29984);
xor UO_633 (O_633,N_29878,N_29912);
or UO_634 (O_634,N_29831,N_29549);
xor UO_635 (O_635,N_29510,N_29995);
nand UO_636 (O_636,N_29972,N_29902);
and UO_637 (O_637,N_29791,N_29724);
or UO_638 (O_638,N_29809,N_29537);
xor UO_639 (O_639,N_29768,N_29505);
nand UO_640 (O_640,N_29810,N_29545);
nor UO_641 (O_641,N_29998,N_29588);
and UO_642 (O_642,N_29745,N_29574);
and UO_643 (O_643,N_29936,N_29758);
nand UO_644 (O_644,N_29862,N_29623);
nand UO_645 (O_645,N_29676,N_29592);
nor UO_646 (O_646,N_29549,N_29926);
and UO_647 (O_647,N_29647,N_29600);
xnor UO_648 (O_648,N_29923,N_29939);
or UO_649 (O_649,N_29993,N_29870);
xor UO_650 (O_650,N_29513,N_29561);
nor UO_651 (O_651,N_29992,N_29586);
nor UO_652 (O_652,N_29712,N_29893);
and UO_653 (O_653,N_29639,N_29755);
nor UO_654 (O_654,N_29764,N_29889);
nand UO_655 (O_655,N_29741,N_29812);
nand UO_656 (O_656,N_29682,N_29670);
nand UO_657 (O_657,N_29707,N_29702);
and UO_658 (O_658,N_29876,N_29696);
and UO_659 (O_659,N_29577,N_29834);
xnor UO_660 (O_660,N_29838,N_29574);
and UO_661 (O_661,N_29622,N_29718);
nor UO_662 (O_662,N_29959,N_29916);
nor UO_663 (O_663,N_29578,N_29660);
or UO_664 (O_664,N_29899,N_29960);
nand UO_665 (O_665,N_29579,N_29737);
or UO_666 (O_666,N_29761,N_29644);
nand UO_667 (O_667,N_29515,N_29886);
and UO_668 (O_668,N_29804,N_29574);
nand UO_669 (O_669,N_29859,N_29959);
nand UO_670 (O_670,N_29889,N_29952);
or UO_671 (O_671,N_29600,N_29868);
or UO_672 (O_672,N_29633,N_29868);
nand UO_673 (O_673,N_29667,N_29703);
nand UO_674 (O_674,N_29660,N_29763);
nand UO_675 (O_675,N_29599,N_29822);
nand UO_676 (O_676,N_29522,N_29922);
nand UO_677 (O_677,N_29924,N_29706);
nand UO_678 (O_678,N_29821,N_29998);
and UO_679 (O_679,N_29993,N_29744);
or UO_680 (O_680,N_29761,N_29542);
nand UO_681 (O_681,N_29835,N_29811);
nor UO_682 (O_682,N_29875,N_29968);
or UO_683 (O_683,N_29999,N_29545);
nand UO_684 (O_684,N_29936,N_29909);
nor UO_685 (O_685,N_29842,N_29875);
or UO_686 (O_686,N_29773,N_29911);
and UO_687 (O_687,N_29715,N_29685);
nor UO_688 (O_688,N_29997,N_29682);
nand UO_689 (O_689,N_29833,N_29555);
nor UO_690 (O_690,N_29695,N_29775);
and UO_691 (O_691,N_29635,N_29701);
xnor UO_692 (O_692,N_29746,N_29717);
nor UO_693 (O_693,N_29621,N_29701);
or UO_694 (O_694,N_29732,N_29673);
nor UO_695 (O_695,N_29579,N_29639);
and UO_696 (O_696,N_29691,N_29701);
nor UO_697 (O_697,N_29602,N_29951);
or UO_698 (O_698,N_29688,N_29860);
xor UO_699 (O_699,N_29670,N_29525);
nor UO_700 (O_700,N_29758,N_29928);
nand UO_701 (O_701,N_29720,N_29777);
nand UO_702 (O_702,N_29641,N_29649);
xnor UO_703 (O_703,N_29880,N_29701);
nand UO_704 (O_704,N_29720,N_29900);
or UO_705 (O_705,N_29813,N_29848);
or UO_706 (O_706,N_29528,N_29623);
nand UO_707 (O_707,N_29912,N_29800);
and UO_708 (O_708,N_29861,N_29594);
and UO_709 (O_709,N_29711,N_29638);
or UO_710 (O_710,N_29526,N_29887);
xnor UO_711 (O_711,N_29659,N_29786);
nand UO_712 (O_712,N_29787,N_29939);
and UO_713 (O_713,N_29967,N_29523);
xnor UO_714 (O_714,N_29589,N_29720);
nand UO_715 (O_715,N_29560,N_29552);
nand UO_716 (O_716,N_29574,N_29847);
nand UO_717 (O_717,N_29530,N_29667);
xor UO_718 (O_718,N_29826,N_29647);
or UO_719 (O_719,N_29870,N_29859);
nand UO_720 (O_720,N_29523,N_29775);
xor UO_721 (O_721,N_29905,N_29759);
or UO_722 (O_722,N_29998,N_29776);
nor UO_723 (O_723,N_29745,N_29612);
and UO_724 (O_724,N_29673,N_29560);
nand UO_725 (O_725,N_29716,N_29986);
nor UO_726 (O_726,N_29580,N_29653);
xor UO_727 (O_727,N_29883,N_29597);
xnor UO_728 (O_728,N_29544,N_29729);
or UO_729 (O_729,N_29998,N_29897);
xor UO_730 (O_730,N_29985,N_29946);
and UO_731 (O_731,N_29809,N_29913);
xor UO_732 (O_732,N_29979,N_29671);
nor UO_733 (O_733,N_29690,N_29698);
xnor UO_734 (O_734,N_29889,N_29507);
nand UO_735 (O_735,N_29935,N_29564);
nand UO_736 (O_736,N_29868,N_29592);
and UO_737 (O_737,N_29848,N_29553);
nand UO_738 (O_738,N_29974,N_29889);
or UO_739 (O_739,N_29876,N_29608);
nand UO_740 (O_740,N_29937,N_29904);
xor UO_741 (O_741,N_29603,N_29679);
xor UO_742 (O_742,N_29888,N_29980);
xnor UO_743 (O_743,N_29984,N_29768);
nand UO_744 (O_744,N_29643,N_29552);
xor UO_745 (O_745,N_29552,N_29877);
xnor UO_746 (O_746,N_29827,N_29837);
and UO_747 (O_747,N_29848,N_29502);
nor UO_748 (O_748,N_29590,N_29674);
nor UO_749 (O_749,N_29735,N_29558);
xnor UO_750 (O_750,N_29878,N_29992);
and UO_751 (O_751,N_29640,N_29804);
nand UO_752 (O_752,N_29782,N_29697);
or UO_753 (O_753,N_29713,N_29514);
nand UO_754 (O_754,N_29653,N_29933);
nor UO_755 (O_755,N_29548,N_29670);
and UO_756 (O_756,N_29825,N_29528);
nand UO_757 (O_757,N_29865,N_29649);
xor UO_758 (O_758,N_29772,N_29816);
nand UO_759 (O_759,N_29685,N_29943);
nor UO_760 (O_760,N_29777,N_29963);
xor UO_761 (O_761,N_29659,N_29741);
or UO_762 (O_762,N_29921,N_29749);
xor UO_763 (O_763,N_29578,N_29976);
xor UO_764 (O_764,N_29753,N_29905);
nand UO_765 (O_765,N_29687,N_29780);
nor UO_766 (O_766,N_29911,N_29628);
and UO_767 (O_767,N_29526,N_29900);
or UO_768 (O_768,N_29727,N_29598);
or UO_769 (O_769,N_29839,N_29552);
xor UO_770 (O_770,N_29650,N_29530);
and UO_771 (O_771,N_29672,N_29725);
and UO_772 (O_772,N_29874,N_29604);
nor UO_773 (O_773,N_29921,N_29523);
xnor UO_774 (O_774,N_29618,N_29987);
nor UO_775 (O_775,N_29851,N_29900);
and UO_776 (O_776,N_29568,N_29720);
or UO_777 (O_777,N_29844,N_29724);
nor UO_778 (O_778,N_29762,N_29767);
and UO_779 (O_779,N_29973,N_29917);
nand UO_780 (O_780,N_29816,N_29594);
xor UO_781 (O_781,N_29698,N_29859);
or UO_782 (O_782,N_29721,N_29535);
nor UO_783 (O_783,N_29851,N_29505);
or UO_784 (O_784,N_29603,N_29614);
or UO_785 (O_785,N_29867,N_29753);
xor UO_786 (O_786,N_29804,N_29988);
or UO_787 (O_787,N_29657,N_29650);
or UO_788 (O_788,N_29989,N_29550);
and UO_789 (O_789,N_29653,N_29501);
and UO_790 (O_790,N_29873,N_29860);
nor UO_791 (O_791,N_29713,N_29519);
or UO_792 (O_792,N_29679,N_29987);
xor UO_793 (O_793,N_29962,N_29501);
nand UO_794 (O_794,N_29952,N_29735);
xor UO_795 (O_795,N_29686,N_29934);
nand UO_796 (O_796,N_29522,N_29980);
nor UO_797 (O_797,N_29665,N_29596);
nor UO_798 (O_798,N_29908,N_29892);
or UO_799 (O_799,N_29520,N_29734);
nor UO_800 (O_800,N_29773,N_29993);
nor UO_801 (O_801,N_29590,N_29974);
nor UO_802 (O_802,N_29576,N_29642);
and UO_803 (O_803,N_29793,N_29503);
or UO_804 (O_804,N_29589,N_29966);
xnor UO_805 (O_805,N_29790,N_29686);
or UO_806 (O_806,N_29579,N_29986);
nand UO_807 (O_807,N_29653,N_29648);
xnor UO_808 (O_808,N_29577,N_29990);
nor UO_809 (O_809,N_29973,N_29968);
and UO_810 (O_810,N_29602,N_29897);
nand UO_811 (O_811,N_29980,N_29606);
or UO_812 (O_812,N_29984,N_29978);
and UO_813 (O_813,N_29633,N_29902);
or UO_814 (O_814,N_29669,N_29681);
and UO_815 (O_815,N_29558,N_29788);
or UO_816 (O_816,N_29653,N_29981);
nand UO_817 (O_817,N_29898,N_29840);
nand UO_818 (O_818,N_29574,N_29935);
nand UO_819 (O_819,N_29511,N_29859);
nand UO_820 (O_820,N_29509,N_29579);
xnor UO_821 (O_821,N_29857,N_29597);
or UO_822 (O_822,N_29810,N_29894);
and UO_823 (O_823,N_29767,N_29847);
nand UO_824 (O_824,N_29959,N_29505);
or UO_825 (O_825,N_29839,N_29696);
xnor UO_826 (O_826,N_29697,N_29854);
and UO_827 (O_827,N_29776,N_29530);
nor UO_828 (O_828,N_29713,N_29900);
nand UO_829 (O_829,N_29938,N_29728);
nand UO_830 (O_830,N_29861,N_29765);
nor UO_831 (O_831,N_29932,N_29665);
nor UO_832 (O_832,N_29891,N_29852);
and UO_833 (O_833,N_29648,N_29955);
xnor UO_834 (O_834,N_29605,N_29669);
nand UO_835 (O_835,N_29984,N_29688);
and UO_836 (O_836,N_29667,N_29794);
nor UO_837 (O_837,N_29508,N_29522);
and UO_838 (O_838,N_29963,N_29697);
and UO_839 (O_839,N_29675,N_29901);
xor UO_840 (O_840,N_29944,N_29786);
xnor UO_841 (O_841,N_29536,N_29516);
nor UO_842 (O_842,N_29691,N_29771);
or UO_843 (O_843,N_29893,N_29760);
nor UO_844 (O_844,N_29981,N_29598);
xor UO_845 (O_845,N_29602,N_29770);
or UO_846 (O_846,N_29573,N_29746);
nor UO_847 (O_847,N_29623,N_29818);
nor UO_848 (O_848,N_29932,N_29672);
nor UO_849 (O_849,N_29722,N_29720);
nand UO_850 (O_850,N_29984,N_29587);
or UO_851 (O_851,N_29693,N_29810);
xnor UO_852 (O_852,N_29988,N_29554);
and UO_853 (O_853,N_29540,N_29904);
nand UO_854 (O_854,N_29649,N_29592);
xor UO_855 (O_855,N_29566,N_29577);
nand UO_856 (O_856,N_29935,N_29741);
or UO_857 (O_857,N_29609,N_29534);
or UO_858 (O_858,N_29998,N_29916);
or UO_859 (O_859,N_29551,N_29989);
and UO_860 (O_860,N_29909,N_29701);
and UO_861 (O_861,N_29757,N_29872);
or UO_862 (O_862,N_29734,N_29693);
and UO_863 (O_863,N_29708,N_29570);
xnor UO_864 (O_864,N_29718,N_29916);
xnor UO_865 (O_865,N_29708,N_29600);
or UO_866 (O_866,N_29548,N_29814);
nor UO_867 (O_867,N_29875,N_29977);
nor UO_868 (O_868,N_29583,N_29672);
nor UO_869 (O_869,N_29879,N_29972);
and UO_870 (O_870,N_29751,N_29535);
and UO_871 (O_871,N_29992,N_29604);
or UO_872 (O_872,N_29745,N_29627);
nor UO_873 (O_873,N_29558,N_29576);
nor UO_874 (O_874,N_29621,N_29755);
or UO_875 (O_875,N_29707,N_29986);
xnor UO_876 (O_876,N_29595,N_29733);
nor UO_877 (O_877,N_29551,N_29976);
or UO_878 (O_878,N_29745,N_29882);
or UO_879 (O_879,N_29804,N_29843);
nor UO_880 (O_880,N_29536,N_29851);
and UO_881 (O_881,N_29924,N_29672);
or UO_882 (O_882,N_29646,N_29722);
and UO_883 (O_883,N_29836,N_29988);
nand UO_884 (O_884,N_29682,N_29762);
and UO_885 (O_885,N_29754,N_29940);
xor UO_886 (O_886,N_29797,N_29724);
nand UO_887 (O_887,N_29994,N_29934);
and UO_888 (O_888,N_29684,N_29952);
nand UO_889 (O_889,N_29739,N_29783);
and UO_890 (O_890,N_29763,N_29530);
or UO_891 (O_891,N_29930,N_29701);
nand UO_892 (O_892,N_29796,N_29643);
nand UO_893 (O_893,N_29745,N_29625);
and UO_894 (O_894,N_29762,N_29774);
nor UO_895 (O_895,N_29774,N_29878);
nand UO_896 (O_896,N_29789,N_29896);
xnor UO_897 (O_897,N_29906,N_29683);
nor UO_898 (O_898,N_29908,N_29508);
nor UO_899 (O_899,N_29702,N_29550);
and UO_900 (O_900,N_29774,N_29633);
nor UO_901 (O_901,N_29772,N_29884);
nand UO_902 (O_902,N_29771,N_29864);
xnor UO_903 (O_903,N_29794,N_29762);
xor UO_904 (O_904,N_29726,N_29908);
nand UO_905 (O_905,N_29627,N_29879);
nand UO_906 (O_906,N_29647,N_29755);
or UO_907 (O_907,N_29762,N_29757);
or UO_908 (O_908,N_29874,N_29711);
or UO_909 (O_909,N_29948,N_29765);
nand UO_910 (O_910,N_29575,N_29551);
nand UO_911 (O_911,N_29623,N_29911);
or UO_912 (O_912,N_29835,N_29790);
and UO_913 (O_913,N_29507,N_29678);
nor UO_914 (O_914,N_29793,N_29993);
or UO_915 (O_915,N_29974,N_29655);
and UO_916 (O_916,N_29913,N_29516);
nand UO_917 (O_917,N_29562,N_29524);
xnor UO_918 (O_918,N_29610,N_29747);
nand UO_919 (O_919,N_29744,N_29745);
nor UO_920 (O_920,N_29838,N_29745);
nor UO_921 (O_921,N_29547,N_29728);
nor UO_922 (O_922,N_29764,N_29725);
or UO_923 (O_923,N_29978,N_29862);
and UO_924 (O_924,N_29765,N_29580);
and UO_925 (O_925,N_29596,N_29832);
xnor UO_926 (O_926,N_29939,N_29713);
xnor UO_927 (O_927,N_29969,N_29815);
xor UO_928 (O_928,N_29692,N_29926);
nand UO_929 (O_929,N_29967,N_29731);
nand UO_930 (O_930,N_29661,N_29998);
and UO_931 (O_931,N_29998,N_29996);
nor UO_932 (O_932,N_29710,N_29882);
or UO_933 (O_933,N_29946,N_29970);
and UO_934 (O_934,N_29901,N_29588);
xnor UO_935 (O_935,N_29542,N_29695);
nand UO_936 (O_936,N_29797,N_29535);
or UO_937 (O_937,N_29747,N_29570);
xnor UO_938 (O_938,N_29767,N_29698);
nor UO_939 (O_939,N_29568,N_29668);
nor UO_940 (O_940,N_29801,N_29634);
xnor UO_941 (O_941,N_29971,N_29545);
xnor UO_942 (O_942,N_29601,N_29941);
nand UO_943 (O_943,N_29697,N_29532);
xor UO_944 (O_944,N_29505,N_29765);
or UO_945 (O_945,N_29913,N_29785);
nor UO_946 (O_946,N_29908,N_29919);
or UO_947 (O_947,N_29550,N_29562);
xnor UO_948 (O_948,N_29672,N_29785);
xnor UO_949 (O_949,N_29613,N_29878);
nor UO_950 (O_950,N_29650,N_29993);
nand UO_951 (O_951,N_29784,N_29863);
nand UO_952 (O_952,N_29597,N_29732);
and UO_953 (O_953,N_29966,N_29516);
or UO_954 (O_954,N_29576,N_29926);
and UO_955 (O_955,N_29668,N_29728);
and UO_956 (O_956,N_29781,N_29816);
xor UO_957 (O_957,N_29761,N_29549);
xnor UO_958 (O_958,N_29843,N_29899);
nand UO_959 (O_959,N_29771,N_29884);
or UO_960 (O_960,N_29610,N_29848);
nor UO_961 (O_961,N_29579,N_29561);
nor UO_962 (O_962,N_29774,N_29720);
or UO_963 (O_963,N_29571,N_29975);
xor UO_964 (O_964,N_29850,N_29737);
and UO_965 (O_965,N_29662,N_29782);
nor UO_966 (O_966,N_29535,N_29628);
xnor UO_967 (O_967,N_29518,N_29976);
nand UO_968 (O_968,N_29510,N_29895);
xnor UO_969 (O_969,N_29807,N_29826);
and UO_970 (O_970,N_29602,N_29771);
nor UO_971 (O_971,N_29912,N_29718);
and UO_972 (O_972,N_29860,N_29517);
or UO_973 (O_973,N_29541,N_29915);
nor UO_974 (O_974,N_29711,N_29763);
xor UO_975 (O_975,N_29863,N_29992);
xnor UO_976 (O_976,N_29978,N_29954);
and UO_977 (O_977,N_29587,N_29956);
xor UO_978 (O_978,N_29528,N_29991);
nand UO_979 (O_979,N_29513,N_29934);
nor UO_980 (O_980,N_29940,N_29770);
nor UO_981 (O_981,N_29609,N_29682);
and UO_982 (O_982,N_29692,N_29765);
nand UO_983 (O_983,N_29992,N_29913);
xor UO_984 (O_984,N_29720,N_29768);
nor UO_985 (O_985,N_29897,N_29854);
or UO_986 (O_986,N_29953,N_29651);
and UO_987 (O_987,N_29580,N_29907);
and UO_988 (O_988,N_29749,N_29585);
nor UO_989 (O_989,N_29863,N_29916);
nor UO_990 (O_990,N_29656,N_29689);
and UO_991 (O_991,N_29508,N_29937);
nand UO_992 (O_992,N_29622,N_29879);
xor UO_993 (O_993,N_29626,N_29584);
and UO_994 (O_994,N_29713,N_29700);
xnor UO_995 (O_995,N_29596,N_29594);
xnor UO_996 (O_996,N_29540,N_29998);
or UO_997 (O_997,N_29997,N_29885);
or UO_998 (O_998,N_29591,N_29913);
nor UO_999 (O_999,N_29954,N_29927);
nor UO_1000 (O_1000,N_29646,N_29830);
xnor UO_1001 (O_1001,N_29529,N_29617);
nor UO_1002 (O_1002,N_29574,N_29984);
nor UO_1003 (O_1003,N_29841,N_29920);
nand UO_1004 (O_1004,N_29944,N_29789);
nand UO_1005 (O_1005,N_29946,N_29728);
and UO_1006 (O_1006,N_29593,N_29792);
nand UO_1007 (O_1007,N_29907,N_29820);
xor UO_1008 (O_1008,N_29997,N_29714);
or UO_1009 (O_1009,N_29845,N_29786);
nor UO_1010 (O_1010,N_29826,N_29673);
or UO_1011 (O_1011,N_29777,N_29820);
nand UO_1012 (O_1012,N_29558,N_29679);
nand UO_1013 (O_1013,N_29517,N_29739);
xor UO_1014 (O_1014,N_29959,N_29652);
nand UO_1015 (O_1015,N_29694,N_29805);
nor UO_1016 (O_1016,N_29684,N_29857);
or UO_1017 (O_1017,N_29670,N_29748);
xnor UO_1018 (O_1018,N_29901,N_29542);
nand UO_1019 (O_1019,N_29969,N_29565);
xnor UO_1020 (O_1020,N_29832,N_29900);
nand UO_1021 (O_1021,N_29796,N_29533);
nand UO_1022 (O_1022,N_29660,N_29866);
xnor UO_1023 (O_1023,N_29992,N_29720);
nor UO_1024 (O_1024,N_29676,N_29820);
xnor UO_1025 (O_1025,N_29562,N_29942);
nor UO_1026 (O_1026,N_29593,N_29904);
or UO_1027 (O_1027,N_29885,N_29589);
nor UO_1028 (O_1028,N_29931,N_29512);
or UO_1029 (O_1029,N_29595,N_29565);
nor UO_1030 (O_1030,N_29968,N_29526);
and UO_1031 (O_1031,N_29919,N_29644);
xnor UO_1032 (O_1032,N_29639,N_29546);
nand UO_1033 (O_1033,N_29916,N_29532);
nor UO_1034 (O_1034,N_29632,N_29980);
xor UO_1035 (O_1035,N_29877,N_29647);
xnor UO_1036 (O_1036,N_29560,N_29997);
or UO_1037 (O_1037,N_29822,N_29710);
nor UO_1038 (O_1038,N_29599,N_29561);
and UO_1039 (O_1039,N_29817,N_29518);
nor UO_1040 (O_1040,N_29760,N_29988);
nor UO_1041 (O_1041,N_29873,N_29547);
nor UO_1042 (O_1042,N_29621,N_29774);
or UO_1043 (O_1043,N_29775,N_29511);
xor UO_1044 (O_1044,N_29865,N_29664);
nor UO_1045 (O_1045,N_29620,N_29804);
xor UO_1046 (O_1046,N_29694,N_29826);
nor UO_1047 (O_1047,N_29968,N_29995);
nand UO_1048 (O_1048,N_29892,N_29515);
and UO_1049 (O_1049,N_29529,N_29670);
nand UO_1050 (O_1050,N_29926,N_29522);
nor UO_1051 (O_1051,N_29504,N_29949);
nand UO_1052 (O_1052,N_29836,N_29556);
nor UO_1053 (O_1053,N_29577,N_29930);
nand UO_1054 (O_1054,N_29548,N_29977);
nand UO_1055 (O_1055,N_29882,N_29805);
or UO_1056 (O_1056,N_29576,N_29783);
nor UO_1057 (O_1057,N_29658,N_29542);
nor UO_1058 (O_1058,N_29888,N_29824);
or UO_1059 (O_1059,N_29935,N_29642);
xnor UO_1060 (O_1060,N_29715,N_29594);
and UO_1061 (O_1061,N_29907,N_29817);
xnor UO_1062 (O_1062,N_29603,N_29573);
nor UO_1063 (O_1063,N_29554,N_29674);
or UO_1064 (O_1064,N_29946,N_29695);
xnor UO_1065 (O_1065,N_29509,N_29933);
xor UO_1066 (O_1066,N_29702,N_29722);
nand UO_1067 (O_1067,N_29953,N_29960);
xor UO_1068 (O_1068,N_29862,N_29537);
or UO_1069 (O_1069,N_29746,N_29935);
nand UO_1070 (O_1070,N_29928,N_29847);
or UO_1071 (O_1071,N_29955,N_29519);
nand UO_1072 (O_1072,N_29795,N_29969);
nor UO_1073 (O_1073,N_29522,N_29733);
nor UO_1074 (O_1074,N_29742,N_29926);
xnor UO_1075 (O_1075,N_29737,N_29769);
nand UO_1076 (O_1076,N_29967,N_29600);
xor UO_1077 (O_1077,N_29812,N_29635);
xnor UO_1078 (O_1078,N_29665,N_29633);
and UO_1079 (O_1079,N_29521,N_29553);
xnor UO_1080 (O_1080,N_29740,N_29799);
and UO_1081 (O_1081,N_29930,N_29552);
xnor UO_1082 (O_1082,N_29912,N_29615);
nand UO_1083 (O_1083,N_29852,N_29841);
xor UO_1084 (O_1084,N_29599,N_29698);
or UO_1085 (O_1085,N_29508,N_29801);
nor UO_1086 (O_1086,N_29858,N_29819);
nor UO_1087 (O_1087,N_29813,N_29833);
or UO_1088 (O_1088,N_29518,N_29592);
or UO_1089 (O_1089,N_29559,N_29532);
xor UO_1090 (O_1090,N_29717,N_29758);
or UO_1091 (O_1091,N_29640,N_29566);
xnor UO_1092 (O_1092,N_29565,N_29814);
or UO_1093 (O_1093,N_29898,N_29623);
nand UO_1094 (O_1094,N_29550,N_29649);
nor UO_1095 (O_1095,N_29979,N_29735);
nor UO_1096 (O_1096,N_29692,N_29792);
nor UO_1097 (O_1097,N_29738,N_29606);
and UO_1098 (O_1098,N_29589,N_29867);
nor UO_1099 (O_1099,N_29712,N_29853);
nor UO_1100 (O_1100,N_29672,N_29566);
xor UO_1101 (O_1101,N_29796,N_29744);
xor UO_1102 (O_1102,N_29810,N_29688);
nor UO_1103 (O_1103,N_29941,N_29511);
nand UO_1104 (O_1104,N_29623,N_29546);
xnor UO_1105 (O_1105,N_29734,N_29847);
and UO_1106 (O_1106,N_29738,N_29948);
nand UO_1107 (O_1107,N_29580,N_29852);
and UO_1108 (O_1108,N_29687,N_29951);
nor UO_1109 (O_1109,N_29729,N_29581);
xor UO_1110 (O_1110,N_29535,N_29629);
and UO_1111 (O_1111,N_29794,N_29976);
and UO_1112 (O_1112,N_29711,N_29984);
nand UO_1113 (O_1113,N_29875,N_29623);
nand UO_1114 (O_1114,N_29511,N_29894);
nor UO_1115 (O_1115,N_29559,N_29622);
nor UO_1116 (O_1116,N_29647,N_29716);
xor UO_1117 (O_1117,N_29950,N_29504);
nor UO_1118 (O_1118,N_29810,N_29561);
nand UO_1119 (O_1119,N_29521,N_29790);
nor UO_1120 (O_1120,N_29821,N_29952);
xor UO_1121 (O_1121,N_29580,N_29720);
xor UO_1122 (O_1122,N_29888,N_29525);
nand UO_1123 (O_1123,N_29777,N_29510);
nand UO_1124 (O_1124,N_29677,N_29510);
or UO_1125 (O_1125,N_29780,N_29629);
xnor UO_1126 (O_1126,N_29646,N_29649);
and UO_1127 (O_1127,N_29656,N_29937);
nor UO_1128 (O_1128,N_29802,N_29924);
nand UO_1129 (O_1129,N_29869,N_29799);
xnor UO_1130 (O_1130,N_29856,N_29582);
xnor UO_1131 (O_1131,N_29509,N_29796);
and UO_1132 (O_1132,N_29736,N_29688);
xnor UO_1133 (O_1133,N_29652,N_29610);
xor UO_1134 (O_1134,N_29838,N_29513);
nor UO_1135 (O_1135,N_29722,N_29730);
nand UO_1136 (O_1136,N_29851,N_29697);
nand UO_1137 (O_1137,N_29910,N_29604);
nor UO_1138 (O_1138,N_29972,N_29614);
nor UO_1139 (O_1139,N_29828,N_29959);
nor UO_1140 (O_1140,N_29687,N_29818);
or UO_1141 (O_1141,N_29806,N_29539);
and UO_1142 (O_1142,N_29771,N_29783);
nor UO_1143 (O_1143,N_29907,N_29700);
xor UO_1144 (O_1144,N_29566,N_29950);
nor UO_1145 (O_1145,N_29947,N_29589);
nor UO_1146 (O_1146,N_29795,N_29553);
nor UO_1147 (O_1147,N_29530,N_29634);
nor UO_1148 (O_1148,N_29949,N_29561);
nor UO_1149 (O_1149,N_29889,N_29965);
or UO_1150 (O_1150,N_29649,N_29914);
or UO_1151 (O_1151,N_29501,N_29587);
and UO_1152 (O_1152,N_29675,N_29859);
or UO_1153 (O_1153,N_29561,N_29836);
or UO_1154 (O_1154,N_29912,N_29924);
and UO_1155 (O_1155,N_29695,N_29534);
and UO_1156 (O_1156,N_29708,N_29610);
nor UO_1157 (O_1157,N_29704,N_29737);
xnor UO_1158 (O_1158,N_29895,N_29827);
nand UO_1159 (O_1159,N_29518,N_29500);
xor UO_1160 (O_1160,N_29751,N_29942);
xor UO_1161 (O_1161,N_29532,N_29558);
or UO_1162 (O_1162,N_29954,N_29647);
nand UO_1163 (O_1163,N_29996,N_29937);
nor UO_1164 (O_1164,N_29544,N_29850);
xor UO_1165 (O_1165,N_29734,N_29580);
xnor UO_1166 (O_1166,N_29545,N_29993);
and UO_1167 (O_1167,N_29682,N_29774);
and UO_1168 (O_1168,N_29922,N_29718);
or UO_1169 (O_1169,N_29901,N_29995);
xnor UO_1170 (O_1170,N_29772,N_29939);
and UO_1171 (O_1171,N_29839,N_29542);
nor UO_1172 (O_1172,N_29993,N_29742);
xnor UO_1173 (O_1173,N_29634,N_29524);
xor UO_1174 (O_1174,N_29513,N_29659);
xnor UO_1175 (O_1175,N_29623,N_29935);
nand UO_1176 (O_1176,N_29505,N_29539);
xnor UO_1177 (O_1177,N_29810,N_29905);
and UO_1178 (O_1178,N_29791,N_29731);
nor UO_1179 (O_1179,N_29529,N_29686);
and UO_1180 (O_1180,N_29674,N_29996);
nand UO_1181 (O_1181,N_29513,N_29747);
nand UO_1182 (O_1182,N_29518,N_29667);
or UO_1183 (O_1183,N_29736,N_29698);
and UO_1184 (O_1184,N_29925,N_29791);
or UO_1185 (O_1185,N_29578,N_29860);
xor UO_1186 (O_1186,N_29791,N_29993);
nand UO_1187 (O_1187,N_29910,N_29719);
nand UO_1188 (O_1188,N_29559,N_29773);
or UO_1189 (O_1189,N_29626,N_29807);
or UO_1190 (O_1190,N_29645,N_29756);
xor UO_1191 (O_1191,N_29506,N_29712);
nor UO_1192 (O_1192,N_29969,N_29573);
or UO_1193 (O_1193,N_29894,N_29862);
xor UO_1194 (O_1194,N_29831,N_29677);
and UO_1195 (O_1195,N_29808,N_29591);
nand UO_1196 (O_1196,N_29914,N_29531);
xnor UO_1197 (O_1197,N_29541,N_29503);
xnor UO_1198 (O_1198,N_29852,N_29809);
xnor UO_1199 (O_1199,N_29654,N_29525);
xor UO_1200 (O_1200,N_29774,N_29988);
nor UO_1201 (O_1201,N_29848,N_29544);
and UO_1202 (O_1202,N_29989,N_29942);
and UO_1203 (O_1203,N_29545,N_29629);
xor UO_1204 (O_1204,N_29616,N_29936);
or UO_1205 (O_1205,N_29560,N_29609);
xnor UO_1206 (O_1206,N_29614,N_29697);
xnor UO_1207 (O_1207,N_29926,N_29646);
and UO_1208 (O_1208,N_29771,N_29998);
and UO_1209 (O_1209,N_29593,N_29832);
nor UO_1210 (O_1210,N_29824,N_29878);
or UO_1211 (O_1211,N_29517,N_29717);
or UO_1212 (O_1212,N_29842,N_29728);
nor UO_1213 (O_1213,N_29950,N_29682);
xnor UO_1214 (O_1214,N_29500,N_29729);
nor UO_1215 (O_1215,N_29507,N_29948);
nor UO_1216 (O_1216,N_29610,N_29855);
or UO_1217 (O_1217,N_29584,N_29814);
nand UO_1218 (O_1218,N_29934,N_29565);
and UO_1219 (O_1219,N_29806,N_29647);
and UO_1220 (O_1220,N_29846,N_29707);
nand UO_1221 (O_1221,N_29797,N_29553);
xor UO_1222 (O_1222,N_29525,N_29872);
or UO_1223 (O_1223,N_29868,N_29598);
nand UO_1224 (O_1224,N_29816,N_29844);
xor UO_1225 (O_1225,N_29636,N_29928);
or UO_1226 (O_1226,N_29772,N_29659);
and UO_1227 (O_1227,N_29725,N_29929);
or UO_1228 (O_1228,N_29931,N_29533);
or UO_1229 (O_1229,N_29770,N_29882);
and UO_1230 (O_1230,N_29794,N_29857);
or UO_1231 (O_1231,N_29777,N_29761);
or UO_1232 (O_1232,N_29802,N_29987);
nor UO_1233 (O_1233,N_29936,N_29517);
or UO_1234 (O_1234,N_29902,N_29840);
nand UO_1235 (O_1235,N_29924,N_29922);
xnor UO_1236 (O_1236,N_29848,N_29706);
xor UO_1237 (O_1237,N_29511,N_29914);
nor UO_1238 (O_1238,N_29670,N_29700);
and UO_1239 (O_1239,N_29909,N_29652);
nor UO_1240 (O_1240,N_29678,N_29816);
or UO_1241 (O_1241,N_29837,N_29600);
xnor UO_1242 (O_1242,N_29736,N_29865);
and UO_1243 (O_1243,N_29703,N_29955);
or UO_1244 (O_1244,N_29676,N_29633);
or UO_1245 (O_1245,N_29981,N_29640);
nand UO_1246 (O_1246,N_29632,N_29561);
nand UO_1247 (O_1247,N_29514,N_29598);
nand UO_1248 (O_1248,N_29803,N_29780);
nor UO_1249 (O_1249,N_29945,N_29824);
or UO_1250 (O_1250,N_29544,N_29682);
nor UO_1251 (O_1251,N_29671,N_29922);
and UO_1252 (O_1252,N_29880,N_29518);
or UO_1253 (O_1253,N_29532,N_29680);
and UO_1254 (O_1254,N_29587,N_29767);
nand UO_1255 (O_1255,N_29560,N_29749);
or UO_1256 (O_1256,N_29678,N_29696);
xor UO_1257 (O_1257,N_29884,N_29702);
xnor UO_1258 (O_1258,N_29755,N_29895);
or UO_1259 (O_1259,N_29543,N_29566);
or UO_1260 (O_1260,N_29691,N_29971);
nor UO_1261 (O_1261,N_29983,N_29881);
or UO_1262 (O_1262,N_29896,N_29861);
and UO_1263 (O_1263,N_29679,N_29721);
and UO_1264 (O_1264,N_29724,N_29554);
nor UO_1265 (O_1265,N_29921,N_29714);
nor UO_1266 (O_1266,N_29969,N_29553);
nor UO_1267 (O_1267,N_29501,N_29676);
or UO_1268 (O_1268,N_29583,N_29731);
or UO_1269 (O_1269,N_29691,N_29570);
nor UO_1270 (O_1270,N_29569,N_29644);
nand UO_1271 (O_1271,N_29926,N_29947);
nor UO_1272 (O_1272,N_29738,N_29769);
nand UO_1273 (O_1273,N_29573,N_29635);
xnor UO_1274 (O_1274,N_29541,N_29724);
and UO_1275 (O_1275,N_29970,N_29711);
or UO_1276 (O_1276,N_29509,N_29979);
and UO_1277 (O_1277,N_29634,N_29863);
xnor UO_1278 (O_1278,N_29657,N_29574);
nor UO_1279 (O_1279,N_29503,N_29604);
and UO_1280 (O_1280,N_29906,N_29927);
or UO_1281 (O_1281,N_29809,N_29951);
xnor UO_1282 (O_1282,N_29541,N_29676);
and UO_1283 (O_1283,N_29598,N_29890);
xor UO_1284 (O_1284,N_29703,N_29678);
and UO_1285 (O_1285,N_29611,N_29870);
nor UO_1286 (O_1286,N_29553,N_29617);
or UO_1287 (O_1287,N_29858,N_29501);
nor UO_1288 (O_1288,N_29664,N_29573);
nand UO_1289 (O_1289,N_29997,N_29782);
xor UO_1290 (O_1290,N_29717,N_29894);
nor UO_1291 (O_1291,N_29857,N_29964);
xor UO_1292 (O_1292,N_29926,N_29709);
nor UO_1293 (O_1293,N_29882,N_29568);
xor UO_1294 (O_1294,N_29822,N_29978);
nand UO_1295 (O_1295,N_29695,N_29610);
and UO_1296 (O_1296,N_29728,N_29932);
nand UO_1297 (O_1297,N_29538,N_29508);
nand UO_1298 (O_1298,N_29981,N_29873);
and UO_1299 (O_1299,N_29847,N_29570);
xor UO_1300 (O_1300,N_29981,N_29945);
and UO_1301 (O_1301,N_29742,N_29744);
nor UO_1302 (O_1302,N_29524,N_29782);
nor UO_1303 (O_1303,N_29671,N_29630);
and UO_1304 (O_1304,N_29886,N_29786);
or UO_1305 (O_1305,N_29849,N_29763);
nor UO_1306 (O_1306,N_29799,N_29667);
nand UO_1307 (O_1307,N_29736,N_29597);
nor UO_1308 (O_1308,N_29932,N_29725);
and UO_1309 (O_1309,N_29665,N_29610);
and UO_1310 (O_1310,N_29576,N_29597);
xnor UO_1311 (O_1311,N_29900,N_29764);
nor UO_1312 (O_1312,N_29570,N_29621);
nand UO_1313 (O_1313,N_29835,N_29721);
and UO_1314 (O_1314,N_29631,N_29886);
xor UO_1315 (O_1315,N_29745,N_29582);
xnor UO_1316 (O_1316,N_29876,N_29661);
nand UO_1317 (O_1317,N_29634,N_29714);
nor UO_1318 (O_1318,N_29751,N_29779);
nor UO_1319 (O_1319,N_29635,N_29990);
or UO_1320 (O_1320,N_29838,N_29608);
xor UO_1321 (O_1321,N_29752,N_29661);
and UO_1322 (O_1322,N_29565,N_29991);
xnor UO_1323 (O_1323,N_29695,N_29892);
and UO_1324 (O_1324,N_29569,N_29783);
and UO_1325 (O_1325,N_29833,N_29741);
and UO_1326 (O_1326,N_29765,N_29912);
and UO_1327 (O_1327,N_29506,N_29628);
nand UO_1328 (O_1328,N_29670,N_29672);
xor UO_1329 (O_1329,N_29944,N_29879);
and UO_1330 (O_1330,N_29923,N_29667);
nor UO_1331 (O_1331,N_29966,N_29556);
xnor UO_1332 (O_1332,N_29749,N_29927);
xor UO_1333 (O_1333,N_29665,N_29784);
nor UO_1334 (O_1334,N_29759,N_29629);
nor UO_1335 (O_1335,N_29860,N_29944);
xnor UO_1336 (O_1336,N_29872,N_29592);
and UO_1337 (O_1337,N_29531,N_29518);
or UO_1338 (O_1338,N_29877,N_29785);
and UO_1339 (O_1339,N_29546,N_29660);
or UO_1340 (O_1340,N_29733,N_29768);
nand UO_1341 (O_1341,N_29923,N_29650);
nor UO_1342 (O_1342,N_29545,N_29706);
and UO_1343 (O_1343,N_29585,N_29565);
nand UO_1344 (O_1344,N_29989,N_29647);
nand UO_1345 (O_1345,N_29741,N_29613);
xnor UO_1346 (O_1346,N_29999,N_29921);
and UO_1347 (O_1347,N_29690,N_29773);
nand UO_1348 (O_1348,N_29615,N_29944);
nor UO_1349 (O_1349,N_29892,N_29643);
xor UO_1350 (O_1350,N_29835,N_29878);
and UO_1351 (O_1351,N_29597,N_29672);
or UO_1352 (O_1352,N_29962,N_29659);
nand UO_1353 (O_1353,N_29827,N_29653);
or UO_1354 (O_1354,N_29987,N_29623);
and UO_1355 (O_1355,N_29953,N_29726);
nand UO_1356 (O_1356,N_29916,N_29761);
or UO_1357 (O_1357,N_29520,N_29986);
or UO_1358 (O_1358,N_29787,N_29507);
and UO_1359 (O_1359,N_29820,N_29520);
nor UO_1360 (O_1360,N_29937,N_29712);
xor UO_1361 (O_1361,N_29839,N_29671);
nor UO_1362 (O_1362,N_29576,N_29640);
nor UO_1363 (O_1363,N_29895,N_29519);
xor UO_1364 (O_1364,N_29825,N_29539);
nor UO_1365 (O_1365,N_29968,N_29518);
nand UO_1366 (O_1366,N_29505,N_29555);
nand UO_1367 (O_1367,N_29610,N_29646);
nand UO_1368 (O_1368,N_29547,N_29544);
nor UO_1369 (O_1369,N_29692,N_29501);
nor UO_1370 (O_1370,N_29957,N_29979);
nor UO_1371 (O_1371,N_29926,N_29772);
or UO_1372 (O_1372,N_29902,N_29988);
and UO_1373 (O_1373,N_29556,N_29518);
and UO_1374 (O_1374,N_29722,N_29728);
xnor UO_1375 (O_1375,N_29716,N_29972);
nor UO_1376 (O_1376,N_29807,N_29785);
or UO_1377 (O_1377,N_29854,N_29963);
nor UO_1378 (O_1378,N_29848,N_29622);
and UO_1379 (O_1379,N_29548,N_29709);
nor UO_1380 (O_1380,N_29512,N_29895);
and UO_1381 (O_1381,N_29541,N_29559);
nand UO_1382 (O_1382,N_29595,N_29702);
nand UO_1383 (O_1383,N_29980,N_29920);
xor UO_1384 (O_1384,N_29898,N_29926);
nand UO_1385 (O_1385,N_29965,N_29883);
and UO_1386 (O_1386,N_29696,N_29675);
and UO_1387 (O_1387,N_29895,N_29571);
xor UO_1388 (O_1388,N_29671,N_29843);
and UO_1389 (O_1389,N_29685,N_29883);
nor UO_1390 (O_1390,N_29860,N_29932);
nor UO_1391 (O_1391,N_29983,N_29538);
and UO_1392 (O_1392,N_29939,N_29999);
and UO_1393 (O_1393,N_29977,N_29793);
and UO_1394 (O_1394,N_29681,N_29735);
or UO_1395 (O_1395,N_29735,N_29699);
and UO_1396 (O_1396,N_29885,N_29916);
and UO_1397 (O_1397,N_29795,N_29997);
and UO_1398 (O_1398,N_29590,N_29563);
xor UO_1399 (O_1399,N_29785,N_29627);
or UO_1400 (O_1400,N_29839,N_29539);
and UO_1401 (O_1401,N_29552,N_29822);
nand UO_1402 (O_1402,N_29714,N_29874);
and UO_1403 (O_1403,N_29612,N_29843);
or UO_1404 (O_1404,N_29631,N_29528);
nor UO_1405 (O_1405,N_29857,N_29949);
nand UO_1406 (O_1406,N_29522,N_29640);
or UO_1407 (O_1407,N_29694,N_29519);
nor UO_1408 (O_1408,N_29614,N_29854);
or UO_1409 (O_1409,N_29619,N_29958);
xor UO_1410 (O_1410,N_29596,N_29794);
nand UO_1411 (O_1411,N_29618,N_29688);
and UO_1412 (O_1412,N_29841,N_29941);
nand UO_1413 (O_1413,N_29523,N_29903);
and UO_1414 (O_1414,N_29845,N_29886);
xor UO_1415 (O_1415,N_29541,N_29610);
nand UO_1416 (O_1416,N_29982,N_29708);
nor UO_1417 (O_1417,N_29677,N_29612);
nor UO_1418 (O_1418,N_29754,N_29728);
xor UO_1419 (O_1419,N_29724,N_29879);
and UO_1420 (O_1420,N_29902,N_29619);
or UO_1421 (O_1421,N_29630,N_29631);
nor UO_1422 (O_1422,N_29645,N_29634);
or UO_1423 (O_1423,N_29690,N_29631);
nand UO_1424 (O_1424,N_29976,N_29613);
and UO_1425 (O_1425,N_29731,N_29922);
and UO_1426 (O_1426,N_29629,N_29908);
xnor UO_1427 (O_1427,N_29598,N_29546);
nand UO_1428 (O_1428,N_29931,N_29545);
nand UO_1429 (O_1429,N_29945,N_29705);
nor UO_1430 (O_1430,N_29972,N_29938);
xnor UO_1431 (O_1431,N_29576,N_29702);
or UO_1432 (O_1432,N_29967,N_29777);
nor UO_1433 (O_1433,N_29869,N_29956);
nand UO_1434 (O_1434,N_29624,N_29781);
or UO_1435 (O_1435,N_29878,N_29579);
xor UO_1436 (O_1436,N_29556,N_29782);
xnor UO_1437 (O_1437,N_29867,N_29579);
nor UO_1438 (O_1438,N_29575,N_29530);
or UO_1439 (O_1439,N_29545,N_29561);
and UO_1440 (O_1440,N_29958,N_29774);
nor UO_1441 (O_1441,N_29715,N_29539);
nand UO_1442 (O_1442,N_29980,N_29504);
nand UO_1443 (O_1443,N_29743,N_29643);
nor UO_1444 (O_1444,N_29907,N_29707);
xnor UO_1445 (O_1445,N_29657,N_29828);
nor UO_1446 (O_1446,N_29741,N_29510);
or UO_1447 (O_1447,N_29751,N_29953);
xnor UO_1448 (O_1448,N_29908,N_29720);
nand UO_1449 (O_1449,N_29874,N_29570);
nor UO_1450 (O_1450,N_29807,N_29712);
and UO_1451 (O_1451,N_29791,N_29616);
nor UO_1452 (O_1452,N_29842,N_29505);
nand UO_1453 (O_1453,N_29687,N_29990);
and UO_1454 (O_1454,N_29827,N_29715);
nor UO_1455 (O_1455,N_29809,N_29807);
and UO_1456 (O_1456,N_29642,N_29928);
nor UO_1457 (O_1457,N_29623,N_29831);
nand UO_1458 (O_1458,N_29608,N_29625);
nor UO_1459 (O_1459,N_29775,N_29881);
nand UO_1460 (O_1460,N_29956,N_29751);
nor UO_1461 (O_1461,N_29835,N_29611);
xor UO_1462 (O_1462,N_29811,N_29981);
nand UO_1463 (O_1463,N_29795,N_29981);
nand UO_1464 (O_1464,N_29821,N_29634);
xnor UO_1465 (O_1465,N_29728,N_29589);
and UO_1466 (O_1466,N_29828,N_29855);
nand UO_1467 (O_1467,N_29809,N_29763);
nand UO_1468 (O_1468,N_29702,N_29876);
nand UO_1469 (O_1469,N_29782,N_29710);
and UO_1470 (O_1470,N_29539,N_29901);
or UO_1471 (O_1471,N_29668,N_29954);
nor UO_1472 (O_1472,N_29774,N_29679);
and UO_1473 (O_1473,N_29561,N_29845);
nor UO_1474 (O_1474,N_29539,N_29573);
nand UO_1475 (O_1475,N_29587,N_29912);
and UO_1476 (O_1476,N_29960,N_29546);
nand UO_1477 (O_1477,N_29565,N_29569);
and UO_1478 (O_1478,N_29975,N_29570);
xnor UO_1479 (O_1479,N_29653,N_29713);
or UO_1480 (O_1480,N_29784,N_29550);
nor UO_1481 (O_1481,N_29962,N_29888);
or UO_1482 (O_1482,N_29936,N_29634);
nand UO_1483 (O_1483,N_29562,N_29884);
and UO_1484 (O_1484,N_29885,N_29854);
and UO_1485 (O_1485,N_29684,N_29958);
or UO_1486 (O_1486,N_29944,N_29791);
or UO_1487 (O_1487,N_29566,N_29702);
nand UO_1488 (O_1488,N_29944,N_29501);
nor UO_1489 (O_1489,N_29535,N_29568);
nor UO_1490 (O_1490,N_29905,N_29795);
nor UO_1491 (O_1491,N_29834,N_29845);
and UO_1492 (O_1492,N_29697,N_29511);
nand UO_1493 (O_1493,N_29783,N_29869);
and UO_1494 (O_1494,N_29768,N_29806);
nor UO_1495 (O_1495,N_29750,N_29721);
and UO_1496 (O_1496,N_29641,N_29991);
or UO_1497 (O_1497,N_29564,N_29991);
xnor UO_1498 (O_1498,N_29793,N_29515);
or UO_1499 (O_1499,N_29700,N_29598);
xnor UO_1500 (O_1500,N_29876,N_29719);
xor UO_1501 (O_1501,N_29600,N_29841);
and UO_1502 (O_1502,N_29603,N_29875);
nor UO_1503 (O_1503,N_29600,N_29550);
xnor UO_1504 (O_1504,N_29657,N_29655);
xnor UO_1505 (O_1505,N_29873,N_29923);
and UO_1506 (O_1506,N_29954,N_29884);
or UO_1507 (O_1507,N_29590,N_29876);
and UO_1508 (O_1508,N_29588,N_29931);
or UO_1509 (O_1509,N_29731,N_29650);
xor UO_1510 (O_1510,N_29683,N_29576);
nand UO_1511 (O_1511,N_29733,N_29701);
xnor UO_1512 (O_1512,N_29723,N_29504);
xnor UO_1513 (O_1513,N_29892,N_29682);
and UO_1514 (O_1514,N_29937,N_29563);
nand UO_1515 (O_1515,N_29678,N_29628);
and UO_1516 (O_1516,N_29768,N_29793);
xor UO_1517 (O_1517,N_29785,N_29864);
xor UO_1518 (O_1518,N_29788,N_29983);
and UO_1519 (O_1519,N_29578,N_29535);
and UO_1520 (O_1520,N_29548,N_29717);
and UO_1521 (O_1521,N_29898,N_29712);
xor UO_1522 (O_1522,N_29511,N_29623);
and UO_1523 (O_1523,N_29519,N_29938);
and UO_1524 (O_1524,N_29600,N_29508);
nor UO_1525 (O_1525,N_29997,N_29511);
nand UO_1526 (O_1526,N_29934,N_29740);
nand UO_1527 (O_1527,N_29578,N_29732);
nor UO_1528 (O_1528,N_29918,N_29944);
nand UO_1529 (O_1529,N_29746,N_29807);
or UO_1530 (O_1530,N_29722,N_29724);
and UO_1531 (O_1531,N_29605,N_29814);
nand UO_1532 (O_1532,N_29949,N_29887);
nand UO_1533 (O_1533,N_29715,N_29705);
and UO_1534 (O_1534,N_29879,N_29826);
nand UO_1535 (O_1535,N_29663,N_29808);
and UO_1536 (O_1536,N_29627,N_29927);
nor UO_1537 (O_1537,N_29917,N_29723);
nand UO_1538 (O_1538,N_29872,N_29818);
and UO_1539 (O_1539,N_29672,N_29917);
nand UO_1540 (O_1540,N_29724,N_29899);
nor UO_1541 (O_1541,N_29621,N_29593);
xnor UO_1542 (O_1542,N_29663,N_29683);
nor UO_1543 (O_1543,N_29792,N_29540);
or UO_1544 (O_1544,N_29955,N_29539);
or UO_1545 (O_1545,N_29824,N_29740);
nor UO_1546 (O_1546,N_29871,N_29914);
and UO_1547 (O_1547,N_29656,N_29692);
xor UO_1548 (O_1548,N_29645,N_29794);
or UO_1549 (O_1549,N_29563,N_29901);
nor UO_1550 (O_1550,N_29703,N_29844);
or UO_1551 (O_1551,N_29736,N_29815);
nand UO_1552 (O_1552,N_29552,N_29708);
nand UO_1553 (O_1553,N_29907,N_29782);
nand UO_1554 (O_1554,N_29943,N_29646);
nand UO_1555 (O_1555,N_29768,N_29659);
xnor UO_1556 (O_1556,N_29814,N_29838);
nand UO_1557 (O_1557,N_29991,N_29883);
nor UO_1558 (O_1558,N_29728,N_29618);
xor UO_1559 (O_1559,N_29612,N_29840);
or UO_1560 (O_1560,N_29949,N_29872);
xor UO_1561 (O_1561,N_29535,N_29630);
or UO_1562 (O_1562,N_29995,N_29878);
nor UO_1563 (O_1563,N_29681,N_29508);
or UO_1564 (O_1564,N_29810,N_29659);
nor UO_1565 (O_1565,N_29657,N_29634);
nor UO_1566 (O_1566,N_29519,N_29964);
xnor UO_1567 (O_1567,N_29526,N_29609);
and UO_1568 (O_1568,N_29796,N_29765);
xnor UO_1569 (O_1569,N_29779,N_29541);
or UO_1570 (O_1570,N_29703,N_29508);
or UO_1571 (O_1571,N_29811,N_29619);
xor UO_1572 (O_1572,N_29766,N_29819);
or UO_1573 (O_1573,N_29995,N_29974);
and UO_1574 (O_1574,N_29596,N_29867);
nor UO_1575 (O_1575,N_29951,N_29969);
nor UO_1576 (O_1576,N_29777,N_29616);
nand UO_1577 (O_1577,N_29902,N_29765);
xnor UO_1578 (O_1578,N_29867,N_29877);
nand UO_1579 (O_1579,N_29529,N_29785);
or UO_1580 (O_1580,N_29827,N_29655);
nor UO_1581 (O_1581,N_29533,N_29682);
or UO_1582 (O_1582,N_29572,N_29840);
nand UO_1583 (O_1583,N_29804,N_29641);
nand UO_1584 (O_1584,N_29989,N_29825);
nor UO_1585 (O_1585,N_29872,N_29510);
xor UO_1586 (O_1586,N_29947,N_29864);
nand UO_1587 (O_1587,N_29841,N_29985);
or UO_1588 (O_1588,N_29745,N_29781);
xnor UO_1589 (O_1589,N_29945,N_29911);
nand UO_1590 (O_1590,N_29638,N_29883);
nor UO_1591 (O_1591,N_29952,N_29725);
xnor UO_1592 (O_1592,N_29925,N_29926);
xor UO_1593 (O_1593,N_29501,N_29645);
nand UO_1594 (O_1594,N_29546,N_29537);
and UO_1595 (O_1595,N_29697,N_29650);
and UO_1596 (O_1596,N_29659,N_29680);
nand UO_1597 (O_1597,N_29601,N_29680);
nand UO_1598 (O_1598,N_29992,N_29866);
nand UO_1599 (O_1599,N_29808,N_29978);
nand UO_1600 (O_1600,N_29929,N_29902);
xor UO_1601 (O_1601,N_29566,N_29927);
nand UO_1602 (O_1602,N_29694,N_29610);
nor UO_1603 (O_1603,N_29877,N_29981);
or UO_1604 (O_1604,N_29848,N_29921);
nand UO_1605 (O_1605,N_29977,N_29659);
or UO_1606 (O_1606,N_29973,N_29765);
and UO_1607 (O_1607,N_29525,N_29820);
or UO_1608 (O_1608,N_29752,N_29960);
nand UO_1609 (O_1609,N_29566,N_29957);
xor UO_1610 (O_1610,N_29907,N_29574);
xnor UO_1611 (O_1611,N_29977,N_29693);
and UO_1612 (O_1612,N_29779,N_29631);
nand UO_1613 (O_1613,N_29994,N_29501);
nor UO_1614 (O_1614,N_29878,N_29783);
nor UO_1615 (O_1615,N_29997,N_29766);
or UO_1616 (O_1616,N_29697,N_29879);
nand UO_1617 (O_1617,N_29629,N_29564);
xnor UO_1618 (O_1618,N_29827,N_29905);
xnor UO_1619 (O_1619,N_29531,N_29819);
and UO_1620 (O_1620,N_29874,N_29674);
or UO_1621 (O_1621,N_29727,N_29976);
nor UO_1622 (O_1622,N_29942,N_29879);
nand UO_1623 (O_1623,N_29889,N_29962);
or UO_1624 (O_1624,N_29637,N_29920);
or UO_1625 (O_1625,N_29814,N_29768);
and UO_1626 (O_1626,N_29581,N_29562);
nand UO_1627 (O_1627,N_29772,N_29954);
xor UO_1628 (O_1628,N_29868,N_29704);
or UO_1629 (O_1629,N_29594,N_29541);
or UO_1630 (O_1630,N_29827,N_29748);
xnor UO_1631 (O_1631,N_29860,N_29625);
and UO_1632 (O_1632,N_29784,N_29953);
and UO_1633 (O_1633,N_29882,N_29896);
xor UO_1634 (O_1634,N_29835,N_29581);
xnor UO_1635 (O_1635,N_29896,N_29776);
and UO_1636 (O_1636,N_29695,N_29898);
nand UO_1637 (O_1637,N_29718,N_29721);
xnor UO_1638 (O_1638,N_29986,N_29560);
or UO_1639 (O_1639,N_29982,N_29653);
nand UO_1640 (O_1640,N_29859,N_29604);
or UO_1641 (O_1641,N_29580,N_29978);
nor UO_1642 (O_1642,N_29794,N_29500);
or UO_1643 (O_1643,N_29581,N_29705);
or UO_1644 (O_1644,N_29979,N_29906);
xnor UO_1645 (O_1645,N_29807,N_29992);
or UO_1646 (O_1646,N_29799,N_29902);
nand UO_1647 (O_1647,N_29743,N_29995);
or UO_1648 (O_1648,N_29826,N_29512);
xnor UO_1649 (O_1649,N_29603,N_29625);
xnor UO_1650 (O_1650,N_29509,N_29821);
xnor UO_1651 (O_1651,N_29722,N_29543);
xor UO_1652 (O_1652,N_29846,N_29958);
nor UO_1653 (O_1653,N_29906,N_29841);
or UO_1654 (O_1654,N_29653,N_29884);
xnor UO_1655 (O_1655,N_29860,N_29700);
and UO_1656 (O_1656,N_29683,N_29510);
or UO_1657 (O_1657,N_29509,N_29727);
nor UO_1658 (O_1658,N_29607,N_29863);
and UO_1659 (O_1659,N_29733,N_29779);
and UO_1660 (O_1660,N_29899,N_29698);
nor UO_1661 (O_1661,N_29501,N_29906);
and UO_1662 (O_1662,N_29871,N_29959);
or UO_1663 (O_1663,N_29881,N_29680);
xnor UO_1664 (O_1664,N_29500,N_29522);
and UO_1665 (O_1665,N_29561,N_29597);
and UO_1666 (O_1666,N_29658,N_29884);
nand UO_1667 (O_1667,N_29865,N_29693);
and UO_1668 (O_1668,N_29574,N_29589);
or UO_1669 (O_1669,N_29954,N_29749);
nor UO_1670 (O_1670,N_29701,N_29787);
xnor UO_1671 (O_1671,N_29807,N_29858);
and UO_1672 (O_1672,N_29848,N_29689);
nand UO_1673 (O_1673,N_29692,N_29567);
xor UO_1674 (O_1674,N_29681,N_29625);
nor UO_1675 (O_1675,N_29764,N_29636);
nor UO_1676 (O_1676,N_29864,N_29805);
xnor UO_1677 (O_1677,N_29935,N_29943);
nor UO_1678 (O_1678,N_29561,N_29628);
and UO_1679 (O_1679,N_29612,N_29918);
and UO_1680 (O_1680,N_29843,N_29785);
xor UO_1681 (O_1681,N_29830,N_29549);
nor UO_1682 (O_1682,N_29727,N_29967);
or UO_1683 (O_1683,N_29678,N_29669);
xnor UO_1684 (O_1684,N_29696,N_29560);
nor UO_1685 (O_1685,N_29845,N_29833);
or UO_1686 (O_1686,N_29598,N_29548);
nand UO_1687 (O_1687,N_29728,N_29732);
nor UO_1688 (O_1688,N_29514,N_29634);
nand UO_1689 (O_1689,N_29587,N_29778);
xor UO_1690 (O_1690,N_29824,N_29692);
nand UO_1691 (O_1691,N_29916,N_29621);
or UO_1692 (O_1692,N_29931,N_29567);
nor UO_1693 (O_1693,N_29754,N_29681);
xor UO_1694 (O_1694,N_29636,N_29741);
xnor UO_1695 (O_1695,N_29588,N_29566);
nand UO_1696 (O_1696,N_29984,N_29562);
xnor UO_1697 (O_1697,N_29859,N_29564);
or UO_1698 (O_1698,N_29707,N_29593);
nor UO_1699 (O_1699,N_29879,N_29884);
nand UO_1700 (O_1700,N_29871,N_29519);
nand UO_1701 (O_1701,N_29609,N_29994);
xnor UO_1702 (O_1702,N_29735,N_29649);
xnor UO_1703 (O_1703,N_29792,N_29732);
and UO_1704 (O_1704,N_29623,N_29728);
xor UO_1705 (O_1705,N_29968,N_29893);
nand UO_1706 (O_1706,N_29691,N_29847);
and UO_1707 (O_1707,N_29909,N_29879);
nor UO_1708 (O_1708,N_29987,N_29762);
and UO_1709 (O_1709,N_29663,N_29713);
and UO_1710 (O_1710,N_29992,N_29939);
nand UO_1711 (O_1711,N_29849,N_29882);
nand UO_1712 (O_1712,N_29841,N_29739);
nor UO_1713 (O_1713,N_29860,N_29613);
or UO_1714 (O_1714,N_29556,N_29788);
nand UO_1715 (O_1715,N_29911,N_29768);
nand UO_1716 (O_1716,N_29826,N_29596);
and UO_1717 (O_1717,N_29561,N_29528);
nor UO_1718 (O_1718,N_29573,N_29764);
and UO_1719 (O_1719,N_29787,N_29876);
xnor UO_1720 (O_1720,N_29788,N_29922);
and UO_1721 (O_1721,N_29799,N_29863);
and UO_1722 (O_1722,N_29565,N_29583);
nand UO_1723 (O_1723,N_29701,N_29605);
xor UO_1724 (O_1724,N_29704,N_29544);
or UO_1725 (O_1725,N_29606,N_29665);
nand UO_1726 (O_1726,N_29939,N_29520);
nor UO_1727 (O_1727,N_29915,N_29512);
or UO_1728 (O_1728,N_29546,N_29939);
or UO_1729 (O_1729,N_29562,N_29777);
nor UO_1730 (O_1730,N_29779,N_29706);
nor UO_1731 (O_1731,N_29770,N_29989);
nor UO_1732 (O_1732,N_29663,N_29859);
xor UO_1733 (O_1733,N_29869,N_29509);
or UO_1734 (O_1734,N_29758,N_29922);
and UO_1735 (O_1735,N_29959,N_29684);
nand UO_1736 (O_1736,N_29984,N_29796);
nand UO_1737 (O_1737,N_29771,N_29708);
xnor UO_1738 (O_1738,N_29602,N_29721);
nand UO_1739 (O_1739,N_29898,N_29680);
and UO_1740 (O_1740,N_29891,N_29650);
nand UO_1741 (O_1741,N_29692,N_29577);
nor UO_1742 (O_1742,N_29610,N_29775);
nor UO_1743 (O_1743,N_29804,N_29674);
and UO_1744 (O_1744,N_29787,N_29602);
nor UO_1745 (O_1745,N_29554,N_29678);
nor UO_1746 (O_1746,N_29675,N_29791);
xnor UO_1747 (O_1747,N_29713,N_29668);
and UO_1748 (O_1748,N_29777,N_29630);
nand UO_1749 (O_1749,N_29752,N_29640);
nand UO_1750 (O_1750,N_29929,N_29895);
or UO_1751 (O_1751,N_29692,N_29548);
nor UO_1752 (O_1752,N_29703,N_29962);
or UO_1753 (O_1753,N_29905,N_29950);
nand UO_1754 (O_1754,N_29631,N_29683);
xnor UO_1755 (O_1755,N_29513,N_29904);
and UO_1756 (O_1756,N_29651,N_29748);
xnor UO_1757 (O_1757,N_29599,N_29595);
xor UO_1758 (O_1758,N_29946,N_29647);
and UO_1759 (O_1759,N_29605,N_29571);
nor UO_1760 (O_1760,N_29749,N_29869);
or UO_1761 (O_1761,N_29658,N_29836);
xor UO_1762 (O_1762,N_29902,N_29863);
xor UO_1763 (O_1763,N_29757,N_29563);
nor UO_1764 (O_1764,N_29577,N_29964);
xor UO_1765 (O_1765,N_29740,N_29500);
xnor UO_1766 (O_1766,N_29675,N_29520);
nand UO_1767 (O_1767,N_29575,N_29833);
xor UO_1768 (O_1768,N_29983,N_29893);
xor UO_1769 (O_1769,N_29702,N_29822);
nand UO_1770 (O_1770,N_29575,N_29949);
or UO_1771 (O_1771,N_29745,N_29648);
nand UO_1772 (O_1772,N_29943,N_29934);
xor UO_1773 (O_1773,N_29666,N_29878);
nor UO_1774 (O_1774,N_29655,N_29893);
or UO_1775 (O_1775,N_29645,N_29706);
nand UO_1776 (O_1776,N_29893,N_29585);
nor UO_1777 (O_1777,N_29544,N_29851);
and UO_1778 (O_1778,N_29541,N_29543);
xnor UO_1779 (O_1779,N_29789,N_29669);
nand UO_1780 (O_1780,N_29915,N_29907);
xnor UO_1781 (O_1781,N_29836,N_29873);
nand UO_1782 (O_1782,N_29974,N_29787);
xnor UO_1783 (O_1783,N_29651,N_29521);
nand UO_1784 (O_1784,N_29587,N_29796);
xor UO_1785 (O_1785,N_29521,N_29559);
nor UO_1786 (O_1786,N_29757,N_29616);
and UO_1787 (O_1787,N_29910,N_29504);
or UO_1788 (O_1788,N_29941,N_29766);
nand UO_1789 (O_1789,N_29720,N_29551);
or UO_1790 (O_1790,N_29850,N_29746);
nor UO_1791 (O_1791,N_29724,N_29992);
nor UO_1792 (O_1792,N_29929,N_29689);
xnor UO_1793 (O_1793,N_29751,N_29544);
and UO_1794 (O_1794,N_29642,N_29877);
nor UO_1795 (O_1795,N_29768,N_29560);
or UO_1796 (O_1796,N_29882,N_29729);
nand UO_1797 (O_1797,N_29849,N_29907);
nor UO_1798 (O_1798,N_29658,N_29876);
or UO_1799 (O_1799,N_29676,N_29707);
or UO_1800 (O_1800,N_29787,N_29702);
and UO_1801 (O_1801,N_29798,N_29767);
or UO_1802 (O_1802,N_29710,N_29684);
xor UO_1803 (O_1803,N_29880,N_29695);
nor UO_1804 (O_1804,N_29869,N_29915);
xnor UO_1805 (O_1805,N_29701,N_29872);
and UO_1806 (O_1806,N_29780,N_29755);
and UO_1807 (O_1807,N_29571,N_29630);
xor UO_1808 (O_1808,N_29916,N_29985);
xnor UO_1809 (O_1809,N_29758,N_29944);
nand UO_1810 (O_1810,N_29813,N_29795);
xor UO_1811 (O_1811,N_29877,N_29737);
nor UO_1812 (O_1812,N_29557,N_29546);
nor UO_1813 (O_1813,N_29912,N_29788);
nor UO_1814 (O_1814,N_29631,N_29586);
nor UO_1815 (O_1815,N_29711,N_29574);
xnor UO_1816 (O_1816,N_29836,N_29742);
xor UO_1817 (O_1817,N_29817,N_29946);
nand UO_1818 (O_1818,N_29667,N_29783);
and UO_1819 (O_1819,N_29601,N_29543);
nand UO_1820 (O_1820,N_29777,N_29996);
or UO_1821 (O_1821,N_29626,N_29629);
or UO_1822 (O_1822,N_29710,N_29516);
nand UO_1823 (O_1823,N_29811,N_29646);
and UO_1824 (O_1824,N_29535,N_29771);
or UO_1825 (O_1825,N_29526,N_29879);
xnor UO_1826 (O_1826,N_29584,N_29685);
and UO_1827 (O_1827,N_29891,N_29994);
nand UO_1828 (O_1828,N_29740,N_29938);
nand UO_1829 (O_1829,N_29986,N_29613);
and UO_1830 (O_1830,N_29865,N_29823);
nand UO_1831 (O_1831,N_29582,N_29768);
and UO_1832 (O_1832,N_29907,N_29742);
nor UO_1833 (O_1833,N_29844,N_29914);
xnor UO_1834 (O_1834,N_29514,N_29729);
and UO_1835 (O_1835,N_29813,N_29789);
and UO_1836 (O_1836,N_29976,N_29939);
or UO_1837 (O_1837,N_29581,N_29829);
and UO_1838 (O_1838,N_29513,N_29673);
nor UO_1839 (O_1839,N_29599,N_29694);
or UO_1840 (O_1840,N_29623,N_29527);
nand UO_1841 (O_1841,N_29740,N_29654);
nor UO_1842 (O_1842,N_29922,N_29926);
nor UO_1843 (O_1843,N_29727,N_29835);
nor UO_1844 (O_1844,N_29941,N_29816);
nor UO_1845 (O_1845,N_29854,N_29816);
or UO_1846 (O_1846,N_29580,N_29696);
xor UO_1847 (O_1847,N_29959,N_29826);
xnor UO_1848 (O_1848,N_29732,N_29608);
and UO_1849 (O_1849,N_29773,N_29588);
nand UO_1850 (O_1850,N_29695,N_29616);
nor UO_1851 (O_1851,N_29658,N_29846);
or UO_1852 (O_1852,N_29824,N_29653);
xor UO_1853 (O_1853,N_29745,N_29646);
or UO_1854 (O_1854,N_29830,N_29781);
nand UO_1855 (O_1855,N_29638,N_29998);
xor UO_1856 (O_1856,N_29983,N_29596);
xor UO_1857 (O_1857,N_29862,N_29521);
nor UO_1858 (O_1858,N_29776,N_29914);
and UO_1859 (O_1859,N_29706,N_29600);
or UO_1860 (O_1860,N_29626,N_29779);
and UO_1861 (O_1861,N_29540,N_29651);
nand UO_1862 (O_1862,N_29783,N_29583);
and UO_1863 (O_1863,N_29637,N_29760);
nand UO_1864 (O_1864,N_29573,N_29859);
and UO_1865 (O_1865,N_29649,N_29636);
nand UO_1866 (O_1866,N_29566,N_29913);
nor UO_1867 (O_1867,N_29970,N_29762);
and UO_1868 (O_1868,N_29764,N_29880);
nand UO_1869 (O_1869,N_29780,N_29741);
xnor UO_1870 (O_1870,N_29684,N_29892);
or UO_1871 (O_1871,N_29585,N_29611);
xor UO_1872 (O_1872,N_29635,N_29530);
nand UO_1873 (O_1873,N_29780,N_29550);
and UO_1874 (O_1874,N_29913,N_29667);
xnor UO_1875 (O_1875,N_29975,N_29834);
xnor UO_1876 (O_1876,N_29913,N_29544);
nand UO_1877 (O_1877,N_29628,N_29613);
and UO_1878 (O_1878,N_29923,N_29767);
nor UO_1879 (O_1879,N_29781,N_29697);
xnor UO_1880 (O_1880,N_29752,N_29864);
xnor UO_1881 (O_1881,N_29664,N_29727);
nand UO_1882 (O_1882,N_29522,N_29585);
xnor UO_1883 (O_1883,N_29578,N_29706);
nand UO_1884 (O_1884,N_29766,N_29588);
nand UO_1885 (O_1885,N_29501,N_29750);
or UO_1886 (O_1886,N_29876,N_29992);
xnor UO_1887 (O_1887,N_29882,N_29793);
nand UO_1888 (O_1888,N_29571,N_29872);
nand UO_1889 (O_1889,N_29554,N_29645);
nand UO_1890 (O_1890,N_29920,N_29558);
and UO_1891 (O_1891,N_29819,N_29667);
nand UO_1892 (O_1892,N_29590,N_29553);
nor UO_1893 (O_1893,N_29690,N_29617);
nor UO_1894 (O_1894,N_29537,N_29745);
or UO_1895 (O_1895,N_29707,N_29715);
nand UO_1896 (O_1896,N_29860,N_29977);
nor UO_1897 (O_1897,N_29562,N_29848);
nand UO_1898 (O_1898,N_29506,N_29509);
nand UO_1899 (O_1899,N_29727,N_29535);
nor UO_1900 (O_1900,N_29966,N_29538);
or UO_1901 (O_1901,N_29565,N_29664);
or UO_1902 (O_1902,N_29555,N_29852);
and UO_1903 (O_1903,N_29767,N_29780);
or UO_1904 (O_1904,N_29763,N_29877);
nor UO_1905 (O_1905,N_29826,N_29666);
xor UO_1906 (O_1906,N_29962,N_29785);
nand UO_1907 (O_1907,N_29768,N_29965);
or UO_1908 (O_1908,N_29628,N_29996);
or UO_1909 (O_1909,N_29791,N_29939);
nor UO_1910 (O_1910,N_29860,N_29608);
nand UO_1911 (O_1911,N_29934,N_29946);
nand UO_1912 (O_1912,N_29970,N_29783);
nor UO_1913 (O_1913,N_29700,N_29751);
nand UO_1914 (O_1914,N_29991,N_29916);
and UO_1915 (O_1915,N_29858,N_29675);
nand UO_1916 (O_1916,N_29605,N_29716);
nand UO_1917 (O_1917,N_29929,N_29897);
nor UO_1918 (O_1918,N_29700,N_29789);
nand UO_1919 (O_1919,N_29744,N_29982);
nor UO_1920 (O_1920,N_29955,N_29801);
or UO_1921 (O_1921,N_29825,N_29505);
or UO_1922 (O_1922,N_29548,N_29737);
nor UO_1923 (O_1923,N_29858,N_29629);
or UO_1924 (O_1924,N_29797,N_29676);
nand UO_1925 (O_1925,N_29796,N_29988);
or UO_1926 (O_1926,N_29577,N_29726);
or UO_1927 (O_1927,N_29577,N_29877);
nor UO_1928 (O_1928,N_29713,N_29722);
nor UO_1929 (O_1929,N_29938,N_29836);
nor UO_1930 (O_1930,N_29723,N_29535);
and UO_1931 (O_1931,N_29599,N_29738);
xnor UO_1932 (O_1932,N_29933,N_29944);
xnor UO_1933 (O_1933,N_29784,N_29992);
and UO_1934 (O_1934,N_29948,N_29526);
or UO_1935 (O_1935,N_29616,N_29528);
nor UO_1936 (O_1936,N_29607,N_29883);
and UO_1937 (O_1937,N_29654,N_29764);
or UO_1938 (O_1938,N_29503,N_29868);
or UO_1939 (O_1939,N_29511,N_29766);
xnor UO_1940 (O_1940,N_29605,N_29690);
and UO_1941 (O_1941,N_29712,N_29743);
nand UO_1942 (O_1942,N_29911,N_29618);
or UO_1943 (O_1943,N_29889,N_29518);
nor UO_1944 (O_1944,N_29921,N_29788);
nand UO_1945 (O_1945,N_29505,N_29575);
xor UO_1946 (O_1946,N_29878,N_29737);
or UO_1947 (O_1947,N_29549,N_29712);
xor UO_1948 (O_1948,N_29965,N_29695);
or UO_1949 (O_1949,N_29608,N_29747);
xor UO_1950 (O_1950,N_29520,N_29773);
nor UO_1951 (O_1951,N_29767,N_29633);
nor UO_1952 (O_1952,N_29919,N_29735);
and UO_1953 (O_1953,N_29848,N_29788);
or UO_1954 (O_1954,N_29810,N_29972);
nand UO_1955 (O_1955,N_29782,N_29668);
xnor UO_1956 (O_1956,N_29722,N_29830);
and UO_1957 (O_1957,N_29881,N_29824);
nand UO_1958 (O_1958,N_29612,N_29900);
and UO_1959 (O_1959,N_29861,N_29637);
nor UO_1960 (O_1960,N_29782,N_29974);
nor UO_1961 (O_1961,N_29850,N_29853);
or UO_1962 (O_1962,N_29648,N_29986);
xnor UO_1963 (O_1963,N_29531,N_29731);
nand UO_1964 (O_1964,N_29810,N_29993);
xor UO_1965 (O_1965,N_29746,N_29894);
nand UO_1966 (O_1966,N_29818,N_29992);
nand UO_1967 (O_1967,N_29760,N_29905);
or UO_1968 (O_1968,N_29575,N_29803);
xnor UO_1969 (O_1969,N_29871,N_29728);
xnor UO_1970 (O_1970,N_29921,N_29665);
and UO_1971 (O_1971,N_29659,N_29661);
nor UO_1972 (O_1972,N_29541,N_29636);
nor UO_1973 (O_1973,N_29794,N_29726);
or UO_1974 (O_1974,N_29670,N_29836);
or UO_1975 (O_1975,N_29911,N_29900);
nand UO_1976 (O_1976,N_29881,N_29822);
and UO_1977 (O_1977,N_29946,N_29563);
xor UO_1978 (O_1978,N_29869,N_29889);
or UO_1979 (O_1979,N_29908,N_29682);
and UO_1980 (O_1980,N_29647,N_29656);
nand UO_1981 (O_1981,N_29756,N_29998);
or UO_1982 (O_1982,N_29743,N_29674);
nand UO_1983 (O_1983,N_29746,N_29708);
nand UO_1984 (O_1984,N_29880,N_29729);
nand UO_1985 (O_1985,N_29997,N_29667);
nand UO_1986 (O_1986,N_29744,N_29688);
nor UO_1987 (O_1987,N_29930,N_29976);
and UO_1988 (O_1988,N_29558,N_29797);
or UO_1989 (O_1989,N_29520,N_29535);
and UO_1990 (O_1990,N_29654,N_29838);
nand UO_1991 (O_1991,N_29878,N_29750);
xnor UO_1992 (O_1992,N_29878,N_29953);
and UO_1993 (O_1993,N_29574,N_29961);
xor UO_1994 (O_1994,N_29507,N_29572);
and UO_1995 (O_1995,N_29972,N_29683);
nor UO_1996 (O_1996,N_29509,N_29532);
or UO_1997 (O_1997,N_29567,N_29905);
nor UO_1998 (O_1998,N_29513,N_29719);
and UO_1999 (O_1999,N_29996,N_29670);
or UO_2000 (O_2000,N_29576,N_29520);
nor UO_2001 (O_2001,N_29700,N_29924);
nand UO_2002 (O_2002,N_29867,N_29773);
nand UO_2003 (O_2003,N_29906,N_29924);
and UO_2004 (O_2004,N_29733,N_29877);
or UO_2005 (O_2005,N_29545,N_29798);
or UO_2006 (O_2006,N_29862,N_29688);
and UO_2007 (O_2007,N_29606,N_29860);
and UO_2008 (O_2008,N_29753,N_29675);
xor UO_2009 (O_2009,N_29536,N_29872);
nor UO_2010 (O_2010,N_29881,N_29544);
xor UO_2011 (O_2011,N_29928,N_29920);
nor UO_2012 (O_2012,N_29720,N_29926);
or UO_2013 (O_2013,N_29975,N_29533);
or UO_2014 (O_2014,N_29776,N_29712);
nand UO_2015 (O_2015,N_29641,N_29648);
nor UO_2016 (O_2016,N_29659,N_29634);
xor UO_2017 (O_2017,N_29833,N_29890);
nand UO_2018 (O_2018,N_29772,N_29865);
nand UO_2019 (O_2019,N_29515,N_29893);
nand UO_2020 (O_2020,N_29633,N_29842);
or UO_2021 (O_2021,N_29823,N_29643);
or UO_2022 (O_2022,N_29812,N_29973);
and UO_2023 (O_2023,N_29968,N_29509);
nor UO_2024 (O_2024,N_29968,N_29751);
xor UO_2025 (O_2025,N_29568,N_29927);
nor UO_2026 (O_2026,N_29981,N_29736);
or UO_2027 (O_2027,N_29703,N_29941);
or UO_2028 (O_2028,N_29563,N_29959);
nand UO_2029 (O_2029,N_29579,N_29924);
nor UO_2030 (O_2030,N_29700,N_29997);
and UO_2031 (O_2031,N_29616,N_29765);
and UO_2032 (O_2032,N_29868,N_29955);
or UO_2033 (O_2033,N_29707,N_29861);
and UO_2034 (O_2034,N_29969,N_29500);
nand UO_2035 (O_2035,N_29930,N_29803);
and UO_2036 (O_2036,N_29675,N_29607);
nor UO_2037 (O_2037,N_29702,N_29901);
and UO_2038 (O_2038,N_29907,N_29674);
and UO_2039 (O_2039,N_29680,N_29820);
nand UO_2040 (O_2040,N_29788,N_29942);
nand UO_2041 (O_2041,N_29897,N_29802);
and UO_2042 (O_2042,N_29685,N_29776);
nand UO_2043 (O_2043,N_29918,N_29845);
xnor UO_2044 (O_2044,N_29986,N_29755);
or UO_2045 (O_2045,N_29879,N_29521);
and UO_2046 (O_2046,N_29684,N_29540);
nor UO_2047 (O_2047,N_29939,N_29631);
nand UO_2048 (O_2048,N_29645,N_29613);
nand UO_2049 (O_2049,N_29888,N_29835);
nor UO_2050 (O_2050,N_29504,N_29564);
nor UO_2051 (O_2051,N_29700,N_29680);
or UO_2052 (O_2052,N_29931,N_29714);
or UO_2053 (O_2053,N_29817,N_29604);
xor UO_2054 (O_2054,N_29954,N_29530);
nor UO_2055 (O_2055,N_29694,N_29550);
or UO_2056 (O_2056,N_29752,N_29756);
and UO_2057 (O_2057,N_29910,N_29501);
xnor UO_2058 (O_2058,N_29720,N_29972);
or UO_2059 (O_2059,N_29857,N_29755);
or UO_2060 (O_2060,N_29895,N_29786);
nor UO_2061 (O_2061,N_29708,N_29865);
nand UO_2062 (O_2062,N_29515,N_29596);
nor UO_2063 (O_2063,N_29905,N_29614);
nand UO_2064 (O_2064,N_29655,N_29739);
or UO_2065 (O_2065,N_29950,N_29635);
and UO_2066 (O_2066,N_29775,N_29589);
xor UO_2067 (O_2067,N_29565,N_29689);
nor UO_2068 (O_2068,N_29929,N_29588);
or UO_2069 (O_2069,N_29732,N_29846);
and UO_2070 (O_2070,N_29936,N_29743);
xnor UO_2071 (O_2071,N_29532,N_29870);
and UO_2072 (O_2072,N_29541,N_29669);
and UO_2073 (O_2073,N_29576,N_29694);
xor UO_2074 (O_2074,N_29796,N_29845);
nor UO_2075 (O_2075,N_29891,N_29761);
and UO_2076 (O_2076,N_29841,N_29687);
nor UO_2077 (O_2077,N_29737,N_29859);
nand UO_2078 (O_2078,N_29978,N_29888);
or UO_2079 (O_2079,N_29952,N_29656);
nor UO_2080 (O_2080,N_29888,N_29876);
nor UO_2081 (O_2081,N_29510,N_29645);
nand UO_2082 (O_2082,N_29897,N_29698);
and UO_2083 (O_2083,N_29648,N_29904);
nand UO_2084 (O_2084,N_29763,N_29671);
xnor UO_2085 (O_2085,N_29864,N_29762);
nand UO_2086 (O_2086,N_29977,N_29513);
or UO_2087 (O_2087,N_29578,N_29544);
nand UO_2088 (O_2088,N_29852,N_29611);
nand UO_2089 (O_2089,N_29944,N_29556);
xor UO_2090 (O_2090,N_29853,N_29695);
nand UO_2091 (O_2091,N_29979,N_29935);
nand UO_2092 (O_2092,N_29574,N_29861);
nor UO_2093 (O_2093,N_29585,N_29667);
or UO_2094 (O_2094,N_29786,N_29651);
nor UO_2095 (O_2095,N_29965,N_29636);
nand UO_2096 (O_2096,N_29606,N_29621);
xnor UO_2097 (O_2097,N_29734,N_29552);
nor UO_2098 (O_2098,N_29693,N_29673);
and UO_2099 (O_2099,N_29954,N_29717);
nand UO_2100 (O_2100,N_29832,N_29720);
nor UO_2101 (O_2101,N_29830,N_29683);
and UO_2102 (O_2102,N_29878,N_29648);
nand UO_2103 (O_2103,N_29975,N_29893);
nor UO_2104 (O_2104,N_29913,N_29756);
nor UO_2105 (O_2105,N_29847,N_29652);
nor UO_2106 (O_2106,N_29815,N_29945);
nor UO_2107 (O_2107,N_29753,N_29605);
xnor UO_2108 (O_2108,N_29878,N_29577);
nor UO_2109 (O_2109,N_29798,N_29980);
and UO_2110 (O_2110,N_29884,N_29744);
nor UO_2111 (O_2111,N_29773,N_29721);
nand UO_2112 (O_2112,N_29970,N_29610);
nand UO_2113 (O_2113,N_29995,N_29912);
and UO_2114 (O_2114,N_29536,N_29750);
nand UO_2115 (O_2115,N_29614,N_29598);
xor UO_2116 (O_2116,N_29782,N_29890);
nor UO_2117 (O_2117,N_29801,N_29575);
and UO_2118 (O_2118,N_29993,N_29997);
nand UO_2119 (O_2119,N_29693,N_29818);
or UO_2120 (O_2120,N_29720,N_29931);
or UO_2121 (O_2121,N_29975,N_29839);
nand UO_2122 (O_2122,N_29654,N_29549);
xor UO_2123 (O_2123,N_29529,N_29911);
and UO_2124 (O_2124,N_29735,N_29955);
or UO_2125 (O_2125,N_29904,N_29569);
nor UO_2126 (O_2126,N_29971,N_29606);
xor UO_2127 (O_2127,N_29841,N_29568);
nand UO_2128 (O_2128,N_29980,N_29987);
xor UO_2129 (O_2129,N_29726,N_29634);
nor UO_2130 (O_2130,N_29808,N_29644);
xnor UO_2131 (O_2131,N_29550,N_29908);
xor UO_2132 (O_2132,N_29655,N_29667);
nor UO_2133 (O_2133,N_29660,N_29526);
xor UO_2134 (O_2134,N_29760,N_29880);
or UO_2135 (O_2135,N_29558,N_29620);
nand UO_2136 (O_2136,N_29653,N_29683);
nand UO_2137 (O_2137,N_29960,N_29703);
or UO_2138 (O_2138,N_29738,N_29530);
and UO_2139 (O_2139,N_29886,N_29936);
and UO_2140 (O_2140,N_29607,N_29657);
and UO_2141 (O_2141,N_29590,N_29517);
and UO_2142 (O_2142,N_29515,N_29789);
or UO_2143 (O_2143,N_29958,N_29967);
xor UO_2144 (O_2144,N_29623,N_29957);
or UO_2145 (O_2145,N_29577,N_29530);
nor UO_2146 (O_2146,N_29552,N_29897);
xor UO_2147 (O_2147,N_29908,N_29806);
or UO_2148 (O_2148,N_29812,N_29967);
nand UO_2149 (O_2149,N_29987,N_29727);
xnor UO_2150 (O_2150,N_29745,N_29857);
xor UO_2151 (O_2151,N_29865,N_29572);
nand UO_2152 (O_2152,N_29644,N_29738);
nand UO_2153 (O_2153,N_29826,N_29595);
or UO_2154 (O_2154,N_29740,N_29990);
nor UO_2155 (O_2155,N_29650,N_29550);
xor UO_2156 (O_2156,N_29734,N_29899);
nor UO_2157 (O_2157,N_29654,N_29773);
nor UO_2158 (O_2158,N_29572,N_29795);
and UO_2159 (O_2159,N_29739,N_29533);
nor UO_2160 (O_2160,N_29502,N_29620);
nand UO_2161 (O_2161,N_29935,N_29625);
xnor UO_2162 (O_2162,N_29521,N_29947);
nand UO_2163 (O_2163,N_29900,N_29577);
xnor UO_2164 (O_2164,N_29712,N_29771);
or UO_2165 (O_2165,N_29682,N_29907);
xnor UO_2166 (O_2166,N_29942,N_29588);
and UO_2167 (O_2167,N_29984,N_29906);
or UO_2168 (O_2168,N_29926,N_29730);
nor UO_2169 (O_2169,N_29822,N_29760);
nor UO_2170 (O_2170,N_29778,N_29630);
or UO_2171 (O_2171,N_29758,N_29734);
or UO_2172 (O_2172,N_29998,N_29847);
xnor UO_2173 (O_2173,N_29846,N_29745);
xnor UO_2174 (O_2174,N_29745,N_29507);
xor UO_2175 (O_2175,N_29988,N_29765);
and UO_2176 (O_2176,N_29652,N_29792);
or UO_2177 (O_2177,N_29677,N_29586);
nor UO_2178 (O_2178,N_29922,N_29851);
or UO_2179 (O_2179,N_29861,N_29940);
nor UO_2180 (O_2180,N_29552,N_29845);
xnor UO_2181 (O_2181,N_29551,N_29951);
nor UO_2182 (O_2182,N_29833,N_29815);
nor UO_2183 (O_2183,N_29845,N_29756);
xor UO_2184 (O_2184,N_29927,N_29720);
or UO_2185 (O_2185,N_29777,N_29582);
xor UO_2186 (O_2186,N_29671,N_29719);
xor UO_2187 (O_2187,N_29810,N_29875);
or UO_2188 (O_2188,N_29970,N_29928);
nand UO_2189 (O_2189,N_29731,N_29604);
and UO_2190 (O_2190,N_29849,N_29520);
or UO_2191 (O_2191,N_29858,N_29836);
nand UO_2192 (O_2192,N_29504,N_29865);
or UO_2193 (O_2193,N_29932,N_29766);
nand UO_2194 (O_2194,N_29590,N_29522);
nor UO_2195 (O_2195,N_29682,N_29987);
xnor UO_2196 (O_2196,N_29609,N_29525);
xor UO_2197 (O_2197,N_29883,N_29522);
and UO_2198 (O_2198,N_29625,N_29967);
nand UO_2199 (O_2199,N_29558,N_29743);
and UO_2200 (O_2200,N_29904,N_29923);
nor UO_2201 (O_2201,N_29641,N_29992);
nor UO_2202 (O_2202,N_29659,N_29575);
or UO_2203 (O_2203,N_29937,N_29517);
xnor UO_2204 (O_2204,N_29863,N_29660);
nor UO_2205 (O_2205,N_29805,N_29657);
and UO_2206 (O_2206,N_29788,N_29846);
nor UO_2207 (O_2207,N_29551,N_29835);
or UO_2208 (O_2208,N_29816,N_29807);
nand UO_2209 (O_2209,N_29966,N_29857);
or UO_2210 (O_2210,N_29691,N_29864);
or UO_2211 (O_2211,N_29709,N_29511);
nand UO_2212 (O_2212,N_29972,N_29532);
nor UO_2213 (O_2213,N_29770,N_29809);
or UO_2214 (O_2214,N_29988,N_29878);
nand UO_2215 (O_2215,N_29987,N_29730);
nand UO_2216 (O_2216,N_29934,N_29838);
and UO_2217 (O_2217,N_29764,N_29693);
or UO_2218 (O_2218,N_29821,N_29738);
nand UO_2219 (O_2219,N_29684,N_29725);
nand UO_2220 (O_2220,N_29575,N_29978);
xor UO_2221 (O_2221,N_29742,N_29770);
xnor UO_2222 (O_2222,N_29626,N_29859);
nor UO_2223 (O_2223,N_29602,N_29643);
nor UO_2224 (O_2224,N_29804,N_29602);
or UO_2225 (O_2225,N_29684,N_29685);
nand UO_2226 (O_2226,N_29996,N_29763);
and UO_2227 (O_2227,N_29788,N_29588);
xor UO_2228 (O_2228,N_29838,N_29983);
nor UO_2229 (O_2229,N_29518,N_29970);
xnor UO_2230 (O_2230,N_29668,N_29971);
nor UO_2231 (O_2231,N_29597,N_29892);
and UO_2232 (O_2232,N_29630,N_29813);
nand UO_2233 (O_2233,N_29967,N_29769);
nor UO_2234 (O_2234,N_29657,N_29715);
or UO_2235 (O_2235,N_29540,N_29539);
xor UO_2236 (O_2236,N_29605,N_29747);
and UO_2237 (O_2237,N_29994,N_29887);
xnor UO_2238 (O_2238,N_29764,N_29939);
nand UO_2239 (O_2239,N_29834,N_29919);
or UO_2240 (O_2240,N_29856,N_29743);
nand UO_2241 (O_2241,N_29598,N_29845);
nand UO_2242 (O_2242,N_29668,N_29601);
and UO_2243 (O_2243,N_29731,N_29842);
nor UO_2244 (O_2244,N_29527,N_29616);
nor UO_2245 (O_2245,N_29500,N_29799);
nor UO_2246 (O_2246,N_29900,N_29817);
xor UO_2247 (O_2247,N_29650,N_29773);
or UO_2248 (O_2248,N_29913,N_29551);
xnor UO_2249 (O_2249,N_29895,N_29642);
nor UO_2250 (O_2250,N_29511,N_29909);
nand UO_2251 (O_2251,N_29734,N_29990);
and UO_2252 (O_2252,N_29782,N_29661);
nor UO_2253 (O_2253,N_29608,N_29840);
xnor UO_2254 (O_2254,N_29816,N_29637);
xnor UO_2255 (O_2255,N_29615,N_29824);
nand UO_2256 (O_2256,N_29987,N_29633);
xnor UO_2257 (O_2257,N_29850,N_29916);
nand UO_2258 (O_2258,N_29805,N_29775);
xnor UO_2259 (O_2259,N_29505,N_29826);
or UO_2260 (O_2260,N_29615,N_29651);
or UO_2261 (O_2261,N_29887,N_29941);
nor UO_2262 (O_2262,N_29708,N_29514);
nand UO_2263 (O_2263,N_29876,N_29910);
or UO_2264 (O_2264,N_29741,N_29941);
nand UO_2265 (O_2265,N_29984,N_29986);
xnor UO_2266 (O_2266,N_29680,N_29511);
nand UO_2267 (O_2267,N_29681,N_29606);
nand UO_2268 (O_2268,N_29504,N_29893);
xor UO_2269 (O_2269,N_29641,N_29704);
or UO_2270 (O_2270,N_29574,N_29668);
xor UO_2271 (O_2271,N_29533,N_29904);
and UO_2272 (O_2272,N_29548,N_29780);
or UO_2273 (O_2273,N_29995,N_29557);
or UO_2274 (O_2274,N_29883,N_29684);
nand UO_2275 (O_2275,N_29841,N_29958);
or UO_2276 (O_2276,N_29546,N_29948);
and UO_2277 (O_2277,N_29947,N_29663);
and UO_2278 (O_2278,N_29663,N_29965);
xnor UO_2279 (O_2279,N_29707,N_29579);
or UO_2280 (O_2280,N_29954,N_29955);
nand UO_2281 (O_2281,N_29904,N_29850);
or UO_2282 (O_2282,N_29907,N_29992);
or UO_2283 (O_2283,N_29995,N_29851);
and UO_2284 (O_2284,N_29682,N_29820);
xnor UO_2285 (O_2285,N_29527,N_29650);
nor UO_2286 (O_2286,N_29535,N_29847);
nor UO_2287 (O_2287,N_29903,N_29531);
or UO_2288 (O_2288,N_29993,N_29645);
nor UO_2289 (O_2289,N_29982,N_29805);
nor UO_2290 (O_2290,N_29848,N_29836);
nand UO_2291 (O_2291,N_29920,N_29710);
nor UO_2292 (O_2292,N_29655,N_29789);
or UO_2293 (O_2293,N_29952,N_29772);
nor UO_2294 (O_2294,N_29829,N_29973);
or UO_2295 (O_2295,N_29556,N_29636);
or UO_2296 (O_2296,N_29955,N_29902);
and UO_2297 (O_2297,N_29595,N_29825);
xnor UO_2298 (O_2298,N_29871,N_29955);
nor UO_2299 (O_2299,N_29804,N_29598);
and UO_2300 (O_2300,N_29744,N_29524);
nor UO_2301 (O_2301,N_29871,N_29774);
xnor UO_2302 (O_2302,N_29742,N_29739);
nor UO_2303 (O_2303,N_29628,N_29767);
nor UO_2304 (O_2304,N_29732,N_29807);
nand UO_2305 (O_2305,N_29873,N_29736);
nor UO_2306 (O_2306,N_29834,N_29989);
nand UO_2307 (O_2307,N_29887,N_29966);
nor UO_2308 (O_2308,N_29662,N_29653);
xor UO_2309 (O_2309,N_29791,N_29652);
xor UO_2310 (O_2310,N_29839,N_29551);
nor UO_2311 (O_2311,N_29780,N_29603);
or UO_2312 (O_2312,N_29719,N_29923);
xnor UO_2313 (O_2313,N_29990,N_29603);
nor UO_2314 (O_2314,N_29601,N_29958);
and UO_2315 (O_2315,N_29925,N_29651);
xnor UO_2316 (O_2316,N_29605,N_29759);
or UO_2317 (O_2317,N_29816,N_29812);
or UO_2318 (O_2318,N_29698,N_29963);
nor UO_2319 (O_2319,N_29890,N_29844);
or UO_2320 (O_2320,N_29771,N_29582);
nor UO_2321 (O_2321,N_29536,N_29767);
and UO_2322 (O_2322,N_29982,N_29662);
and UO_2323 (O_2323,N_29739,N_29956);
nor UO_2324 (O_2324,N_29864,N_29626);
and UO_2325 (O_2325,N_29673,N_29919);
xnor UO_2326 (O_2326,N_29695,N_29648);
nand UO_2327 (O_2327,N_29622,N_29595);
nor UO_2328 (O_2328,N_29767,N_29751);
or UO_2329 (O_2329,N_29792,N_29856);
nor UO_2330 (O_2330,N_29646,N_29929);
or UO_2331 (O_2331,N_29761,N_29699);
nand UO_2332 (O_2332,N_29911,N_29820);
nor UO_2333 (O_2333,N_29621,N_29573);
or UO_2334 (O_2334,N_29757,N_29961);
nor UO_2335 (O_2335,N_29534,N_29862);
nor UO_2336 (O_2336,N_29639,N_29606);
and UO_2337 (O_2337,N_29739,N_29558);
nand UO_2338 (O_2338,N_29794,N_29954);
xor UO_2339 (O_2339,N_29741,N_29971);
xnor UO_2340 (O_2340,N_29844,N_29982);
or UO_2341 (O_2341,N_29854,N_29818);
xnor UO_2342 (O_2342,N_29502,N_29842);
or UO_2343 (O_2343,N_29881,N_29602);
xor UO_2344 (O_2344,N_29964,N_29659);
nand UO_2345 (O_2345,N_29618,N_29929);
and UO_2346 (O_2346,N_29975,N_29512);
nand UO_2347 (O_2347,N_29865,N_29688);
nand UO_2348 (O_2348,N_29585,N_29750);
xnor UO_2349 (O_2349,N_29895,N_29721);
nor UO_2350 (O_2350,N_29511,N_29841);
and UO_2351 (O_2351,N_29647,N_29986);
or UO_2352 (O_2352,N_29711,N_29514);
nor UO_2353 (O_2353,N_29604,N_29584);
and UO_2354 (O_2354,N_29614,N_29552);
xor UO_2355 (O_2355,N_29932,N_29500);
and UO_2356 (O_2356,N_29520,N_29886);
xor UO_2357 (O_2357,N_29819,N_29977);
nand UO_2358 (O_2358,N_29933,N_29910);
xnor UO_2359 (O_2359,N_29646,N_29719);
and UO_2360 (O_2360,N_29967,N_29517);
and UO_2361 (O_2361,N_29809,N_29629);
or UO_2362 (O_2362,N_29913,N_29770);
and UO_2363 (O_2363,N_29788,N_29851);
xor UO_2364 (O_2364,N_29709,N_29603);
or UO_2365 (O_2365,N_29564,N_29805);
xor UO_2366 (O_2366,N_29800,N_29661);
or UO_2367 (O_2367,N_29518,N_29902);
nand UO_2368 (O_2368,N_29555,N_29622);
nand UO_2369 (O_2369,N_29701,N_29972);
nand UO_2370 (O_2370,N_29651,N_29731);
and UO_2371 (O_2371,N_29535,N_29812);
xnor UO_2372 (O_2372,N_29520,N_29934);
nand UO_2373 (O_2373,N_29609,N_29502);
and UO_2374 (O_2374,N_29888,N_29547);
and UO_2375 (O_2375,N_29756,N_29972);
or UO_2376 (O_2376,N_29514,N_29919);
nand UO_2377 (O_2377,N_29867,N_29736);
xor UO_2378 (O_2378,N_29937,N_29685);
or UO_2379 (O_2379,N_29866,N_29740);
or UO_2380 (O_2380,N_29778,N_29681);
and UO_2381 (O_2381,N_29740,N_29630);
xnor UO_2382 (O_2382,N_29937,N_29924);
xor UO_2383 (O_2383,N_29640,N_29724);
xor UO_2384 (O_2384,N_29994,N_29967);
nor UO_2385 (O_2385,N_29511,N_29813);
nand UO_2386 (O_2386,N_29760,N_29907);
nor UO_2387 (O_2387,N_29935,N_29666);
nand UO_2388 (O_2388,N_29742,N_29673);
nand UO_2389 (O_2389,N_29821,N_29748);
nand UO_2390 (O_2390,N_29558,N_29824);
nand UO_2391 (O_2391,N_29768,N_29895);
nand UO_2392 (O_2392,N_29673,N_29631);
or UO_2393 (O_2393,N_29925,N_29566);
or UO_2394 (O_2394,N_29527,N_29597);
nor UO_2395 (O_2395,N_29517,N_29943);
nand UO_2396 (O_2396,N_29838,N_29642);
or UO_2397 (O_2397,N_29910,N_29595);
nand UO_2398 (O_2398,N_29803,N_29670);
nand UO_2399 (O_2399,N_29806,N_29761);
xor UO_2400 (O_2400,N_29866,N_29579);
xnor UO_2401 (O_2401,N_29592,N_29973);
nand UO_2402 (O_2402,N_29628,N_29965);
xor UO_2403 (O_2403,N_29983,N_29895);
xor UO_2404 (O_2404,N_29711,N_29570);
or UO_2405 (O_2405,N_29780,N_29511);
nor UO_2406 (O_2406,N_29714,N_29622);
nor UO_2407 (O_2407,N_29756,N_29706);
and UO_2408 (O_2408,N_29866,N_29936);
nor UO_2409 (O_2409,N_29653,N_29868);
and UO_2410 (O_2410,N_29708,N_29726);
nand UO_2411 (O_2411,N_29578,N_29678);
or UO_2412 (O_2412,N_29612,N_29995);
xnor UO_2413 (O_2413,N_29534,N_29522);
nor UO_2414 (O_2414,N_29714,N_29579);
nor UO_2415 (O_2415,N_29530,N_29719);
xnor UO_2416 (O_2416,N_29907,N_29670);
xnor UO_2417 (O_2417,N_29995,N_29822);
nor UO_2418 (O_2418,N_29860,N_29719);
and UO_2419 (O_2419,N_29677,N_29811);
xor UO_2420 (O_2420,N_29601,N_29700);
and UO_2421 (O_2421,N_29978,N_29530);
nor UO_2422 (O_2422,N_29804,N_29569);
xnor UO_2423 (O_2423,N_29568,N_29850);
and UO_2424 (O_2424,N_29967,N_29975);
nand UO_2425 (O_2425,N_29984,N_29845);
nand UO_2426 (O_2426,N_29919,N_29945);
xnor UO_2427 (O_2427,N_29531,N_29675);
nor UO_2428 (O_2428,N_29775,N_29803);
and UO_2429 (O_2429,N_29954,N_29502);
nand UO_2430 (O_2430,N_29782,N_29686);
or UO_2431 (O_2431,N_29565,N_29884);
xnor UO_2432 (O_2432,N_29553,N_29547);
or UO_2433 (O_2433,N_29731,N_29564);
nor UO_2434 (O_2434,N_29915,N_29830);
nand UO_2435 (O_2435,N_29823,N_29994);
nand UO_2436 (O_2436,N_29976,N_29573);
xnor UO_2437 (O_2437,N_29944,N_29504);
and UO_2438 (O_2438,N_29546,N_29841);
or UO_2439 (O_2439,N_29951,N_29545);
xnor UO_2440 (O_2440,N_29888,N_29517);
nor UO_2441 (O_2441,N_29568,N_29872);
xor UO_2442 (O_2442,N_29726,N_29926);
or UO_2443 (O_2443,N_29719,N_29751);
or UO_2444 (O_2444,N_29722,N_29634);
or UO_2445 (O_2445,N_29621,N_29794);
xnor UO_2446 (O_2446,N_29681,N_29918);
or UO_2447 (O_2447,N_29937,N_29778);
xnor UO_2448 (O_2448,N_29770,N_29803);
nor UO_2449 (O_2449,N_29859,N_29846);
and UO_2450 (O_2450,N_29957,N_29563);
or UO_2451 (O_2451,N_29646,N_29557);
and UO_2452 (O_2452,N_29563,N_29760);
xor UO_2453 (O_2453,N_29896,N_29711);
nor UO_2454 (O_2454,N_29731,N_29716);
or UO_2455 (O_2455,N_29898,N_29530);
xnor UO_2456 (O_2456,N_29697,N_29671);
nand UO_2457 (O_2457,N_29869,N_29520);
nand UO_2458 (O_2458,N_29521,N_29794);
xor UO_2459 (O_2459,N_29551,N_29892);
xor UO_2460 (O_2460,N_29999,N_29544);
nand UO_2461 (O_2461,N_29809,N_29910);
or UO_2462 (O_2462,N_29660,N_29945);
nor UO_2463 (O_2463,N_29875,N_29847);
nor UO_2464 (O_2464,N_29863,N_29619);
nor UO_2465 (O_2465,N_29659,N_29738);
or UO_2466 (O_2466,N_29792,N_29528);
xor UO_2467 (O_2467,N_29952,N_29828);
and UO_2468 (O_2468,N_29578,N_29973);
and UO_2469 (O_2469,N_29816,N_29539);
nor UO_2470 (O_2470,N_29936,N_29975);
or UO_2471 (O_2471,N_29955,N_29880);
nor UO_2472 (O_2472,N_29932,N_29788);
or UO_2473 (O_2473,N_29617,N_29917);
nor UO_2474 (O_2474,N_29791,N_29760);
and UO_2475 (O_2475,N_29620,N_29888);
xnor UO_2476 (O_2476,N_29934,N_29589);
xnor UO_2477 (O_2477,N_29932,N_29534);
and UO_2478 (O_2478,N_29763,N_29864);
and UO_2479 (O_2479,N_29968,N_29780);
or UO_2480 (O_2480,N_29671,N_29910);
nor UO_2481 (O_2481,N_29564,N_29706);
nor UO_2482 (O_2482,N_29576,N_29556);
nor UO_2483 (O_2483,N_29534,N_29963);
nand UO_2484 (O_2484,N_29955,N_29737);
or UO_2485 (O_2485,N_29878,N_29532);
nand UO_2486 (O_2486,N_29981,N_29783);
or UO_2487 (O_2487,N_29911,N_29946);
nor UO_2488 (O_2488,N_29678,N_29803);
and UO_2489 (O_2489,N_29952,N_29590);
or UO_2490 (O_2490,N_29810,N_29675);
xnor UO_2491 (O_2491,N_29809,N_29657);
or UO_2492 (O_2492,N_29902,N_29971);
and UO_2493 (O_2493,N_29529,N_29692);
and UO_2494 (O_2494,N_29826,N_29910);
nor UO_2495 (O_2495,N_29952,N_29557);
or UO_2496 (O_2496,N_29604,N_29803);
nand UO_2497 (O_2497,N_29684,N_29586);
xor UO_2498 (O_2498,N_29872,N_29937);
or UO_2499 (O_2499,N_29626,N_29886);
nor UO_2500 (O_2500,N_29629,N_29707);
nor UO_2501 (O_2501,N_29997,N_29627);
or UO_2502 (O_2502,N_29711,N_29746);
nor UO_2503 (O_2503,N_29755,N_29584);
and UO_2504 (O_2504,N_29881,N_29549);
and UO_2505 (O_2505,N_29948,N_29641);
and UO_2506 (O_2506,N_29847,N_29522);
and UO_2507 (O_2507,N_29920,N_29974);
nand UO_2508 (O_2508,N_29631,N_29773);
nand UO_2509 (O_2509,N_29848,N_29698);
and UO_2510 (O_2510,N_29949,N_29914);
nand UO_2511 (O_2511,N_29534,N_29665);
or UO_2512 (O_2512,N_29538,N_29763);
nand UO_2513 (O_2513,N_29968,N_29512);
or UO_2514 (O_2514,N_29739,N_29697);
xnor UO_2515 (O_2515,N_29665,N_29780);
or UO_2516 (O_2516,N_29578,N_29944);
xnor UO_2517 (O_2517,N_29911,N_29742);
and UO_2518 (O_2518,N_29720,N_29614);
nor UO_2519 (O_2519,N_29945,N_29765);
and UO_2520 (O_2520,N_29755,N_29825);
nor UO_2521 (O_2521,N_29983,N_29757);
xnor UO_2522 (O_2522,N_29639,N_29750);
nand UO_2523 (O_2523,N_29857,N_29790);
nand UO_2524 (O_2524,N_29736,N_29774);
xor UO_2525 (O_2525,N_29527,N_29694);
and UO_2526 (O_2526,N_29820,N_29671);
and UO_2527 (O_2527,N_29787,N_29814);
or UO_2528 (O_2528,N_29657,N_29551);
nor UO_2529 (O_2529,N_29729,N_29787);
xnor UO_2530 (O_2530,N_29720,N_29890);
nand UO_2531 (O_2531,N_29954,N_29548);
or UO_2532 (O_2532,N_29712,N_29709);
and UO_2533 (O_2533,N_29676,N_29683);
nand UO_2534 (O_2534,N_29536,N_29506);
or UO_2535 (O_2535,N_29819,N_29915);
nor UO_2536 (O_2536,N_29550,N_29623);
nand UO_2537 (O_2537,N_29681,N_29886);
or UO_2538 (O_2538,N_29913,N_29714);
nand UO_2539 (O_2539,N_29999,N_29823);
nor UO_2540 (O_2540,N_29728,N_29528);
nand UO_2541 (O_2541,N_29774,N_29906);
nand UO_2542 (O_2542,N_29824,N_29880);
nand UO_2543 (O_2543,N_29863,N_29652);
nand UO_2544 (O_2544,N_29687,N_29811);
xor UO_2545 (O_2545,N_29554,N_29560);
xnor UO_2546 (O_2546,N_29873,N_29864);
xnor UO_2547 (O_2547,N_29600,N_29715);
nand UO_2548 (O_2548,N_29784,N_29673);
and UO_2549 (O_2549,N_29757,N_29804);
or UO_2550 (O_2550,N_29895,N_29692);
and UO_2551 (O_2551,N_29847,N_29800);
nor UO_2552 (O_2552,N_29947,N_29690);
xnor UO_2553 (O_2553,N_29580,N_29859);
nor UO_2554 (O_2554,N_29956,N_29673);
nor UO_2555 (O_2555,N_29702,N_29524);
xor UO_2556 (O_2556,N_29614,N_29829);
or UO_2557 (O_2557,N_29608,N_29922);
xnor UO_2558 (O_2558,N_29612,N_29645);
nor UO_2559 (O_2559,N_29500,N_29770);
xnor UO_2560 (O_2560,N_29948,N_29867);
or UO_2561 (O_2561,N_29736,N_29606);
nand UO_2562 (O_2562,N_29599,N_29741);
and UO_2563 (O_2563,N_29831,N_29843);
nand UO_2564 (O_2564,N_29716,N_29995);
nor UO_2565 (O_2565,N_29829,N_29505);
or UO_2566 (O_2566,N_29734,N_29994);
xor UO_2567 (O_2567,N_29786,N_29682);
nor UO_2568 (O_2568,N_29923,N_29814);
nor UO_2569 (O_2569,N_29637,N_29669);
or UO_2570 (O_2570,N_29713,N_29875);
nor UO_2571 (O_2571,N_29611,N_29613);
nor UO_2572 (O_2572,N_29661,N_29701);
or UO_2573 (O_2573,N_29799,N_29943);
and UO_2574 (O_2574,N_29868,N_29631);
and UO_2575 (O_2575,N_29984,N_29930);
xnor UO_2576 (O_2576,N_29930,N_29591);
and UO_2577 (O_2577,N_29770,N_29646);
nand UO_2578 (O_2578,N_29604,N_29665);
nand UO_2579 (O_2579,N_29683,N_29884);
or UO_2580 (O_2580,N_29947,N_29545);
and UO_2581 (O_2581,N_29742,N_29599);
or UO_2582 (O_2582,N_29626,N_29568);
xor UO_2583 (O_2583,N_29897,N_29531);
nand UO_2584 (O_2584,N_29738,N_29510);
xnor UO_2585 (O_2585,N_29976,N_29975);
and UO_2586 (O_2586,N_29656,N_29760);
or UO_2587 (O_2587,N_29815,N_29782);
xnor UO_2588 (O_2588,N_29943,N_29697);
xor UO_2589 (O_2589,N_29724,N_29524);
and UO_2590 (O_2590,N_29846,N_29538);
xor UO_2591 (O_2591,N_29691,N_29591);
xnor UO_2592 (O_2592,N_29747,N_29737);
xor UO_2593 (O_2593,N_29750,N_29903);
or UO_2594 (O_2594,N_29780,N_29923);
or UO_2595 (O_2595,N_29508,N_29981);
nand UO_2596 (O_2596,N_29984,N_29793);
nor UO_2597 (O_2597,N_29929,N_29706);
nand UO_2598 (O_2598,N_29508,N_29828);
nand UO_2599 (O_2599,N_29835,N_29725);
xnor UO_2600 (O_2600,N_29585,N_29511);
xnor UO_2601 (O_2601,N_29672,N_29649);
nand UO_2602 (O_2602,N_29842,N_29931);
or UO_2603 (O_2603,N_29968,N_29595);
nand UO_2604 (O_2604,N_29631,N_29598);
xor UO_2605 (O_2605,N_29575,N_29576);
nand UO_2606 (O_2606,N_29582,N_29669);
or UO_2607 (O_2607,N_29620,N_29932);
nand UO_2608 (O_2608,N_29894,N_29901);
and UO_2609 (O_2609,N_29859,N_29980);
nor UO_2610 (O_2610,N_29807,N_29594);
and UO_2611 (O_2611,N_29923,N_29955);
and UO_2612 (O_2612,N_29968,N_29500);
and UO_2613 (O_2613,N_29618,N_29895);
nand UO_2614 (O_2614,N_29531,N_29617);
and UO_2615 (O_2615,N_29648,N_29568);
or UO_2616 (O_2616,N_29811,N_29836);
or UO_2617 (O_2617,N_29987,N_29601);
or UO_2618 (O_2618,N_29586,N_29823);
xor UO_2619 (O_2619,N_29628,N_29878);
or UO_2620 (O_2620,N_29559,N_29795);
nor UO_2621 (O_2621,N_29809,N_29818);
or UO_2622 (O_2622,N_29900,N_29645);
or UO_2623 (O_2623,N_29735,N_29575);
and UO_2624 (O_2624,N_29661,N_29730);
xnor UO_2625 (O_2625,N_29746,N_29841);
nor UO_2626 (O_2626,N_29543,N_29868);
xnor UO_2627 (O_2627,N_29801,N_29743);
nand UO_2628 (O_2628,N_29651,N_29973);
or UO_2629 (O_2629,N_29829,N_29708);
xor UO_2630 (O_2630,N_29713,N_29539);
or UO_2631 (O_2631,N_29708,N_29819);
and UO_2632 (O_2632,N_29687,N_29722);
and UO_2633 (O_2633,N_29994,N_29789);
nand UO_2634 (O_2634,N_29523,N_29944);
or UO_2635 (O_2635,N_29795,N_29612);
xnor UO_2636 (O_2636,N_29842,N_29753);
and UO_2637 (O_2637,N_29748,N_29574);
or UO_2638 (O_2638,N_29640,N_29754);
xnor UO_2639 (O_2639,N_29523,N_29860);
or UO_2640 (O_2640,N_29544,N_29583);
and UO_2641 (O_2641,N_29736,N_29563);
nor UO_2642 (O_2642,N_29604,N_29606);
nand UO_2643 (O_2643,N_29919,N_29755);
or UO_2644 (O_2644,N_29554,N_29990);
nand UO_2645 (O_2645,N_29595,N_29905);
and UO_2646 (O_2646,N_29897,N_29783);
xor UO_2647 (O_2647,N_29972,N_29896);
or UO_2648 (O_2648,N_29928,N_29647);
nor UO_2649 (O_2649,N_29597,N_29794);
nor UO_2650 (O_2650,N_29689,N_29516);
nor UO_2651 (O_2651,N_29672,N_29861);
nor UO_2652 (O_2652,N_29805,N_29641);
and UO_2653 (O_2653,N_29582,N_29523);
nor UO_2654 (O_2654,N_29902,N_29777);
nor UO_2655 (O_2655,N_29957,N_29535);
or UO_2656 (O_2656,N_29623,N_29912);
xnor UO_2657 (O_2657,N_29622,N_29915);
nor UO_2658 (O_2658,N_29854,N_29892);
nor UO_2659 (O_2659,N_29933,N_29992);
xor UO_2660 (O_2660,N_29536,N_29544);
xnor UO_2661 (O_2661,N_29938,N_29939);
nand UO_2662 (O_2662,N_29634,N_29923);
xor UO_2663 (O_2663,N_29670,N_29976);
and UO_2664 (O_2664,N_29965,N_29685);
xor UO_2665 (O_2665,N_29935,N_29525);
and UO_2666 (O_2666,N_29724,N_29957);
or UO_2667 (O_2667,N_29854,N_29654);
and UO_2668 (O_2668,N_29870,N_29634);
xor UO_2669 (O_2669,N_29511,N_29962);
or UO_2670 (O_2670,N_29833,N_29898);
and UO_2671 (O_2671,N_29921,N_29860);
nor UO_2672 (O_2672,N_29958,N_29970);
and UO_2673 (O_2673,N_29986,N_29780);
nor UO_2674 (O_2674,N_29712,N_29867);
and UO_2675 (O_2675,N_29784,N_29561);
nor UO_2676 (O_2676,N_29571,N_29929);
xnor UO_2677 (O_2677,N_29793,N_29578);
and UO_2678 (O_2678,N_29558,N_29663);
or UO_2679 (O_2679,N_29561,N_29718);
or UO_2680 (O_2680,N_29787,N_29629);
nor UO_2681 (O_2681,N_29865,N_29745);
nor UO_2682 (O_2682,N_29723,N_29741);
or UO_2683 (O_2683,N_29514,N_29997);
nor UO_2684 (O_2684,N_29587,N_29708);
xnor UO_2685 (O_2685,N_29918,N_29854);
and UO_2686 (O_2686,N_29876,N_29813);
nor UO_2687 (O_2687,N_29717,N_29667);
and UO_2688 (O_2688,N_29652,N_29724);
and UO_2689 (O_2689,N_29806,N_29901);
nand UO_2690 (O_2690,N_29898,N_29659);
nor UO_2691 (O_2691,N_29986,N_29906);
xnor UO_2692 (O_2692,N_29654,N_29783);
and UO_2693 (O_2693,N_29775,N_29739);
or UO_2694 (O_2694,N_29589,N_29646);
nand UO_2695 (O_2695,N_29880,N_29969);
nor UO_2696 (O_2696,N_29848,N_29638);
nor UO_2697 (O_2697,N_29858,N_29919);
or UO_2698 (O_2698,N_29907,N_29680);
xor UO_2699 (O_2699,N_29830,N_29834);
and UO_2700 (O_2700,N_29785,N_29995);
xnor UO_2701 (O_2701,N_29766,N_29582);
or UO_2702 (O_2702,N_29981,N_29926);
xor UO_2703 (O_2703,N_29585,N_29519);
nor UO_2704 (O_2704,N_29883,N_29871);
or UO_2705 (O_2705,N_29522,N_29717);
nor UO_2706 (O_2706,N_29937,N_29732);
xor UO_2707 (O_2707,N_29978,N_29930);
nand UO_2708 (O_2708,N_29708,N_29831);
xnor UO_2709 (O_2709,N_29893,N_29703);
nand UO_2710 (O_2710,N_29623,N_29986);
or UO_2711 (O_2711,N_29750,N_29529);
xnor UO_2712 (O_2712,N_29960,N_29701);
nor UO_2713 (O_2713,N_29609,N_29641);
and UO_2714 (O_2714,N_29564,N_29542);
nor UO_2715 (O_2715,N_29634,N_29806);
nor UO_2716 (O_2716,N_29909,N_29987);
xnor UO_2717 (O_2717,N_29769,N_29622);
and UO_2718 (O_2718,N_29850,N_29833);
or UO_2719 (O_2719,N_29616,N_29746);
or UO_2720 (O_2720,N_29885,N_29533);
and UO_2721 (O_2721,N_29503,N_29762);
nand UO_2722 (O_2722,N_29681,N_29869);
nand UO_2723 (O_2723,N_29682,N_29538);
xor UO_2724 (O_2724,N_29661,N_29738);
xor UO_2725 (O_2725,N_29556,N_29726);
and UO_2726 (O_2726,N_29572,N_29960);
nor UO_2727 (O_2727,N_29985,N_29792);
nor UO_2728 (O_2728,N_29776,N_29803);
xnor UO_2729 (O_2729,N_29982,N_29968);
nor UO_2730 (O_2730,N_29853,N_29924);
xnor UO_2731 (O_2731,N_29759,N_29758);
and UO_2732 (O_2732,N_29519,N_29922);
nand UO_2733 (O_2733,N_29833,N_29687);
nand UO_2734 (O_2734,N_29991,N_29554);
nor UO_2735 (O_2735,N_29692,N_29658);
and UO_2736 (O_2736,N_29805,N_29906);
nand UO_2737 (O_2737,N_29571,N_29990);
or UO_2738 (O_2738,N_29759,N_29548);
nand UO_2739 (O_2739,N_29505,N_29846);
nor UO_2740 (O_2740,N_29992,N_29764);
and UO_2741 (O_2741,N_29675,N_29824);
and UO_2742 (O_2742,N_29523,N_29751);
and UO_2743 (O_2743,N_29593,N_29584);
nand UO_2744 (O_2744,N_29733,N_29992);
nor UO_2745 (O_2745,N_29802,N_29501);
xor UO_2746 (O_2746,N_29763,N_29780);
and UO_2747 (O_2747,N_29675,N_29939);
nor UO_2748 (O_2748,N_29954,N_29721);
and UO_2749 (O_2749,N_29672,N_29603);
nand UO_2750 (O_2750,N_29882,N_29524);
nand UO_2751 (O_2751,N_29852,N_29595);
nor UO_2752 (O_2752,N_29690,N_29668);
or UO_2753 (O_2753,N_29833,N_29776);
nand UO_2754 (O_2754,N_29586,N_29696);
xor UO_2755 (O_2755,N_29502,N_29811);
nand UO_2756 (O_2756,N_29705,N_29936);
or UO_2757 (O_2757,N_29740,N_29948);
or UO_2758 (O_2758,N_29852,N_29516);
nand UO_2759 (O_2759,N_29517,N_29574);
and UO_2760 (O_2760,N_29545,N_29868);
or UO_2761 (O_2761,N_29823,N_29591);
nand UO_2762 (O_2762,N_29792,N_29775);
or UO_2763 (O_2763,N_29777,N_29530);
nor UO_2764 (O_2764,N_29659,N_29846);
nor UO_2765 (O_2765,N_29847,N_29765);
nand UO_2766 (O_2766,N_29571,N_29996);
xor UO_2767 (O_2767,N_29916,N_29877);
nor UO_2768 (O_2768,N_29835,N_29655);
nor UO_2769 (O_2769,N_29543,N_29912);
nand UO_2770 (O_2770,N_29552,N_29757);
or UO_2771 (O_2771,N_29621,N_29991);
xor UO_2772 (O_2772,N_29841,N_29993);
nand UO_2773 (O_2773,N_29792,N_29933);
and UO_2774 (O_2774,N_29685,N_29587);
and UO_2775 (O_2775,N_29930,N_29751);
or UO_2776 (O_2776,N_29602,N_29750);
nor UO_2777 (O_2777,N_29679,N_29935);
xor UO_2778 (O_2778,N_29786,N_29862);
xnor UO_2779 (O_2779,N_29728,N_29885);
or UO_2780 (O_2780,N_29971,N_29833);
or UO_2781 (O_2781,N_29852,N_29696);
and UO_2782 (O_2782,N_29652,N_29988);
nand UO_2783 (O_2783,N_29667,N_29519);
nand UO_2784 (O_2784,N_29508,N_29913);
or UO_2785 (O_2785,N_29693,N_29829);
or UO_2786 (O_2786,N_29633,N_29588);
nor UO_2787 (O_2787,N_29802,N_29751);
nand UO_2788 (O_2788,N_29798,N_29969);
and UO_2789 (O_2789,N_29988,N_29808);
or UO_2790 (O_2790,N_29718,N_29523);
and UO_2791 (O_2791,N_29621,N_29997);
xor UO_2792 (O_2792,N_29547,N_29733);
and UO_2793 (O_2793,N_29864,N_29565);
nor UO_2794 (O_2794,N_29791,N_29796);
and UO_2795 (O_2795,N_29565,N_29819);
nand UO_2796 (O_2796,N_29824,N_29999);
and UO_2797 (O_2797,N_29821,N_29651);
xnor UO_2798 (O_2798,N_29948,N_29636);
and UO_2799 (O_2799,N_29846,N_29843);
nor UO_2800 (O_2800,N_29793,N_29811);
nor UO_2801 (O_2801,N_29788,N_29719);
nor UO_2802 (O_2802,N_29571,N_29799);
and UO_2803 (O_2803,N_29859,N_29689);
or UO_2804 (O_2804,N_29670,N_29649);
and UO_2805 (O_2805,N_29726,N_29544);
nand UO_2806 (O_2806,N_29973,N_29632);
nand UO_2807 (O_2807,N_29898,N_29681);
nor UO_2808 (O_2808,N_29721,N_29698);
nor UO_2809 (O_2809,N_29833,N_29591);
nand UO_2810 (O_2810,N_29761,N_29803);
nor UO_2811 (O_2811,N_29553,N_29970);
nor UO_2812 (O_2812,N_29727,N_29821);
nand UO_2813 (O_2813,N_29751,N_29693);
and UO_2814 (O_2814,N_29597,N_29674);
xor UO_2815 (O_2815,N_29733,N_29686);
xnor UO_2816 (O_2816,N_29719,N_29995);
nand UO_2817 (O_2817,N_29681,N_29580);
nor UO_2818 (O_2818,N_29983,N_29733);
or UO_2819 (O_2819,N_29808,N_29627);
and UO_2820 (O_2820,N_29681,N_29583);
and UO_2821 (O_2821,N_29673,N_29600);
and UO_2822 (O_2822,N_29879,N_29567);
xnor UO_2823 (O_2823,N_29852,N_29980);
or UO_2824 (O_2824,N_29558,N_29818);
and UO_2825 (O_2825,N_29936,N_29944);
xor UO_2826 (O_2826,N_29633,N_29831);
or UO_2827 (O_2827,N_29768,N_29511);
nor UO_2828 (O_2828,N_29716,N_29696);
nand UO_2829 (O_2829,N_29920,N_29883);
xnor UO_2830 (O_2830,N_29918,N_29582);
xor UO_2831 (O_2831,N_29635,N_29550);
or UO_2832 (O_2832,N_29521,N_29965);
nand UO_2833 (O_2833,N_29501,N_29629);
or UO_2834 (O_2834,N_29669,N_29627);
nand UO_2835 (O_2835,N_29775,N_29726);
and UO_2836 (O_2836,N_29692,N_29996);
nand UO_2837 (O_2837,N_29852,N_29795);
xor UO_2838 (O_2838,N_29872,N_29907);
xnor UO_2839 (O_2839,N_29613,N_29653);
and UO_2840 (O_2840,N_29812,N_29966);
or UO_2841 (O_2841,N_29617,N_29569);
nand UO_2842 (O_2842,N_29533,N_29769);
nor UO_2843 (O_2843,N_29543,N_29809);
nor UO_2844 (O_2844,N_29874,N_29939);
xor UO_2845 (O_2845,N_29751,N_29940);
and UO_2846 (O_2846,N_29678,N_29542);
and UO_2847 (O_2847,N_29546,N_29587);
and UO_2848 (O_2848,N_29914,N_29588);
nor UO_2849 (O_2849,N_29593,N_29550);
xor UO_2850 (O_2850,N_29638,N_29932);
and UO_2851 (O_2851,N_29987,N_29848);
nor UO_2852 (O_2852,N_29745,N_29795);
and UO_2853 (O_2853,N_29651,N_29853);
and UO_2854 (O_2854,N_29534,N_29985);
or UO_2855 (O_2855,N_29624,N_29615);
and UO_2856 (O_2856,N_29778,N_29546);
or UO_2857 (O_2857,N_29967,N_29902);
nor UO_2858 (O_2858,N_29886,N_29687);
nor UO_2859 (O_2859,N_29622,N_29763);
nor UO_2860 (O_2860,N_29625,N_29859);
xor UO_2861 (O_2861,N_29894,N_29647);
xor UO_2862 (O_2862,N_29579,N_29585);
nor UO_2863 (O_2863,N_29717,N_29858);
or UO_2864 (O_2864,N_29902,N_29714);
nand UO_2865 (O_2865,N_29562,N_29920);
and UO_2866 (O_2866,N_29657,N_29618);
or UO_2867 (O_2867,N_29531,N_29663);
xnor UO_2868 (O_2868,N_29949,N_29790);
nand UO_2869 (O_2869,N_29821,N_29633);
nor UO_2870 (O_2870,N_29668,N_29623);
nand UO_2871 (O_2871,N_29718,N_29654);
nor UO_2872 (O_2872,N_29962,N_29601);
xor UO_2873 (O_2873,N_29864,N_29842);
nand UO_2874 (O_2874,N_29977,N_29745);
and UO_2875 (O_2875,N_29531,N_29536);
and UO_2876 (O_2876,N_29833,N_29565);
nand UO_2877 (O_2877,N_29923,N_29970);
nand UO_2878 (O_2878,N_29949,N_29501);
and UO_2879 (O_2879,N_29714,N_29767);
xor UO_2880 (O_2880,N_29943,N_29565);
or UO_2881 (O_2881,N_29798,N_29708);
and UO_2882 (O_2882,N_29502,N_29662);
or UO_2883 (O_2883,N_29649,N_29602);
nand UO_2884 (O_2884,N_29902,N_29539);
or UO_2885 (O_2885,N_29897,N_29837);
or UO_2886 (O_2886,N_29650,N_29514);
nand UO_2887 (O_2887,N_29874,N_29549);
xor UO_2888 (O_2888,N_29567,N_29964);
and UO_2889 (O_2889,N_29775,N_29784);
xor UO_2890 (O_2890,N_29881,N_29770);
xor UO_2891 (O_2891,N_29687,N_29653);
nand UO_2892 (O_2892,N_29782,N_29919);
nor UO_2893 (O_2893,N_29542,N_29871);
nand UO_2894 (O_2894,N_29892,N_29795);
xnor UO_2895 (O_2895,N_29849,N_29559);
nand UO_2896 (O_2896,N_29576,N_29636);
nor UO_2897 (O_2897,N_29661,N_29599);
nor UO_2898 (O_2898,N_29838,N_29545);
xnor UO_2899 (O_2899,N_29668,N_29711);
nand UO_2900 (O_2900,N_29932,N_29757);
nor UO_2901 (O_2901,N_29890,N_29969);
and UO_2902 (O_2902,N_29744,N_29795);
and UO_2903 (O_2903,N_29574,N_29698);
or UO_2904 (O_2904,N_29592,N_29935);
nand UO_2905 (O_2905,N_29693,N_29804);
xor UO_2906 (O_2906,N_29757,N_29985);
and UO_2907 (O_2907,N_29663,N_29930);
and UO_2908 (O_2908,N_29616,N_29769);
nand UO_2909 (O_2909,N_29569,N_29861);
and UO_2910 (O_2910,N_29548,N_29629);
and UO_2911 (O_2911,N_29626,N_29942);
nor UO_2912 (O_2912,N_29687,N_29977);
nand UO_2913 (O_2913,N_29654,N_29951);
nand UO_2914 (O_2914,N_29671,N_29942);
nand UO_2915 (O_2915,N_29970,N_29819);
xnor UO_2916 (O_2916,N_29646,N_29957);
or UO_2917 (O_2917,N_29544,N_29730);
or UO_2918 (O_2918,N_29873,N_29790);
and UO_2919 (O_2919,N_29530,N_29658);
or UO_2920 (O_2920,N_29529,N_29862);
nor UO_2921 (O_2921,N_29915,N_29800);
or UO_2922 (O_2922,N_29926,N_29979);
nor UO_2923 (O_2923,N_29804,N_29549);
nand UO_2924 (O_2924,N_29758,N_29518);
xnor UO_2925 (O_2925,N_29924,N_29814);
nand UO_2926 (O_2926,N_29946,N_29522);
xor UO_2927 (O_2927,N_29853,N_29985);
or UO_2928 (O_2928,N_29868,N_29909);
nor UO_2929 (O_2929,N_29948,N_29907);
and UO_2930 (O_2930,N_29751,N_29790);
nand UO_2931 (O_2931,N_29583,N_29769);
nor UO_2932 (O_2932,N_29571,N_29639);
xor UO_2933 (O_2933,N_29802,N_29916);
or UO_2934 (O_2934,N_29920,N_29828);
nor UO_2935 (O_2935,N_29652,N_29746);
and UO_2936 (O_2936,N_29740,N_29668);
nand UO_2937 (O_2937,N_29558,N_29607);
nand UO_2938 (O_2938,N_29541,N_29819);
xor UO_2939 (O_2939,N_29907,N_29526);
nand UO_2940 (O_2940,N_29526,N_29720);
and UO_2941 (O_2941,N_29567,N_29619);
nor UO_2942 (O_2942,N_29564,N_29757);
and UO_2943 (O_2943,N_29594,N_29706);
and UO_2944 (O_2944,N_29816,N_29581);
nand UO_2945 (O_2945,N_29804,N_29756);
xnor UO_2946 (O_2946,N_29607,N_29925);
nor UO_2947 (O_2947,N_29669,N_29650);
nor UO_2948 (O_2948,N_29733,N_29993);
nand UO_2949 (O_2949,N_29587,N_29597);
and UO_2950 (O_2950,N_29902,N_29758);
or UO_2951 (O_2951,N_29851,N_29636);
and UO_2952 (O_2952,N_29912,N_29506);
nand UO_2953 (O_2953,N_29772,N_29973);
and UO_2954 (O_2954,N_29549,N_29653);
nand UO_2955 (O_2955,N_29624,N_29603);
nand UO_2956 (O_2956,N_29853,N_29997);
and UO_2957 (O_2957,N_29616,N_29570);
nand UO_2958 (O_2958,N_29563,N_29813);
xnor UO_2959 (O_2959,N_29860,N_29962);
or UO_2960 (O_2960,N_29642,N_29801);
nor UO_2961 (O_2961,N_29511,N_29799);
or UO_2962 (O_2962,N_29580,N_29511);
nor UO_2963 (O_2963,N_29609,N_29784);
nand UO_2964 (O_2964,N_29698,N_29958);
or UO_2965 (O_2965,N_29838,N_29923);
xnor UO_2966 (O_2966,N_29789,N_29900);
xnor UO_2967 (O_2967,N_29863,N_29663);
nor UO_2968 (O_2968,N_29833,N_29787);
nor UO_2969 (O_2969,N_29508,N_29919);
and UO_2970 (O_2970,N_29758,N_29822);
xnor UO_2971 (O_2971,N_29996,N_29687);
or UO_2972 (O_2972,N_29905,N_29899);
nand UO_2973 (O_2973,N_29924,N_29506);
nand UO_2974 (O_2974,N_29696,N_29634);
nor UO_2975 (O_2975,N_29926,N_29661);
nor UO_2976 (O_2976,N_29569,N_29738);
nand UO_2977 (O_2977,N_29779,N_29993);
nand UO_2978 (O_2978,N_29931,N_29759);
nor UO_2979 (O_2979,N_29691,N_29739);
nor UO_2980 (O_2980,N_29517,N_29551);
or UO_2981 (O_2981,N_29658,N_29708);
or UO_2982 (O_2982,N_29650,N_29548);
or UO_2983 (O_2983,N_29545,N_29631);
nor UO_2984 (O_2984,N_29639,N_29914);
xor UO_2985 (O_2985,N_29515,N_29540);
nand UO_2986 (O_2986,N_29573,N_29523);
and UO_2987 (O_2987,N_29663,N_29656);
and UO_2988 (O_2988,N_29537,N_29752);
nor UO_2989 (O_2989,N_29947,N_29883);
nor UO_2990 (O_2990,N_29677,N_29854);
and UO_2991 (O_2991,N_29589,N_29610);
nand UO_2992 (O_2992,N_29861,N_29661);
or UO_2993 (O_2993,N_29539,N_29710);
nor UO_2994 (O_2994,N_29539,N_29795);
xnor UO_2995 (O_2995,N_29954,N_29720);
nand UO_2996 (O_2996,N_29675,N_29805);
nor UO_2997 (O_2997,N_29533,N_29535);
nand UO_2998 (O_2998,N_29777,N_29560);
xor UO_2999 (O_2999,N_29642,N_29599);
and UO_3000 (O_3000,N_29594,N_29686);
xor UO_3001 (O_3001,N_29844,N_29747);
and UO_3002 (O_3002,N_29939,N_29703);
nor UO_3003 (O_3003,N_29587,N_29519);
or UO_3004 (O_3004,N_29743,N_29773);
or UO_3005 (O_3005,N_29946,N_29597);
and UO_3006 (O_3006,N_29656,N_29564);
nor UO_3007 (O_3007,N_29860,N_29820);
and UO_3008 (O_3008,N_29968,N_29552);
nor UO_3009 (O_3009,N_29623,N_29624);
xor UO_3010 (O_3010,N_29581,N_29653);
nor UO_3011 (O_3011,N_29563,N_29823);
xnor UO_3012 (O_3012,N_29861,N_29629);
xnor UO_3013 (O_3013,N_29634,N_29711);
nand UO_3014 (O_3014,N_29740,N_29816);
or UO_3015 (O_3015,N_29684,N_29681);
nand UO_3016 (O_3016,N_29799,N_29563);
nand UO_3017 (O_3017,N_29979,N_29982);
and UO_3018 (O_3018,N_29604,N_29572);
or UO_3019 (O_3019,N_29962,N_29692);
xor UO_3020 (O_3020,N_29706,N_29518);
nor UO_3021 (O_3021,N_29973,N_29971);
nand UO_3022 (O_3022,N_29891,N_29878);
and UO_3023 (O_3023,N_29816,N_29507);
nor UO_3024 (O_3024,N_29854,N_29753);
nand UO_3025 (O_3025,N_29617,N_29525);
or UO_3026 (O_3026,N_29944,N_29686);
and UO_3027 (O_3027,N_29818,N_29804);
xor UO_3028 (O_3028,N_29507,N_29938);
xor UO_3029 (O_3029,N_29596,N_29898);
nand UO_3030 (O_3030,N_29992,N_29500);
xnor UO_3031 (O_3031,N_29994,N_29827);
xnor UO_3032 (O_3032,N_29792,N_29839);
nor UO_3033 (O_3033,N_29995,N_29755);
nand UO_3034 (O_3034,N_29892,N_29863);
xor UO_3035 (O_3035,N_29540,N_29774);
nand UO_3036 (O_3036,N_29840,N_29711);
nor UO_3037 (O_3037,N_29634,N_29703);
xnor UO_3038 (O_3038,N_29915,N_29913);
nor UO_3039 (O_3039,N_29990,N_29941);
xnor UO_3040 (O_3040,N_29622,N_29992);
xor UO_3041 (O_3041,N_29775,N_29777);
and UO_3042 (O_3042,N_29860,N_29534);
nor UO_3043 (O_3043,N_29599,N_29756);
or UO_3044 (O_3044,N_29729,N_29740);
xnor UO_3045 (O_3045,N_29671,N_29766);
xor UO_3046 (O_3046,N_29541,N_29603);
xor UO_3047 (O_3047,N_29937,N_29682);
nor UO_3048 (O_3048,N_29738,N_29529);
xnor UO_3049 (O_3049,N_29731,N_29956);
or UO_3050 (O_3050,N_29990,N_29758);
and UO_3051 (O_3051,N_29537,N_29914);
or UO_3052 (O_3052,N_29917,N_29596);
and UO_3053 (O_3053,N_29552,N_29876);
nand UO_3054 (O_3054,N_29903,N_29850);
and UO_3055 (O_3055,N_29514,N_29535);
or UO_3056 (O_3056,N_29825,N_29816);
xnor UO_3057 (O_3057,N_29731,N_29957);
or UO_3058 (O_3058,N_29848,N_29591);
or UO_3059 (O_3059,N_29745,N_29851);
or UO_3060 (O_3060,N_29616,N_29786);
xnor UO_3061 (O_3061,N_29781,N_29791);
nand UO_3062 (O_3062,N_29882,N_29608);
nand UO_3063 (O_3063,N_29596,N_29626);
and UO_3064 (O_3064,N_29834,N_29671);
or UO_3065 (O_3065,N_29753,N_29870);
or UO_3066 (O_3066,N_29936,N_29651);
nand UO_3067 (O_3067,N_29985,N_29631);
nand UO_3068 (O_3068,N_29669,N_29933);
or UO_3069 (O_3069,N_29926,N_29744);
nor UO_3070 (O_3070,N_29720,N_29868);
and UO_3071 (O_3071,N_29906,N_29706);
or UO_3072 (O_3072,N_29594,N_29592);
nor UO_3073 (O_3073,N_29579,N_29732);
or UO_3074 (O_3074,N_29924,N_29732);
xnor UO_3075 (O_3075,N_29895,N_29546);
xor UO_3076 (O_3076,N_29882,N_29945);
and UO_3077 (O_3077,N_29839,N_29599);
nor UO_3078 (O_3078,N_29676,N_29544);
nand UO_3079 (O_3079,N_29971,N_29997);
or UO_3080 (O_3080,N_29987,N_29800);
and UO_3081 (O_3081,N_29613,N_29985);
and UO_3082 (O_3082,N_29854,N_29600);
nand UO_3083 (O_3083,N_29754,N_29750);
nor UO_3084 (O_3084,N_29826,N_29953);
and UO_3085 (O_3085,N_29956,N_29932);
or UO_3086 (O_3086,N_29884,N_29540);
or UO_3087 (O_3087,N_29544,N_29650);
nand UO_3088 (O_3088,N_29908,N_29961);
xor UO_3089 (O_3089,N_29864,N_29717);
or UO_3090 (O_3090,N_29901,N_29572);
nand UO_3091 (O_3091,N_29833,N_29516);
and UO_3092 (O_3092,N_29753,N_29902);
and UO_3093 (O_3093,N_29525,N_29805);
and UO_3094 (O_3094,N_29563,N_29718);
or UO_3095 (O_3095,N_29749,N_29558);
nand UO_3096 (O_3096,N_29926,N_29907);
or UO_3097 (O_3097,N_29730,N_29913);
or UO_3098 (O_3098,N_29546,N_29605);
xor UO_3099 (O_3099,N_29534,N_29708);
nor UO_3100 (O_3100,N_29845,N_29696);
xnor UO_3101 (O_3101,N_29830,N_29566);
nand UO_3102 (O_3102,N_29725,N_29692);
nand UO_3103 (O_3103,N_29849,N_29689);
and UO_3104 (O_3104,N_29963,N_29636);
or UO_3105 (O_3105,N_29508,N_29943);
nor UO_3106 (O_3106,N_29613,N_29623);
and UO_3107 (O_3107,N_29905,N_29836);
nand UO_3108 (O_3108,N_29715,N_29937);
and UO_3109 (O_3109,N_29686,N_29653);
and UO_3110 (O_3110,N_29798,N_29898);
and UO_3111 (O_3111,N_29945,N_29516);
and UO_3112 (O_3112,N_29635,N_29586);
nor UO_3113 (O_3113,N_29633,N_29867);
and UO_3114 (O_3114,N_29600,N_29876);
and UO_3115 (O_3115,N_29608,N_29818);
nor UO_3116 (O_3116,N_29559,N_29667);
or UO_3117 (O_3117,N_29763,N_29593);
nand UO_3118 (O_3118,N_29545,N_29550);
nor UO_3119 (O_3119,N_29980,N_29653);
or UO_3120 (O_3120,N_29966,N_29975);
nand UO_3121 (O_3121,N_29798,N_29719);
and UO_3122 (O_3122,N_29747,N_29555);
nor UO_3123 (O_3123,N_29612,N_29708);
and UO_3124 (O_3124,N_29623,N_29741);
and UO_3125 (O_3125,N_29860,N_29696);
nand UO_3126 (O_3126,N_29609,N_29857);
xnor UO_3127 (O_3127,N_29669,N_29972);
or UO_3128 (O_3128,N_29545,N_29575);
or UO_3129 (O_3129,N_29710,N_29873);
or UO_3130 (O_3130,N_29842,N_29635);
xor UO_3131 (O_3131,N_29794,N_29622);
xor UO_3132 (O_3132,N_29856,N_29552);
and UO_3133 (O_3133,N_29702,N_29902);
or UO_3134 (O_3134,N_29885,N_29625);
nor UO_3135 (O_3135,N_29828,N_29918);
nor UO_3136 (O_3136,N_29565,N_29998);
nand UO_3137 (O_3137,N_29566,N_29962);
nor UO_3138 (O_3138,N_29577,N_29849);
and UO_3139 (O_3139,N_29919,N_29866);
or UO_3140 (O_3140,N_29885,N_29744);
xor UO_3141 (O_3141,N_29912,N_29535);
nand UO_3142 (O_3142,N_29569,N_29743);
or UO_3143 (O_3143,N_29560,N_29789);
and UO_3144 (O_3144,N_29755,N_29829);
nor UO_3145 (O_3145,N_29873,N_29814);
nor UO_3146 (O_3146,N_29894,N_29838);
or UO_3147 (O_3147,N_29599,N_29916);
nor UO_3148 (O_3148,N_29664,N_29784);
nand UO_3149 (O_3149,N_29791,N_29632);
nand UO_3150 (O_3150,N_29813,N_29712);
or UO_3151 (O_3151,N_29914,N_29770);
nand UO_3152 (O_3152,N_29920,N_29930);
nand UO_3153 (O_3153,N_29511,N_29599);
xor UO_3154 (O_3154,N_29767,N_29575);
xor UO_3155 (O_3155,N_29987,N_29681);
nor UO_3156 (O_3156,N_29564,N_29974);
or UO_3157 (O_3157,N_29506,N_29943);
nand UO_3158 (O_3158,N_29999,N_29998);
xnor UO_3159 (O_3159,N_29785,N_29901);
or UO_3160 (O_3160,N_29735,N_29809);
xnor UO_3161 (O_3161,N_29558,N_29526);
nor UO_3162 (O_3162,N_29575,N_29555);
or UO_3163 (O_3163,N_29598,N_29941);
and UO_3164 (O_3164,N_29870,N_29983);
nand UO_3165 (O_3165,N_29967,N_29791);
and UO_3166 (O_3166,N_29855,N_29754);
xnor UO_3167 (O_3167,N_29654,N_29717);
or UO_3168 (O_3168,N_29688,N_29683);
nor UO_3169 (O_3169,N_29587,N_29729);
and UO_3170 (O_3170,N_29958,N_29567);
and UO_3171 (O_3171,N_29587,N_29591);
and UO_3172 (O_3172,N_29913,N_29511);
and UO_3173 (O_3173,N_29922,N_29900);
nand UO_3174 (O_3174,N_29505,N_29730);
or UO_3175 (O_3175,N_29551,N_29554);
or UO_3176 (O_3176,N_29580,N_29783);
xor UO_3177 (O_3177,N_29699,N_29720);
or UO_3178 (O_3178,N_29825,N_29517);
nor UO_3179 (O_3179,N_29960,N_29748);
nor UO_3180 (O_3180,N_29827,N_29696);
or UO_3181 (O_3181,N_29770,N_29928);
xnor UO_3182 (O_3182,N_29734,N_29543);
xor UO_3183 (O_3183,N_29731,N_29784);
nand UO_3184 (O_3184,N_29758,N_29586);
or UO_3185 (O_3185,N_29540,N_29804);
nand UO_3186 (O_3186,N_29971,N_29667);
and UO_3187 (O_3187,N_29613,N_29906);
or UO_3188 (O_3188,N_29801,N_29520);
nand UO_3189 (O_3189,N_29744,N_29957);
and UO_3190 (O_3190,N_29846,N_29589);
nand UO_3191 (O_3191,N_29892,N_29719);
and UO_3192 (O_3192,N_29946,N_29851);
nor UO_3193 (O_3193,N_29575,N_29745);
nand UO_3194 (O_3194,N_29953,N_29565);
or UO_3195 (O_3195,N_29598,N_29622);
nor UO_3196 (O_3196,N_29881,N_29804);
and UO_3197 (O_3197,N_29820,N_29813);
or UO_3198 (O_3198,N_29684,N_29660);
xor UO_3199 (O_3199,N_29961,N_29585);
xnor UO_3200 (O_3200,N_29903,N_29997);
nor UO_3201 (O_3201,N_29967,N_29538);
or UO_3202 (O_3202,N_29864,N_29582);
nor UO_3203 (O_3203,N_29843,N_29856);
xor UO_3204 (O_3204,N_29650,N_29794);
and UO_3205 (O_3205,N_29759,N_29783);
xnor UO_3206 (O_3206,N_29647,N_29590);
or UO_3207 (O_3207,N_29957,N_29516);
xnor UO_3208 (O_3208,N_29633,N_29804);
and UO_3209 (O_3209,N_29797,N_29845);
or UO_3210 (O_3210,N_29636,N_29611);
and UO_3211 (O_3211,N_29836,N_29861);
and UO_3212 (O_3212,N_29952,N_29674);
nor UO_3213 (O_3213,N_29836,N_29879);
nor UO_3214 (O_3214,N_29690,N_29807);
nand UO_3215 (O_3215,N_29859,N_29782);
nand UO_3216 (O_3216,N_29771,N_29662);
or UO_3217 (O_3217,N_29846,N_29632);
nor UO_3218 (O_3218,N_29792,N_29735);
or UO_3219 (O_3219,N_29805,N_29809);
or UO_3220 (O_3220,N_29944,N_29576);
and UO_3221 (O_3221,N_29728,N_29545);
and UO_3222 (O_3222,N_29966,N_29692);
nor UO_3223 (O_3223,N_29988,N_29720);
nand UO_3224 (O_3224,N_29742,N_29596);
nand UO_3225 (O_3225,N_29640,N_29652);
nand UO_3226 (O_3226,N_29629,N_29648);
or UO_3227 (O_3227,N_29783,N_29903);
and UO_3228 (O_3228,N_29700,N_29671);
nor UO_3229 (O_3229,N_29786,N_29755);
nor UO_3230 (O_3230,N_29742,N_29985);
nor UO_3231 (O_3231,N_29616,N_29751);
xor UO_3232 (O_3232,N_29592,N_29749);
and UO_3233 (O_3233,N_29580,N_29915);
xnor UO_3234 (O_3234,N_29618,N_29788);
xnor UO_3235 (O_3235,N_29840,N_29884);
nor UO_3236 (O_3236,N_29725,N_29891);
nor UO_3237 (O_3237,N_29938,N_29533);
and UO_3238 (O_3238,N_29936,N_29744);
xnor UO_3239 (O_3239,N_29838,N_29527);
nand UO_3240 (O_3240,N_29728,N_29704);
and UO_3241 (O_3241,N_29932,N_29944);
and UO_3242 (O_3242,N_29634,N_29907);
or UO_3243 (O_3243,N_29766,N_29998);
nand UO_3244 (O_3244,N_29683,N_29924);
xor UO_3245 (O_3245,N_29875,N_29596);
nor UO_3246 (O_3246,N_29955,N_29865);
and UO_3247 (O_3247,N_29723,N_29746);
nand UO_3248 (O_3248,N_29999,N_29533);
or UO_3249 (O_3249,N_29752,N_29666);
nand UO_3250 (O_3250,N_29922,N_29647);
nand UO_3251 (O_3251,N_29755,N_29551);
xor UO_3252 (O_3252,N_29865,N_29731);
nor UO_3253 (O_3253,N_29866,N_29515);
or UO_3254 (O_3254,N_29845,N_29765);
or UO_3255 (O_3255,N_29789,N_29885);
and UO_3256 (O_3256,N_29855,N_29940);
xor UO_3257 (O_3257,N_29755,N_29586);
xnor UO_3258 (O_3258,N_29878,N_29663);
or UO_3259 (O_3259,N_29723,N_29800);
and UO_3260 (O_3260,N_29640,N_29505);
nor UO_3261 (O_3261,N_29819,N_29632);
nor UO_3262 (O_3262,N_29847,N_29741);
and UO_3263 (O_3263,N_29592,N_29746);
nor UO_3264 (O_3264,N_29506,N_29743);
nand UO_3265 (O_3265,N_29555,N_29961);
nand UO_3266 (O_3266,N_29638,N_29583);
and UO_3267 (O_3267,N_29832,N_29923);
or UO_3268 (O_3268,N_29605,N_29721);
and UO_3269 (O_3269,N_29961,N_29923);
and UO_3270 (O_3270,N_29927,N_29563);
nand UO_3271 (O_3271,N_29833,N_29601);
nor UO_3272 (O_3272,N_29977,N_29786);
nand UO_3273 (O_3273,N_29983,N_29684);
xnor UO_3274 (O_3274,N_29720,N_29801);
and UO_3275 (O_3275,N_29791,N_29806);
and UO_3276 (O_3276,N_29528,N_29857);
nor UO_3277 (O_3277,N_29991,N_29516);
nor UO_3278 (O_3278,N_29907,N_29677);
xnor UO_3279 (O_3279,N_29636,N_29542);
xnor UO_3280 (O_3280,N_29992,N_29838);
xor UO_3281 (O_3281,N_29573,N_29580);
or UO_3282 (O_3282,N_29791,N_29913);
and UO_3283 (O_3283,N_29633,N_29976);
xor UO_3284 (O_3284,N_29506,N_29697);
xnor UO_3285 (O_3285,N_29682,N_29878);
nor UO_3286 (O_3286,N_29571,N_29842);
nand UO_3287 (O_3287,N_29970,N_29594);
or UO_3288 (O_3288,N_29659,N_29735);
xor UO_3289 (O_3289,N_29548,N_29821);
or UO_3290 (O_3290,N_29923,N_29734);
or UO_3291 (O_3291,N_29714,N_29979);
and UO_3292 (O_3292,N_29515,N_29815);
or UO_3293 (O_3293,N_29504,N_29568);
and UO_3294 (O_3294,N_29983,N_29577);
or UO_3295 (O_3295,N_29911,N_29712);
or UO_3296 (O_3296,N_29613,N_29890);
nor UO_3297 (O_3297,N_29517,N_29556);
and UO_3298 (O_3298,N_29889,N_29500);
xnor UO_3299 (O_3299,N_29738,N_29791);
nor UO_3300 (O_3300,N_29818,N_29935);
and UO_3301 (O_3301,N_29985,N_29827);
and UO_3302 (O_3302,N_29938,N_29790);
nand UO_3303 (O_3303,N_29940,N_29677);
nor UO_3304 (O_3304,N_29537,N_29730);
or UO_3305 (O_3305,N_29943,N_29927);
nor UO_3306 (O_3306,N_29710,N_29622);
nand UO_3307 (O_3307,N_29783,N_29884);
nor UO_3308 (O_3308,N_29871,N_29762);
and UO_3309 (O_3309,N_29737,N_29676);
or UO_3310 (O_3310,N_29579,N_29759);
and UO_3311 (O_3311,N_29788,N_29647);
xnor UO_3312 (O_3312,N_29855,N_29968);
xor UO_3313 (O_3313,N_29519,N_29973);
nor UO_3314 (O_3314,N_29959,N_29772);
and UO_3315 (O_3315,N_29504,N_29567);
xor UO_3316 (O_3316,N_29893,N_29819);
and UO_3317 (O_3317,N_29514,N_29593);
xnor UO_3318 (O_3318,N_29908,N_29660);
xnor UO_3319 (O_3319,N_29611,N_29759);
nand UO_3320 (O_3320,N_29739,N_29689);
nand UO_3321 (O_3321,N_29791,N_29513);
nand UO_3322 (O_3322,N_29554,N_29778);
and UO_3323 (O_3323,N_29516,N_29749);
or UO_3324 (O_3324,N_29508,N_29764);
xor UO_3325 (O_3325,N_29971,N_29895);
xnor UO_3326 (O_3326,N_29866,N_29995);
nor UO_3327 (O_3327,N_29987,N_29824);
nand UO_3328 (O_3328,N_29699,N_29725);
or UO_3329 (O_3329,N_29874,N_29521);
xor UO_3330 (O_3330,N_29534,N_29888);
xnor UO_3331 (O_3331,N_29583,N_29878);
or UO_3332 (O_3332,N_29917,N_29662);
or UO_3333 (O_3333,N_29803,N_29854);
and UO_3334 (O_3334,N_29587,N_29515);
and UO_3335 (O_3335,N_29900,N_29683);
or UO_3336 (O_3336,N_29848,N_29970);
or UO_3337 (O_3337,N_29736,N_29932);
nor UO_3338 (O_3338,N_29979,N_29629);
xnor UO_3339 (O_3339,N_29589,N_29975);
nor UO_3340 (O_3340,N_29520,N_29501);
nand UO_3341 (O_3341,N_29955,N_29647);
nand UO_3342 (O_3342,N_29943,N_29953);
nand UO_3343 (O_3343,N_29623,N_29917);
and UO_3344 (O_3344,N_29716,N_29828);
and UO_3345 (O_3345,N_29704,N_29649);
and UO_3346 (O_3346,N_29516,N_29840);
or UO_3347 (O_3347,N_29798,N_29723);
or UO_3348 (O_3348,N_29966,N_29636);
or UO_3349 (O_3349,N_29964,N_29700);
nand UO_3350 (O_3350,N_29971,N_29802);
nand UO_3351 (O_3351,N_29551,N_29540);
xnor UO_3352 (O_3352,N_29643,N_29947);
xnor UO_3353 (O_3353,N_29748,N_29890);
nor UO_3354 (O_3354,N_29515,N_29913);
and UO_3355 (O_3355,N_29518,N_29615);
and UO_3356 (O_3356,N_29789,N_29916);
xnor UO_3357 (O_3357,N_29968,N_29752);
xor UO_3358 (O_3358,N_29544,N_29906);
nor UO_3359 (O_3359,N_29794,N_29607);
xor UO_3360 (O_3360,N_29818,N_29672);
and UO_3361 (O_3361,N_29741,N_29634);
or UO_3362 (O_3362,N_29989,N_29537);
or UO_3363 (O_3363,N_29613,N_29604);
or UO_3364 (O_3364,N_29731,N_29579);
xor UO_3365 (O_3365,N_29725,N_29828);
nor UO_3366 (O_3366,N_29628,N_29772);
or UO_3367 (O_3367,N_29641,N_29936);
nor UO_3368 (O_3368,N_29868,N_29586);
or UO_3369 (O_3369,N_29554,N_29919);
xor UO_3370 (O_3370,N_29984,N_29598);
and UO_3371 (O_3371,N_29608,N_29678);
and UO_3372 (O_3372,N_29569,N_29729);
xor UO_3373 (O_3373,N_29993,N_29510);
xnor UO_3374 (O_3374,N_29968,N_29563);
nand UO_3375 (O_3375,N_29735,N_29999);
nor UO_3376 (O_3376,N_29752,N_29692);
and UO_3377 (O_3377,N_29984,N_29669);
and UO_3378 (O_3378,N_29637,N_29733);
and UO_3379 (O_3379,N_29784,N_29697);
nor UO_3380 (O_3380,N_29913,N_29993);
nor UO_3381 (O_3381,N_29820,N_29974);
and UO_3382 (O_3382,N_29674,N_29562);
xnor UO_3383 (O_3383,N_29684,N_29704);
and UO_3384 (O_3384,N_29547,N_29599);
nand UO_3385 (O_3385,N_29845,N_29912);
xnor UO_3386 (O_3386,N_29751,N_29534);
nor UO_3387 (O_3387,N_29653,N_29867);
nor UO_3388 (O_3388,N_29500,N_29632);
nand UO_3389 (O_3389,N_29935,N_29883);
or UO_3390 (O_3390,N_29626,N_29793);
and UO_3391 (O_3391,N_29959,N_29522);
or UO_3392 (O_3392,N_29711,N_29565);
xor UO_3393 (O_3393,N_29903,N_29886);
or UO_3394 (O_3394,N_29562,N_29560);
or UO_3395 (O_3395,N_29961,N_29707);
nand UO_3396 (O_3396,N_29582,N_29692);
nand UO_3397 (O_3397,N_29527,N_29859);
nor UO_3398 (O_3398,N_29901,N_29593);
nand UO_3399 (O_3399,N_29599,N_29507);
xor UO_3400 (O_3400,N_29812,N_29512);
nand UO_3401 (O_3401,N_29576,N_29768);
xnor UO_3402 (O_3402,N_29810,N_29678);
nand UO_3403 (O_3403,N_29920,N_29590);
nor UO_3404 (O_3404,N_29733,N_29945);
or UO_3405 (O_3405,N_29725,N_29841);
nand UO_3406 (O_3406,N_29833,N_29854);
xor UO_3407 (O_3407,N_29728,N_29705);
or UO_3408 (O_3408,N_29755,N_29966);
xnor UO_3409 (O_3409,N_29843,N_29580);
and UO_3410 (O_3410,N_29873,N_29795);
or UO_3411 (O_3411,N_29688,N_29537);
nor UO_3412 (O_3412,N_29961,N_29952);
nand UO_3413 (O_3413,N_29838,N_29857);
or UO_3414 (O_3414,N_29817,N_29774);
or UO_3415 (O_3415,N_29948,N_29746);
or UO_3416 (O_3416,N_29983,N_29756);
nor UO_3417 (O_3417,N_29729,N_29536);
and UO_3418 (O_3418,N_29892,N_29528);
and UO_3419 (O_3419,N_29555,N_29879);
and UO_3420 (O_3420,N_29881,N_29914);
and UO_3421 (O_3421,N_29664,N_29895);
nand UO_3422 (O_3422,N_29727,N_29826);
nor UO_3423 (O_3423,N_29976,N_29908);
and UO_3424 (O_3424,N_29639,N_29614);
nor UO_3425 (O_3425,N_29799,N_29675);
and UO_3426 (O_3426,N_29834,N_29623);
xnor UO_3427 (O_3427,N_29719,N_29609);
xnor UO_3428 (O_3428,N_29540,N_29678);
nor UO_3429 (O_3429,N_29528,N_29627);
or UO_3430 (O_3430,N_29993,N_29825);
nand UO_3431 (O_3431,N_29594,N_29611);
nor UO_3432 (O_3432,N_29593,N_29911);
nand UO_3433 (O_3433,N_29755,N_29757);
and UO_3434 (O_3434,N_29917,N_29791);
nor UO_3435 (O_3435,N_29546,N_29907);
nor UO_3436 (O_3436,N_29569,N_29690);
or UO_3437 (O_3437,N_29870,N_29891);
and UO_3438 (O_3438,N_29505,N_29787);
nand UO_3439 (O_3439,N_29548,N_29667);
nand UO_3440 (O_3440,N_29642,N_29574);
nand UO_3441 (O_3441,N_29873,N_29916);
or UO_3442 (O_3442,N_29727,N_29960);
nor UO_3443 (O_3443,N_29828,N_29860);
xor UO_3444 (O_3444,N_29887,N_29713);
nand UO_3445 (O_3445,N_29833,N_29795);
xor UO_3446 (O_3446,N_29725,N_29707);
and UO_3447 (O_3447,N_29969,N_29584);
and UO_3448 (O_3448,N_29711,N_29880);
nand UO_3449 (O_3449,N_29827,N_29571);
or UO_3450 (O_3450,N_29745,N_29914);
nand UO_3451 (O_3451,N_29775,N_29848);
or UO_3452 (O_3452,N_29665,N_29620);
or UO_3453 (O_3453,N_29541,N_29867);
xor UO_3454 (O_3454,N_29793,N_29669);
nor UO_3455 (O_3455,N_29672,N_29614);
xnor UO_3456 (O_3456,N_29507,N_29705);
nand UO_3457 (O_3457,N_29543,N_29650);
nand UO_3458 (O_3458,N_29634,N_29736);
nor UO_3459 (O_3459,N_29907,N_29938);
and UO_3460 (O_3460,N_29666,N_29568);
nor UO_3461 (O_3461,N_29852,N_29702);
nand UO_3462 (O_3462,N_29615,N_29888);
xnor UO_3463 (O_3463,N_29634,N_29897);
nand UO_3464 (O_3464,N_29631,N_29754);
xor UO_3465 (O_3465,N_29755,N_29519);
or UO_3466 (O_3466,N_29726,N_29538);
and UO_3467 (O_3467,N_29649,N_29558);
or UO_3468 (O_3468,N_29919,N_29540);
and UO_3469 (O_3469,N_29635,N_29847);
xor UO_3470 (O_3470,N_29860,N_29644);
xnor UO_3471 (O_3471,N_29859,N_29710);
or UO_3472 (O_3472,N_29503,N_29666);
and UO_3473 (O_3473,N_29803,N_29960);
or UO_3474 (O_3474,N_29945,N_29725);
nor UO_3475 (O_3475,N_29891,N_29745);
xor UO_3476 (O_3476,N_29693,N_29755);
nor UO_3477 (O_3477,N_29569,N_29917);
nor UO_3478 (O_3478,N_29609,N_29976);
or UO_3479 (O_3479,N_29766,N_29668);
xor UO_3480 (O_3480,N_29572,N_29824);
and UO_3481 (O_3481,N_29961,N_29636);
nor UO_3482 (O_3482,N_29817,N_29845);
nor UO_3483 (O_3483,N_29875,N_29598);
nand UO_3484 (O_3484,N_29621,N_29905);
nor UO_3485 (O_3485,N_29864,N_29663);
or UO_3486 (O_3486,N_29946,N_29922);
nor UO_3487 (O_3487,N_29901,N_29928);
and UO_3488 (O_3488,N_29517,N_29723);
nor UO_3489 (O_3489,N_29901,N_29529);
nor UO_3490 (O_3490,N_29757,N_29555);
xnor UO_3491 (O_3491,N_29675,N_29714);
or UO_3492 (O_3492,N_29739,N_29540);
nand UO_3493 (O_3493,N_29691,N_29906);
nor UO_3494 (O_3494,N_29743,N_29691);
nor UO_3495 (O_3495,N_29874,N_29863);
nor UO_3496 (O_3496,N_29870,N_29554);
nor UO_3497 (O_3497,N_29975,N_29712);
xnor UO_3498 (O_3498,N_29860,N_29771);
xor UO_3499 (O_3499,N_29661,N_29938);
endmodule