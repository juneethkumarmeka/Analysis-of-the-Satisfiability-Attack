module basic_750_5000_1000_5_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_594,In_412);
nor U1 (N_1,In_558,In_646);
nand U2 (N_2,In_458,In_358);
nand U3 (N_3,In_562,In_53);
or U4 (N_4,In_566,In_693);
or U5 (N_5,In_213,In_507);
and U6 (N_6,In_694,In_99);
nor U7 (N_7,In_433,In_407);
or U8 (N_8,In_712,In_255);
nor U9 (N_9,In_557,In_378);
and U10 (N_10,In_253,In_573);
xnor U11 (N_11,In_595,In_263);
and U12 (N_12,In_181,In_219);
nor U13 (N_13,In_245,In_674);
nor U14 (N_14,In_70,In_110);
nor U15 (N_15,In_454,In_576);
nor U16 (N_16,In_277,In_715);
or U17 (N_17,In_603,In_88);
or U18 (N_18,In_406,In_740);
or U19 (N_19,In_626,In_442);
or U20 (N_20,In_112,In_288);
nand U21 (N_21,In_12,In_105);
nor U22 (N_22,In_249,In_119);
or U23 (N_23,In_50,In_178);
or U24 (N_24,In_14,In_260);
nand U25 (N_25,In_68,In_164);
and U26 (N_26,In_191,In_92);
nand U27 (N_27,In_203,In_738);
or U28 (N_28,In_739,In_415);
and U29 (N_29,In_103,In_609);
nor U30 (N_30,In_652,In_536);
or U31 (N_31,In_294,In_328);
or U32 (N_32,In_259,In_138);
nor U33 (N_33,In_79,In_610);
nor U34 (N_34,In_123,In_656);
nand U35 (N_35,In_32,In_354);
nor U36 (N_36,In_719,In_23);
nand U37 (N_37,In_657,In_720);
or U38 (N_38,In_71,In_227);
and U39 (N_39,In_15,In_612);
and U40 (N_40,In_379,In_311);
or U41 (N_41,In_539,In_645);
and U42 (N_42,In_630,In_198);
nor U43 (N_43,In_727,In_350);
or U44 (N_44,In_301,In_93);
nand U45 (N_45,In_672,In_220);
xor U46 (N_46,In_96,In_601);
or U47 (N_47,In_347,In_139);
nor U48 (N_48,In_560,In_0);
nor U49 (N_49,In_469,In_450);
nor U50 (N_50,In_737,In_546);
and U51 (N_51,In_239,In_658);
or U52 (N_52,In_401,In_729);
and U53 (N_53,In_532,In_503);
or U54 (N_54,In_383,In_335);
and U55 (N_55,In_614,In_592);
nor U56 (N_56,In_184,In_207);
or U57 (N_57,In_555,In_486);
or U58 (N_58,In_64,In_188);
nand U59 (N_59,In_212,In_726);
or U60 (N_60,In_586,In_685);
or U61 (N_61,In_686,In_129);
and U62 (N_62,In_522,In_28);
nor U63 (N_63,In_448,In_159);
nor U64 (N_64,In_228,In_535);
and U65 (N_65,In_437,In_638);
or U66 (N_66,In_63,In_393);
and U67 (N_67,In_215,In_19);
or U68 (N_68,In_517,In_77);
and U69 (N_69,In_167,In_363);
nand U70 (N_70,In_380,In_473);
and U71 (N_71,In_598,In_366);
and U72 (N_72,In_183,In_474);
nand U73 (N_73,In_514,In_137);
and U74 (N_74,In_484,In_297);
nand U75 (N_75,In_35,In_196);
and U76 (N_76,In_143,In_650);
or U77 (N_77,In_571,In_244);
and U78 (N_78,In_548,In_281);
or U79 (N_79,In_154,In_695);
or U80 (N_80,In_736,In_216);
nor U81 (N_81,In_190,In_156);
nor U82 (N_82,In_243,In_3);
nor U83 (N_83,In_37,In_318);
or U84 (N_84,In_648,In_420);
and U85 (N_85,In_563,In_118);
nand U86 (N_86,In_16,In_635);
and U87 (N_87,In_660,In_290);
or U88 (N_88,In_195,In_404);
nand U89 (N_89,In_459,In_682);
nand U90 (N_90,In_482,In_722);
or U91 (N_91,In_287,In_157);
or U92 (N_92,In_218,In_31);
nand U93 (N_93,In_743,In_606);
or U94 (N_94,In_531,In_394);
nand U95 (N_95,In_233,In_422);
and U96 (N_96,In_189,In_483);
and U97 (N_97,In_307,In_644);
or U98 (N_98,In_599,In_545);
nand U99 (N_99,In_206,In_197);
or U100 (N_100,In_440,In_174);
or U101 (N_101,In_647,In_126);
and U102 (N_102,In_374,In_411);
nand U103 (N_103,In_225,In_247);
nand U104 (N_104,In_240,In_149);
and U105 (N_105,In_276,In_632);
or U106 (N_106,In_567,In_106);
xnor U107 (N_107,In_526,In_707);
or U108 (N_108,In_516,In_359);
nand U109 (N_109,In_403,In_543);
nor U110 (N_110,In_730,In_279);
nand U111 (N_111,In_29,In_510);
nor U112 (N_112,In_339,In_529);
or U113 (N_113,In_349,In_67);
or U114 (N_114,In_701,In_716);
and U115 (N_115,In_631,In_55);
nand U116 (N_116,In_177,In_187);
and U117 (N_117,In_629,In_564);
nor U118 (N_118,In_170,In_7);
nand U119 (N_119,In_390,In_130);
nand U120 (N_120,In_742,In_34);
and U121 (N_121,In_271,In_713);
xnor U122 (N_122,In_201,In_725);
and U123 (N_123,In_425,In_361);
nand U124 (N_124,In_579,In_127);
nor U125 (N_125,In_659,In_222);
nor U126 (N_126,In_231,In_210);
nand U127 (N_127,In_661,In_398);
or U128 (N_128,In_534,In_278);
or U129 (N_129,In_549,In_597);
and U130 (N_130,In_698,In_365);
nor U131 (N_131,In_423,In_85);
nor U132 (N_132,In_264,In_302);
and U133 (N_133,In_33,In_10);
nand U134 (N_134,In_100,In_395);
or U135 (N_135,In_296,In_224);
nand U136 (N_136,In_321,In_9);
and U137 (N_137,In_747,In_97);
and U138 (N_138,In_111,In_27);
nor U139 (N_139,In_475,In_43);
or U140 (N_140,In_460,In_688);
nand U141 (N_141,In_465,In_286);
or U142 (N_142,In_495,In_320);
or U143 (N_143,In_42,In_690);
and U144 (N_144,In_133,In_581);
and U145 (N_145,In_387,In_551);
xor U146 (N_146,In_351,In_17);
nor U147 (N_147,In_687,In_509);
nor U148 (N_148,In_4,In_691);
xnor U149 (N_149,In_257,In_434);
or U150 (N_150,In_357,In_541);
and U151 (N_151,In_427,In_508);
nor U152 (N_152,In_678,In_405);
or U153 (N_153,In_455,In_39);
nand U154 (N_154,In_325,In_410);
and U155 (N_155,In_462,In_500);
or U156 (N_156,In_41,In_283);
or U157 (N_157,In_709,In_499);
and U158 (N_158,In_40,In_641);
or U159 (N_159,In_270,In_73);
or U160 (N_160,In_82,In_699);
and U161 (N_161,In_221,In_578);
nor U162 (N_162,In_51,In_329);
nor U163 (N_163,In_104,In_413);
nor U164 (N_164,In_449,In_700);
nand U165 (N_165,In_356,In_147);
and U166 (N_166,In_616,In_223);
nand U167 (N_167,In_236,In_131);
or U168 (N_168,In_5,In_205);
nand U169 (N_169,In_511,In_368);
or U170 (N_170,In_141,In_204);
nand U171 (N_171,In_280,In_346);
and U172 (N_172,In_731,In_128);
or U173 (N_173,In_65,In_538);
nand U174 (N_174,In_266,In_445);
or U175 (N_175,In_81,In_340);
or U176 (N_176,In_303,In_319);
nor U177 (N_177,In_671,In_663);
or U178 (N_178,In_692,In_113);
nand U179 (N_179,In_336,In_735);
nor U180 (N_180,In_467,In_91);
or U181 (N_181,In_424,In_36);
nand U182 (N_182,In_684,In_337);
nor U183 (N_183,In_705,In_584);
and U184 (N_184,In_45,In_618);
nand U185 (N_185,In_386,In_176);
or U186 (N_186,In_62,In_444);
and U187 (N_187,In_76,In_25);
and U188 (N_188,In_642,In_491);
nor U189 (N_189,In_275,In_324);
and U190 (N_190,In_284,In_679);
and U191 (N_191,In_285,In_140);
or U192 (N_192,In_670,In_464);
nor U193 (N_193,In_680,In_314);
or U194 (N_194,In_282,In_57);
and U195 (N_195,In_565,In_162);
and U196 (N_196,In_1,In_744);
and U197 (N_197,In_478,In_6);
and U198 (N_198,In_733,In_590);
nand U199 (N_199,In_317,In_417);
or U200 (N_200,In_388,In_683);
nor U201 (N_201,In_323,In_367);
and U202 (N_202,In_74,In_497);
or U203 (N_203,In_636,In_362);
xor U204 (N_204,In_498,In_291);
or U205 (N_205,In_18,In_577);
nand U206 (N_206,In_135,In_217);
nand U207 (N_207,In_116,In_504);
nand U208 (N_208,In_226,In_588);
nor U209 (N_209,In_496,In_211);
and U210 (N_210,In_298,In_418);
nand U211 (N_211,In_621,In_268);
or U212 (N_212,In_521,In_145);
or U213 (N_213,In_554,In_471);
and U214 (N_214,In_721,In_430);
nand U215 (N_215,In_515,In_250);
nor U216 (N_216,In_265,In_269);
nor U217 (N_217,In_108,In_615);
nor U218 (N_218,In_466,In_477);
or U219 (N_219,In_408,In_341);
or U220 (N_220,In_668,In_355);
nand U221 (N_221,In_468,In_664);
or U222 (N_222,In_171,In_429);
and U223 (N_223,In_527,In_476);
nor U224 (N_224,In_107,In_414);
nand U225 (N_225,In_728,In_300);
and U226 (N_226,In_26,In_561);
nand U227 (N_227,In_540,In_348);
and U228 (N_228,In_666,In_193);
nor U229 (N_229,In_710,In_622);
and U230 (N_230,In_272,In_593);
nand U231 (N_231,In_559,In_375);
nor U232 (N_232,In_242,In_2);
nand U233 (N_233,In_547,In_256);
or U234 (N_234,In_24,In_61);
or U235 (N_235,In_186,In_152);
and U236 (N_236,In_463,In_182);
or U237 (N_237,In_80,In_261);
xor U238 (N_238,In_506,In_345);
and U239 (N_239,In_47,In_583);
and U240 (N_240,In_185,In_155);
nand U241 (N_241,In_436,In_708);
or U242 (N_242,In_158,In_640);
nor U243 (N_243,In_479,In_132);
nand U244 (N_244,In_304,In_397);
nand U245 (N_245,In_432,In_550);
or U246 (N_246,In_501,In_741);
nor U247 (N_247,In_98,In_489);
nor U248 (N_248,In_370,In_146);
and U249 (N_249,In_246,In_617);
and U250 (N_250,In_518,In_274);
nor U251 (N_251,In_734,In_173);
and U252 (N_252,In_267,In_421);
or U253 (N_253,In_519,In_381);
nor U254 (N_254,In_21,In_125);
or U255 (N_255,In_711,In_675);
nand U256 (N_256,In_306,In_717);
xnor U257 (N_257,In_627,In_487);
nor U258 (N_258,In_530,In_343);
or U259 (N_259,In_673,In_293);
and U260 (N_260,In_447,In_214);
nand U261 (N_261,In_600,In_60);
and U262 (N_262,In_456,In_585);
nor U263 (N_263,In_78,In_101);
or U264 (N_264,In_299,In_46);
nand U265 (N_265,In_704,In_655);
or U266 (N_266,In_689,In_435);
or U267 (N_267,In_575,In_52);
nand U268 (N_268,In_706,In_409);
or U269 (N_269,In_331,In_371);
nor U270 (N_270,In_192,In_625);
and U271 (N_271,In_537,In_124);
or U272 (N_272,In_724,In_443);
nand U273 (N_273,In_238,In_502);
and U274 (N_274,In_373,In_122);
nand U275 (N_275,In_179,In_230);
nor U276 (N_276,In_544,In_69);
and U277 (N_277,In_634,In_669);
nor U278 (N_278,In_38,In_117);
nor U279 (N_279,In_382,In_392);
or U280 (N_280,In_94,In_121);
nor U281 (N_281,In_485,In_142);
nor U282 (N_282,In_396,In_322);
nor U283 (N_283,In_254,In_248);
nand U284 (N_284,In_574,In_20);
xor U285 (N_285,In_513,In_651);
and U286 (N_286,In_95,In_22);
or U287 (N_287,In_653,In_326);
nor U288 (N_288,In_732,In_505);
nor U289 (N_289,In_533,In_419);
and U290 (N_290,In_718,In_151);
xor U291 (N_291,In_258,In_385);
nor U292 (N_292,In_237,In_470);
or U293 (N_293,In_384,In_480);
nor U294 (N_294,In_611,In_589);
or U295 (N_295,In_439,In_490);
nor U296 (N_296,In_49,In_89);
and U297 (N_297,In_332,In_662);
nor U298 (N_298,In_524,In_613);
nand U299 (N_299,In_369,In_667);
and U300 (N_300,In_461,In_569);
nor U301 (N_301,In_623,In_607);
nand U302 (N_302,In_702,In_234);
and U303 (N_303,In_552,In_344);
or U304 (N_304,In_628,In_54);
or U305 (N_305,In_570,In_637);
or U306 (N_306,In_66,In_180);
and U307 (N_307,In_209,In_426);
and U308 (N_308,In_208,In_639);
nand U309 (N_309,In_457,In_310);
nor U310 (N_310,In_372,In_619);
nand U311 (N_311,In_745,In_169);
or U312 (N_312,In_488,In_316);
and U313 (N_313,In_90,In_165);
nor U314 (N_314,In_229,In_148);
or U315 (N_315,In_161,In_289);
nor U316 (N_316,In_441,In_313);
nand U317 (N_317,In_451,In_714);
and U318 (N_318,In_523,In_59);
nor U319 (N_319,In_528,In_746);
nand U320 (N_320,In_30,In_232);
or U321 (N_321,In_696,In_153);
and U322 (N_322,In_525,In_72);
nand U323 (N_323,In_481,In_494);
and U324 (N_324,In_360,In_199);
nand U325 (N_325,In_572,In_472);
or U326 (N_326,In_602,In_391);
xnor U327 (N_327,In_172,In_308);
and U328 (N_328,In_431,In_723);
and U329 (N_329,In_115,In_163);
nor U330 (N_330,In_334,In_13);
nand U331 (N_331,In_333,In_377);
or U332 (N_332,In_633,In_512);
or U333 (N_333,In_262,In_428);
nor U334 (N_334,In_86,In_150);
or U335 (N_335,In_352,In_399);
nor U336 (N_336,In_677,In_200);
nor U337 (N_337,In_315,In_654);
nand U338 (N_338,In_620,In_376);
nand U339 (N_339,In_312,In_273);
or U340 (N_340,In_175,In_202);
or U341 (N_341,In_241,In_703);
and U342 (N_342,In_568,In_166);
nand U343 (N_343,In_136,In_330);
and U344 (N_344,In_649,In_48);
nor U345 (N_345,In_587,In_416);
xor U346 (N_346,In_605,In_748);
nor U347 (N_347,In_114,In_102);
and U348 (N_348,In_327,In_643);
nor U349 (N_349,In_292,In_305);
or U350 (N_350,In_520,In_542);
or U351 (N_351,In_84,In_252);
nand U352 (N_352,In_342,In_83);
nand U353 (N_353,In_402,In_553);
and U354 (N_354,In_11,In_446);
and U355 (N_355,In_295,In_452);
or U356 (N_356,In_160,In_580);
or U357 (N_357,In_400,In_8);
nand U358 (N_358,In_251,In_604);
xor U359 (N_359,In_608,In_665);
or U360 (N_360,In_582,In_87);
and U361 (N_361,In_364,In_44);
nor U362 (N_362,In_624,In_168);
and U363 (N_363,In_453,In_75);
and U364 (N_364,In_353,In_492);
nand U365 (N_365,In_438,In_194);
or U366 (N_366,In_58,In_556);
and U367 (N_367,In_596,In_338);
nor U368 (N_368,In_681,In_749);
or U369 (N_369,In_109,In_676);
nand U370 (N_370,In_235,In_697);
nor U371 (N_371,In_493,In_134);
nand U372 (N_372,In_309,In_144);
nand U373 (N_373,In_120,In_389);
nand U374 (N_374,In_56,In_591);
nor U375 (N_375,In_364,In_481);
or U376 (N_376,In_438,In_96);
and U377 (N_377,In_157,In_649);
and U378 (N_378,In_507,In_643);
or U379 (N_379,In_445,In_361);
or U380 (N_380,In_67,In_725);
nand U381 (N_381,In_581,In_482);
and U382 (N_382,In_707,In_120);
or U383 (N_383,In_71,In_441);
nor U384 (N_384,In_465,In_108);
nand U385 (N_385,In_363,In_439);
nor U386 (N_386,In_30,In_362);
and U387 (N_387,In_236,In_298);
and U388 (N_388,In_709,In_473);
or U389 (N_389,In_344,In_616);
or U390 (N_390,In_640,In_219);
nand U391 (N_391,In_435,In_618);
or U392 (N_392,In_229,In_190);
nor U393 (N_393,In_463,In_459);
nor U394 (N_394,In_626,In_216);
nor U395 (N_395,In_31,In_470);
and U396 (N_396,In_119,In_83);
or U397 (N_397,In_600,In_145);
and U398 (N_398,In_643,In_648);
nor U399 (N_399,In_428,In_484);
or U400 (N_400,In_300,In_729);
nand U401 (N_401,In_637,In_616);
and U402 (N_402,In_147,In_128);
and U403 (N_403,In_415,In_268);
nand U404 (N_404,In_159,In_290);
nand U405 (N_405,In_439,In_207);
and U406 (N_406,In_514,In_191);
and U407 (N_407,In_135,In_403);
or U408 (N_408,In_94,In_290);
nor U409 (N_409,In_454,In_688);
and U410 (N_410,In_239,In_630);
nor U411 (N_411,In_146,In_219);
nor U412 (N_412,In_606,In_228);
nand U413 (N_413,In_29,In_160);
nor U414 (N_414,In_74,In_73);
and U415 (N_415,In_538,In_137);
and U416 (N_416,In_332,In_369);
and U417 (N_417,In_372,In_120);
nand U418 (N_418,In_394,In_217);
nor U419 (N_419,In_343,In_580);
and U420 (N_420,In_454,In_224);
nand U421 (N_421,In_456,In_665);
and U422 (N_422,In_373,In_223);
xnor U423 (N_423,In_99,In_50);
nor U424 (N_424,In_708,In_300);
nor U425 (N_425,In_81,In_488);
or U426 (N_426,In_538,In_309);
or U427 (N_427,In_291,In_623);
and U428 (N_428,In_320,In_612);
or U429 (N_429,In_151,In_289);
nand U430 (N_430,In_178,In_424);
nand U431 (N_431,In_268,In_166);
and U432 (N_432,In_406,In_617);
or U433 (N_433,In_283,In_127);
nor U434 (N_434,In_727,In_527);
or U435 (N_435,In_222,In_661);
and U436 (N_436,In_542,In_154);
nor U437 (N_437,In_597,In_258);
nor U438 (N_438,In_283,In_219);
or U439 (N_439,In_170,In_601);
or U440 (N_440,In_435,In_576);
nor U441 (N_441,In_5,In_501);
or U442 (N_442,In_388,In_105);
or U443 (N_443,In_387,In_607);
xnor U444 (N_444,In_525,In_1);
xnor U445 (N_445,In_563,In_140);
or U446 (N_446,In_419,In_637);
nor U447 (N_447,In_224,In_90);
and U448 (N_448,In_635,In_583);
or U449 (N_449,In_28,In_345);
or U450 (N_450,In_304,In_632);
and U451 (N_451,In_425,In_194);
and U452 (N_452,In_209,In_171);
or U453 (N_453,In_223,In_15);
nand U454 (N_454,In_665,In_649);
nand U455 (N_455,In_172,In_670);
nand U456 (N_456,In_351,In_160);
or U457 (N_457,In_533,In_554);
nor U458 (N_458,In_323,In_112);
nand U459 (N_459,In_314,In_699);
nor U460 (N_460,In_614,In_518);
nand U461 (N_461,In_725,In_27);
nand U462 (N_462,In_702,In_241);
nand U463 (N_463,In_47,In_293);
or U464 (N_464,In_743,In_456);
and U465 (N_465,In_280,In_685);
nand U466 (N_466,In_706,In_41);
and U467 (N_467,In_474,In_9);
nand U468 (N_468,In_161,In_561);
nand U469 (N_469,In_374,In_543);
or U470 (N_470,In_171,In_718);
nor U471 (N_471,In_739,In_45);
and U472 (N_472,In_245,In_382);
and U473 (N_473,In_80,In_537);
nor U474 (N_474,In_437,In_443);
and U475 (N_475,In_107,In_652);
nor U476 (N_476,In_22,In_591);
or U477 (N_477,In_183,In_98);
and U478 (N_478,In_339,In_240);
nor U479 (N_479,In_211,In_29);
nor U480 (N_480,In_268,In_531);
nand U481 (N_481,In_699,In_496);
nor U482 (N_482,In_647,In_43);
nor U483 (N_483,In_736,In_722);
nand U484 (N_484,In_80,In_15);
and U485 (N_485,In_707,In_433);
or U486 (N_486,In_506,In_647);
nor U487 (N_487,In_456,In_736);
xor U488 (N_488,In_168,In_285);
nor U489 (N_489,In_65,In_328);
nor U490 (N_490,In_25,In_493);
nand U491 (N_491,In_206,In_7);
nand U492 (N_492,In_659,In_594);
and U493 (N_493,In_221,In_47);
or U494 (N_494,In_445,In_2);
or U495 (N_495,In_260,In_230);
nor U496 (N_496,In_389,In_205);
nor U497 (N_497,In_691,In_306);
nor U498 (N_498,In_272,In_433);
or U499 (N_499,In_292,In_554);
and U500 (N_500,In_507,In_4);
nor U501 (N_501,In_551,In_617);
or U502 (N_502,In_409,In_402);
xnor U503 (N_503,In_180,In_113);
nand U504 (N_504,In_17,In_465);
and U505 (N_505,In_34,In_316);
and U506 (N_506,In_206,In_186);
nand U507 (N_507,In_120,In_11);
or U508 (N_508,In_7,In_564);
nor U509 (N_509,In_564,In_529);
or U510 (N_510,In_276,In_377);
and U511 (N_511,In_159,In_277);
nand U512 (N_512,In_154,In_434);
nand U513 (N_513,In_519,In_160);
nor U514 (N_514,In_160,In_495);
or U515 (N_515,In_592,In_169);
nand U516 (N_516,In_465,In_481);
nor U517 (N_517,In_81,In_112);
and U518 (N_518,In_218,In_409);
nand U519 (N_519,In_1,In_22);
or U520 (N_520,In_337,In_489);
or U521 (N_521,In_633,In_681);
nand U522 (N_522,In_522,In_75);
or U523 (N_523,In_64,In_450);
nand U524 (N_524,In_83,In_207);
and U525 (N_525,In_304,In_357);
xor U526 (N_526,In_677,In_142);
or U527 (N_527,In_19,In_594);
nor U528 (N_528,In_310,In_74);
and U529 (N_529,In_395,In_250);
or U530 (N_530,In_683,In_41);
and U531 (N_531,In_205,In_449);
nand U532 (N_532,In_26,In_166);
and U533 (N_533,In_390,In_510);
nand U534 (N_534,In_350,In_347);
nand U535 (N_535,In_188,In_627);
and U536 (N_536,In_619,In_349);
and U537 (N_537,In_454,In_517);
and U538 (N_538,In_610,In_454);
nor U539 (N_539,In_134,In_706);
nand U540 (N_540,In_119,In_487);
nor U541 (N_541,In_723,In_257);
nand U542 (N_542,In_371,In_367);
and U543 (N_543,In_190,In_651);
or U544 (N_544,In_560,In_169);
or U545 (N_545,In_262,In_277);
and U546 (N_546,In_150,In_169);
nor U547 (N_547,In_466,In_675);
nand U548 (N_548,In_396,In_111);
or U549 (N_549,In_82,In_409);
nand U550 (N_550,In_355,In_46);
and U551 (N_551,In_425,In_221);
nor U552 (N_552,In_544,In_699);
and U553 (N_553,In_695,In_428);
or U554 (N_554,In_481,In_424);
nand U555 (N_555,In_28,In_97);
or U556 (N_556,In_601,In_337);
and U557 (N_557,In_64,In_306);
xor U558 (N_558,In_484,In_23);
nand U559 (N_559,In_309,In_653);
nor U560 (N_560,In_480,In_390);
nor U561 (N_561,In_635,In_368);
and U562 (N_562,In_316,In_466);
or U563 (N_563,In_265,In_87);
xnor U564 (N_564,In_242,In_615);
and U565 (N_565,In_350,In_619);
or U566 (N_566,In_422,In_354);
and U567 (N_567,In_117,In_185);
nor U568 (N_568,In_94,In_349);
or U569 (N_569,In_24,In_525);
and U570 (N_570,In_355,In_657);
or U571 (N_571,In_538,In_542);
nor U572 (N_572,In_437,In_642);
and U573 (N_573,In_545,In_605);
nand U574 (N_574,In_154,In_699);
and U575 (N_575,In_106,In_708);
or U576 (N_576,In_498,In_493);
and U577 (N_577,In_352,In_278);
nor U578 (N_578,In_654,In_120);
and U579 (N_579,In_19,In_633);
or U580 (N_580,In_123,In_125);
and U581 (N_581,In_453,In_648);
or U582 (N_582,In_482,In_648);
nor U583 (N_583,In_58,In_395);
nor U584 (N_584,In_367,In_365);
nor U585 (N_585,In_44,In_524);
xnor U586 (N_586,In_26,In_695);
and U587 (N_587,In_73,In_16);
nand U588 (N_588,In_147,In_223);
or U589 (N_589,In_510,In_527);
or U590 (N_590,In_171,In_104);
or U591 (N_591,In_512,In_188);
or U592 (N_592,In_53,In_696);
or U593 (N_593,In_317,In_455);
or U594 (N_594,In_697,In_727);
nand U595 (N_595,In_264,In_103);
or U596 (N_596,In_356,In_704);
or U597 (N_597,In_411,In_172);
nor U598 (N_598,In_171,In_410);
and U599 (N_599,In_470,In_661);
and U600 (N_600,In_554,In_432);
nor U601 (N_601,In_396,In_120);
or U602 (N_602,In_502,In_655);
or U603 (N_603,In_575,In_663);
or U604 (N_604,In_388,In_734);
nand U605 (N_605,In_338,In_307);
or U606 (N_606,In_516,In_481);
and U607 (N_607,In_308,In_151);
or U608 (N_608,In_74,In_91);
or U609 (N_609,In_514,In_503);
nand U610 (N_610,In_333,In_516);
nand U611 (N_611,In_62,In_54);
or U612 (N_612,In_156,In_277);
nand U613 (N_613,In_621,In_251);
xor U614 (N_614,In_387,In_602);
nor U615 (N_615,In_622,In_56);
nand U616 (N_616,In_651,In_502);
and U617 (N_617,In_322,In_704);
and U618 (N_618,In_61,In_466);
and U619 (N_619,In_660,In_721);
or U620 (N_620,In_559,In_416);
or U621 (N_621,In_179,In_282);
or U622 (N_622,In_344,In_254);
nand U623 (N_623,In_258,In_151);
nand U624 (N_624,In_617,In_600);
nand U625 (N_625,In_78,In_345);
nor U626 (N_626,In_313,In_221);
or U627 (N_627,In_334,In_273);
nand U628 (N_628,In_717,In_329);
or U629 (N_629,In_491,In_464);
nor U630 (N_630,In_603,In_245);
nand U631 (N_631,In_718,In_475);
nor U632 (N_632,In_309,In_591);
nand U633 (N_633,In_571,In_190);
nand U634 (N_634,In_206,In_271);
nand U635 (N_635,In_345,In_572);
and U636 (N_636,In_176,In_392);
nand U637 (N_637,In_109,In_445);
and U638 (N_638,In_325,In_601);
nor U639 (N_639,In_91,In_560);
or U640 (N_640,In_371,In_313);
or U641 (N_641,In_300,In_594);
nor U642 (N_642,In_294,In_376);
or U643 (N_643,In_130,In_366);
xnor U644 (N_644,In_106,In_739);
nor U645 (N_645,In_194,In_472);
nand U646 (N_646,In_175,In_716);
and U647 (N_647,In_687,In_588);
or U648 (N_648,In_576,In_607);
or U649 (N_649,In_693,In_304);
nor U650 (N_650,In_426,In_671);
nor U651 (N_651,In_41,In_526);
nor U652 (N_652,In_535,In_380);
xnor U653 (N_653,In_590,In_631);
and U654 (N_654,In_213,In_271);
nor U655 (N_655,In_471,In_242);
nand U656 (N_656,In_569,In_23);
and U657 (N_657,In_77,In_10);
or U658 (N_658,In_640,In_188);
and U659 (N_659,In_564,In_31);
and U660 (N_660,In_479,In_437);
or U661 (N_661,In_141,In_34);
nand U662 (N_662,In_541,In_747);
nor U663 (N_663,In_108,In_448);
nand U664 (N_664,In_479,In_189);
or U665 (N_665,In_668,In_689);
nor U666 (N_666,In_365,In_586);
nor U667 (N_667,In_480,In_112);
nand U668 (N_668,In_412,In_742);
or U669 (N_669,In_308,In_157);
nor U670 (N_670,In_681,In_632);
and U671 (N_671,In_143,In_330);
or U672 (N_672,In_52,In_229);
nor U673 (N_673,In_342,In_720);
nand U674 (N_674,In_489,In_659);
and U675 (N_675,In_55,In_683);
and U676 (N_676,In_693,In_390);
nand U677 (N_677,In_425,In_517);
nor U678 (N_678,In_311,In_635);
nand U679 (N_679,In_436,In_282);
and U680 (N_680,In_190,In_368);
nand U681 (N_681,In_357,In_495);
or U682 (N_682,In_260,In_271);
nor U683 (N_683,In_116,In_279);
and U684 (N_684,In_290,In_84);
nor U685 (N_685,In_381,In_105);
nand U686 (N_686,In_423,In_356);
or U687 (N_687,In_632,In_462);
nand U688 (N_688,In_88,In_731);
nand U689 (N_689,In_572,In_275);
nand U690 (N_690,In_199,In_504);
nand U691 (N_691,In_687,In_199);
or U692 (N_692,In_365,In_288);
nor U693 (N_693,In_569,In_624);
and U694 (N_694,In_42,In_513);
nand U695 (N_695,In_226,In_186);
nor U696 (N_696,In_475,In_114);
nand U697 (N_697,In_628,In_277);
nand U698 (N_698,In_576,In_661);
and U699 (N_699,In_92,In_344);
nor U700 (N_700,In_672,In_443);
nor U701 (N_701,In_14,In_151);
nor U702 (N_702,In_219,In_732);
and U703 (N_703,In_701,In_402);
nand U704 (N_704,In_542,In_1);
nor U705 (N_705,In_485,In_640);
nor U706 (N_706,In_667,In_694);
and U707 (N_707,In_504,In_734);
nor U708 (N_708,In_400,In_108);
and U709 (N_709,In_74,In_476);
or U710 (N_710,In_63,In_557);
nand U711 (N_711,In_345,In_713);
or U712 (N_712,In_61,In_645);
nor U713 (N_713,In_606,In_80);
nand U714 (N_714,In_511,In_506);
nor U715 (N_715,In_739,In_666);
nand U716 (N_716,In_495,In_633);
and U717 (N_717,In_412,In_280);
nand U718 (N_718,In_380,In_252);
nand U719 (N_719,In_687,In_667);
or U720 (N_720,In_7,In_319);
nor U721 (N_721,In_102,In_115);
nand U722 (N_722,In_432,In_439);
nand U723 (N_723,In_90,In_271);
xnor U724 (N_724,In_511,In_233);
and U725 (N_725,In_42,In_504);
nand U726 (N_726,In_303,In_674);
nand U727 (N_727,In_238,In_450);
nor U728 (N_728,In_598,In_403);
nor U729 (N_729,In_75,In_359);
nand U730 (N_730,In_415,In_732);
xor U731 (N_731,In_32,In_424);
nor U732 (N_732,In_149,In_595);
and U733 (N_733,In_262,In_626);
or U734 (N_734,In_533,In_168);
nor U735 (N_735,In_716,In_15);
or U736 (N_736,In_356,In_267);
nor U737 (N_737,In_15,In_24);
and U738 (N_738,In_721,In_140);
or U739 (N_739,In_690,In_160);
nor U740 (N_740,In_13,In_470);
or U741 (N_741,In_21,In_328);
nand U742 (N_742,In_541,In_479);
and U743 (N_743,In_413,In_677);
or U744 (N_744,In_494,In_417);
nor U745 (N_745,In_744,In_302);
xor U746 (N_746,In_424,In_646);
and U747 (N_747,In_705,In_188);
and U748 (N_748,In_176,In_664);
or U749 (N_749,In_213,In_496);
nand U750 (N_750,In_318,In_593);
nor U751 (N_751,In_7,In_35);
or U752 (N_752,In_597,In_224);
and U753 (N_753,In_150,In_65);
nor U754 (N_754,In_380,In_136);
nor U755 (N_755,In_460,In_218);
and U756 (N_756,In_277,In_413);
and U757 (N_757,In_369,In_61);
and U758 (N_758,In_643,In_652);
or U759 (N_759,In_395,In_636);
nand U760 (N_760,In_728,In_122);
nand U761 (N_761,In_650,In_225);
or U762 (N_762,In_605,In_215);
nand U763 (N_763,In_185,In_468);
and U764 (N_764,In_85,In_392);
nand U765 (N_765,In_190,In_348);
nor U766 (N_766,In_387,In_431);
and U767 (N_767,In_409,In_607);
and U768 (N_768,In_180,In_57);
and U769 (N_769,In_410,In_351);
nor U770 (N_770,In_375,In_707);
and U771 (N_771,In_264,In_29);
nor U772 (N_772,In_544,In_119);
nand U773 (N_773,In_317,In_533);
nor U774 (N_774,In_499,In_635);
and U775 (N_775,In_502,In_261);
nor U776 (N_776,In_705,In_420);
nor U777 (N_777,In_188,In_501);
or U778 (N_778,In_82,In_669);
or U779 (N_779,In_199,In_312);
or U780 (N_780,In_384,In_120);
and U781 (N_781,In_55,In_699);
and U782 (N_782,In_327,In_701);
nand U783 (N_783,In_556,In_338);
and U784 (N_784,In_60,In_337);
and U785 (N_785,In_716,In_271);
nor U786 (N_786,In_599,In_657);
and U787 (N_787,In_424,In_443);
nand U788 (N_788,In_517,In_688);
nand U789 (N_789,In_458,In_371);
or U790 (N_790,In_563,In_310);
or U791 (N_791,In_110,In_62);
nand U792 (N_792,In_428,In_615);
nor U793 (N_793,In_189,In_411);
and U794 (N_794,In_16,In_474);
or U795 (N_795,In_349,In_577);
nor U796 (N_796,In_132,In_2);
nand U797 (N_797,In_221,In_718);
nand U798 (N_798,In_179,In_541);
nand U799 (N_799,In_485,In_662);
or U800 (N_800,In_453,In_444);
and U801 (N_801,In_388,In_722);
nand U802 (N_802,In_90,In_619);
nand U803 (N_803,In_144,In_664);
nor U804 (N_804,In_310,In_273);
nand U805 (N_805,In_212,In_415);
or U806 (N_806,In_496,In_22);
or U807 (N_807,In_453,In_499);
or U808 (N_808,In_665,In_590);
and U809 (N_809,In_730,In_207);
nand U810 (N_810,In_522,In_355);
nand U811 (N_811,In_601,In_468);
and U812 (N_812,In_315,In_282);
or U813 (N_813,In_511,In_120);
or U814 (N_814,In_328,In_114);
or U815 (N_815,In_423,In_205);
nand U816 (N_816,In_687,In_261);
nand U817 (N_817,In_673,In_272);
nor U818 (N_818,In_544,In_457);
and U819 (N_819,In_151,In_197);
xor U820 (N_820,In_79,In_661);
and U821 (N_821,In_669,In_535);
nor U822 (N_822,In_207,In_166);
and U823 (N_823,In_287,In_269);
or U824 (N_824,In_248,In_469);
and U825 (N_825,In_195,In_671);
nor U826 (N_826,In_571,In_257);
or U827 (N_827,In_397,In_494);
nand U828 (N_828,In_129,In_749);
and U829 (N_829,In_209,In_490);
and U830 (N_830,In_363,In_381);
or U831 (N_831,In_488,In_442);
and U832 (N_832,In_182,In_500);
or U833 (N_833,In_116,In_84);
nor U834 (N_834,In_339,In_317);
and U835 (N_835,In_474,In_632);
nor U836 (N_836,In_292,In_80);
or U837 (N_837,In_688,In_357);
nor U838 (N_838,In_643,In_480);
and U839 (N_839,In_82,In_507);
nor U840 (N_840,In_446,In_595);
and U841 (N_841,In_87,In_505);
nor U842 (N_842,In_647,In_738);
nand U843 (N_843,In_187,In_438);
or U844 (N_844,In_520,In_174);
and U845 (N_845,In_555,In_681);
and U846 (N_846,In_599,In_366);
and U847 (N_847,In_170,In_238);
nor U848 (N_848,In_476,In_612);
xor U849 (N_849,In_396,In_627);
nor U850 (N_850,In_71,In_279);
nand U851 (N_851,In_678,In_742);
or U852 (N_852,In_327,In_220);
and U853 (N_853,In_629,In_274);
nand U854 (N_854,In_334,In_201);
or U855 (N_855,In_532,In_79);
or U856 (N_856,In_1,In_499);
and U857 (N_857,In_208,In_543);
and U858 (N_858,In_617,In_540);
xnor U859 (N_859,In_21,In_650);
or U860 (N_860,In_579,In_292);
and U861 (N_861,In_296,In_678);
nand U862 (N_862,In_583,In_28);
or U863 (N_863,In_344,In_112);
and U864 (N_864,In_189,In_96);
and U865 (N_865,In_152,In_639);
nand U866 (N_866,In_534,In_48);
nand U867 (N_867,In_258,In_511);
nand U868 (N_868,In_575,In_284);
nor U869 (N_869,In_674,In_70);
or U870 (N_870,In_567,In_93);
and U871 (N_871,In_585,In_238);
nor U872 (N_872,In_583,In_214);
or U873 (N_873,In_446,In_43);
or U874 (N_874,In_190,In_333);
nand U875 (N_875,In_287,In_443);
and U876 (N_876,In_687,In_196);
nor U877 (N_877,In_267,In_451);
or U878 (N_878,In_144,In_125);
nand U879 (N_879,In_394,In_99);
nand U880 (N_880,In_39,In_339);
nor U881 (N_881,In_722,In_317);
and U882 (N_882,In_266,In_162);
or U883 (N_883,In_248,In_163);
or U884 (N_884,In_480,In_78);
nand U885 (N_885,In_101,In_112);
nand U886 (N_886,In_126,In_317);
nand U887 (N_887,In_637,In_645);
nand U888 (N_888,In_287,In_607);
nand U889 (N_889,In_214,In_484);
nor U890 (N_890,In_379,In_104);
and U891 (N_891,In_393,In_356);
nor U892 (N_892,In_83,In_664);
and U893 (N_893,In_665,In_173);
or U894 (N_894,In_533,In_538);
and U895 (N_895,In_589,In_145);
nand U896 (N_896,In_515,In_590);
or U897 (N_897,In_180,In_326);
and U898 (N_898,In_620,In_452);
or U899 (N_899,In_660,In_105);
and U900 (N_900,In_53,In_530);
nor U901 (N_901,In_81,In_52);
or U902 (N_902,In_552,In_264);
nor U903 (N_903,In_179,In_672);
and U904 (N_904,In_338,In_726);
and U905 (N_905,In_491,In_479);
or U906 (N_906,In_116,In_388);
and U907 (N_907,In_11,In_116);
or U908 (N_908,In_120,In_563);
and U909 (N_909,In_746,In_229);
nand U910 (N_910,In_388,In_711);
and U911 (N_911,In_256,In_316);
nand U912 (N_912,In_414,In_641);
nand U913 (N_913,In_673,In_206);
nand U914 (N_914,In_689,In_135);
nor U915 (N_915,In_437,In_136);
and U916 (N_916,In_198,In_230);
or U917 (N_917,In_526,In_673);
nand U918 (N_918,In_122,In_688);
or U919 (N_919,In_515,In_511);
or U920 (N_920,In_476,In_429);
or U921 (N_921,In_198,In_545);
or U922 (N_922,In_533,In_124);
nand U923 (N_923,In_674,In_107);
nor U924 (N_924,In_305,In_83);
nor U925 (N_925,In_691,In_46);
or U926 (N_926,In_316,In_467);
nor U927 (N_927,In_63,In_16);
nand U928 (N_928,In_310,In_712);
xnor U929 (N_929,In_280,In_244);
xor U930 (N_930,In_286,In_227);
nor U931 (N_931,In_232,In_495);
or U932 (N_932,In_527,In_180);
nor U933 (N_933,In_690,In_126);
and U934 (N_934,In_336,In_42);
or U935 (N_935,In_503,In_466);
or U936 (N_936,In_218,In_45);
and U937 (N_937,In_0,In_70);
nand U938 (N_938,In_393,In_470);
nor U939 (N_939,In_236,In_660);
nand U940 (N_940,In_415,In_736);
nor U941 (N_941,In_151,In_403);
or U942 (N_942,In_462,In_295);
nor U943 (N_943,In_559,In_488);
or U944 (N_944,In_714,In_705);
nand U945 (N_945,In_546,In_334);
nor U946 (N_946,In_639,In_515);
nor U947 (N_947,In_255,In_449);
nor U948 (N_948,In_466,In_731);
or U949 (N_949,In_191,In_176);
and U950 (N_950,In_47,In_522);
or U951 (N_951,In_244,In_563);
or U952 (N_952,In_274,In_546);
and U953 (N_953,In_157,In_475);
and U954 (N_954,In_305,In_12);
nor U955 (N_955,In_227,In_693);
or U956 (N_956,In_353,In_104);
and U957 (N_957,In_388,In_296);
and U958 (N_958,In_318,In_123);
or U959 (N_959,In_625,In_363);
or U960 (N_960,In_708,In_738);
nor U961 (N_961,In_461,In_735);
nand U962 (N_962,In_559,In_168);
or U963 (N_963,In_556,In_537);
nand U964 (N_964,In_434,In_339);
and U965 (N_965,In_452,In_190);
nor U966 (N_966,In_538,In_717);
or U967 (N_967,In_429,In_693);
nand U968 (N_968,In_5,In_352);
and U969 (N_969,In_159,In_236);
nand U970 (N_970,In_716,In_595);
nor U971 (N_971,In_549,In_141);
nor U972 (N_972,In_135,In_402);
nor U973 (N_973,In_183,In_734);
or U974 (N_974,In_585,In_131);
nand U975 (N_975,In_51,In_614);
and U976 (N_976,In_340,In_691);
and U977 (N_977,In_274,In_285);
or U978 (N_978,In_104,In_44);
nor U979 (N_979,In_677,In_82);
and U980 (N_980,In_411,In_321);
nor U981 (N_981,In_97,In_355);
nand U982 (N_982,In_514,In_583);
nand U983 (N_983,In_145,In_83);
or U984 (N_984,In_77,In_619);
and U985 (N_985,In_268,In_467);
or U986 (N_986,In_675,In_190);
nor U987 (N_987,In_553,In_181);
nor U988 (N_988,In_161,In_278);
and U989 (N_989,In_14,In_132);
or U990 (N_990,In_124,In_125);
or U991 (N_991,In_33,In_446);
or U992 (N_992,In_449,In_393);
nor U993 (N_993,In_524,In_133);
nor U994 (N_994,In_610,In_691);
or U995 (N_995,In_238,In_169);
or U996 (N_996,In_549,In_347);
and U997 (N_997,In_306,In_280);
nor U998 (N_998,In_195,In_202);
nor U999 (N_999,In_51,In_98);
or U1000 (N_1000,N_489,N_534);
and U1001 (N_1001,N_712,N_513);
and U1002 (N_1002,N_479,N_425);
and U1003 (N_1003,N_692,N_501);
or U1004 (N_1004,N_683,N_438);
or U1005 (N_1005,N_987,N_848);
or U1006 (N_1006,N_257,N_923);
nor U1007 (N_1007,N_263,N_540);
nor U1008 (N_1008,N_889,N_665);
nand U1009 (N_1009,N_57,N_51);
nor U1010 (N_1010,N_484,N_111);
nand U1011 (N_1011,N_556,N_217);
or U1012 (N_1012,N_364,N_41);
nand U1013 (N_1013,N_106,N_478);
or U1014 (N_1014,N_812,N_695);
nand U1015 (N_1015,N_197,N_509);
nand U1016 (N_1016,N_814,N_678);
nor U1017 (N_1017,N_351,N_633);
nand U1018 (N_1018,N_519,N_175);
xnor U1019 (N_1019,N_123,N_897);
nand U1020 (N_1020,N_223,N_24);
or U1021 (N_1021,N_718,N_754);
xnor U1022 (N_1022,N_492,N_433);
nor U1023 (N_1023,N_903,N_562);
nor U1024 (N_1024,N_370,N_729);
nor U1025 (N_1025,N_236,N_115);
nand U1026 (N_1026,N_886,N_73);
nor U1027 (N_1027,N_944,N_42);
or U1028 (N_1028,N_136,N_505);
and U1029 (N_1029,N_885,N_777);
and U1030 (N_1030,N_837,N_358);
nand U1031 (N_1031,N_843,N_663);
xnor U1032 (N_1032,N_486,N_644);
nor U1033 (N_1033,N_634,N_259);
xor U1034 (N_1034,N_823,N_635);
nor U1035 (N_1035,N_912,N_803);
xor U1036 (N_1036,N_183,N_563);
nor U1037 (N_1037,N_746,N_439);
nand U1038 (N_1038,N_228,N_258);
and U1039 (N_1039,N_272,N_165);
or U1040 (N_1040,N_961,N_442);
nand U1041 (N_1041,N_871,N_378);
or U1042 (N_1042,N_300,N_347);
nand U1043 (N_1043,N_649,N_977);
and U1044 (N_1044,N_161,N_291);
or U1045 (N_1045,N_594,N_753);
nor U1046 (N_1046,N_415,N_604);
nand U1047 (N_1047,N_884,N_137);
or U1048 (N_1048,N_572,N_834);
nand U1049 (N_1049,N_227,N_164);
or U1050 (N_1050,N_846,N_857);
nor U1051 (N_1051,N_577,N_172);
and U1052 (N_1052,N_968,N_25);
or U1053 (N_1053,N_743,N_598);
or U1054 (N_1054,N_87,N_770);
nor U1055 (N_1055,N_781,N_606);
nor U1056 (N_1056,N_662,N_715);
or U1057 (N_1057,N_946,N_945);
nand U1058 (N_1058,N_617,N_178);
nand U1059 (N_1059,N_711,N_219);
nand U1060 (N_1060,N_129,N_660);
nand U1061 (N_1061,N_995,N_811);
nor U1062 (N_1062,N_369,N_826);
xor U1063 (N_1063,N_174,N_639);
nand U1064 (N_1064,N_459,N_50);
nand U1065 (N_1065,N_21,N_608);
nand U1066 (N_1066,N_798,N_354);
and U1067 (N_1067,N_531,N_307);
and U1068 (N_1068,N_1,N_842);
nand U1069 (N_1069,N_595,N_497);
nand U1070 (N_1070,N_708,N_93);
or U1071 (N_1071,N_864,N_116);
xnor U1072 (N_1072,N_702,N_778);
or U1073 (N_1073,N_216,N_933);
nand U1074 (N_1074,N_282,N_52);
nor U1075 (N_1075,N_560,N_108);
or U1076 (N_1076,N_867,N_973);
or U1077 (N_1077,N_749,N_963);
nor U1078 (N_1078,N_851,N_265);
or U1079 (N_1079,N_461,N_422);
xor U1080 (N_1080,N_416,N_221);
nand U1081 (N_1081,N_631,N_186);
or U1082 (N_1082,N_460,N_187);
and U1083 (N_1083,N_671,N_703);
nor U1084 (N_1084,N_140,N_601);
or U1085 (N_1085,N_940,N_986);
and U1086 (N_1086,N_862,N_276);
nand U1087 (N_1087,N_239,N_962);
or U1088 (N_1088,N_975,N_687);
nand U1089 (N_1089,N_905,N_853);
and U1090 (N_1090,N_523,N_773);
nor U1091 (N_1091,N_85,N_592);
nand U1092 (N_1092,N_481,N_555);
and U1093 (N_1093,N_679,N_177);
and U1094 (N_1094,N_584,N_602);
nand U1095 (N_1095,N_440,N_487);
nor U1096 (N_1096,N_135,N_569);
nand U1097 (N_1097,N_371,N_261);
nand U1098 (N_1098,N_830,N_0);
nor U1099 (N_1099,N_648,N_386);
and U1100 (N_1100,N_532,N_689);
nand U1101 (N_1101,N_407,N_469);
nor U1102 (N_1102,N_810,N_482);
or U1103 (N_1103,N_820,N_318);
nor U1104 (N_1104,N_201,N_965);
and U1105 (N_1105,N_338,N_767);
and U1106 (N_1106,N_822,N_76);
nor U1107 (N_1107,N_697,N_854);
nor U1108 (N_1108,N_794,N_713);
nand U1109 (N_1109,N_881,N_898);
nor U1110 (N_1110,N_654,N_467);
or U1111 (N_1111,N_349,N_793);
nand U1112 (N_1112,N_567,N_225);
nor U1113 (N_1113,N_808,N_657);
or U1114 (N_1114,N_141,N_143);
xnor U1115 (N_1115,N_868,N_974);
nor U1116 (N_1116,N_199,N_355);
nor U1117 (N_1117,N_262,N_22);
and U1118 (N_1118,N_816,N_499);
nor U1119 (N_1119,N_458,N_53);
or U1120 (N_1120,N_647,N_163);
or U1121 (N_1121,N_270,N_833);
nor U1122 (N_1122,N_296,N_67);
and U1123 (N_1123,N_651,N_151);
or U1124 (N_1124,N_421,N_858);
or U1125 (N_1125,N_443,N_786);
and U1126 (N_1126,N_142,N_312);
nand U1127 (N_1127,N_894,N_930);
and U1128 (N_1128,N_526,N_879);
nor U1129 (N_1129,N_967,N_17);
or U1130 (N_1130,N_795,N_105);
nand U1131 (N_1131,N_74,N_472);
or U1132 (N_1132,N_324,N_326);
or U1133 (N_1133,N_475,N_60);
or U1134 (N_1134,N_906,N_491);
or U1135 (N_1135,N_942,N_511);
and U1136 (N_1136,N_740,N_235);
nand U1137 (N_1137,N_6,N_131);
nand U1138 (N_1138,N_207,N_78);
nor U1139 (N_1139,N_688,N_504);
nor U1140 (N_1140,N_189,N_206);
or U1141 (N_1141,N_809,N_892);
or U1142 (N_1142,N_550,N_676);
and U1143 (N_1143,N_88,N_690);
and U1144 (N_1144,N_668,N_670);
and U1145 (N_1145,N_391,N_138);
nor U1146 (N_1146,N_368,N_20);
nand U1147 (N_1147,N_935,N_8);
or U1148 (N_1148,N_185,N_280);
nand U1149 (N_1149,N_79,N_976);
and U1150 (N_1150,N_149,N_171);
or U1151 (N_1151,N_922,N_917);
nand U1152 (N_1152,N_909,N_144);
or U1153 (N_1153,N_620,N_941);
nand U1154 (N_1154,N_612,N_546);
nand U1155 (N_1155,N_30,N_981);
and U1156 (N_1156,N_992,N_464);
or U1157 (N_1157,N_653,N_423);
or U1158 (N_1158,N_485,N_39);
or U1159 (N_1159,N_520,N_698);
nand U1160 (N_1160,N_474,N_998);
and U1161 (N_1161,N_27,N_457);
nor U1162 (N_1162,N_339,N_605);
nor U1163 (N_1163,N_730,N_441);
and U1164 (N_1164,N_94,N_112);
nor U1165 (N_1165,N_335,N_376);
and U1166 (N_1166,N_719,N_506);
nand U1167 (N_1167,N_191,N_516);
nand U1168 (N_1168,N_515,N_15);
nor U1169 (N_1169,N_251,N_547);
nor U1170 (N_1170,N_915,N_452);
or U1171 (N_1171,N_267,N_203);
nand U1172 (N_1172,N_673,N_694);
or U1173 (N_1173,N_72,N_230);
and U1174 (N_1174,N_564,N_752);
nor U1175 (N_1175,N_264,N_736);
or U1176 (N_1176,N_931,N_463);
and U1177 (N_1177,N_359,N_855);
xor U1178 (N_1178,N_395,N_529);
nand U1179 (N_1179,N_828,N_924);
or U1180 (N_1180,N_345,N_63);
nand U1181 (N_1181,N_224,N_342);
nor U1182 (N_1182,N_632,N_346);
or U1183 (N_1183,N_782,N_677);
nand U1184 (N_1184,N_575,N_701);
nand U1185 (N_1185,N_542,N_603);
nand U1186 (N_1186,N_852,N_84);
and U1187 (N_1187,N_286,N_28);
and U1188 (N_1188,N_54,N_934);
or U1189 (N_1189,N_313,N_284);
xnor U1190 (N_1190,N_69,N_290);
and U1191 (N_1191,N_951,N_29);
nand U1192 (N_1192,N_252,N_530);
nor U1193 (N_1193,N_748,N_597);
and U1194 (N_1194,N_23,N_658);
and U1195 (N_1195,N_538,N_574);
nand U1196 (N_1196,N_785,N_396);
nor U1197 (N_1197,N_302,N_587);
or U1198 (N_1198,N_431,N_989);
nand U1199 (N_1199,N_993,N_916);
nor U1200 (N_1200,N_950,N_751);
nand U1201 (N_1201,N_675,N_71);
or U1202 (N_1202,N_797,N_95);
and U1203 (N_1203,N_738,N_938);
or U1204 (N_1204,N_321,N_622);
xnor U1205 (N_1205,N_873,N_732);
xnor U1206 (N_1206,N_503,N_292);
or U1207 (N_1207,N_860,N_250);
nand U1208 (N_1208,N_825,N_907);
xor U1209 (N_1209,N_727,N_133);
nand U1210 (N_1210,N_124,N_763);
xnor U1211 (N_1211,N_836,N_323);
and U1212 (N_1212,N_621,N_213);
or U1213 (N_1213,N_70,N_446);
or U1214 (N_1214,N_322,N_218);
nand U1215 (N_1215,N_101,N_194);
xnor U1216 (N_1216,N_401,N_205);
nand U1217 (N_1217,N_704,N_896);
nand U1218 (N_1218,N_308,N_103);
nor U1219 (N_1219,N_222,N_705);
nand U1220 (N_1220,N_999,N_669);
and U1221 (N_1221,N_710,N_367);
nand U1222 (N_1222,N_343,N_616);
and U1223 (N_1223,N_181,N_996);
or U1224 (N_1224,N_229,N_383);
nor U1225 (N_1225,N_269,N_192);
and U1226 (N_1226,N_919,N_780);
and U1227 (N_1227,N_429,N_380);
and U1228 (N_1228,N_527,N_588);
and U1229 (N_1229,N_180,N_744);
or U1230 (N_1230,N_581,N_971);
nand U1231 (N_1231,N_182,N_958);
nand U1232 (N_1232,N_533,N_91);
and U1233 (N_1233,N_589,N_611);
or U1234 (N_1234,N_900,N_747);
and U1235 (N_1235,N_121,N_271);
or U1236 (N_1236,N_361,N_476);
nor U1237 (N_1237,N_646,N_878);
nor U1238 (N_1238,N_585,N_193);
or U1239 (N_1239,N_398,N_435);
xor U1240 (N_1240,N_561,N_334);
and U1241 (N_1241,N_758,N_430);
nand U1242 (N_1242,N_273,N_256);
nand U1243 (N_1243,N_377,N_921);
and U1244 (N_1244,N_424,N_314);
nand U1245 (N_1245,N_394,N_173);
or U1246 (N_1246,N_248,N_984);
or U1247 (N_1247,N_382,N_661);
or U1248 (N_1248,N_988,N_162);
or U1249 (N_1249,N_184,N_211);
nor U1250 (N_1250,N_806,N_813);
nor U1251 (N_1251,N_99,N_568);
nor U1252 (N_1252,N_553,N_215);
or U1253 (N_1253,N_949,N_447);
nand U1254 (N_1254,N_918,N_283);
or U1255 (N_1255,N_437,N_139);
and U1256 (N_1256,N_643,N_590);
nand U1257 (N_1257,N_824,N_525);
or U1258 (N_1258,N_887,N_9);
or U1259 (N_1259,N_693,N_249);
nand U1260 (N_1260,N_56,N_68);
nand U1261 (N_1261,N_130,N_412);
and U1262 (N_1262,N_49,N_957);
and U1263 (N_1263,N_920,N_666);
or U1264 (N_1264,N_35,N_496);
or U1265 (N_1265,N_609,N_925);
and U1266 (N_1266,N_47,N_208);
nand U1267 (N_1267,N_707,N_776);
or U1268 (N_1268,N_883,N_477);
and U1269 (N_1269,N_948,N_462);
nor U1270 (N_1270,N_895,N_381);
nand U1271 (N_1271,N_154,N_619);
nand U1272 (N_1272,N_874,N_169);
nor U1273 (N_1273,N_210,N_869);
nor U1274 (N_1274,N_11,N_397);
and U1275 (N_1275,N_991,N_762);
nand U1276 (N_1276,N_389,N_839);
or U1277 (N_1277,N_309,N_295);
or U1278 (N_1278,N_45,N_787);
nand U1279 (N_1279,N_667,N_624);
nand U1280 (N_1280,N_937,N_521);
nor U1281 (N_1281,N_253,N_287);
or U1282 (N_1282,N_348,N_146);
and U1283 (N_1283,N_859,N_510);
and U1284 (N_1284,N_861,N_331);
nor U1285 (N_1285,N_982,N_445);
and U1286 (N_1286,N_681,N_387);
or U1287 (N_1287,N_628,N_537);
nand U1288 (N_1288,N_847,N_43);
nand U1289 (N_1289,N_456,N_195);
and U1290 (N_1290,N_128,N_317);
nand U1291 (N_1291,N_234,N_279);
and U1292 (N_1292,N_414,N_36);
or U1293 (N_1293,N_548,N_627);
or U1294 (N_1294,N_913,N_686);
nor U1295 (N_1295,N_630,N_233);
and U1296 (N_1296,N_92,N_582);
nor U1297 (N_1297,N_303,N_304);
or U1298 (N_1298,N_40,N_266);
and U1299 (N_1299,N_327,N_200);
nand U1300 (N_1300,N_3,N_330);
nand U1301 (N_1301,N_125,N_706);
nand U1302 (N_1302,N_202,N_278);
and U1303 (N_1303,N_850,N_720);
and U1304 (N_1304,N_642,N_466);
xor U1305 (N_1305,N_725,N_388);
nor U1306 (N_1306,N_932,N_204);
or U1307 (N_1307,N_403,N_583);
or U1308 (N_1308,N_888,N_148);
and U1309 (N_1309,N_32,N_344);
xor U1310 (N_1310,N_220,N_427);
xor U1311 (N_1311,N_14,N_576);
nand U1312 (N_1312,N_927,N_928);
nand U1313 (N_1313,N_818,N_237);
and U1314 (N_1314,N_379,N_779);
or U1315 (N_1315,N_882,N_305);
nand U1316 (N_1316,N_578,N_607);
or U1317 (N_1317,N_432,N_801);
and U1318 (N_1318,N_939,N_498);
or U1319 (N_1319,N_288,N_315);
and U1320 (N_1320,N_512,N_89);
or U1321 (N_1321,N_904,N_7);
nand U1322 (N_1322,N_13,N_363);
nand U1323 (N_1323,N_319,N_539);
nor U1324 (N_1324,N_332,N_788);
nor U1325 (N_1325,N_341,N_514);
or U1326 (N_1326,N_856,N_952);
or U1327 (N_1327,N_274,N_297);
nor U1328 (N_1328,N_970,N_483);
nor U1329 (N_1329,N_411,N_366);
nand U1330 (N_1330,N_557,N_413);
and U1331 (N_1331,N_800,N_268);
or U1332 (N_1332,N_34,N_699);
nand U1333 (N_1333,N_306,N_728);
nor U1334 (N_1334,N_910,N_245);
or U1335 (N_1335,N_77,N_277);
nand U1336 (N_1336,N_109,N_807);
or U1337 (N_1337,N_929,N_774);
or U1338 (N_1338,N_337,N_783);
nor U1339 (N_1339,N_880,N_275);
or U1340 (N_1340,N_769,N_374);
or U1341 (N_1341,N_739,N_426);
or U1342 (N_1342,N_65,N_645);
nor U1343 (N_1343,N_618,N_159);
nor U1344 (N_1344,N_983,N_565);
nor U1345 (N_1345,N_471,N_750);
nor U1346 (N_1346,N_102,N_152);
nor U1347 (N_1347,N_978,N_62);
nor U1348 (N_1348,N_723,N_100);
nand U1349 (N_1349,N_132,N_247);
nor U1350 (N_1350,N_114,N_418);
and U1351 (N_1351,N_357,N_58);
nand U1352 (N_1352,N_480,N_490);
nand U1353 (N_1353,N_325,N_473);
nand U1354 (N_1354,N_5,N_238);
or U1355 (N_1355,N_353,N_59);
or U1356 (N_1356,N_953,N_827);
nor U1357 (N_1357,N_289,N_495);
or U1358 (N_1358,N_741,N_872);
nand U1359 (N_1359,N_299,N_404);
or U1360 (N_1360,N_419,N_866);
nor U1361 (N_1361,N_243,N_734);
or U1362 (N_1362,N_908,N_761);
and U1363 (N_1363,N_449,N_468);
nor U1364 (N_1364,N_637,N_493);
and U1365 (N_1365,N_680,N_402);
and U1366 (N_1366,N_716,N_766);
and U1367 (N_1367,N_409,N_2);
xor U1368 (N_1368,N_375,N_488);
and U1369 (N_1369,N_759,N_19);
nor U1370 (N_1370,N_802,N_641);
nand U1371 (N_1371,N_771,N_37);
or U1372 (N_1372,N_650,N_549);
or U1373 (N_1373,N_507,N_966);
nor U1374 (N_1374,N_936,N_494);
and U1375 (N_1375,N_198,N_333);
and U1376 (N_1376,N_110,N_454);
xor U1377 (N_1377,N_293,N_384);
xor U1378 (N_1378,N_652,N_685);
and U1379 (N_1379,N_55,N_815);
nand U1380 (N_1380,N_768,N_571);
nand U1381 (N_1381,N_231,N_254);
nor U1382 (N_1382,N_914,N_260);
nor U1383 (N_1383,N_899,N_157);
and U1384 (N_1384,N_400,N_522);
or U1385 (N_1385,N_96,N_947);
xor U1386 (N_1386,N_870,N_544);
or U1387 (N_1387,N_4,N_61);
xor U1388 (N_1388,N_551,N_891);
nand U1389 (N_1389,N_190,N_535);
and U1390 (N_1390,N_792,N_311);
xnor U1391 (N_1391,N_420,N_742);
or U1392 (N_1392,N_757,N_610);
nand U1393 (N_1393,N_726,N_156);
nor U1394 (N_1394,N_969,N_294);
and U1395 (N_1395,N_682,N_586);
or U1396 (N_1396,N_244,N_636);
nor U1397 (N_1397,N_528,N_518);
or U1398 (N_1398,N_902,N_242);
or U1399 (N_1399,N_117,N_959);
nor U1400 (N_1400,N_596,N_791);
nand U1401 (N_1401,N_819,N_118);
nand U1402 (N_1402,N_448,N_120);
and U1403 (N_1403,N_552,N_558);
and U1404 (N_1404,N_876,N_80);
nor U1405 (N_1405,N_392,N_717);
and U1406 (N_1406,N_434,N_745);
nand U1407 (N_1407,N_700,N_393);
nand U1408 (N_1408,N_122,N_580);
xnor U1409 (N_1409,N_696,N_508);
or U1410 (N_1410,N_804,N_674);
and U1411 (N_1411,N_799,N_980);
and U1412 (N_1412,N_784,N_241);
nor U1413 (N_1413,N_593,N_298);
and U1414 (N_1414,N_545,N_838);
nand U1415 (N_1415,N_664,N_10);
nand U1416 (N_1416,N_579,N_212);
or U1417 (N_1417,N_450,N_240);
and U1418 (N_1418,N_901,N_285);
nand U1419 (N_1419,N_166,N_328);
nand U1420 (N_1420,N_691,N_417);
nor U1421 (N_1421,N_453,N_390);
nor U1422 (N_1422,N_44,N_226);
nand U1423 (N_1423,N_640,N_844);
nor U1424 (N_1424,N_147,N_86);
nor U1425 (N_1425,N_408,N_352);
or U1426 (N_1426,N_470,N_764);
nand U1427 (N_1427,N_990,N_840);
nand U1428 (N_1428,N_623,N_75);
or U1429 (N_1429,N_722,N_893);
or U1430 (N_1430,N_543,N_659);
and U1431 (N_1431,N_18,N_107);
nor U1432 (N_1432,N_329,N_209);
nand U1433 (N_1433,N_731,N_789);
or U1434 (N_1434,N_829,N_790);
nand U1435 (N_1435,N_817,N_721);
and U1436 (N_1436,N_541,N_428);
or U1437 (N_1437,N_145,N_943);
nand U1438 (N_1438,N_656,N_153);
or U1439 (N_1439,N_655,N_566);
and U1440 (N_1440,N_985,N_176);
and U1441 (N_1441,N_436,N_755);
nor U1442 (N_1442,N_517,N_119);
nor U1443 (N_1443,N_38,N_765);
or U1444 (N_1444,N_835,N_12);
and U1445 (N_1445,N_849,N_626);
and U1446 (N_1446,N_831,N_911);
nor U1447 (N_1447,N_559,N_724);
or U1448 (N_1448,N_841,N_877);
nand U1449 (N_1449,N_570,N_90);
and U1450 (N_1450,N_954,N_246);
and U1451 (N_1451,N_772,N_179);
nand U1452 (N_1452,N_890,N_214);
nor U1453 (N_1453,N_994,N_336);
and U1454 (N_1454,N_33,N_502);
and U1455 (N_1455,N_805,N_629);
nor U1456 (N_1456,N_733,N_97);
xnor U1457 (N_1457,N_64,N_500);
nor U1458 (N_1458,N_625,N_113);
nand U1459 (N_1459,N_126,N_158);
or U1460 (N_1460,N_672,N_255);
or U1461 (N_1461,N_845,N_340);
nand U1462 (N_1462,N_573,N_196);
and U1463 (N_1463,N_760,N_83);
or U1464 (N_1464,N_168,N_796);
nand U1465 (N_1465,N_356,N_600);
and U1466 (N_1466,N_863,N_26);
nand U1467 (N_1467,N_46,N_964);
and U1468 (N_1468,N_320,N_955);
nand U1469 (N_1469,N_455,N_997);
and U1470 (N_1470,N_832,N_82);
nand U1471 (N_1471,N_385,N_714);
nor U1472 (N_1472,N_709,N_188);
and U1473 (N_1473,N_98,N_775);
nand U1474 (N_1474,N_66,N_81);
nand U1475 (N_1475,N_614,N_405);
nor U1476 (N_1476,N_373,N_591);
and U1477 (N_1477,N_465,N_865);
nand U1478 (N_1478,N_615,N_127);
nand U1479 (N_1479,N_160,N_737);
nand U1480 (N_1480,N_350,N_956);
or U1481 (N_1481,N_972,N_735);
nand U1482 (N_1482,N_316,N_167);
nand U1483 (N_1483,N_756,N_536);
nor U1484 (N_1484,N_170,N_613);
and U1485 (N_1485,N_451,N_365);
or U1486 (N_1486,N_134,N_875);
nand U1487 (N_1487,N_232,N_360);
or U1488 (N_1488,N_554,N_821);
and U1489 (N_1489,N_399,N_48);
and U1490 (N_1490,N_406,N_16);
xnor U1491 (N_1491,N_104,N_684);
or U1492 (N_1492,N_301,N_926);
nand U1493 (N_1493,N_638,N_524);
nor U1494 (N_1494,N_979,N_31);
nand U1495 (N_1495,N_599,N_310);
nand U1496 (N_1496,N_410,N_444);
or U1497 (N_1497,N_960,N_281);
nand U1498 (N_1498,N_372,N_155);
nor U1499 (N_1499,N_150,N_362);
or U1500 (N_1500,N_427,N_936);
and U1501 (N_1501,N_686,N_817);
nand U1502 (N_1502,N_585,N_347);
and U1503 (N_1503,N_955,N_493);
and U1504 (N_1504,N_558,N_913);
xor U1505 (N_1505,N_374,N_289);
and U1506 (N_1506,N_940,N_180);
nor U1507 (N_1507,N_445,N_527);
and U1508 (N_1508,N_240,N_293);
nand U1509 (N_1509,N_877,N_110);
nand U1510 (N_1510,N_884,N_930);
nand U1511 (N_1511,N_368,N_561);
nand U1512 (N_1512,N_732,N_273);
or U1513 (N_1513,N_168,N_5);
nand U1514 (N_1514,N_643,N_916);
or U1515 (N_1515,N_19,N_82);
and U1516 (N_1516,N_151,N_708);
or U1517 (N_1517,N_729,N_177);
nor U1518 (N_1518,N_413,N_126);
nor U1519 (N_1519,N_953,N_829);
xor U1520 (N_1520,N_89,N_326);
and U1521 (N_1521,N_960,N_647);
and U1522 (N_1522,N_16,N_453);
and U1523 (N_1523,N_603,N_115);
nand U1524 (N_1524,N_566,N_215);
or U1525 (N_1525,N_233,N_391);
nor U1526 (N_1526,N_237,N_644);
nor U1527 (N_1527,N_165,N_95);
xnor U1528 (N_1528,N_83,N_885);
and U1529 (N_1529,N_596,N_646);
or U1530 (N_1530,N_102,N_928);
or U1531 (N_1531,N_286,N_191);
or U1532 (N_1532,N_982,N_117);
xor U1533 (N_1533,N_496,N_412);
or U1534 (N_1534,N_778,N_5);
and U1535 (N_1535,N_337,N_439);
nor U1536 (N_1536,N_82,N_984);
nor U1537 (N_1537,N_430,N_884);
nor U1538 (N_1538,N_418,N_275);
nand U1539 (N_1539,N_481,N_783);
nor U1540 (N_1540,N_786,N_213);
nand U1541 (N_1541,N_21,N_448);
xnor U1542 (N_1542,N_632,N_581);
nand U1543 (N_1543,N_467,N_891);
nand U1544 (N_1544,N_510,N_542);
and U1545 (N_1545,N_729,N_235);
and U1546 (N_1546,N_332,N_196);
nand U1547 (N_1547,N_954,N_790);
or U1548 (N_1548,N_147,N_73);
and U1549 (N_1549,N_382,N_300);
or U1550 (N_1550,N_787,N_195);
xor U1551 (N_1551,N_472,N_943);
nor U1552 (N_1552,N_661,N_535);
nor U1553 (N_1553,N_304,N_714);
nand U1554 (N_1554,N_811,N_462);
and U1555 (N_1555,N_39,N_22);
nand U1556 (N_1556,N_170,N_11);
and U1557 (N_1557,N_305,N_531);
nand U1558 (N_1558,N_887,N_978);
or U1559 (N_1559,N_834,N_624);
nor U1560 (N_1560,N_33,N_161);
and U1561 (N_1561,N_289,N_58);
nand U1562 (N_1562,N_12,N_468);
nand U1563 (N_1563,N_646,N_210);
nand U1564 (N_1564,N_789,N_38);
nand U1565 (N_1565,N_162,N_769);
and U1566 (N_1566,N_452,N_541);
nor U1567 (N_1567,N_977,N_680);
nand U1568 (N_1568,N_831,N_110);
or U1569 (N_1569,N_846,N_836);
nand U1570 (N_1570,N_338,N_176);
nand U1571 (N_1571,N_255,N_884);
and U1572 (N_1572,N_660,N_236);
nand U1573 (N_1573,N_271,N_321);
or U1574 (N_1574,N_30,N_729);
and U1575 (N_1575,N_419,N_962);
nand U1576 (N_1576,N_957,N_146);
nand U1577 (N_1577,N_152,N_287);
xor U1578 (N_1578,N_717,N_138);
nand U1579 (N_1579,N_93,N_289);
nor U1580 (N_1580,N_899,N_150);
nand U1581 (N_1581,N_136,N_784);
or U1582 (N_1582,N_693,N_153);
nand U1583 (N_1583,N_493,N_878);
nor U1584 (N_1584,N_782,N_774);
or U1585 (N_1585,N_890,N_751);
nand U1586 (N_1586,N_187,N_194);
nor U1587 (N_1587,N_806,N_362);
nand U1588 (N_1588,N_282,N_800);
and U1589 (N_1589,N_25,N_562);
nand U1590 (N_1590,N_812,N_269);
nand U1591 (N_1591,N_31,N_321);
and U1592 (N_1592,N_959,N_221);
nor U1593 (N_1593,N_512,N_730);
nand U1594 (N_1594,N_726,N_964);
xor U1595 (N_1595,N_882,N_257);
or U1596 (N_1596,N_158,N_87);
nor U1597 (N_1597,N_846,N_333);
and U1598 (N_1598,N_332,N_480);
nand U1599 (N_1599,N_810,N_235);
nand U1600 (N_1600,N_35,N_964);
or U1601 (N_1601,N_863,N_817);
or U1602 (N_1602,N_658,N_757);
and U1603 (N_1603,N_918,N_161);
nand U1604 (N_1604,N_481,N_860);
nor U1605 (N_1605,N_277,N_35);
xnor U1606 (N_1606,N_777,N_469);
and U1607 (N_1607,N_496,N_612);
or U1608 (N_1608,N_346,N_289);
or U1609 (N_1609,N_321,N_546);
or U1610 (N_1610,N_840,N_266);
or U1611 (N_1611,N_919,N_157);
xnor U1612 (N_1612,N_262,N_764);
and U1613 (N_1613,N_441,N_194);
and U1614 (N_1614,N_807,N_748);
or U1615 (N_1615,N_466,N_885);
and U1616 (N_1616,N_623,N_889);
and U1617 (N_1617,N_802,N_475);
nor U1618 (N_1618,N_966,N_429);
nand U1619 (N_1619,N_164,N_624);
nor U1620 (N_1620,N_980,N_860);
and U1621 (N_1621,N_898,N_806);
or U1622 (N_1622,N_403,N_670);
nand U1623 (N_1623,N_896,N_352);
nand U1624 (N_1624,N_177,N_441);
and U1625 (N_1625,N_588,N_287);
and U1626 (N_1626,N_7,N_533);
and U1627 (N_1627,N_773,N_802);
or U1628 (N_1628,N_788,N_906);
and U1629 (N_1629,N_167,N_145);
and U1630 (N_1630,N_925,N_498);
nand U1631 (N_1631,N_662,N_659);
and U1632 (N_1632,N_552,N_56);
nand U1633 (N_1633,N_598,N_944);
nand U1634 (N_1634,N_243,N_92);
nand U1635 (N_1635,N_960,N_503);
or U1636 (N_1636,N_756,N_626);
nand U1637 (N_1637,N_548,N_43);
and U1638 (N_1638,N_953,N_799);
nand U1639 (N_1639,N_261,N_515);
or U1640 (N_1640,N_854,N_416);
and U1641 (N_1641,N_61,N_903);
xnor U1642 (N_1642,N_66,N_804);
and U1643 (N_1643,N_373,N_531);
nor U1644 (N_1644,N_778,N_135);
nor U1645 (N_1645,N_922,N_820);
nor U1646 (N_1646,N_860,N_936);
and U1647 (N_1647,N_921,N_597);
and U1648 (N_1648,N_664,N_972);
and U1649 (N_1649,N_610,N_765);
nand U1650 (N_1650,N_959,N_326);
or U1651 (N_1651,N_280,N_109);
nor U1652 (N_1652,N_140,N_112);
and U1653 (N_1653,N_738,N_541);
nor U1654 (N_1654,N_515,N_563);
and U1655 (N_1655,N_362,N_369);
nand U1656 (N_1656,N_970,N_404);
nor U1657 (N_1657,N_141,N_310);
and U1658 (N_1658,N_100,N_591);
nor U1659 (N_1659,N_751,N_112);
or U1660 (N_1660,N_664,N_8);
nand U1661 (N_1661,N_107,N_968);
xor U1662 (N_1662,N_388,N_959);
or U1663 (N_1663,N_40,N_134);
nand U1664 (N_1664,N_810,N_952);
nand U1665 (N_1665,N_182,N_778);
and U1666 (N_1666,N_600,N_349);
and U1667 (N_1667,N_257,N_635);
nand U1668 (N_1668,N_439,N_496);
and U1669 (N_1669,N_775,N_791);
nand U1670 (N_1670,N_628,N_732);
and U1671 (N_1671,N_674,N_324);
and U1672 (N_1672,N_401,N_202);
nand U1673 (N_1673,N_48,N_419);
nor U1674 (N_1674,N_19,N_918);
nand U1675 (N_1675,N_657,N_434);
and U1676 (N_1676,N_33,N_879);
or U1677 (N_1677,N_732,N_4);
nand U1678 (N_1678,N_191,N_335);
and U1679 (N_1679,N_15,N_135);
or U1680 (N_1680,N_617,N_147);
or U1681 (N_1681,N_57,N_820);
nor U1682 (N_1682,N_946,N_285);
and U1683 (N_1683,N_404,N_142);
nor U1684 (N_1684,N_247,N_413);
xnor U1685 (N_1685,N_856,N_302);
or U1686 (N_1686,N_982,N_417);
nor U1687 (N_1687,N_729,N_377);
xnor U1688 (N_1688,N_566,N_945);
nor U1689 (N_1689,N_20,N_437);
and U1690 (N_1690,N_171,N_408);
and U1691 (N_1691,N_1,N_350);
nor U1692 (N_1692,N_900,N_421);
nand U1693 (N_1693,N_374,N_719);
nor U1694 (N_1694,N_662,N_178);
nand U1695 (N_1695,N_235,N_764);
nand U1696 (N_1696,N_145,N_272);
and U1697 (N_1697,N_628,N_892);
or U1698 (N_1698,N_971,N_547);
nor U1699 (N_1699,N_758,N_914);
or U1700 (N_1700,N_415,N_728);
and U1701 (N_1701,N_634,N_228);
or U1702 (N_1702,N_205,N_999);
and U1703 (N_1703,N_218,N_458);
or U1704 (N_1704,N_93,N_433);
nand U1705 (N_1705,N_71,N_841);
and U1706 (N_1706,N_567,N_445);
nor U1707 (N_1707,N_617,N_78);
nor U1708 (N_1708,N_322,N_991);
and U1709 (N_1709,N_920,N_54);
and U1710 (N_1710,N_771,N_411);
nor U1711 (N_1711,N_857,N_140);
nor U1712 (N_1712,N_341,N_633);
and U1713 (N_1713,N_527,N_477);
and U1714 (N_1714,N_14,N_183);
nand U1715 (N_1715,N_920,N_182);
or U1716 (N_1716,N_545,N_222);
or U1717 (N_1717,N_490,N_576);
or U1718 (N_1718,N_133,N_541);
and U1719 (N_1719,N_57,N_843);
nand U1720 (N_1720,N_478,N_169);
and U1721 (N_1721,N_396,N_370);
or U1722 (N_1722,N_465,N_666);
or U1723 (N_1723,N_956,N_183);
nand U1724 (N_1724,N_365,N_699);
nand U1725 (N_1725,N_448,N_505);
and U1726 (N_1726,N_9,N_728);
nand U1727 (N_1727,N_439,N_109);
nor U1728 (N_1728,N_225,N_502);
and U1729 (N_1729,N_603,N_130);
and U1730 (N_1730,N_209,N_135);
nor U1731 (N_1731,N_614,N_561);
and U1732 (N_1732,N_915,N_895);
nand U1733 (N_1733,N_561,N_362);
or U1734 (N_1734,N_672,N_985);
and U1735 (N_1735,N_394,N_956);
and U1736 (N_1736,N_305,N_283);
nand U1737 (N_1737,N_7,N_199);
and U1738 (N_1738,N_784,N_504);
nor U1739 (N_1739,N_673,N_442);
nand U1740 (N_1740,N_49,N_761);
or U1741 (N_1741,N_413,N_851);
or U1742 (N_1742,N_989,N_451);
nor U1743 (N_1743,N_805,N_748);
and U1744 (N_1744,N_262,N_131);
nand U1745 (N_1745,N_422,N_415);
and U1746 (N_1746,N_638,N_533);
nor U1747 (N_1747,N_560,N_146);
nand U1748 (N_1748,N_767,N_837);
nor U1749 (N_1749,N_641,N_884);
nand U1750 (N_1750,N_555,N_759);
nor U1751 (N_1751,N_193,N_983);
and U1752 (N_1752,N_38,N_790);
nor U1753 (N_1753,N_677,N_70);
or U1754 (N_1754,N_943,N_113);
nand U1755 (N_1755,N_948,N_424);
nand U1756 (N_1756,N_553,N_587);
nor U1757 (N_1757,N_519,N_638);
nand U1758 (N_1758,N_780,N_842);
nor U1759 (N_1759,N_876,N_252);
or U1760 (N_1760,N_424,N_178);
nand U1761 (N_1761,N_107,N_791);
nor U1762 (N_1762,N_978,N_236);
xnor U1763 (N_1763,N_892,N_177);
xor U1764 (N_1764,N_656,N_387);
and U1765 (N_1765,N_459,N_599);
nand U1766 (N_1766,N_89,N_409);
nor U1767 (N_1767,N_358,N_782);
or U1768 (N_1768,N_461,N_489);
nor U1769 (N_1769,N_467,N_850);
nand U1770 (N_1770,N_187,N_434);
and U1771 (N_1771,N_781,N_762);
or U1772 (N_1772,N_234,N_567);
nor U1773 (N_1773,N_1,N_8);
or U1774 (N_1774,N_369,N_562);
nor U1775 (N_1775,N_158,N_845);
and U1776 (N_1776,N_7,N_166);
nand U1777 (N_1777,N_971,N_12);
or U1778 (N_1778,N_843,N_13);
nand U1779 (N_1779,N_409,N_946);
or U1780 (N_1780,N_979,N_310);
nor U1781 (N_1781,N_45,N_463);
and U1782 (N_1782,N_858,N_910);
or U1783 (N_1783,N_937,N_526);
nand U1784 (N_1784,N_334,N_420);
and U1785 (N_1785,N_930,N_844);
or U1786 (N_1786,N_256,N_277);
or U1787 (N_1787,N_959,N_717);
nor U1788 (N_1788,N_59,N_678);
and U1789 (N_1789,N_480,N_402);
or U1790 (N_1790,N_888,N_126);
nor U1791 (N_1791,N_169,N_743);
nand U1792 (N_1792,N_602,N_969);
and U1793 (N_1793,N_764,N_453);
or U1794 (N_1794,N_217,N_896);
nor U1795 (N_1795,N_499,N_762);
nor U1796 (N_1796,N_829,N_35);
or U1797 (N_1797,N_502,N_664);
nor U1798 (N_1798,N_824,N_937);
and U1799 (N_1799,N_861,N_249);
or U1800 (N_1800,N_263,N_60);
nand U1801 (N_1801,N_727,N_316);
or U1802 (N_1802,N_133,N_977);
and U1803 (N_1803,N_970,N_790);
nand U1804 (N_1804,N_955,N_615);
or U1805 (N_1805,N_135,N_265);
nor U1806 (N_1806,N_128,N_279);
nand U1807 (N_1807,N_468,N_370);
nor U1808 (N_1808,N_896,N_677);
and U1809 (N_1809,N_379,N_744);
and U1810 (N_1810,N_282,N_211);
xor U1811 (N_1811,N_978,N_385);
xnor U1812 (N_1812,N_243,N_180);
nand U1813 (N_1813,N_372,N_117);
and U1814 (N_1814,N_727,N_382);
nand U1815 (N_1815,N_364,N_278);
or U1816 (N_1816,N_910,N_576);
or U1817 (N_1817,N_993,N_30);
nor U1818 (N_1818,N_755,N_650);
and U1819 (N_1819,N_206,N_413);
and U1820 (N_1820,N_313,N_846);
and U1821 (N_1821,N_354,N_463);
nor U1822 (N_1822,N_811,N_133);
or U1823 (N_1823,N_751,N_400);
nor U1824 (N_1824,N_983,N_820);
and U1825 (N_1825,N_179,N_135);
or U1826 (N_1826,N_759,N_296);
and U1827 (N_1827,N_208,N_333);
or U1828 (N_1828,N_546,N_335);
and U1829 (N_1829,N_221,N_715);
nor U1830 (N_1830,N_358,N_249);
or U1831 (N_1831,N_704,N_135);
nand U1832 (N_1832,N_495,N_376);
nor U1833 (N_1833,N_333,N_201);
nand U1834 (N_1834,N_0,N_111);
nor U1835 (N_1835,N_448,N_777);
and U1836 (N_1836,N_444,N_766);
and U1837 (N_1837,N_502,N_380);
and U1838 (N_1838,N_749,N_886);
nor U1839 (N_1839,N_658,N_834);
and U1840 (N_1840,N_953,N_966);
and U1841 (N_1841,N_12,N_814);
and U1842 (N_1842,N_525,N_250);
nand U1843 (N_1843,N_58,N_906);
nand U1844 (N_1844,N_323,N_636);
or U1845 (N_1845,N_333,N_959);
or U1846 (N_1846,N_300,N_928);
nor U1847 (N_1847,N_609,N_995);
nor U1848 (N_1848,N_479,N_937);
nand U1849 (N_1849,N_751,N_495);
nor U1850 (N_1850,N_167,N_866);
or U1851 (N_1851,N_825,N_978);
or U1852 (N_1852,N_439,N_434);
and U1853 (N_1853,N_948,N_742);
nor U1854 (N_1854,N_880,N_674);
and U1855 (N_1855,N_704,N_795);
or U1856 (N_1856,N_273,N_21);
and U1857 (N_1857,N_11,N_987);
nand U1858 (N_1858,N_699,N_846);
and U1859 (N_1859,N_389,N_328);
xnor U1860 (N_1860,N_342,N_588);
or U1861 (N_1861,N_279,N_9);
nand U1862 (N_1862,N_237,N_991);
or U1863 (N_1863,N_817,N_236);
and U1864 (N_1864,N_339,N_276);
nand U1865 (N_1865,N_659,N_740);
and U1866 (N_1866,N_270,N_396);
and U1867 (N_1867,N_741,N_959);
and U1868 (N_1868,N_636,N_846);
and U1869 (N_1869,N_903,N_860);
xor U1870 (N_1870,N_326,N_358);
or U1871 (N_1871,N_833,N_82);
and U1872 (N_1872,N_128,N_65);
nand U1873 (N_1873,N_397,N_659);
and U1874 (N_1874,N_445,N_77);
nor U1875 (N_1875,N_415,N_892);
nor U1876 (N_1876,N_271,N_642);
nor U1877 (N_1877,N_268,N_607);
and U1878 (N_1878,N_116,N_832);
nor U1879 (N_1879,N_356,N_984);
or U1880 (N_1880,N_234,N_626);
nand U1881 (N_1881,N_909,N_377);
or U1882 (N_1882,N_381,N_761);
nor U1883 (N_1883,N_735,N_386);
and U1884 (N_1884,N_75,N_484);
nand U1885 (N_1885,N_950,N_891);
xnor U1886 (N_1886,N_791,N_513);
or U1887 (N_1887,N_174,N_547);
nor U1888 (N_1888,N_339,N_674);
nor U1889 (N_1889,N_246,N_874);
nand U1890 (N_1890,N_692,N_675);
nand U1891 (N_1891,N_131,N_340);
nor U1892 (N_1892,N_630,N_168);
nor U1893 (N_1893,N_370,N_559);
or U1894 (N_1894,N_481,N_292);
and U1895 (N_1895,N_475,N_438);
nand U1896 (N_1896,N_492,N_798);
and U1897 (N_1897,N_881,N_687);
and U1898 (N_1898,N_143,N_284);
nor U1899 (N_1899,N_307,N_312);
nand U1900 (N_1900,N_907,N_524);
nand U1901 (N_1901,N_571,N_696);
nor U1902 (N_1902,N_728,N_228);
and U1903 (N_1903,N_551,N_982);
nand U1904 (N_1904,N_505,N_282);
or U1905 (N_1905,N_89,N_734);
or U1906 (N_1906,N_641,N_488);
nor U1907 (N_1907,N_506,N_187);
and U1908 (N_1908,N_202,N_930);
nand U1909 (N_1909,N_940,N_842);
nand U1910 (N_1910,N_394,N_242);
or U1911 (N_1911,N_641,N_303);
nor U1912 (N_1912,N_827,N_583);
xor U1913 (N_1913,N_780,N_442);
or U1914 (N_1914,N_463,N_108);
or U1915 (N_1915,N_453,N_75);
or U1916 (N_1916,N_508,N_352);
or U1917 (N_1917,N_108,N_335);
or U1918 (N_1918,N_946,N_835);
and U1919 (N_1919,N_88,N_327);
nand U1920 (N_1920,N_942,N_460);
nand U1921 (N_1921,N_60,N_865);
nor U1922 (N_1922,N_780,N_713);
nand U1923 (N_1923,N_852,N_533);
or U1924 (N_1924,N_339,N_176);
nand U1925 (N_1925,N_703,N_666);
or U1926 (N_1926,N_567,N_75);
nor U1927 (N_1927,N_268,N_78);
nor U1928 (N_1928,N_632,N_542);
and U1929 (N_1929,N_112,N_883);
nand U1930 (N_1930,N_394,N_759);
and U1931 (N_1931,N_376,N_721);
nand U1932 (N_1932,N_720,N_781);
and U1933 (N_1933,N_112,N_172);
nor U1934 (N_1934,N_574,N_198);
nand U1935 (N_1935,N_145,N_927);
and U1936 (N_1936,N_155,N_109);
and U1937 (N_1937,N_382,N_713);
and U1938 (N_1938,N_248,N_145);
nor U1939 (N_1939,N_868,N_446);
nand U1940 (N_1940,N_800,N_649);
or U1941 (N_1941,N_806,N_785);
xor U1942 (N_1942,N_551,N_230);
and U1943 (N_1943,N_594,N_931);
and U1944 (N_1944,N_820,N_568);
and U1945 (N_1945,N_362,N_179);
nand U1946 (N_1946,N_922,N_791);
or U1947 (N_1947,N_529,N_750);
nand U1948 (N_1948,N_752,N_283);
xnor U1949 (N_1949,N_778,N_240);
nand U1950 (N_1950,N_14,N_682);
and U1951 (N_1951,N_541,N_534);
or U1952 (N_1952,N_228,N_953);
or U1953 (N_1953,N_377,N_929);
nand U1954 (N_1954,N_701,N_938);
or U1955 (N_1955,N_649,N_741);
nand U1956 (N_1956,N_735,N_776);
or U1957 (N_1957,N_281,N_536);
and U1958 (N_1958,N_111,N_848);
nand U1959 (N_1959,N_443,N_679);
nand U1960 (N_1960,N_990,N_111);
and U1961 (N_1961,N_451,N_995);
or U1962 (N_1962,N_271,N_730);
nor U1963 (N_1963,N_159,N_379);
nand U1964 (N_1964,N_875,N_318);
and U1965 (N_1965,N_586,N_614);
and U1966 (N_1966,N_380,N_716);
and U1967 (N_1967,N_811,N_663);
or U1968 (N_1968,N_980,N_570);
and U1969 (N_1969,N_425,N_69);
xor U1970 (N_1970,N_383,N_238);
or U1971 (N_1971,N_942,N_655);
and U1972 (N_1972,N_650,N_986);
or U1973 (N_1973,N_83,N_92);
nand U1974 (N_1974,N_917,N_61);
nor U1975 (N_1975,N_808,N_733);
nor U1976 (N_1976,N_171,N_872);
nor U1977 (N_1977,N_24,N_705);
and U1978 (N_1978,N_982,N_81);
and U1979 (N_1979,N_364,N_857);
nor U1980 (N_1980,N_932,N_289);
or U1981 (N_1981,N_436,N_182);
nor U1982 (N_1982,N_598,N_850);
nor U1983 (N_1983,N_878,N_185);
and U1984 (N_1984,N_617,N_910);
nor U1985 (N_1985,N_619,N_460);
or U1986 (N_1986,N_911,N_439);
or U1987 (N_1987,N_303,N_418);
and U1988 (N_1988,N_161,N_694);
nor U1989 (N_1989,N_579,N_445);
and U1990 (N_1990,N_604,N_6);
and U1991 (N_1991,N_242,N_481);
nand U1992 (N_1992,N_529,N_992);
nand U1993 (N_1993,N_755,N_35);
nor U1994 (N_1994,N_380,N_401);
nor U1995 (N_1995,N_69,N_442);
and U1996 (N_1996,N_153,N_657);
nor U1997 (N_1997,N_994,N_835);
nand U1998 (N_1998,N_94,N_363);
or U1999 (N_1999,N_410,N_705);
nand U2000 (N_2000,N_1061,N_1633);
and U2001 (N_2001,N_1110,N_1941);
nand U2002 (N_2002,N_1226,N_1240);
or U2003 (N_2003,N_1290,N_1643);
or U2004 (N_2004,N_1391,N_1315);
nand U2005 (N_2005,N_1943,N_1053);
and U2006 (N_2006,N_1779,N_1004);
nor U2007 (N_2007,N_1371,N_1994);
nor U2008 (N_2008,N_1449,N_1539);
or U2009 (N_2009,N_1854,N_1613);
nand U2010 (N_2010,N_1585,N_1015);
nand U2011 (N_2011,N_1795,N_1051);
xnor U2012 (N_2012,N_1114,N_1563);
nor U2013 (N_2013,N_1988,N_1363);
or U2014 (N_2014,N_1626,N_1444);
nor U2015 (N_2015,N_1178,N_1870);
or U2016 (N_2016,N_1509,N_1582);
nand U2017 (N_2017,N_1171,N_1274);
or U2018 (N_2018,N_1596,N_1491);
or U2019 (N_2019,N_1791,N_1901);
and U2020 (N_2020,N_1070,N_1561);
and U2021 (N_2021,N_1484,N_1165);
nand U2022 (N_2022,N_1570,N_1669);
nor U2023 (N_2023,N_1587,N_1798);
xor U2024 (N_2024,N_1551,N_1929);
or U2025 (N_2025,N_1604,N_1326);
and U2026 (N_2026,N_1193,N_1662);
or U2027 (N_2027,N_1856,N_1222);
and U2028 (N_2028,N_1523,N_1871);
and U2029 (N_2029,N_1574,N_1461);
nand U2030 (N_2030,N_1517,N_1223);
or U2031 (N_2031,N_1900,N_1298);
nor U2032 (N_2032,N_1269,N_1725);
or U2033 (N_2033,N_1914,N_1873);
and U2034 (N_2034,N_1378,N_1620);
nand U2035 (N_2035,N_1147,N_1595);
or U2036 (N_2036,N_1323,N_1243);
nand U2037 (N_2037,N_1097,N_1251);
nor U2038 (N_2038,N_1899,N_1977);
nand U2039 (N_2039,N_1266,N_1438);
and U2040 (N_2040,N_1526,N_1804);
nand U2041 (N_2041,N_1212,N_1228);
nor U2042 (N_2042,N_1621,N_1191);
nor U2043 (N_2043,N_1064,N_1541);
nand U2044 (N_2044,N_1842,N_1992);
and U2045 (N_2045,N_1625,N_1005);
or U2046 (N_2046,N_1122,N_1489);
nor U2047 (N_2047,N_1336,N_1978);
nor U2048 (N_2048,N_1105,N_1826);
and U2049 (N_2049,N_1088,N_1289);
and U2050 (N_2050,N_1908,N_1014);
nand U2051 (N_2051,N_1384,N_1263);
and U2052 (N_2052,N_1395,N_1163);
or U2053 (N_2053,N_1698,N_1809);
and U2054 (N_2054,N_1537,N_1608);
nand U2055 (N_2055,N_1867,N_1667);
nor U2056 (N_2056,N_1514,N_1916);
nor U2057 (N_2057,N_1721,N_1982);
nor U2058 (N_2058,N_1880,N_1696);
nor U2059 (N_2059,N_1821,N_1155);
or U2060 (N_2060,N_1360,N_1749);
or U2061 (N_2061,N_1600,N_1174);
nor U2062 (N_2062,N_1388,N_1717);
nor U2063 (N_2063,N_1383,N_1035);
nor U2064 (N_2064,N_1262,N_1028);
or U2065 (N_2065,N_1022,N_1271);
nor U2066 (N_2066,N_1258,N_1907);
or U2067 (N_2067,N_1960,N_1961);
or U2068 (N_2068,N_1148,N_1018);
nand U2069 (N_2069,N_1709,N_1134);
or U2070 (N_2070,N_1328,N_1065);
nor U2071 (N_2071,N_1936,N_1543);
or U2072 (N_2072,N_1707,N_1670);
or U2073 (N_2073,N_1758,N_1934);
nand U2074 (N_2074,N_1536,N_1851);
nor U2075 (N_2075,N_1353,N_1957);
or U2076 (N_2076,N_1632,N_1349);
or U2077 (N_2077,N_1589,N_1132);
or U2078 (N_2078,N_1091,N_1457);
and U2079 (N_2079,N_1882,N_1970);
nand U2080 (N_2080,N_1149,N_1739);
nand U2081 (N_2081,N_1843,N_1127);
nor U2082 (N_2082,N_1689,N_1664);
nand U2083 (N_2083,N_1614,N_1676);
or U2084 (N_2084,N_1468,N_1953);
nand U2085 (N_2085,N_1711,N_1179);
nor U2086 (N_2086,N_1233,N_1265);
or U2087 (N_2087,N_1547,N_1708);
nor U2088 (N_2088,N_1838,N_1902);
nor U2089 (N_2089,N_1682,N_1442);
and U2090 (N_2090,N_1086,N_1277);
nor U2091 (N_2091,N_1974,N_1690);
nand U2092 (N_2092,N_1488,N_1525);
xnor U2093 (N_2093,N_1412,N_1590);
nor U2094 (N_2094,N_1032,N_1405);
or U2095 (N_2095,N_1074,N_1607);
nand U2096 (N_2096,N_1466,N_1714);
nor U2097 (N_2097,N_1622,N_1888);
nor U2098 (N_2098,N_1511,N_1441);
or U2099 (N_2099,N_1087,N_1630);
and U2100 (N_2100,N_1747,N_1469);
nor U2101 (N_2101,N_1531,N_1048);
nor U2102 (N_2102,N_1783,N_1672);
and U2103 (N_2103,N_1432,N_1577);
or U2104 (N_2104,N_1121,N_1242);
or U2105 (N_2105,N_1403,N_1860);
and U2106 (N_2106,N_1340,N_1325);
or U2107 (N_2107,N_1636,N_1093);
nor U2108 (N_2108,N_1557,N_1701);
and U2109 (N_2109,N_1638,N_1656);
nor U2110 (N_2110,N_1849,N_1055);
nor U2111 (N_2111,N_1748,N_1231);
nand U2112 (N_2112,N_1910,N_1092);
or U2113 (N_2113,N_1423,N_1275);
nand U2114 (N_2114,N_1117,N_1524);
and U2115 (N_2115,N_1955,N_1320);
nand U2116 (N_2116,N_1026,N_1213);
nand U2117 (N_2117,N_1245,N_1085);
or U2118 (N_2118,N_1877,N_1562);
or U2119 (N_2119,N_1344,N_1164);
nor U2120 (N_2120,N_1396,N_1575);
or U2121 (N_2121,N_1131,N_1244);
nand U2122 (N_2122,N_1042,N_1218);
nor U2123 (N_2123,N_1678,N_1368);
nand U2124 (N_2124,N_1780,N_1508);
and U2125 (N_2125,N_1790,N_1406);
nand U2126 (N_2126,N_1852,N_1774);
or U2127 (N_2127,N_1715,N_1935);
and U2128 (N_2128,N_1654,N_1499);
and U2129 (N_2129,N_1306,N_1834);
nor U2130 (N_2130,N_1544,N_1528);
nor U2131 (N_2131,N_1822,N_1685);
or U2132 (N_2132,N_1675,N_1199);
or U2133 (N_2133,N_1983,N_1576);
nor U2134 (N_2134,N_1189,N_1844);
nor U2135 (N_2135,N_1335,N_1972);
nor U2136 (N_2136,N_1920,N_1981);
and U2137 (N_2137,N_1422,N_1505);
nor U2138 (N_2138,N_1366,N_1000);
nand U2139 (N_2139,N_1002,N_1694);
nor U2140 (N_2140,N_1776,N_1280);
nor U2141 (N_2141,N_1080,N_1476);
and U2142 (N_2142,N_1592,N_1765);
and U2143 (N_2143,N_1940,N_1376);
nor U2144 (N_2144,N_1796,N_1426);
xnor U2145 (N_2145,N_1173,N_1470);
nand U2146 (N_2146,N_1175,N_1415);
nand U2147 (N_2147,N_1889,N_1425);
nor U2148 (N_2148,N_1635,N_1357);
or U2149 (N_2149,N_1788,N_1845);
nor U2150 (N_2150,N_1052,N_1706);
or U2151 (N_2151,N_1285,N_1818);
or U2152 (N_2152,N_1201,N_1886);
or U2153 (N_2153,N_1309,N_1753);
nor U2154 (N_2154,N_1374,N_1713);
nand U2155 (N_2155,N_1408,N_1658);
nor U2156 (N_2156,N_1247,N_1639);
xnor U2157 (N_2157,N_1008,N_1593);
and U2158 (N_2158,N_1436,N_1400);
nand U2159 (N_2159,N_1581,N_1996);
and U2160 (N_2160,N_1569,N_1098);
nor U2161 (N_2161,N_1997,N_1786);
nand U2162 (N_2162,N_1304,N_1964);
nor U2163 (N_2163,N_1450,N_1949);
nand U2164 (N_2164,N_1912,N_1785);
nand U2165 (N_2165,N_1364,N_1471);
nand U2166 (N_2166,N_1361,N_1120);
nand U2167 (N_2167,N_1712,N_1876);
nor U2168 (N_2168,N_1282,N_1154);
or U2169 (N_2169,N_1160,N_1389);
and U2170 (N_2170,N_1166,N_1159);
nor U2171 (N_2171,N_1588,N_1399);
nand U2172 (N_2172,N_1520,N_1971);
nor U2173 (N_2173,N_1027,N_1238);
and U2174 (N_2174,N_1980,N_1502);
and U2175 (N_2175,N_1872,N_1560);
and U2176 (N_2176,N_1062,N_1661);
nor U2177 (N_2177,N_1808,N_1874);
or U2178 (N_2178,N_1657,N_1659);
nor U2179 (N_2179,N_1460,N_1533);
or U2180 (N_2180,N_1730,N_1688);
nor U2181 (N_2181,N_1623,N_1665);
or U2182 (N_2182,N_1096,N_1299);
nand U2183 (N_2183,N_1078,N_1136);
nand U2184 (N_2184,N_1564,N_1073);
nor U2185 (N_2185,N_1261,N_1465);
and U2186 (N_2186,N_1865,N_1229);
or U2187 (N_2187,N_1904,N_1392);
nand U2188 (N_2188,N_1601,N_1516);
or U2189 (N_2189,N_1927,N_1938);
nand U2190 (N_2190,N_1816,N_1653);
or U2191 (N_2191,N_1823,N_1033);
nand U2192 (N_2192,N_1710,N_1501);
and U2193 (N_2193,N_1703,N_1979);
or U2194 (N_2194,N_1031,N_1759);
nand U2195 (N_2195,N_1732,N_1507);
and U2196 (N_2196,N_1177,N_1833);
and U2197 (N_2197,N_1291,N_1922);
and U2198 (N_2198,N_1631,N_1369);
nor U2199 (N_2199,N_1068,N_1681);
nor U2200 (N_2200,N_1354,N_1337);
nor U2201 (N_2201,N_1735,N_1649);
xnor U2202 (N_2202,N_1385,N_1478);
nand U2203 (N_2203,N_1820,N_1755);
or U2204 (N_2204,N_1503,N_1702);
and U2205 (N_2205,N_1025,N_1375);
or U2206 (N_2206,N_1294,N_1249);
or U2207 (N_2207,N_1090,N_1113);
nand U2208 (N_2208,N_1512,N_1750);
nor U2209 (N_2209,N_1252,N_1553);
nor U2210 (N_2210,N_1495,N_1220);
and U2211 (N_2211,N_1118,N_1719);
nor U2212 (N_2212,N_1124,N_1778);
and U2213 (N_2213,N_1006,N_1855);
and U2214 (N_2214,N_1281,N_1677);
nand U2215 (N_2215,N_1846,N_1924);
nand U2216 (N_2216,N_1792,N_1775);
and U2217 (N_2217,N_1430,N_1411);
and U2218 (N_2218,N_1102,N_1518);
or U2219 (N_2219,N_1918,N_1045);
nor U2220 (N_2220,N_1339,N_1571);
or U2221 (N_2221,N_1738,N_1370);
or U2222 (N_2222,N_1158,N_1781);
nor U2223 (N_2223,N_1766,N_1187);
and U2224 (N_2224,N_1342,N_1319);
or U2225 (N_2225,N_1991,N_1329);
and U2226 (N_2226,N_1419,N_1651);
nand U2227 (N_2227,N_1506,N_1869);
nor U2228 (N_2228,N_1321,N_1350);
and U2229 (N_2229,N_1767,N_1009);
or U2230 (N_2230,N_1602,N_1194);
nand U2231 (N_2231,N_1530,N_1861);
or U2232 (N_2232,N_1546,N_1417);
or U2233 (N_2233,N_1697,N_1453);
or U2234 (N_2234,N_1390,N_1255);
nor U2235 (N_2235,N_1905,N_1038);
and U2236 (N_2236,N_1202,N_1515);
nand U2237 (N_2237,N_1568,N_1944);
nor U2238 (N_2238,N_1030,N_1799);
nand U2239 (N_2239,N_1742,N_1756);
and U2240 (N_2240,N_1379,N_1579);
and U2241 (N_2241,N_1761,N_1496);
and U2242 (N_2242,N_1203,N_1167);
and U2243 (N_2243,N_1236,N_1216);
or U2244 (N_2244,N_1868,N_1040);
nor U2245 (N_2245,N_1402,N_1176);
nor U2246 (N_2246,N_1292,N_1057);
or U2247 (N_2247,N_1836,N_1067);
nand U2248 (N_2248,N_1076,N_1327);
nor U2249 (N_2249,N_1987,N_1183);
and U2250 (N_2250,N_1807,N_1017);
and U2251 (N_2251,N_1278,N_1410);
nor U2252 (N_2252,N_1217,N_1937);
nor U2253 (N_2253,N_1204,N_1288);
and U2254 (N_2254,N_1398,N_1023);
or U2255 (N_2255,N_1161,N_1214);
and U2256 (N_2256,N_1356,N_1906);
nor U2257 (N_2257,N_1296,N_1485);
nor U2258 (N_2258,N_1140,N_1377);
and U2259 (N_2259,N_1883,N_1825);
or U2260 (N_2260,N_1976,N_1850);
nand U2261 (N_2261,N_1655,N_1162);
nor U2262 (N_2262,N_1831,N_1692);
nand U2263 (N_2263,N_1380,N_1443);
and U2264 (N_2264,N_1235,N_1745);
nand U2265 (N_2265,N_1351,N_1684);
nor U2266 (N_2266,N_1001,N_1984);
nand U2267 (N_2267,N_1801,N_1172);
xor U2268 (N_2268,N_1046,N_1232);
nor U2269 (N_2269,N_1011,N_1185);
nor U2270 (N_2270,N_1594,N_1827);
nor U2271 (N_2271,N_1211,N_1897);
or U2272 (N_2272,N_1966,N_1986);
nand U2273 (N_2273,N_1777,N_1915);
or U2274 (N_2274,N_1683,N_1112);
or U2275 (N_2275,N_1726,N_1119);
nand U2276 (N_2276,N_1673,N_1230);
nor U2277 (N_2277,N_1013,N_1610);
or U2278 (N_2278,N_1858,N_1881);
nor U2279 (N_2279,N_1760,N_1990);
nand U2280 (N_2280,N_1305,N_1464);
xor U2281 (N_2281,N_1597,N_1660);
or U2282 (N_2282,N_1892,N_1728);
and U2283 (N_2283,N_1695,N_1373);
nand U2284 (N_2284,N_1141,N_1451);
and U2285 (N_2285,N_1687,N_1890);
nor U2286 (N_2286,N_1959,N_1884);
nor U2287 (N_2287,N_1797,N_1050);
nor U2288 (N_2288,N_1313,N_1210);
or U2289 (N_2289,N_1493,N_1763);
nand U2290 (N_2290,N_1168,N_1487);
or U2291 (N_2291,N_1479,N_1157);
nand U2292 (N_2292,N_1930,N_1772);
nor U2293 (N_2293,N_1347,N_1534);
xor U2294 (N_2294,N_1522,N_1181);
and U2295 (N_2295,N_1599,N_1567);
and U2296 (N_2296,N_1839,N_1021);
and U2297 (N_2297,N_1059,N_1066);
or U2298 (N_2298,N_1129,N_1650);
or U2299 (N_2299,N_1513,N_1572);
xnor U2300 (N_2300,N_1762,N_1215);
and U2301 (N_2301,N_1490,N_1985);
and U2302 (N_2302,N_1752,N_1704);
nand U2303 (N_2303,N_1652,N_1751);
nor U2304 (N_2304,N_1500,N_1629);
and U2305 (N_2305,N_1605,N_1558);
nand U2306 (N_2306,N_1421,N_1404);
or U2307 (N_2307,N_1693,N_1699);
nor U2308 (N_2308,N_1477,N_1205);
and U2309 (N_2309,N_1722,N_1942);
nand U2310 (N_2310,N_1063,N_1773);
or U2311 (N_2311,N_1878,N_1334);
nor U2312 (N_2312,N_1951,N_1475);
nor U2313 (N_2313,N_1740,N_1967);
nor U2314 (N_2314,N_1737,N_1115);
and U2315 (N_2315,N_1627,N_1770);
nand U2316 (N_2316,N_1318,N_1452);
nand U2317 (N_2317,N_1548,N_1239);
and U2318 (N_2318,N_1283,N_1103);
nand U2319 (N_2319,N_1666,N_1819);
and U2320 (N_2320,N_1019,N_1089);
or U2321 (N_2321,N_1771,N_1169);
and U2322 (N_2322,N_1857,N_1903);
nand U2323 (N_2323,N_1504,N_1542);
and U2324 (N_2324,N_1101,N_1617);
nand U2325 (N_2325,N_1381,N_1056);
and U2326 (N_2326,N_1812,N_1246);
or U2327 (N_2327,N_1387,N_1474);
and U2328 (N_2328,N_1427,N_1946);
or U2329 (N_2329,N_1192,N_1919);
and U2330 (N_2330,N_1555,N_1219);
or U2331 (N_2331,N_1150,N_1724);
nand U2332 (N_2332,N_1358,N_1931);
and U2333 (N_2333,N_1793,N_1133);
and U2334 (N_2334,N_1257,N_1439);
or U2335 (N_2335,N_1029,N_1445);
nor U2336 (N_2336,N_1447,N_1100);
or U2337 (N_2337,N_1151,N_1260);
and U2338 (N_2338,N_1895,N_1206);
nor U2339 (N_2339,N_1322,N_1221);
or U2340 (N_2340,N_1853,N_1691);
or U2341 (N_2341,N_1311,N_1303);
nand U2342 (N_2342,N_1648,N_1948);
or U2343 (N_2343,N_1300,N_1705);
nor U2344 (N_2344,N_1898,N_1923);
nand U2345 (N_2345,N_1253,N_1896);
and U2346 (N_2346,N_1611,N_1824);
or U2347 (N_2347,N_1184,N_1301);
nand U2348 (N_2348,N_1433,N_1768);
and U2349 (N_2349,N_1913,N_1287);
nand U2350 (N_2350,N_1312,N_1123);
nand U2351 (N_2351,N_1583,N_1142);
and U2352 (N_2352,N_1295,N_1429);
or U2353 (N_2353,N_1723,N_1606);
or U2354 (N_2354,N_1810,N_1448);
or U2355 (N_2355,N_1359,N_1828);
nand U2356 (N_2356,N_1586,N_1346);
or U2357 (N_2357,N_1521,N_1473);
nand U2358 (N_2358,N_1414,N_1847);
nor U2359 (N_2359,N_1866,N_1463);
nand U2360 (N_2360,N_1111,N_1081);
nand U2361 (N_2361,N_1925,N_1307);
nand U2362 (N_2362,N_1386,N_1787);
nand U2363 (N_2363,N_1538,N_1891);
nand U2364 (N_2364,N_1352,N_1481);
nor U2365 (N_2365,N_1794,N_1805);
and U2366 (N_2366,N_1440,N_1324);
and U2367 (N_2367,N_1044,N_1146);
or U2368 (N_2368,N_1182,N_1248);
and U2369 (N_2369,N_1529,N_1663);
nand U2370 (N_2370,N_1273,N_1227);
nand U2371 (N_2371,N_1224,N_1279);
nor U2372 (N_2372,N_1727,N_1104);
nor U2373 (N_2373,N_1126,N_1435);
or U2374 (N_2374,N_1815,N_1973);
nor U2375 (N_2375,N_1911,N_1556);
or U2376 (N_2376,N_1003,N_1459);
nand U2377 (N_2377,N_1079,N_1863);
nand U2378 (N_2378,N_1734,N_1879);
nor U2379 (N_2379,N_1535,N_1993);
and U2380 (N_2380,N_1145,N_1641);
nor U2381 (N_2381,N_1813,N_1094);
nor U2382 (N_2382,N_1928,N_1498);
or U2383 (N_2383,N_1393,N_1130);
nor U2384 (N_2384,N_1237,N_1041);
or U2385 (N_2385,N_1036,N_1921);
nand U2386 (N_2386,N_1264,N_1950);
or U2387 (N_2387,N_1945,N_1071);
or U2388 (N_2388,N_1999,N_1348);
nand U2389 (N_2389,N_1559,N_1420);
or U2390 (N_2390,N_1718,N_1144);
and U2391 (N_2391,N_1268,N_1109);
nor U2392 (N_2392,N_1338,N_1254);
or U2393 (N_2393,N_1225,N_1143);
nor U2394 (N_2394,N_1998,N_1345);
nand U2395 (N_2395,N_1720,N_1566);
or U2396 (N_2396,N_1286,N_1975);
or U2397 (N_2397,N_1084,N_1272);
or U2398 (N_2398,N_1413,N_1060);
and U2399 (N_2399,N_1108,N_1989);
or U2400 (N_2400,N_1107,N_1716);
or U2401 (N_2401,N_1619,N_1198);
nand U2402 (N_2402,N_1077,N_1744);
nor U2403 (N_2403,N_1917,N_1332);
or U2404 (N_2404,N_1310,N_1106);
or U2405 (N_2405,N_1397,N_1082);
nor U2406 (N_2406,N_1640,N_1598);
xnor U2407 (N_2407,N_1782,N_1848);
nand U2408 (N_2408,N_1519,N_1746);
nand U2409 (N_2409,N_1965,N_1138);
or U2410 (N_2410,N_1156,N_1527);
nand U2411 (N_2411,N_1811,N_1754);
and U2412 (N_2412,N_1188,N_1200);
and U2413 (N_2413,N_1552,N_1037);
and U2414 (N_2414,N_1012,N_1424);
nand U2415 (N_2415,N_1069,N_1618);
or U2416 (N_2416,N_1963,N_1401);
or U2417 (N_2417,N_1624,N_1365);
or U2418 (N_2418,N_1428,N_1736);
nand U2419 (N_2419,N_1209,N_1840);
or U2420 (N_2420,N_1195,N_1947);
and U2421 (N_2421,N_1969,N_1540);
or U2422 (N_2422,N_1671,N_1197);
and U2423 (N_2423,N_1190,N_1125);
nor U2424 (N_2424,N_1462,N_1314);
nand U2425 (N_2425,N_1784,N_1409);
or U2426 (N_2426,N_1647,N_1532);
nor U2427 (N_2427,N_1668,N_1330);
or U2428 (N_2428,N_1612,N_1584);
or U2429 (N_2429,N_1802,N_1859);
or U2430 (N_2430,N_1446,N_1153);
or U2431 (N_2431,N_1829,N_1016);
nor U2432 (N_2432,N_1939,N_1580);
nor U2433 (N_2433,N_1616,N_1995);
or U2434 (N_2434,N_1565,N_1909);
nand U2435 (N_2435,N_1480,N_1297);
nor U2436 (N_2436,N_1894,N_1467);
or U2437 (N_2437,N_1591,N_1454);
nor U2438 (N_2438,N_1550,N_1039);
nor U2439 (N_2439,N_1700,N_1455);
and U2440 (N_2440,N_1072,N_1276);
nand U2441 (N_2441,N_1789,N_1431);
nor U2442 (N_2442,N_1293,N_1757);
or U2443 (N_2443,N_1054,N_1554);
and U2444 (N_2444,N_1510,N_1817);
or U2445 (N_2445,N_1099,N_1302);
nand U2446 (N_2446,N_1208,N_1020);
nor U2447 (N_2447,N_1058,N_1926);
nor U2448 (N_2448,N_1615,N_1733);
or U2449 (N_2449,N_1731,N_1047);
nand U2450 (N_2450,N_1196,N_1887);
xor U2451 (N_2451,N_1010,N_1308);
nand U2452 (N_2452,N_1241,N_1180);
nor U2453 (N_2453,N_1492,N_1885);
nand U2454 (N_2454,N_1437,N_1549);
nand U2455 (N_2455,N_1603,N_1256);
nand U2456 (N_2456,N_1637,N_1095);
nor U2457 (N_2457,N_1135,N_1394);
nand U2458 (N_2458,N_1644,N_1116);
xor U2459 (N_2459,N_1418,N_1316);
or U2460 (N_2460,N_1083,N_1609);
xor U2461 (N_2461,N_1954,N_1331);
nand U2462 (N_2462,N_1952,N_1482);
nand U2463 (N_2463,N_1686,N_1545);
nor U2464 (N_2464,N_1494,N_1367);
nand U2465 (N_2465,N_1800,N_1835);
nand U2466 (N_2466,N_1139,N_1284);
nor U2467 (N_2467,N_1932,N_1472);
or U2468 (N_2468,N_1341,N_1862);
and U2469 (N_2469,N_1958,N_1729);
nor U2470 (N_2470,N_1832,N_1933);
nor U2471 (N_2471,N_1207,N_1968);
and U2472 (N_2472,N_1764,N_1259);
nor U2473 (N_2473,N_1007,N_1837);
nor U2474 (N_2474,N_1814,N_1634);
nand U2475 (N_2475,N_1841,N_1458);
or U2476 (N_2476,N_1317,N_1573);
or U2477 (N_2477,N_1628,N_1674);
nand U2478 (N_2478,N_1642,N_1578);
xor U2479 (N_2479,N_1343,N_1679);
and U2480 (N_2480,N_1962,N_1830);
nand U2481 (N_2481,N_1250,N_1234);
nor U2482 (N_2482,N_1049,N_1355);
nand U2483 (N_2483,N_1875,N_1267);
nand U2484 (N_2484,N_1137,N_1407);
and U2485 (N_2485,N_1483,N_1741);
nor U2486 (N_2486,N_1680,N_1434);
nand U2487 (N_2487,N_1372,N_1893);
nor U2488 (N_2488,N_1186,N_1416);
or U2489 (N_2489,N_1333,N_1956);
or U2490 (N_2490,N_1270,N_1646);
and U2491 (N_2491,N_1486,N_1043);
nand U2492 (N_2492,N_1152,N_1497);
nand U2493 (N_2493,N_1769,N_1806);
nor U2494 (N_2494,N_1645,N_1362);
nand U2495 (N_2495,N_1034,N_1743);
nor U2496 (N_2496,N_1803,N_1170);
nand U2497 (N_2497,N_1382,N_1128);
and U2498 (N_2498,N_1075,N_1024);
xor U2499 (N_2499,N_1864,N_1456);
xor U2500 (N_2500,N_1173,N_1412);
or U2501 (N_2501,N_1371,N_1646);
nand U2502 (N_2502,N_1719,N_1975);
and U2503 (N_2503,N_1577,N_1373);
xnor U2504 (N_2504,N_1541,N_1075);
xor U2505 (N_2505,N_1114,N_1448);
and U2506 (N_2506,N_1235,N_1635);
nand U2507 (N_2507,N_1669,N_1338);
and U2508 (N_2508,N_1767,N_1702);
nor U2509 (N_2509,N_1484,N_1228);
or U2510 (N_2510,N_1137,N_1327);
and U2511 (N_2511,N_1444,N_1235);
nand U2512 (N_2512,N_1669,N_1733);
or U2513 (N_2513,N_1875,N_1679);
and U2514 (N_2514,N_1674,N_1192);
or U2515 (N_2515,N_1835,N_1329);
nor U2516 (N_2516,N_1328,N_1913);
and U2517 (N_2517,N_1932,N_1945);
nor U2518 (N_2518,N_1968,N_1060);
nand U2519 (N_2519,N_1960,N_1687);
nor U2520 (N_2520,N_1561,N_1280);
nor U2521 (N_2521,N_1942,N_1887);
nand U2522 (N_2522,N_1410,N_1003);
nor U2523 (N_2523,N_1976,N_1635);
and U2524 (N_2524,N_1005,N_1077);
and U2525 (N_2525,N_1228,N_1140);
nand U2526 (N_2526,N_1407,N_1781);
or U2527 (N_2527,N_1815,N_1573);
and U2528 (N_2528,N_1787,N_1003);
nand U2529 (N_2529,N_1307,N_1213);
nor U2530 (N_2530,N_1734,N_1847);
and U2531 (N_2531,N_1738,N_1261);
nor U2532 (N_2532,N_1427,N_1076);
nand U2533 (N_2533,N_1174,N_1134);
nor U2534 (N_2534,N_1598,N_1220);
and U2535 (N_2535,N_1184,N_1651);
nor U2536 (N_2536,N_1757,N_1561);
or U2537 (N_2537,N_1485,N_1879);
xnor U2538 (N_2538,N_1210,N_1738);
or U2539 (N_2539,N_1588,N_1440);
and U2540 (N_2540,N_1176,N_1447);
and U2541 (N_2541,N_1675,N_1028);
and U2542 (N_2542,N_1333,N_1972);
nand U2543 (N_2543,N_1928,N_1381);
nor U2544 (N_2544,N_1419,N_1443);
nand U2545 (N_2545,N_1459,N_1850);
or U2546 (N_2546,N_1280,N_1357);
nor U2547 (N_2547,N_1796,N_1166);
nand U2548 (N_2548,N_1618,N_1885);
and U2549 (N_2549,N_1612,N_1138);
or U2550 (N_2550,N_1479,N_1729);
nand U2551 (N_2551,N_1490,N_1707);
nor U2552 (N_2552,N_1710,N_1128);
nor U2553 (N_2553,N_1236,N_1776);
nand U2554 (N_2554,N_1090,N_1700);
nor U2555 (N_2555,N_1805,N_1713);
and U2556 (N_2556,N_1320,N_1499);
nand U2557 (N_2557,N_1484,N_1098);
and U2558 (N_2558,N_1460,N_1435);
nor U2559 (N_2559,N_1789,N_1487);
xor U2560 (N_2560,N_1449,N_1096);
or U2561 (N_2561,N_1998,N_1492);
and U2562 (N_2562,N_1354,N_1502);
xor U2563 (N_2563,N_1499,N_1998);
nor U2564 (N_2564,N_1455,N_1411);
and U2565 (N_2565,N_1778,N_1092);
nor U2566 (N_2566,N_1012,N_1062);
and U2567 (N_2567,N_1538,N_1476);
and U2568 (N_2568,N_1647,N_1978);
and U2569 (N_2569,N_1458,N_1152);
nand U2570 (N_2570,N_1010,N_1562);
and U2571 (N_2571,N_1096,N_1762);
nand U2572 (N_2572,N_1891,N_1420);
and U2573 (N_2573,N_1137,N_1873);
nand U2574 (N_2574,N_1288,N_1548);
nor U2575 (N_2575,N_1908,N_1564);
or U2576 (N_2576,N_1357,N_1679);
nor U2577 (N_2577,N_1688,N_1394);
nand U2578 (N_2578,N_1013,N_1800);
nand U2579 (N_2579,N_1965,N_1389);
and U2580 (N_2580,N_1062,N_1328);
nor U2581 (N_2581,N_1274,N_1294);
nand U2582 (N_2582,N_1667,N_1941);
and U2583 (N_2583,N_1894,N_1337);
nand U2584 (N_2584,N_1906,N_1414);
or U2585 (N_2585,N_1801,N_1472);
or U2586 (N_2586,N_1705,N_1061);
and U2587 (N_2587,N_1875,N_1773);
nand U2588 (N_2588,N_1670,N_1580);
and U2589 (N_2589,N_1682,N_1848);
xor U2590 (N_2590,N_1985,N_1161);
nand U2591 (N_2591,N_1801,N_1988);
nand U2592 (N_2592,N_1203,N_1738);
nor U2593 (N_2593,N_1286,N_1721);
and U2594 (N_2594,N_1037,N_1268);
nor U2595 (N_2595,N_1948,N_1266);
and U2596 (N_2596,N_1220,N_1352);
and U2597 (N_2597,N_1726,N_1037);
and U2598 (N_2598,N_1116,N_1134);
nand U2599 (N_2599,N_1249,N_1112);
or U2600 (N_2600,N_1052,N_1518);
nand U2601 (N_2601,N_1065,N_1176);
or U2602 (N_2602,N_1459,N_1955);
or U2603 (N_2603,N_1399,N_1330);
or U2604 (N_2604,N_1652,N_1003);
nand U2605 (N_2605,N_1111,N_1065);
nor U2606 (N_2606,N_1195,N_1930);
nand U2607 (N_2607,N_1734,N_1039);
and U2608 (N_2608,N_1826,N_1749);
or U2609 (N_2609,N_1003,N_1524);
nand U2610 (N_2610,N_1066,N_1361);
nor U2611 (N_2611,N_1197,N_1904);
nand U2612 (N_2612,N_1614,N_1718);
nor U2613 (N_2613,N_1595,N_1504);
or U2614 (N_2614,N_1521,N_1738);
or U2615 (N_2615,N_1943,N_1938);
and U2616 (N_2616,N_1071,N_1115);
nor U2617 (N_2617,N_1145,N_1318);
nand U2618 (N_2618,N_1915,N_1016);
xor U2619 (N_2619,N_1038,N_1857);
xnor U2620 (N_2620,N_1960,N_1569);
and U2621 (N_2621,N_1959,N_1746);
or U2622 (N_2622,N_1964,N_1732);
nor U2623 (N_2623,N_1675,N_1727);
nor U2624 (N_2624,N_1821,N_1357);
nor U2625 (N_2625,N_1200,N_1888);
nand U2626 (N_2626,N_1926,N_1848);
nand U2627 (N_2627,N_1194,N_1775);
nand U2628 (N_2628,N_1122,N_1838);
and U2629 (N_2629,N_1827,N_1576);
nor U2630 (N_2630,N_1648,N_1606);
and U2631 (N_2631,N_1406,N_1309);
or U2632 (N_2632,N_1409,N_1501);
nand U2633 (N_2633,N_1104,N_1916);
nand U2634 (N_2634,N_1144,N_1167);
nor U2635 (N_2635,N_1516,N_1644);
nand U2636 (N_2636,N_1297,N_1032);
or U2637 (N_2637,N_1442,N_1584);
nand U2638 (N_2638,N_1702,N_1739);
nand U2639 (N_2639,N_1702,N_1722);
and U2640 (N_2640,N_1425,N_1126);
nand U2641 (N_2641,N_1385,N_1989);
or U2642 (N_2642,N_1209,N_1015);
or U2643 (N_2643,N_1449,N_1828);
nor U2644 (N_2644,N_1725,N_1526);
and U2645 (N_2645,N_1833,N_1813);
nor U2646 (N_2646,N_1897,N_1706);
and U2647 (N_2647,N_1740,N_1248);
nand U2648 (N_2648,N_1303,N_1875);
nor U2649 (N_2649,N_1849,N_1344);
nand U2650 (N_2650,N_1904,N_1799);
xnor U2651 (N_2651,N_1041,N_1885);
nor U2652 (N_2652,N_1181,N_1139);
or U2653 (N_2653,N_1363,N_1407);
nand U2654 (N_2654,N_1385,N_1003);
and U2655 (N_2655,N_1974,N_1732);
nor U2656 (N_2656,N_1409,N_1822);
or U2657 (N_2657,N_1617,N_1192);
nand U2658 (N_2658,N_1952,N_1741);
nand U2659 (N_2659,N_1989,N_1220);
and U2660 (N_2660,N_1548,N_1161);
and U2661 (N_2661,N_1115,N_1469);
or U2662 (N_2662,N_1476,N_1239);
or U2663 (N_2663,N_1917,N_1575);
or U2664 (N_2664,N_1518,N_1173);
nor U2665 (N_2665,N_1817,N_1453);
nand U2666 (N_2666,N_1682,N_1642);
or U2667 (N_2667,N_1461,N_1903);
and U2668 (N_2668,N_1387,N_1160);
nor U2669 (N_2669,N_1061,N_1024);
nand U2670 (N_2670,N_1000,N_1064);
or U2671 (N_2671,N_1339,N_1329);
or U2672 (N_2672,N_1525,N_1354);
or U2673 (N_2673,N_1735,N_1781);
nor U2674 (N_2674,N_1683,N_1125);
nand U2675 (N_2675,N_1962,N_1657);
or U2676 (N_2676,N_1677,N_1906);
or U2677 (N_2677,N_1668,N_1741);
and U2678 (N_2678,N_1004,N_1825);
nor U2679 (N_2679,N_1920,N_1490);
nor U2680 (N_2680,N_1192,N_1080);
nor U2681 (N_2681,N_1349,N_1066);
nand U2682 (N_2682,N_1362,N_1341);
and U2683 (N_2683,N_1114,N_1378);
xnor U2684 (N_2684,N_1183,N_1742);
nor U2685 (N_2685,N_1599,N_1243);
and U2686 (N_2686,N_1133,N_1080);
and U2687 (N_2687,N_1002,N_1334);
or U2688 (N_2688,N_1678,N_1940);
or U2689 (N_2689,N_1371,N_1656);
and U2690 (N_2690,N_1161,N_1493);
or U2691 (N_2691,N_1579,N_1553);
nor U2692 (N_2692,N_1902,N_1316);
or U2693 (N_2693,N_1752,N_1242);
or U2694 (N_2694,N_1827,N_1009);
and U2695 (N_2695,N_1564,N_1271);
or U2696 (N_2696,N_1059,N_1449);
and U2697 (N_2697,N_1672,N_1362);
nand U2698 (N_2698,N_1362,N_1225);
nand U2699 (N_2699,N_1837,N_1473);
and U2700 (N_2700,N_1151,N_1131);
nor U2701 (N_2701,N_1435,N_1712);
or U2702 (N_2702,N_1072,N_1363);
or U2703 (N_2703,N_1299,N_1868);
nor U2704 (N_2704,N_1292,N_1501);
nand U2705 (N_2705,N_1028,N_1285);
and U2706 (N_2706,N_1925,N_1321);
and U2707 (N_2707,N_1169,N_1903);
nand U2708 (N_2708,N_1972,N_1167);
and U2709 (N_2709,N_1961,N_1402);
nor U2710 (N_2710,N_1288,N_1113);
and U2711 (N_2711,N_1887,N_1135);
and U2712 (N_2712,N_1522,N_1056);
nor U2713 (N_2713,N_1086,N_1821);
nor U2714 (N_2714,N_1505,N_1540);
xnor U2715 (N_2715,N_1352,N_1083);
nor U2716 (N_2716,N_1354,N_1383);
nand U2717 (N_2717,N_1490,N_1501);
and U2718 (N_2718,N_1526,N_1984);
nand U2719 (N_2719,N_1058,N_1637);
or U2720 (N_2720,N_1061,N_1682);
and U2721 (N_2721,N_1370,N_1590);
or U2722 (N_2722,N_1675,N_1911);
nand U2723 (N_2723,N_1103,N_1135);
or U2724 (N_2724,N_1891,N_1616);
nand U2725 (N_2725,N_1097,N_1270);
nor U2726 (N_2726,N_1871,N_1265);
or U2727 (N_2727,N_1141,N_1649);
nor U2728 (N_2728,N_1807,N_1645);
nand U2729 (N_2729,N_1439,N_1697);
nor U2730 (N_2730,N_1411,N_1897);
and U2731 (N_2731,N_1917,N_1896);
or U2732 (N_2732,N_1150,N_1573);
nor U2733 (N_2733,N_1865,N_1256);
nand U2734 (N_2734,N_1791,N_1004);
nand U2735 (N_2735,N_1612,N_1910);
or U2736 (N_2736,N_1367,N_1711);
and U2737 (N_2737,N_1409,N_1958);
and U2738 (N_2738,N_1759,N_1799);
or U2739 (N_2739,N_1522,N_1292);
nor U2740 (N_2740,N_1161,N_1163);
nand U2741 (N_2741,N_1785,N_1963);
nor U2742 (N_2742,N_1969,N_1370);
or U2743 (N_2743,N_1015,N_1357);
nor U2744 (N_2744,N_1940,N_1402);
nor U2745 (N_2745,N_1422,N_1269);
and U2746 (N_2746,N_1764,N_1300);
or U2747 (N_2747,N_1183,N_1581);
or U2748 (N_2748,N_1389,N_1633);
and U2749 (N_2749,N_1353,N_1863);
and U2750 (N_2750,N_1272,N_1819);
or U2751 (N_2751,N_1408,N_1768);
nand U2752 (N_2752,N_1411,N_1955);
and U2753 (N_2753,N_1717,N_1399);
or U2754 (N_2754,N_1110,N_1824);
or U2755 (N_2755,N_1534,N_1331);
nand U2756 (N_2756,N_1651,N_1894);
nor U2757 (N_2757,N_1948,N_1644);
or U2758 (N_2758,N_1903,N_1569);
or U2759 (N_2759,N_1907,N_1277);
and U2760 (N_2760,N_1047,N_1946);
nor U2761 (N_2761,N_1817,N_1074);
and U2762 (N_2762,N_1726,N_1926);
and U2763 (N_2763,N_1397,N_1907);
and U2764 (N_2764,N_1867,N_1289);
nor U2765 (N_2765,N_1399,N_1476);
nand U2766 (N_2766,N_1456,N_1746);
and U2767 (N_2767,N_1972,N_1356);
xor U2768 (N_2768,N_1882,N_1311);
nor U2769 (N_2769,N_1120,N_1158);
nand U2770 (N_2770,N_1894,N_1066);
or U2771 (N_2771,N_1139,N_1615);
and U2772 (N_2772,N_1271,N_1709);
and U2773 (N_2773,N_1744,N_1963);
or U2774 (N_2774,N_1807,N_1696);
nand U2775 (N_2775,N_1700,N_1687);
nand U2776 (N_2776,N_1479,N_1666);
or U2777 (N_2777,N_1856,N_1051);
nor U2778 (N_2778,N_1403,N_1465);
nor U2779 (N_2779,N_1418,N_1595);
and U2780 (N_2780,N_1451,N_1292);
nor U2781 (N_2781,N_1988,N_1864);
nor U2782 (N_2782,N_1363,N_1429);
xnor U2783 (N_2783,N_1827,N_1172);
nor U2784 (N_2784,N_1500,N_1777);
and U2785 (N_2785,N_1868,N_1775);
or U2786 (N_2786,N_1155,N_1584);
and U2787 (N_2787,N_1484,N_1400);
and U2788 (N_2788,N_1660,N_1573);
nand U2789 (N_2789,N_1517,N_1123);
or U2790 (N_2790,N_1909,N_1056);
nand U2791 (N_2791,N_1263,N_1734);
nand U2792 (N_2792,N_1789,N_1961);
and U2793 (N_2793,N_1298,N_1193);
and U2794 (N_2794,N_1071,N_1320);
and U2795 (N_2795,N_1455,N_1426);
nand U2796 (N_2796,N_1454,N_1617);
nand U2797 (N_2797,N_1984,N_1804);
nor U2798 (N_2798,N_1526,N_1649);
and U2799 (N_2799,N_1277,N_1626);
nand U2800 (N_2800,N_1842,N_1054);
and U2801 (N_2801,N_1902,N_1670);
nor U2802 (N_2802,N_1626,N_1264);
nand U2803 (N_2803,N_1416,N_1787);
and U2804 (N_2804,N_1548,N_1258);
or U2805 (N_2805,N_1992,N_1461);
and U2806 (N_2806,N_1154,N_1704);
or U2807 (N_2807,N_1402,N_1661);
or U2808 (N_2808,N_1143,N_1353);
and U2809 (N_2809,N_1969,N_1415);
and U2810 (N_2810,N_1027,N_1144);
nand U2811 (N_2811,N_1665,N_1410);
or U2812 (N_2812,N_1505,N_1021);
and U2813 (N_2813,N_1954,N_1320);
nor U2814 (N_2814,N_1403,N_1371);
and U2815 (N_2815,N_1133,N_1953);
or U2816 (N_2816,N_1948,N_1087);
nand U2817 (N_2817,N_1442,N_1708);
and U2818 (N_2818,N_1526,N_1231);
or U2819 (N_2819,N_1921,N_1389);
nand U2820 (N_2820,N_1932,N_1087);
nand U2821 (N_2821,N_1574,N_1804);
nor U2822 (N_2822,N_1205,N_1638);
and U2823 (N_2823,N_1698,N_1601);
or U2824 (N_2824,N_1045,N_1528);
or U2825 (N_2825,N_1969,N_1191);
nor U2826 (N_2826,N_1561,N_1367);
nand U2827 (N_2827,N_1752,N_1984);
and U2828 (N_2828,N_1593,N_1789);
or U2829 (N_2829,N_1215,N_1492);
nor U2830 (N_2830,N_1314,N_1569);
and U2831 (N_2831,N_1487,N_1586);
nand U2832 (N_2832,N_1890,N_1721);
nand U2833 (N_2833,N_1177,N_1055);
and U2834 (N_2834,N_1264,N_1277);
or U2835 (N_2835,N_1895,N_1033);
or U2836 (N_2836,N_1162,N_1775);
nand U2837 (N_2837,N_1299,N_1126);
nand U2838 (N_2838,N_1090,N_1414);
nand U2839 (N_2839,N_1024,N_1021);
nor U2840 (N_2840,N_1189,N_1675);
and U2841 (N_2841,N_1050,N_1982);
nor U2842 (N_2842,N_1557,N_1773);
or U2843 (N_2843,N_1807,N_1536);
nand U2844 (N_2844,N_1135,N_1719);
or U2845 (N_2845,N_1993,N_1996);
nand U2846 (N_2846,N_1865,N_1382);
or U2847 (N_2847,N_1201,N_1896);
and U2848 (N_2848,N_1078,N_1448);
and U2849 (N_2849,N_1724,N_1514);
or U2850 (N_2850,N_1644,N_1658);
nand U2851 (N_2851,N_1381,N_1879);
nor U2852 (N_2852,N_1312,N_1130);
and U2853 (N_2853,N_1866,N_1808);
nand U2854 (N_2854,N_1150,N_1084);
nor U2855 (N_2855,N_1814,N_1030);
or U2856 (N_2856,N_1359,N_1471);
nand U2857 (N_2857,N_1759,N_1422);
and U2858 (N_2858,N_1794,N_1835);
xor U2859 (N_2859,N_1318,N_1024);
or U2860 (N_2860,N_1487,N_1262);
nand U2861 (N_2861,N_1320,N_1397);
and U2862 (N_2862,N_1114,N_1777);
or U2863 (N_2863,N_1381,N_1358);
nor U2864 (N_2864,N_1142,N_1351);
nor U2865 (N_2865,N_1699,N_1490);
and U2866 (N_2866,N_1196,N_1920);
or U2867 (N_2867,N_1152,N_1158);
nor U2868 (N_2868,N_1478,N_1346);
nor U2869 (N_2869,N_1352,N_1667);
or U2870 (N_2870,N_1941,N_1636);
nand U2871 (N_2871,N_1420,N_1906);
nor U2872 (N_2872,N_1791,N_1353);
and U2873 (N_2873,N_1945,N_1280);
nor U2874 (N_2874,N_1602,N_1964);
nand U2875 (N_2875,N_1365,N_1800);
nand U2876 (N_2876,N_1868,N_1733);
nand U2877 (N_2877,N_1585,N_1805);
or U2878 (N_2878,N_1678,N_1636);
nand U2879 (N_2879,N_1778,N_1532);
xnor U2880 (N_2880,N_1903,N_1452);
nor U2881 (N_2881,N_1604,N_1808);
nand U2882 (N_2882,N_1996,N_1606);
or U2883 (N_2883,N_1206,N_1608);
and U2884 (N_2884,N_1796,N_1955);
and U2885 (N_2885,N_1797,N_1862);
or U2886 (N_2886,N_1570,N_1352);
or U2887 (N_2887,N_1995,N_1396);
nor U2888 (N_2888,N_1950,N_1341);
and U2889 (N_2889,N_1818,N_1353);
nand U2890 (N_2890,N_1291,N_1112);
and U2891 (N_2891,N_1005,N_1958);
and U2892 (N_2892,N_1136,N_1604);
and U2893 (N_2893,N_1376,N_1143);
and U2894 (N_2894,N_1859,N_1705);
nand U2895 (N_2895,N_1349,N_1734);
nand U2896 (N_2896,N_1429,N_1413);
nand U2897 (N_2897,N_1290,N_1571);
or U2898 (N_2898,N_1389,N_1307);
or U2899 (N_2899,N_1523,N_1739);
or U2900 (N_2900,N_1145,N_1778);
and U2901 (N_2901,N_1598,N_1423);
nor U2902 (N_2902,N_1826,N_1766);
nand U2903 (N_2903,N_1459,N_1714);
or U2904 (N_2904,N_1720,N_1914);
and U2905 (N_2905,N_1318,N_1504);
or U2906 (N_2906,N_1620,N_1929);
nor U2907 (N_2907,N_1538,N_1015);
or U2908 (N_2908,N_1904,N_1127);
nand U2909 (N_2909,N_1995,N_1161);
and U2910 (N_2910,N_1131,N_1991);
nand U2911 (N_2911,N_1770,N_1851);
nor U2912 (N_2912,N_1163,N_1439);
and U2913 (N_2913,N_1753,N_1166);
nand U2914 (N_2914,N_1725,N_1651);
nand U2915 (N_2915,N_1163,N_1044);
and U2916 (N_2916,N_1626,N_1293);
or U2917 (N_2917,N_1122,N_1548);
nand U2918 (N_2918,N_1055,N_1346);
and U2919 (N_2919,N_1956,N_1332);
and U2920 (N_2920,N_1446,N_1268);
or U2921 (N_2921,N_1331,N_1931);
nand U2922 (N_2922,N_1082,N_1249);
or U2923 (N_2923,N_1249,N_1938);
nor U2924 (N_2924,N_1891,N_1095);
or U2925 (N_2925,N_1288,N_1987);
nor U2926 (N_2926,N_1538,N_1943);
nand U2927 (N_2927,N_1322,N_1189);
or U2928 (N_2928,N_1835,N_1539);
nand U2929 (N_2929,N_1500,N_1687);
and U2930 (N_2930,N_1536,N_1897);
nor U2931 (N_2931,N_1453,N_1234);
nor U2932 (N_2932,N_1506,N_1968);
and U2933 (N_2933,N_1685,N_1403);
and U2934 (N_2934,N_1532,N_1252);
nand U2935 (N_2935,N_1319,N_1736);
nor U2936 (N_2936,N_1450,N_1954);
or U2937 (N_2937,N_1380,N_1653);
nor U2938 (N_2938,N_1144,N_1481);
nor U2939 (N_2939,N_1782,N_1280);
nand U2940 (N_2940,N_1995,N_1543);
nor U2941 (N_2941,N_1097,N_1512);
and U2942 (N_2942,N_1241,N_1206);
or U2943 (N_2943,N_1378,N_1092);
and U2944 (N_2944,N_1754,N_1396);
and U2945 (N_2945,N_1135,N_1785);
and U2946 (N_2946,N_1824,N_1384);
nand U2947 (N_2947,N_1321,N_1694);
nand U2948 (N_2948,N_1999,N_1046);
nor U2949 (N_2949,N_1188,N_1159);
and U2950 (N_2950,N_1618,N_1913);
nor U2951 (N_2951,N_1920,N_1254);
or U2952 (N_2952,N_1001,N_1106);
nand U2953 (N_2953,N_1921,N_1423);
nand U2954 (N_2954,N_1296,N_1881);
nand U2955 (N_2955,N_1917,N_1139);
nand U2956 (N_2956,N_1862,N_1531);
nand U2957 (N_2957,N_1284,N_1385);
and U2958 (N_2958,N_1666,N_1307);
nand U2959 (N_2959,N_1622,N_1119);
or U2960 (N_2960,N_1177,N_1652);
nor U2961 (N_2961,N_1924,N_1891);
and U2962 (N_2962,N_1087,N_1124);
or U2963 (N_2963,N_1039,N_1383);
nand U2964 (N_2964,N_1635,N_1471);
or U2965 (N_2965,N_1456,N_1001);
and U2966 (N_2966,N_1135,N_1761);
nand U2967 (N_2967,N_1955,N_1365);
and U2968 (N_2968,N_1022,N_1708);
nand U2969 (N_2969,N_1075,N_1921);
or U2970 (N_2970,N_1218,N_1258);
or U2971 (N_2971,N_1742,N_1116);
nand U2972 (N_2972,N_1219,N_1949);
and U2973 (N_2973,N_1654,N_1421);
or U2974 (N_2974,N_1537,N_1270);
nand U2975 (N_2975,N_1513,N_1157);
and U2976 (N_2976,N_1089,N_1448);
nor U2977 (N_2977,N_1424,N_1269);
or U2978 (N_2978,N_1497,N_1306);
xor U2979 (N_2979,N_1349,N_1501);
and U2980 (N_2980,N_1584,N_1066);
nor U2981 (N_2981,N_1060,N_1393);
and U2982 (N_2982,N_1429,N_1210);
nor U2983 (N_2983,N_1883,N_1195);
nand U2984 (N_2984,N_1233,N_1089);
nor U2985 (N_2985,N_1432,N_1388);
nor U2986 (N_2986,N_1377,N_1066);
nor U2987 (N_2987,N_1820,N_1867);
or U2988 (N_2988,N_1090,N_1380);
and U2989 (N_2989,N_1877,N_1831);
nor U2990 (N_2990,N_1394,N_1459);
or U2991 (N_2991,N_1294,N_1306);
and U2992 (N_2992,N_1271,N_1894);
xnor U2993 (N_2993,N_1481,N_1502);
nand U2994 (N_2994,N_1327,N_1116);
or U2995 (N_2995,N_1740,N_1281);
or U2996 (N_2996,N_1839,N_1345);
nand U2997 (N_2997,N_1759,N_1358);
nand U2998 (N_2998,N_1347,N_1590);
or U2999 (N_2999,N_1850,N_1205);
and U3000 (N_3000,N_2023,N_2356);
and U3001 (N_3001,N_2516,N_2351);
xor U3002 (N_3002,N_2521,N_2820);
nand U3003 (N_3003,N_2988,N_2380);
and U3004 (N_3004,N_2155,N_2900);
or U3005 (N_3005,N_2305,N_2086);
xnor U3006 (N_3006,N_2314,N_2401);
nor U3007 (N_3007,N_2689,N_2211);
nor U3008 (N_3008,N_2686,N_2447);
and U3009 (N_3009,N_2428,N_2239);
and U3010 (N_3010,N_2697,N_2242);
nand U3011 (N_3011,N_2137,N_2912);
and U3012 (N_3012,N_2021,N_2538);
and U3013 (N_3013,N_2745,N_2321);
and U3014 (N_3014,N_2678,N_2633);
or U3015 (N_3015,N_2092,N_2814);
nor U3016 (N_3016,N_2306,N_2655);
and U3017 (N_3017,N_2354,N_2691);
and U3018 (N_3018,N_2634,N_2954);
and U3019 (N_3019,N_2492,N_2527);
nand U3020 (N_3020,N_2225,N_2790);
or U3021 (N_3021,N_2709,N_2270);
and U3022 (N_3022,N_2374,N_2440);
nand U3023 (N_3023,N_2475,N_2404);
nand U3024 (N_3024,N_2570,N_2536);
nand U3025 (N_3025,N_2661,N_2542);
nor U3026 (N_3026,N_2108,N_2269);
and U3027 (N_3027,N_2600,N_2808);
nand U3028 (N_3028,N_2220,N_2638);
nor U3029 (N_3029,N_2913,N_2559);
and U3030 (N_3030,N_2131,N_2977);
and U3031 (N_3031,N_2961,N_2624);
and U3032 (N_3032,N_2048,N_2959);
nor U3033 (N_3033,N_2972,N_2489);
nand U3034 (N_3034,N_2857,N_2387);
nor U3035 (N_3035,N_2552,N_2893);
or U3036 (N_3036,N_2484,N_2293);
nor U3037 (N_3037,N_2282,N_2585);
nor U3038 (N_3038,N_2568,N_2158);
nor U3039 (N_3039,N_2557,N_2353);
xor U3040 (N_3040,N_2813,N_2718);
and U3041 (N_3041,N_2599,N_2271);
nor U3042 (N_3042,N_2199,N_2236);
xor U3043 (N_3043,N_2402,N_2554);
nand U3044 (N_3044,N_2160,N_2576);
nand U3045 (N_3045,N_2856,N_2839);
or U3046 (N_3046,N_2964,N_2509);
and U3047 (N_3047,N_2513,N_2304);
or U3048 (N_3048,N_2241,N_2965);
nand U3049 (N_3049,N_2230,N_2692);
nand U3050 (N_3050,N_2317,N_2300);
nand U3051 (N_3051,N_2760,N_2165);
nand U3052 (N_3052,N_2435,N_2099);
or U3053 (N_3053,N_2997,N_2560);
nor U3054 (N_3054,N_2501,N_2342);
nand U3055 (N_3055,N_2916,N_2938);
nor U3056 (N_3056,N_2382,N_2748);
or U3057 (N_3057,N_2188,N_2334);
nor U3058 (N_3058,N_2641,N_2054);
and U3059 (N_3059,N_2053,N_2962);
nand U3060 (N_3060,N_2181,N_2076);
and U3061 (N_3061,N_2528,N_2672);
nand U3062 (N_3062,N_2622,N_2135);
or U3063 (N_3063,N_2246,N_2629);
and U3064 (N_3064,N_2882,N_2326);
nor U3065 (N_3065,N_2545,N_2684);
and U3066 (N_3066,N_2454,N_2470);
xor U3067 (N_3067,N_2022,N_2788);
nor U3068 (N_3068,N_2381,N_2315);
nor U3069 (N_3069,N_2819,N_2416);
nor U3070 (N_3070,N_2039,N_2118);
or U3071 (N_3071,N_2892,N_2504);
nand U3072 (N_3072,N_2758,N_2966);
or U3073 (N_3073,N_2045,N_2761);
or U3074 (N_3074,N_2187,N_2647);
nor U3075 (N_3075,N_2297,N_2247);
nand U3076 (N_3076,N_2734,N_2073);
nand U3077 (N_3077,N_2915,N_2606);
nand U3078 (N_3078,N_2415,N_2001);
or U3079 (N_3079,N_2040,N_2626);
nand U3080 (N_3080,N_2384,N_2620);
and U3081 (N_3081,N_2403,N_2098);
or U3082 (N_3082,N_2074,N_2782);
and U3083 (N_3083,N_2574,N_2083);
nand U3084 (N_3084,N_2170,N_2849);
nand U3085 (N_3085,N_2172,N_2979);
and U3086 (N_3086,N_2291,N_2324);
or U3087 (N_3087,N_2990,N_2422);
or U3088 (N_3088,N_2350,N_2320);
and U3089 (N_3089,N_2095,N_2936);
and U3090 (N_3090,N_2658,N_2056);
and U3091 (N_3091,N_2737,N_2925);
nand U3092 (N_3092,N_2649,N_2227);
nor U3093 (N_3093,N_2609,N_2464);
or U3094 (N_3094,N_2153,N_2329);
nand U3095 (N_3095,N_2847,N_2526);
and U3096 (N_3096,N_2453,N_2698);
nor U3097 (N_3097,N_2205,N_2340);
nand U3098 (N_3098,N_2926,N_2590);
and U3099 (N_3099,N_2244,N_2343);
and U3100 (N_3100,N_2569,N_2399);
nor U3101 (N_3101,N_2414,N_2749);
or U3102 (N_3102,N_2166,N_2100);
nand U3103 (N_3103,N_2676,N_2087);
and U3104 (N_3104,N_2327,N_2630);
xnor U3105 (N_3105,N_2763,N_2046);
or U3106 (N_3106,N_2379,N_2460);
or U3107 (N_3107,N_2645,N_2112);
or U3108 (N_3108,N_2935,N_2002);
nor U3109 (N_3109,N_2774,N_2794);
nor U3110 (N_3110,N_2250,N_2715);
or U3111 (N_3111,N_2840,N_2871);
or U3112 (N_3112,N_2529,N_2923);
nand U3113 (N_3113,N_2796,N_2174);
and U3114 (N_3114,N_2855,N_2822);
nor U3115 (N_3115,N_2369,N_2419);
and U3116 (N_3116,N_2746,N_2911);
and U3117 (N_3117,N_2011,N_2178);
nand U3118 (N_3118,N_2996,N_2807);
and U3119 (N_3119,N_2680,N_2156);
nand U3120 (N_3120,N_2117,N_2891);
or U3121 (N_3121,N_2660,N_2206);
xnor U3122 (N_3122,N_2821,N_2832);
nand U3123 (N_3123,N_2260,N_2062);
and U3124 (N_3124,N_2522,N_2503);
nor U3125 (N_3125,N_2751,N_2555);
and U3126 (N_3126,N_2251,N_2496);
and U3127 (N_3127,N_2104,N_2614);
or U3128 (N_3128,N_2082,N_2601);
nand U3129 (N_3129,N_2121,N_2427);
or U3130 (N_3130,N_2989,N_2115);
nor U3131 (N_3131,N_2514,N_2922);
nor U3132 (N_3132,N_2096,N_2420);
xor U3133 (N_3133,N_2025,N_2237);
or U3134 (N_3134,N_2278,N_2478);
nand U3135 (N_3135,N_2548,N_2481);
nor U3136 (N_3136,N_2815,N_2258);
nor U3137 (N_3137,N_2063,N_2721);
nor U3138 (N_3138,N_2279,N_2307);
nand U3139 (N_3139,N_2009,N_2603);
nor U3140 (N_3140,N_2951,N_2147);
or U3141 (N_3141,N_2640,N_2969);
nor U3142 (N_3142,N_2176,N_2543);
and U3143 (N_3143,N_2049,N_2488);
and U3144 (N_3144,N_2345,N_2332);
or U3145 (N_3145,N_2927,N_2311);
nor U3146 (N_3146,N_2373,N_2519);
nor U3147 (N_3147,N_2703,N_2993);
and U3148 (N_3148,N_2248,N_2862);
or U3149 (N_3149,N_2066,N_2755);
nand U3150 (N_3150,N_2224,N_2852);
nand U3151 (N_3151,N_2704,N_2101);
nor U3152 (N_3152,N_2941,N_2446);
and U3153 (N_3153,N_2722,N_2602);
nor U3154 (N_3154,N_2143,N_2587);
or U3155 (N_3155,N_2879,N_2854);
and U3156 (N_3156,N_2970,N_2508);
and U3157 (N_3157,N_2673,N_2204);
and U3158 (N_3158,N_2567,N_2268);
or U3159 (N_3159,N_2303,N_2865);
or U3160 (N_3160,N_2395,N_2799);
xor U3161 (N_3161,N_2418,N_2594);
nor U3162 (N_3162,N_2823,N_2675);
and U3163 (N_3163,N_2877,N_2598);
or U3164 (N_3164,N_2141,N_2829);
nor U3165 (N_3165,N_2383,N_2531);
and U3166 (N_3166,N_2967,N_2360);
nor U3167 (N_3167,N_2439,N_2848);
and U3168 (N_3168,N_2215,N_2836);
nor U3169 (N_3169,N_2093,N_2408);
nand U3170 (N_3170,N_2319,N_2006);
or U3171 (N_3171,N_2253,N_2605);
nand U3172 (N_3172,N_2263,N_2842);
and U3173 (N_3173,N_2671,N_2019);
and U3174 (N_3174,N_2400,N_2541);
and U3175 (N_3175,N_2608,N_2449);
nor U3176 (N_3176,N_2889,N_2667);
nor U3177 (N_3177,N_2267,N_2929);
nand U3178 (N_3178,N_2586,N_2029);
and U3179 (N_3179,N_2679,N_2287);
nor U3180 (N_3180,N_2752,N_2824);
nand U3181 (N_3181,N_2057,N_2412);
nand U3182 (N_3182,N_2370,N_2284);
or U3183 (N_3183,N_2637,N_2072);
or U3184 (N_3184,N_2851,N_2471);
nand U3185 (N_3185,N_2249,N_2525);
or U3186 (N_3186,N_2195,N_2766);
nor U3187 (N_3187,N_2580,N_2068);
nor U3188 (N_3188,N_2308,N_2845);
nor U3189 (N_3189,N_2597,N_2750);
or U3190 (N_3190,N_2533,N_2331);
nand U3191 (N_3191,N_2059,N_2981);
nor U3192 (N_3192,N_2802,N_2907);
nand U3193 (N_3193,N_2222,N_2575);
nor U3194 (N_3194,N_2274,N_2659);
nor U3195 (N_3195,N_2299,N_2480);
or U3196 (N_3196,N_2716,N_2785);
and U3197 (N_3197,N_2391,N_2456);
nand U3198 (N_3198,N_2151,N_2301);
nor U3199 (N_3199,N_2264,N_2589);
nor U3200 (N_3200,N_2051,N_2860);
nand U3201 (N_3201,N_2731,N_2775);
or U3202 (N_3202,N_2119,N_2372);
and U3203 (N_3203,N_2789,N_2757);
or U3204 (N_3204,N_2359,N_2458);
or U3205 (N_3205,N_2732,N_2357);
nor U3206 (N_3206,N_2201,N_2719);
or U3207 (N_3207,N_2266,N_2825);
or U3208 (N_3208,N_2561,N_2050);
nand U3209 (N_3209,N_2393,N_2411);
nor U3210 (N_3210,N_2210,N_2708);
nand U3211 (N_3211,N_2896,N_2336);
and U3212 (N_3212,N_2726,N_2127);
or U3213 (N_3213,N_2706,N_2656);
xnor U3214 (N_3214,N_2777,N_2450);
nor U3215 (N_3215,N_2347,N_2872);
and U3216 (N_3216,N_2619,N_2012);
or U3217 (N_3217,N_2505,N_2474);
nor U3218 (N_3218,N_2621,N_2956);
nor U3219 (N_3219,N_2459,N_2910);
or U3220 (N_3220,N_2610,N_2067);
nor U3221 (N_3221,N_2413,N_2125);
nand U3222 (N_3222,N_2358,N_2710);
and U3223 (N_3223,N_2764,N_2133);
nor U3224 (N_3224,N_2060,N_2218);
and U3225 (N_3225,N_2994,N_2540);
xnor U3226 (N_3226,N_2566,N_2801);
nand U3227 (N_3227,N_2616,N_2216);
and U3228 (N_3228,N_2874,N_2390);
nand U3229 (N_3229,N_2363,N_2759);
or U3230 (N_3230,N_2000,N_2762);
xor U3231 (N_3231,N_2203,N_2613);
nand U3232 (N_3232,N_2998,N_2036);
or U3233 (N_3233,N_2070,N_2903);
or U3234 (N_3234,N_2940,N_2438);
nand U3235 (N_3235,N_2114,N_2277);
or U3236 (N_3236,N_2681,N_2429);
and U3237 (N_3237,N_2102,N_2385);
and U3238 (N_3238,N_2939,N_2577);
nor U3239 (N_3239,N_2946,N_2725);
or U3240 (N_3240,N_2469,N_2448);
or U3241 (N_3241,N_2344,N_2787);
nand U3242 (N_3242,N_2631,N_2739);
nor U3243 (N_3243,N_2375,N_2983);
and U3244 (N_3244,N_2714,N_2804);
or U3245 (N_3245,N_2265,N_2564);
or U3246 (N_3246,N_2423,N_2713);
nor U3247 (N_3247,N_2743,N_2221);
or U3248 (N_3248,N_2583,N_2890);
xnor U3249 (N_3249,N_2677,N_2674);
and U3250 (N_3250,N_2261,N_2873);
nor U3251 (N_3251,N_2611,N_2506);
nand U3252 (N_3252,N_2535,N_2846);
or U3253 (N_3253,N_2843,N_2733);
or U3254 (N_3254,N_2349,N_2200);
nor U3255 (N_3255,N_2779,N_2955);
and U3256 (N_3256,N_2957,N_2835);
or U3257 (N_3257,N_2933,N_2693);
nor U3258 (N_3258,N_2867,N_2768);
and U3259 (N_3259,N_2861,N_2431);
nand U3260 (N_3260,N_2549,N_2126);
nand U3261 (N_3261,N_2409,N_2717);
or U3262 (N_3262,N_2858,N_2736);
nand U3263 (N_3263,N_2361,N_2335);
nor U3264 (N_3264,N_2537,N_2784);
and U3265 (N_3265,N_2666,N_2652);
xor U3266 (N_3266,N_2240,N_2798);
or U3267 (N_3267,N_2280,N_2037);
nand U3268 (N_3268,N_2088,N_2812);
and U3269 (N_3269,N_2662,N_2213);
or U3270 (N_3270,N_2288,N_2985);
and U3271 (N_3271,N_2163,N_2604);
and U3272 (N_3272,N_2052,N_2417);
or U3273 (N_3273,N_2883,N_2032);
and U3274 (N_3274,N_2235,N_2312);
nand U3275 (N_3275,N_2497,N_2124);
and U3276 (N_3276,N_2364,N_2130);
or U3277 (N_3277,N_2931,N_2573);
and U3278 (N_3278,N_2313,N_2971);
nor U3279 (N_3279,N_2744,N_2817);
or U3280 (N_3280,N_2534,N_2139);
nor U3281 (N_3281,N_2337,N_2781);
or U3282 (N_3282,N_2974,N_2878);
or U3283 (N_3283,N_2058,N_2175);
and U3284 (N_3284,N_2272,N_2255);
nor U3285 (N_3285,N_2097,N_2302);
nor U3286 (N_3286,N_2436,N_2167);
and U3287 (N_3287,N_2657,N_2193);
or U3288 (N_3288,N_2665,N_2368);
or U3289 (N_3289,N_2451,N_2027);
and U3290 (N_3290,N_2226,N_2999);
nor U3291 (N_3291,N_2844,N_2491);
or U3292 (N_3292,N_2517,N_2180);
or U3293 (N_3293,N_2323,N_2984);
nor U3294 (N_3294,N_2378,N_2389);
nor U3295 (N_3295,N_2171,N_2355);
nor U3296 (N_3296,N_2243,N_2198);
or U3297 (N_3297,N_2229,N_2132);
xnor U3298 (N_3298,N_2795,N_2930);
or U3299 (N_3299,N_2105,N_2982);
and U3300 (N_3300,N_2079,N_2123);
nand U3301 (N_3301,N_2367,N_2341);
and U3302 (N_3302,N_2864,N_2191);
nor U3303 (N_3303,N_2003,N_2376);
or U3304 (N_3304,N_2394,N_2701);
nand U3305 (N_3305,N_2421,N_2887);
nor U3306 (N_3306,N_2562,N_2034);
and U3307 (N_3307,N_2841,N_2273);
nor U3308 (N_3308,N_2008,N_2806);
nand U3309 (N_3309,N_2651,N_2473);
nor U3310 (N_3310,N_2122,N_2146);
and U3311 (N_3311,N_2081,N_2909);
or U3312 (N_3312,N_2285,N_2581);
nor U3313 (N_3313,N_2905,N_2138);
xnor U3314 (N_3314,N_2038,N_2884);
and U3315 (N_3315,N_2120,N_2047);
nor U3316 (N_3316,N_2833,N_2477);
and U3317 (N_3317,N_2699,N_2077);
nand U3318 (N_3318,N_2712,N_2546);
xnor U3319 (N_3319,N_2924,N_2392);
nand U3320 (N_3320,N_2705,N_2043);
or U3321 (N_3321,N_2510,N_2544);
nor U3322 (N_3322,N_2828,N_2209);
nor U3323 (N_3323,N_2149,N_2711);
xnor U3324 (N_3324,N_2588,N_2623);
nor U3325 (N_3325,N_2283,N_2441);
nor U3326 (N_3326,N_2007,N_2500);
nand U3327 (N_3327,N_2579,N_2030);
xor U3328 (N_3328,N_2430,N_2452);
or U3329 (N_3329,N_2129,N_2238);
nand U3330 (N_3330,N_2257,N_2457);
nor U3331 (N_3331,N_2978,N_2702);
nor U3332 (N_3332,N_2767,N_2695);
nand U3333 (N_3333,N_2182,N_2869);
or U3334 (N_3334,N_2352,N_2868);
nand U3335 (N_3335,N_2031,N_2770);
and U3336 (N_3336,N_2830,N_2639);
nor U3337 (N_3337,N_2948,N_2479);
nor U3338 (N_3338,N_2042,N_2553);
nor U3339 (N_3339,N_2897,N_2952);
nor U3340 (N_3340,N_2424,N_2811);
or U3341 (N_3341,N_2793,N_2729);
and U3342 (N_3342,N_2837,N_2859);
nor U3343 (N_3343,N_2189,N_2918);
and U3344 (N_3344,N_2863,N_2906);
and U3345 (N_3345,N_2885,N_2532);
or U3346 (N_3346,N_2720,N_2366);
nand U3347 (N_3347,N_2013,N_2208);
or U3348 (N_3348,N_2650,N_2362);
or U3349 (N_3349,N_2168,N_2466);
and U3350 (N_3350,N_2571,N_2017);
nand U3351 (N_3351,N_2018,N_2898);
nand U3352 (N_3352,N_2875,N_2472);
or U3353 (N_3353,N_2563,N_2128);
and U3354 (N_3354,N_2944,N_2894);
and U3355 (N_3355,N_2333,N_2520);
or U3356 (N_3356,N_2730,N_2850);
and U3357 (N_3357,N_2330,N_2084);
nand U3358 (N_3358,N_2467,N_2584);
xnor U3359 (N_3359,N_2325,N_2578);
nand U3360 (N_3360,N_2556,N_2294);
nand U3361 (N_3361,N_2190,N_2202);
or U3362 (N_3362,N_2365,N_2089);
and U3363 (N_3363,N_2953,N_2618);
or U3364 (N_3364,N_2328,N_2914);
and U3365 (N_3365,N_2476,N_2463);
nand U3366 (N_3366,N_2169,N_2738);
or U3367 (N_3367,N_2765,N_2668);
or U3368 (N_3368,N_2065,N_2632);
or U3369 (N_3369,N_2783,N_2499);
nor U3370 (N_3370,N_2116,N_2186);
and U3371 (N_3371,N_2157,N_2196);
or U3372 (N_3372,N_2826,N_2539);
and U3373 (N_3373,N_2377,N_2346);
nand U3374 (N_3374,N_2724,N_2524);
or U3375 (N_3375,N_2776,N_2809);
and U3376 (N_3376,N_2643,N_2075);
nor U3377 (N_3377,N_2292,N_2061);
or U3378 (N_3378,N_2986,N_2976);
or U3379 (N_3379,N_2735,N_2173);
nor U3380 (N_3380,N_2803,N_2932);
nor U3381 (N_3381,N_2485,N_2164);
and U3382 (N_3382,N_2968,N_2465);
or U3383 (N_3383,N_2800,N_2853);
nand U3384 (N_3384,N_2033,N_2487);
nor U3385 (N_3385,N_2742,N_2192);
or U3386 (N_3386,N_2425,N_2483);
and U3387 (N_3387,N_2917,N_2490);
and U3388 (N_3388,N_2498,N_2339);
and U3389 (N_3389,N_2035,N_2444);
and U3390 (N_3390,N_2627,N_2904);
and U3391 (N_3391,N_2664,N_2947);
nor U3392 (N_3392,N_2309,N_2593);
or U3393 (N_3393,N_2442,N_2407);
nand U3394 (N_3394,N_2572,N_2565);
nand U3395 (N_3395,N_2295,N_2612);
nor U3396 (N_3396,N_2493,N_2973);
nor U3397 (N_3397,N_2773,N_2014);
and U3398 (N_3398,N_2682,N_2886);
nor U3399 (N_3399,N_2512,N_2296);
and U3400 (N_3400,N_2223,N_2895);
and U3401 (N_3401,N_2024,N_2870);
or U3402 (N_3402,N_2145,N_2792);
nor U3403 (N_3403,N_2669,N_2142);
and U3404 (N_3404,N_2310,N_2461);
and U3405 (N_3405,N_2184,N_2595);
nand U3406 (N_3406,N_2942,N_2410);
nand U3407 (N_3407,N_2318,N_2831);
or U3408 (N_3408,N_2592,N_2016);
nor U3409 (N_3409,N_2992,N_2044);
nand U3410 (N_3410,N_2607,N_2502);
nand U3411 (N_3411,N_2080,N_2110);
and U3412 (N_3412,N_2880,N_2960);
nand U3413 (N_3413,N_2107,N_2183);
nand U3414 (N_3414,N_2111,N_2094);
xnor U3415 (N_3415,N_2432,N_2338);
nor U3416 (N_3416,N_2615,N_2834);
nor U3417 (N_3417,N_2069,N_2636);
nor U3418 (N_3418,N_2754,N_2728);
nor U3419 (N_3419,N_2004,N_2197);
or U3420 (N_3420,N_2109,N_2975);
nand U3421 (N_3421,N_2217,N_2426);
nand U3422 (N_3422,N_2262,N_2005);
nor U3423 (N_3423,N_2219,N_2908);
nand U3424 (N_3424,N_2140,N_2443);
or U3425 (N_3425,N_2797,N_2259);
xnor U3426 (N_3426,N_2136,N_2995);
nand U3427 (N_3427,N_2159,N_2214);
nand U3428 (N_3428,N_2617,N_2397);
nor U3429 (N_3429,N_2298,N_2495);
or U3430 (N_3430,N_2388,N_2635);
nand U3431 (N_3431,N_2769,N_2434);
nor U3432 (N_3432,N_2228,N_2462);
xnor U3433 (N_3433,N_2596,N_2551);
or U3434 (N_3434,N_2161,N_2591);
and U3435 (N_3435,N_2547,N_2991);
nor U3436 (N_3436,N_2254,N_2179);
and U3437 (N_3437,N_2753,N_2015);
and U3438 (N_3438,N_2177,N_2185);
nor U3439 (N_3439,N_2276,N_2644);
and U3440 (N_3440,N_2106,N_2433);
nand U3441 (N_3441,N_2888,N_2690);
and U3442 (N_3442,N_2289,N_2286);
nand U3443 (N_3443,N_2928,N_2950);
nand U3444 (N_3444,N_2234,N_2778);
or U3445 (N_3445,N_2683,N_2945);
or U3446 (N_3446,N_2281,N_2064);
nand U3447 (N_3447,N_2154,N_2091);
or U3448 (N_3448,N_2515,N_2980);
or U3449 (N_3449,N_2685,N_2902);
nand U3450 (N_3450,N_2756,N_2398);
or U3451 (N_3451,N_2468,N_2558);
nor U3452 (N_3452,N_2899,N_2881);
nor U3453 (N_3453,N_2041,N_2207);
nand U3454 (N_3454,N_2771,N_2919);
nand U3455 (N_3455,N_2405,N_2780);
nand U3456 (N_3456,N_2010,N_2486);
nor U3457 (N_3457,N_2322,N_2071);
nand U3458 (N_3458,N_2921,N_2838);
nor U3459 (N_3459,N_2642,N_2482);
nand U3460 (N_3460,N_2511,N_2085);
nor U3461 (N_3461,N_2648,N_2943);
nand U3462 (N_3462,N_2371,N_2507);
nor U3463 (N_3463,N_2134,N_2090);
and U3464 (N_3464,N_2818,N_2152);
and U3465 (N_3465,N_2148,N_2740);
nand U3466 (N_3466,N_2348,N_2687);
and U3467 (N_3467,N_2920,N_2582);
or U3468 (N_3468,N_2316,N_2876);
nor U3469 (N_3469,N_2805,N_2518);
nand U3470 (N_3470,N_2113,N_2901);
nor U3471 (N_3471,N_2162,N_2055);
xor U3472 (N_3472,N_2396,N_2625);
nor U3473 (N_3473,N_2290,N_2020);
or U3474 (N_3474,N_2026,N_2646);
or U3475 (N_3475,N_2252,N_2530);
and U3476 (N_3476,N_2455,N_2963);
and U3477 (N_3477,N_2233,N_2232);
nor U3478 (N_3478,N_2934,N_2550);
nand U3479 (N_3479,N_2707,N_2144);
or U3480 (N_3480,N_2663,N_2700);
nor U3481 (N_3481,N_2256,N_2523);
or U3482 (N_3482,N_2406,N_2866);
or U3483 (N_3483,N_2816,N_2437);
and U3484 (N_3484,N_2628,N_2949);
and U3485 (N_3485,N_2670,N_2150);
and U3486 (N_3486,N_2654,N_2791);
or U3487 (N_3487,N_2078,N_2747);
nand U3488 (N_3488,N_2810,N_2696);
or U3489 (N_3489,N_2028,N_2827);
nor U3490 (N_3490,N_2741,N_2987);
and U3491 (N_3491,N_2723,N_2445);
nor U3492 (N_3492,N_2694,N_2386);
and U3493 (N_3493,N_2772,N_2494);
or U3494 (N_3494,N_2245,N_2688);
and U3495 (N_3495,N_2212,N_2653);
or U3496 (N_3496,N_2103,N_2937);
nand U3497 (N_3497,N_2786,N_2275);
nand U3498 (N_3498,N_2727,N_2231);
nand U3499 (N_3499,N_2194,N_2958);
nor U3500 (N_3500,N_2711,N_2868);
or U3501 (N_3501,N_2860,N_2814);
or U3502 (N_3502,N_2197,N_2419);
nor U3503 (N_3503,N_2964,N_2683);
nor U3504 (N_3504,N_2753,N_2619);
nand U3505 (N_3505,N_2428,N_2620);
and U3506 (N_3506,N_2843,N_2080);
or U3507 (N_3507,N_2051,N_2137);
or U3508 (N_3508,N_2895,N_2974);
nand U3509 (N_3509,N_2836,N_2802);
nand U3510 (N_3510,N_2343,N_2160);
and U3511 (N_3511,N_2044,N_2997);
nor U3512 (N_3512,N_2703,N_2811);
nor U3513 (N_3513,N_2762,N_2299);
and U3514 (N_3514,N_2928,N_2527);
or U3515 (N_3515,N_2173,N_2935);
nand U3516 (N_3516,N_2532,N_2874);
nor U3517 (N_3517,N_2412,N_2530);
nor U3518 (N_3518,N_2312,N_2037);
nand U3519 (N_3519,N_2074,N_2265);
nand U3520 (N_3520,N_2554,N_2379);
nor U3521 (N_3521,N_2474,N_2135);
nor U3522 (N_3522,N_2149,N_2240);
nor U3523 (N_3523,N_2850,N_2977);
and U3524 (N_3524,N_2210,N_2642);
or U3525 (N_3525,N_2406,N_2214);
or U3526 (N_3526,N_2377,N_2181);
nor U3527 (N_3527,N_2458,N_2070);
and U3528 (N_3528,N_2465,N_2335);
and U3529 (N_3529,N_2791,N_2490);
and U3530 (N_3530,N_2761,N_2752);
nand U3531 (N_3531,N_2388,N_2695);
and U3532 (N_3532,N_2640,N_2524);
and U3533 (N_3533,N_2390,N_2855);
or U3534 (N_3534,N_2720,N_2649);
and U3535 (N_3535,N_2056,N_2878);
nor U3536 (N_3536,N_2716,N_2134);
nor U3537 (N_3537,N_2603,N_2502);
or U3538 (N_3538,N_2889,N_2683);
and U3539 (N_3539,N_2976,N_2349);
or U3540 (N_3540,N_2220,N_2263);
or U3541 (N_3541,N_2982,N_2369);
nor U3542 (N_3542,N_2331,N_2037);
and U3543 (N_3543,N_2430,N_2679);
and U3544 (N_3544,N_2447,N_2842);
or U3545 (N_3545,N_2266,N_2042);
and U3546 (N_3546,N_2235,N_2826);
nand U3547 (N_3547,N_2916,N_2921);
and U3548 (N_3548,N_2769,N_2860);
and U3549 (N_3549,N_2151,N_2947);
or U3550 (N_3550,N_2684,N_2094);
and U3551 (N_3551,N_2517,N_2552);
nor U3552 (N_3552,N_2667,N_2115);
or U3553 (N_3553,N_2391,N_2751);
and U3554 (N_3554,N_2512,N_2374);
nor U3555 (N_3555,N_2594,N_2602);
or U3556 (N_3556,N_2903,N_2889);
nor U3557 (N_3557,N_2506,N_2421);
nor U3558 (N_3558,N_2983,N_2693);
or U3559 (N_3559,N_2219,N_2422);
nor U3560 (N_3560,N_2623,N_2131);
nand U3561 (N_3561,N_2257,N_2859);
nor U3562 (N_3562,N_2047,N_2670);
xor U3563 (N_3563,N_2715,N_2008);
or U3564 (N_3564,N_2979,N_2962);
nor U3565 (N_3565,N_2172,N_2791);
nor U3566 (N_3566,N_2196,N_2793);
and U3567 (N_3567,N_2569,N_2395);
and U3568 (N_3568,N_2186,N_2873);
or U3569 (N_3569,N_2732,N_2873);
nor U3570 (N_3570,N_2783,N_2133);
or U3571 (N_3571,N_2340,N_2893);
or U3572 (N_3572,N_2847,N_2557);
or U3573 (N_3573,N_2993,N_2718);
nand U3574 (N_3574,N_2870,N_2800);
nor U3575 (N_3575,N_2910,N_2130);
or U3576 (N_3576,N_2294,N_2337);
nand U3577 (N_3577,N_2348,N_2831);
nor U3578 (N_3578,N_2149,N_2376);
or U3579 (N_3579,N_2930,N_2155);
nor U3580 (N_3580,N_2905,N_2272);
nand U3581 (N_3581,N_2913,N_2832);
nand U3582 (N_3582,N_2862,N_2725);
nor U3583 (N_3583,N_2391,N_2589);
nor U3584 (N_3584,N_2053,N_2449);
and U3585 (N_3585,N_2748,N_2648);
nand U3586 (N_3586,N_2417,N_2388);
and U3587 (N_3587,N_2778,N_2282);
or U3588 (N_3588,N_2386,N_2626);
and U3589 (N_3589,N_2019,N_2176);
or U3590 (N_3590,N_2341,N_2893);
or U3591 (N_3591,N_2725,N_2496);
nor U3592 (N_3592,N_2137,N_2842);
nor U3593 (N_3593,N_2271,N_2707);
nor U3594 (N_3594,N_2194,N_2423);
or U3595 (N_3595,N_2305,N_2690);
nor U3596 (N_3596,N_2340,N_2447);
nand U3597 (N_3597,N_2510,N_2549);
and U3598 (N_3598,N_2649,N_2098);
and U3599 (N_3599,N_2109,N_2342);
nor U3600 (N_3600,N_2355,N_2476);
or U3601 (N_3601,N_2443,N_2296);
or U3602 (N_3602,N_2393,N_2901);
and U3603 (N_3603,N_2455,N_2721);
or U3604 (N_3604,N_2145,N_2033);
and U3605 (N_3605,N_2219,N_2359);
nand U3606 (N_3606,N_2612,N_2828);
and U3607 (N_3607,N_2363,N_2025);
and U3608 (N_3608,N_2241,N_2421);
or U3609 (N_3609,N_2149,N_2745);
and U3610 (N_3610,N_2126,N_2320);
and U3611 (N_3611,N_2065,N_2880);
nor U3612 (N_3612,N_2277,N_2306);
and U3613 (N_3613,N_2851,N_2870);
nor U3614 (N_3614,N_2759,N_2037);
or U3615 (N_3615,N_2373,N_2379);
nand U3616 (N_3616,N_2396,N_2827);
nor U3617 (N_3617,N_2389,N_2569);
nand U3618 (N_3618,N_2730,N_2969);
nor U3619 (N_3619,N_2409,N_2999);
nor U3620 (N_3620,N_2071,N_2697);
nor U3621 (N_3621,N_2791,N_2288);
nand U3622 (N_3622,N_2089,N_2527);
xnor U3623 (N_3623,N_2000,N_2382);
nand U3624 (N_3624,N_2331,N_2720);
or U3625 (N_3625,N_2881,N_2553);
or U3626 (N_3626,N_2240,N_2191);
nand U3627 (N_3627,N_2250,N_2532);
and U3628 (N_3628,N_2344,N_2889);
and U3629 (N_3629,N_2497,N_2770);
or U3630 (N_3630,N_2934,N_2688);
nand U3631 (N_3631,N_2550,N_2355);
or U3632 (N_3632,N_2390,N_2741);
nand U3633 (N_3633,N_2868,N_2603);
nand U3634 (N_3634,N_2797,N_2565);
nor U3635 (N_3635,N_2182,N_2725);
or U3636 (N_3636,N_2374,N_2966);
nand U3637 (N_3637,N_2027,N_2445);
nand U3638 (N_3638,N_2942,N_2992);
nand U3639 (N_3639,N_2356,N_2306);
nand U3640 (N_3640,N_2179,N_2911);
nor U3641 (N_3641,N_2875,N_2965);
nand U3642 (N_3642,N_2342,N_2892);
or U3643 (N_3643,N_2720,N_2845);
nor U3644 (N_3644,N_2533,N_2670);
nor U3645 (N_3645,N_2984,N_2378);
or U3646 (N_3646,N_2561,N_2645);
nand U3647 (N_3647,N_2504,N_2589);
and U3648 (N_3648,N_2604,N_2119);
nand U3649 (N_3649,N_2190,N_2243);
and U3650 (N_3650,N_2219,N_2060);
or U3651 (N_3651,N_2343,N_2982);
nand U3652 (N_3652,N_2623,N_2692);
and U3653 (N_3653,N_2314,N_2776);
nor U3654 (N_3654,N_2394,N_2903);
and U3655 (N_3655,N_2809,N_2236);
nand U3656 (N_3656,N_2949,N_2597);
or U3657 (N_3657,N_2856,N_2875);
nor U3658 (N_3658,N_2408,N_2348);
nand U3659 (N_3659,N_2792,N_2054);
nor U3660 (N_3660,N_2934,N_2988);
or U3661 (N_3661,N_2737,N_2882);
nor U3662 (N_3662,N_2705,N_2444);
nor U3663 (N_3663,N_2398,N_2470);
nand U3664 (N_3664,N_2573,N_2722);
and U3665 (N_3665,N_2785,N_2956);
and U3666 (N_3666,N_2865,N_2683);
nor U3667 (N_3667,N_2947,N_2147);
nor U3668 (N_3668,N_2650,N_2810);
nand U3669 (N_3669,N_2683,N_2370);
xnor U3670 (N_3670,N_2779,N_2634);
nand U3671 (N_3671,N_2893,N_2185);
nand U3672 (N_3672,N_2409,N_2890);
nor U3673 (N_3673,N_2171,N_2798);
or U3674 (N_3674,N_2243,N_2689);
nand U3675 (N_3675,N_2268,N_2765);
nand U3676 (N_3676,N_2879,N_2843);
nand U3677 (N_3677,N_2661,N_2829);
or U3678 (N_3678,N_2722,N_2416);
nand U3679 (N_3679,N_2350,N_2662);
nand U3680 (N_3680,N_2485,N_2810);
nand U3681 (N_3681,N_2732,N_2633);
nand U3682 (N_3682,N_2611,N_2935);
nand U3683 (N_3683,N_2774,N_2618);
nor U3684 (N_3684,N_2879,N_2703);
or U3685 (N_3685,N_2812,N_2730);
nand U3686 (N_3686,N_2508,N_2817);
or U3687 (N_3687,N_2344,N_2530);
and U3688 (N_3688,N_2859,N_2265);
nand U3689 (N_3689,N_2096,N_2668);
nand U3690 (N_3690,N_2311,N_2088);
nand U3691 (N_3691,N_2034,N_2909);
nor U3692 (N_3692,N_2126,N_2484);
or U3693 (N_3693,N_2032,N_2363);
nand U3694 (N_3694,N_2890,N_2021);
nand U3695 (N_3695,N_2170,N_2174);
and U3696 (N_3696,N_2920,N_2897);
or U3697 (N_3697,N_2723,N_2976);
nor U3698 (N_3698,N_2809,N_2272);
nor U3699 (N_3699,N_2042,N_2776);
nor U3700 (N_3700,N_2532,N_2974);
xnor U3701 (N_3701,N_2142,N_2474);
or U3702 (N_3702,N_2696,N_2930);
and U3703 (N_3703,N_2941,N_2719);
or U3704 (N_3704,N_2560,N_2451);
or U3705 (N_3705,N_2175,N_2969);
nor U3706 (N_3706,N_2065,N_2953);
and U3707 (N_3707,N_2288,N_2065);
nor U3708 (N_3708,N_2720,N_2575);
or U3709 (N_3709,N_2277,N_2998);
nand U3710 (N_3710,N_2514,N_2486);
and U3711 (N_3711,N_2593,N_2713);
nand U3712 (N_3712,N_2138,N_2827);
and U3713 (N_3713,N_2527,N_2342);
or U3714 (N_3714,N_2264,N_2064);
and U3715 (N_3715,N_2872,N_2351);
and U3716 (N_3716,N_2911,N_2006);
nor U3717 (N_3717,N_2367,N_2264);
or U3718 (N_3718,N_2518,N_2690);
nand U3719 (N_3719,N_2033,N_2962);
or U3720 (N_3720,N_2295,N_2756);
nand U3721 (N_3721,N_2596,N_2455);
nor U3722 (N_3722,N_2896,N_2511);
or U3723 (N_3723,N_2378,N_2300);
nor U3724 (N_3724,N_2269,N_2442);
or U3725 (N_3725,N_2169,N_2672);
or U3726 (N_3726,N_2714,N_2972);
and U3727 (N_3727,N_2037,N_2819);
nand U3728 (N_3728,N_2437,N_2671);
nand U3729 (N_3729,N_2860,N_2462);
nand U3730 (N_3730,N_2452,N_2209);
and U3731 (N_3731,N_2723,N_2519);
and U3732 (N_3732,N_2146,N_2953);
or U3733 (N_3733,N_2173,N_2805);
and U3734 (N_3734,N_2835,N_2978);
nand U3735 (N_3735,N_2940,N_2970);
and U3736 (N_3736,N_2701,N_2131);
or U3737 (N_3737,N_2233,N_2520);
or U3738 (N_3738,N_2358,N_2169);
nor U3739 (N_3739,N_2957,N_2320);
nor U3740 (N_3740,N_2093,N_2021);
nor U3741 (N_3741,N_2366,N_2726);
and U3742 (N_3742,N_2236,N_2209);
nand U3743 (N_3743,N_2707,N_2628);
and U3744 (N_3744,N_2829,N_2071);
xnor U3745 (N_3745,N_2829,N_2781);
nor U3746 (N_3746,N_2906,N_2598);
or U3747 (N_3747,N_2961,N_2212);
nand U3748 (N_3748,N_2864,N_2098);
and U3749 (N_3749,N_2049,N_2725);
and U3750 (N_3750,N_2605,N_2609);
or U3751 (N_3751,N_2894,N_2367);
nor U3752 (N_3752,N_2850,N_2227);
and U3753 (N_3753,N_2866,N_2478);
or U3754 (N_3754,N_2157,N_2803);
nor U3755 (N_3755,N_2682,N_2295);
nor U3756 (N_3756,N_2009,N_2907);
and U3757 (N_3757,N_2355,N_2951);
and U3758 (N_3758,N_2459,N_2560);
nor U3759 (N_3759,N_2755,N_2329);
or U3760 (N_3760,N_2346,N_2566);
nand U3761 (N_3761,N_2076,N_2496);
and U3762 (N_3762,N_2729,N_2765);
nor U3763 (N_3763,N_2160,N_2715);
xnor U3764 (N_3764,N_2938,N_2342);
and U3765 (N_3765,N_2574,N_2886);
or U3766 (N_3766,N_2956,N_2949);
nand U3767 (N_3767,N_2026,N_2918);
or U3768 (N_3768,N_2482,N_2306);
nor U3769 (N_3769,N_2297,N_2551);
and U3770 (N_3770,N_2097,N_2518);
nand U3771 (N_3771,N_2594,N_2147);
and U3772 (N_3772,N_2778,N_2312);
or U3773 (N_3773,N_2452,N_2618);
nand U3774 (N_3774,N_2234,N_2995);
nor U3775 (N_3775,N_2816,N_2481);
nand U3776 (N_3776,N_2666,N_2865);
or U3777 (N_3777,N_2726,N_2100);
nor U3778 (N_3778,N_2536,N_2124);
nor U3779 (N_3779,N_2463,N_2662);
nand U3780 (N_3780,N_2925,N_2203);
nand U3781 (N_3781,N_2744,N_2078);
nand U3782 (N_3782,N_2339,N_2333);
nor U3783 (N_3783,N_2458,N_2571);
nor U3784 (N_3784,N_2444,N_2666);
and U3785 (N_3785,N_2063,N_2049);
nor U3786 (N_3786,N_2606,N_2046);
xor U3787 (N_3787,N_2818,N_2732);
or U3788 (N_3788,N_2184,N_2087);
nor U3789 (N_3789,N_2846,N_2464);
nand U3790 (N_3790,N_2142,N_2502);
nand U3791 (N_3791,N_2931,N_2725);
nor U3792 (N_3792,N_2876,N_2235);
or U3793 (N_3793,N_2523,N_2685);
and U3794 (N_3794,N_2213,N_2970);
xnor U3795 (N_3795,N_2551,N_2782);
nand U3796 (N_3796,N_2071,N_2194);
nor U3797 (N_3797,N_2539,N_2476);
xor U3798 (N_3798,N_2360,N_2153);
or U3799 (N_3799,N_2616,N_2254);
or U3800 (N_3800,N_2172,N_2567);
nor U3801 (N_3801,N_2309,N_2235);
nand U3802 (N_3802,N_2236,N_2890);
and U3803 (N_3803,N_2928,N_2608);
xnor U3804 (N_3804,N_2573,N_2248);
nor U3805 (N_3805,N_2456,N_2568);
and U3806 (N_3806,N_2022,N_2688);
nand U3807 (N_3807,N_2374,N_2933);
and U3808 (N_3808,N_2909,N_2586);
nand U3809 (N_3809,N_2621,N_2573);
and U3810 (N_3810,N_2759,N_2928);
nor U3811 (N_3811,N_2869,N_2636);
nor U3812 (N_3812,N_2943,N_2609);
and U3813 (N_3813,N_2983,N_2617);
nand U3814 (N_3814,N_2889,N_2201);
and U3815 (N_3815,N_2735,N_2107);
xor U3816 (N_3816,N_2110,N_2605);
nor U3817 (N_3817,N_2265,N_2504);
nor U3818 (N_3818,N_2738,N_2540);
xnor U3819 (N_3819,N_2347,N_2689);
or U3820 (N_3820,N_2496,N_2665);
nand U3821 (N_3821,N_2968,N_2670);
and U3822 (N_3822,N_2910,N_2774);
nor U3823 (N_3823,N_2395,N_2178);
or U3824 (N_3824,N_2524,N_2822);
nand U3825 (N_3825,N_2276,N_2856);
and U3826 (N_3826,N_2909,N_2305);
nor U3827 (N_3827,N_2931,N_2058);
nor U3828 (N_3828,N_2560,N_2384);
nor U3829 (N_3829,N_2826,N_2782);
xor U3830 (N_3830,N_2783,N_2049);
and U3831 (N_3831,N_2735,N_2603);
and U3832 (N_3832,N_2968,N_2690);
nand U3833 (N_3833,N_2982,N_2212);
and U3834 (N_3834,N_2370,N_2386);
and U3835 (N_3835,N_2970,N_2150);
nand U3836 (N_3836,N_2108,N_2647);
and U3837 (N_3837,N_2860,N_2708);
nand U3838 (N_3838,N_2306,N_2059);
nand U3839 (N_3839,N_2733,N_2050);
and U3840 (N_3840,N_2934,N_2931);
nor U3841 (N_3841,N_2818,N_2262);
nand U3842 (N_3842,N_2106,N_2922);
and U3843 (N_3843,N_2590,N_2655);
or U3844 (N_3844,N_2687,N_2501);
and U3845 (N_3845,N_2001,N_2089);
nor U3846 (N_3846,N_2497,N_2485);
and U3847 (N_3847,N_2635,N_2254);
xor U3848 (N_3848,N_2286,N_2272);
nand U3849 (N_3849,N_2934,N_2913);
nand U3850 (N_3850,N_2683,N_2088);
nand U3851 (N_3851,N_2217,N_2271);
nor U3852 (N_3852,N_2304,N_2413);
or U3853 (N_3853,N_2104,N_2090);
or U3854 (N_3854,N_2135,N_2870);
nor U3855 (N_3855,N_2584,N_2671);
or U3856 (N_3856,N_2704,N_2332);
nor U3857 (N_3857,N_2238,N_2672);
nor U3858 (N_3858,N_2857,N_2258);
and U3859 (N_3859,N_2625,N_2249);
and U3860 (N_3860,N_2409,N_2581);
and U3861 (N_3861,N_2157,N_2694);
or U3862 (N_3862,N_2487,N_2595);
nor U3863 (N_3863,N_2996,N_2180);
nor U3864 (N_3864,N_2955,N_2678);
or U3865 (N_3865,N_2999,N_2562);
or U3866 (N_3866,N_2636,N_2542);
nand U3867 (N_3867,N_2633,N_2411);
nor U3868 (N_3868,N_2344,N_2944);
nand U3869 (N_3869,N_2926,N_2783);
nor U3870 (N_3870,N_2981,N_2741);
nand U3871 (N_3871,N_2664,N_2976);
nor U3872 (N_3872,N_2960,N_2567);
and U3873 (N_3873,N_2669,N_2785);
nor U3874 (N_3874,N_2949,N_2927);
or U3875 (N_3875,N_2780,N_2997);
or U3876 (N_3876,N_2011,N_2847);
nand U3877 (N_3877,N_2735,N_2211);
or U3878 (N_3878,N_2016,N_2034);
nor U3879 (N_3879,N_2026,N_2228);
and U3880 (N_3880,N_2112,N_2922);
and U3881 (N_3881,N_2053,N_2085);
nor U3882 (N_3882,N_2332,N_2135);
or U3883 (N_3883,N_2116,N_2903);
and U3884 (N_3884,N_2801,N_2654);
nand U3885 (N_3885,N_2083,N_2499);
and U3886 (N_3886,N_2756,N_2144);
nand U3887 (N_3887,N_2830,N_2755);
nand U3888 (N_3888,N_2311,N_2242);
and U3889 (N_3889,N_2769,N_2281);
and U3890 (N_3890,N_2080,N_2352);
and U3891 (N_3891,N_2816,N_2777);
or U3892 (N_3892,N_2376,N_2719);
nand U3893 (N_3893,N_2940,N_2523);
nand U3894 (N_3894,N_2715,N_2630);
or U3895 (N_3895,N_2660,N_2079);
and U3896 (N_3896,N_2868,N_2907);
nand U3897 (N_3897,N_2472,N_2846);
nand U3898 (N_3898,N_2182,N_2820);
or U3899 (N_3899,N_2310,N_2935);
nor U3900 (N_3900,N_2729,N_2863);
nor U3901 (N_3901,N_2766,N_2084);
or U3902 (N_3902,N_2526,N_2730);
or U3903 (N_3903,N_2638,N_2972);
and U3904 (N_3904,N_2133,N_2411);
and U3905 (N_3905,N_2376,N_2079);
nor U3906 (N_3906,N_2159,N_2397);
nor U3907 (N_3907,N_2698,N_2132);
nor U3908 (N_3908,N_2009,N_2927);
nand U3909 (N_3909,N_2584,N_2201);
and U3910 (N_3910,N_2901,N_2011);
and U3911 (N_3911,N_2599,N_2557);
nor U3912 (N_3912,N_2526,N_2483);
or U3913 (N_3913,N_2110,N_2292);
nor U3914 (N_3914,N_2436,N_2741);
nand U3915 (N_3915,N_2296,N_2692);
or U3916 (N_3916,N_2918,N_2946);
and U3917 (N_3917,N_2797,N_2666);
and U3918 (N_3918,N_2705,N_2566);
and U3919 (N_3919,N_2804,N_2167);
nand U3920 (N_3920,N_2928,N_2707);
nor U3921 (N_3921,N_2212,N_2269);
nor U3922 (N_3922,N_2443,N_2467);
or U3923 (N_3923,N_2679,N_2416);
or U3924 (N_3924,N_2000,N_2907);
nand U3925 (N_3925,N_2826,N_2131);
or U3926 (N_3926,N_2795,N_2609);
or U3927 (N_3927,N_2681,N_2537);
and U3928 (N_3928,N_2429,N_2745);
and U3929 (N_3929,N_2872,N_2021);
xnor U3930 (N_3930,N_2490,N_2511);
nand U3931 (N_3931,N_2518,N_2804);
nand U3932 (N_3932,N_2414,N_2017);
or U3933 (N_3933,N_2222,N_2095);
and U3934 (N_3934,N_2069,N_2727);
xnor U3935 (N_3935,N_2305,N_2147);
xnor U3936 (N_3936,N_2979,N_2233);
or U3937 (N_3937,N_2192,N_2890);
nor U3938 (N_3938,N_2448,N_2189);
nand U3939 (N_3939,N_2686,N_2832);
nor U3940 (N_3940,N_2244,N_2013);
and U3941 (N_3941,N_2404,N_2789);
nand U3942 (N_3942,N_2197,N_2156);
and U3943 (N_3943,N_2626,N_2802);
or U3944 (N_3944,N_2958,N_2660);
or U3945 (N_3945,N_2567,N_2228);
and U3946 (N_3946,N_2335,N_2471);
nand U3947 (N_3947,N_2265,N_2562);
and U3948 (N_3948,N_2154,N_2338);
nor U3949 (N_3949,N_2533,N_2879);
nand U3950 (N_3950,N_2969,N_2695);
nor U3951 (N_3951,N_2589,N_2831);
or U3952 (N_3952,N_2066,N_2354);
and U3953 (N_3953,N_2883,N_2627);
and U3954 (N_3954,N_2922,N_2373);
or U3955 (N_3955,N_2706,N_2477);
nor U3956 (N_3956,N_2552,N_2314);
and U3957 (N_3957,N_2307,N_2280);
or U3958 (N_3958,N_2434,N_2647);
nor U3959 (N_3959,N_2868,N_2630);
nor U3960 (N_3960,N_2168,N_2766);
or U3961 (N_3961,N_2615,N_2440);
nor U3962 (N_3962,N_2911,N_2684);
or U3963 (N_3963,N_2613,N_2749);
nor U3964 (N_3964,N_2032,N_2485);
or U3965 (N_3965,N_2529,N_2720);
and U3966 (N_3966,N_2775,N_2031);
or U3967 (N_3967,N_2987,N_2067);
nor U3968 (N_3968,N_2905,N_2775);
or U3969 (N_3969,N_2009,N_2040);
nand U3970 (N_3970,N_2445,N_2505);
or U3971 (N_3971,N_2538,N_2712);
and U3972 (N_3972,N_2935,N_2270);
nor U3973 (N_3973,N_2672,N_2717);
or U3974 (N_3974,N_2909,N_2463);
nand U3975 (N_3975,N_2280,N_2125);
or U3976 (N_3976,N_2727,N_2112);
and U3977 (N_3977,N_2451,N_2797);
nor U3978 (N_3978,N_2264,N_2998);
or U3979 (N_3979,N_2802,N_2269);
nor U3980 (N_3980,N_2171,N_2448);
and U3981 (N_3981,N_2372,N_2918);
nand U3982 (N_3982,N_2010,N_2911);
and U3983 (N_3983,N_2485,N_2010);
or U3984 (N_3984,N_2893,N_2921);
nor U3985 (N_3985,N_2607,N_2714);
or U3986 (N_3986,N_2345,N_2174);
and U3987 (N_3987,N_2520,N_2742);
and U3988 (N_3988,N_2025,N_2592);
nor U3989 (N_3989,N_2853,N_2537);
and U3990 (N_3990,N_2564,N_2560);
nor U3991 (N_3991,N_2019,N_2502);
nor U3992 (N_3992,N_2589,N_2017);
nand U3993 (N_3993,N_2798,N_2861);
xor U3994 (N_3994,N_2575,N_2114);
nand U3995 (N_3995,N_2911,N_2564);
nor U3996 (N_3996,N_2620,N_2340);
nand U3997 (N_3997,N_2927,N_2386);
and U3998 (N_3998,N_2367,N_2284);
nand U3999 (N_3999,N_2529,N_2107);
or U4000 (N_4000,N_3174,N_3779);
and U4001 (N_4001,N_3180,N_3326);
nor U4002 (N_4002,N_3507,N_3784);
nor U4003 (N_4003,N_3868,N_3246);
nor U4004 (N_4004,N_3707,N_3661);
and U4005 (N_4005,N_3242,N_3215);
or U4006 (N_4006,N_3420,N_3586);
nor U4007 (N_4007,N_3184,N_3310);
or U4008 (N_4008,N_3293,N_3378);
nand U4009 (N_4009,N_3013,N_3313);
and U4010 (N_4010,N_3706,N_3190);
nor U4011 (N_4011,N_3883,N_3499);
nand U4012 (N_4012,N_3544,N_3773);
or U4013 (N_4013,N_3510,N_3672);
or U4014 (N_4014,N_3280,N_3655);
or U4015 (N_4015,N_3135,N_3537);
or U4016 (N_4016,N_3610,N_3910);
nand U4017 (N_4017,N_3475,N_3627);
and U4018 (N_4018,N_3723,N_3011);
and U4019 (N_4019,N_3120,N_3224);
or U4020 (N_4020,N_3940,N_3423);
and U4021 (N_4021,N_3817,N_3907);
nand U4022 (N_4022,N_3097,N_3149);
nand U4023 (N_4023,N_3440,N_3838);
or U4024 (N_4024,N_3298,N_3702);
or U4025 (N_4025,N_3249,N_3799);
nand U4026 (N_4026,N_3680,N_3696);
or U4027 (N_4027,N_3901,N_3018);
and U4028 (N_4028,N_3296,N_3049);
and U4029 (N_4029,N_3364,N_3098);
nand U4030 (N_4030,N_3549,N_3558);
or U4031 (N_4031,N_3321,N_3769);
and U4032 (N_4032,N_3593,N_3287);
and U4033 (N_4033,N_3487,N_3887);
and U4034 (N_4034,N_3162,N_3413);
nor U4035 (N_4035,N_3330,N_3971);
nor U4036 (N_4036,N_3419,N_3976);
and U4037 (N_4037,N_3067,N_3460);
nand U4038 (N_4038,N_3917,N_3704);
and U4039 (N_4039,N_3875,N_3343);
nor U4040 (N_4040,N_3541,N_3151);
or U4041 (N_4041,N_3990,N_3227);
or U4042 (N_4042,N_3152,N_3676);
nand U4043 (N_4043,N_3922,N_3974);
or U4044 (N_4044,N_3625,N_3979);
and U4045 (N_4045,N_3456,N_3466);
nand U4046 (N_4046,N_3240,N_3041);
xor U4047 (N_4047,N_3303,N_3134);
xnor U4048 (N_4048,N_3394,N_3520);
and U4049 (N_4049,N_3618,N_3830);
nand U4050 (N_4050,N_3569,N_3252);
or U4051 (N_4051,N_3919,N_3764);
nand U4052 (N_4052,N_3128,N_3412);
and U4053 (N_4053,N_3457,N_3436);
and U4054 (N_4054,N_3331,N_3027);
or U4055 (N_4055,N_3775,N_3344);
nor U4056 (N_4056,N_3671,N_3173);
and U4057 (N_4057,N_3991,N_3847);
nand U4058 (N_4058,N_3103,N_3845);
nand U4059 (N_4059,N_3122,N_3382);
nand U4060 (N_4060,N_3973,N_3984);
nand U4061 (N_4061,N_3898,N_3894);
or U4062 (N_4062,N_3132,N_3709);
nor U4063 (N_4063,N_3124,N_3346);
nor U4064 (N_4064,N_3908,N_3309);
nor U4065 (N_4065,N_3892,N_3731);
nor U4066 (N_4066,N_3725,N_3471);
and U4067 (N_4067,N_3599,N_3981);
or U4068 (N_4068,N_3074,N_3719);
nor U4069 (N_4069,N_3634,N_3489);
and U4070 (N_4070,N_3673,N_3038);
and U4071 (N_4071,N_3685,N_3031);
or U4072 (N_4072,N_3314,N_3464);
nand U4073 (N_4073,N_3588,N_3029);
and U4074 (N_4074,N_3145,N_3543);
and U4075 (N_4075,N_3862,N_3708);
and U4076 (N_4076,N_3159,N_3563);
or U4077 (N_4077,N_3010,N_3664);
or U4078 (N_4078,N_3478,N_3276);
and U4079 (N_4079,N_3086,N_3484);
or U4080 (N_4080,N_3051,N_3161);
nand U4081 (N_4081,N_3465,N_3737);
nor U4082 (N_4082,N_3131,N_3866);
and U4083 (N_4083,N_3800,N_3669);
or U4084 (N_4084,N_3636,N_3444);
or U4085 (N_4085,N_3983,N_3207);
nand U4086 (N_4086,N_3283,N_3656);
nor U4087 (N_4087,N_3753,N_3076);
nand U4088 (N_4088,N_3323,N_3893);
nor U4089 (N_4089,N_3441,N_3209);
nand U4090 (N_4090,N_3886,N_3720);
nand U4091 (N_4091,N_3951,N_3823);
and U4092 (N_4092,N_3089,N_3579);
nand U4093 (N_4093,N_3325,N_3212);
and U4094 (N_4094,N_3975,N_3153);
nand U4095 (N_4095,N_3551,N_3062);
or U4096 (N_4096,N_3175,N_3552);
and U4097 (N_4097,N_3793,N_3117);
and U4098 (N_4098,N_3196,N_3649);
or U4099 (N_4099,N_3009,N_3306);
xnor U4100 (N_4100,N_3626,N_3255);
and U4101 (N_4101,N_3926,N_3026);
nor U4102 (N_4102,N_3597,N_3547);
and U4103 (N_4103,N_3874,N_3002);
or U4104 (N_4104,N_3424,N_3949);
xor U4105 (N_4105,N_3494,N_3366);
or U4106 (N_4106,N_3872,N_3846);
or U4107 (N_4107,N_3241,N_3824);
nor U4108 (N_4108,N_3046,N_3305);
and U4109 (N_4109,N_3234,N_3607);
nor U4110 (N_4110,N_3019,N_3477);
nor U4111 (N_4111,N_3654,N_3495);
or U4112 (N_4112,N_3094,N_3187);
nand U4113 (N_4113,N_3534,N_3396);
nor U4114 (N_4114,N_3197,N_3929);
or U4115 (N_4115,N_3311,N_3994);
or U4116 (N_4116,N_3783,N_3788);
nor U4117 (N_4117,N_3090,N_3611);
nand U4118 (N_4118,N_3904,N_3210);
nor U4119 (N_4119,N_3329,N_3055);
or U4120 (N_4120,N_3913,N_3623);
nand U4121 (N_4121,N_3455,N_3877);
or U4122 (N_4122,N_3127,N_3256);
and U4123 (N_4123,N_3759,N_3405);
or U4124 (N_4124,N_3250,N_3577);
nor U4125 (N_4125,N_3622,N_3620);
or U4126 (N_4126,N_3641,N_3275);
and U4127 (N_4127,N_3039,N_3550);
nor U4128 (N_4128,N_3267,N_3107);
nor U4129 (N_4129,N_3400,N_3679);
and U4130 (N_4130,N_3934,N_3591);
nor U4131 (N_4131,N_3381,N_3531);
and U4132 (N_4132,N_3884,N_3065);
and U4133 (N_4133,N_3048,N_3452);
or U4134 (N_4134,N_3570,N_3142);
and U4135 (N_4135,N_3658,N_3372);
or U4136 (N_4136,N_3938,N_3269);
nand U4137 (N_4137,N_3118,N_3391);
and U4138 (N_4138,N_3512,N_3492);
nand U4139 (N_4139,N_3485,N_3431);
or U4140 (N_4140,N_3113,N_3063);
or U4141 (N_4141,N_3612,N_3722);
nor U4142 (N_4142,N_3081,N_3223);
or U4143 (N_4143,N_3402,N_3843);
or U4144 (N_4144,N_3491,N_3189);
nor U4145 (N_4145,N_3941,N_3606);
nand U4146 (N_4146,N_3980,N_3746);
nand U4147 (N_4147,N_3615,N_3932);
nand U4148 (N_4148,N_3384,N_3699);
nor U4149 (N_4149,N_3944,N_3416);
and U4150 (N_4150,N_3965,N_3853);
or U4151 (N_4151,N_3802,N_3380);
xor U4152 (N_4152,N_3070,N_3827);
nand U4153 (N_4153,N_3337,N_3479);
nor U4154 (N_4154,N_3933,N_3012);
nand U4155 (N_4155,N_3168,N_3792);
nand U4156 (N_4156,N_3397,N_3272);
nor U4157 (N_4157,N_3590,N_3312);
nand U4158 (N_4158,N_3459,N_3101);
or U4159 (N_4159,N_3871,N_3835);
nand U4160 (N_4160,N_3342,N_3849);
nor U4161 (N_4161,N_3756,N_3740);
or U4162 (N_4162,N_3542,N_3767);
or U4163 (N_4163,N_3624,N_3301);
or U4164 (N_4164,N_3111,N_3943);
xnor U4165 (N_4165,N_3273,N_3995);
or U4166 (N_4166,N_3408,N_3203);
nor U4167 (N_4167,N_3829,N_3840);
nor U4168 (N_4168,N_3185,N_3748);
nor U4169 (N_4169,N_3595,N_3750);
nand U4170 (N_4170,N_3855,N_3869);
nor U4171 (N_4171,N_3523,N_3468);
nand U4172 (N_4172,N_3996,N_3739);
nand U4173 (N_4173,N_3890,N_3208);
or U4174 (N_4174,N_3566,N_3476);
or U4175 (N_4175,N_3682,N_3059);
and U4176 (N_4176,N_3870,N_3368);
or U4177 (N_4177,N_3946,N_3918);
and U4178 (N_4178,N_3345,N_3064);
or U4179 (N_4179,N_3515,N_3742);
and U4180 (N_4180,N_3147,N_3714);
or U4181 (N_4181,N_3964,N_3498);
or U4182 (N_4182,N_3474,N_3220);
and U4183 (N_4183,N_3571,N_3473);
and U4184 (N_4184,N_3482,N_3148);
and U4185 (N_4185,N_3832,N_3888);
or U4186 (N_4186,N_3422,N_3506);
or U4187 (N_4187,N_3016,N_3809);
nor U4188 (N_4188,N_3322,N_3916);
or U4189 (N_4189,N_3387,N_3317);
nand U4190 (N_4190,N_3490,N_3072);
and U4191 (N_4191,N_3529,N_3628);
nand U4192 (N_4192,N_3257,N_3229);
and U4193 (N_4193,N_3160,N_3514);
xor U4194 (N_4194,N_3519,N_3294);
nand U4195 (N_4195,N_3297,N_3666);
nand U4196 (N_4196,N_3078,N_3088);
and U4197 (N_4197,N_3896,N_3864);
or U4198 (N_4198,N_3211,N_3677);
nor U4199 (N_4199,N_3967,N_3106);
nor U4200 (N_4200,N_3369,N_3355);
or U4201 (N_4201,N_3822,N_3948);
nor U4202 (N_4202,N_3539,N_3277);
nor U4203 (N_4203,N_3766,N_3760);
or U4204 (N_4204,N_3710,N_3988);
or U4205 (N_4205,N_3966,N_3114);
xor U4206 (N_4206,N_3526,N_3956);
nor U4207 (N_4207,N_3839,N_3998);
and U4208 (N_4208,N_3481,N_3260);
nand U4209 (N_4209,N_3021,N_3808);
nor U4210 (N_4210,N_3540,N_3417);
and U4211 (N_4211,N_3825,N_3375);
nand U4212 (N_4212,N_3504,N_3333);
nor U4213 (N_4213,N_3819,N_3911);
and U4214 (N_4214,N_3613,N_3407);
and U4215 (N_4215,N_3087,N_3365);
and U4216 (N_4216,N_3906,N_3172);
nor U4217 (N_4217,N_3942,N_3925);
or U4218 (N_4218,N_3001,N_3061);
nor U4219 (N_4219,N_3015,N_3797);
nand U4220 (N_4220,N_3259,N_3741);
or U4221 (N_4221,N_3181,N_3388);
nand U4222 (N_4222,N_3583,N_3557);
and U4223 (N_4223,N_3195,N_3617);
and U4224 (N_4224,N_3139,N_3667);
nor U4225 (N_4225,N_3000,N_3379);
nor U4226 (N_4226,N_3360,N_3361);
or U4227 (N_4227,N_3427,N_3865);
nor U4228 (N_4228,N_3598,N_3376);
nor U4229 (N_4229,N_3430,N_3453);
and U4230 (N_4230,N_3036,N_3339);
or U4231 (N_4231,N_3435,N_3828);
and U4232 (N_4232,N_3977,N_3924);
nor U4233 (N_4233,N_3447,N_3768);
and U4234 (N_4234,N_3217,N_3434);
nor U4235 (N_4235,N_3713,N_3497);
and U4236 (N_4236,N_3426,N_3521);
xor U4237 (N_4237,N_3858,N_3262);
or U4238 (N_4238,N_3157,N_3794);
xnor U4239 (N_4239,N_3957,N_3584);
and U4240 (N_4240,N_3581,N_3650);
nand U4241 (N_4241,N_3488,N_3082);
nand U4242 (N_4242,N_3289,N_3804);
or U4243 (N_4243,N_3318,N_3385);
nor U4244 (N_4244,N_3782,N_3616);
or U4245 (N_4245,N_3406,N_3700);
nor U4246 (N_4246,N_3171,N_3528);
nand U4247 (N_4247,N_3660,N_3861);
xor U4248 (N_4248,N_3020,N_3080);
nor U4249 (N_4249,N_3102,N_3561);
or U4250 (N_4250,N_3439,N_3353);
or U4251 (N_4251,N_3263,N_3837);
nor U4252 (N_4252,N_3878,N_3167);
and U4253 (N_4253,N_3638,N_3500);
or U4254 (N_4254,N_3158,N_3221);
nor U4255 (N_4255,N_3633,N_3762);
and U4256 (N_4256,N_3176,N_3023);
nand U4257 (N_4257,N_3282,N_3604);
nand U4258 (N_4258,N_3678,N_3204);
nor U4259 (N_4259,N_3022,N_3787);
and U4260 (N_4260,N_3812,N_3042);
or U4261 (N_4261,N_3692,N_3596);
nand U4262 (N_4262,N_3017,N_3724);
nor U4263 (N_4263,N_3104,N_3445);
or U4264 (N_4264,N_3054,N_3150);
nand U4265 (N_4265,N_3050,N_3693);
and U4266 (N_4266,N_3178,N_3216);
or U4267 (N_4267,N_3774,N_3553);
nor U4268 (N_4268,N_3791,N_3371);
nand U4269 (N_4269,N_3580,N_3469);
nand U4270 (N_4270,N_3047,N_3073);
and U4271 (N_4271,N_3575,N_3032);
nand U4272 (N_4272,N_3589,N_3170);
nor U4273 (N_4273,N_3816,N_3605);
nand U4274 (N_4274,N_3443,N_3686);
and U4275 (N_4275,N_3805,N_3429);
nand U4276 (N_4276,N_3776,N_3527);
nor U4277 (N_4277,N_3806,N_3244);
nor U4278 (N_4278,N_3137,N_3433);
and U4279 (N_4279,N_3645,N_3328);
or U4280 (N_4280,N_3651,N_3729);
or U4281 (N_4281,N_3425,N_3952);
and U4282 (N_4282,N_3218,N_3718);
and U4283 (N_4283,N_3903,N_3136);
or U4284 (N_4284,N_3844,N_3524);
nor U4285 (N_4285,N_3530,N_3790);
nand U4286 (N_4286,N_3014,N_3125);
nand U4287 (N_4287,N_3662,N_3066);
nand U4288 (N_4288,N_3254,N_3997);
nor U4289 (N_4289,N_3505,N_3642);
or U4290 (N_4290,N_3133,N_3327);
and U4291 (N_4291,N_3785,N_3352);
or U4292 (N_4292,N_3228,N_3335);
nand U4293 (N_4293,N_3576,N_3857);
nand U4294 (N_4294,N_3274,N_3268);
or U4295 (N_4295,N_3921,N_3349);
xor U4296 (N_4296,N_3232,N_3694);
and U4297 (N_4297,N_3451,N_3989);
or U4298 (N_4298,N_3084,N_3357);
or U4299 (N_4299,N_3291,N_3535);
and U4300 (N_4300,N_3532,N_3121);
nand U4301 (N_4301,N_3233,N_3186);
and U4302 (N_4302,N_3193,N_3226);
nand U4303 (N_4303,N_3116,N_3603);
and U4304 (N_4304,N_3691,N_3126);
nor U4305 (N_4305,N_3914,N_3467);
nand U4306 (N_4306,N_3115,N_3213);
nand U4307 (N_4307,N_3716,N_3005);
nand U4308 (N_4308,N_3630,N_3960);
or U4309 (N_4309,N_3068,N_3592);
and U4310 (N_4310,N_3177,N_3730);
nand U4311 (N_4311,N_3091,N_3745);
nand U4312 (N_4312,N_3647,N_3545);
nand U4313 (N_4313,N_3567,N_3920);
or U4314 (N_4314,N_3747,N_3214);
or U4315 (N_4315,N_3572,N_3119);
and U4316 (N_4316,N_3744,N_3867);
and U4317 (N_4317,N_3715,N_3814);
or U4318 (N_4318,N_3688,N_3421);
or U4319 (N_4319,N_3736,N_3194);
or U4320 (N_4320,N_3450,N_3334);
nand U4321 (N_4321,N_3155,N_3681);
or U4322 (N_4322,N_3732,N_3554);
or U4323 (N_4323,N_3939,N_3284);
nand U4324 (N_4324,N_3734,N_3992);
nor U4325 (N_4325,N_3961,N_3299);
nor U4326 (N_4326,N_3237,N_3958);
or U4327 (N_4327,N_3045,N_3202);
and U4328 (N_4328,N_3972,N_3290);
and U4329 (N_4329,N_3937,N_3449);
xor U4330 (N_4330,N_3164,N_3689);
or U4331 (N_4331,N_3415,N_3351);
nor U4332 (N_4332,N_3728,N_3144);
and U4333 (N_4333,N_3780,N_3442);
and U4334 (N_4334,N_3235,N_3140);
xor U4335 (N_4335,N_3856,N_3559);
nand U4336 (N_4336,N_3743,N_3945);
or U4337 (N_4337,N_3999,N_3936);
or U4338 (N_4338,N_3205,N_3985);
nand U4339 (N_4339,N_3432,N_3428);
and U4340 (N_4340,N_3850,N_3950);
or U4341 (N_4341,N_3281,N_3876);
nor U4342 (N_4342,N_3698,N_3758);
xor U4343 (N_4343,N_3033,N_3548);
and U4344 (N_4344,N_3796,N_3562);
nand U4345 (N_4345,N_3373,N_3383);
and U4346 (N_4346,N_3880,N_3079);
nand U4347 (N_4347,N_3879,N_3332);
nand U4348 (N_4348,N_3953,N_3286);
nand U4349 (N_4349,N_3600,N_3602);
nor U4350 (N_4350,N_3362,N_3755);
or U4351 (N_4351,N_3789,N_3270);
or U4352 (N_4352,N_3652,N_3927);
nor U4353 (N_4353,N_3993,N_3414);
and U4354 (N_4354,N_3601,N_3219);
nand U4355 (N_4355,N_3462,N_3818);
or U4356 (N_4356,N_3963,N_3644);
or U4357 (N_4357,N_3182,N_3711);
or U4358 (N_4358,N_3508,N_3931);
nor U4359 (N_4359,N_3165,N_3071);
nor U4360 (N_4360,N_3243,N_3037);
or U4361 (N_4361,N_3472,N_3201);
or U4362 (N_4362,N_3771,N_3969);
nor U4363 (N_4363,N_3770,N_3555);
nor U4364 (N_4364,N_3982,N_3821);
nand U4365 (N_4365,N_3619,N_3820);
nand U4366 (N_4366,N_3668,N_3757);
nand U4367 (N_4367,N_3044,N_3188);
and U4368 (N_4368,N_3356,N_3024);
or U4369 (N_4369,N_3859,N_3665);
nor U4370 (N_4370,N_3112,N_3810);
nand U4371 (N_4371,N_3536,N_3986);
or U4372 (N_4372,N_3522,N_3486);
nand U4373 (N_4373,N_3348,N_3848);
or U4374 (N_4374,N_3712,N_3928);
nand U4375 (N_4375,N_3409,N_3860);
nand U4376 (N_4376,N_3034,N_3643);
nand U4377 (N_4377,N_3105,N_3826);
nand U4378 (N_4378,N_3899,N_3721);
nand U4379 (N_4379,N_3110,N_3873);
nor U4380 (N_4380,N_3096,N_3463);
nor U4381 (N_4381,N_3546,N_3253);
or U4382 (N_4382,N_3222,N_3781);
nor U4383 (N_4383,N_3503,N_3653);
or U4384 (N_4384,N_3438,N_3245);
and U4385 (N_4385,N_3803,N_3295);
nand U4386 (N_4386,N_3386,N_3726);
nor U4387 (N_4387,N_3302,N_3836);
nor U4388 (N_4388,N_3754,N_3060);
or U4389 (N_4389,N_3621,N_3261);
nand U4390 (N_4390,N_3889,N_3320);
or U4391 (N_4391,N_3053,N_3513);
nor U4392 (N_4392,N_3639,N_3798);
nand U4393 (N_4393,N_3006,N_3842);
and U4394 (N_4394,N_3518,N_3891);
and U4395 (N_4395,N_3930,N_3959);
nand U4396 (N_4396,N_3377,N_3900);
nor U4397 (N_4397,N_3304,N_3882);
nor U4398 (N_4398,N_3501,N_3568);
nand U4399 (N_4399,N_3483,N_3786);
and U4400 (N_4400,N_3092,N_3565);
nand U4401 (N_4401,N_3717,N_3437);
nor U4402 (N_4402,N_3727,N_3367);
or U4403 (N_4403,N_3265,N_3831);
and U4404 (N_4404,N_3480,N_3030);
nand U4405 (N_4405,N_3292,N_3765);
or U4406 (N_4406,N_3266,N_3278);
or U4407 (N_4407,N_3703,N_3239);
nor U4408 (N_4408,N_3470,N_3003);
nand U4409 (N_4409,N_3493,N_3230);
nand U4410 (N_4410,N_3895,N_3648);
or U4411 (N_4411,N_3285,N_3264);
nand U4412 (N_4412,N_3538,N_3008);
xnor U4413 (N_4413,N_3403,N_3083);
nand U4414 (N_4414,N_3578,N_3683);
nand U4415 (N_4415,N_3594,N_3043);
and U4416 (N_4416,N_3390,N_3347);
or U4417 (N_4417,N_3684,N_3923);
and U4418 (N_4418,N_3517,N_3614);
or U4419 (N_4419,N_3851,N_3251);
nor U4420 (N_4420,N_3813,N_3632);
nor U4421 (N_4421,N_3968,N_3778);
nor U4422 (N_4422,N_3404,N_3815);
or U4423 (N_4423,N_3056,N_3069);
nor U4424 (N_4424,N_3609,N_3947);
or U4425 (N_4425,N_3341,N_3454);
nand U4426 (N_4426,N_3129,N_3978);
nand U4427 (N_4427,N_3040,N_3970);
nor U4428 (N_4428,N_3085,N_3516);
and U4429 (N_4429,N_3733,N_3834);
nor U4430 (N_4430,N_3509,N_3640);
and U4431 (N_4431,N_3247,N_3511);
and U4432 (N_4432,N_3962,N_3659);
and U4433 (N_4433,N_3749,N_3987);
and U4434 (N_4434,N_3279,N_3735);
and U4435 (N_4435,N_3675,N_3763);
nand U4436 (N_4436,N_3752,N_3025);
nor U4437 (N_4437,N_3075,N_3587);
nand U4438 (N_4438,N_3695,N_3881);
nand U4439 (N_4439,N_3663,N_3496);
nor U4440 (N_4440,N_3761,N_3448);
nor U4441 (N_4441,N_3801,N_3183);
and U4442 (N_4442,N_3392,N_3582);
and U4443 (N_4443,N_3004,N_3401);
or U4444 (N_4444,N_3007,N_3143);
and U4445 (N_4445,N_3608,N_3954);
nand U4446 (N_4446,N_3225,N_3350);
or U4447 (N_4447,N_3912,N_3697);
nor U4448 (N_4448,N_3316,N_3411);
nand U4449 (N_4449,N_3095,N_3300);
nand U4450 (N_4450,N_3446,N_3035);
or U4451 (N_4451,N_3169,N_3358);
nor U4452 (N_4452,N_3154,N_3751);
nor U4453 (N_4453,N_3458,N_3093);
nor U4454 (N_4454,N_3108,N_3410);
and U4455 (N_4455,N_3146,N_3585);
nor U4456 (N_4456,N_3374,N_3674);
or U4457 (N_4457,N_3206,N_3885);
and U4458 (N_4458,N_3238,N_3336);
or U4459 (N_4459,N_3123,N_3099);
nor U4460 (N_4460,N_3863,N_3399);
or U4461 (N_4461,N_3258,N_3738);
nand U4462 (N_4462,N_3057,N_3395);
or U4463 (N_4463,N_3166,N_3179);
or U4464 (N_4464,N_3191,N_3690);
nand U4465 (N_4465,N_3198,N_3854);
or U4466 (N_4466,N_3841,N_3109);
nor U4467 (N_4467,N_3955,N_3687);
nor U4468 (N_4468,N_3915,N_3398);
nor U4469 (N_4469,N_3077,N_3338);
nand U4470 (N_4470,N_3288,N_3058);
nand U4471 (N_4471,N_3935,N_3156);
nand U4472 (N_4472,N_3701,N_3130);
nor U4473 (N_4473,N_3833,N_3574);
and U4474 (N_4474,N_3461,N_3271);
nor U4475 (N_4475,N_3141,N_3852);
nand U4476 (N_4476,N_3370,N_3631);
xor U4477 (N_4477,N_3807,N_3200);
xnor U4478 (N_4478,N_3307,N_3705);
or U4479 (N_4479,N_3308,N_3772);
or U4480 (N_4480,N_3248,N_3138);
and U4481 (N_4481,N_3163,N_3028);
and U4482 (N_4482,N_3635,N_3573);
and U4483 (N_4483,N_3670,N_3359);
nor U4484 (N_4484,N_3560,N_3909);
and U4485 (N_4485,N_3389,N_3811);
nor U4486 (N_4486,N_3052,N_3657);
or U4487 (N_4487,N_3556,N_3192);
or U4488 (N_4488,N_3646,N_3525);
or U4489 (N_4489,N_3905,N_3777);
nand U4490 (N_4490,N_3354,N_3393);
nor U4491 (N_4491,N_3315,N_3231);
xnor U4492 (N_4492,N_3319,N_3564);
and U4493 (N_4493,N_3199,N_3324);
and U4494 (N_4494,N_3795,N_3902);
or U4495 (N_4495,N_3100,N_3363);
nor U4496 (N_4496,N_3502,N_3533);
and U4497 (N_4497,N_3637,N_3629);
nand U4498 (N_4498,N_3236,N_3418);
or U4499 (N_4499,N_3897,N_3340);
and U4500 (N_4500,N_3430,N_3227);
or U4501 (N_4501,N_3687,N_3124);
and U4502 (N_4502,N_3845,N_3413);
or U4503 (N_4503,N_3988,N_3540);
and U4504 (N_4504,N_3645,N_3700);
nand U4505 (N_4505,N_3078,N_3691);
and U4506 (N_4506,N_3636,N_3354);
and U4507 (N_4507,N_3215,N_3851);
or U4508 (N_4508,N_3251,N_3859);
and U4509 (N_4509,N_3854,N_3016);
and U4510 (N_4510,N_3486,N_3672);
nor U4511 (N_4511,N_3570,N_3891);
nand U4512 (N_4512,N_3307,N_3197);
or U4513 (N_4513,N_3837,N_3853);
and U4514 (N_4514,N_3799,N_3001);
or U4515 (N_4515,N_3971,N_3195);
nor U4516 (N_4516,N_3942,N_3780);
nand U4517 (N_4517,N_3447,N_3307);
nand U4518 (N_4518,N_3919,N_3387);
or U4519 (N_4519,N_3633,N_3049);
and U4520 (N_4520,N_3545,N_3483);
or U4521 (N_4521,N_3976,N_3492);
nand U4522 (N_4522,N_3322,N_3475);
nand U4523 (N_4523,N_3640,N_3256);
or U4524 (N_4524,N_3298,N_3621);
nand U4525 (N_4525,N_3999,N_3263);
nand U4526 (N_4526,N_3860,N_3313);
nor U4527 (N_4527,N_3928,N_3752);
and U4528 (N_4528,N_3559,N_3351);
and U4529 (N_4529,N_3289,N_3465);
xor U4530 (N_4530,N_3638,N_3786);
or U4531 (N_4531,N_3962,N_3239);
and U4532 (N_4532,N_3107,N_3811);
and U4533 (N_4533,N_3918,N_3486);
and U4534 (N_4534,N_3516,N_3672);
or U4535 (N_4535,N_3734,N_3115);
or U4536 (N_4536,N_3308,N_3409);
or U4537 (N_4537,N_3855,N_3247);
nand U4538 (N_4538,N_3139,N_3002);
nor U4539 (N_4539,N_3337,N_3032);
nor U4540 (N_4540,N_3579,N_3000);
and U4541 (N_4541,N_3551,N_3528);
nand U4542 (N_4542,N_3009,N_3915);
nor U4543 (N_4543,N_3494,N_3034);
or U4544 (N_4544,N_3724,N_3380);
nor U4545 (N_4545,N_3284,N_3120);
nor U4546 (N_4546,N_3975,N_3952);
or U4547 (N_4547,N_3126,N_3889);
nor U4548 (N_4548,N_3427,N_3337);
nor U4549 (N_4549,N_3942,N_3997);
and U4550 (N_4550,N_3321,N_3211);
and U4551 (N_4551,N_3767,N_3586);
nor U4552 (N_4552,N_3512,N_3468);
nand U4553 (N_4553,N_3233,N_3316);
nand U4554 (N_4554,N_3379,N_3817);
and U4555 (N_4555,N_3491,N_3026);
nand U4556 (N_4556,N_3996,N_3532);
nand U4557 (N_4557,N_3757,N_3387);
xnor U4558 (N_4558,N_3963,N_3371);
nor U4559 (N_4559,N_3908,N_3491);
nand U4560 (N_4560,N_3129,N_3803);
or U4561 (N_4561,N_3660,N_3450);
nand U4562 (N_4562,N_3121,N_3641);
or U4563 (N_4563,N_3879,N_3087);
nand U4564 (N_4564,N_3471,N_3981);
and U4565 (N_4565,N_3578,N_3524);
or U4566 (N_4566,N_3275,N_3639);
or U4567 (N_4567,N_3513,N_3283);
xnor U4568 (N_4568,N_3148,N_3328);
nand U4569 (N_4569,N_3267,N_3995);
and U4570 (N_4570,N_3075,N_3179);
or U4571 (N_4571,N_3091,N_3176);
nor U4572 (N_4572,N_3478,N_3201);
nand U4573 (N_4573,N_3606,N_3251);
or U4574 (N_4574,N_3088,N_3999);
nand U4575 (N_4575,N_3988,N_3131);
and U4576 (N_4576,N_3648,N_3464);
and U4577 (N_4577,N_3299,N_3235);
or U4578 (N_4578,N_3498,N_3419);
xnor U4579 (N_4579,N_3235,N_3222);
nor U4580 (N_4580,N_3141,N_3004);
and U4581 (N_4581,N_3021,N_3248);
nor U4582 (N_4582,N_3878,N_3685);
or U4583 (N_4583,N_3713,N_3766);
nor U4584 (N_4584,N_3826,N_3031);
or U4585 (N_4585,N_3304,N_3161);
and U4586 (N_4586,N_3657,N_3310);
or U4587 (N_4587,N_3140,N_3504);
nand U4588 (N_4588,N_3030,N_3532);
nor U4589 (N_4589,N_3542,N_3350);
or U4590 (N_4590,N_3816,N_3449);
and U4591 (N_4591,N_3342,N_3017);
nor U4592 (N_4592,N_3284,N_3753);
and U4593 (N_4593,N_3316,N_3222);
nor U4594 (N_4594,N_3078,N_3837);
nor U4595 (N_4595,N_3282,N_3850);
nor U4596 (N_4596,N_3425,N_3267);
nand U4597 (N_4597,N_3281,N_3476);
or U4598 (N_4598,N_3553,N_3614);
nand U4599 (N_4599,N_3264,N_3445);
or U4600 (N_4600,N_3139,N_3017);
nand U4601 (N_4601,N_3848,N_3487);
or U4602 (N_4602,N_3575,N_3547);
and U4603 (N_4603,N_3293,N_3279);
or U4604 (N_4604,N_3851,N_3434);
and U4605 (N_4605,N_3732,N_3194);
or U4606 (N_4606,N_3322,N_3463);
nand U4607 (N_4607,N_3024,N_3224);
nor U4608 (N_4608,N_3709,N_3682);
or U4609 (N_4609,N_3856,N_3688);
nand U4610 (N_4610,N_3365,N_3648);
nand U4611 (N_4611,N_3643,N_3469);
nand U4612 (N_4612,N_3821,N_3721);
nor U4613 (N_4613,N_3685,N_3141);
or U4614 (N_4614,N_3705,N_3134);
nand U4615 (N_4615,N_3289,N_3028);
nand U4616 (N_4616,N_3399,N_3305);
nand U4617 (N_4617,N_3760,N_3018);
nor U4618 (N_4618,N_3550,N_3501);
or U4619 (N_4619,N_3442,N_3499);
nand U4620 (N_4620,N_3963,N_3431);
and U4621 (N_4621,N_3852,N_3347);
or U4622 (N_4622,N_3249,N_3316);
nand U4623 (N_4623,N_3333,N_3531);
nor U4624 (N_4624,N_3252,N_3649);
and U4625 (N_4625,N_3053,N_3153);
nor U4626 (N_4626,N_3812,N_3846);
and U4627 (N_4627,N_3233,N_3909);
and U4628 (N_4628,N_3826,N_3238);
nand U4629 (N_4629,N_3098,N_3198);
and U4630 (N_4630,N_3001,N_3817);
and U4631 (N_4631,N_3109,N_3449);
nor U4632 (N_4632,N_3681,N_3975);
and U4633 (N_4633,N_3186,N_3266);
and U4634 (N_4634,N_3681,N_3817);
nand U4635 (N_4635,N_3652,N_3385);
and U4636 (N_4636,N_3670,N_3949);
and U4637 (N_4637,N_3094,N_3597);
nor U4638 (N_4638,N_3866,N_3879);
nor U4639 (N_4639,N_3292,N_3489);
or U4640 (N_4640,N_3908,N_3712);
and U4641 (N_4641,N_3810,N_3361);
nor U4642 (N_4642,N_3761,N_3675);
nand U4643 (N_4643,N_3086,N_3754);
or U4644 (N_4644,N_3565,N_3401);
nand U4645 (N_4645,N_3846,N_3104);
nand U4646 (N_4646,N_3840,N_3506);
or U4647 (N_4647,N_3401,N_3940);
nand U4648 (N_4648,N_3979,N_3074);
or U4649 (N_4649,N_3593,N_3873);
or U4650 (N_4650,N_3378,N_3395);
nand U4651 (N_4651,N_3226,N_3153);
nand U4652 (N_4652,N_3687,N_3804);
xor U4653 (N_4653,N_3558,N_3758);
or U4654 (N_4654,N_3797,N_3937);
nand U4655 (N_4655,N_3357,N_3076);
nand U4656 (N_4656,N_3556,N_3454);
nor U4657 (N_4657,N_3703,N_3680);
nand U4658 (N_4658,N_3300,N_3787);
and U4659 (N_4659,N_3287,N_3203);
or U4660 (N_4660,N_3664,N_3987);
or U4661 (N_4661,N_3187,N_3495);
nor U4662 (N_4662,N_3519,N_3862);
nor U4663 (N_4663,N_3478,N_3785);
or U4664 (N_4664,N_3529,N_3895);
nand U4665 (N_4665,N_3352,N_3582);
and U4666 (N_4666,N_3511,N_3153);
or U4667 (N_4667,N_3601,N_3098);
nand U4668 (N_4668,N_3986,N_3491);
nor U4669 (N_4669,N_3594,N_3830);
or U4670 (N_4670,N_3926,N_3592);
nand U4671 (N_4671,N_3537,N_3709);
or U4672 (N_4672,N_3573,N_3513);
nor U4673 (N_4673,N_3245,N_3987);
nor U4674 (N_4674,N_3138,N_3322);
or U4675 (N_4675,N_3764,N_3556);
nand U4676 (N_4676,N_3130,N_3212);
and U4677 (N_4677,N_3539,N_3623);
nand U4678 (N_4678,N_3071,N_3066);
and U4679 (N_4679,N_3318,N_3204);
and U4680 (N_4680,N_3046,N_3833);
nand U4681 (N_4681,N_3377,N_3780);
or U4682 (N_4682,N_3172,N_3140);
and U4683 (N_4683,N_3341,N_3281);
and U4684 (N_4684,N_3651,N_3512);
or U4685 (N_4685,N_3013,N_3032);
nor U4686 (N_4686,N_3660,N_3734);
and U4687 (N_4687,N_3714,N_3838);
and U4688 (N_4688,N_3257,N_3069);
nand U4689 (N_4689,N_3622,N_3758);
nor U4690 (N_4690,N_3898,N_3646);
nor U4691 (N_4691,N_3401,N_3798);
nand U4692 (N_4692,N_3466,N_3707);
nor U4693 (N_4693,N_3018,N_3636);
nand U4694 (N_4694,N_3794,N_3142);
and U4695 (N_4695,N_3155,N_3593);
nor U4696 (N_4696,N_3705,N_3846);
nand U4697 (N_4697,N_3813,N_3211);
nor U4698 (N_4698,N_3547,N_3503);
xor U4699 (N_4699,N_3267,N_3758);
and U4700 (N_4700,N_3198,N_3310);
nor U4701 (N_4701,N_3951,N_3428);
nand U4702 (N_4702,N_3040,N_3926);
and U4703 (N_4703,N_3757,N_3566);
nand U4704 (N_4704,N_3551,N_3956);
or U4705 (N_4705,N_3699,N_3788);
or U4706 (N_4706,N_3666,N_3862);
nand U4707 (N_4707,N_3965,N_3609);
nand U4708 (N_4708,N_3950,N_3557);
nand U4709 (N_4709,N_3177,N_3115);
and U4710 (N_4710,N_3156,N_3547);
nor U4711 (N_4711,N_3191,N_3144);
and U4712 (N_4712,N_3078,N_3570);
or U4713 (N_4713,N_3562,N_3077);
and U4714 (N_4714,N_3935,N_3542);
or U4715 (N_4715,N_3344,N_3856);
xor U4716 (N_4716,N_3004,N_3417);
nor U4717 (N_4717,N_3829,N_3620);
or U4718 (N_4718,N_3220,N_3903);
or U4719 (N_4719,N_3754,N_3955);
or U4720 (N_4720,N_3529,N_3697);
nand U4721 (N_4721,N_3140,N_3170);
and U4722 (N_4722,N_3075,N_3709);
nand U4723 (N_4723,N_3855,N_3959);
and U4724 (N_4724,N_3668,N_3936);
nand U4725 (N_4725,N_3963,N_3353);
nand U4726 (N_4726,N_3021,N_3318);
or U4727 (N_4727,N_3559,N_3890);
nor U4728 (N_4728,N_3878,N_3246);
and U4729 (N_4729,N_3227,N_3009);
nor U4730 (N_4730,N_3159,N_3700);
and U4731 (N_4731,N_3008,N_3707);
nor U4732 (N_4732,N_3479,N_3981);
and U4733 (N_4733,N_3850,N_3748);
nor U4734 (N_4734,N_3024,N_3929);
nand U4735 (N_4735,N_3618,N_3305);
or U4736 (N_4736,N_3687,N_3244);
nor U4737 (N_4737,N_3798,N_3192);
nand U4738 (N_4738,N_3651,N_3425);
nand U4739 (N_4739,N_3180,N_3127);
and U4740 (N_4740,N_3399,N_3323);
and U4741 (N_4741,N_3224,N_3057);
and U4742 (N_4742,N_3643,N_3115);
nand U4743 (N_4743,N_3163,N_3187);
nand U4744 (N_4744,N_3369,N_3174);
nor U4745 (N_4745,N_3826,N_3866);
nand U4746 (N_4746,N_3757,N_3081);
or U4747 (N_4747,N_3698,N_3433);
xor U4748 (N_4748,N_3959,N_3910);
or U4749 (N_4749,N_3137,N_3744);
and U4750 (N_4750,N_3496,N_3113);
nor U4751 (N_4751,N_3992,N_3556);
nand U4752 (N_4752,N_3086,N_3704);
nor U4753 (N_4753,N_3369,N_3427);
nand U4754 (N_4754,N_3959,N_3478);
or U4755 (N_4755,N_3218,N_3396);
nor U4756 (N_4756,N_3798,N_3732);
or U4757 (N_4757,N_3573,N_3238);
nor U4758 (N_4758,N_3930,N_3436);
or U4759 (N_4759,N_3741,N_3366);
or U4760 (N_4760,N_3892,N_3234);
or U4761 (N_4761,N_3009,N_3341);
nor U4762 (N_4762,N_3419,N_3116);
nor U4763 (N_4763,N_3738,N_3819);
or U4764 (N_4764,N_3390,N_3595);
nand U4765 (N_4765,N_3987,N_3900);
and U4766 (N_4766,N_3496,N_3296);
xnor U4767 (N_4767,N_3268,N_3895);
nand U4768 (N_4768,N_3168,N_3954);
nor U4769 (N_4769,N_3596,N_3755);
nor U4770 (N_4770,N_3382,N_3238);
nand U4771 (N_4771,N_3518,N_3358);
nor U4772 (N_4772,N_3035,N_3402);
nor U4773 (N_4773,N_3427,N_3694);
and U4774 (N_4774,N_3927,N_3417);
and U4775 (N_4775,N_3281,N_3404);
and U4776 (N_4776,N_3475,N_3302);
or U4777 (N_4777,N_3093,N_3230);
and U4778 (N_4778,N_3560,N_3872);
nand U4779 (N_4779,N_3127,N_3384);
or U4780 (N_4780,N_3510,N_3781);
nor U4781 (N_4781,N_3881,N_3311);
and U4782 (N_4782,N_3892,N_3511);
nor U4783 (N_4783,N_3568,N_3190);
nor U4784 (N_4784,N_3144,N_3744);
and U4785 (N_4785,N_3775,N_3665);
and U4786 (N_4786,N_3846,N_3446);
or U4787 (N_4787,N_3238,N_3568);
nand U4788 (N_4788,N_3232,N_3001);
nand U4789 (N_4789,N_3703,N_3427);
nand U4790 (N_4790,N_3420,N_3053);
nor U4791 (N_4791,N_3342,N_3260);
or U4792 (N_4792,N_3274,N_3745);
and U4793 (N_4793,N_3302,N_3441);
nor U4794 (N_4794,N_3866,N_3150);
or U4795 (N_4795,N_3362,N_3909);
or U4796 (N_4796,N_3654,N_3548);
nand U4797 (N_4797,N_3418,N_3889);
or U4798 (N_4798,N_3540,N_3609);
and U4799 (N_4799,N_3409,N_3161);
nor U4800 (N_4800,N_3949,N_3548);
and U4801 (N_4801,N_3663,N_3057);
nand U4802 (N_4802,N_3693,N_3836);
or U4803 (N_4803,N_3829,N_3741);
and U4804 (N_4804,N_3047,N_3560);
nor U4805 (N_4805,N_3688,N_3480);
and U4806 (N_4806,N_3549,N_3135);
nor U4807 (N_4807,N_3695,N_3427);
and U4808 (N_4808,N_3362,N_3732);
nand U4809 (N_4809,N_3036,N_3836);
or U4810 (N_4810,N_3290,N_3672);
nor U4811 (N_4811,N_3194,N_3585);
or U4812 (N_4812,N_3302,N_3914);
or U4813 (N_4813,N_3610,N_3970);
and U4814 (N_4814,N_3228,N_3509);
or U4815 (N_4815,N_3927,N_3438);
and U4816 (N_4816,N_3971,N_3983);
nand U4817 (N_4817,N_3882,N_3456);
nand U4818 (N_4818,N_3134,N_3004);
nand U4819 (N_4819,N_3124,N_3327);
or U4820 (N_4820,N_3469,N_3924);
nor U4821 (N_4821,N_3250,N_3679);
nand U4822 (N_4822,N_3176,N_3880);
nor U4823 (N_4823,N_3467,N_3665);
and U4824 (N_4824,N_3071,N_3151);
or U4825 (N_4825,N_3794,N_3871);
and U4826 (N_4826,N_3681,N_3097);
nor U4827 (N_4827,N_3995,N_3422);
nand U4828 (N_4828,N_3912,N_3988);
nand U4829 (N_4829,N_3481,N_3458);
nand U4830 (N_4830,N_3604,N_3938);
or U4831 (N_4831,N_3200,N_3260);
or U4832 (N_4832,N_3727,N_3277);
or U4833 (N_4833,N_3894,N_3037);
nand U4834 (N_4834,N_3427,N_3101);
or U4835 (N_4835,N_3945,N_3298);
nor U4836 (N_4836,N_3948,N_3877);
nor U4837 (N_4837,N_3059,N_3315);
and U4838 (N_4838,N_3809,N_3049);
nor U4839 (N_4839,N_3186,N_3401);
nor U4840 (N_4840,N_3999,N_3804);
xor U4841 (N_4841,N_3697,N_3428);
and U4842 (N_4842,N_3693,N_3913);
nor U4843 (N_4843,N_3706,N_3444);
nand U4844 (N_4844,N_3956,N_3563);
and U4845 (N_4845,N_3099,N_3559);
nand U4846 (N_4846,N_3084,N_3953);
nor U4847 (N_4847,N_3246,N_3308);
nor U4848 (N_4848,N_3778,N_3569);
nand U4849 (N_4849,N_3380,N_3831);
or U4850 (N_4850,N_3010,N_3261);
nand U4851 (N_4851,N_3866,N_3938);
nor U4852 (N_4852,N_3355,N_3507);
or U4853 (N_4853,N_3543,N_3057);
nor U4854 (N_4854,N_3615,N_3199);
nor U4855 (N_4855,N_3883,N_3536);
nor U4856 (N_4856,N_3582,N_3089);
nand U4857 (N_4857,N_3018,N_3468);
or U4858 (N_4858,N_3976,N_3993);
nand U4859 (N_4859,N_3498,N_3667);
nor U4860 (N_4860,N_3785,N_3488);
or U4861 (N_4861,N_3311,N_3330);
nor U4862 (N_4862,N_3070,N_3118);
or U4863 (N_4863,N_3966,N_3170);
and U4864 (N_4864,N_3546,N_3500);
or U4865 (N_4865,N_3990,N_3423);
nand U4866 (N_4866,N_3740,N_3265);
nor U4867 (N_4867,N_3370,N_3137);
nor U4868 (N_4868,N_3071,N_3486);
nand U4869 (N_4869,N_3420,N_3242);
nand U4870 (N_4870,N_3571,N_3891);
xnor U4871 (N_4871,N_3187,N_3830);
or U4872 (N_4872,N_3608,N_3618);
or U4873 (N_4873,N_3424,N_3624);
xor U4874 (N_4874,N_3758,N_3935);
nor U4875 (N_4875,N_3216,N_3639);
or U4876 (N_4876,N_3723,N_3630);
nor U4877 (N_4877,N_3865,N_3260);
and U4878 (N_4878,N_3778,N_3587);
nand U4879 (N_4879,N_3969,N_3479);
xor U4880 (N_4880,N_3534,N_3288);
nand U4881 (N_4881,N_3109,N_3559);
and U4882 (N_4882,N_3582,N_3834);
nand U4883 (N_4883,N_3425,N_3199);
nor U4884 (N_4884,N_3090,N_3936);
xor U4885 (N_4885,N_3140,N_3175);
nor U4886 (N_4886,N_3036,N_3934);
nand U4887 (N_4887,N_3575,N_3503);
and U4888 (N_4888,N_3430,N_3861);
nand U4889 (N_4889,N_3128,N_3719);
and U4890 (N_4890,N_3153,N_3004);
and U4891 (N_4891,N_3630,N_3632);
and U4892 (N_4892,N_3110,N_3915);
nor U4893 (N_4893,N_3087,N_3929);
and U4894 (N_4894,N_3379,N_3083);
or U4895 (N_4895,N_3101,N_3664);
nor U4896 (N_4896,N_3756,N_3611);
and U4897 (N_4897,N_3150,N_3798);
nand U4898 (N_4898,N_3953,N_3649);
xor U4899 (N_4899,N_3871,N_3717);
and U4900 (N_4900,N_3970,N_3062);
nor U4901 (N_4901,N_3831,N_3927);
nand U4902 (N_4902,N_3868,N_3047);
or U4903 (N_4903,N_3227,N_3091);
and U4904 (N_4904,N_3909,N_3341);
nand U4905 (N_4905,N_3092,N_3749);
nand U4906 (N_4906,N_3877,N_3814);
xor U4907 (N_4907,N_3656,N_3338);
and U4908 (N_4908,N_3849,N_3180);
and U4909 (N_4909,N_3165,N_3623);
and U4910 (N_4910,N_3097,N_3053);
and U4911 (N_4911,N_3739,N_3224);
or U4912 (N_4912,N_3476,N_3161);
and U4913 (N_4913,N_3307,N_3065);
nor U4914 (N_4914,N_3852,N_3741);
nor U4915 (N_4915,N_3111,N_3792);
and U4916 (N_4916,N_3204,N_3508);
nor U4917 (N_4917,N_3892,N_3133);
nand U4918 (N_4918,N_3889,N_3460);
and U4919 (N_4919,N_3521,N_3745);
nor U4920 (N_4920,N_3223,N_3262);
nand U4921 (N_4921,N_3575,N_3339);
nand U4922 (N_4922,N_3570,N_3733);
and U4923 (N_4923,N_3722,N_3998);
and U4924 (N_4924,N_3277,N_3245);
nor U4925 (N_4925,N_3848,N_3276);
nor U4926 (N_4926,N_3532,N_3617);
nor U4927 (N_4927,N_3654,N_3710);
nand U4928 (N_4928,N_3838,N_3456);
or U4929 (N_4929,N_3610,N_3268);
nand U4930 (N_4930,N_3825,N_3980);
or U4931 (N_4931,N_3443,N_3306);
and U4932 (N_4932,N_3967,N_3643);
and U4933 (N_4933,N_3305,N_3599);
nand U4934 (N_4934,N_3938,N_3336);
and U4935 (N_4935,N_3395,N_3159);
nand U4936 (N_4936,N_3258,N_3381);
or U4937 (N_4937,N_3295,N_3689);
nand U4938 (N_4938,N_3844,N_3053);
and U4939 (N_4939,N_3345,N_3789);
or U4940 (N_4940,N_3620,N_3665);
or U4941 (N_4941,N_3011,N_3187);
and U4942 (N_4942,N_3197,N_3164);
xnor U4943 (N_4943,N_3085,N_3539);
and U4944 (N_4944,N_3434,N_3627);
and U4945 (N_4945,N_3612,N_3892);
xnor U4946 (N_4946,N_3071,N_3502);
or U4947 (N_4947,N_3366,N_3890);
and U4948 (N_4948,N_3147,N_3288);
and U4949 (N_4949,N_3257,N_3344);
nor U4950 (N_4950,N_3828,N_3256);
and U4951 (N_4951,N_3574,N_3114);
nand U4952 (N_4952,N_3015,N_3722);
nand U4953 (N_4953,N_3720,N_3810);
nor U4954 (N_4954,N_3974,N_3547);
nor U4955 (N_4955,N_3129,N_3690);
nand U4956 (N_4956,N_3942,N_3286);
or U4957 (N_4957,N_3219,N_3706);
or U4958 (N_4958,N_3234,N_3695);
and U4959 (N_4959,N_3436,N_3069);
or U4960 (N_4960,N_3843,N_3161);
nor U4961 (N_4961,N_3265,N_3359);
nand U4962 (N_4962,N_3235,N_3297);
nor U4963 (N_4963,N_3555,N_3664);
nor U4964 (N_4964,N_3151,N_3959);
or U4965 (N_4965,N_3936,N_3124);
and U4966 (N_4966,N_3915,N_3315);
nand U4967 (N_4967,N_3705,N_3137);
nand U4968 (N_4968,N_3874,N_3121);
nor U4969 (N_4969,N_3191,N_3044);
nor U4970 (N_4970,N_3988,N_3549);
nand U4971 (N_4971,N_3877,N_3443);
nand U4972 (N_4972,N_3093,N_3429);
or U4973 (N_4973,N_3961,N_3438);
and U4974 (N_4974,N_3399,N_3286);
and U4975 (N_4975,N_3754,N_3108);
and U4976 (N_4976,N_3815,N_3597);
and U4977 (N_4977,N_3360,N_3991);
nor U4978 (N_4978,N_3880,N_3140);
or U4979 (N_4979,N_3018,N_3940);
or U4980 (N_4980,N_3615,N_3455);
and U4981 (N_4981,N_3895,N_3994);
and U4982 (N_4982,N_3002,N_3192);
nor U4983 (N_4983,N_3558,N_3031);
and U4984 (N_4984,N_3731,N_3164);
or U4985 (N_4985,N_3485,N_3532);
nor U4986 (N_4986,N_3688,N_3971);
xor U4987 (N_4987,N_3663,N_3078);
nand U4988 (N_4988,N_3012,N_3451);
and U4989 (N_4989,N_3285,N_3926);
nor U4990 (N_4990,N_3117,N_3162);
nor U4991 (N_4991,N_3985,N_3577);
nand U4992 (N_4992,N_3360,N_3169);
and U4993 (N_4993,N_3035,N_3729);
nand U4994 (N_4994,N_3737,N_3262);
nor U4995 (N_4995,N_3831,N_3991);
or U4996 (N_4996,N_3466,N_3309);
xnor U4997 (N_4997,N_3025,N_3136);
nor U4998 (N_4998,N_3235,N_3123);
or U4999 (N_4999,N_3499,N_3076);
or UO_0 (O_0,N_4368,N_4477);
or UO_1 (O_1,N_4841,N_4800);
and UO_2 (O_2,N_4309,N_4732);
nor UO_3 (O_3,N_4527,N_4925);
nand UO_4 (O_4,N_4748,N_4337);
or UO_5 (O_5,N_4495,N_4150);
and UO_6 (O_6,N_4422,N_4213);
or UO_7 (O_7,N_4632,N_4525);
nor UO_8 (O_8,N_4733,N_4012);
and UO_9 (O_9,N_4242,N_4194);
nand UO_10 (O_10,N_4342,N_4420);
or UO_11 (O_11,N_4146,N_4860);
nand UO_12 (O_12,N_4695,N_4131);
or UO_13 (O_13,N_4757,N_4161);
and UO_14 (O_14,N_4284,N_4238);
nor UO_15 (O_15,N_4974,N_4159);
nor UO_16 (O_16,N_4214,N_4389);
and UO_17 (O_17,N_4931,N_4363);
and UO_18 (O_18,N_4351,N_4911);
or UO_19 (O_19,N_4057,N_4714);
and UO_20 (O_20,N_4723,N_4809);
nor UO_21 (O_21,N_4643,N_4324);
nand UO_22 (O_22,N_4487,N_4502);
and UO_23 (O_23,N_4443,N_4429);
nand UO_24 (O_24,N_4290,N_4038);
nor UO_25 (O_25,N_4188,N_4927);
nand UO_26 (O_26,N_4271,N_4036);
nor UO_27 (O_27,N_4541,N_4153);
nor UO_28 (O_28,N_4582,N_4893);
or UO_29 (O_29,N_4503,N_4580);
or UO_30 (O_30,N_4303,N_4829);
or UO_31 (O_31,N_4781,N_4787);
or UO_32 (O_32,N_4965,N_4382);
and UO_33 (O_33,N_4500,N_4837);
or UO_34 (O_34,N_4745,N_4967);
or UO_35 (O_35,N_4231,N_4239);
and UO_36 (O_36,N_4418,N_4071);
and UO_37 (O_37,N_4707,N_4544);
nand UO_38 (O_38,N_4205,N_4882);
nand UO_39 (O_39,N_4996,N_4097);
and UO_40 (O_40,N_4570,N_4111);
nand UO_41 (O_41,N_4497,N_4456);
or UO_42 (O_42,N_4144,N_4210);
nor UO_43 (O_43,N_4653,N_4622);
and UO_44 (O_44,N_4921,N_4450);
nor UO_45 (O_45,N_4407,N_4658);
and UO_46 (O_46,N_4591,N_4050);
and UO_47 (O_47,N_4721,N_4319);
nor UO_48 (O_48,N_4042,N_4133);
and UO_49 (O_49,N_4986,N_4275);
or UO_50 (O_50,N_4228,N_4143);
nand UO_51 (O_51,N_4181,N_4127);
nand UO_52 (O_52,N_4372,N_4762);
nand UO_53 (O_53,N_4227,N_4908);
nor UO_54 (O_54,N_4964,N_4857);
or UO_55 (O_55,N_4813,N_4003);
nor UO_56 (O_56,N_4509,N_4252);
or UO_57 (O_57,N_4192,N_4076);
nand UO_58 (O_58,N_4014,N_4444);
and UO_59 (O_59,N_4453,N_4427);
and UO_60 (O_60,N_4025,N_4620);
or UO_61 (O_61,N_4824,N_4321);
or UO_62 (O_62,N_4631,N_4177);
nor UO_63 (O_63,N_4668,N_4564);
or UO_64 (O_64,N_4114,N_4508);
and UO_65 (O_65,N_4362,N_4627);
and UO_66 (O_66,N_4322,N_4777);
or UO_67 (O_67,N_4918,N_4356);
nand UO_68 (O_68,N_4152,N_4796);
nor UO_69 (O_69,N_4330,N_4089);
and UO_70 (O_70,N_4718,N_4528);
nor UO_71 (O_71,N_4128,N_4229);
and UO_72 (O_72,N_4391,N_4613);
nor UO_73 (O_73,N_4867,N_4053);
or UO_74 (O_74,N_4215,N_4990);
and UO_75 (O_75,N_4838,N_4577);
nand UO_76 (O_76,N_4682,N_4460);
nor UO_77 (O_77,N_4393,N_4346);
nor UO_78 (O_78,N_4780,N_4191);
and UO_79 (O_79,N_4415,N_4123);
or UO_80 (O_80,N_4889,N_4056);
nor UO_81 (O_81,N_4307,N_4994);
or UO_82 (O_82,N_4295,N_4088);
or UO_83 (O_83,N_4696,N_4514);
nor UO_84 (O_84,N_4575,N_4232);
or UO_85 (O_85,N_4440,N_4872);
and UO_86 (O_86,N_4080,N_4786);
xor UO_87 (O_87,N_4226,N_4736);
nand UO_88 (O_88,N_4834,N_4431);
nor UO_89 (O_89,N_4300,N_4886);
and UO_90 (O_90,N_4955,N_4505);
and UO_91 (O_91,N_4022,N_4568);
or UO_92 (O_92,N_4712,N_4166);
nand UO_93 (O_93,N_4864,N_4155);
nor UO_94 (O_94,N_4173,N_4944);
or UO_95 (O_95,N_4428,N_4753);
nor UO_96 (O_96,N_4851,N_4469);
or UO_97 (O_97,N_4017,N_4016);
or UO_98 (O_98,N_4065,N_4545);
nand UO_99 (O_99,N_4654,N_4963);
nor UO_100 (O_100,N_4353,N_4028);
or UO_101 (O_101,N_4280,N_4744);
nand UO_102 (O_102,N_4381,N_4576);
nand UO_103 (O_103,N_4984,N_4385);
nor UO_104 (O_104,N_4616,N_4833);
or UO_105 (O_105,N_4988,N_4052);
xnor UO_106 (O_106,N_4865,N_4105);
or UO_107 (O_107,N_4218,N_4660);
nor UO_108 (O_108,N_4416,N_4141);
nor UO_109 (O_109,N_4818,N_4675);
and UO_110 (O_110,N_4002,N_4273);
nand UO_111 (O_111,N_4184,N_4709);
nand UO_112 (O_112,N_4629,N_4225);
and UO_113 (O_113,N_4788,N_4451);
and UO_114 (O_114,N_4399,N_4198);
nor UO_115 (O_115,N_4673,N_4083);
nand UO_116 (O_116,N_4187,N_4852);
or UO_117 (O_117,N_4145,N_4426);
nor UO_118 (O_118,N_4434,N_4529);
nand UO_119 (O_119,N_4490,N_4815);
or UO_120 (O_120,N_4458,N_4532);
and UO_121 (O_121,N_4684,N_4806);
nor UO_122 (O_122,N_4007,N_4727);
nand UO_123 (O_123,N_4211,N_4171);
nand UO_124 (O_124,N_4909,N_4315);
or UO_125 (O_125,N_4236,N_4033);
nand UO_126 (O_126,N_4015,N_4785);
nor UO_127 (O_127,N_4004,N_4738);
xor UO_128 (O_128,N_4726,N_4929);
and UO_129 (O_129,N_4890,N_4926);
nand UO_130 (O_130,N_4085,N_4983);
nor UO_131 (O_131,N_4339,N_4384);
nand UO_132 (O_132,N_4976,N_4896);
nand UO_133 (O_133,N_4596,N_4095);
nor UO_134 (O_134,N_4072,N_4068);
nand UO_135 (O_135,N_4092,N_4581);
or UO_136 (O_136,N_4357,N_4661);
or UO_137 (O_137,N_4801,N_4438);
and UO_138 (O_138,N_4794,N_4621);
and UO_139 (O_139,N_4817,N_4607);
nand UO_140 (O_140,N_4104,N_4109);
nor UO_141 (O_141,N_4987,N_4183);
and UO_142 (O_142,N_4482,N_4037);
nand UO_143 (O_143,N_4196,N_4135);
and UO_144 (O_144,N_4485,N_4790);
or UO_145 (O_145,N_4405,N_4822);
or UO_146 (O_146,N_4708,N_4553);
or UO_147 (O_147,N_4245,N_4219);
or UO_148 (O_148,N_4916,N_4945);
nor UO_149 (O_149,N_4840,N_4592);
and UO_150 (O_150,N_4255,N_4612);
and UO_151 (O_151,N_4871,N_4234);
nor UO_152 (O_152,N_4008,N_4101);
and UO_153 (O_153,N_4628,N_4463);
nor UO_154 (O_154,N_4314,N_4262);
and UO_155 (O_155,N_4870,N_4151);
or UO_156 (O_156,N_4040,N_4774);
nor UO_157 (O_157,N_4048,N_4947);
and UO_158 (O_158,N_4470,N_4206);
or UO_159 (O_159,N_4973,N_4064);
and UO_160 (O_160,N_4681,N_4350);
or UO_161 (O_161,N_4378,N_4797);
or UO_162 (O_162,N_4062,N_4137);
nor UO_163 (O_163,N_4881,N_4977);
nand UO_164 (O_164,N_4783,N_4634);
or UO_165 (O_165,N_4536,N_4140);
nand UO_166 (O_166,N_4334,N_4594);
or UO_167 (O_167,N_4432,N_4139);
nor UO_168 (O_168,N_4934,N_4803);
or UO_169 (O_169,N_4812,N_4699);
nand UO_170 (O_170,N_4784,N_4473);
nand UO_171 (O_171,N_4656,N_4878);
or UO_172 (O_172,N_4782,N_4396);
and UO_173 (O_173,N_4539,N_4449);
or UO_174 (O_174,N_4240,N_4808);
nor UO_175 (O_175,N_4625,N_4876);
nor UO_176 (O_176,N_4154,N_4020);
nor UO_177 (O_177,N_4247,N_4730);
nor UO_178 (O_178,N_4531,N_4676);
or UO_179 (O_179,N_4633,N_4630);
and UO_180 (O_180,N_4483,N_4717);
or UO_181 (O_181,N_4390,N_4107);
or UO_182 (O_182,N_4667,N_4941);
and UO_183 (O_183,N_4367,N_4799);
nand UO_184 (O_184,N_4488,N_4202);
nand UO_185 (O_185,N_4162,N_4725);
nor UO_186 (O_186,N_4999,N_4193);
and UO_187 (O_187,N_4603,N_4826);
or UO_188 (O_188,N_4602,N_4519);
nor UO_189 (O_189,N_4601,N_4742);
nor UO_190 (O_190,N_4058,N_4816);
or UO_191 (O_191,N_4773,N_4641);
nor UO_192 (O_192,N_4026,N_4827);
nand UO_193 (O_193,N_4567,N_4116);
nand UO_194 (O_194,N_4398,N_4222);
and UO_195 (O_195,N_4679,N_4253);
nor UO_196 (O_196,N_4254,N_4626);
nor UO_197 (O_197,N_4044,N_4383);
nand UO_198 (O_198,N_4597,N_4566);
nor UO_199 (O_199,N_4365,N_4775);
and UO_200 (O_200,N_4935,N_4433);
or UO_201 (O_201,N_4515,N_4689);
nor UO_202 (O_202,N_4542,N_4165);
nor UO_203 (O_203,N_4891,N_4523);
nand UO_204 (O_204,N_4377,N_4494);
nand UO_205 (O_205,N_4939,N_4261);
nor UO_206 (O_206,N_4855,N_4070);
nand UO_207 (O_207,N_4618,N_4244);
nor UO_208 (O_208,N_4397,N_4583);
nor UO_209 (O_209,N_4129,N_4493);
nor UO_210 (O_210,N_4138,N_4340);
nand UO_211 (O_211,N_4358,N_4705);
nor UO_212 (O_212,N_4847,N_4359);
and UO_213 (O_213,N_4454,N_4952);
or UO_214 (O_214,N_4169,N_4595);
or UO_215 (O_215,N_4966,N_4659);
nand UO_216 (O_216,N_4992,N_4543);
nand UO_217 (O_217,N_4124,N_4185);
or UO_218 (O_218,N_4106,N_4474);
nand UO_219 (O_219,N_4610,N_4501);
xor UO_220 (O_220,N_4031,N_4301);
nor UO_221 (O_221,N_4928,N_4480);
and UO_222 (O_222,N_4655,N_4018);
nand UO_223 (O_223,N_4924,N_4086);
or UO_224 (O_224,N_4619,N_4197);
nand UO_225 (O_225,N_4555,N_4703);
nor UO_226 (O_226,N_4327,N_4765);
nand UO_227 (O_227,N_4289,N_4439);
and UO_228 (O_228,N_4204,N_4175);
and UO_229 (O_229,N_4035,N_4572);
xnor UO_230 (O_230,N_4376,N_4323);
and UO_231 (O_231,N_4027,N_4291);
and UO_232 (O_232,N_4554,N_4671);
nor UO_233 (O_233,N_4073,N_4912);
nor UO_234 (O_234,N_4856,N_4233);
nor UO_235 (O_235,N_4112,N_4954);
and UO_236 (O_236,N_4691,N_4969);
or UO_237 (O_237,N_4286,N_4549);
or UO_238 (O_238,N_4122,N_4863);
xor UO_239 (O_239,N_4574,N_4805);
and UO_240 (O_240,N_4795,N_4306);
nor UO_241 (O_241,N_4164,N_4190);
xnor UO_242 (O_242,N_4614,N_4930);
nor UO_243 (O_243,N_4267,N_4825);
and UO_244 (O_244,N_4571,N_4513);
or UO_245 (O_245,N_4221,N_4972);
and UO_246 (O_246,N_4836,N_4103);
or UO_247 (O_247,N_4237,N_4318);
nor UO_248 (O_248,N_4646,N_4063);
nor UO_249 (O_249,N_4979,N_4666);
or UO_250 (O_250,N_4913,N_4821);
and UO_251 (O_251,N_4904,N_4650);
or UO_252 (O_252,N_4546,N_4264);
nor UO_253 (O_253,N_4403,N_4932);
nand UO_254 (O_254,N_4537,N_4149);
nand UO_255 (O_255,N_4352,N_4120);
nor UO_256 (O_256,N_4710,N_4600);
or UO_257 (O_257,N_4258,N_4586);
or UO_258 (O_258,N_4338,N_4409);
nor UO_259 (O_259,N_4388,N_4716);
and UO_260 (O_260,N_4875,N_4640);
nand UO_261 (O_261,N_4452,N_4305);
and UO_262 (O_262,N_4496,N_4345);
nand UO_263 (O_263,N_4968,N_4302);
or UO_264 (O_264,N_4995,N_4764);
and UO_265 (O_265,N_4760,N_4134);
or UO_266 (O_266,N_4142,N_4110);
nor UO_267 (O_267,N_4688,N_4437);
and UO_268 (O_268,N_4425,N_4579);
and UO_269 (O_269,N_4936,N_4364);
nor UO_270 (O_270,N_4749,N_4157);
nand UO_271 (O_271,N_4678,N_4859);
or UO_272 (O_272,N_4078,N_4556);
nand UO_273 (O_273,N_4522,N_4844);
nor UO_274 (O_274,N_4615,N_4804);
or UO_275 (O_275,N_4895,N_4410);
and UO_276 (O_276,N_4598,N_4938);
nor UO_277 (O_277,N_4333,N_4702);
and UO_278 (O_278,N_4414,N_4670);
nand UO_279 (O_279,N_4313,N_4858);
nand UO_280 (O_280,N_4066,N_4960);
or UO_281 (O_281,N_4902,N_4569);
nor UO_282 (O_282,N_4098,N_4959);
xor UO_283 (O_283,N_4693,N_4186);
nor UO_284 (O_284,N_4810,N_4259);
or UO_285 (O_285,N_4997,N_4224);
nand UO_286 (O_286,N_4683,N_4520);
and UO_287 (O_287,N_4332,N_4779);
and UO_288 (O_288,N_4958,N_4680);
and UO_289 (O_289,N_4713,N_4189);
nand UO_290 (O_290,N_4272,N_4094);
or UO_291 (O_291,N_4923,N_4498);
xnor UO_292 (O_292,N_4850,N_4652);
or UO_293 (O_293,N_4329,N_4701);
or UO_294 (O_294,N_4132,N_4386);
and UO_295 (O_295,N_4814,N_4516);
and UO_296 (O_296,N_4970,N_4687);
nand UO_297 (O_297,N_4282,N_4769);
and UO_298 (O_298,N_4663,N_4336);
and UO_299 (O_299,N_4914,N_4811);
or UO_300 (O_300,N_4069,N_4354);
or UO_301 (O_301,N_4669,N_4512);
or UO_302 (O_302,N_4770,N_4866);
nand UO_303 (O_303,N_4030,N_4328);
and UO_304 (O_304,N_4167,N_4465);
or UO_305 (O_305,N_4310,N_4412);
nand UO_306 (O_306,N_4442,N_4754);
nor UO_307 (O_307,N_4756,N_4090);
nor UO_308 (O_308,N_4751,N_4763);
nand UO_309 (O_309,N_4557,N_4013);
or UO_310 (O_310,N_4046,N_4119);
and UO_311 (O_311,N_4989,N_4355);
or UO_312 (O_312,N_4606,N_4125);
or UO_313 (O_313,N_4251,N_4534);
nor UO_314 (O_314,N_4373,N_4919);
and UO_315 (O_315,N_4395,N_4755);
nand UO_316 (O_316,N_4611,N_4371);
nand UO_317 (O_317,N_4906,N_4686);
and UO_318 (O_318,N_4894,N_4343);
nand UO_319 (O_319,N_4957,N_4903);
or UO_320 (O_320,N_4526,N_4010);
nor UO_321 (O_321,N_4468,N_4467);
nand UO_322 (O_322,N_4049,N_4820);
and UO_323 (O_323,N_4647,N_4750);
nor UO_324 (O_324,N_4943,N_4081);
nor UO_325 (O_325,N_4366,N_4294);
or UO_326 (O_326,N_4486,N_4406);
nand UO_327 (O_327,N_4320,N_4915);
nand UO_328 (O_328,N_4005,N_4802);
or UO_329 (O_329,N_4061,N_4517);
nand UO_330 (O_330,N_4423,N_4521);
or UO_331 (O_331,N_4248,N_4293);
and UO_332 (O_332,N_4304,N_4156);
nor UO_333 (O_333,N_4243,N_4113);
nand UO_334 (O_334,N_4369,N_4475);
nor UO_335 (O_335,N_4277,N_4341);
or UO_336 (O_336,N_4148,N_4953);
nand UO_337 (O_337,N_4436,N_4511);
nor UO_338 (O_338,N_4873,N_4920);
or UO_339 (O_339,N_4807,N_4067);
nand UO_340 (O_340,N_4160,N_4768);
nor UO_341 (O_341,N_4380,N_4108);
nand UO_342 (O_342,N_4715,N_4182);
nor UO_343 (O_343,N_4249,N_4846);
and UO_344 (O_344,N_4082,N_4547);
and UO_345 (O_345,N_4698,N_4692);
nand UO_346 (O_346,N_4349,N_4880);
and UO_347 (O_347,N_4819,N_4484);
nor UO_348 (O_348,N_4370,N_4000);
and UO_349 (O_349,N_4901,N_4441);
or UO_350 (O_350,N_4766,N_4117);
or UO_351 (O_351,N_4874,N_4019);
or UO_352 (O_352,N_4985,N_4344);
nor UO_353 (O_353,N_4981,N_4637);
and UO_354 (O_354,N_4793,N_4402);
and UO_355 (O_355,N_4897,N_4848);
xor UO_356 (O_356,N_4734,N_4424);
and UO_357 (O_357,N_4608,N_4464);
nor UO_358 (O_358,N_4664,N_4455);
and UO_359 (O_359,N_4032,N_4533);
nor UO_360 (O_360,N_4778,N_4642);
nor UO_361 (O_361,N_4023,N_4998);
and UO_362 (O_362,N_4281,N_4690);
nand UO_363 (O_363,N_4212,N_4518);
nor UO_364 (O_364,N_4636,N_4179);
and UO_365 (O_365,N_4492,N_4297);
nand UO_366 (O_366,N_4203,N_4335);
and UO_367 (O_367,N_4263,N_4223);
nand UO_368 (O_368,N_4674,N_4317);
nand UO_369 (O_369,N_4685,N_4538);
or UO_370 (O_370,N_4843,N_4375);
or UO_371 (O_371,N_4937,N_4201);
and UO_372 (O_372,N_4348,N_4563);
nor UO_373 (O_373,N_4900,N_4216);
and UO_374 (O_374,N_4605,N_4694);
nor UO_375 (O_375,N_4722,N_4946);
nand UO_376 (O_376,N_4311,N_4158);
and UO_377 (O_377,N_4623,N_4269);
or UO_378 (O_378,N_4180,N_4609);
or UO_379 (O_379,N_4411,N_4540);
and UO_380 (O_380,N_4728,N_4457);
and UO_381 (O_381,N_4408,N_4933);
nand UO_382 (O_382,N_4853,N_4325);
nand UO_383 (O_383,N_4835,N_4499);
or UO_384 (O_384,N_4791,N_4948);
nand UO_385 (O_385,N_4059,N_4472);
or UO_386 (O_386,N_4230,N_4208);
and UO_387 (O_387,N_4892,N_4102);
nand UO_388 (O_388,N_4430,N_4172);
nor UO_389 (O_389,N_4093,N_4831);
nor UO_390 (O_390,N_4126,N_4772);
or UO_391 (O_391,N_4740,N_4459);
nand UO_392 (O_392,N_4700,N_4697);
and UO_393 (O_393,N_4100,N_4256);
and UO_394 (O_394,N_4752,N_4077);
nand UO_395 (O_395,N_4624,N_4001);
or UO_396 (O_396,N_4758,N_4392);
nand UO_397 (O_397,N_4055,N_4510);
or UO_398 (O_398,N_4551,N_4462);
or UO_399 (O_399,N_4400,N_4832);
and UO_400 (O_400,N_4299,N_4746);
nor UO_401 (O_401,N_4504,N_4885);
nor UO_402 (O_402,N_4879,N_4278);
nand UO_403 (O_403,N_4877,N_4949);
or UO_404 (O_404,N_4374,N_4711);
and UO_405 (O_405,N_4798,N_4009);
nand UO_406 (O_406,N_4651,N_4163);
nand UO_407 (O_407,N_4195,N_4079);
nand UO_408 (O_408,N_4849,N_4471);
nand UO_409 (O_409,N_4387,N_4199);
nor UO_410 (O_410,N_4250,N_4021);
nor UO_411 (O_411,N_4975,N_4604);
nand UO_412 (O_412,N_4034,N_4417);
and UO_413 (O_413,N_4029,N_4617);
nand UO_414 (O_414,N_4445,N_4771);
and UO_415 (O_415,N_4447,N_4446);
or UO_416 (O_416,N_4584,N_4888);
or UO_417 (O_417,N_4743,N_4266);
or UO_418 (O_418,N_4401,N_4011);
nand UO_419 (O_419,N_4558,N_4361);
and UO_420 (O_420,N_4130,N_4993);
nor UO_421 (O_421,N_4121,N_4479);
and UO_422 (O_422,N_4298,N_4524);
or UO_423 (O_423,N_4147,N_4170);
and UO_424 (O_424,N_4039,N_4276);
nand UO_425 (O_425,N_4489,N_4560);
nand UO_426 (O_426,N_4246,N_4379);
nor UO_427 (O_427,N_4991,N_4060);
and UO_428 (O_428,N_4466,N_4115);
nor UO_429 (O_429,N_4448,N_4260);
nor UO_430 (O_430,N_4074,N_4731);
or UO_431 (O_431,N_4176,N_4257);
and UO_432 (O_432,N_4747,N_4235);
nand UO_433 (O_433,N_4823,N_4862);
or UO_434 (O_434,N_4506,N_4980);
nor UO_435 (O_435,N_4207,N_4599);
nand UO_436 (O_436,N_4719,N_4887);
nand UO_437 (O_437,N_4220,N_4869);
and UO_438 (O_438,N_4905,N_4168);
nand UO_439 (O_439,N_4645,N_4279);
and UO_440 (O_440,N_4308,N_4565);
or UO_441 (O_441,N_4561,N_4724);
or UO_442 (O_442,N_4476,N_4562);
and UO_443 (O_443,N_4638,N_4550);
nor UO_444 (O_444,N_4209,N_4435);
and UO_445 (O_445,N_4741,N_4587);
nand UO_446 (O_446,N_4585,N_4507);
and UO_447 (O_447,N_4917,N_4789);
xnor UO_448 (O_448,N_4830,N_4761);
and UO_449 (O_449,N_4296,N_4404);
and UO_450 (O_450,N_4047,N_4665);
nor UO_451 (O_451,N_4644,N_4978);
nand UO_452 (O_452,N_4739,N_4178);
xor UO_453 (O_453,N_4961,N_4360);
nand UO_454 (O_454,N_4677,N_4720);
xor UO_455 (O_455,N_4593,N_4288);
nand UO_456 (O_456,N_4922,N_4729);
and UO_457 (O_457,N_4589,N_4737);
and UO_458 (O_458,N_4951,N_4043);
and UO_459 (O_459,N_4861,N_4635);
nor UO_460 (O_460,N_4828,N_4971);
and UO_461 (O_461,N_4950,N_4639);
or UO_462 (O_462,N_4842,N_4530);
nor UO_463 (O_463,N_4845,N_4898);
or UO_464 (O_464,N_4421,N_4099);
and UO_465 (O_465,N_4854,N_4578);
and UO_466 (O_466,N_4910,N_4956);
nor UO_467 (O_467,N_4312,N_4942);
nand UO_468 (O_468,N_4759,N_4241);
and UO_469 (O_469,N_4649,N_4274);
nand UO_470 (O_470,N_4962,N_4268);
nor UO_471 (O_471,N_4096,N_4478);
nor UO_472 (O_472,N_4006,N_4648);
nand UO_473 (O_473,N_4839,N_4347);
or UO_474 (O_474,N_4174,N_4657);
or UO_475 (O_475,N_4868,N_4326);
or UO_476 (O_476,N_4899,N_4907);
and UO_477 (O_477,N_4461,N_4045);
nand UO_478 (O_478,N_4491,N_4075);
nor UO_479 (O_479,N_4287,N_4481);
nor UO_480 (O_480,N_4559,N_4940);
nor UO_481 (O_481,N_4552,N_4792);
nor UO_482 (O_482,N_4041,N_4087);
nand UO_483 (O_483,N_4270,N_4413);
and UO_484 (O_484,N_4285,N_4200);
nor UO_485 (O_485,N_4283,N_4884);
nand UO_486 (O_486,N_4118,N_4776);
or UO_487 (O_487,N_4091,N_4767);
or UO_488 (O_488,N_4292,N_4706);
or UO_489 (O_489,N_4419,N_4672);
nand UO_490 (O_490,N_4982,N_4883);
nor UO_491 (O_491,N_4735,N_4265);
and UO_492 (O_492,N_4024,N_4051);
and UO_493 (O_493,N_4590,N_4535);
or UO_494 (O_494,N_4662,N_4548);
and UO_495 (O_495,N_4394,N_4331);
and UO_496 (O_496,N_4573,N_4588);
nand UO_497 (O_497,N_4084,N_4704);
nor UO_498 (O_498,N_4136,N_4316);
nand UO_499 (O_499,N_4217,N_4054);
or UO_500 (O_500,N_4576,N_4614);
or UO_501 (O_501,N_4936,N_4097);
nand UO_502 (O_502,N_4887,N_4526);
or UO_503 (O_503,N_4187,N_4855);
and UO_504 (O_504,N_4462,N_4999);
nand UO_505 (O_505,N_4125,N_4087);
or UO_506 (O_506,N_4887,N_4100);
xor UO_507 (O_507,N_4868,N_4851);
xor UO_508 (O_508,N_4935,N_4106);
nand UO_509 (O_509,N_4668,N_4598);
nand UO_510 (O_510,N_4376,N_4773);
or UO_511 (O_511,N_4039,N_4639);
nand UO_512 (O_512,N_4176,N_4351);
and UO_513 (O_513,N_4635,N_4951);
nor UO_514 (O_514,N_4806,N_4570);
nor UO_515 (O_515,N_4337,N_4221);
and UO_516 (O_516,N_4082,N_4898);
or UO_517 (O_517,N_4495,N_4551);
nor UO_518 (O_518,N_4202,N_4551);
and UO_519 (O_519,N_4480,N_4705);
or UO_520 (O_520,N_4699,N_4230);
nor UO_521 (O_521,N_4306,N_4904);
nand UO_522 (O_522,N_4576,N_4677);
nand UO_523 (O_523,N_4860,N_4089);
or UO_524 (O_524,N_4524,N_4611);
nor UO_525 (O_525,N_4487,N_4811);
nor UO_526 (O_526,N_4354,N_4983);
and UO_527 (O_527,N_4463,N_4950);
and UO_528 (O_528,N_4249,N_4697);
and UO_529 (O_529,N_4092,N_4938);
nor UO_530 (O_530,N_4335,N_4042);
and UO_531 (O_531,N_4266,N_4766);
nor UO_532 (O_532,N_4874,N_4633);
and UO_533 (O_533,N_4476,N_4744);
nor UO_534 (O_534,N_4602,N_4393);
nand UO_535 (O_535,N_4041,N_4001);
nand UO_536 (O_536,N_4027,N_4082);
and UO_537 (O_537,N_4293,N_4426);
or UO_538 (O_538,N_4906,N_4994);
or UO_539 (O_539,N_4439,N_4674);
or UO_540 (O_540,N_4357,N_4542);
or UO_541 (O_541,N_4820,N_4677);
nand UO_542 (O_542,N_4484,N_4838);
nor UO_543 (O_543,N_4355,N_4027);
or UO_544 (O_544,N_4732,N_4008);
nand UO_545 (O_545,N_4207,N_4921);
nor UO_546 (O_546,N_4083,N_4208);
nand UO_547 (O_547,N_4447,N_4958);
nor UO_548 (O_548,N_4609,N_4983);
nand UO_549 (O_549,N_4033,N_4002);
or UO_550 (O_550,N_4642,N_4056);
nand UO_551 (O_551,N_4898,N_4496);
and UO_552 (O_552,N_4482,N_4064);
or UO_553 (O_553,N_4730,N_4809);
or UO_554 (O_554,N_4165,N_4387);
nor UO_555 (O_555,N_4563,N_4452);
or UO_556 (O_556,N_4161,N_4648);
or UO_557 (O_557,N_4373,N_4022);
nand UO_558 (O_558,N_4775,N_4163);
nor UO_559 (O_559,N_4230,N_4596);
or UO_560 (O_560,N_4911,N_4144);
nor UO_561 (O_561,N_4497,N_4945);
nor UO_562 (O_562,N_4133,N_4222);
and UO_563 (O_563,N_4892,N_4952);
or UO_564 (O_564,N_4374,N_4588);
nand UO_565 (O_565,N_4189,N_4996);
and UO_566 (O_566,N_4526,N_4004);
and UO_567 (O_567,N_4805,N_4462);
nand UO_568 (O_568,N_4822,N_4641);
and UO_569 (O_569,N_4274,N_4660);
nor UO_570 (O_570,N_4461,N_4682);
and UO_571 (O_571,N_4586,N_4789);
nand UO_572 (O_572,N_4940,N_4584);
or UO_573 (O_573,N_4623,N_4220);
nor UO_574 (O_574,N_4347,N_4844);
and UO_575 (O_575,N_4518,N_4922);
nand UO_576 (O_576,N_4730,N_4120);
nor UO_577 (O_577,N_4231,N_4251);
or UO_578 (O_578,N_4211,N_4436);
or UO_579 (O_579,N_4230,N_4490);
nor UO_580 (O_580,N_4794,N_4619);
nand UO_581 (O_581,N_4494,N_4359);
and UO_582 (O_582,N_4058,N_4911);
nand UO_583 (O_583,N_4990,N_4077);
or UO_584 (O_584,N_4519,N_4331);
or UO_585 (O_585,N_4401,N_4411);
or UO_586 (O_586,N_4631,N_4565);
nand UO_587 (O_587,N_4192,N_4305);
xnor UO_588 (O_588,N_4088,N_4464);
nor UO_589 (O_589,N_4412,N_4419);
nor UO_590 (O_590,N_4290,N_4823);
and UO_591 (O_591,N_4350,N_4745);
and UO_592 (O_592,N_4390,N_4951);
and UO_593 (O_593,N_4639,N_4558);
nor UO_594 (O_594,N_4374,N_4948);
nor UO_595 (O_595,N_4961,N_4286);
nor UO_596 (O_596,N_4998,N_4258);
or UO_597 (O_597,N_4796,N_4252);
and UO_598 (O_598,N_4795,N_4891);
and UO_599 (O_599,N_4867,N_4858);
and UO_600 (O_600,N_4128,N_4286);
nor UO_601 (O_601,N_4996,N_4876);
xnor UO_602 (O_602,N_4761,N_4962);
or UO_603 (O_603,N_4893,N_4471);
nor UO_604 (O_604,N_4488,N_4265);
or UO_605 (O_605,N_4622,N_4445);
nand UO_606 (O_606,N_4828,N_4301);
nand UO_607 (O_607,N_4628,N_4178);
nand UO_608 (O_608,N_4731,N_4540);
or UO_609 (O_609,N_4699,N_4514);
nand UO_610 (O_610,N_4927,N_4137);
nand UO_611 (O_611,N_4441,N_4767);
nand UO_612 (O_612,N_4306,N_4924);
nor UO_613 (O_613,N_4303,N_4895);
nand UO_614 (O_614,N_4997,N_4209);
nand UO_615 (O_615,N_4878,N_4329);
nand UO_616 (O_616,N_4277,N_4045);
and UO_617 (O_617,N_4692,N_4614);
or UO_618 (O_618,N_4221,N_4378);
and UO_619 (O_619,N_4865,N_4226);
or UO_620 (O_620,N_4756,N_4409);
or UO_621 (O_621,N_4534,N_4348);
nand UO_622 (O_622,N_4327,N_4655);
or UO_623 (O_623,N_4148,N_4325);
nor UO_624 (O_624,N_4140,N_4839);
and UO_625 (O_625,N_4390,N_4597);
or UO_626 (O_626,N_4182,N_4382);
nand UO_627 (O_627,N_4204,N_4856);
or UO_628 (O_628,N_4277,N_4970);
or UO_629 (O_629,N_4698,N_4062);
nand UO_630 (O_630,N_4332,N_4482);
or UO_631 (O_631,N_4343,N_4239);
nand UO_632 (O_632,N_4449,N_4892);
or UO_633 (O_633,N_4227,N_4772);
and UO_634 (O_634,N_4366,N_4690);
nor UO_635 (O_635,N_4195,N_4723);
nand UO_636 (O_636,N_4980,N_4552);
or UO_637 (O_637,N_4427,N_4400);
or UO_638 (O_638,N_4427,N_4607);
nor UO_639 (O_639,N_4996,N_4602);
nand UO_640 (O_640,N_4187,N_4183);
and UO_641 (O_641,N_4777,N_4132);
or UO_642 (O_642,N_4497,N_4148);
nand UO_643 (O_643,N_4546,N_4477);
nor UO_644 (O_644,N_4782,N_4677);
or UO_645 (O_645,N_4689,N_4362);
nand UO_646 (O_646,N_4430,N_4713);
nor UO_647 (O_647,N_4063,N_4660);
nor UO_648 (O_648,N_4066,N_4271);
and UO_649 (O_649,N_4992,N_4134);
nor UO_650 (O_650,N_4994,N_4160);
nor UO_651 (O_651,N_4161,N_4904);
nand UO_652 (O_652,N_4698,N_4435);
nor UO_653 (O_653,N_4707,N_4958);
and UO_654 (O_654,N_4262,N_4101);
and UO_655 (O_655,N_4288,N_4241);
or UO_656 (O_656,N_4517,N_4611);
nand UO_657 (O_657,N_4817,N_4523);
nor UO_658 (O_658,N_4682,N_4993);
and UO_659 (O_659,N_4186,N_4169);
or UO_660 (O_660,N_4690,N_4992);
nor UO_661 (O_661,N_4808,N_4539);
nand UO_662 (O_662,N_4240,N_4905);
or UO_663 (O_663,N_4307,N_4906);
nand UO_664 (O_664,N_4881,N_4181);
or UO_665 (O_665,N_4321,N_4240);
nor UO_666 (O_666,N_4508,N_4006);
or UO_667 (O_667,N_4196,N_4194);
or UO_668 (O_668,N_4705,N_4978);
or UO_669 (O_669,N_4505,N_4280);
nand UO_670 (O_670,N_4301,N_4899);
nand UO_671 (O_671,N_4202,N_4210);
nor UO_672 (O_672,N_4158,N_4978);
or UO_673 (O_673,N_4121,N_4977);
nand UO_674 (O_674,N_4105,N_4051);
or UO_675 (O_675,N_4887,N_4722);
nand UO_676 (O_676,N_4526,N_4000);
and UO_677 (O_677,N_4213,N_4227);
nand UO_678 (O_678,N_4191,N_4441);
nand UO_679 (O_679,N_4647,N_4068);
and UO_680 (O_680,N_4005,N_4111);
nand UO_681 (O_681,N_4502,N_4025);
or UO_682 (O_682,N_4906,N_4815);
or UO_683 (O_683,N_4998,N_4402);
nand UO_684 (O_684,N_4425,N_4737);
and UO_685 (O_685,N_4740,N_4873);
or UO_686 (O_686,N_4555,N_4219);
and UO_687 (O_687,N_4481,N_4903);
nor UO_688 (O_688,N_4416,N_4628);
and UO_689 (O_689,N_4226,N_4046);
nand UO_690 (O_690,N_4893,N_4126);
and UO_691 (O_691,N_4075,N_4098);
or UO_692 (O_692,N_4941,N_4336);
nand UO_693 (O_693,N_4312,N_4525);
nor UO_694 (O_694,N_4538,N_4419);
nor UO_695 (O_695,N_4939,N_4548);
or UO_696 (O_696,N_4601,N_4917);
nor UO_697 (O_697,N_4974,N_4306);
nand UO_698 (O_698,N_4072,N_4013);
nor UO_699 (O_699,N_4879,N_4343);
nand UO_700 (O_700,N_4066,N_4317);
or UO_701 (O_701,N_4426,N_4496);
nand UO_702 (O_702,N_4685,N_4325);
nor UO_703 (O_703,N_4822,N_4667);
nand UO_704 (O_704,N_4984,N_4074);
nor UO_705 (O_705,N_4785,N_4070);
nand UO_706 (O_706,N_4123,N_4622);
or UO_707 (O_707,N_4167,N_4912);
and UO_708 (O_708,N_4476,N_4865);
and UO_709 (O_709,N_4242,N_4197);
or UO_710 (O_710,N_4820,N_4604);
nor UO_711 (O_711,N_4192,N_4691);
nand UO_712 (O_712,N_4938,N_4703);
nand UO_713 (O_713,N_4697,N_4152);
or UO_714 (O_714,N_4845,N_4785);
and UO_715 (O_715,N_4044,N_4759);
nor UO_716 (O_716,N_4274,N_4232);
nor UO_717 (O_717,N_4527,N_4234);
and UO_718 (O_718,N_4747,N_4817);
or UO_719 (O_719,N_4320,N_4488);
or UO_720 (O_720,N_4495,N_4791);
or UO_721 (O_721,N_4698,N_4344);
nand UO_722 (O_722,N_4253,N_4801);
nor UO_723 (O_723,N_4286,N_4406);
and UO_724 (O_724,N_4958,N_4504);
or UO_725 (O_725,N_4201,N_4296);
nor UO_726 (O_726,N_4278,N_4894);
nand UO_727 (O_727,N_4202,N_4485);
nand UO_728 (O_728,N_4260,N_4074);
or UO_729 (O_729,N_4194,N_4745);
nand UO_730 (O_730,N_4761,N_4788);
nor UO_731 (O_731,N_4077,N_4010);
nor UO_732 (O_732,N_4594,N_4996);
and UO_733 (O_733,N_4235,N_4298);
nand UO_734 (O_734,N_4304,N_4368);
or UO_735 (O_735,N_4969,N_4403);
nand UO_736 (O_736,N_4797,N_4864);
nor UO_737 (O_737,N_4604,N_4487);
nor UO_738 (O_738,N_4364,N_4739);
nand UO_739 (O_739,N_4200,N_4852);
or UO_740 (O_740,N_4431,N_4216);
nand UO_741 (O_741,N_4489,N_4220);
or UO_742 (O_742,N_4214,N_4190);
or UO_743 (O_743,N_4232,N_4959);
and UO_744 (O_744,N_4371,N_4568);
or UO_745 (O_745,N_4493,N_4228);
and UO_746 (O_746,N_4409,N_4961);
and UO_747 (O_747,N_4789,N_4396);
xnor UO_748 (O_748,N_4420,N_4143);
and UO_749 (O_749,N_4301,N_4328);
nor UO_750 (O_750,N_4502,N_4956);
nor UO_751 (O_751,N_4297,N_4021);
nand UO_752 (O_752,N_4380,N_4396);
and UO_753 (O_753,N_4108,N_4941);
nor UO_754 (O_754,N_4601,N_4202);
nand UO_755 (O_755,N_4375,N_4946);
or UO_756 (O_756,N_4068,N_4489);
or UO_757 (O_757,N_4453,N_4474);
nand UO_758 (O_758,N_4891,N_4022);
and UO_759 (O_759,N_4759,N_4836);
and UO_760 (O_760,N_4272,N_4072);
or UO_761 (O_761,N_4412,N_4263);
or UO_762 (O_762,N_4978,N_4496);
nand UO_763 (O_763,N_4993,N_4890);
nor UO_764 (O_764,N_4290,N_4196);
nand UO_765 (O_765,N_4613,N_4382);
nor UO_766 (O_766,N_4114,N_4140);
or UO_767 (O_767,N_4885,N_4890);
nor UO_768 (O_768,N_4530,N_4109);
and UO_769 (O_769,N_4480,N_4053);
nand UO_770 (O_770,N_4181,N_4413);
nand UO_771 (O_771,N_4353,N_4280);
nor UO_772 (O_772,N_4154,N_4031);
nand UO_773 (O_773,N_4526,N_4922);
and UO_774 (O_774,N_4355,N_4806);
and UO_775 (O_775,N_4536,N_4839);
and UO_776 (O_776,N_4488,N_4465);
xnor UO_777 (O_777,N_4533,N_4416);
nand UO_778 (O_778,N_4647,N_4025);
or UO_779 (O_779,N_4296,N_4705);
nand UO_780 (O_780,N_4558,N_4910);
nor UO_781 (O_781,N_4021,N_4513);
nand UO_782 (O_782,N_4865,N_4146);
nor UO_783 (O_783,N_4248,N_4857);
nor UO_784 (O_784,N_4286,N_4615);
or UO_785 (O_785,N_4047,N_4734);
and UO_786 (O_786,N_4136,N_4529);
nor UO_787 (O_787,N_4231,N_4040);
or UO_788 (O_788,N_4416,N_4220);
nor UO_789 (O_789,N_4445,N_4040);
and UO_790 (O_790,N_4336,N_4294);
nand UO_791 (O_791,N_4567,N_4155);
nor UO_792 (O_792,N_4741,N_4081);
and UO_793 (O_793,N_4805,N_4493);
xor UO_794 (O_794,N_4636,N_4816);
nand UO_795 (O_795,N_4236,N_4049);
and UO_796 (O_796,N_4752,N_4361);
or UO_797 (O_797,N_4885,N_4949);
nor UO_798 (O_798,N_4005,N_4838);
nor UO_799 (O_799,N_4396,N_4600);
nor UO_800 (O_800,N_4357,N_4656);
and UO_801 (O_801,N_4655,N_4068);
nand UO_802 (O_802,N_4478,N_4705);
nand UO_803 (O_803,N_4943,N_4255);
nand UO_804 (O_804,N_4021,N_4974);
and UO_805 (O_805,N_4402,N_4364);
nand UO_806 (O_806,N_4853,N_4196);
nor UO_807 (O_807,N_4922,N_4277);
and UO_808 (O_808,N_4591,N_4707);
and UO_809 (O_809,N_4370,N_4520);
nand UO_810 (O_810,N_4302,N_4476);
nor UO_811 (O_811,N_4678,N_4774);
or UO_812 (O_812,N_4970,N_4482);
and UO_813 (O_813,N_4323,N_4094);
nand UO_814 (O_814,N_4296,N_4457);
nand UO_815 (O_815,N_4886,N_4640);
nor UO_816 (O_816,N_4872,N_4495);
nand UO_817 (O_817,N_4598,N_4200);
or UO_818 (O_818,N_4220,N_4129);
nand UO_819 (O_819,N_4907,N_4908);
nor UO_820 (O_820,N_4583,N_4831);
nand UO_821 (O_821,N_4940,N_4460);
and UO_822 (O_822,N_4802,N_4464);
nand UO_823 (O_823,N_4040,N_4186);
nand UO_824 (O_824,N_4503,N_4059);
nand UO_825 (O_825,N_4654,N_4363);
nand UO_826 (O_826,N_4947,N_4691);
nor UO_827 (O_827,N_4732,N_4603);
and UO_828 (O_828,N_4900,N_4388);
or UO_829 (O_829,N_4475,N_4589);
and UO_830 (O_830,N_4169,N_4380);
and UO_831 (O_831,N_4193,N_4530);
and UO_832 (O_832,N_4400,N_4509);
nor UO_833 (O_833,N_4752,N_4249);
or UO_834 (O_834,N_4403,N_4215);
nor UO_835 (O_835,N_4454,N_4762);
nor UO_836 (O_836,N_4354,N_4281);
nor UO_837 (O_837,N_4105,N_4989);
nor UO_838 (O_838,N_4010,N_4045);
or UO_839 (O_839,N_4860,N_4349);
nor UO_840 (O_840,N_4689,N_4477);
or UO_841 (O_841,N_4992,N_4013);
and UO_842 (O_842,N_4531,N_4692);
nand UO_843 (O_843,N_4087,N_4238);
or UO_844 (O_844,N_4376,N_4407);
nor UO_845 (O_845,N_4110,N_4547);
nand UO_846 (O_846,N_4839,N_4297);
or UO_847 (O_847,N_4247,N_4211);
nand UO_848 (O_848,N_4616,N_4398);
or UO_849 (O_849,N_4718,N_4381);
nand UO_850 (O_850,N_4524,N_4857);
and UO_851 (O_851,N_4749,N_4659);
and UO_852 (O_852,N_4568,N_4904);
or UO_853 (O_853,N_4825,N_4922);
and UO_854 (O_854,N_4456,N_4176);
or UO_855 (O_855,N_4660,N_4940);
nor UO_856 (O_856,N_4424,N_4200);
nor UO_857 (O_857,N_4399,N_4957);
nand UO_858 (O_858,N_4300,N_4165);
nor UO_859 (O_859,N_4653,N_4723);
or UO_860 (O_860,N_4523,N_4274);
nor UO_861 (O_861,N_4838,N_4187);
and UO_862 (O_862,N_4714,N_4703);
and UO_863 (O_863,N_4810,N_4598);
nor UO_864 (O_864,N_4636,N_4364);
nand UO_865 (O_865,N_4211,N_4210);
xor UO_866 (O_866,N_4727,N_4691);
nand UO_867 (O_867,N_4207,N_4874);
nor UO_868 (O_868,N_4493,N_4327);
or UO_869 (O_869,N_4427,N_4548);
or UO_870 (O_870,N_4662,N_4009);
nand UO_871 (O_871,N_4351,N_4675);
or UO_872 (O_872,N_4093,N_4240);
and UO_873 (O_873,N_4007,N_4113);
nor UO_874 (O_874,N_4117,N_4206);
and UO_875 (O_875,N_4318,N_4639);
nor UO_876 (O_876,N_4143,N_4116);
xnor UO_877 (O_877,N_4305,N_4684);
or UO_878 (O_878,N_4692,N_4250);
nor UO_879 (O_879,N_4431,N_4923);
or UO_880 (O_880,N_4312,N_4357);
nand UO_881 (O_881,N_4628,N_4439);
and UO_882 (O_882,N_4933,N_4422);
xnor UO_883 (O_883,N_4580,N_4472);
nand UO_884 (O_884,N_4761,N_4309);
nor UO_885 (O_885,N_4736,N_4439);
nor UO_886 (O_886,N_4444,N_4953);
or UO_887 (O_887,N_4735,N_4796);
nor UO_888 (O_888,N_4372,N_4593);
nand UO_889 (O_889,N_4298,N_4083);
and UO_890 (O_890,N_4046,N_4047);
and UO_891 (O_891,N_4770,N_4514);
nor UO_892 (O_892,N_4573,N_4972);
or UO_893 (O_893,N_4466,N_4817);
nor UO_894 (O_894,N_4141,N_4738);
nand UO_895 (O_895,N_4750,N_4627);
nand UO_896 (O_896,N_4162,N_4203);
nand UO_897 (O_897,N_4385,N_4025);
or UO_898 (O_898,N_4195,N_4139);
or UO_899 (O_899,N_4444,N_4748);
and UO_900 (O_900,N_4834,N_4390);
nand UO_901 (O_901,N_4949,N_4581);
or UO_902 (O_902,N_4792,N_4047);
xor UO_903 (O_903,N_4757,N_4351);
nor UO_904 (O_904,N_4267,N_4413);
and UO_905 (O_905,N_4359,N_4393);
and UO_906 (O_906,N_4633,N_4439);
or UO_907 (O_907,N_4454,N_4490);
nor UO_908 (O_908,N_4837,N_4179);
nand UO_909 (O_909,N_4800,N_4751);
and UO_910 (O_910,N_4139,N_4232);
nor UO_911 (O_911,N_4605,N_4230);
nor UO_912 (O_912,N_4506,N_4542);
nor UO_913 (O_913,N_4530,N_4084);
and UO_914 (O_914,N_4449,N_4719);
nor UO_915 (O_915,N_4830,N_4966);
nand UO_916 (O_916,N_4320,N_4000);
nand UO_917 (O_917,N_4601,N_4980);
xor UO_918 (O_918,N_4051,N_4710);
nor UO_919 (O_919,N_4446,N_4277);
and UO_920 (O_920,N_4362,N_4075);
and UO_921 (O_921,N_4154,N_4697);
nand UO_922 (O_922,N_4822,N_4824);
and UO_923 (O_923,N_4793,N_4670);
or UO_924 (O_924,N_4533,N_4124);
nand UO_925 (O_925,N_4460,N_4768);
nand UO_926 (O_926,N_4540,N_4002);
nand UO_927 (O_927,N_4005,N_4554);
nor UO_928 (O_928,N_4356,N_4345);
nor UO_929 (O_929,N_4329,N_4706);
nand UO_930 (O_930,N_4826,N_4766);
nand UO_931 (O_931,N_4331,N_4830);
nor UO_932 (O_932,N_4299,N_4141);
nand UO_933 (O_933,N_4771,N_4515);
xor UO_934 (O_934,N_4098,N_4594);
and UO_935 (O_935,N_4090,N_4765);
nor UO_936 (O_936,N_4817,N_4863);
or UO_937 (O_937,N_4713,N_4546);
or UO_938 (O_938,N_4939,N_4122);
and UO_939 (O_939,N_4203,N_4132);
and UO_940 (O_940,N_4404,N_4134);
nor UO_941 (O_941,N_4391,N_4671);
and UO_942 (O_942,N_4674,N_4177);
nand UO_943 (O_943,N_4839,N_4443);
or UO_944 (O_944,N_4581,N_4552);
or UO_945 (O_945,N_4356,N_4917);
and UO_946 (O_946,N_4645,N_4718);
and UO_947 (O_947,N_4247,N_4322);
nor UO_948 (O_948,N_4241,N_4304);
xor UO_949 (O_949,N_4436,N_4485);
nand UO_950 (O_950,N_4236,N_4496);
and UO_951 (O_951,N_4052,N_4145);
and UO_952 (O_952,N_4429,N_4576);
nor UO_953 (O_953,N_4801,N_4453);
nor UO_954 (O_954,N_4763,N_4305);
nand UO_955 (O_955,N_4797,N_4577);
nand UO_956 (O_956,N_4386,N_4211);
or UO_957 (O_957,N_4968,N_4379);
nor UO_958 (O_958,N_4423,N_4364);
and UO_959 (O_959,N_4623,N_4573);
and UO_960 (O_960,N_4031,N_4392);
nand UO_961 (O_961,N_4193,N_4127);
xnor UO_962 (O_962,N_4133,N_4678);
or UO_963 (O_963,N_4586,N_4607);
or UO_964 (O_964,N_4778,N_4159);
or UO_965 (O_965,N_4248,N_4556);
nor UO_966 (O_966,N_4105,N_4660);
or UO_967 (O_967,N_4283,N_4201);
nand UO_968 (O_968,N_4595,N_4853);
or UO_969 (O_969,N_4757,N_4619);
nor UO_970 (O_970,N_4213,N_4724);
or UO_971 (O_971,N_4137,N_4297);
nor UO_972 (O_972,N_4991,N_4599);
or UO_973 (O_973,N_4982,N_4042);
or UO_974 (O_974,N_4613,N_4047);
and UO_975 (O_975,N_4468,N_4814);
nand UO_976 (O_976,N_4865,N_4530);
or UO_977 (O_977,N_4008,N_4813);
or UO_978 (O_978,N_4610,N_4645);
nor UO_979 (O_979,N_4215,N_4735);
and UO_980 (O_980,N_4573,N_4279);
nand UO_981 (O_981,N_4853,N_4796);
and UO_982 (O_982,N_4401,N_4225);
nand UO_983 (O_983,N_4952,N_4189);
and UO_984 (O_984,N_4786,N_4776);
or UO_985 (O_985,N_4769,N_4486);
nand UO_986 (O_986,N_4164,N_4084);
nor UO_987 (O_987,N_4430,N_4738);
and UO_988 (O_988,N_4788,N_4182);
nor UO_989 (O_989,N_4610,N_4643);
and UO_990 (O_990,N_4660,N_4411);
and UO_991 (O_991,N_4975,N_4758);
and UO_992 (O_992,N_4535,N_4144);
or UO_993 (O_993,N_4680,N_4705);
nand UO_994 (O_994,N_4141,N_4994);
and UO_995 (O_995,N_4167,N_4573);
nor UO_996 (O_996,N_4350,N_4001);
nor UO_997 (O_997,N_4291,N_4684);
or UO_998 (O_998,N_4221,N_4799);
nand UO_999 (O_999,N_4065,N_4055);
endmodule