module basic_2500_25000_3000_10_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_2128,In_357);
or U1 (N_1,In_110,In_2393);
nor U2 (N_2,In_342,In_1041);
nor U3 (N_3,In_734,In_1535);
and U4 (N_4,In_1264,In_864);
or U5 (N_5,In_1141,In_1721);
nand U6 (N_6,In_1104,In_2295);
or U7 (N_7,In_788,In_1150);
and U8 (N_8,In_1910,In_33);
xnor U9 (N_9,In_1094,In_1427);
nor U10 (N_10,In_2084,In_1415);
nand U11 (N_11,In_438,In_1877);
and U12 (N_12,In_486,In_1968);
and U13 (N_13,In_1582,In_2306);
or U14 (N_14,In_254,In_1078);
nor U15 (N_15,In_896,In_1620);
nor U16 (N_16,In_759,In_525);
nand U17 (N_17,In_693,In_2422);
nand U18 (N_18,In_284,In_395);
nor U19 (N_19,In_1419,In_1562);
nand U20 (N_20,In_2257,In_1510);
xor U21 (N_21,In_546,In_2056);
nor U22 (N_22,In_1011,In_1730);
and U23 (N_23,In_2485,In_1692);
and U24 (N_24,In_1956,In_2308);
nand U25 (N_25,In_1804,In_1564);
and U26 (N_26,In_2279,In_1318);
nand U27 (N_27,In_1227,In_1711);
xnor U28 (N_28,In_823,In_319);
xor U29 (N_29,In_1075,In_1890);
nor U30 (N_30,In_2112,In_1892);
or U31 (N_31,In_1256,In_54);
nand U32 (N_32,In_819,In_905);
and U33 (N_33,In_1845,In_185);
or U34 (N_34,In_2424,In_1604);
nor U35 (N_35,In_1611,In_1600);
and U36 (N_36,In_2102,In_692);
or U37 (N_37,In_1576,In_1990);
or U38 (N_38,In_721,In_2009);
and U39 (N_39,In_296,In_1848);
and U40 (N_40,In_850,In_746);
nand U41 (N_41,In_1004,In_423);
nor U42 (N_42,In_573,In_2367);
or U43 (N_43,In_1856,In_786);
nor U44 (N_44,In_508,In_1977);
xnor U45 (N_45,In_1158,In_1667);
and U46 (N_46,In_93,In_455);
or U47 (N_47,In_38,In_2234);
nand U48 (N_48,In_2423,In_1286);
nand U49 (N_49,In_410,In_1393);
nor U50 (N_50,In_1097,In_1043);
nand U51 (N_51,In_2085,In_876);
xor U52 (N_52,In_676,In_50);
xnor U53 (N_53,In_750,In_2473);
xor U54 (N_54,In_49,In_1112);
or U55 (N_55,In_2203,In_2125);
nor U56 (N_56,In_725,In_190);
or U57 (N_57,In_2383,In_944);
nor U58 (N_58,In_1357,In_1241);
or U59 (N_59,In_2478,In_86);
and U60 (N_60,In_394,In_368);
nand U61 (N_61,In_527,In_1223);
xor U62 (N_62,In_1090,In_2205);
nand U63 (N_63,In_2036,In_1450);
or U64 (N_64,In_581,In_562);
nor U65 (N_65,In_1115,In_1009);
and U66 (N_66,In_1735,In_1580);
nor U67 (N_67,In_1723,In_891);
xnor U68 (N_68,In_2122,In_1777);
or U69 (N_69,In_640,In_2280);
and U70 (N_70,In_208,In_1740);
nand U71 (N_71,In_200,In_334);
nand U72 (N_72,In_658,In_990);
nand U73 (N_73,In_491,In_1146);
xor U74 (N_74,In_881,In_2208);
and U75 (N_75,In_2063,In_2090);
or U76 (N_76,In_2166,In_1841);
xor U77 (N_77,In_2227,In_1581);
or U78 (N_78,In_1032,In_2159);
nand U79 (N_79,In_417,In_2161);
and U80 (N_80,In_1081,In_1317);
and U81 (N_81,In_187,In_1280);
nand U82 (N_82,In_605,In_1636);
nand U83 (N_83,In_1125,In_2369);
or U84 (N_84,In_2148,In_660);
nor U85 (N_85,In_579,In_1034);
nor U86 (N_86,In_463,In_1706);
or U87 (N_87,In_1861,In_9);
nand U88 (N_88,In_1356,In_530);
nor U89 (N_89,In_1281,In_2034);
nor U90 (N_90,In_2456,In_94);
or U91 (N_91,In_2450,In_739);
nor U92 (N_92,In_2150,In_1405);
xnor U93 (N_93,In_2167,In_2057);
xor U94 (N_94,In_726,In_2066);
or U95 (N_95,In_1132,In_1635);
and U96 (N_96,In_1336,In_415);
or U97 (N_97,In_2300,In_413);
nor U98 (N_98,In_481,In_2312);
nor U99 (N_99,In_1020,In_89);
nor U100 (N_100,In_576,In_569);
and U101 (N_101,In_2173,In_1451);
nand U102 (N_102,In_470,In_419);
nand U103 (N_103,In_362,In_162);
nor U104 (N_104,In_1985,In_1271);
nor U105 (N_105,In_1443,In_1481);
nor U106 (N_106,In_754,In_697);
nor U107 (N_107,In_2024,In_2105);
or U108 (N_108,In_426,In_1249);
and U109 (N_109,In_2183,In_2322);
nand U110 (N_110,In_1549,In_442);
and U111 (N_111,In_2494,In_1261);
nand U112 (N_112,In_965,In_1325);
xnor U113 (N_113,In_2339,In_1616);
or U114 (N_114,In_2490,In_1370);
and U115 (N_115,In_2468,In_1805);
nor U116 (N_116,In_281,In_260);
xor U117 (N_117,In_854,In_996);
and U118 (N_118,In_580,In_1755);
xnor U119 (N_119,In_1683,In_425);
and U120 (N_120,In_2427,In_2259);
nor U121 (N_121,In_1769,In_1203);
or U122 (N_122,In_288,In_351);
or U123 (N_123,In_150,In_774);
xor U124 (N_124,In_1137,In_2343);
nand U125 (N_125,In_1063,In_540);
nor U126 (N_126,In_2398,In_1434);
and U127 (N_127,In_1901,In_2470);
xnor U128 (N_128,In_2457,In_632);
nand U129 (N_129,In_364,In_1383);
or U130 (N_130,In_495,In_2239);
and U131 (N_131,In_521,In_1028);
nand U132 (N_132,In_1821,In_129);
nor U133 (N_133,In_259,In_1399);
or U134 (N_134,In_1416,In_1029);
xor U135 (N_135,In_636,In_2083);
or U136 (N_136,In_873,In_1529);
or U137 (N_137,In_517,In_720);
nand U138 (N_138,In_1829,In_1301);
nand U139 (N_139,In_2124,In_1888);
or U140 (N_140,In_1152,In_1536);
xor U141 (N_141,In_1088,In_2484);
and U142 (N_142,In_704,In_2314);
nand U143 (N_143,In_700,In_1981);
and U144 (N_144,In_299,In_1646);
or U145 (N_145,In_336,In_2168);
or U146 (N_146,In_1147,In_1543);
nand U147 (N_147,In_1190,In_287);
nor U148 (N_148,In_890,In_1698);
nand U149 (N_149,In_2164,In_1639);
nand U150 (N_150,In_1082,In_166);
xnor U151 (N_151,In_144,In_432);
or U152 (N_152,In_1052,In_1423);
or U153 (N_153,In_1701,In_1362);
nand U154 (N_154,In_225,In_329);
xnor U155 (N_155,In_2242,In_1975);
and U156 (N_156,In_16,In_1970);
nand U157 (N_157,In_2170,In_1313);
xnor U158 (N_158,In_1632,In_724);
or U159 (N_159,In_1940,In_679);
or U160 (N_160,In_651,In_2100);
and U161 (N_161,In_1103,In_1629);
or U162 (N_162,In_2440,In_258);
or U163 (N_163,In_2345,In_1623);
and U164 (N_164,In_1793,In_743);
or U165 (N_165,In_1656,In_2233);
nor U166 (N_166,In_39,In_1479);
nor U167 (N_167,In_2237,In_169);
nor U168 (N_168,In_51,In_1534);
nand U169 (N_169,In_2176,In_1111);
or U170 (N_170,In_807,In_1284);
xor U171 (N_171,In_1889,In_857);
and U172 (N_172,In_184,In_353);
nand U173 (N_173,In_1411,In_1380);
nor U174 (N_174,In_2248,In_1283);
or U175 (N_175,In_1588,In_1236);
or U176 (N_176,In_1074,In_1798);
xnor U177 (N_177,In_1538,In_1684);
or U178 (N_178,In_23,In_469);
nor U179 (N_179,In_1678,In_1893);
xor U180 (N_180,In_1900,In_1060);
or U181 (N_181,In_1748,In_2344);
nand U182 (N_182,In_99,In_1865);
xor U183 (N_183,In_584,In_279);
or U184 (N_184,In_65,In_2048);
xnor U185 (N_185,In_454,In_1106);
or U186 (N_186,In_793,In_1351);
nor U187 (N_187,In_796,In_1225);
xor U188 (N_188,In_1941,In_2191);
or U189 (N_189,In_108,In_783);
and U190 (N_190,In_1929,In_1922);
and U191 (N_191,In_2018,In_1775);
nand U192 (N_192,In_338,In_799);
nor U193 (N_193,In_1187,In_993);
and U194 (N_194,In_804,In_252);
nor U195 (N_195,In_1188,In_1213);
and U196 (N_196,In_2082,In_1566);
nor U197 (N_197,In_1191,In_2454);
xnor U198 (N_198,In_1988,In_2416);
xnor U199 (N_199,In_2304,In_775);
nor U200 (N_200,In_1521,In_2462);
nor U201 (N_201,In_2061,In_1686);
xnor U202 (N_202,In_1739,In_749);
xor U203 (N_203,In_1100,In_1449);
nand U204 (N_204,In_106,In_677);
or U205 (N_205,In_979,In_1770);
or U206 (N_206,In_1853,In_1453);
nor U207 (N_207,In_1499,In_479);
nand U208 (N_208,In_852,In_1989);
or U209 (N_209,In_1508,In_1007);
nor U210 (N_210,In_1110,In_808);
nand U211 (N_211,In_303,In_963);
xor U212 (N_212,In_1816,In_2118);
xor U213 (N_213,In_1420,In_85);
nor U214 (N_214,In_1824,In_1209);
or U215 (N_215,In_790,In_2436);
xnor U216 (N_216,In_1477,In_1161);
or U217 (N_217,In_1745,In_2178);
nor U218 (N_218,In_191,In_1354);
nor U219 (N_219,In_1350,In_203);
nand U220 (N_220,In_1355,In_2253);
xnor U221 (N_221,In_949,In_1907);
and U222 (N_222,In_2390,In_639);
nand U223 (N_223,In_2111,In_2324);
xor U224 (N_224,In_1307,In_1918);
or U225 (N_225,In_966,In_459);
or U226 (N_226,In_1488,In_1466);
or U227 (N_227,In_1118,In_1114);
or U228 (N_228,In_2081,In_585);
xnor U229 (N_229,In_1098,In_533);
and U230 (N_230,In_510,In_895);
nand U231 (N_231,In_1234,In_923);
nor U232 (N_232,In_451,In_2165);
or U233 (N_233,In_2493,In_1432);
nand U234 (N_234,In_142,In_2220);
nor U235 (N_235,In_452,In_1906);
nor U236 (N_236,In_1182,In_1064);
nor U237 (N_237,In_172,In_275);
or U238 (N_238,In_812,In_645);
and U239 (N_239,In_1257,In_2350);
nand U240 (N_240,In_1135,In_1145);
xor U241 (N_241,In_2366,In_877);
nand U242 (N_242,In_1168,In_2192);
nor U243 (N_243,In_331,In_1596);
nor U244 (N_244,In_907,In_1612);
and U245 (N_245,In_936,In_251);
nand U246 (N_246,In_1278,In_557);
and U247 (N_247,In_524,In_1820);
or U248 (N_248,In_1859,In_407);
xnor U249 (N_249,In_1177,In_1672);
and U250 (N_250,In_2041,In_2087);
nand U251 (N_251,In_816,In_1838);
xor U252 (N_252,In_1458,In_1676);
nor U253 (N_253,In_2264,In_1523);
nor U254 (N_254,In_1468,In_1130);
and U255 (N_255,In_2254,In_1050);
or U256 (N_256,In_542,In_305);
or U257 (N_257,In_2269,In_1167);
xor U258 (N_258,In_128,In_732);
nand U259 (N_259,In_1903,In_95);
and U260 (N_260,In_1830,In_2483);
and U261 (N_261,In_929,In_602);
xor U262 (N_262,In_125,In_1323);
xnor U263 (N_263,In_1952,In_738);
or U264 (N_264,In_1418,In_1899);
nor U265 (N_265,In_682,In_96);
nor U266 (N_266,In_274,In_780);
or U267 (N_267,In_2160,In_827);
nor U268 (N_268,In_483,In_1183);
or U269 (N_269,In_863,In_2311);
and U270 (N_270,In_1270,In_1377);
xnor U271 (N_271,In_430,In_712);
or U272 (N_272,In_1300,In_803);
or U273 (N_273,In_1487,In_104);
nand U274 (N_274,In_587,In_1069);
nand U275 (N_275,In_2005,In_1665);
nor U276 (N_276,In_371,In_1363);
nor U277 (N_277,In_1882,In_1799);
nand U278 (N_278,In_1659,In_885);
nand U279 (N_279,In_2114,In_1996);
or U280 (N_280,In_1983,In_77);
nor U281 (N_281,In_56,In_1012);
and U282 (N_282,In_942,In_691);
nor U283 (N_283,In_293,In_868);
nand U284 (N_284,In_15,In_2219);
nand U285 (N_285,In_2467,In_897);
nand U286 (N_286,In_814,In_1444);
xor U287 (N_287,In_1083,In_1429);
or U288 (N_288,In_26,In_53);
nand U289 (N_289,In_1279,In_1459);
nor U290 (N_290,In_1540,In_969);
nand U291 (N_291,In_887,In_2400);
nor U292 (N_292,In_2039,In_2241);
xnor U293 (N_293,In_2000,In_647);
nor U294 (N_294,In_625,In_2073);
nor U295 (N_295,In_2333,In_2397);
nor U296 (N_296,In_1276,In_131);
nand U297 (N_297,In_286,In_1606);
or U298 (N_298,In_773,In_559);
and U299 (N_299,In_867,In_2441);
nand U300 (N_300,In_127,In_1719);
and U301 (N_301,In_219,In_2007);
or U302 (N_302,In_291,In_1265);
nand U303 (N_303,In_927,In_1093);
or U304 (N_304,In_1653,In_729);
nand U305 (N_305,In_2271,In_839);
nor U306 (N_306,In_307,In_1781);
nand U307 (N_307,In_2135,In_1197);
nand U308 (N_308,In_809,In_1785);
xor U309 (N_309,In_1320,In_2052);
xor U310 (N_310,In_244,In_63);
xor U311 (N_311,In_256,In_789);
nand U312 (N_312,In_1762,In_2446);
nor U313 (N_313,In_1019,In_1978);
and U314 (N_314,In_1868,In_1953);
xor U315 (N_315,In_18,In_1976);
xor U316 (N_316,In_711,In_1319);
nand U317 (N_317,In_2348,In_263);
nor U318 (N_318,In_13,In_2449);
and U319 (N_319,In_741,In_1341);
nor U320 (N_320,In_1396,In_1085);
and U321 (N_321,In_447,In_1916);
nand U322 (N_322,In_1476,In_1718);
xnor U323 (N_323,In_669,In_2117);
and U324 (N_324,In_2008,In_114);
or U325 (N_325,In_1537,In_1036);
and U326 (N_326,In_2182,In_2051);
nand U327 (N_327,In_363,In_1303);
or U328 (N_328,In_935,In_1920);
nor U329 (N_329,In_2194,In_1293);
or U330 (N_330,In_843,In_2316);
or U331 (N_331,In_2381,In_2079);
or U332 (N_332,In_1483,In_6);
or U333 (N_333,In_44,In_1517);
and U334 (N_334,In_683,In_380);
nand U335 (N_335,In_1758,In_1206);
xor U336 (N_336,In_1601,In_2472);
nand U337 (N_337,In_332,In_234);
xnor U338 (N_338,In_235,In_543);
nand U339 (N_339,In_341,In_986);
xnor U340 (N_340,In_1773,In_2213);
xor U341 (N_341,In_629,In_242);
or U342 (N_342,In_1169,In_80);
nor U343 (N_343,In_1710,In_2101);
xnor U344 (N_344,In_462,In_1017);
nand U345 (N_345,In_2266,In_1447);
xor U346 (N_346,In_502,In_2228);
xnor U347 (N_347,In_1473,In_1475);
or U348 (N_348,In_2292,In_285);
or U349 (N_349,In_1984,In_1251);
and U350 (N_350,In_1084,In_2064);
nor U351 (N_351,In_1259,In_2389);
or U352 (N_352,In_1024,In_2133);
and U353 (N_353,In_1035,In_321);
xnor U354 (N_354,In_2108,In_1732);
nor U355 (N_355,In_312,In_1008);
nor U356 (N_356,In_2116,In_2238);
nand U357 (N_357,In_811,In_504);
xor U358 (N_358,In_1408,In_500);
nand U359 (N_359,In_141,In_795);
nor U360 (N_360,In_1156,In_690);
nor U361 (N_361,In_798,In_678);
xnor U362 (N_362,In_1912,In_390);
nand U363 (N_363,In_236,In_1018);
or U364 (N_364,In_1042,In_1682);
nor U365 (N_365,In_1885,In_201);
xor U366 (N_366,In_1496,In_1438);
and U367 (N_367,In_1954,In_1511);
nand U368 (N_368,In_1772,In_506);
nor U369 (N_369,In_914,In_392);
nor U370 (N_370,In_2169,In_424);
nand U371 (N_371,In_1717,In_2226);
or U372 (N_372,In_673,In_1224);
and U373 (N_373,In_2268,In_2492);
xor U374 (N_374,In_2476,In_1237);
nand U375 (N_375,In_1938,In_615);
or U376 (N_376,In_822,In_352);
nand U377 (N_377,In_2037,In_177);
and U378 (N_378,In_1514,In_633);
nor U379 (N_379,In_1797,In_1911);
or U380 (N_380,In_2442,In_1609);
nor U381 (N_381,In_590,In_46);
or U382 (N_382,In_431,In_994);
nor U383 (N_383,In_889,In_461);
or U384 (N_384,In_1054,In_1960);
xnor U385 (N_385,In_1179,In_1253);
nand U386 (N_386,In_689,In_784);
and U387 (N_387,In_1121,In_1555);
nor U388 (N_388,In_474,In_978);
xnor U389 (N_389,In_1851,In_670);
and U390 (N_390,In_2179,In_2359);
nor U391 (N_391,In_1352,In_1460);
nor U392 (N_392,In_1565,In_70);
or U393 (N_393,In_1812,In_1749);
or U394 (N_394,In_1518,In_2458);
and U395 (N_395,In_544,In_206);
xor U396 (N_396,In_345,In_952);
or U397 (N_397,In_1136,In_1490);
or U398 (N_398,In_2362,In_2255);
xnor U399 (N_399,In_2099,In_627);
or U400 (N_400,In_1801,In_523);
or U401 (N_401,In_1747,In_2187);
nor U402 (N_402,In_947,In_381);
nor U403 (N_403,In_1057,In_115);
nand U404 (N_404,In_320,In_901);
xor U405 (N_405,In_1171,In_964);
nor U406 (N_406,In_1212,In_1462);
or U407 (N_407,In_249,In_1248);
or U408 (N_408,In_2055,In_358);
xor U409 (N_409,In_2399,In_866);
xor U410 (N_410,In_865,In_1578);
nand U411 (N_411,In_1010,In_1969);
nand U412 (N_412,In_1869,In_72);
and U413 (N_413,In_975,In_2469);
and U414 (N_414,In_2258,In_1982);
and U415 (N_415,In_21,In_2368);
and U416 (N_416,In_117,In_2356);
xor U417 (N_417,In_2092,In_103);
or U418 (N_418,In_1108,In_3);
or U419 (N_419,In_1379,In_253);
xor U420 (N_420,In_40,In_1633);
nor U421 (N_421,In_1592,In_1756);
nand U422 (N_422,In_982,In_4);
xnor U423 (N_423,In_2282,In_1767);
xor U424 (N_424,In_718,In_2156);
or U425 (N_425,In_83,In_1229);
or U426 (N_426,In_1016,In_2218);
nor U427 (N_427,In_988,In_1788);
and U428 (N_428,In_499,In_385);
nand U429 (N_429,In_372,In_1005);
nand U430 (N_430,In_2001,In_448);
or U431 (N_431,In_1180,In_1298);
xnor U432 (N_432,In_204,In_1129);
and U433 (N_433,In_482,In_1840);
or U434 (N_434,In_2405,In_326);
or U435 (N_435,In_195,In_176);
nor U436 (N_436,In_1149,In_346);
xnor U437 (N_437,In_2412,In_1096);
or U438 (N_438,In_904,In_1366);
nand U439 (N_439,In_2331,In_1328);
nor U440 (N_440,In_2070,In_421);
and U441 (N_441,In_548,In_250);
nand U442 (N_442,In_551,In_2106);
or U443 (N_443,In_912,In_1172);
and U444 (N_444,In_84,In_1049);
xor U445 (N_445,In_731,In_597);
nor U446 (N_446,In_282,In_1768);
nand U447 (N_447,In_384,In_2236);
and U448 (N_448,In_1673,In_411);
xnor U449 (N_449,In_1406,In_902);
or U450 (N_450,In_1160,In_958);
nor U451 (N_451,In_939,In_2223);
nor U452 (N_452,In_503,In_140);
nand U453 (N_453,In_1000,In_2270);
nand U454 (N_454,In_1232,In_1071);
nor U455 (N_455,In_1943,In_648);
nand U456 (N_456,In_674,In_1857);
xor U457 (N_457,In_715,In_1963);
and U458 (N_458,In_240,In_2360);
xor U459 (N_459,In_324,In_1515);
nor U460 (N_460,In_492,In_1095);
nor U461 (N_461,In_107,In_122);
nor U462 (N_462,In_2216,In_1478);
nor U463 (N_463,In_2050,In_1046);
nand U464 (N_464,In_2038,In_2317);
and U465 (N_465,In_1441,In_2373);
nand U466 (N_466,In_552,In_133);
xor U467 (N_467,In_2355,In_2157);
nand U468 (N_468,In_1372,In_389);
nand U469 (N_469,In_2047,In_1860);
nor U470 (N_470,In_566,In_1647);
nor U471 (N_471,In_1999,In_1586);
xor U472 (N_472,In_2026,In_1164);
nand U473 (N_473,In_1512,In_2141);
and U474 (N_474,In_1624,In_2217);
xor U475 (N_475,In_1198,In_671);
nand U476 (N_476,In_834,In_100);
xnor U477 (N_477,In_498,In_374);
or U478 (N_478,In_649,In_1597);
nand U479 (N_479,In_1944,In_2013);
nor U480 (N_480,In_1200,In_1573);
nor U481 (N_481,In_1353,In_2480);
or U482 (N_482,In_1503,In_59);
xor U483 (N_483,In_2154,In_22);
or U484 (N_484,In_1827,In_2021);
nand U485 (N_485,In_1734,In_1077);
nor U486 (N_486,In_913,In_1163);
nand U487 (N_487,In_105,In_268);
xnor U488 (N_488,In_1329,In_1087);
nor U489 (N_489,In_2302,In_875);
or U490 (N_490,In_170,In_337);
or U491 (N_491,In_1384,In_2175);
and U492 (N_492,In_2411,In_1282);
xor U493 (N_493,In_1634,In_1359);
and U494 (N_494,In_1022,In_62);
nand U495 (N_495,In_1516,In_393);
and U496 (N_496,In_132,In_1737);
or U497 (N_497,In_1658,In_227);
nor U498 (N_498,In_2303,In_2380);
nand U499 (N_499,In_2463,In_160);
xnor U500 (N_500,In_932,In_592);
and U501 (N_501,In_189,In_1852);
or U502 (N_502,In_1437,In_872);
nand U503 (N_503,In_2019,In_2017);
or U504 (N_504,In_2180,In_1891);
xnor U505 (N_505,In_835,In_2471);
nand U506 (N_506,In_1570,In_436);
xnor U507 (N_507,In_2137,In_1974);
xnor U508 (N_508,In_484,In_1839);
and U509 (N_509,In_685,In_261);
nor U510 (N_510,In_886,In_1925);
xnor U511 (N_511,In_1288,In_1433);
nand U512 (N_512,In_445,In_29);
and U513 (N_513,In_1709,In_628);
xor U514 (N_514,In_2325,In_1302);
and U515 (N_515,In_821,In_1655);
and U516 (N_516,In_642,In_1360);
or U517 (N_517,In_1548,In_622);
nand U518 (N_518,In_1738,In_2305);
and U519 (N_519,In_1844,In_1752);
nand U520 (N_520,In_2077,In_574);
nor U521 (N_521,In_930,In_737);
nand U522 (N_522,In_238,In_1365);
nor U523 (N_523,In_2177,In_1173);
or U524 (N_524,In_2145,In_2287);
and U525 (N_525,In_138,In_1645);
or U526 (N_526,In_2414,In_1073);
nand U527 (N_527,In_870,In_2376);
nor U528 (N_528,In_791,In_1875);
or U529 (N_529,In_614,In_1247);
xnor U530 (N_530,In_1277,In_1378);
nand U531 (N_531,In_350,In_1470);
or U532 (N_532,In_437,In_1065);
and U533 (N_533,In_2146,In_1375);
xor U534 (N_534,In_742,In_680);
and U535 (N_535,In_2429,In_1165);
or U536 (N_536,In_918,In_2088);
xnor U537 (N_537,In_1961,In_903);
xnor U538 (N_538,In_475,In_139);
or U539 (N_539,In_817,In_488);
and U540 (N_540,In_333,In_2251);
and U541 (N_541,In_1242,In_215);
and U542 (N_542,In_847,In_760);
xnor U543 (N_543,In_757,In_2294);
and U544 (N_544,In_2072,In_1671);
nand U545 (N_545,In_239,In_2244);
nand U546 (N_546,In_1546,In_2378);
nand U547 (N_547,In_1927,In_920);
or U548 (N_548,In_2252,In_661);
or U549 (N_549,In_1822,In_1832);
nor U550 (N_550,In_1235,In_1571);
or U551 (N_551,In_621,In_1442);
nand U552 (N_552,In_1792,In_443);
and U553 (N_553,In_1669,In_2439);
and U554 (N_554,In_2455,In_313);
or U555 (N_555,In_43,In_157);
and U556 (N_556,In_2155,In_909);
xor U557 (N_557,In_2201,In_2197);
nand U558 (N_558,In_2016,In_2044);
nand U559 (N_559,In_57,In_2447);
nand U560 (N_560,In_1599,In_1385);
xor U561 (N_561,In_787,In_977);
nand U562 (N_562,In_1579,In_1327);
or U563 (N_563,In_1560,In_1299);
xor U564 (N_564,In_570,In_938);
or U565 (N_565,In_1708,In_2418);
and U566 (N_566,In_1880,In_946);
nand U567 (N_567,In_1520,In_2354);
or U568 (N_568,In_1993,In_74);
nor U569 (N_569,In_2262,In_1215);
or U570 (N_570,In_1404,In_135);
nand U571 (N_571,In_1105,In_1628);
nor U572 (N_572,In_830,In_1810);
xnor U573 (N_573,In_727,In_826);
nand U574 (N_574,In_1184,In_2033);
and U575 (N_575,In_1491,In_1465);
xnor U576 (N_576,In_340,In_1502);
nand U577 (N_577,In_607,In_858);
or U578 (N_578,In_174,In_1649);
xnor U579 (N_579,In_458,In_2126);
nand U580 (N_580,In_1568,In_1705);
and U581 (N_581,In_1558,In_1670);
and U582 (N_582,In_1210,In_740);
nor U583 (N_583,In_2121,In_2172);
nor U584 (N_584,In_1871,In_2207);
nor U585 (N_585,In_1687,In_450);
nand U586 (N_586,In_391,In_879);
and U587 (N_587,In_999,In_1506);
and U588 (N_588,In_515,In_440);
xnor U589 (N_589,In_1674,In_761);
xor U590 (N_590,In_435,In_971);
or U591 (N_591,In_355,In_1766);
nand U592 (N_592,In_1275,In_11);
nor U593 (N_593,In_377,In_2435);
and U594 (N_594,In_531,In_116);
nor U595 (N_595,In_1783,In_1312);
or U596 (N_596,In_1837,In_134);
nor U597 (N_597,In_2181,In_588);
nand U598 (N_598,In_186,In_1290);
or U599 (N_599,In_2210,In_841);
or U600 (N_600,In_433,In_97);
xnor U601 (N_601,In_1045,In_2093);
nand U602 (N_602,In_1726,In_90);
nor U603 (N_603,In_953,In_776);
nor U604 (N_604,In_2346,In_453);
nand U605 (N_605,In_753,In_2406);
xnor U606 (N_606,In_266,In_1831);
nor U607 (N_607,In_467,In_1688);
nor U608 (N_608,In_2448,In_779);
xor U609 (N_609,In_1026,In_130);
xnor U610 (N_610,In_2347,In_2263);
nor U611 (N_611,In_1819,In_2235);
and U612 (N_612,In_1176,In_68);
nand U613 (N_613,In_2080,In_1193);
and U614 (N_614,In_832,In_1836);
nor U615 (N_615,In_1031,In_64);
or U616 (N_616,In_1643,In_2426);
nor U617 (N_617,In_1858,In_1902);
xnor U618 (N_618,In_806,In_507);
nand U619 (N_619,In_2139,In_152);
nor U620 (N_620,In_1128,In_2212);
nand U621 (N_621,In_1808,In_1426);
or U622 (N_622,In_387,In_1979);
nor U623 (N_623,In_1333,In_1694);
or U624 (N_624,In_518,In_1339);
nor U625 (N_625,In_2027,In_968);
nor U626 (N_626,In_643,In_2069);
nor U627 (N_627,In_295,In_555);
or U628 (N_628,In_1134,In_257);
and U629 (N_629,In_1140,In_2384);
or U630 (N_630,In_153,In_1056);
nor U631 (N_631,In_327,In_418);
nor U632 (N_632,In_1240,In_378);
nor U633 (N_633,In_2482,In_2012);
and U634 (N_634,In_1614,In_124);
or U635 (N_635,In_624,In_173);
nor U636 (N_636,In_289,In_631);
and U637 (N_637,In_1668,In_1957);
nor U638 (N_638,In_457,In_1039);
xnor U639 (N_639,In_2459,In_2289);
nor U640 (N_640,In_81,In_35);
or U641 (N_641,In_1040,In_752);
nand U642 (N_642,In_987,In_1545);
and U643 (N_643,In_770,In_1998);
nand U644 (N_644,In_801,In_1689);
nor U645 (N_645,In_194,In_196);
and U646 (N_646,In_1507,In_2022);
and U647 (N_647,In_2499,In_1304);
xnor U648 (N_648,In_1931,In_598);
nor U649 (N_649,In_1314,In_1809);
nor U650 (N_650,In_956,In_735);
xor U651 (N_651,In_1924,In_1347);
nor U652 (N_652,In_2049,In_308);
nand U653 (N_653,In_589,In_126);
and U654 (N_654,In_983,In_1870);
nor U655 (N_655,In_1500,In_892);
or U656 (N_656,In_985,In_1338);
nor U657 (N_657,In_10,In_976);
and U658 (N_658,In_2123,In_961);
xnor U659 (N_659,In_539,In_1166);
nor U660 (N_660,In_1594,In_1218);
or U661 (N_661,In_1068,In_1344);
nor U662 (N_662,In_1625,In_917);
nand U663 (N_663,In_664,In_339);
or U664 (N_664,In_1712,In_1876);
nor U665 (N_665,In_1245,In_1728);
and U666 (N_666,In_2318,In_1417);
nand U667 (N_667,In_2420,In_612);
nand U668 (N_668,In_2415,In_2377);
xor U669 (N_669,In_2460,In_2096);
and U670 (N_670,In_2115,In_2029);
or U671 (N_671,In_810,In_224);
xor U672 (N_672,In_1262,In_2290);
xor U673 (N_673,In_846,In_883);
or U674 (N_674,In_1021,In_849);
nor U675 (N_675,In_2281,In_717);
xnor U676 (N_676,In_1474,In_1080);
nor U677 (N_677,In_755,In_2195);
or U678 (N_678,In_957,In_1124);
nand U679 (N_679,In_2310,In_1864);
or U680 (N_680,In_538,In_1873);
xnor U681 (N_681,In_156,In_1895);
and U682 (N_682,In_2131,In_2014);
or U683 (N_683,In_1332,In_1531);
xnor U684 (N_684,In_1308,In_25);
nor U685 (N_685,In_733,In_2059);
xnor U686 (N_686,In_1412,In_1942);
xnor U687 (N_687,In_82,In_1445);
or U688 (N_688,In_2260,In_1850);
nor U689 (N_689,In_2046,In_202);
nand U690 (N_690,In_509,In_2437);
and U691 (N_691,In_42,In_2385);
and U692 (N_692,In_565,In_1846);
nand U693 (N_693,In_2120,In_1714);
or U694 (N_694,In_2320,In_2342);
and U695 (N_695,In_311,In_1196);
nand U696 (N_696,In_373,In_1204);
nor U697 (N_697,In_2284,In_1753);
nor U698 (N_698,In_487,In_2174);
or U699 (N_699,In_2094,In_2358);
and U700 (N_700,In_427,In_1519);
nor U701 (N_701,In_659,In_2428);
nand U702 (N_702,In_514,In_98);
nand U703 (N_703,In_845,In_1572);
nor U704 (N_704,In_1725,In_306);
xor U705 (N_705,In_1269,In_599);
or U706 (N_706,In_2497,In_232);
and U707 (N_707,In_2158,In_1055);
xnor U708 (N_708,In_217,In_1919);
or U709 (N_709,In_69,In_1872);
or U710 (N_710,In_1553,In_309);
nor U711 (N_711,In_2229,In_1791);
nor U712 (N_712,In_119,In_277);
nand U713 (N_713,In_1162,In_1002);
and U714 (N_714,In_1681,In_520);
xnor U715 (N_715,In_991,In_1928);
and U716 (N_716,In_553,In_608);
or U717 (N_717,In_1113,In_136);
and U718 (N_718,In_703,In_751);
and U719 (N_719,In_1070,In_1343);
xnor U720 (N_720,In_2132,In_298);
and U721 (N_721,In_1471,In_1677);
and U722 (N_722,In_1127,In_802);
and U723 (N_723,In_2147,In_1527);
nand U724 (N_724,In_167,In_2394);
or U725 (N_725,In_2104,In_596);
and U726 (N_726,In_290,In_1116);
or U727 (N_727,In_2286,In_1843);
nand U728 (N_728,In_2357,In_2095);
nand U729 (N_729,In_2189,In_1066);
or U730 (N_730,In_1346,In_1642);
nand U731 (N_731,In_2109,In_61);
nor U732 (N_732,In_76,In_434);
nor U733 (N_733,In_1648,In_1222);
nand U734 (N_734,In_972,In_1255);
or U735 (N_735,In_273,In_2443);
nor U736 (N_736,In_2250,In_2185);
and U737 (N_737,In_1556,In_522);
nand U738 (N_738,In_898,In_650);
xor U739 (N_739,In_1881,In_874);
nor U740 (N_740,In_1492,In_1980);
xor U741 (N_741,In_472,In_1746);
nand U742 (N_742,In_67,In_404);
nor U743 (N_743,In_1446,In_1216);
nor U744 (N_744,In_1794,In_855);
and U745 (N_745,In_1644,In_1238);
and U746 (N_746,In_37,In_2091);
and U747 (N_747,In_2240,In_1589);
nand U748 (N_748,In_1847,In_149);
or U749 (N_749,In_118,In_1440);
nand U750 (N_750,In_516,In_1806);
and U751 (N_751,In_560,In_2110);
or U752 (N_752,In_264,In_513);
or U753 (N_753,In_2011,In_2298);
or U754 (N_754,In_88,In_1513);
nand U755 (N_755,In_851,In_2032);
and U756 (N_756,In_2136,In_300);
xor U757 (N_757,In_681,In_1274);
nor U758 (N_758,In_31,In_400);
or U759 (N_759,In_2143,In_1436);
or U760 (N_760,In_283,In_954);
xnor U761 (N_761,In_1401,In_1154);
nor U762 (N_762,In_2315,In_388);
xor U763 (N_763,In_900,In_1003);
xnor U764 (N_764,In_2365,In_1398);
and U765 (N_765,In_974,In_653);
or U766 (N_766,In_1842,In_728);
nand U767 (N_767,In_493,In_2204);
nor U768 (N_768,In_785,In_1435);
nor U769 (N_769,In_2144,In_2015);
and U770 (N_770,In_1194,In_2487);
xor U771 (N_771,In_2444,In_2464);
and U772 (N_772,In_1208,In_2004);
or U773 (N_773,In_2278,In_471);
nor U774 (N_774,In_2434,In_223);
nor U775 (N_775,In_1774,In_940);
nand U776 (N_776,In_1971,In_1120);
nor U777 (N_777,In_1525,In_2198);
xnor U778 (N_778,In_2243,In_1109);
and U779 (N_779,In_2477,In_1915);
or U780 (N_780,In_406,In_594);
and U781 (N_781,In_1664,In_878);
and U782 (N_782,In_2296,In_2193);
nor U783 (N_783,In_155,In_1731);
nor U784 (N_784,In_209,In_713);
and U785 (N_785,In_1467,In_941);
and U786 (N_786,In_571,In_1273);
and U787 (N_787,In_265,In_349);
nor U788 (N_788,In_1425,In_998);
and U789 (N_789,In_1486,In_1874);
nand U790 (N_790,In_1170,In_468);
xor U791 (N_791,In_756,In_330);
nor U792 (N_792,In_1144,In_477);
xor U793 (N_793,In_1898,In_2074);
xnor U794 (N_794,In_2498,In_1771);
or U795 (N_795,In_2293,In_1884);
or U796 (N_796,In_1214,In_269);
or U797 (N_797,In_638,In_1650);
nor U798 (N_798,In_1652,In_981);
and U799 (N_799,In_2379,In_1896);
and U800 (N_800,In_2188,In_2361);
or U801 (N_801,In_412,In_2335);
and U802 (N_802,In_193,In_2410);
xor U803 (N_803,In_716,In_1330);
or U804 (N_804,In_2421,In_2299);
and U805 (N_805,In_1700,In_1522);
nand U806 (N_806,In_1407,In_1250);
and U807 (N_807,In_824,In_366);
nor U808 (N_808,In_1763,In_1724);
nand U809 (N_809,In_583,In_233);
xor U810 (N_810,In_1,In_1729);
nand U811 (N_811,In_2276,In_2247);
xor U812 (N_812,In_646,In_1722);
xnor U813 (N_813,In_997,In_314);
nor U814 (N_814,In_245,In_2391);
and U815 (N_815,In_2404,In_561);
xor U816 (N_816,In_840,In_229);
nand U817 (N_817,In_1693,In_2249);
xnor U818 (N_818,In_1913,In_1533);
nor U819 (N_819,In_613,In_2352);
nor U820 (N_820,In_2138,In_79);
or U821 (N_821,In_2382,In_1157);
nand U822 (N_822,In_1260,In_2370);
nor U823 (N_823,In_684,In_1524);
nor U824 (N_824,In_2030,In_1185);
and U825 (N_825,In_1454,In_1750);
or U826 (N_826,In_464,In_771);
nor U827 (N_827,In_1991,In_2401);
nand U828 (N_828,In_2273,In_536);
or U829 (N_829,In_1569,In_1660);
and U830 (N_830,In_2023,In_401);
xnor U831 (N_831,In_558,In_1815);
nand U832 (N_832,In_2042,In_414);
nor U833 (N_833,In_541,In_1243);
nand U834 (N_834,In_600,In_2113);
xnor U835 (N_835,In_1813,In_1139);
or U836 (N_836,In_1062,In_1239);
or U837 (N_837,In_2387,In_1030);
nor U838 (N_838,In_1727,In_2327);
and U839 (N_839,In_1754,In_2285);
nand U840 (N_840,In_2283,In_317);
nand U841 (N_841,In_402,In_2328);
nand U842 (N_842,In_1230,In_1541);
nor U843 (N_843,In_354,In_2245);
or U844 (N_844,In_161,In_1263);
nand U845 (N_845,In_547,In_496);
nor U846 (N_846,In_1862,In_1391);
xor U847 (N_847,In_1703,In_1715);
or U848 (N_848,In_1937,In_429);
or U849 (N_849,In_382,In_1939);
or U850 (N_850,In_1457,In_1220);
xor U851 (N_851,In_1219,In_212);
nand U852 (N_852,In_582,In_1690);
nor U853 (N_853,In_1713,In_950);
xnor U854 (N_854,In_1485,In_1390);
nand U855 (N_855,In_667,In_489);
and U856 (N_856,In_1640,In_348);
nand U857 (N_857,In_480,In_2452);
xor U858 (N_858,In_2232,In_1122);
nor U859 (N_859,In_328,In_1504);
or U860 (N_860,In_2313,In_663);
nor U861 (N_861,In_210,In_34);
nor U862 (N_862,In_2291,In_2265);
nor U863 (N_863,In_316,In_931);
and U864 (N_864,In_747,In_1297);
xor U865 (N_865,In_1567,In_1439);
nor U866 (N_866,In_304,In_397);
and U867 (N_867,In_101,In_884);
nand U868 (N_868,In_1807,In_1086);
nand U869 (N_869,In_1131,In_27);
nor U870 (N_870,In_1489,In_563);
and U871 (N_871,In_688,In_2163);
and U872 (N_872,In_1638,In_465);
and U873 (N_873,In_356,In_1367);
xor U874 (N_874,In_637,In_768);
and U875 (N_875,In_2496,In_1825);
nand U876 (N_876,In_1917,In_967);
nor U877 (N_877,In_831,In_910);
nor U878 (N_878,In_1472,In_1526);
and U879 (N_879,In_860,In_937);
nor U880 (N_880,In_705,In_1102);
nor U881 (N_881,In_441,In_1863);
xnor U882 (N_882,In_478,In_1618);
or U883 (N_883,In_1138,In_2272);
nor U884 (N_884,In_41,In_28);
nand U885 (N_885,In_1544,In_665);
nand U886 (N_886,In_554,In_928);
or U887 (N_887,In_2332,In_270);
nand U888 (N_888,In_1936,In_2098);
nor U889 (N_889,In_1047,In_112);
nor U890 (N_890,In_1226,In_1598);
and U891 (N_891,In_2408,In_2107);
or U892 (N_892,In_294,In_960);
nand U893 (N_893,In_1296,In_1654);
nor U894 (N_894,In_1494,In_2003);
nand U895 (N_895,In_1285,In_1972);
nor U896 (N_896,In_1493,In_405);
nand U897 (N_897,In_1879,In_369);
and U898 (N_898,In_66,In_696);
xnor U899 (N_899,In_323,In_1776);
or U900 (N_900,In_813,In_335);
nand U901 (N_901,In_1322,In_1866);
xor U902 (N_902,In_147,In_528);
nor U903 (N_903,In_241,In_1697);
or U904 (N_904,In_1376,In_1315);
nand U905 (N_905,In_1736,In_2341);
xnor U906 (N_906,In_1295,In_71);
nor U907 (N_907,In_2364,In_2215);
nor U908 (N_908,In_604,In_490);
nand U909 (N_909,In_1886,In_1409);
or U910 (N_910,In_1342,In_47);
nor U911 (N_911,In_2413,In_1617);
xor U912 (N_912,In_1563,In_893);
and U913 (N_913,In_30,In_1258);
and U914 (N_914,In_2319,In_828);
xnor U915 (N_915,In_188,In_1751);
and U916 (N_916,In_2431,In_1532);
nor U917 (N_917,In_73,In_2006);
nor U918 (N_918,In_2231,In_2190);
nand U919 (N_919,In_2129,In_610);
or U920 (N_920,In_221,In_1765);
nand U921 (N_921,In_322,In_1189);
nor U922 (N_922,In_800,In_1246);
nand U923 (N_923,In_1244,In_325);
and U924 (N_924,In_2288,In_8);
and U925 (N_925,In_121,In_1661);
nand U926 (N_926,In_143,In_2403);
nor U927 (N_927,In_723,In_1371);
nor U928 (N_928,In_1006,In_934);
nor U929 (N_929,In_1720,In_1211);
and U930 (N_930,In_485,In_1782);
nor U931 (N_931,In_745,In_1530);
nor U932 (N_932,In_922,In_1394);
xor U933 (N_933,In_1337,In_1796);
nand U934 (N_934,In_1431,In_111);
and U935 (N_935,In_2353,In_2089);
nand U936 (N_936,In_2334,In_1340);
and U937 (N_937,In_2301,In_945);
nor U938 (N_938,In_2119,In_92);
nor U939 (N_939,In_641,In_1951);
and U940 (N_940,In_1966,In_652);
nand U941 (N_941,In_36,In_398);
and U942 (N_942,In_262,In_276);
nand U943 (N_943,In_1221,In_449);
and U944 (N_944,In_2430,In_601);
or U945 (N_945,In_1704,In_1666);
or U946 (N_946,In_2045,In_164);
and U947 (N_947,In_1908,In_719);
nor U948 (N_948,In_2256,In_871);
nand U949 (N_949,In_2209,In_1349);
and U950 (N_950,In_1178,In_1117);
and U951 (N_951,In_2323,In_2433);
nand U952 (N_952,In_1038,In_1945);
nand U953 (N_953,In_375,In_1897);
xnor U954 (N_954,In_159,In_888);
nor U955 (N_955,In_1691,In_609);
nand U956 (N_956,In_192,In_2337);
nor U957 (N_957,In_1575,In_2224);
nand U958 (N_958,In_842,In_2372);
xnor U959 (N_959,In_1987,In_695);
or U960 (N_960,In_318,In_1883);
and U961 (N_961,In_2495,In_519);
nor U962 (N_962,In_1076,In_1584);
xor U963 (N_963,In_137,In_1464);
nand U964 (N_964,In_1023,In_1309);
xor U965 (N_965,In_409,In_19);
or U966 (N_966,In_1015,In_178);
and U967 (N_967,In_422,In_181);
nand U968 (N_968,In_1386,In_1744);
xnor U969 (N_969,In_1759,In_1388);
nand U970 (N_970,In_1287,In_815);
xnor U971 (N_971,In_0,In_657);
nor U972 (N_972,In_995,In_1657);
and U973 (N_973,In_545,In_1795);
or U974 (N_974,In_171,In_1266);
xor U975 (N_975,In_32,In_2222);
and U976 (N_976,In_1855,In_2196);
and U977 (N_977,In_766,In_970);
xnor U978 (N_978,In_1967,In_420);
or U979 (N_979,In_1610,In_1778);
nor U980 (N_980,In_466,In_1835);
and U981 (N_981,In_91,In_532);
and U982 (N_982,In_505,In_428);
nand U983 (N_983,In_916,In_1946);
or U984 (N_984,In_1590,In_1680);
nand U985 (N_985,In_45,In_292);
nand U986 (N_986,In_619,In_2474);
nand U987 (N_987,In_1498,In_1619);
xnor U988 (N_988,In_1790,In_2491);
nand U989 (N_989,In_880,In_1382);
xor U990 (N_990,In_1585,In_278);
nor U991 (N_991,In_383,In_1374);
and U992 (N_992,In_230,In_1413);
xnor U993 (N_993,In_2153,In_2392);
and U994 (N_994,In_1192,In_2438);
xnor U995 (N_995,In_568,In_87);
or U996 (N_996,In_1577,In_1217);
nor U997 (N_997,In_2386,In_820);
nor U998 (N_998,In_1119,In_2127);
nand U999 (N_999,In_2068,In_1817);
nand U1000 (N_1000,In_1932,In_399);
xnor U1001 (N_1001,In_113,In_1914);
and U1002 (N_1002,In_586,In_1800);
or U1003 (N_1003,In_1986,In_512);
or U1004 (N_1004,In_347,In_675);
or U1005 (N_1005,In_1651,In_1201);
xor U1006 (N_1006,In_1615,In_1292);
nor U1007 (N_1007,In_862,In_630);
or U1008 (N_1008,In_501,In_634);
and U1009 (N_1009,In_2130,In_1887);
xnor U1010 (N_1010,In_906,In_17);
and U1011 (N_1011,In_2246,In_1552);
nor U1012 (N_1012,In_702,In_1133);
or U1013 (N_1013,In_782,In_1373);
nor U1014 (N_1014,In_710,In_915);
nand U1015 (N_1015,In_1631,In_1014);
nor U1016 (N_1016,In_616,In_744);
xnor U1017 (N_1017,In_899,In_1641);
or U1018 (N_1018,In_962,In_825);
nand U1019 (N_1019,In_1025,In_1072);
xnor U1020 (N_1020,In_2230,In_1828);
nand U1021 (N_1021,In_1495,In_60);
or U1022 (N_1022,In_1602,In_123);
xnor U1023 (N_1023,In_591,In_1463);
nor U1024 (N_1024,In_158,In_207);
or U1025 (N_1025,In_1331,In_148);
or U1026 (N_1026,In_1482,In_2058);
and U1027 (N_1027,In_1501,In_1605);
xnor U1028 (N_1028,In_2211,In_694);
xor U1029 (N_1029,In_2417,In_280);
and U1030 (N_1030,In_984,In_617);
or U1031 (N_1031,In_662,In_2461);
and U1032 (N_1032,In_1780,In_1174);
nor U1033 (N_1033,In_359,In_933);
nand U1034 (N_1034,In_1155,In_12);
xor U1035 (N_1035,In_549,In_1079);
xor U1036 (N_1036,In_2,In_894);
nor U1037 (N_1037,In_1368,In_777);
or U1038 (N_1038,In_367,In_2395);
or U1039 (N_1039,In_1143,In_1834);
nand U1040 (N_1040,In_473,In_1345);
nor U1041 (N_1041,In_1089,In_623);
nand U1042 (N_1042,In_2076,In_861);
and U1043 (N_1043,In_758,In_1637);
or U1044 (N_1044,In_762,In_2206);
xnor U1045 (N_1045,In_2453,In_1310);
and U1046 (N_1046,In_1202,In_2407);
or U1047 (N_1047,In_408,In_297);
and U1048 (N_1048,In_1696,In_848);
or U1049 (N_1049,In_1743,In_2261);
nor U1050 (N_1050,In_272,In_1959);
nor U1051 (N_1051,In_1764,In_1291);
xnor U1052 (N_1052,In_722,In_1994);
nor U1053 (N_1053,In_534,In_1484);
and U1054 (N_1054,In_1542,In_2152);
nand U1055 (N_1055,In_1402,In_1608);
nand U1056 (N_1056,In_1833,In_1364);
nand U1057 (N_1057,In_1935,In_1099);
xnor U1058 (N_1058,In_1361,In_2488);
or U1059 (N_1059,In_386,In_343);
xnor U1060 (N_1060,In_48,In_948);
xnor U1061 (N_1061,In_792,In_2297);
and U1062 (N_1062,In_926,In_1316);
and U1063 (N_1063,In_2071,In_2274);
nand U1064 (N_1064,In_1613,In_2486);
or U1065 (N_1065,In_1228,In_1311);
and U1066 (N_1066,In_1930,In_1195);
and U1067 (N_1067,In_151,In_1947);
nor U1068 (N_1068,In_2321,In_2134);
and U1069 (N_1069,In_243,In_730);
nor U1070 (N_1070,In_2481,In_220);
xnor U1071 (N_1071,In_1294,In_1268);
and U1072 (N_1072,In_635,In_1326);
nor U1073 (N_1073,In_2475,In_955);
nand U1074 (N_1074,In_1926,In_2028);
or U1075 (N_1075,In_2065,In_1267);
nor U1076 (N_1076,In_370,In_2103);
and U1077 (N_1077,In_1997,In_2043);
xor U1078 (N_1078,In_1324,In_2053);
nand U1079 (N_1079,In_216,In_921);
nor U1080 (N_1080,In_1306,In_2035);
xnor U1081 (N_1081,In_1027,In_154);
nand U1082 (N_1082,In_2267,In_654);
and U1083 (N_1083,In_2349,In_686);
nand U1084 (N_1084,In_1591,In_620);
nand U1085 (N_1085,In_2419,In_1051);
and U1086 (N_1086,In_526,In_365);
nand U1087 (N_1087,In_818,In_226);
nor U1088 (N_1088,In_1554,In_1955);
and U1089 (N_1089,In_781,In_213);
nand U1090 (N_1090,In_1392,In_379);
and U1091 (N_1091,In_1452,In_1962);
nand U1092 (N_1092,In_497,In_1621);
nor U1093 (N_1093,In_572,In_980);
and U1094 (N_1094,In_794,In_1001);
nand U1095 (N_1095,In_1037,In_837);
or U1096 (N_1096,In_797,In_1811);
nand U1097 (N_1097,In_255,In_535);
xor U1098 (N_1098,In_439,In_75);
nand U1099 (N_1099,In_1814,In_247);
xor U1100 (N_1100,In_1547,In_765);
and U1101 (N_1101,In_146,In_2140);
and U1102 (N_1102,In_714,In_2031);
and U1103 (N_1103,In_2086,In_564);
and U1104 (N_1104,In_165,In_1153);
and U1105 (N_1105,In_1335,In_1058);
and U1106 (N_1106,In_315,In_644);
xor U1107 (N_1107,In_175,In_246);
nor U1108 (N_1108,In_1695,In_1679);
or U1109 (N_1109,In_1272,In_1334);
nor U1110 (N_1110,In_55,In_593);
nand U1111 (N_1111,In_1505,In_1397);
and U1112 (N_1112,In_1395,In_805);
or U1113 (N_1113,In_511,In_1551);
nand U1114 (N_1114,In_361,In_595);
nand U1115 (N_1115,In_1233,In_575);
nor U1116 (N_1116,In_1707,In_179);
and U1117 (N_1117,In_78,In_1205);
and U1118 (N_1118,In_1181,In_1148);
xor U1119 (N_1119,In_767,In_2326);
or U1120 (N_1120,In_1787,In_764);
or U1121 (N_1121,In_1550,In_924);
nor U1122 (N_1122,In_959,In_2336);
nand U1123 (N_1123,In_1595,In_763);
nand U1124 (N_1124,In_344,In_668);
and U1125 (N_1125,In_1175,In_1142);
nand U1126 (N_1126,In_556,In_1403);
xor U1127 (N_1127,In_2489,In_1091);
xor U1128 (N_1128,In_1107,In_836);
xnor U1129 (N_1129,In_908,In_360);
nor U1130 (N_1130,In_1849,In_24);
nor U1131 (N_1131,In_550,In_1622);
nand U1132 (N_1132,In_2225,In_769);
nand U1133 (N_1133,In_2186,In_2432);
and U1134 (N_1134,In_1716,In_2451);
nand U1135 (N_1135,In_2067,In_460);
and U1136 (N_1136,In_1092,In_1733);
xnor U1137 (N_1137,In_231,In_1934);
and U1138 (N_1138,In_606,In_925);
xnor U1139 (N_1139,In_2200,In_1958);
or U1140 (N_1140,In_163,In_1867);
and U1141 (N_1141,In_1826,In_1321);
and U1142 (N_1142,In_1480,In_687);
xnor U1143 (N_1143,In_2402,In_1033);
nand U1144 (N_1144,In_2396,In_911);
and U1145 (N_1145,In_2307,In_1528);
or U1146 (N_1146,In_1101,In_1761);
and U1147 (N_1147,In_2214,In_52);
or U1148 (N_1148,In_1964,In_109);
and U1149 (N_1149,In_709,In_1878);
nor U1150 (N_1150,In_1779,In_707);
nand U1151 (N_1151,In_271,In_2340);
xnor U1152 (N_1152,In_102,In_302);
or U1153 (N_1153,In_1430,In_197);
nor U1154 (N_1154,In_205,In_1818);
nor U1155 (N_1155,In_1053,In_2054);
nand U1156 (N_1156,In_1389,In_1539);
and U1157 (N_1157,In_2409,In_199);
xnor U1158 (N_1158,In_1905,In_2202);
nor U1159 (N_1159,In_1387,In_1973);
nor U1160 (N_1160,In_611,In_1422);
or U1161 (N_1161,In_1497,In_1561);
or U1162 (N_1162,In_989,In_1059);
nand U1163 (N_1163,In_1802,In_672);
nand U1164 (N_1164,In_882,In_706);
and U1165 (N_1165,In_1061,In_2097);
xor U1166 (N_1166,In_198,In_844);
or U1167 (N_1167,In_1992,In_2388);
xnor U1168 (N_1168,In_1593,In_578);
nor U1169 (N_1169,In_1424,In_1923);
or U1170 (N_1170,In_376,In_494);
or U1171 (N_1171,In_1469,In_2275);
xnor U1172 (N_1172,In_1854,In_1231);
nand U1173 (N_1173,In_2466,In_403);
nand U1174 (N_1174,In_1559,In_1786);
nand U1175 (N_1175,In_973,In_1965);
and U1176 (N_1176,In_736,In_2162);
or U1177 (N_1177,In_856,In_1789);
nand U1178 (N_1178,In_145,In_1933);
xnor U1179 (N_1179,In_237,In_1904);
and U1180 (N_1180,In_14,In_1305);
nand U1181 (N_1181,In_1358,In_772);
nor U1182 (N_1182,In_2330,In_1151);
nor U1183 (N_1183,In_699,In_1894);
nand U1184 (N_1184,In_2375,In_1949);
or U1185 (N_1185,In_1685,In_1603);
nand U1186 (N_1186,In_456,In_1909);
nand U1187 (N_1187,In_992,In_1199);
and U1188 (N_1188,In_698,In_656);
and U1189 (N_1189,In_577,In_2351);
or U1190 (N_1190,In_1067,In_1741);
nor U1191 (N_1191,In_1410,In_1583);
nand U1192 (N_1192,In_1509,In_2149);
or U1193 (N_1193,In_1289,In_2184);
nor U1194 (N_1194,In_1126,In_2425);
nor U1195 (N_1195,In_2002,In_1702);
or U1196 (N_1196,In_248,In_1626);
or U1197 (N_1197,In_222,In_20);
nand U1198 (N_1198,In_1254,In_1044);
xor U1199 (N_1199,In_2199,In_267);
xnor U1200 (N_1200,In_2479,In_2020);
nor U1201 (N_1201,In_1760,In_310);
nor U1202 (N_1202,In_2078,In_2060);
and U1203 (N_1203,In_2465,In_666);
nand U1204 (N_1204,In_2075,In_1428);
nand U1205 (N_1205,In_537,In_869);
xnor U1206 (N_1206,In_1742,In_919);
and U1207 (N_1207,In_180,In_748);
xnor U1208 (N_1208,In_1013,In_2010);
nor U1209 (N_1209,In_1252,In_1414);
and U1210 (N_1210,In_58,In_618);
xor U1211 (N_1211,In_603,In_1048);
and U1212 (N_1212,In_2338,In_2309);
nor U1213 (N_1213,In_1675,In_1455);
and U1214 (N_1214,In_301,In_183);
xor U1215 (N_1215,In_2171,In_859);
nand U1216 (N_1216,In_2371,In_228);
nor U1217 (N_1217,In_2374,In_444);
nand U1218 (N_1218,In_446,In_7);
xor U1219 (N_1219,In_1699,In_567);
nand U1220 (N_1220,In_214,In_626);
nor U1221 (N_1221,In_655,In_476);
xor U1222 (N_1222,In_1630,In_2363);
nand U1223 (N_1223,In_182,In_1574);
nand U1224 (N_1224,In_1627,In_2277);
nand U1225 (N_1225,In_2025,In_1207);
and U1226 (N_1226,In_1757,In_218);
or U1227 (N_1227,In_708,In_1663);
or U1228 (N_1228,In_2445,In_701);
and U1229 (N_1229,In_2142,In_1123);
xor U1230 (N_1230,In_1557,In_1823);
or U1231 (N_1231,In_829,In_1995);
nand U1232 (N_1232,In_1448,In_1803);
nor U1233 (N_1233,In_1159,In_1456);
nand U1234 (N_1234,In_951,In_778);
nand U1235 (N_1235,In_1587,In_833);
xnor U1236 (N_1236,In_396,In_1369);
nor U1237 (N_1237,In_943,In_168);
and U1238 (N_1238,In_1421,In_853);
xor U1239 (N_1239,In_2040,In_1921);
nor U1240 (N_1240,In_120,In_2062);
nand U1241 (N_1241,In_838,In_529);
and U1242 (N_1242,In_416,In_1400);
or U1243 (N_1243,In_1950,In_1461);
and U1244 (N_1244,In_2151,In_1784);
nand U1245 (N_1245,In_1186,In_2329);
or U1246 (N_1246,In_1348,In_1607);
xor U1247 (N_1247,In_5,In_1662);
or U1248 (N_1248,In_1948,In_2221);
nand U1249 (N_1249,In_211,In_1381);
nor U1250 (N_1250,In_2016,In_1803);
nor U1251 (N_1251,In_773,In_1802);
xnor U1252 (N_1252,In_1247,In_1663);
nor U1253 (N_1253,In_2050,In_1563);
nor U1254 (N_1254,In_1611,In_988);
xnor U1255 (N_1255,In_398,In_2480);
nand U1256 (N_1256,In_1947,In_1597);
nand U1257 (N_1257,In_1117,In_261);
nand U1258 (N_1258,In_1005,In_540);
xor U1259 (N_1259,In_1042,In_921);
or U1260 (N_1260,In_1386,In_1481);
xor U1261 (N_1261,In_1458,In_2243);
nor U1262 (N_1262,In_1119,In_1115);
xnor U1263 (N_1263,In_828,In_2286);
and U1264 (N_1264,In_1433,In_1568);
nor U1265 (N_1265,In_2199,In_1620);
nand U1266 (N_1266,In_2073,In_780);
nor U1267 (N_1267,In_291,In_1616);
or U1268 (N_1268,In_2197,In_1989);
xor U1269 (N_1269,In_1281,In_349);
nand U1270 (N_1270,In_235,In_1984);
xor U1271 (N_1271,In_172,In_892);
nand U1272 (N_1272,In_1930,In_2495);
or U1273 (N_1273,In_1773,In_311);
nand U1274 (N_1274,In_926,In_2437);
and U1275 (N_1275,In_1363,In_610);
nand U1276 (N_1276,In_660,In_2400);
and U1277 (N_1277,In_1414,In_2260);
nand U1278 (N_1278,In_806,In_1685);
nand U1279 (N_1279,In_72,In_2334);
or U1280 (N_1280,In_23,In_1644);
xor U1281 (N_1281,In_1060,In_1658);
xor U1282 (N_1282,In_1160,In_1772);
or U1283 (N_1283,In_663,In_1043);
and U1284 (N_1284,In_2238,In_2153);
and U1285 (N_1285,In_1401,In_106);
nor U1286 (N_1286,In_72,In_1157);
and U1287 (N_1287,In_2037,In_2455);
xnor U1288 (N_1288,In_845,In_2207);
and U1289 (N_1289,In_1932,In_1645);
and U1290 (N_1290,In_2224,In_1555);
xnor U1291 (N_1291,In_2094,In_1095);
or U1292 (N_1292,In_2196,In_1988);
and U1293 (N_1293,In_2398,In_503);
or U1294 (N_1294,In_728,In_205);
nor U1295 (N_1295,In_98,In_258);
xnor U1296 (N_1296,In_2038,In_993);
nand U1297 (N_1297,In_681,In_737);
nand U1298 (N_1298,In_1662,In_2445);
and U1299 (N_1299,In_852,In_823);
xnor U1300 (N_1300,In_1052,In_2456);
nor U1301 (N_1301,In_19,In_1246);
xnor U1302 (N_1302,In_1544,In_1321);
nand U1303 (N_1303,In_1707,In_971);
or U1304 (N_1304,In_975,In_2320);
or U1305 (N_1305,In_496,In_1533);
nor U1306 (N_1306,In_1292,In_2060);
nand U1307 (N_1307,In_52,In_2415);
or U1308 (N_1308,In_2294,In_1989);
and U1309 (N_1309,In_959,In_2076);
nand U1310 (N_1310,In_1312,In_1966);
or U1311 (N_1311,In_2413,In_1155);
and U1312 (N_1312,In_1685,In_1557);
and U1313 (N_1313,In_1262,In_120);
nand U1314 (N_1314,In_1342,In_901);
nor U1315 (N_1315,In_1061,In_1091);
xor U1316 (N_1316,In_1044,In_1268);
xnor U1317 (N_1317,In_34,In_1837);
and U1318 (N_1318,In_1365,In_1754);
or U1319 (N_1319,In_1954,In_721);
xnor U1320 (N_1320,In_2160,In_2107);
xnor U1321 (N_1321,In_1323,In_534);
and U1322 (N_1322,In_1540,In_1078);
xor U1323 (N_1323,In_1071,In_2241);
xor U1324 (N_1324,In_1836,In_353);
nand U1325 (N_1325,In_2200,In_121);
xor U1326 (N_1326,In_589,In_677);
nor U1327 (N_1327,In_1380,In_1544);
nor U1328 (N_1328,In_1632,In_1343);
nand U1329 (N_1329,In_313,In_455);
nand U1330 (N_1330,In_757,In_740);
xnor U1331 (N_1331,In_135,In_867);
and U1332 (N_1332,In_267,In_2010);
xnor U1333 (N_1333,In_537,In_1740);
and U1334 (N_1334,In_2318,In_1931);
nor U1335 (N_1335,In_318,In_209);
nand U1336 (N_1336,In_217,In_1960);
nor U1337 (N_1337,In_1005,In_1380);
xor U1338 (N_1338,In_810,In_808);
or U1339 (N_1339,In_1100,In_1451);
xnor U1340 (N_1340,In_1503,In_2285);
or U1341 (N_1341,In_626,In_2215);
nor U1342 (N_1342,In_2440,In_2377);
xnor U1343 (N_1343,In_993,In_327);
or U1344 (N_1344,In_137,In_165);
or U1345 (N_1345,In_1642,In_1714);
and U1346 (N_1346,In_404,In_1197);
and U1347 (N_1347,In_1755,In_520);
or U1348 (N_1348,In_711,In_1043);
and U1349 (N_1349,In_879,In_2343);
or U1350 (N_1350,In_2215,In_417);
nand U1351 (N_1351,In_2417,In_345);
xnor U1352 (N_1352,In_1270,In_1415);
xnor U1353 (N_1353,In_984,In_669);
or U1354 (N_1354,In_488,In_885);
or U1355 (N_1355,In_2348,In_403);
nor U1356 (N_1356,In_677,In_2408);
nand U1357 (N_1357,In_1245,In_513);
and U1358 (N_1358,In_1158,In_359);
nor U1359 (N_1359,In_1513,In_1889);
xor U1360 (N_1360,In_1470,In_1427);
and U1361 (N_1361,In_1601,In_154);
xor U1362 (N_1362,In_1815,In_1167);
nor U1363 (N_1363,In_1224,In_2163);
xor U1364 (N_1364,In_836,In_1490);
xnor U1365 (N_1365,In_2159,In_1293);
nand U1366 (N_1366,In_1428,In_765);
and U1367 (N_1367,In_1080,In_718);
or U1368 (N_1368,In_1767,In_2312);
xor U1369 (N_1369,In_397,In_1987);
nand U1370 (N_1370,In_156,In_2186);
or U1371 (N_1371,In_1959,In_1017);
xnor U1372 (N_1372,In_1488,In_828);
nor U1373 (N_1373,In_1096,In_1248);
nand U1374 (N_1374,In_1345,In_1574);
xnor U1375 (N_1375,In_2202,In_758);
xnor U1376 (N_1376,In_1726,In_954);
xor U1377 (N_1377,In_423,In_2263);
nor U1378 (N_1378,In_622,In_2384);
xor U1379 (N_1379,In_635,In_1778);
nor U1380 (N_1380,In_123,In_673);
nor U1381 (N_1381,In_2302,In_749);
or U1382 (N_1382,In_972,In_1935);
nor U1383 (N_1383,In_1074,In_941);
or U1384 (N_1384,In_62,In_1886);
and U1385 (N_1385,In_759,In_409);
xnor U1386 (N_1386,In_2078,In_294);
and U1387 (N_1387,In_2355,In_559);
nand U1388 (N_1388,In_905,In_1842);
xnor U1389 (N_1389,In_1772,In_1150);
xor U1390 (N_1390,In_1549,In_658);
nand U1391 (N_1391,In_1013,In_891);
nand U1392 (N_1392,In_1714,In_2071);
and U1393 (N_1393,In_1394,In_1922);
nor U1394 (N_1394,In_1375,In_1438);
or U1395 (N_1395,In_1323,In_157);
and U1396 (N_1396,In_1900,In_1270);
or U1397 (N_1397,In_1895,In_2100);
nand U1398 (N_1398,In_60,In_1031);
and U1399 (N_1399,In_2009,In_2042);
or U1400 (N_1400,In_1664,In_2081);
xnor U1401 (N_1401,In_200,In_1430);
and U1402 (N_1402,In_2470,In_506);
xor U1403 (N_1403,In_11,In_1317);
nand U1404 (N_1404,In_1856,In_586);
or U1405 (N_1405,In_293,In_257);
nand U1406 (N_1406,In_597,In_21);
nor U1407 (N_1407,In_2420,In_1399);
and U1408 (N_1408,In_1094,In_1659);
nor U1409 (N_1409,In_1693,In_1655);
or U1410 (N_1410,In_1028,In_227);
nand U1411 (N_1411,In_0,In_1645);
nor U1412 (N_1412,In_164,In_589);
or U1413 (N_1413,In_1093,In_2025);
and U1414 (N_1414,In_1239,In_808);
xor U1415 (N_1415,In_1275,In_1344);
and U1416 (N_1416,In_503,In_167);
nand U1417 (N_1417,In_2138,In_1739);
xor U1418 (N_1418,In_2257,In_1603);
or U1419 (N_1419,In_1688,In_1355);
nand U1420 (N_1420,In_2268,In_1449);
and U1421 (N_1421,In_1372,In_768);
nand U1422 (N_1422,In_831,In_363);
nor U1423 (N_1423,In_1099,In_984);
and U1424 (N_1424,In_1677,In_1278);
and U1425 (N_1425,In_2190,In_643);
nand U1426 (N_1426,In_1444,In_1723);
and U1427 (N_1427,In_2193,In_892);
xor U1428 (N_1428,In_1743,In_767);
and U1429 (N_1429,In_708,In_924);
xnor U1430 (N_1430,In_9,In_1002);
or U1431 (N_1431,In_115,In_1727);
nor U1432 (N_1432,In_2021,In_1489);
and U1433 (N_1433,In_1764,In_1854);
or U1434 (N_1434,In_2377,In_631);
and U1435 (N_1435,In_2330,In_22);
nand U1436 (N_1436,In_1756,In_910);
and U1437 (N_1437,In_2199,In_293);
or U1438 (N_1438,In_1786,In_770);
and U1439 (N_1439,In_577,In_1705);
xor U1440 (N_1440,In_240,In_139);
and U1441 (N_1441,In_2010,In_938);
or U1442 (N_1442,In_961,In_931);
or U1443 (N_1443,In_592,In_2439);
xor U1444 (N_1444,In_824,In_1346);
or U1445 (N_1445,In_278,In_211);
and U1446 (N_1446,In_463,In_1947);
xor U1447 (N_1447,In_1726,In_230);
and U1448 (N_1448,In_691,In_924);
nor U1449 (N_1449,In_1774,In_826);
nor U1450 (N_1450,In_1269,In_38);
nand U1451 (N_1451,In_1876,In_332);
nand U1452 (N_1452,In_125,In_1509);
nand U1453 (N_1453,In_2003,In_1267);
and U1454 (N_1454,In_1205,In_626);
or U1455 (N_1455,In_1530,In_1064);
nand U1456 (N_1456,In_2252,In_2281);
nor U1457 (N_1457,In_453,In_2403);
or U1458 (N_1458,In_720,In_877);
nor U1459 (N_1459,In_408,In_1254);
nand U1460 (N_1460,In_161,In_1445);
xor U1461 (N_1461,In_2147,In_91);
and U1462 (N_1462,In_1864,In_927);
nor U1463 (N_1463,In_2260,In_2290);
nor U1464 (N_1464,In_44,In_388);
and U1465 (N_1465,In_111,In_808);
nor U1466 (N_1466,In_2458,In_1010);
and U1467 (N_1467,In_517,In_2155);
or U1468 (N_1468,In_486,In_512);
nor U1469 (N_1469,In_1169,In_480);
nor U1470 (N_1470,In_246,In_1261);
and U1471 (N_1471,In_1359,In_1693);
xor U1472 (N_1472,In_2468,In_232);
or U1473 (N_1473,In_1137,In_1227);
nand U1474 (N_1474,In_1138,In_1895);
and U1475 (N_1475,In_935,In_1192);
or U1476 (N_1476,In_2311,In_761);
or U1477 (N_1477,In_311,In_2192);
nor U1478 (N_1478,In_430,In_719);
xnor U1479 (N_1479,In_1504,In_796);
and U1480 (N_1480,In_2065,In_2309);
nand U1481 (N_1481,In_2403,In_1965);
nand U1482 (N_1482,In_2230,In_1216);
xor U1483 (N_1483,In_683,In_717);
or U1484 (N_1484,In_621,In_1991);
or U1485 (N_1485,In_539,In_1951);
or U1486 (N_1486,In_2315,In_714);
nand U1487 (N_1487,In_2071,In_2264);
or U1488 (N_1488,In_1375,In_72);
or U1489 (N_1489,In_1715,In_138);
nand U1490 (N_1490,In_2141,In_2131);
nor U1491 (N_1491,In_563,In_1445);
and U1492 (N_1492,In_2064,In_2413);
and U1493 (N_1493,In_1588,In_175);
or U1494 (N_1494,In_1598,In_741);
nor U1495 (N_1495,In_1010,In_365);
nor U1496 (N_1496,In_1606,In_623);
nor U1497 (N_1497,In_745,In_1454);
xnor U1498 (N_1498,In_1816,In_946);
nand U1499 (N_1499,In_1258,In_1279);
xor U1500 (N_1500,In_1823,In_1959);
and U1501 (N_1501,In_1343,In_1671);
or U1502 (N_1502,In_48,In_1141);
nor U1503 (N_1503,In_452,In_643);
and U1504 (N_1504,In_489,In_915);
nor U1505 (N_1505,In_42,In_1627);
and U1506 (N_1506,In_1963,In_1523);
nand U1507 (N_1507,In_378,In_945);
and U1508 (N_1508,In_2245,In_1622);
xor U1509 (N_1509,In_101,In_159);
and U1510 (N_1510,In_1760,In_297);
or U1511 (N_1511,In_591,In_2246);
or U1512 (N_1512,In_816,In_1757);
xor U1513 (N_1513,In_1051,In_1663);
nor U1514 (N_1514,In_805,In_806);
nor U1515 (N_1515,In_1873,In_2132);
nand U1516 (N_1516,In_1942,In_1554);
nor U1517 (N_1517,In_347,In_2302);
xor U1518 (N_1518,In_1466,In_1625);
and U1519 (N_1519,In_1801,In_1061);
nor U1520 (N_1520,In_962,In_704);
and U1521 (N_1521,In_2351,In_1787);
and U1522 (N_1522,In_66,In_1431);
or U1523 (N_1523,In_1954,In_1584);
xnor U1524 (N_1524,In_1511,In_937);
nor U1525 (N_1525,In_146,In_1602);
nor U1526 (N_1526,In_1200,In_1624);
nor U1527 (N_1527,In_552,In_393);
or U1528 (N_1528,In_1275,In_1351);
and U1529 (N_1529,In_1503,In_1568);
and U1530 (N_1530,In_914,In_2382);
xor U1531 (N_1531,In_2187,In_1557);
or U1532 (N_1532,In_883,In_2114);
and U1533 (N_1533,In_872,In_1063);
nand U1534 (N_1534,In_264,In_807);
and U1535 (N_1535,In_2133,In_1421);
nor U1536 (N_1536,In_1967,In_167);
or U1537 (N_1537,In_2027,In_139);
nand U1538 (N_1538,In_47,In_199);
xor U1539 (N_1539,In_985,In_1264);
or U1540 (N_1540,In_1246,In_2059);
or U1541 (N_1541,In_454,In_179);
nor U1542 (N_1542,In_755,In_2220);
or U1543 (N_1543,In_150,In_1539);
and U1544 (N_1544,In_1527,In_1768);
and U1545 (N_1545,In_281,In_798);
xnor U1546 (N_1546,In_990,In_1686);
or U1547 (N_1547,In_1110,In_1217);
nor U1548 (N_1548,In_1755,In_1314);
or U1549 (N_1549,In_1964,In_977);
and U1550 (N_1550,In_2278,In_1728);
or U1551 (N_1551,In_500,In_1650);
nor U1552 (N_1552,In_1679,In_362);
and U1553 (N_1553,In_2106,In_2360);
and U1554 (N_1554,In_1095,In_157);
nand U1555 (N_1555,In_1284,In_1884);
nor U1556 (N_1556,In_475,In_1218);
nand U1557 (N_1557,In_2068,In_1227);
nand U1558 (N_1558,In_971,In_1115);
nor U1559 (N_1559,In_1374,In_2006);
xor U1560 (N_1560,In_1428,In_1254);
nor U1561 (N_1561,In_2297,In_1182);
and U1562 (N_1562,In_2406,In_389);
xor U1563 (N_1563,In_990,In_1042);
and U1564 (N_1564,In_1070,In_1372);
nand U1565 (N_1565,In_381,In_999);
nand U1566 (N_1566,In_1623,In_2381);
xor U1567 (N_1567,In_72,In_2274);
or U1568 (N_1568,In_420,In_2282);
nor U1569 (N_1569,In_1444,In_1186);
or U1570 (N_1570,In_1149,In_1707);
nor U1571 (N_1571,In_389,In_369);
or U1572 (N_1572,In_9,In_2323);
nor U1573 (N_1573,In_2340,In_58);
xor U1574 (N_1574,In_1263,In_2108);
and U1575 (N_1575,In_2143,In_1334);
nand U1576 (N_1576,In_1652,In_1821);
and U1577 (N_1577,In_927,In_2481);
nor U1578 (N_1578,In_1352,In_15);
xor U1579 (N_1579,In_2300,In_1031);
or U1580 (N_1580,In_335,In_2190);
and U1581 (N_1581,In_882,In_1702);
nand U1582 (N_1582,In_186,In_2117);
and U1583 (N_1583,In_88,In_2346);
and U1584 (N_1584,In_1890,In_1699);
or U1585 (N_1585,In_2338,In_2259);
xnor U1586 (N_1586,In_721,In_2350);
nor U1587 (N_1587,In_2200,In_569);
nor U1588 (N_1588,In_800,In_665);
or U1589 (N_1589,In_1649,In_375);
and U1590 (N_1590,In_257,In_1524);
xor U1591 (N_1591,In_62,In_2079);
and U1592 (N_1592,In_1153,In_276);
nor U1593 (N_1593,In_686,In_1449);
nand U1594 (N_1594,In_748,In_1820);
and U1595 (N_1595,In_2178,In_677);
or U1596 (N_1596,In_2466,In_2294);
nor U1597 (N_1597,In_1781,In_540);
or U1598 (N_1598,In_984,In_326);
xor U1599 (N_1599,In_54,In_2236);
nand U1600 (N_1600,In_2081,In_657);
and U1601 (N_1601,In_93,In_2370);
xor U1602 (N_1602,In_2475,In_1413);
nor U1603 (N_1603,In_587,In_1082);
xnor U1604 (N_1604,In_2296,In_1444);
nor U1605 (N_1605,In_314,In_351);
xor U1606 (N_1606,In_613,In_1980);
or U1607 (N_1607,In_2151,In_795);
or U1608 (N_1608,In_1592,In_1124);
nand U1609 (N_1609,In_288,In_436);
nor U1610 (N_1610,In_1251,In_2436);
nor U1611 (N_1611,In_1096,In_482);
and U1612 (N_1612,In_591,In_182);
nor U1613 (N_1613,In_1757,In_1591);
nand U1614 (N_1614,In_1019,In_1290);
or U1615 (N_1615,In_1718,In_1383);
nand U1616 (N_1616,In_785,In_2285);
xor U1617 (N_1617,In_2403,In_1356);
and U1618 (N_1618,In_1898,In_397);
xnor U1619 (N_1619,In_43,In_115);
xnor U1620 (N_1620,In_792,In_1801);
and U1621 (N_1621,In_1271,In_1198);
nand U1622 (N_1622,In_825,In_1228);
xor U1623 (N_1623,In_579,In_614);
nor U1624 (N_1624,In_1748,In_1919);
and U1625 (N_1625,In_943,In_942);
nand U1626 (N_1626,In_816,In_409);
nand U1627 (N_1627,In_956,In_733);
xnor U1628 (N_1628,In_1682,In_1554);
and U1629 (N_1629,In_1332,In_1945);
and U1630 (N_1630,In_1167,In_877);
xor U1631 (N_1631,In_119,In_19);
or U1632 (N_1632,In_1798,In_99);
nand U1633 (N_1633,In_344,In_1704);
and U1634 (N_1634,In_2146,In_1965);
nor U1635 (N_1635,In_1904,In_1312);
or U1636 (N_1636,In_119,In_1175);
nor U1637 (N_1637,In_736,In_964);
or U1638 (N_1638,In_2197,In_1651);
xor U1639 (N_1639,In_862,In_524);
nor U1640 (N_1640,In_2123,In_2481);
and U1641 (N_1641,In_1260,In_1584);
and U1642 (N_1642,In_1174,In_2229);
xor U1643 (N_1643,In_1840,In_1091);
and U1644 (N_1644,In_827,In_1167);
xnor U1645 (N_1645,In_395,In_2354);
or U1646 (N_1646,In_546,In_1005);
nor U1647 (N_1647,In_471,In_2480);
or U1648 (N_1648,In_1260,In_1044);
nor U1649 (N_1649,In_1076,In_1175);
xor U1650 (N_1650,In_2138,In_1503);
nor U1651 (N_1651,In_651,In_973);
and U1652 (N_1652,In_881,In_1384);
or U1653 (N_1653,In_775,In_94);
nand U1654 (N_1654,In_1698,In_1704);
nand U1655 (N_1655,In_1683,In_634);
nand U1656 (N_1656,In_1603,In_1208);
nand U1657 (N_1657,In_1333,In_795);
and U1658 (N_1658,In_315,In_1296);
nand U1659 (N_1659,In_609,In_754);
nand U1660 (N_1660,In_2130,In_2285);
xor U1661 (N_1661,In_1641,In_797);
or U1662 (N_1662,In_1970,In_707);
xor U1663 (N_1663,In_1974,In_498);
or U1664 (N_1664,In_201,In_720);
nand U1665 (N_1665,In_335,In_439);
nor U1666 (N_1666,In_835,In_2465);
nand U1667 (N_1667,In_2141,In_2463);
and U1668 (N_1668,In_2266,In_538);
or U1669 (N_1669,In_2011,In_997);
xnor U1670 (N_1670,In_1718,In_842);
nand U1671 (N_1671,In_1173,In_1102);
xnor U1672 (N_1672,In_2083,In_64);
or U1673 (N_1673,In_1970,In_449);
nand U1674 (N_1674,In_1437,In_220);
and U1675 (N_1675,In_2435,In_656);
xnor U1676 (N_1676,In_723,In_300);
xor U1677 (N_1677,In_662,In_582);
nand U1678 (N_1678,In_1213,In_1792);
nor U1679 (N_1679,In_50,In_488);
xor U1680 (N_1680,In_560,In_358);
or U1681 (N_1681,In_259,In_1874);
or U1682 (N_1682,In_362,In_932);
xor U1683 (N_1683,In_897,In_1222);
nand U1684 (N_1684,In_1819,In_1250);
and U1685 (N_1685,In_148,In_1549);
or U1686 (N_1686,In_2295,In_1816);
and U1687 (N_1687,In_1304,In_1038);
and U1688 (N_1688,In_505,In_1631);
or U1689 (N_1689,In_791,In_75);
nand U1690 (N_1690,In_1314,In_2288);
nand U1691 (N_1691,In_933,In_608);
or U1692 (N_1692,In_850,In_2455);
nor U1693 (N_1693,In_1371,In_1123);
nand U1694 (N_1694,In_361,In_967);
xor U1695 (N_1695,In_2493,In_2319);
nor U1696 (N_1696,In_826,In_2184);
nor U1697 (N_1697,In_984,In_1813);
or U1698 (N_1698,In_1918,In_382);
and U1699 (N_1699,In_2308,In_701);
nand U1700 (N_1700,In_1196,In_542);
xnor U1701 (N_1701,In_629,In_2117);
nand U1702 (N_1702,In_449,In_2000);
nand U1703 (N_1703,In_646,In_1448);
and U1704 (N_1704,In_1359,In_1570);
nor U1705 (N_1705,In_200,In_757);
xnor U1706 (N_1706,In_1193,In_2014);
nand U1707 (N_1707,In_1618,In_1512);
nor U1708 (N_1708,In_1925,In_1887);
xnor U1709 (N_1709,In_2369,In_305);
and U1710 (N_1710,In_2073,In_879);
or U1711 (N_1711,In_2085,In_1352);
or U1712 (N_1712,In_8,In_1624);
nand U1713 (N_1713,In_253,In_1354);
xor U1714 (N_1714,In_744,In_1152);
xnor U1715 (N_1715,In_1770,In_1710);
or U1716 (N_1716,In_1994,In_2268);
nor U1717 (N_1717,In_401,In_2317);
nand U1718 (N_1718,In_2359,In_1678);
and U1719 (N_1719,In_887,In_1029);
and U1720 (N_1720,In_1444,In_212);
or U1721 (N_1721,In_940,In_1838);
and U1722 (N_1722,In_1885,In_667);
nand U1723 (N_1723,In_304,In_763);
xnor U1724 (N_1724,In_889,In_1608);
or U1725 (N_1725,In_1679,In_291);
and U1726 (N_1726,In_1145,In_2107);
nor U1727 (N_1727,In_1975,In_1679);
nor U1728 (N_1728,In_1114,In_34);
xor U1729 (N_1729,In_243,In_252);
or U1730 (N_1730,In_1374,In_1700);
or U1731 (N_1731,In_1565,In_1396);
nand U1732 (N_1732,In_711,In_605);
nor U1733 (N_1733,In_1085,In_673);
nor U1734 (N_1734,In_1453,In_1329);
or U1735 (N_1735,In_182,In_1697);
xnor U1736 (N_1736,In_2404,In_2486);
nor U1737 (N_1737,In_370,In_906);
nand U1738 (N_1738,In_659,In_2001);
nand U1739 (N_1739,In_2262,In_464);
and U1740 (N_1740,In_2158,In_1634);
or U1741 (N_1741,In_2275,In_2075);
xor U1742 (N_1742,In_1010,In_1212);
nand U1743 (N_1743,In_1774,In_706);
and U1744 (N_1744,In_1715,In_1023);
or U1745 (N_1745,In_1733,In_2106);
and U1746 (N_1746,In_220,In_1375);
and U1747 (N_1747,In_573,In_2172);
and U1748 (N_1748,In_552,In_734);
nor U1749 (N_1749,In_775,In_1448);
nor U1750 (N_1750,In_379,In_458);
or U1751 (N_1751,In_2385,In_1304);
and U1752 (N_1752,In_296,In_546);
or U1753 (N_1753,In_792,In_1748);
and U1754 (N_1754,In_1332,In_1706);
or U1755 (N_1755,In_1550,In_1989);
and U1756 (N_1756,In_2024,In_1671);
nand U1757 (N_1757,In_857,In_2001);
or U1758 (N_1758,In_1710,In_1032);
or U1759 (N_1759,In_2149,In_1137);
or U1760 (N_1760,In_2253,In_321);
nand U1761 (N_1761,In_591,In_483);
nor U1762 (N_1762,In_447,In_500);
xnor U1763 (N_1763,In_851,In_1198);
and U1764 (N_1764,In_2177,In_569);
nand U1765 (N_1765,In_1271,In_1487);
xor U1766 (N_1766,In_1917,In_1350);
xor U1767 (N_1767,In_513,In_1182);
and U1768 (N_1768,In_1342,In_1647);
and U1769 (N_1769,In_2403,In_2199);
nand U1770 (N_1770,In_905,In_894);
xnor U1771 (N_1771,In_2325,In_1174);
nand U1772 (N_1772,In_308,In_1849);
nor U1773 (N_1773,In_1087,In_1656);
nand U1774 (N_1774,In_706,In_1668);
nand U1775 (N_1775,In_1851,In_1343);
xor U1776 (N_1776,In_393,In_755);
nor U1777 (N_1777,In_429,In_860);
xnor U1778 (N_1778,In_1978,In_52);
nand U1779 (N_1779,In_2440,In_856);
nor U1780 (N_1780,In_1338,In_2440);
or U1781 (N_1781,In_266,In_534);
xor U1782 (N_1782,In_962,In_1685);
nand U1783 (N_1783,In_180,In_625);
or U1784 (N_1784,In_2400,In_1759);
xor U1785 (N_1785,In_2381,In_1199);
or U1786 (N_1786,In_2065,In_1002);
nand U1787 (N_1787,In_1658,In_164);
or U1788 (N_1788,In_61,In_51);
or U1789 (N_1789,In_2294,In_1143);
nand U1790 (N_1790,In_849,In_1591);
or U1791 (N_1791,In_997,In_1644);
and U1792 (N_1792,In_479,In_2190);
nor U1793 (N_1793,In_55,In_977);
xnor U1794 (N_1794,In_1505,In_1386);
and U1795 (N_1795,In_211,In_1960);
nand U1796 (N_1796,In_577,In_567);
nor U1797 (N_1797,In_2035,In_642);
nor U1798 (N_1798,In_29,In_2460);
nand U1799 (N_1799,In_1188,In_2375);
or U1800 (N_1800,In_1276,In_950);
and U1801 (N_1801,In_2057,In_1224);
xor U1802 (N_1802,In_2428,In_1144);
and U1803 (N_1803,In_385,In_377);
nor U1804 (N_1804,In_403,In_2260);
nor U1805 (N_1805,In_453,In_817);
or U1806 (N_1806,In_873,In_132);
or U1807 (N_1807,In_1461,In_586);
xnor U1808 (N_1808,In_1658,In_252);
and U1809 (N_1809,In_593,In_382);
xnor U1810 (N_1810,In_1238,In_964);
nand U1811 (N_1811,In_61,In_239);
or U1812 (N_1812,In_2259,In_2061);
nor U1813 (N_1813,In_1798,In_2278);
and U1814 (N_1814,In_1309,In_1526);
nand U1815 (N_1815,In_1238,In_719);
nand U1816 (N_1816,In_2267,In_2017);
nor U1817 (N_1817,In_2456,In_1460);
nor U1818 (N_1818,In_502,In_1366);
nand U1819 (N_1819,In_2127,In_2313);
or U1820 (N_1820,In_741,In_1306);
or U1821 (N_1821,In_2343,In_1026);
nand U1822 (N_1822,In_11,In_2483);
and U1823 (N_1823,In_2299,In_388);
nor U1824 (N_1824,In_201,In_673);
and U1825 (N_1825,In_1782,In_452);
xnor U1826 (N_1826,In_1575,In_483);
or U1827 (N_1827,In_359,In_1225);
nor U1828 (N_1828,In_1237,In_200);
xnor U1829 (N_1829,In_1572,In_976);
and U1830 (N_1830,In_379,In_1818);
nor U1831 (N_1831,In_2306,In_1697);
xnor U1832 (N_1832,In_1742,In_222);
xnor U1833 (N_1833,In_1098,In_756);
and U1834 (N_1834,In_983,In_260);
nand U1835 (N_1835,In_511,In_1146);
nand U1836 (N_1836,In_308,In_887);
xor U1837 (N_1837,In_699,In_2401);
and U1838 (N_1838,In_193,In_166);
and U1839 (N_1839,In_816,In_2155);
nand U1840 (N_1840,In_2164,In_1785);
xor U1841 (N_1841,In_714,In_1527);
or U1842 (N_1842,In_1166,In_2102);
nor U1843 (N_1843,In_1452,In_1670);
and U1844 (N_1844,In_485,In_488);
or U1845 (N_1845,In_628,In_658);
nand U1846 (N_1846,In_1074,In_824);
nor U1847 (N_1847,In_645,In_1237);
xor U1848 (N_1848,In_835,In_450);
nor U1849 (N_1849,In_21,In_1475);
or U1850 (N_1850,In_2107,In_1237);
or U1851 (N_1851,In_227,In_1808);
nand U1852 (N_1852,In_889,In_1696);
or U1853 (N_1853,In_2107,In_1919);
xnor U1854 (N_1854,In_1725,In_419);
nor U1855 (N_1855,In_1790,In_2186);
and U1856 (N_1856,In_848,In_1907);
or U1857 (N_1857,In_1915,In_1354);
nand U1858 (N_1858,In_1905,In_1900);
and U1859 (N_1859,In_1843,In_1513);
nand U1860 (N_1860,In_2389,In_2492);
and U1861 (N_1861,In_2193,In_2323);
nand U1862 (N_1862,In_2258,In_552);
xnor U1863 (N_1863,In_413,In_1029);
xnor U1864 (N_1864,In_2180,In_442);
xnor U1865 (N_1865,In_1516,In_1083);
nand U1866 (N_1866,In_376,In_1181);
nand U1867 (N_1867,In_2327,In_2402);
or U1868 (N_1868,In_295,In_548);
nor U1869 (N_1869,In_2354,In_836);
or U1870 (N_1870,In_1693,In_2369);
nor U1871 (N_1871,In_2261,In_1061);
nor U1872 (N_1872,In_914,In_1100);
nor U1873 (N_1873,In_1456,In_1573);
nor U1874 (N_1874,In_1,In_282);
nand U1875 (N_1875,In_1864,In_235);
nor U1876 (N_1876,In_1808,In_962);
xnor U1877 (N_1877,In_2357,In_41);
and U1878 (N_1878,In_1441,In_1359);
nand U1879 (N_1879,In_2258,In_757);
nor U1880 (N_1880,In_310,In_228);
xor U1881 (N_1881,In_65,In_1790);
xnor U1882 (N_1882,In_1699,In_1658);
nand U1883 (N_1883,In_1419,In_920);
nand U1884 (N_1884,In_398,In_2218);
or U1885 (N_1885,In_2268,In_1155);
nand U1886 (N_1886,In_1798,In_812);
nand U1887 (N_1887,In_1367,In_1175);
or U1888 (N_1888,In_664,In_1097);
and U1889 (N_1889,In_785,In_2142);
nand U1890 (N_1890,In_582,In_871);
or U1891 (N_1891,In_1946,In_559);
and U1892 (N_1892,In_1805,In_392);
nand U1893 (N_1893,In_1230,In_1705);
and U1894 (N_1894,In_1856,In_2396);
nand U1895 (N_1895,In_2485,In_1240);
or U1896 (N_1896,In_1424,In_108);
nand U1897 (N_1897,In_727,In_866);
or U1898 (N_1898,In_97,In_800);
nand U1899 (N_1899,In_572,In_1608);
and U1900 (N_1900,In_921,In_710);
xor U1901 (N_1901,In_59,In_332);
xnor U1902 (N_1902,In_2271,In_1950);
and U1903 (N_1903,In_956,In_917);
or U1904 (N_1904,In_556,In_262);
nor U1905 (N_1905,In_1352,In_826);
xor U1906 (N_1906,In_1871,In_2277);
nand U1907 (N_1907,In_72,In_448);
or U1908 (N_1908,In_2476,In_1127);
nor U1909 (N_1909,In_2288,In_838);
or U1910 (N_1910,In_7,In_766);
nand U1911 (N_1911,In_1946,In_2366);
nor U1912 (N_1912,In_218,In_1152);
and U1913 (N_1913,In_1175,In_535);
nand U1914 (N_1914,In_2003,In_2442);
xnor U1915 (N_1915,In_2468,In_559);
xor U1916 (N_1916,In_217,In_1068);
and U1917 (N_1917,In_741,In_1171);
xnor U1918 (N_1918,In_123,In_32);
and U1919 (N_1919,In_163,In_2349);
xnor U1920 (N_1920,In_319,In_2004);
nand U1921 (N_1921,In_2321,In_1678);
or U1922 (N_1922,In_100,In_2197);
nand U1923 (N_1923,In_749,In_1279);
and U1924 (N_1924,In_870,In_1602);
nand U1925 (N_1925,In_143,In_1085);
xnor U1926 (N_1926,In_679,In_195);
nor U1927 (N_1927,In_597,In_2456);
nor U1928 (N_1928,In_49,In_1351);
nor U1929 (N_1929,In_1140,In_1190);
and U1930 (N_1930,In_1307,In_2234);
and U1931 (N_1931,In_193,In_8);
and U1932 (N_1932,In_902,In_1367);
and U1933 (N_1933,In_1675,In_859);
xnor U1934 (N_1934,In_2389,In_2103);
nand U1935 (N_1935,In_1966,In_306);
nor U1936 (N_1936,In_1717,In_1544);
xnor U1937 (N_1937,In_2283,In_1331);
xor U1938 (N_1938,In_2108,In_2228);
or U1939 (N_1939,In_980,In_282);
or U1940 (N_1940,In_2461,In_414);
and U1941 (N_1941,In_617,In_35);
or U1942 (N_1942,In_1917,In_1885);
nand U1943 (N_1943,In_2489,In_197);
and U1944 (N_1944,In_1090,In_118);
or U1945 (N_1945,In_1942,In_1250);
or U1946 (N_1946,In_230,In_1015);
xnor U1947 (N_1947,In_1286,In_2172);
or U1948 (N_1948,In_158,In_2388);
nand U1949 (N_1949,In_1350,In_50);
nand U1950 (N_1950,In_2325,In_888);
nand U1951 (N_1951,In_793,In_410);
or U1952 (N_1952,In_456,In_1962);
nand U1953 (N_1953,In_2335,In_2298);
nand U1954 (N_1954,In_1155,In_377);
nand U1955 (N_1955,In_124,In_1490);
nand U1956 (N_1956,In_702,In_2467);
and U1957 (N_1957,In_1017,In_792);
nand U1958 (N_1958,In_766,In_765);
and U1959 (N_1959,In_983,In_2278);
xnor U1960 (N_1960,In_1583,In_2121);
xnor U1961 (N_1961,In_218,In_2296);
nor U1962 (N_1962,In_2414,In_1520);
nor U1963 (N_1963,In_2112,In_2495);
nand U1964 (N_1964,In_2084,In_1401);
xnor U1965 (N_1965,In_1106,In_463);
or U1966 (N_1966,In_398,In_2447);
nor U1967 (N_1967,In_2141,In_869);
and U1968 (N_1968,In_740,In_1890);
xor U1969 (N_1969,In_314,In_1154);
xnor U1970 (N_1970,In_1213,In_1100);
or U1971 (N_1971,In_1780,In_1751);
xor U1972 (N_1972,In_819,In_2310);
nor U1973 (N_1973,In_1195,In_2002);
or U1974 (N_1974,In_2195,In_864);
xnor U1975 (N_1975,In_2326,In_72);
or U1976 (N_1976,In_1508,In_253);
or U1977 (N_1977,In_2105,In_981);
or U1978 (N_1978,In_1211,In_2169);
nand U1979 (N_1979,In_759,In_1742);
nor U1980 (N_1980,In_2357,In_876);
nand U1981 (N_1981,In_1097,In_1546);
xnor U1982 (N_1982,In_1623,In_2019);
or U1983 (N_1983,In_2213,In_1978);
nand U1984 (N_1984,In_1959,In_368);
and U1985 (N_1985,In_2301,In_982);
nand U1986 (N_1986,In_216,In_200);
nand U1987 (N_1987,In_97,In_664);
nor U1988 (N_1988,In_1665,In_1060);
xor U1989 (N_1989,In_2003,In_1226);
xnor U1990 (N_1990,In_1339,In_163);
nor U1991 (N_1991,In_1541,In_1812);
and U1992 (N_1992,In_2139,In_192);
nand U1993 (N_1993,In_1318,In_742);
xor U1994 (N_1994,In_1139,In_371);
nor U1995 (N_1995,In_356,In_530);
and U1996 (N_1996,In_2283,In_2224);
xnor U1997 (N_1997,In_1850,In_303);
nand U1998 (N_1998,In_2143,In_471);
nor U1999 (N_1999,In_2279,In_324);
or U2000 (N_2000,In_691,In_259);
or U2001 (N_2001,In_2227,In_2039);
nand U2002 (N_2002,In_163,In_439);
xnor U2003 (N_2003,In_2452,In_1564);
xor U2004 (N_2004,In_1473,In_1103);
or U2005 (N_2005,In_290,In_1802);
nor U2006 (N_2006,In_812,In_999);
xor U2007 (N_2007,In_346,In_2301);
xor U2008 (N_2008,In_635,In_1158);
nor U2009 (N_2009,In_2361,In_574);
and U2010 (N_2010,In_1255,In_896);
or U2011 (N_2011,In_2078,In_11);
nor U2012 (N_2012,In_508,In_316);
nand U2013 (N_2013,In_869,In_327);
xnor U2014 (N_2014,In_993,In_2451);
xor U2015 (N_2015,In_713,In_721);
xor U2016 (N_2016,In_1898,In_326);
nor U2017 (N_2017,In_1068,In_1375);
or U2018 (N_2018,In_325,In_2103);
or U2019 (N_2019,In_2412,In_1367);
and U2020 (N_2020,In_401,In_354);
nand U2021 (N_2021,In_1593,In_1893);
or U2022 (N_2022,In_37,In_1814);
nand U2023 (N_2023,In_507,In_1588);
nand U2024 (N_2024,In_1014,In_1975);
nor U2025 (N_2025,In_2059,In_1760);
and U2026 (N_2026,In_524,In_271);
and U2027 (N_2027,In_1301,In_1851);
nor U2028 (N_2028,In_2053,In_980);
nor U2029 (N_2029,In_1215,In_2298);
or U2030 (N_2030,In_2242,In_1368);
nand U2031 (N_2031,In_897,In_2291);
or U2032 (N_2032,In_1598,In_738);
nor U2033 (N_2033,In_1968,In_1459);
nor U2034 (N_2034,In_1770,In_2175);
nand U2035 (N_2035,In_930,In_625);
or U2036 (N_2036,In_921,In_809);
or U2037 (N_2037,In_1162,In_1603);
or U2038 (N_2038,In_1238,In_858);
and U2039 (N_2039,In_241,In_93);
nor U2040 (N_2040,In_1744,In_1549);
nand U2041 (N_2041,In_2126,In_1261);
nand U2042 (N_2042,In_1366,In_2304);
nand U2043 (N_2043,In_1194,In_2371);
nand U2044 (N_2044,In_417,In_811);
or U2045 (N_2045,In_1163,In_1434);
nor U2046 (N_2046,In_1271,In_36);
nand U2047 (N_2047,In_1431,In_383);
nor U2048 (N_2048,In_2480,In_1249);
nand U2049 (N_2049,In_1350,In_359);
or U2050 (N_2050,In_871,In_246);
nand U2051 (N_2051,In_2182,In_1873);
xor U2052 (N_2052,In_1631,In_2395);
or U2053 (N_2053,In_560,In_302);
and U2054 (N_2054,In_2350,In_822);
nand U2055 (N_2055,In_1982,In_1655);
nor U2056 (N_2056,In_858,In_1011);
nor U2057 (N_2057,In_1756,In_1605);
and U2058 (N_2058,In_1482,In_1193);
nor U2059 (N_2059,In_1884,In_225);
and U2060 (N_2060,In_972,In_639);
xnor U2061 (N_2061,In_1866,In_185);
and U2062 (N_2062,In_1657,In_1211);
nand U2063 (N_2063,In_779,In_81);
nor U2064 (N_2064,In_122,In_51);
nor U2065 (N_2065,In_2480,In_238);
and U2066 (N_2066,In_2084,In_2398);
nor U2067 (N_2067,In_2171,In_999);
nor U2068 (N_2068,In_1988,In_457);
nor U2069 (N_2069,In_1160,In_75);
nor U2070 (N_2070,In_113,In_476);
nor U2071 (N_2071,In_1290,In_307);
xnor U2072 (N_2072,In_892,In_1313);
nor U2073 (N_2073,In_1475,In_1068);
nand U2074 (N_2074,In_1789,In_2384);
nand U2075 (N_2075,In_2,In_1385);
nor U2076 (N_2076,In_259,In_311);
xnor U2077 (N_2077,In_990,In_1001);
xor U2078 (N_2078,In_43,In_756);
nand U2079 (N_2079,In_544,In_808);
nor U2080 (N_2080,In_1973,In_198);
or U2081 (N_2081,In_231,In_2133);
and U2082 (N_2082,In_644,In_1889);
nor U2083 (N_2083,In_2098,In_731);
or U2084 (N_2084,In_2394,In_224);
nor U2085 (N_2085,In_672,In_1375);
and U2086 (N_2086,In_1352,In_496);
xor U2087 (N_2087,In_174,In_2249);
and U2088 (N_2088,In_1484,In_1669);
or U2089 (N_2089,In_180,In_1683);
nor U2090 (N_2090,In_1109,In_1557);
xnor U2091 (N_2091,In_515,In_12);
nor U2092 (N_2092,In_343,In_10);
and U2093 (N_2093,In_2402,In_952);
nand U2094 (N_2094,In_1267,In_83);
and U2095 (N_2095,In_2133,In_667);
xor U2096 (N_2096,In_1278,In_111);
nor U2097 (N_2097,In_657,In_1324);
xnor U2098 (N_2098,In_1104,In_619);
or U2099 (N_2099,In_1522,In_90);
or U2100 (N_2100,In_1152,In_129);
nand U2101 (N_2101,In_1514,In_2394);
or U2102 (N_2102,In_1452,In_2459);
xor U2103 (N_2103,In_203,In_1268);
and U2104 (N_2104,In_637,In_211);
nand U2105 (N_2105,In_1166,In_2428);
xnor U2106 (N_2106,In_66,In_1053);
nand U2107 (N_2107,In_1403,In_1668);
nor U2108 (N_2108,In_479,In_493);
and U2109 (N_2109,In_464,In_221);
or U2110 (N_2110,In_1746,In_2339);
or U2111 (N_2111,In_2150,In_529);
nand U2112 (N_2112,In_1890,In_1616);
or U2113 (N_2113,In_1255,In_1781);
nor U2114 (N_2114,In_1203,In_2128);
nand U2115 (N_2115,In_1679,In_915);
xnor U2116 (N_2116,In_517,In_43);
nand U2117 (N_2117,In_1392,In_440);
nand U2118 (N_2118,In_1961,In_682);
nor U2119 (N_2119,In_283,In_1190);
nand U2120 (N_2120,In_1135,In_180);
or U2121 (N_2121,In_2214,In_978);
and U2122 (N_2122,In_2392,In_374);
nor U2123 (N_2123,In_1926,In_250);
or U2124 (N_2124,In_1245,In_1904);
nor U2125 (N_2125,In_471,In_2132);
nor U2126 (N_2126,In_1166,In_921);
xor U2127 (N_2127,In_512,In_1592);
or U2128 (N_2128,In_1971,In_563);
nor U2129 (N_2129,In_510,In_745);
nand U2130 (N_2130,In_478,In_322);
nand U2131 (N_2131,In_170,In_1780);
or U2132 (N_2132,In_963,In_1053);
and U2133 (N_2133,In_656,In_614);
xor U2134 (N_2134,In_1526,In_86);
xnor U2135 (N_2135,In_1919,In_2250);
and U2136 (N_2136,In_1804,In_1281);
nand U2137 (N_2137,In_374,In_276);
or U2138 (N_2138,In_667,In_456);
or U2139 (N_2139,In_1861,In_2220);
xor U2140 (N_2140,In_763,In_255);
nor U2141 (N_2141,In_410,In_2024);
xnor U2142 (N_2142,In_561,In_934);
nor U2143 (N_2143,In_1792,In_1484);
nand U2144 (N_2144,In_664,In_1806);
and U2145 (N_2145,In_985,In_206);
nor U2146 (N_2146,In_1315,In_1174);
or U2147 (N_2147,In_643,In_341);
or U2148 (N_2148,In_327,In_441);
xor U2149 (N_2149,In_1122,In_721);
xnor U2150 (N_2150,In_2001,In_43);
or U2151 (N_2151,In_1902,In_202);
xor U2152 (N_2152,In_1417,In_2220);
xor U2153 (N_2153,In_2219,In_1166);
nand U2154 (N_2154,In_776,In_1883);
or U2155 (N_2155,In_170,In_2121);
nand U2156 (N_2156,In_2124,In_877);
nand U2157 (N_2157,In_122,In_2003);
or U2158 (N_2158,In_1364,In_165);
nand U2159 (N_2159,In_520,In_335);
and U2160 (N_2160,In_379,In_1959);
and U2161 (N_2161,In_910,In_948);
nand U2162 (N_2162,In_725,In_636);
xnor U2163 (N_2163,In_43,In_677);
xor U2164 (N_2164,In_2183,In_2158);
nand U2165 (N_2165,In_1551,In_355);
nor U2166 (N_2166,In_1152,In_977);
xnor U2167 (N_2167,In_1813,In_1177);
nor U2168 (N_2168,In_2040,In_1);
xnor U2169 (N_2169,In_18,In_1922);
nor U2170 (N_2170,In_1316,In_1896);
nor U2171 (N_2171,In_22,In_2093);
nand U2172 (N_2172,In_1290,In_11);
xor U2173 (N_2173,In_2211,In_187);
nor U2174 (N_2174,In_501,In_2428);
or U2175 (N_2175,In_91,In_1708);
nand U2176 (N_2176,In_766,In_2337);
nor U2177 (N_2177,In_853,In_2384);
or U2178 (N_2178,In_1044,In_2204);
xor U2179 (N_2179,In_1254,In_1457);
nand U2180 (N_2180,In_2049,In_208);
nor U2181 (N_2181,In_301,In_1613);
nor U2182 (N_2182,In_825,In_1930);
and U2183 (N_2183,In_2197,In_1393);
xnor U2184 (N_2184,In_1306,In_773);
or U2185 (N_2185,In_970,In_670);
nor U2186 (N_2186,In_413,In_21);
or U2187 (N_2187,In_1542,In_1554);
nor U2188 (N_2188,In_1034,In_1278);
nand U2189 (N_2189,In_776,In_1531);
xor U2190 (N_2190,In_526,In_1918);
nor U2191 (N_2191,In_1477,In_211);
nor U2192 (N_2192,In_776,In_402);
and U2193 (N_2193,In_1098,In_1255);
or U2194 (N_2194,In_222,In_1129);
and U2195 (N_2195,In_533,In_164);
nor U2196 (N_2196,In_2005,In_1555);
xnor U2197 (N_2197,In_773,In_1435);
or U2198 (N_2198,In_987,In_1770);
xnor U2199 (N_2199,In_795,In_2375);
nor U2200 (N_2200,In_149,In_2385);
xor U2201 (N_2201,In_16,In_96);
or U2202 (N_2202,In_1932,In_2430);
nor U2203 (N_2203,In_1242,In_682);
or U2204 (N_2204,In_595,In_1604);
nand U2205 (N_2205,In_1297,In_1182);
xor U2206 (N_2206,In_1111,In_490);
nor U2207 (N_2207,In_130,In_1637);
xnor U2208 (N_2208,In_697,In_2266);
or U2209 (N_2209,In_80,In_450);
and U2210 (N_2210,In_2449,In_403);
or U2211 (N_2211,In_1626,In_1426);
or U2212 (N_2212,In_1634,In_658);
or U2213 (N_2213,In_1525,In_2239);
nor U2214 (N_2214,In_1721,In_299);
and U2215 (N_2215,In_2401,In_2222);
or U2216 (N_2216,In_266,In_1103);
nand U2217 (N_2217,In_662,In_1384);
nor U2218 (N_2218,In_2458,In_104);
nand U2219 (N_2219,In_677,In_679);
or U2220 (N_2220,In_1690,In_2099);
xnor U2221 (N_2221,In_1635,In_1468);
xor U2222 (N_2222,In_251,In_127);
or U2223 (N_2223,In_45,In_1552);
nor U2224 (N_2224,In_534,In_1128);
xnor U2225 (N_2225,In_732,In_1979);
nand U2226 (N_2226,In_1190,In_2171);
and U2227 (N_2227,In_1302,In_1312);
or U2228 (N_2228,In_509,In_1895);
nand U2229 (N_2229,In_988,In_814);
nand U2230 (N_2230,In_2335,In_1649);
or U2231 (N_2231,In_114,In_2009);
nand U2232 (N_2232,In_2236,In_307);
nor U2233 (N_2233,In_1958,In_1936);
and U2234 (N_2234,In_1434,In_1334);
xnor U2235 (N_2235,In_649,In_1910);
nand U2236 (N_2236,In_296,In_2006);
or U2237 (N_2237,In_440,In_1901);
or U2238 (N_2238,In_1741,In_809);
or U2239 (N_2239,In_2270,In_572);
nor U2240 (N_2240,In_760,In_1569);
or U2241 (N_2241,In_1024,In_859);
and U2242 (N_2242,In_918,In_922);
or U2243 (N_2243,In_1704,In_206);
and U2244 (N_2244,In_1968,In_2260);
or U2245 (N_2245,In_2084,In_1450);
xor U2246 (N_2246,In_2045,In_1088);
or U2247 (N_2247,In_1155,In_759);
and U2248 (N_2248,In_829,In_1987);
xor U2249 (N_2249,In_1415,In_617);
xor U2250 (N_2250,In_2150,In_1782);
or U2251 (N_2251,In_1616,In_1847);
nor U2252 (N_2252,In_624,In_1047);
nand U2253 (N_2253,In_1717,In_1204);
nand U2254 (N_2254,In_1329,In_1887);
nor U2255 (N_2255,In_1640,In_1130);
nor U2256 (N_2256,In_1106,In_1667);
and U2257 (N_2257,In_3,In_1142);
xor U2258 (N_2258,In_1167,In_1010);
nand U2259 (N_2259,In_1366,In_880);
nor U2260 (N_2260,In_1415,In_2117);
nor U2261 (N_2261,In_907,In_2031);
and U2262 (N_2262,In_1543,In_987);
nand U2263 (N_2263,In_721,In_2083);
xor U2264 (N_2264,In_2158,In_1179);
or U2265 (N_2265,In_246,In_627);
nand U2266 (N_2266,In_380,In_1958);
nand U2267 (N_2267,In_1788,In_596);
and U2268 (N_2268,In_682,In_162);
nor U2269 (N_2269,In_1603,In_1015);
xnor U2270 (N_2270,In_1958,In_1521);
xor U2271 (N_2271,In_1496,In_965);
nor U2272 (N_2272,In_1859,In_155);
nand U2273 (N_2273,In_820,In_2322);
and U2274 (N_2274,In_1057,In_362);
nor U2275 (N_2275,In_1372,In_968);
xor U2276 (N_2276,In_1590,In_29);
nor U2277 (N_2277,In_414,In_1840);
nand U2278 (N_2278,In_1468,In_2264);
nor U2279 (N_2279,In_1939,In_2073);
or U2280 (N_2280,In_415,In_817);
nand U2281 (N_2281,In_358,In_1382);
and U2282 (N_2282,In_558,In_1449);
and U2283 (N_2283,In_412,In_1332);
and U2284 (N_2284,In_2447,In_1785);
nor U2285 (N_2285,In_79,In_193);
and U2286 (N_2286,In_321,In_2304);
nor U2287 (N_2287,In_871,In_719);
xnor U2288 (N_2288,In_651,In_1980);
or U2289 (N_2289,In_587,In_1994);
or U2290 (N_2290,In_969,In_27);
nor U2291 (N_2291,In_248,In_1881);
and U2292 (N_2292,In_2183,In_394);
and U2293 (N_2293,In_1832,In_296);
nor U2294 (N_2294,In_489,In_2216);
nand U2295 (N_2295,In_1821,In_483);
and U2296 (N_2296,In_960,In_1547);
xnor U2297 (N_2297,In_819,In_826);
and U2298 (N_2298,In_13,In_2256);
or U2299 (N_2299,In_2380,In_1604);
xnor U2300 (N_2300,In_2364,In_1644);
nand U2301 (N_2301,In_903,In_927);
or U2302 (N_2302,In_464,In_796);
and U2303 (N_2303,In_1084,In_23);
xnor U2304 (N_2304,In_987,In_227);
xnor U2305 (N_2305,In_788,In_1848);
nor U2306 (N_2306,In_362,In_1724);
or U2307 (N_2307,In_520,In_2455);
and U2308 (N_2308,In_1696,In_1450);
xnor U2309 (N_2309,In_2467,In_1354);
nand U2310 (N_2310,In_321,In_2479);
nor U2311 (N_2311,In_618,In_1835);
and U2312 (N_2312,In_1063,In_271);
or U2313 (N_2313,In_2090,In_2094);
nand U2314 (N_2314,In_1911,In_252);
nand U2315 (N_2315,In_2416,In_1022);
nand U2316 (N_2316,In_887,In_2241);
or U2317 (N_2317,In_2131,In_1474);
nor U2318 (N_2318,In_617,In_2116);
nand U2319 (N_2319,In_437,In_212);
or U2320 (N_2320,In_762,In_1380);
xor U2321 (N_2321,In_465,In_872);
nand U2322 (N_2322,In_179,In_259);
xor U2323 (N_2323,In_2233,In_1764);
nor U2324 (N_2324,In_911,In_1012);
and U2325 (N_2325,In_917,In_1059);
or U2326 (N_2326,In_1523,In_1863);
xnor U2327 (N_2327,In_2024,In_2364);
xor U2328 (N_2328,In_1826,In_1381);
and U2329 (N_2329,In_1007,In_1060);
xor U2330 (N_2330,In_736,In_69);
or U2331 (N_2331,In_1620,In_840);
or U2332 (N_2332,In_1982,In_34);
or U2333 (N_2333,In_1245,In_146);
or U2334 (N_2334,In_2422,In_101);
nand U2335 (N_2335,In_1576,In_1130);
xor U2336 (N_2336,In_2306,In_2135);
and U2337 (N_2337,In_2172,In_812);
and U2338 (N_2338,In_1432,In_2334);
and U2339 (N_2339,In_1399,In_407);
nand U2340 (N_2340,In_1762,In_2002);
or U2341 (N_2341,In_455,In_1428);
nor U2342 (N_2342,In_2286,In_2107);
and U2343 (N_2343,In_166,In_1367);
xor U2344 (N_2344,In_1121,In_1041);
nor U2345 (N_2345,In_2238,In_1257);
nand U2346 (N_2346,In_1395,In_865);
or U2347 (N_2347,In_1867,In_1227);
or U2348 (N_2348,In_2024,In_1728);
xnor U2349 (N_2349,In_270,In_1749);
nor U2350 (N_2350,In_1170,In_1872);
xnor U2351 (N_2351,In_634,In_454);
xnor U2352 (N_2352,In_903,In_601);
xnor U2353 (N_2353,In_1359,In_2042);
nor U2354 (N_2354,In_1429,In_1039);
nand U2355 (N_2355,In_818,In_762);
or U2356 (N_2356,In_802,In_985);
nand U2357 (N_2357,In_934,In_1677);
nor U2358 (N_2358,In_2256,In_431);
or U2359 (N_2359,In_1838,In_478);
and U2360 (N_2360,In_1623,In_886);
nand U2361 (N_2361,In_272,In_419);
nor U2362 (N_2362,In_2462,In_91);
and U2363 (N_2363,In_561,In_1791);
xnor U2364 (N_2364,In_608,In_920);
or U2365 (N_2365,In_2179,In_1575);
nand U2366 (N_2366,In_2159,In_2193);
nor U2367 (N_2367,In_675,In_2097);
nand U2368 (N_2368,In_2020,In_1202);
and U2369 (N_2369,In_522,In_2335);
and U2370 (N_2370,In_1727,In_2321);
or U2371 (N_2371,In_1732,In_1605);
or U2372 (N_2372,In_1826,In_2358);
xor U2373 (N_2373,In_1205,In_1435);
and U2374 (N_2374,In_686,In_1099);
and U2375 (N_2375,In_331,In_1417);
or U2376 (N_2376,In_560,In_1724);
nand U2377 (N_2377,In_385,In_479);
or U2378 (N_2378,In_51,In_1595);
and U2379 (N_2379,In_2113,In_342);
nand U2380 (N_2380,In_1653,In_948);
nand U2381 (N_2381,In_2357,In_1461);
or U2382 (N_2382,In_2185,In_1935);
or U2383 (N_2383,In_454,In_1081);
and U2384 (N_2384,In_1818,In_577);
nand U2385 (N_2385,In_2046,In_1970);
and U2386 (N_2386,In_1077,In_2041);
nand U2387 (N_2387,In_167,In_1267);
nand U2388 (N_2388,In_1472,In_1530);
nor U2389 (N_2389,In_379,In_770);
and U2390 (N_2390,In_329,In_894);
nand U2391 (N_2391,In_1896,In_1066);
and U2392 (N_2392,In_1273,In_1456);
xnor U2393 (N_2393,In_2043,In_1424);
or U2394 (N_2394,In_885,In_518);
or U2395 (N_2395,In_818,In_1486);
or U2396 (N_2396,In_156,In_1837);
nand U2397 (N_2397,In_2241,In_1625);
xor U2398 (N_2398,In_397,In_1463);
nor U2399 (N_2399,In_1248,In_96);
or U2400 (N_2400,In_1244,In_927);
xor U2401 (N_2401,In_124,In_1744);
or U2402 (N_2402,In_1683,In_2349);
nor U2403 (N_2403,In_2395,In_1410);
nor U2404 (N_2404,In_892,In_1619);
or U2405 (N_2405,In_356,In_1898);
and U2406 (N_2406,In_1846,In_1056);
and U2407 (N_2407,In_923,In_2318);
nor U2408 (N_2408,In_1127,In_1858);
or U2409 (N_2409,In_501,In_1828);
xnor U2410 (N_2410,In_2202,In_1755);
xor U2411 (N_2411,In_2467,In_987);
xor U2412 (N_2412,In_780,In_1231);
and U2413 (N_2413,In_1605,In_1180);
nand U2414 (N_2414,In_1491,In_635);
xor U2415 (N_2415,In_1208,In_815);
or U2416 (N_2416,In_1258,In_2267);
and U2417 (N_2417,In_1125,In_2119);
nor U2418 (N_2418,In_1688,In_411);
or U2419 (N_2419,In_1574,In_1605);
nor U2420 (N_2420,In_1866,In_860);
and U2421 (N_2421,In_2469,In_949);
nor U2422 (N_2422,In_381,In_2114);
and U2423 (N_2423,In_529,In_1876);
and U2424 (N_2424,In_32,In_205);
nand U2425 (N_2425,In_2108,In_358);
nand U2426 (N_2426,In_1495,In_501);
xor U2427 (N_2427,In_1241,In_1579);
nor U2428 (N_2428,In_748,In_686);
nand U2429 (N_2429,In_1745,In_1577);
or U2430 (N_2430,In_1889,In_1214);
and U2431 (N_2431,In_53,In_2367);
and U2432 (N_2432,In_1956,In_535);
and U2433 (N_2433,In_1466,In_1077);
and U2434 (N_2434,In_1472,In_1905);
nand U2435 (N_2435,In_2224,In_1896);
or U2436 (N_2436,In_136,In_1433);
nand U2437 (N_2437,In_758,In_822);
nand U2438 (N_2438,In_711,In_752);
and U2439 (N_2439,In_418,In_2361);
xor U2440 (N_2440,In_2466,In_864);
and U2441 (N_2441,In_889,In_1857);
xnor U2442 (N_2442,In_1662,In_349);
xnor U2443 (N_2443,In_1799,In_1711);
nand U2444 (N_2444,In_1340,In_831);
xnor U2445 (N_2445,In_2074,In_1796);
or U2446 (N_2446,In_273,In_726);
nand U2447 (N_2447,In_2482,In_879);
and U2448 (N_2448,In_252,In_2398);
nor U2449 (N_2449,In_2463,In_435);
nor U2450 (N_2450,In_104,In_1578);
nand U2451 (N_2451,In_2488,In_1182);
or U2452 (N_2452,In_2455,In_1600);
or U2453 (N_2453,In_691,In_638);
nor U2454 (N_2454,In_2052,In_224);
or U2455 (N_2455,In_2081,In_1806);
or U2456 (N_2456,In_74,In_1911);
and U2457 (N_2457,In_62,In_223);
and U2458 (N_2458,In_1684,In_127);
or U2459 (N_2459,In_447,In_517);
or U2460 (N_2460,In_953,In_1522);
or U2461 (N_2461,In_2210,In_1755);
or U2462 (N_2462,In_495,In_1147);
nand U2463 (N_2463,In_489,In_1749);
xnor U2464 (N_2464,In_1884,In_553);
and U2465 (N_2465,In_520,In_592);
nand U2466 (N_2466,In_626,In_533);
nand U2467 (N_2467,In_370,In_98);
xor U2468 (N_2468,In_2135,In_964);
nor U2469 (N_2469,In_429,In_2199);
xor U2470 (N_2470,In_446,In_1106);
nor U2471 (N_2471,In_333,In_1688);
or U2472 (N_2472,In_49,In_417);
xor U2473 (N_2473,In_2140,In_860);
xnor U2474 (N_2474,In_692,In_2395);
and U2475 (N_2475,In_1617,In_2186);
nand U2476 (N_2476,In_1453,In_1693);
xnor U2477 (N_2477,In_1539,In_1152);
xnor U2478 (N_2478,In_2092,In_1537);
nand U2479 (N_2479,In_558,In_1240);
nor U2480 (N_2480,In_1853,In_1886);
nor U2481 (N_2481,In_556,In_628);
nand U2482 (N_2482,In_1647,In_2185);
and U2483 (N_2483,In_1114,In_1985);
or U2484 (N_2484,In_1210,In_1700);
xor U2485 (N_2485,In_1992,In_772);
and U2486 (N_2486,In_1198,In_2391);
nand U2487 (N_2487,In_619,In_1258);
and U2488 (N_2488,In_102,In_1278);
and U2489 (N_2489,In_2209,In_1966);
and U2490 (N_2490,In_151,In_2482);
nand U2491 (N_2491,In_210,In_1603);
nand U2492 (N_2492,In_1061,In_966);
nand U2493 (N_2493,In_2143,In_2059);
nor U2494 (N_2494,In_670,In_1847);
nand U2495 (N_2495,In_1320,In_219);
nand U2496 (N_2496,In_1082,In_456);
or U2497 (N_2497,In_178,In_1769);
xnor U2498 (N_2498,In_1332,In_521);
nand U2499 (N_2499,In_61,In_2275);
nand U2500 (N_2500,N_1105,N_1425);
nor U2501 (N_2501,N_1397,N_851);
xor U2502 (N_2502,N_2271,N_40);
nand U2503 (N_2503,N_90,N_684);
and U2504 (N_2504,N_1324,N_1378);
and U2505 (N_2505,N_384,N_1242);
or U2506 (N_2506,N_1849,N_1075);
nor U2507 (N_2507,N_1808,N_1902);
nor U2508 (N_2508,N_2294,N_2014);
nor U2509 (N_2509,N_86,N_2045);
nor U2510 (N_2510,N_1540,N_1614);
and U2511 (N_2511,N_1405,N_1409);
nand U2512 (N_2512,N_2453,N_1975);
nand U2513 (N_2513,N_2024,N_125);
nand U2514 (N_2514,N_301,N_1213);
nor U2515 (N_2515,N_1644,N_2410);
or U2516 (N_2516,N_2197,N_83);
nor U2517 (N_2517,N_1571,N_264);
or U2518 (N_2518,N_1311,N_1946);
or U2519 (N_2519,N_1699,N_571);
or U2520 (N_2520,N_49,N_2223);
nor U2521 (N_2521,N_1132,N_1532);
or U2522 (N_2522,N_2140,N_1720);
and U2523 (N_2523,N_2021,N_2230);
and U2524 (N_2524,N_1257,N_149);
and U2525 (N_2525,N_2037,N_1286);
nand U2526 (N_2526,N_1044,N_2084);
nor U2527 (N_2527,N_1868,N_1756);
nand U2528 (N_2528,N_630,N_1907);
nand U2529 (N_2529,N_74,N_2270);
nand U2530 (N_2530,N_1106,N_65);
nor U2531 (N_2531,N_1154,N_1917);
xnor U2532 (N_2532,N_1028,N_898);
xnor U2533 (N_2533,N_1578,N_1003);
nand U2534 (N_2534,N_1847,N_1771);
and U2535 (N_2535,N_931,N_2411);
nor U2536 (N_2536,N_913,N_192);
nor U2537 (N_2537,N_2201,N_1527);
nand U2538 (N_2538,N_990,N_1231);
or U2539 (N_2539,N_126,N_1101);
nor U2540 (N_2540,N_1635,N_1321);
xnor U2541 (N_2541,N_2452,N_1099);
nor U2542 (N_2542,N_1663,N_191);
xnor U2543 (N_2543,N_1862,N_381);
nor U2544 (N_2544,N_1108,N_594);
nor U2545 (N_2545,N_521,N_2485);
nor U2546 (N_2546,N_878,N_1455);
or U2547 (N_2547,N_1301,N_600);
and U2548 (N_2548,N_2254,N_967);
nand U2549 (N_2549,N_2320,N_2013);
or U2550 (N_2550,N_661,N_813);
or U2551 (N_2551,N_429,N_518);
xnor U2552 (N_2552,N_1310,N_812);
xnor U2553 (N_2553,N_1822,N_665);
nand U2554 (N_2554,N_1131,N_1402);
nand U2555 (N_2555,N_441,N_275);
or U2556 (N_2556,N_585,N_918);
nand U2557 (N_2557,N_500,N_1208);
or U2558 (N_2558,N_958,N_1201);
and U2559 (N_2559,N_2180,N_1550);
nand U2560 (N_2560,N_2279,N_1485);
nor U2561 (N_2561,N_1495,N_2354);
nand U2562 (N_2562,N_1173,N_2399);
nand U2563 (N_2563,N_117,N_347);
nand U2564 (N_2564,N_1037,N_2095);
nor U2565 (N_2565,N_1512,N_775);
nand U2566 (N_2566,N_971,N_1556);
and U2567 (N_2567,N_448,N_2184);
or U2568 (N_2568,N_440,N_2402);
or U2569 (N_2569,N_1423,N_499);
or U2570 (N_2570,N_1992,N_262);
xnor U2571 (N_2571,N_830,N_1785);
nand U2572 (N_2572,N_21,N_1394);
nand U2573 (N_2573,N_1458,N_1240);
nand U2574 (N_2574,N_1912,N_758);
nor U2575 (N_2575,N_866,N_576);
nor U2576 (N_2576,N_2303,N_1831);
nand U2577 (N_2577,N_686,N_1491);
and U2578 (N_2578,N_1941,N_635);
or U2579 (N_2579,N_1668,N_614);
xor U2580 (N_2580,N_496,N_471);
and U2581 (N_2581,N_2128,N_260);
and U2582 (N_2582,N_1953,N_552);
or U2583 (N_2583,N_351,N_1928);
xnor U2584 (N_2584,N_1006,N_2169);
and U2585 (N_2585,N_2359,N_879);
xnor U2586 (N_2586,N_1730,N_1565);
xor U2587 (N_2587,N_422,N_1178);
nor U2588 (N_2588,N_488,N_999);
nor U2589 (N_2589,N_357,N_487);
and U2590 (N_2590,N_2446,N_2383);
nor U2591 (N_2591,N_657,N_2390);
nor U2592 (N_2592,N_1329,N_1032);
xnor U2593 (N_2593,N_1399,N_162);
xor U2594 (N_2594,N_1770,N_1783);
nand U2595 (N_2595,N_2412,N_1288);
nand U2596 (N_2596,N_2031,N_2034);
nor U2597 (N_2597,N_724,N_826);
nor U2598 (N_2598,N_1843,N_829);
xor U2599 (N_2599,N_1384,N_2490);
or U2600 (N_2600,N_281,N_757);
or U2601 (N_2601,N_2454,N_1176);
xor U2602 (N_2602,N_29,N_1277);
nand U2603 (N_2603,N_2160,N_1990);
and U2604 (N_2604,N_2398,N_2442);
nor U2605 (N_2605,N_966,N_823);
nor U2606 (N_2606,N_368,N_1871);
nand U2607 (N_2607,N_1905,N_1183);
nand U2608 (N_2608,N_911,N_1833);
nand U2609 (N_2609,N_1219,N_315);
nand U2610 (N_2610,N_490,N_222);
nand U2611 (N_2611,N_326,N_1657);
or U2612 (N_2612,N_166,N_2121);
or U2613 (N_2613,N_1389,N_842);
nor U2614 (N_2614,N_1093,N_160);
nand U2615 (N_2615,N_1189,N_1387);
nand U2616 (N_2616,N_1145,N_1320);
or U2617 (N_2617,N_921,N_1563);
xnor U2618 (N_2618,N_602,N_401);
and U2619 (N_2619,N_1625,N_182);
xor U2620 (N_2620,N_1471,N_1169);
or U2621 (N_2621,N_1237,N_133);
or U2622 (N_2622,N_2185,N_1944);
nand U2623 (N_2623,N_2264,N_2311);
or U2624 (N_2624,N_556,N_1197);
or U2625 (N_2625,N_104,N_863);
xor U2626 (N_2626,N_456,N_982);
nand U2627 (N_2627,N_867,N_330);
nor U2628 (N_2628,N_916,N_450);
xor U2629 (N_2629,N_466,N_2081);
xor U2630 (N_2630,N_1365,N_1890);
xor U2631 (N_2631,N_1008,N_2335);
nand U2632 (N_2632,N_2478,N_20);
and U2633 (N_2633,N_1517,N_1129);
nor U2634 (N_2634,N_1791,N_719);
nand U2635 (N_2635,N_1906,N_1504);
or U2636 (N_2636,N_1782,N_1306);
or U2637 (N_2637,N_547,N_1470);
nand U2638 (N_2638,N_1830,N_1066);
nor U2639 (N_2639,N_1124,N_1986);
nand U2640 (N_2640,N_1874,N_721);
nor U2641 (N_2641,N_93,N_409);
or U2642 (N_2642,N_962,N_1530);
and U2643 (N_2643,N_572,N_1104);
or U2644 (N_2644,N_1741,N_1943);
nor U2645 (N_2645,N_1837,N_2124);
and U2646 (N_2646,N_212,N_1865);
nand U2647 (N_2647,N_1621,N_1376);
xnor U2648 (N_2648,N_324,N_1174);
xor U2649 (N_2649,N_1056,N_204);
or U2650 (N_2650,N_2167,N_1701);
and U2651 (N_2651,N_1395,N_1279);
or U2652 (N_2652,N_716,N_1422);
or U2653 (N_2653,N_1980,N_2087);
xor U2654 (N_2654,N_1616,N_687);
or U2655 (N_2655,N_871,N_1887);
xnor U2656 (N_2656,N_1924,N_1893);
and U2657 (N_2657,N_2208,N_700);
nand U2658 (N_2658,N_1448,N_1745);
xor U2659 (N_2659,N_1936,N_1048);
or U2660 (N_2660,N_1244,N_1488);
xor U2661 (N_2661,N_1337,N_2377);
nor U2662 (N_2662,N_185,N_523);
or U2663 (N_2663,N_2206,N_625);
or U2664 (N_2664,N_905,N_1053);
or U2665 (N_2665,N_1536,N_1866);
and U2666 (N_2666,N_112,N_2198);
nand U2667 (N_2667,N_819,N_987);
nand U2668 (N_2668,N_1267,N_751);
xnor U2669 (N_2669,N_291,N_2257);
xnor U2670 (N_2670,N_1526,N_1648);
nand U2671 (N_2671,N_2434,N_1272);
xnor U2672 (N_2672,N_1679,N_106);
xor U2673 (N_2673,N_1476,N_1004);
xor U2674 (N_2674,N_1241,N_1554);
nand U2675 (N_2675,N_1025,N_1680);
xor U2676 (N_2676,N_2115,N_411);
xor U2677 (N_2677,N_235,N_2414);
nor U2678 (N_2678,N_1092,N_1913);
nor U2679 (N_2679,N_1243,N_1019);
and U2680 (N_2680,N_553,N_1147);
and U2681 (N_2681,N_1901,N_588);
xor U2682 (N_2682,N_459,N_2375);
nand U2683 (N_2683,N_304,N_2464);
nand U2684 (N_2684,N_1542,N_135);
and U2685 (N_2685,N_814,N_203);
or U2686 (N_2686,N_1418,N_855);
or U2687 (N_2687,N_2236,N_712);
nor U2688 (N_2688,N_2226,N_1031);
or U2689 (N_2689,N_749,N_1665);
nand U2690 (N_2690,N_37,N_654);
or U2691 (N_2691,N_1546,N_2248);
nand U2692 (N_2692,N_1118,N_1850);
and U2693 (N_2693,N_802,N_1691);
nand U2694 (N_2694,N_1718,N_1065);
xnor U2695 (N_2695,N_1146,N_877);
nor U2696 (N_2696,N_1689,N_1962);
nand U2697 (N_2697,N_2176,N_1584);
nor U2698 (N_2698,N_662,N_2360);
nor U2699 (N_2699,N_1144,N_1360);
nor U2700 (N_2700,N_1411,N_1851);
nand U2701 (N_2701,N_1179,N_831);
nand U2702 (N_2702,N_525,N_992);
and U2703 (N_2703,N_590,N_428);
or U2704 (N_2704,N_2437,N_178);
or U2705 (N_2705,N_385,N_2018);
nand U2706 (N_2706,N_472,N_1891);
nor U2707 (N_2707,N_954,N_984);
nor U2708 (N_2708,N_2344,N_559);
nor U2709 (N_2709,N_1282,N_2302);
xnor U2710 (N_2710,N_52,N_1062);
and U2711 (N_2711,N_2090,N_1463);
and U2712 (N_2712,N_1723,N_2225);
or U2713 (N_2713,N_551,N_467);
xor U2714 (N_2714,N_1192,N_2425);
nand U2715 (N_2715,N_1172,N_1915);
xor U2716 (N_2716,N_2165,N_101);
nor U2717 (N_2717,N_198,N_312);
nor U2718 (N_2718,N_1230,N_2307);
nand U2719 (N_2719,N_1452,N_1073);
and U2720 (N_2720,N_1807,N_2119);
or U2721 (N_2721,N_298,N_1007);
and U2722 (N_2722,N_1572,N_1030);
xnor U2723 (N_2723,N_682,N_2445);
xor U2724 (N_2724,N_10,N_822);
and U2725 (N_2725,N_583,N_1327);
nand U2726 (N_2726,N_2181,N_1894);
nor U2727 (N_2727,N_2083,N_24);
nand U2728 (N_2728,N_451,N_2423);
xor U2729 (N_2729,N_1352,N_1731);
or U2730 (N_2730,N_161,N_900);
nor U2731 (N_2731,N_2373,N_2483);
or U2732 (N_2732,N_1513,N_2186);
and U2733 (N_2733,N_978,N_2409);
nand U2734 (N_2734,N_850,N_1743);
xor U2735 (N_2735,N_2178,N_295);
nand U2736 (N_2736,N_1567,N_2238);
xor U2737 (N_2737,N_1564,N_1607);
nor U2738 (N_2738,N_142,N_736);
nor U2739 (N_2739,N_663,N_2155);
and U2740 (N_2740,N_80,N_1303);
nand U2741 (N_2741,N_270,N_1878);
or U2742 (N_2742,N_1520,N_693);
nand U2743 (N_2743,N_604,N_225);
nor U2744 (N_2744,N_1670,N_68);
xnor U2745 (N_2745,N_329,N_2154);
nor U2746 (N_2746,N_1225,N_2417);
xor U2747 (N_2747,N_1253,N_2156);
xnor U2748 (N_2748,N_710,N_405);
and U2749 (N_2749,N_857,N_1149);
xor U2750 (N_2750,N_2227,N_2202);
xor U2751 (N_2751,N_1459,N_948);
or U2752 (N_2752,N_1710,N_1909);
nor U2753 (N_2753,N_1400,N_1061);
nor U2754 (N_2754,N_915,N_1610);
xor U2755 (N_2755,N_2372,N_2144);
xor U2756 (N_2756,N_1350,N_1000);
nor U2757 (N_2757,N_263,N_766);
and U2758 (N_2758,N_2350,N_2448);
nor U2759 (N_2759,N_1515,N_1182);
and U2760 (N_2760,N_189,N_322);
xor U2761 (N_2761,N_1134,N_765);
xnor U2762 (N_2762,N_36,N_591);
and U2763 (N_2763,N_1194,N_1292);
or U2764 (N_2764,N_1033,N_1826);
or U2765 (N_2765,N_337,N_2132);
nor U2766 (N_2766,N_2138,N_752);
nand U2767 (N_2767,N_1739,N_1074);
or U2768 (N_2768,N_1744,N_1406);
and U2769 (N_2769,N_1507,N_251);
or U2770 (N_2770,N_582,N_2346);
or U2771 (N_2771,N_1187,N_720);
and U2772 (N_2772,N_239,N_926);
or U2773 (N_2773,N_1768,N_1503);
xnor U2774 (N_2774,N_1587,N_1976);
xor U2775 (N_2775,N_649,N_2053);
xnor U2776 (N_2776,N_1102,N_753);
or U2777 (N_2777,N_1199,N_2370);
nor U2778 (N_2778,N_668,N_1346);
and U2779 (N_2779,N_1140,N_2241);
or U2780 (N_2780,N_942,N_60);
and U2781 (N_2781,N_1840,N_2097);
nand U2782 (N_2782,N_2430,N_904);
or U2783 (N_2783,N_803,N_2352);
nor U2784 (N_2784,N_2322,N_1261);
nor U2785 (N_2785,N_1640,N_2127);
nand U2786 (N_2786,N_435,N_229);
and U2787 (N_2787,N_2030,N_240);
xor U2788 (N_2788,N_961,N_1070);
or U2789 (N_2789,N_2317,N_792);
nor U2790 (N_2790,N_728,N_1753);
nand U2791 (N_2791,N_430,N_387);
nand U2792 (N_2792,N_159,N_542);
or U2793 (N_2793,N_1045,N_1354);
xor U2794 (N_2794,N_1466,N_1068);
or U2795 (N_2795,N_1934,N_1895);
and U2796 (N_2796,N_1453,N_1800);
nor U2797 (N_2797,N_1995,N_314);
or U2798 (N_2798,N_1612,N_2111);
xnor U2799 (N_2799,N_2382,N_417);
nor U2800 (N_2800,N_1064,N_2469);
and U2801 (N_2801,N_1022,N_534);
nand U2802 (N_2802,N_2331,N_1393);
nand U2803 (N_2803,N_2462,N_1383);
nand U2804 (N_2804,N_416,N_1165);
and U2805 (N_2805,N_1776,N_1930);
nor U2806 (N_2806,N_2476,N_163);
xor U2807 (N_2807,N_2285,N_1265);
or U2808 (N_2808,N_1712,N_2336);
nand U2809 (N_2809,N_1467,N_2432);
nor U2810 (N_2810,N_1672,N_1855);
xor U2811 (N_2811,N_664,N_545);
nor U2812 (N_2812,N_550,N_1100);
nand U2813 (N_2813,N_1658,N_2357);
nor U2814 (N_2814,N_1939,N_619);
and U2815 (N_2815,N_2460,N_1523);
xor U2816 (N_2816,N_1886,N_1666);
and U2817 (N_2817,N_1643,N_2195);
nor U2818 (N_2818,N_1835,N_1859);
xnor U2819 (N_2819,N_1561,N_2096);
nor U2820 (N_2820,N_638,N_1198);
xor U2821 (N_2821,N_1287,N_2422);
or U2822 (N_2822,N_660,N_2055);
nor U2823 (N_2823,N_2300,N_2282);
or U2824 (N_2824,N_1150,N_296);
or U2825 (N_2825,N_343,N_784);
xor U2826 (N_2826,N_17,N_759);
or U2827 (N_2827,N_612,N_566);
or U2828 (N_2828,N_1298,N_461);
nand U2829 (N_2829,N_2190,N_1212);
and U2830 (N_2830,N_1325,N_2351);
or U2831 (N_2831,N_1846,N_2209);
nand U2832 (N_2832,N_214,N_50);
nand U2833 (N_2833,N_1275,N_586);
nand U2834 (N_2834,N_1763,N_308);
xor U2835 (N_2835,N_1366,N_2228);
xor U2836 (N_2836,N_640,N_1656);
xor U2837 (N_2837,N_2353,N_2116);
and U2838 (N_2838,N_1649,N_769);
xor U2839 (N_2839,N_1401,N_2072);
or U2840 (N_2840,N_2301,N_933);
and U2841 (N_2841,N_1864,N_1332);
xnor U2842 (N_2842,N_1775,N_1605);
nand U2843 (N_2843,N_1338,N_383);
and U2844 (N_2844,N_1618,N_891);
and U2845 (N_2845,N_883,N_48);
xor U2846 (N_2846,N_530,N_2249);
nor U2847 (N_2847,N_951,N_474);
nor U2848 (N_2848,N_1996,N_1693);
nor U2849 (N_2849,N_1997,N_102);
nand U2850 (N_2850,N_1426,N_620);
nor U2851 (N_2851,N_1067,N_2468);
or U2852 (N_2852,N_1040,N_509);
or U2853 (N_2853,N_2405,N_2444);
nand U2854 (N_2854,N_2361,N_1398);
and U2855 (N_2855,N_398,N_1318);
nor U2856 (N_2856,N_1234,N_1499);
and U2857 (N_2857,N_669,N_725);
nor U2858 (N_2858,N_893,N_1494);
xnor U2859 (N_2859,N_1857,N_965);
nand U2860 (N_2860,N_15,N_2214);
xnor U2861 (N_2861,N_2449,N_1942);
nand U2862 (N_2862,N_1081,N_2416);
xnor U2863 (N_2863,N_470,N_1012);
nand U2864 (N_2864,N_828,N_1266);
nor U2865 (N_2865,N_1415,N_183);
nand U2866 (N_2866,N_152,N_1188);
or U2867 (N_2867,N_2137,N_1562);
nand U2868 (N_2868,N_2232,N_390);
and U2869 (N_2869,N_1017,N_1974);
nand U2870 (N_2870,N_1603,N_1164);
xnor U2871 (N_2871,N_1109,N_1602);
nand U2872 (N_2872,N_672,N_841);
or U2873 (N_2873,N_1137,N_1246);
and U2874 (N_2874,N_364,N_699);
nand U2875 (N_2875,N_205,N_1681);
or U2876 (N_2876,N_678,N_2349);
nand U2877 (N_2877,N_278,N_1335);
nor U2878 (N_2878,N_12,N_696);
nor U2879 (N_2879,N_1881,N_1421);
nor U2880 (N_2880,N_1715,N_318);
xor U2881 (N_2881,N_890,N_341);
or U2882 (N_2882,N_7,N_2080);
or U2883 (N_2883,N_2146,N_202);
xnor U2884 (N_2884,N_895,N_2028);
nand U2885 (N_2885,N_1589,N_292);
nand U2886 (N_2886,N_1464,N_2158);
nand U2887 (N_2887,N_811,N_998);
or U2888 (N_2888,N_835,N_1594);
nor U2889 (N_2889,N_917,N_1058);
xor U2890 (N_2890,N_1049,N_2170);
and U2891 (N_2891,N_276,N_2493);
nand U2892 (N_2892,N_1799,N_1334);
nor U2893 (N_2893,N_484,N_748);
xnor U2894 (N_2894,N_1889,N_1412);
xnor U2895 (N_2895,N_1343,N_976);
nand U2896 (N_2896,N_1461,N_1071);
or U2897 (N_2897,N_1323,N_1035);
nor U2898 (N_2898,N_762,N_656);
nor U2899 (N_2899,N_473,N_558);
nand U2900 (N_2900,N_285,N_1856);
xnor U2901 (N_2901,N_1873,N_869);
and U2902 (N_2902,N_676,N_1965);
and U2903 (N_2903,N_476,N_87);
nor U2904 (N_2904,N_28,N_1623);
nor U2905 (N_2905,N_1671,N_360);
nor U2906 (N_2906,N_2441,N_1861);
nor U2907 (N_2907,N_1255,N_146);
xnor U2908 (N_2908,N_8,N_194);
xor U2909 (N_2909,N_616,N_2059);
xnor U2910 (N_2910,N_1449,N_1970);
nor U2911 (N_2911,N_1755,N_889);
nor U2912 (N_2912,N_1591,N_2193);
or U2913 (N_2913,N_613,N_772);
nand U2914 (N_2914,N_592,N_2288);
and U2915 (N_2915,N_702,N_1410);
nand U2916 (N_2916,N_1940,N_30);
nor U2917 (N_2917,N_1500,N_912);
and U2918 (N_2918,N_1259,N_2110);
nand U2919 (N_2919,N_711,N_46);
or U2920 (N_2920,N_968,N_2340);
or U2921 (N_2921,N_914,N_2192);
xnor U2922 (N_2922,N_653,N_2025);
nor U2923 (N_2923,N_750,N_1372);
nand U2924 (N_2924,N_601,N_2321);
or U2925 (N_2925,N_2187,N_497);
or U2926 (N_2926,N_524,N_1604);
or U2927 (N_2927,N_1722,N_1299);
xnor U2928 (N_2928,N_406,N_833);
and U2929 (N_2929,N_375,N_2079);
or U2930 (N_2930,N_642,N_23);
and U2931 (N_2931,N_1424,N_1686);
nand U2932 (N_2932,N_888,N_1795);
or U2933 (N_2933,N_1609,N_2039);
nand U2934 (N_2934,N_1456,N_271);
and U2935 (N_2935,N_336,N_1597);
and U2936 (N_2936,N_369,N_902);
and U2937 (N_2937,N_1828,N_892);
and U2938 (N_2938,N_674,N_1283);
and U2939 (N_2939,N_1063,N_1392);
and U2940 (N_2940,N_1796,N_1043);
xnor U2941 (N_2941,N_305,N_1186);
nor U2942 (N_2942,N_1832,N_209);
and U2943 (N_2943,N_1114,N_354);
and U2944 (N_2944,N_1949,N_408);
xor U2945 (N_2945,N_1420,N_703);
or U2946 (N_2946,N_2172,N_937);
nand U2947 (N_2947,N_1695,N_731);
nand U2948 (N_2948,N_1543,N_206);
nand U2949 (N_2949,N_2329,N_1727);
nor U2950 (N_2950,N_1854,N_564);
and U2951 (N_2951,N_947,N_1364);
and U2952 (N_2952,N_1447,N_2296);
or U2953 (N_2953,N_2269,N_1460);
xor U2954 (N_2954,N_977,N_1304);
and U2955 (N_2955,N_2290,N_2457);
xor U2956 (N_2956,N_2112,N_1433);
nand U2957 (N_2957,N_632,N_565);
nand U2958 (N_2958,N_1501,N_84);
xnor U2959 (N_2959,N_2343,N_213);
and U2960 (N_2960,N_1780,N_493);
nor U2961 (N_2961,N_2036,N_929);
or U2962 (N_2962,N_2345,N_771);
xor U2963 (N_2963,N_151,N_1836);
nor U2964 (N_2964,N_2488,N_389);
xnor U2965 (N_2965,N_963,N_1682);
and U2966 (N_2966,N_1051,N_1489);
xnor U2967 (N_2967,N_1362,N_2207);
xor U2968 (N_2968,N_64,N_216);
nor U2969 (N_2969,N_1593,N_503);
nand U2970 (N_2970,N_2211,N_1687);
nor U2971 (N_2971,N_1396,N_115);
or U2972 (N_2972,N_870,N_1711);
or U2973 (N_2973,N_243,N_33);
nand U2974 (N_2974,N_2348,N_2094);
xor U2975 (N_2975,N_1271,N_174);
nand U2976 (N_2976,N_1370,N_453);
and U2977 (N_2977,N_1956,N_598);
nand U2978 (N_2978,N_568,N_1300);
or U2979 (N_2979,N_1803,N_936);
nor U2980 (N_2980,N_1232,N_2103);
nor U2981 (N_2981,N_2009,N_412);
xnor U2982 (N_2982,N_1652,N_128);
xor U2983 (N_2983,N_1380,N_338);
nand U2984 (N_2984,N_274,N_1709);
and U2985 (N_2985,N_2293,N_739);
nand U2986 (N_2986,N_745,N_2489);
or U2987 (N_2987,N_1059,N_1737);
or U2988 (N_2988,N_2265,N_1445);
or U2989 (N_2989,N_426,N_1586);
and U2990 (N_2990,N_373,N_2050);
nor U2991 (N_2991,N_1631,N_907);
and U2992 (N_2992,N_498,N_1202);
or U2993 (N_2993,N_111,N_223);
nor U2994 (N_2994,N_420,N_494);
nand U2995 (N_2995,N_1457,N_2327);
or U2996 (N_2996,N_1087,N_2404);
xor U2997 (N_2997,N_254,N_1369);
xor U2998 (N_2998,N_580,N_876);
or U2999 (N_2999,N_1312,N_513);
nand U3000 (N_3000,N_1293,N_2125);
and U3001 (N_3001,N_647,N_927);
and U3002 (N_3002,N_366,N_231);
nor U3003 (N_3003,N_2438,N_2066);
or U3004 (N_3004,N_1998,N_395);
or U3005 (N_3005,N_70,N_516);
or U3006 (N_3006,N_2129,N_574);
xor U3007 (N_3007,N_579,N_145);
and U3008 (N_3008,N_31,N_455);
nand U3009 (N_3009,N_1223,N_1291);
xnor U3010 (N_3010,N_1929,N_2306);
nand U3011 (N_3011,N_201,N_1606);
xor U3012 (N_3012,N_1437,N_247);
and U3013 (N_3013,N_1027,N_284);
nor U3014 (N_3014,N_439,N_1585);
or U3015 (N_3015,N_1967,N_167);
nor U3016 (N_3016,N_779,N_2260);
nor U3017 (N_3017,N_2243,N_622);
and U3018 (N_3018,N_1853,N_1309);
and U3019 (N_3019,N_1883,N_639);
or U3020 (N_3020,N_2316,N_655);
nor U3021 (N_3021,N_1838,N_349);
xor U3022 (N_3022,N_2047,N_1789);
nor U3023 (N_3023,N_1079,N_1294);
nand U3024 (N_3024,N_2466,N_717);
or U3025 (N_3025,N_539,N_1440);
xnor U3026 (N_3026,N_1898,N_1772);
xor U3027 (N_3027,N_1802,N_2374);
nand U3028 (N_3028,N_1361,N_449);
nand U3029 (N_3029,N_1875,N_952);
and U3030 (N_3030,N_1764,N_1575);
or U3031 (N_3031,N_123,N_554);
or U3032 (N_3032,N_2149,N_2308);
nor U3033 (N_3033,N_973,N_2484);
and U3034 (N_3034,N_722,N_1948);
and U3035 (N_3035,N_2280,N_460);
nor U3036 (N_3036,N_1381,N_2250);
or U3037 (N_3037,N_1496,N_2251);
and U3038 (N_3038,N_14,N_1841);
or U3039 (N_3039,N_1014,N_570);
nor U3040 (N_3040,N_587,N_2171);
and U3041 (N_3041,N_1493,N_2439);
nor U3042 (N_3042,N_943,N_1227);
nor U3043 (N_3043,N_1475,N_362);
nand U3044 (N_3044,N_981,N_1641);
nor U3045 (N_3045,N_78,N_1762);
and U3046 (N_3046,N_515,N_2486);
nand U3047 (N_3047,N_1834,N_746);
or U3048 (N_3048,N_980,N_882);
or U3049 (N_3049,N_2048,N_705);
nor U3050 (N_3050,N_2042,N_136);
xnor U3051 (N_3051,N_543,N_2380);
nor U3052 (N_3052,N_1094,N_1193);
or U3053 (N_3053,N_1982,N_230);
and U3054 (N_3054,N_934,N_2063);
nand U3055 (N_3055,N_1115,N_1884);
nand U3056 (N_3056,N_1175,N_709);
nand U3057 (N_3057,N_740,N_2276);
nand U3058 (N_3058,N_2255,N_1914);
and U3059 (N_3059,N_1076,N_371);
nand U3060 (N_3060,N_1617,N_190);
xnor U3061 (N_3061,N_1206,N_1158);
or U3062 (N_3062,N_708,N_47);
xnor U3063 (N_3063,N_98,N_2341);
xnor U3064 (N_3064,N_256,N_2075);
nor U3065 (N_3065,N_520,N_1704);
nand U3066 (N_3066,N_1136,N_1978);
nor U3067 (N_3067,N_2135,N_1746);
nand U3068 (N_3068,N_1698,N_704);
nor U3069 (N_3069,N_1664,N_2070);
or U3070 (N_3070,N_150,N_1794);
nand U3071 (N_3071,N_2164,N_581);
xor U3072 (N_3072,N_2355,N_454);
xnor U3073 (N_3073,N_141,N_2440);
xnor U3074 (N_3074,N_1,N_561);
nor U3075 (N_3075,N_257,N_548);
nor U3076 (N_3076,N_1307,N_2256);
nand U3077 (N_3077,N_1233,N_868);
nor U3078 (N_3078,N_1702,N_2487);
nand U3079 (N_3079,N_2235,N_79);
or U3080 (N_3080,N_846,N_1221);
xor U3081 (N_3081,N_1142,N_1024);
or U3082 (N_3082,N_1340,N_754);
and U3083 (N_3083,N_2213,N_226);
and U3084 (N_3084,N_1462,N_1600);
nor U3085 (N_3085,N_540,N_137);
and U3086 (N_3086,N_1708,N_2106);
or U3087 (N_3087,N_1126,N_1817);
nand U3088 (N_3088,N_789,N_1825);
nor U3089 (N_3089,N_1792,N_334);
or U3090 (N_3090,N_2379,N_1903);
xnor U3091 (N_3091,N_730,N_1305);
nand U3092 (N_3092,N_1778,N_391);
or U3093 (N_3093,N_1880,N_1633);
nor U3094 (N_3094,N_2049,N_1729);
xor U3095 (N_3095,N_627,N_675);
or U3096 (N_3096,N_2408,N_1055);
nor U3097 (N_3097,N_2458,N_2054);
nor U3098 (N_3098,N_2314,N_1683);
nor U3099 (N_3099,N_1313,N_501);
nand U3100 (N_3100,N_1011,N_9);
or U3101 (N_3101,N_2007,N_994);
nor U3102 (N_3102,N_925,N_634);
nand U3103 (N_3103,N_1373,N_538);
and U3104 (N_3104,N_1427,N_238);
or U3105 (N_3105,N_1547,N_2407);
or U3106 (N_3106,N_2245,N_2283);
nand U3107 (N_3107,N_2347,N_2391);
nand U3108 (N_3108,N_1773,N_2363);
and U3109 (N_3109,N_1528,N_58);
and U3110 (N_3110,N_1482,N_1654);
and U3111 (N_3111,N_2093,N_1688);
nand U3112 (N_3112,N_1931,N_234);
and U3113 (N_3113,N_155,N_1879);
xor U3114 (N_3114,N_2284,N_2065);
or U3115 (N_3115,N_932,N_2342);
and U3116 (N_3116,N_2289,N_56);
and U3117 (N_3117,N_1767,N_575);
nand U3118 (N_3118,N_1443,N_1029);
or U3119 (N_3119,N_2074,N_1568);
nor U3120 (N_3120,N_332,N_348);
nand U3121 (N_3121,N_1858,N_852);
xnor U3122 (N_3122,N_1694,N_1863);
and U3123 (N_3123,N_1296,N_795);
xnor U3124 (N_3124,N_1010,N_1904);
nand U3125 (N_3125,N_2189,N_1353);
nor U3126 (N_3126,N_1787,N_2141);
nor U3127 (N_3127,N_2118,N_805);
or U3128 (N_3128,N_532,N_277);
and U3129 (N_3129,N_444,N_2498);
nor U3130 (N_3130,N_228,N_431);
xor U3131 (N_3131,N_2461,N_1541);
nand U3132 (N_3132,N_1820,N_2191);
nand U3133 (N_3133,N_1829,N_2062);
or U3134 (N_3134,N_1660,N_199);
nor U3135 (N_3135,N_447,N_2313);
xnor U3136 (N_3136,N_1347,N_886);
or U3137 (N_3137,N_806,N_2210);
or U3138 (N_3138,N_217,N_1926);
and U3139 (N_3139,N_4,N_637);
xnor U3140 (N_3140,N_560,N_2261);
or U3141 (N_3141,N_2401,N_727);
or U3142 (N_3142,N_608,N_1374);
and U3143 (N_3143,N_2499,N_363);
nand U3144 (N_3144,N_2085,N_1156);
and U3145 (N_3145,N_1662,N_1957);
nor U3146 (N_3146,N_1509,N_1148);
and U3147 (N_3147,N_290,N_818);
xor U3148 (N_3148,N_1958,N_793);
or U3149 (N_3149,N_679,N_599);
nor U3150 (N_3150,N_1774,N_1263);
and U3151 (N_3151,N_1368,N_1359);
xnor U3152 (N_3152,N_1379,N_1050);
nor U3153 (N_3153,N_1637,N_744);
and U3154 (N_3154,N_1516,N_935);
or U3155 (N_3155,N_2000,N_11);
nor U3156 (N_3156,N_648,N_1973);
and U3157 (N_3157,N_733,N_2233);
and U3158 (N_3158,N_376,N_2029);
nand U3159 (N_3159,N_1057,N_1434);
xnor U3160 (N_3160,N_1228,N_1581);
nor U3161 (N_3161,N_1431,N_1908);
xnor U3162 (N_3162,N_517,N_219);
nand U3163 (N_3163,N_519,N_1921);
xor U3164 (N_3164,N_2153,N_261);
or U3165 (N_3165,N_741,N_1673);
and U3166 (N_3166,N_1220,N_2397);
nand U3167 (N_3167,N_2392,N_258);
xor U3168 (N_3168,N_1439,N_2330);
and U3169 (N_3169,N_808,N_2447);
nand U3170 (N_3170,N_1117,N_1531);
and U3171 (N_3171,N_69,N_860);
xor U3172 (N_3172,N_1082,N_2002);
nand U3173 (N_3173,N_791,N_844);
nand U3174 (N_3174,N_164,N_134);
nor U3175 (N_3175,N_1638,N_241);
xor U3176 (N_3176,N_595,N_89);
and U3177 (N_3177,N_1155,N_1249);
or U3178 (N_3178,N_1248,N_1180);
nand U3179 (N_3179,N_2456,N_1506);
or U3180 (N_3180,N_2339,N_970);
nor U3181 (N_3181,N_1927,N_379);
xnor U3182 (N_3182,N_1899,N_1734);
nor U3183 (N_3183,N_631,N_2060);
nand U3184 (N_3184,N_2413,N_252);
or U3185 (N_3185,N_2113,N_1922);
xor U3186 (N_3186,N_2471,N_2200);
nor U3187 (N_3187,N_1278,N_1235);
or U3188 (N_3188,N_196,N_1385);
nor U3189 (N_3189,N_1716,N_2386);
and U3190 (N_3190,N_1264,N_280);
nor U3191 (N_3191,N_1416,N_1450);
and U3192 (N_3192,N_1548,N_1153);
or U3193 (N_3193,N_2133,N_2281);
or U3194 (N_3194,N_974,N_1357);
nor U3195 (N_3195,N_2263,N_1205);
xnor U3196 (N_3196,N_861,N_755);
or U3197 (N_3197,N_2323,N_633);
or U3198 (N_3198,N_945,N_815);
and U3199 (N_3199,N_923,N_197);
and U3200 (N_3200,N_1436,N_1636);
or U3201 (N_3201,N_253,N_2384);
nor U3202 (N_3202,N_1419,N_1166);
and U3203 (N_3203,N_1328,N_386);
xnor U3204 (N_3204,N_2091,N_1678);
or U3205 (N_3205,N_848,N_2136);
nand U3206 (N_3206,N_1993,N_1121);
xor U3207 (N_3207,N_394,N_1474);
nor U3208 (N_3208,N_53,N_2041);
nor U3209 (N_3209,N_997,N_1814);
nand U3210 (N_3210,N_1315,N_403);
nand U3211 (N_3211,N_1968,N_414);
nor U3212 (N_3212,N_313,N_1812);
nand U3213 (N_3213,N_169,N_825);
xor U3214 (N_3214,N_1122,N_181);
xnor U3215 (N_3215,N_51,N_2267);
or U3216 (N_3216,N_153,N_939);
nand U3217 (N_3217,N_45,N_1954);
and U3218 (N_3218,N_1615,N_404);
xnor U3219 (N_3219,N_2328,N_489);
and U3220 (N_3220,N_1650,N_140);
nor U3221 (N_3221,N_1130,N_767);
xnor U3222 (N_3222,N_2315,N_41);
and U3223 (N_3223,N_1280,N_361);
or U3224 (N_3224,N_1821,N_107);
and U3225 (N_3225,N_1285,N_2120);
and U3226 (N_3226,N_1816,N_732);
xor U3227 (N_3227,N_906,N_1218);
nor U3228 (N_3228,N_1444,N_1167);
xor U3229 (N_3229,N_1583,N_991);
xor U3230 (N_3230,N_701,N_1386);
nand U3231 (N_3231,N_743,N_319);
and U3232 (N_3232,N_2131,N_1181);
and U3233 (N_3233,N_2204,N_157);
xor U3234 (N_3234,N_1435,N_2292);
or U3235 (N_3235,N_688,N_940);
nor U3236 (N_3236,N_1119,N_2385);
xor U3237 (N_3237,N_402,N_1157);
nor U3238 (N_3238,N_641,N_62);
xor U3239 (N_3239,N_667,N_2455);
nor U3240 (N_3240,N_1091,N_1598);
nand U3241 (N_3241,N_874,N_1196);
or U3242 (N_3242,N_2395,N_55);
nand U3243 (N_3243,N_22,N_611);
xor U3244 (N_3244,N_2123,N_845);
nor U3245 (N_3245,N_287,N_221);
and U3246 (N_3246,N_1534,N_506);
nor U3247 (N_3247,N_1983,N_457);
xnor U3248 (N_3248,N_250,N_1713);
and U3249 (N_3249,N_1341,N_2088);
nor U3250 (N_3250,N_356,N_677);
and U3251 (N_3251,N_1777,N_706);
or U3252 (N_3252,N_1524,N_816);
nand U3253 (N_3253,N_432,N_666);
nor U3254 (N_3254,N_171,N_1811);
or U3255 (N_3255,N_442,N_1023);
xnor U3256 (N_3256,N_2015,N_2108);
nand U3257 (N_3257,N_2494,N_2337);
nand U3258 (N_3258,N_790,N_1200);
xor U3259 (N_3259,N_355,N_1797);
and U3260 (N_3260,N_2064,N_2092);
xnor U3261 (N_3261,N_901,N_569);
nand U3262 (N_3262,N_1111,N_302);
nor U3263 (N_3263,N_1209,N_1159);
nor U3264 (N_3264,N_885,N_2179);
xnor U3265 (N_3265,N_986,N_956);
and U3266 (N_3266,N_413,N_207);
nor U3267 (N_3267,N_2277,N_421);
nor U3268 (N_3268,N_44,N_1502);
and U3269 (N_3269,N_2067,N_2073);
or U3270 (N_3270,N_1331,N_536);
xor U3271 (N_3271,N_1726,N_1498);
or U3272 (N_3272,N_1185,N_2421);
nor U3273 (N_3273,N_1981,N_1599);
nand U3274 (N_3274,N_1964,N_2117);
nor U3275 (N_3275,N_377,N_18);
or U3276 (N_3276,N_2061,N_67);
or U3277 (N_3277,N_2450,N_1870);
xor U3278 (N_3278,N_138,N_735);
and U3279 (N_3279,N_782,N_1882);
xnor U3280 (N_3280,N_2046,N_1977);
or U3281 (N_3281,N_2032,N_445);
or U3282 (N_3282,N_899,N_742);
and U3283 (N_3283,N_780,N_862);
and U3284 (N_3284,N_563,N_1522);
nand U3285 (N_3285,N_1947,N_1518);
or U3286 (N_3286,N_1473,N_91);
nor U3287 (N_3287,N_788,N_1539);
or U3288 (N_3288,N_651,N_787);
or U3289 (N_3289,N_2152,N_81);
xnor U3290 (N_3290,N_2086,N_2217);
nor U3291 (N_3291,N_2221,N_526);
nand U3292 (N_3292,N_770,N_1659);
and U3293 (N_3293,N_2431,N_2010);
nor U3294 (N_3294,N_61,N_438);
nor U3295 (N_3295,N_903,N_2100);
and U3296 (N_3296,N_464,N_303);
and U3297 (N_3297,N_859,N_1852);
nor U3298 (N_3298,N_266,N_1754);
xnor U3299 (N_3299,N_1054,N_1971);
and U3300 (N_3300,N_265,N_1015);
or U3301 (N_3301,N_2022,N_1521);
and U3302 (N_3302,N_282,N_95);
nor U3303 (N_3303,N_0,N_2305);
xnor U3304 (N_3304,N_2428,N_504);
and U3305 (N_3305,N_1592,N_245);
xnor U3306 (N_3306,N_1611,N_1239);
nor U3307 (N_3307,N_624,N_2071);
nand U3308 (N_3308,N_910,N_1214);
nor U3309 (N_3309,N_2231,N_1308);
nor U3310 (N_3310,N_2429,N_1707);
and U3311 (N_3311,N_1446,N_43);
and U3312 (N_3312,N_691,N_1569);
xnor U3313 (N_3313,N_1845,N_2324);
xor U3314 (N_3314,N_2027,N_2470);
xor U3315 (N_3315,N_1078,N_1892);
and U3316 (N_3316,N_737,N_2388);
and U3317 (N_3317,N_1417,N_1692);
xor U3318 (N_3318,N_400,N_1016);
and U3319 (N_3319,N_2258,N_1951);
nand U3320 (N_3320,N_1302,N_573);
nor U3321 (N_3321,N_1557,N_1706);
nand U3322 (N_3322,N_1002,N_397);
xor U3323 (N_3323,N_269,N_2182);
or U3324 (N_3324,N_1559,N_177);
and U3325 (N_3325,N_922,N_2435);
xnor U3326 (N_3326,N_132,N_1959);
xor U3327 (N_3327,N_680,N_1481);
and U3328 (N_3328,N_399,N_27);
xor U3329 (N_3329,N_1999,N_85);
xnor U3330 (N_3330,N_2188,N_1582);
nor U3331 (N_3331,N_865,N_1620);
and U3332 (N_3332,N_2139,N_1724);
xnor U3333 (N_3333,N_609,N_1624);
xnor U3334 (N_3334,N_458,N_1268);
xor U3335 (N_3335,N_1210,N_1207);
nand U3336 (N_3336,N_374,N_670);
or U3337 (N_3337,N_1510,N_1250);
or U3338 (N_3338,N_407,N_26);
xor U3339 (N_3339,N_2219,N_1195);
nor U3340 (N_3340,N_410,N_75);
nand U3341 (N_3341,N_114,N_1088);
nor U3342 (N_3342,N_19,N_1684);
or U3343 (N_3343,N_1558,N_1628);
or U3344 (N_3344,N_297,N_1289);
or U3345 (N_3345,N_2274,N_786);
and U3346 (N_3346,N_1083,N_1404);
or U3347 (N_3347,N_872,N_685);
nand U3348 (N_3348,N_2272,N_827);
nand U3349 (N_3349,N_5,N_1490);
or U3350 (N_3350,N_1039,N_854);
xor U3351 (N_3351,N_1991,N_1626);
nor U3352 (N_3352,N_1786,N_2089);
nand U3353 (N_3353,N_1877,N_2237);
nand U3354 (N_3354,N_148,N_2114);
nand U3355 (N_3355,N_840,N_1985);
and U3356 (N_3356,N_801,N_2162);
xor U3357 (N_3357,N_1969,N_1590);
nor U3358 (N_3358,N_1336,N_692);
or U3359 (N_3359,N_1738,N_689);
or U3360 (N_3360,N_1254,N_2497);
nand U3361 (N_3361,N_2362,N_2326);
and U3362 (N_3362,N_1651,N_2403);
xor U3363 (N_3363,N_1143,N_1390);
nand U3364 (N_3364,N_2400,N_1211);
nor U3365 (N_3365,N_34,N_388);
xnor U3366 (N_3366,N_985,N_1925);
and U3367 (N_3367,N_120,N_1560);
nand U3368 (N_3368,N_535,N_979);
and U3369 (N_3369,N_1596,N_1486);
nand U3370 (N_3370,N_617,N_2130);
nor U3371 (N_3371,N_794,N_723);
nand U3372 (N_3372,N_577,N_734);
xnor U3373 (N_3373,N_1538,N_1103);
and U3374 (N_3374,N_1963,N_352);
nand U3375 (N_3375,N_2268,N_2332);
or U3376 (N_3376,N_2239,N_1086);
xor U3377 (N_3377,N_1162,N_1622);
or U3378 (N_3378,N_1765,N_1141);
xnor U3379 (N_3379,N_1685,N_2376);
and U3380 (N_3380,N_508,N_1098);
xor U3381 (N_3381,N_2016,N_1919);
nand U3382 (N_3382,N_1735,N_636);
nor U3383 (N_3383,N_187,N_2387);
xor U3384 (N_3384,N_1645,N_2415);
nand U3385 (N_3385,N_2159,N_1824);
nor U3386 (N_3386,N_930,N_320);
xor U3387 (N_3387,N_116,N_2006);
xnor U3388 (N_3388,N_437,N_1733);
nand U3389 (N_3389,N_995,N_16);
nor U3390 (N_3390,N_1508,N_96);
nand U3391 (N_3391,N_2069,N_2058);
nor U3392 (N_3392,N_25,N_122);
and U3393 (N_3393,N_1112,N_1818);
or U3394 (N_3394,N_2150,N_1133);
nand U3395 (N_3395,N_1413,N_1465);
xor U3396 (N_3396,N_1151,N_537);
or U3397 (N_3397,N_1896,N_1013);
xnor U3398 (N_3398,N_1867,N_300);
or U3399 (N_3399,N_2224,N_1632);
xor U3400 (N_3400,N_2420,N_2480);
nor U3401 (N_3401,N_1355,N_378);
xnor U3402 (N_3402,N_964,N_2364);
nand U3403 (N_3403,N_2266,N_32);
or U3404 (N_3404,N_887,N_928);
nor U3405 (N_3405,N_1095,N_176);
or U3406 (N_3406,N_847,N_2371);
xnor U3407 (N_3407,N_2334,N_1696);
and U3408 (N_3408,N_783,N_249);
and U3409 (N_3409,N_436,N_1042);
nand U3410 (N_3410,N_1123,N_1987);
nor U3411 (N_3411,N_94,N_2109);
and U3412 (N_3412,N_179,N_1989);
nor U3413 (N_3413,N_2393,N_2299);
or U3414 (N_3414,N_1258,N_2240);
xor U3415 (N_3415,N_1177,N_2076);
xnor U3416 (N_3416,N_105,N_2474);
nor U3417 (N_3417,N_1920,N_2436);
nor U3418 (N_3418,N_957,N_346);
xor U3419 (N_3419,N_2298,N_293);
xor U3420 (N_3420,N_671,N_1363);
nand U3421 (N_3421,N_452,N_345);
nor U3422 (N_3422,N_218,N_1487);
or U3423 (N_3423,N_1190,N_63);
nand U3424 (N_3424,N_124,N_475);
xnor U3425 (N_3425,N_156,N_960);
or U3426 (N_3426,N_629,N_1096);
nand U3427 (N_3427,N_776,N_184);
or U3428 (N_3428,N_809,N_1348);
nor U3429 (N_3429,N_1748,N_983);
or U3430 (N_3430,N_1403,N_1752);
nand U3431 (N_3431,N_2312,N_2168);
or U3432 (N_3432,N_1472,N_1675);
nor U3433 (N_3433,N_1408,N_72);
and U3434 (N_3434,N_2389,N_589);
xnor U3435 (N_3435,N_975,N_1160);
xnor U3436 (N_3436,N_2325,N_168);
nor U3437 (N_3437,N_1085,N_1256);
xor U3438 (N_3438,N_1036,N_1168);
xnor U3439 (N_3439,N_1034,N_1356);
nand U3440 (N_3440,N_2253,N_549);
or U3441 (N_3441,N_729,N_584);
xnor U3442 (N_3442,N_529,N_764);
xor U3443 (N_3443,N_1480,N_715);
or U3444 (N_3444,N_1697,N_645);
and U3445 (N_3445,N_1020,N_988);
nand U3446 (N_3446,N_646,N_1911);
xnor U3447 (N_3447,N_2433,N_2278);
and U3448 (N_3448,N_1674,N_695);
nand U3449 (N_3449,N_1576,N_2333);
and U3450 (N_3450,N_1761,N_1579);
nor U3451 (N_3451,N_1544,N_1247);
or U3452 (N_3452,N_327,N_1842);
and U3453 (N_3453,N_1813,N_2004);
nor U3454 (N_3454,N_77,N_2381);
and U3455 (N_3455,N_834,N_193);
or U3456 (N_3456,N_2012,N_2005);
nor U3457 (N_3457,N_1442,N_1760);
and U3458 (N_3458,N_1497,N_2481);
xor U3459 (N_3459,N_713,N_1819);
or U3460 (N_3460,N_707,N_100);
nand U3461 (N_3461,N_2244,N_502);
nor U3462 (N_3462,N_2319,N_1552);
nor U3463 (N_3463,N_555,N_71);
and U3464 (N_3464,N_796,N_1284);
and U3465 (N_3465,N_1815,N_1069);
nand U3466 (N_3466,N_1757,N_1204);
or U3467 (N_3467,N_147,N_681);
and U3468 (N_3468,N_2338,N_2259);
or U3469 (N_3469,N_1391,N_2495);
and U3470 (N_3470,N_1700,N_1545);
nor U3471 (N_3471,N_1566,N_154);
xor U3472 (N_3472,N_1001,N_1629);
nand U3473 (N_3473,N_1345,N_2451);
nand U3474 (N_3474,N_1747,N_2477);
xor U3475 (N_3475,N_2356,N_821);
xnor U3476 (N_3476,N_1736,N_172);
nor U3477 (N_3477,N_188,N_1469);
xor U3478 (N_3478,N_1367,N_507);
nand U3479 (N_3479,N_1732,N_832);
and U3480 (N_3480,N_121,N_82);
and U3481 (N_3481,N_233,N_2467);
and U3482 (N_3482,N_1653,N_1125);
xor U3483 (N_3483,N_419,N_2011);
nand U3484 (N_3484,N_2482,N_1407);
or U3485 (N_3485,N_1297,N_1529);
xor U3486 (N_3486,N_1533,N_38);
nand U3487 (N_3487,N_220,N_511);
nor U3488 (N_3488,N_880,N_659);
or U3489 (N_3489,N_1046,N_353);
xor U3490 (N_3490,N_606,N_3);
nand U3491 (N_3491,N_2151,N_2218);
nand U3492 (N_3492,N_1988,N_562);
xor U3493 (N_3493,N_1937,N_2183);
xor U3494 (N_3494,N_768,N_1222);
or U3495 (N_3495,N_283,N_2099);
xnor U3496 (N_3496,N_924,N_2107);
nor U3497 (N_3497,N_2143,N_694);
nor U3498 (N_3498,N_2082,N_186);
and U3499 (N_3499,N_1290,N_1721);
nor U3500 (N_3500,N_1251,N_1238);
or U3501 (N_3501,N_959,N_881);
nor U3502 (N_3502,N_596,N_2148);
xnor U3503 (N_3503,N_1749,N_423);
xnor U3504 (N_3504,N_2246,N_272);
xnor U3505 (N_3505,N_1430,N_485);
nand U3506 (N_3506,N_747,N_533);
nand U3507 (N_3507,N_483,N_92);
or U3508 (N_3508,N_359,N_1910);
nor U3509 (N_3509,N_1839,N_1484);
nand U3510 (N_3510,N_1860,N_482);
and U3511 (N_3511,N_372,N_1161);
and U3512 (N_3512,N_644,N_2175);
and U3513 (N_3513,N_1492,N_1537);
nand U3514 (N_3514,N_57,N_2247);
nand U3515 (N_3515,N_130,N_173);
and U3516 (N_3516,N_726,N_2252);
xor U3517 (N_3517,N_335,N_481);
nor U3518 (N_3518,N_1703,N_774);
nand U3519 (N_3519,N_2443,N_797);
and U3520 (N_3520,N_920,N_1972);
nand U3521 (N_3521,N_1217,N_1740);
nand U3522 (N_3522,N_1120,N_2396);
xor U3523 (N_3523,N_2234,N_2019);
xor U3524 (N_3524,N_208,N_824);
xnor U3525 (N_3525,N_510,N_328);
nor U3526 (N_3526,N_2419,N_2463);
and U3527 (N_3527,N_2044,N_180);
xnor U3528 (N_3528,N_2098,N_365);
and U3529 (N_3529,N_1918,N_2304);
xnor U3530 (N_3530,N_139,N_1326);
nor U3531 (N_3531,N_1676,N_248);
and U3532 (N_3532,N_544,N_1823);
or U3533 (N_3533,N_1994,N_603);
xor U3534 (N_3534,N_1170,N_289);
or U3535 (N_3535,N_1351,N_1938);
and U3536 (N_3536,N_944,N_242);
xnor U3537 (N_3537,N_2023,N_607);
or U3538 (N_3538,N_1077,N_1955);
nand U3539 (N_3539,N_2275,N_1428);
nand U3540 (N_3540,N_2366,N_2077);
and U3541 (N_3541,N_1477,N_628);
nand U3542 (N_3542,N_615,N_760);
nand U3543 (N_3543,N_1642,N_1138);
or U3544 (N_3544,N_2216,N_1869);
and U3545 (N_3545,N_1330,N_996);
nor U3546 (N_3546,N_446,N_843);
xnor U3547 (N_3547,N_781,N_237);
or U3548 (N_3548,N_2212,N_972);
nor U3549 (N_3549,N_2078,N_683);
and U3550 (N_3550,N_227,N_316);
or U3551 (N_3551,N_492,N_1226);
xnor U3552 (N_3552,N_1950,N_839);
nor U3553 (N_3553,N_1052,N_103);
nand U3554 (N_3554,N_1750,N_2142);
or U3555 (N_3555,N_1152,N_875);
and U3556 (N_3556,N_392,N_478);
nand U3557 (N_3557,N_1634,N_2220);
or U3558 (N_3558,N_618,N_1779);
or U3559 (N_3559,N_1319,N_333);
nor U3560 (N_3560,N_1979,N_1897);
and U3561 (N_3561,N_110,N_2229);
nand U3562 (N_3562,N_1519,N_2472);
and U3563 (N_3563,N_1574,N_255);
or U3564 (N_3564,N_1705,N_1952);
and U3565 (N_3565,N_690,N_1163);
nand U3566 (N_3566,N_131,N_2008);
xnor U3567 (N_3567,N_718,N_2365);
and U3568 (N_3568,N_468,N_989);
and U3569 (N_3569,N_756,N_118);
nor U3570 (N_3570,N_1269,N_2242);
nor U3571 (N_3571,N_1344,N_1549);
and U3572 (N_3572,N_224,N_528);
nand U3573 (N_3573,N_1276,N_425);
and U3574 (N_3574,N_1719,N_469);
and U3575 (N_3575,N_259,N_1317);
nor U3576 (N_3576,N_1798,N_2122);
xnor U3577 (N_3577,N_2056,N_2161);
xnor U3578 (N_3578,N_279,N_331);
nand U3579 (N_3579,N_165,N_273);
or U3580 (N_3580,N_288,N_673);
and U3581 (N_3581,N_738,N_1382);
xnor U3582 (N_3582,N_2222,N_1758);
nand U3583 (N_3583,N_97,N_1714);
xnor U3584 (N_3584,N_465,N_1801);
nor U3585 (N_3585,N_113,N_505);
and U3586 (N_3586,N_1759,N_546);
nand U3587 (N_3587,N_955,N_170);
nand U3588 (N_3588,N_873,N_1097);
xor U3589 (N_3589,N_1639,N_1961);
or U3590 (N_3590,N_443,N_1677);
or U3591 (N_3591,N_480,N_864);
xnor U3592 (N_3592,N_6,N_1804);
and U3593 (N_3593,N_1295,N_1038);
xor U3594 (N_3594,N_567,N_2174);
nor U3595 (N_3595,N_2479,N_158);
nor U3596 (N_3596,N_339,N_1260);
or U3597 (N_3597,N_380,N_1072);
nor U3598 (N_3598,N_1766,N_2003);
and U3599 (N_3599,N_2367,N_1414);
xnor U3600 (N_3600,N_59,N_1535);
nand U3601 (N_3601,N_2287,N_2203);
and U3602 (N_3602,N_541,N_1646);
nor U3603 (N_3603,N_1377,N_2475);
and U3604 (N_3604,N_894,N_479);
nor U3605 (N_3605,N_1478,N_1375);
or U3606 (N_3606,N_1888,N_853);
nor U3607 (N_3607,N_1827,N_1441);
nand U3608 (N_3608,N_953,N_773);
and U3609 (N_3609,N_1844,N_2465);
nand U3610 (N_3610,N_2459,N_2473);
or U3611 (N_3611,N_418,N_477);
xnor U3612 (N_3612,N_817,N_2273);
nand U3613 (N_3613,N_652,N_2215);
or U3614 (N_3614,N_1349,N_1274);
nor U3615 (N_3615,N_1742,N_1135);
or U3616 (N_3616,N_42,N_427);
xnor U3617 (N_3617,N_2001,N_1468);
nand U3618 (N_3618,N_1935,N_99);
or U3619 (N_3619,N_13,N_697);
xor U3620 (N_3620,N_268,N_344);
or U3621 (N_3621,N_605,N_309);
or U3622 (N_3622,N_1333,N_1432);
nand U3623 (N_3623,N_1781,N_73);
nor U3624 (N_3624,N_2134,N_244);
nor U3625 (N_3625,N_593,N_88);
and U3626 (N_3626,N_2310,N_1848);
and U3627 (N_3627,N_2491,N_1236);
nand U3628 (N_3628,N_993,N_2318);
xnor U3629 (N_3629,N_119,N_1588);
nor U3630 (N_3630,N_323,N_434);
xor U3631 (N_3631,N_127,N_2424);
nand U3632 (N_3632,N_317,N_1191);
nand U3633 (N_3633,N_1570,N_200);
xnor U3634 (N_3634,N_621,N_1806);
and U3635 (N_3635,N_777,N_1788);
or U3636 (N_3636,N_54,N_1060);
xor U3637 (N_3637,N_286,N_2297);
nand U3638 (N_3638,N_1128,N_1505);
or U3639 (N_3639,N_1139,N_950);
nand U3640 (N_3640,N_2026,N_938);
and U3641 (N_3641,N_2199,N_1810);
xor U3642 (N_3642,N_2358,N_2033);
nand U3643 (N_3643,N_626,N_1026);
xor U3644 (N_3644,N_1454,N_623);
xnor U3645 (N_3645,N_1751,N_2068);
and U3646 (N_3646,N_2038,N_837);
or U3647 (N_3647,N_2043,N_1511);
or U3648 (N_3648,N_2040,N_531);
nor U3649 (N_3649,N_2309,N_1553);
xnor U3650 (N_3650,N_1009,N_1371);
xnor U3651 (N_3651,N_1717,N_1661);
nor U3652 (N_3652,N_798,N_1655);
nor U3653 (N_3653,N_897,N_1116);
nand U3654 (N_3654,N_1316,N_1113);
nand U3655 (N_3655,N_2496,N_578);
nor U3656 (N_3656,N_325,N_393);
or U3657 (N_3657,N_1358,N_236);
and U3658 (N_3658,N_232,N_307);
nand U3659 (N_3659,N_2052,N_396);
nand U3660 (N_3660,N_1171,N_299);
xor U3661 (N_3661,N_658,N_306);
or U3662 (N_3662,N_1339,N_129);
nor U3663 (N_3663,N_2163,N_1224);
xnor U3664 (N_3664,N_2426,N_1252);
xor U3665 (N_3665,N_2173,N_919);
nor U3666 (N_3666,N_350,N_949);
xor U3667 (N_3667,N_267,N_1047);
nor U3668 (N_3668,N_807,N_1966);
and U3669 (N_3669,N_1784,N_1525);
and U3670 (N_3670,N_1438,N_1080);
nor U3671 (N_3671,N_495,N_2369);
nand U3672 (N_3672,N_2105,N_433);
and U3673 (N_3673,N_1041,N_2147);
nand U3674 (N_3674,N_1322,N_2418);
xnor U3675 (N_3675,N_2,N_2102);
nand U3676 (N_3676,N_2286,N_1690);
nor U3677 (N_3677,N_820,N_778);
xor U3678 (N_3678,N_370,N_941);
nor U3679 (N_3679,N_1084,N_2196);
or U3680 (N_3680,N_2035,N_610);
and U3681 (N_3681,N_1769,N_2166);
xnor U3682 (N_3682,N_1960,N_1577);
nor U3683 (N_3683,N_1608,N_527);
xor U3684 (N_3684,N_838,N_1876);
or U3685 (N_3685,N_1089,N_415);
and U3686 (N_3686,N_514,N_1669);
nand U3687 (N_3687,N_1872,N_2205);
or U3688 (N_3688,N_1573,N_2368);
and U3689 (N_3689,N_643,N_66);
or U3690 (N_3690,N_2406,N_799);
or U3691 (N_3691,N_1728,N_2427);
or U3692 (N_3692,N_491,N_1900);
and U3693 (N_3693,N_1479,N_522);
or U3694 (N_3694,N_211,N_1933);
or U3695 (N_3695,N_908,N_1342);
xor U3696 (N_3696,N_2126,N_1203);
xnor U3697 (N_3697,N_1429,N_2057);
nor U3698 (N_3698,N_557,N_800);
xor U3699 (N_3699,N_1483,N_1388);
or U3700 (N_3700,N_108,N_2194);
xor U3701 (N_3701,N_1184,N_1595);
nand U3702 (N_3702,N_76,N_1805);
nor U3703 (N_3703,N_1601,N_856);
and U3704 (N_3704,N_714,N_340);
xor U3705 (N_3705,N_1314,N_761);
and U3706 (N_3706,N_1262,N_810);
or U3707 (N_3707,N_1923,N_1793);
xnor U3708 (N_3708,N_2262,N_1270);
or U3709 (N_3709,N_2020,N_1021);
xor U3710 (N_3710,N_512,N_1245);
nand U3711 (N_3711,N_2177,N_1451);
or U3712 (N_3712,N_311,N_2394);
and U3713 (N_3713,N_1647,N_1613);
and U3714 (N_3714,N_143,N_849);
nand U3715 (N_3715,N_294,N_2101);
and U3716 (N_3716,N_1127,N_884);
or U3717 (N_3717,N_763,N_462);
nor U3718 (N_3718,N_969,N_1090);
and U3719 (N_3719,N_2017,N_1555);
or U3720 (N_3720,N_1619,N_1514);
or U3721 (N_3721,N_109,N_1229);
nor U3722 (N_3722,N_785,N_2291);
and U3723 (N_3723,N_144,N_896);
xnor U3724 (N_3724,N_804,N_210);
xnor U3725 (N_3725,N_946,N_358);
or U3726 (N_3726,N_1790,N_698);
nand U3727 (N_3727,N_1984,N_2145);
nand U3728 (N_3728,N_836,N_2051);
xnor U3729 (N_3729,N_382,N_1281);
and U3730 (N_3730,N_1667,N_1107);
nor U3731 (N_3731,N_1580,N_1809);
xnor U3732 (N_3732,N_463,N_35);
or U3733 (N_3733,N_195,N_1005);
nor U3734 (N_3734,N_2295,N_215);
nand U3735 (N_3735,N_39,N_310);
nor U3736 (N_3736,N_246,N_2104);
xnor U3737 (N_3737,N_1916,N_367);
nand U3738 (N_3738,N_175,N_858);
nand U3739 (N_3739,N_1932,N_486);
xnor U3740 (N_3740,N_909,N_1885);
xor U3741 (N_3741,N_321,N_1215);
xnor U3742 (N_3742,N_1018,N_1945);
or U3743 (N_3743,N_597,N_2492);
nand U3744 (N_3744,N_1216,N_1551);
and U3745 (N_3745,N_650,N_1110);
nor U3746 (N_3746,N_2378,N_342);
nor U3747 (N_3747,N_1630,N_1273);
xor U3748 (N_3748,N_2157,N_424);
nor U3749 (N_3749,N_1627,N_1725);
or U3750 (N_3750,N_2132,N_1705);
and U3751 (N_3751,N_296,N_444);
nor U3752 (N_3752,N_1629,N_1184);
and U3753 (N_3753,N_1799,N_597);
xnor U3754 (N_3754,N_2375,N_2096);
or U3755 (N_3755,N_2430,N_2124);
or U3756 (N_3756,N_108,N_1201);
xor U3757 (N_3757,N_579,N_472);
nor U3758 (N_3758,N_118,N_2064);
nor U3759 (N_3759,N_743,N_1694);
and U3760 (N_3760,N_2425,N_1087);
nand U3761 (N_3761,N_2057,N_1094);
or U3762 (N_3762,N_699,N_307);
nor U3763 (N_3763,N_139,N_729);
xor U3764 (N_3764,N_656,N_79);
nand U3765 (N_3765,N_2468,N_211);
or U3766 (N_3766,N_2077,N_2047);
nor U3767 (N_3767,N_325,N_1952);
nand U3768 (N_3768,N_17,N_361);
or U3769 (N_3769,N_923,N_1036);
and U3770 (N_3770,N_1553,N_2400);
nand U3771 (N_3771,N_1155,N_1534);
xor U3772 (N_3772,N_460,N_566);
xnor U3773 (N_3773,N_107,N_1945);
xnor U3774 (N_3774,N_1411,N_2404);
nand U3775 (N_3775,N_863,N_32);
xnor U3776 (N_3776,N_935,N_1259);
nand U3777 (N_3777,N_388,N_2413);
or U3778 (N_3778,N_29,N_2200);
nand U3779 (N_3779,N_1540,N_1818);
and U3780 (N_3780,N_2349,N_1983);
xnor U3781 (N_3781,N_608,N_755);
or U3782 (N_3782,N_1546,N_996);
nor U3783 (N_3783,N_758,N_1125);
or U3784 (N_3784,N_1692,N_2340);
and U3785 (N_3785,N_470,N_1643);
nor U3786 (N_3786,N_1634,N_659);
nand U3787 (N_3787,N_2479,N_2030);
and U3788 (N_3788,N_2168,N_1580);
or U3789 (N_3789,N_2331,N_802);
nor U3790 (N_3790,N_722,N_1141);
xnor U3791 (N_3791,N_637,N_147);
nor U3792 (N_3792,N_601,N_2198);
or U3793 (N_3793,N_226,N_871);
nor U3794 (N_3794,N_220,N_1587);
nor U3795 (N_3795,N_1105,N_1258);
or U3796 (N_3796,N_186,N_364);
xnor U3797 (N_3797,N_634,N_917);
xor U3798 (N_3798,N_1962,N_1185);
nand U3799 (N_3799,N_1395,N_276);
nand U3800 (N_3800,N_1717,N_1956);
nor U3801 (N_3801,N_1250,N_934);
or U3802 (N_3802,N_1898,N_922);
and U3803 (N_3803,N_2013,N_1221);
or U3804 (N_3804,N_344,N_2019);
and U3805 (N_3805,N_1041,N_1628);
xnor U3806 (N_3806,N_1924,N_1756);
and U3807 (N_3807,N_32,N_1730);
and U3808 (N_3808,N_2143,N_979);
or U3809 (N_3809,N_1424,N_523);
and U3810 (N_3810,N_1764,N_2465);
nor U3811 (N_3811,N_1517,N_882);
nand U3812 (N_3812,N_256,N_123);
nand U3813 (N_3813,N_111,N_1723);
nor U3814 (N_3814,N_1059,N_1657);
and U3815 (N_3815,N_7,N_1952);
nor U3816 (N_3816,N_548,N_1062);
and U3817 (N_3817,N_31,N_461);
nand U3818 (N_3818,N_2296,N_242);
nand U3819 (N_3819,N_16,N_865);
or U3820 (N_3820,N_1795,N_30);
and U3821 (N_3821,N_1993,N_1567);
or U3822 (N_3822,N_777,N_1387);
xor U3823 (N_3823,N_660,N_1444);
or U3824 (N_3824,N_1692,N_940);
nand U3825 (N_3825,N_2437,N_2495);
and U3826 (N_3826,N_2410,N_1337);
nor U3827 (N_3827,N_129,N_1871);
xor U3828 (N_3828,N_697,N_2305);
xor U3829 (N_3829,N_1738,N_1961);
nand U3830 (N_3830,N_2067,N_2145);
or U3831 (N_3831,N_702,N_1701);
nand U3832 (N_3832,N_2040,N_1945);
nor U3833 (N_3833,N_834,N_984);
and U3834 (N_3834,N_1036,N_395);
nor U3835 (N_3835,N_1062,N_281);
nor U3836 (N_3836,N_1995,N_734);
nor U3837 (N_3837,N_1936,N_186);
and U3838 (N_3838,N_2034,N_199);
xnor U3839 (N_3839,N_1237,N_314);
nand U3840 (N_3840,N_1464,N_1439);
nor U3841 (N_3841,N_682,N_1290);
nor U3842 (N_3842,N_2057,N_2471);
and U3843 (N_3843,N_1468,N_202);
or U3844 (N_3844,N_17,N_1252);
or U3845 (N_3845,N_203,N_2447);
nor U3846 (N_3846,N_2391,N_226);
nand U3847 (N_3847,N_1990,N_2138);
nor U3848 (N_3848,N_1105,N_1482);
or U3849 (N_3849,N_1462,N_734);
or U3850 (N_3850,N_2040,N_338);
nor U3851 (N_3851,N_569,N_73);
nor U3852 (N_3852,N_2284,N_719);
or U3853 (N_3853,N_1155,N_397);
xnor U3854 (N_3854,N_1531,N_1053);
nor U3855 (N_3855,N_693,N_1724);
nor U3856 (N_3856,N_369,N_1001);
nor U3857 (N_3857,N_1497,N_2049);
or U3858 (N_3858,N_2078,N_880);
xor U3859 (N_3859,N_1260,N_948);
nor U3860 (N_3860,N_737,N_2414);
nor U3861 (N_3861,N_1050,N_986);
xor U3862 (N_3862,N_606,N_372);
nor U3863 (N_3863,N_1521,N_1734);
xnor U3864 (N_3864,N_1322,N_2118);
or U3865 (N_3865,N_1127,N_32);
and U3866 (N_3866,N_147,N_1);
xnor U3867 (N_3867,N_1174,N_1268);
nand U3868 (N_3868,N_829,N_2159);
and U3869 (N_3869,N_1614,N_2006);
nand U3870 (N_3870,N_119,N_1186);
nand U3871 (N_3871,N_542,N_2001);
xnor U3872 (N_3872,N_1395,N_227);
xnor U3873 (N_3873,N_1144,N_539);
nor U3874 (N_3874,N_1733,N_1594);
and U3875 (N_3875,N_2318,N_1665);
and U3876 (N_3876,N_699,N_102);
xnor U3877 (N_3877,N_261,N_275);
xor U3878 (N_3878,N_2126,N_1815);
nand U3879 (N_3879,N_382,N_1029);
xor U3880 (N_3880,N_1894,N_454);
or U3881 (N_3881,N_1241,N_1331);
xnor U3882 (N_3882,N_1720,N_1648);
or U3883 (N_3883,N_15,N_1451);
nand U3884 (N_3884,N_437,N_1611);
xor U3885 (N_3885,N_263,N_2204);
and U3886 (N_3886,N_204,N_1154);
nand U3887 (N_3887,N_1335,N_292);
nand U3888 (N_3888,N_842,N_649);
and U3889 (N_3889,N_447,N_58);
nand U3890 (N_3890,N_1969,N_425);
xor U3891 (N_3891,N_1540,N_1950);
xor U3892 (N_3892,N_812,N_250);
and U3893 (N_3893,N_1750,N_2019);
nand U3894 (N_3894,N_1135,N_2202);
xor U3895 (N_3895,N_222,N_254);
nand U3896 (N_3896,N_1081,N_2460);
nand U3897 (N_3897,N_610,N_959);
or U3898 (N_3898,N_1469,N_1179);
xor U3899 (N_3899,N_1264,N_2377);
nand U3900 (N_3900,N_2268,N_2045);
xnor U3901 (N_3901,N_1511,N_777);
nand U3902 (N_3902,N_1830,N_2438);
nor U3903 (N_3903,N_109,N_1392);
or U3904 (N_3904,N_1373,N_1271);
xor U3905 (N_3905,N_373,N_2003);
nor U3906 (N_3906,N_2151,N_1034);
or U3907 (N_3907,N_1538,N_1695);
xor U3908 (N_3908,N_1580,N_558);
nand U3909 (N_3909,N_470,N_2339);
xnor U3910 (N_3910,N_175,N_954);
xor U3911 (N_3911,N_1599,N_982);
or U3912 (N_3912,N_1968,N_892);
nand U3913 (N_3913,N_2373,N_807);
xnor U3914 (N_3914,N_1355,N_448);
or U3915 (N_3915,N_2257,N_1171);
and U3916 (N_3916,N_346,N_1017);
nor U3917 (N_3917,N_684,N_2302);
nand U3918 (N_3918,N_2162,N_1929);
and U3919 (N_3919,N_2060,N_798);
nor U3920 (N_3920,N_2321,N_1056);
and U3921 (N_3921,N_1938,N_120);
or U3922 (N_3922,N_899,N_2207);
nand U3923 (N_3923,N_1898,N_1673);
xnor U3924 (N_3924,N_265,N_482);
xor U3925 (N_3925,N_855,N_2050);
xor U3926 (N_3926,N_326,N_1953);
or U3927 (N_3927,N_1143,N_338);
nand U3928 (N_3928,N_1597,N_403);
or U3929 (N_3929,N_1340,N_1933);
and U3930 (N_3930,N_1808,N_1545);
nor U3931 (N_3931,N_2048,N_243);
nor U3932 (N_3932,N_484,N_649);
nand U3933 (N_3933,N_1320,N_1778);
or U3934 (N_3934,N_1032,N_1188);
nor U3935 (N_3935,N_747,N_716);
xor U3936 (N_3936,N_407,N_625);
nor U3937 (N_3937,N_1784,N_810);
and U3938 (N_3938,N_541,N_2002);
and U3939 (N_3939,N_1505,N_889);
or U3940 (N_3940,N_603,N_441);
nor U3941 (N_3941,N_1837,N_915);
or U3942 (N_3942,N_1110,N_268);
or U3943 (N_3943,N_2231,N_354);
xor U3944 (N_3944,N_487,N_1923);
nand U3945 (N_3945,N_2220,N_1398);
or U3946 (N_3946,N_1368,N_1711);
and U3947 (N_3947,N_1505,N_1848);
and U3948 (N_3948,N_221,N_1213);
and U3949 (N_3949,N_2060,N_1965);
or U3950 (N_3950,N_2427,N_2377);
and U3951 (N_3951,N_1112,N_87);
or U3952 (N_3952,N_2155,N_1422);
xor U3953 (N_3953,N_1435,N_1698);
xor U3954 (N_3954,N_1870,N_1562);
nor U3955 (N_3955,N_333,N_2141);
nor U3956 (N_3956,N_1637,N_1160);
nor U3957 (N_3957,N_880,N_954);
nor U3958 (N_3958,N_2230,N_1720);
xor U3959 (N_3959,N_1365,N_2470);
xnor U3960 (N_3960,N_1759,N_757);
and U3961 (N_3961,N_2164,N_2136);
and U3962 (N_3962,N_2421,N_1963);
or U3963 (N_3963,N_32,N_1883);
and U3964 (N_3964,N_1389,N_22);
nand U3965 (N_3965,N_1485,N_149);
nor U3966 (N_3966,N_1710,N_1882);
nand U3967 (N_3967,N_873,N_1837);
nand U3968 (N_3968,N_49,N_734);
nor U3969 (N_3969,N_154,N_1901);
or U3970 (N_3970,N_1153,N_1592);
and U3971 (N_3971,N_1506,N_27);
nor U3972 (N_3972,N_2155,N_1131);
and U3973 (N_3973,N_2158,N_2426);
xnor U3974 (N_3974,N_409,N_626);
nor U3975 (N_3975,N_782,N_894);
nor U3976 (N_3976,N_862,N_1535);
xor U3977 (N_3977,N_171,N_1668);
or U3978 (N_3978,N_1253,N_1913);
nand U3979 (N_3979,N_2055,N_676);
xnor U3980 (N_3980,N_464,N_863);
xnor U3981 (N_3981,N_832,N_635);
and U3982 (N_3982,N_1824,N_801);
nor U3983 (N_3983,N_2235,N_2080);
xnor U3984 (N_3984,N_1532,N_2107);
and U3985 (N_3985,N_2161,N_1742);
xor U3986 (N_3986,N_144,N_1949);
and U3987 (N_3987,N_2378,N_1131);
nand U3988 (N_3988,N_2266,N_627);
and U3989 (N_3989,N_578,N_237);
xnor U3990 (N_3990,N_2236,N_608);
or U3991 (N_3991,N_235,N_1665);
nor U3992 (N_3992,N_2040,N_2237);
nand U3993 (N_3993,N_786,N_48);
or U3994 (N_3994,N_2149,N_912);
nor U3995 (N_3995,N_314,N_995);
nand U3996 (N_3996,N_541,N_1520);
and U3997 (N_3997,N_960,N_1515);
nand U3998 (N_3998,N_1775,N_1475);
or U3999 (N_3999,N_2019,N_2295);
and U4000 (N_4000,N_1503,N_591);
or U4001 (N_4001,N_2186,N_384);
and U4002 (N_4002,N_277,N_416);
xor U4003 (N_4003,N_2360,N_5);
and U4004 (N_4004,N_1037,N_1000);
and U4005 (N_4005,N_760,N_780);
nor U4006 (N_4006,N_1912,N_2380);
nand U4007 (N_4007,N_1183,N_951);
nor U4008 (N_4008,N_1331,N_682);
xnor U4009 (N_4009,N_307,N_1234);
nor U4010 (N_4010,N_1727,N_953);
or U4011 (N_4011,N_2074,N_160);
or U4012 (N_4012,N_1405,N_1933);
nand U4013 (N_4013,N_330,N_1791);
xnor U4014 (N_4014,N_1601,N_2037);
xnor U4015 (N_4015,N_691,N_2137);
nand U4016 (N_4016,N_581,N_1983);
nand U4017 (N_4017,N_1525,N_199);
and U4018 (N_4018,N_2160,N_476);
nand U4019 (N_4019,N_1452,N_2113);
nand U4020 (N_4020,N_2467,N_2006);
or U4021 (N_4021,N_411,N_1455);
xor U4022 (N_4022,N_1291,N_1503);
or U4023 (N_4023,N_1145,N_1093);
or U4024 (N_4024,N_1503,N_2474);
xnor U4025 (N_4025,N_2273,N_1301);
or U4026 (N_4026,N_572,N_2460);
nand U4027 (N_4027,N_1360,N_1963);
nand U4028 (N_4028,N_614,N_2120);
nor U4029 (N_4029,N_338,N_1424);
nor U4030 (N_4030,N_1977,N_2396);
and U4031 (N_4031,N_2371,N_1964);
or U4032 (N_4032,N_2260,N_682);
and U4033 (N_4033,N_780,N_1252);
xnor U4034 (N_4034,N_966,N_1214);
nor U4035 (N_4035,N_2324,N_2445);
nor U4036 (N_4036,N_821,N_1040);
and U4037 (N_4037,N_1744,N_1264);
and U4038 (N_4038,N_1847,N_1628);
and U4039 (N_4039,N_1047,N_1537);
and U4040 (N_4040,N_5,N_480);
nor U4041 (N_4041,N_413,N_2);
xnor U4042 (N_4042,N_1718,N_1260);
or U4043 (N_4043,N_1563,N_1962);
and U4044 (N_4044,N_614,N_1139);
or U4045 (N_4045,N_145,N_612);
nand U4046 (N_4046,N_2051,N_462);
or U4047 (N_4047,N_339,N_2281);
and U4048 (N_4048,N_2000,N_1562);
nand U4049 (N_4049,N_225,N_1238);
nor U4050 (N_4050,N_1636,N_1071);
or U4051 (N_4051,N_2016,N_1041);
xor U4052 (N_4052,N_1210,N_333);
nor U4053 (N_4053,N_2272,N_2168);
nand U4054 (N_4054,N_1322,N_294);
and U4055 (N_4055,N_380,N_976);
xnor U4056 (N_4056,N_434,N_80);
or U4057 (N_4057,N_361,N_936);
nor U4058 (N_4058,N_1124,N_295);
nand U4059 (N_4059,N_1085,N_481);
or U4060 (N_4060,N_1128,N_792);
nand U4061 (N_4061,N_505,N_1794);
nor U4062 (N_4062,N_2323,N_1615);
or U4063 (N_4063,N_886,N_727);
nor U4064 (N_4064,N_1845,N_1839);
nor U4065 (N_4065,N_219,N_279);
and U4066 (N_4066,N_2017,N_1390);
or U4067 (N_4067,N_1212,N_1055);
and U4068 (N_4068,N_1252,N_2422);
or U4069 (N_4069,N_704,N_1325);
nand U4070 (N_4070,N_1245,N_1667);
nand U4071 (N_4071,N_1661,N_2172);
xnor U4072 (N_4072,N_2310,N_1048);
xnor U4073 (N_4073,N_1464,N_1733);
and U4074 (N_4074,N_822,N_2409);
xnor U4075 (N_4075,N_2174,N_2433);
nor U4076 (N_4076,N_323,N_780);
and U4077 (N_4077,N_1674,N_2262);
and U4078 (N_4078,N_478,N_2493);
or U4079 (N_4079,N_1168,N_1161);
nand U4080 (N_4080,N_817,N_656);
or U4081 (N_4081,N_883,N_1709);
nand U4082 (N_4082,N_925,N_2094);
nor U4083 (N_4083,N_466,N_1979);
xor U4084 (N_4084,N_2035,N_719);
and U4085 (N_4085,N_67,N_2303);
or U4086 (N_4086,N_954,N_1120);
nand U4087 (N_4087,N_6,N_671);
nand U4088 (N_4088,N_110,N_1125);
nor U4089 (N_4089,N_946,N_1093);
xnor U4090 (N_4090,N_2465,N_1690);
xor U4091 (N_4091,N_1664,N_1229);
nand U4092 (N_4092,N_522,N_1188);
xor U4093 (N_4093,N_734,N_721);
nor U4094 (N_4094,N_364,N_2077);
xnor U4095 (N_4095,N_375,N_1327);
nand U4096 (N_4096,N_56,N_86);
or U4097 (N_4097,N_1476,N_1630);
xnor U4098 (N_4098,N_181,N_1613);
and U4099 (N_4099,N_171,N_944);
nor U4100 (N_4100,N_1027,N_763);
or U4101 (N_4101,N_936,N_2096);
nand U4102 (N_4102,N_1871,N_2045);
and U4103 (N_4103,N_2065,N_710);
and U4104 (N_4104,N_563,N_1164);
nor U4105 (N_4105,N_1417,N_2142);
nand U4106 (N_4106,N_1088,N_909);
nor U4107 (N_4107,N_1451,N_1211);
nand U4108 (N_4108,N_2249,N_1299);
and U4109 (N_4109,N_2306,N_2434);
xor U4110 (N_4110,N_21,N_2394);
xnor U4111 (N_4111,N_1776,N_2040);
or U4112 (N_4112,N_982,N_628);
and U4113 (N_4113,N_811,N_1817);
nand U4114 (N_4114,N_224,N_1948);
and U4115 (N_4115,N_1051,N_1901);
xnor U4116 (N_4116,N_1635,N_2402);
nand U4117 (N_4117,N_1551,N_2219);
xnor U4118 (N_4118,N_1906,N_119);
xnor U4119 (N_4119,N_1203,N_512);
nor U4120 (N_4120,N_895,N_718);
and U4121 (N_4121,N_114,N_344);
nor U4122 (N_4122,N_479,N_737);
and U4123 (N_4123,N_1114,N_2293);
nand U4124 (N_4124,N_410,N_429);
xor U4125 (N_4125,N_655,N_1462);
xor U4126 (N_4126,N_521,N_2403);
or U4127 (N_4127,N_539,N_2173);
nand U4128 (N_4128,N_3,N_854);
nor U4129 (N_4129,N_764,N_65);
xor U4130 (N_4130,N_2022,N_992);
xor U4131 (N_4131,N_1615,N_1290);
nand U4132 (N_4132,N_1600,N_2196);
nand U4133 (N_4133,N_462,N_1411);
nor U4134 (N_4134,N_2321,N_396);
and U4135 (N_4135,N_1697,N_1579);
nor U4136 (N_4136,N_1378,N_733);
and U4137 (N_4137,N_2030,N_2095);
nor U4138 (N_4138,N_715,N_2329);
and U4139 (N_4139,N_911,N_1424);
and U4140 (N_4140,N_649,N_2147);
and U4141 (N_4141,N_2071,N_1378);
or U4142 (N_4142,N_187,N_509);
nor U4143 (N_4143,N_528,N_88);
xor U4144 (N_4144,N_1647,N_1080);
or U4145 (N_4145,N_203,N_2091);
xnor U4146 (N_4146,N_858,N_1538);
nand U4147 (N_4147,N_2443,N_2453);
or U4148 (N_4148,N_1219,N_2238);
or U4149 (N_4149,N_54,N_2193);
nor U4150 (N_4150,N_829,N_2307);
xor U4151 (N_4151,N_1037,N_1102);
xor U4152 (N_4152,N_862,N_2267);
or U4153 (N_4153,N_955,N_1441);
and U4154 (N_4154,N_1178,N_503);
xnor U4155 (N_4155,N_1099,N_702);
and U4156 (N_4156,N_1502,N_1914);
nand U4157 (N_4157,N_947,N_1439);
xnor U4158 (N_4158,N_120,N_2203);
and U4159 (N_4159,N_883,N_604);
nor U4160 (N_4160,N_2135,N_401);
xnor U4161 (N_4161,N_599,N_421);
or U4162 (N_4162,N_1376,N_1603);
xnor U4163 (N_4163,N_2173,N_2469);
or U4164 (N_4164,N_198,N_2357);
and U4165 (N_4165,N_656,N_1849);
nand U4166 (N_4166,N_306,N_1822);
or U4167 (N_4167,N_41,N_452);
nand U4168 (N_4168,N_59,N_777);
and U4169 (N_4169,N_1656,N_609);
nand U4170 (N_4170,N_118,N_429);
and U4171 (N_4171,N_341,N_167);
and U4172 (N_4172,N_1967,N_1385);
nor U4173 (N_4173,N_1143,N_2097);
nand U4174 (N_4174,N_603,N_1254);
nor U4175 (N_4175,N_1083,N_1469);
and U4176 (N_4176,N_965,N_1363);
xor U4177 (N_4177,N_2280,N_645);
and U4178 (N_4178,N_962,N_2086);
nand U4179 (N_4179,N_1619,N_421);
nand U4180 (N_4180,N_631,N_143);
and U4181 (N_4181,N_1914,N_2183);
xor U4182 (N_4182,N_720,N_167);
or U4183 (N_4183,N_975,N_2453);
xnor U4184 (N_4184,N_2203,N_1493);
xor U4185 (N_4185,N_134,N_1447);
nand U4186 (N_4186,N_1380,N_1530);
and U4187 (N_4187,N_2357,N_1683);
xor U4188 (N_4188,N_1828,N_1470);
and U4189 (N_4189,N_1299,N_473);
nor U4190 (N_4190,N_1524,N_1637);
and U4191 (N_4191,N_2004,N_2438);
xnor U4192 (N_4192,N_2038,N_644);
nand U4193 (N_4193,N_1437,N_1136);
nand U4194 (N_4194,N_495,N_13);
xor U4195 (N_4195,N_657,N_1203);
nor U4196 (N_4196,N_978,N_333);
nand U4197 (N_4197,N_515,N_990);
nand U4198 (N_4198,N_1146,N_1378);
and U4199 (N_4199,N_300,N_1682);
and U4200 (N_4200,N_2119,N_2498);
or U4201 (N_4201,N_255,N_1146);
and U4202 (N_4202,N_133,N_803);
nand U4203 (N_4203,N_643,N_1557);
and U4204 (N_4204,N_76,N_1258);
and U4205 (N_4205,N_209,N_2388);
xnor U4206 (N_4206,N_1862,N_1790);
or U4207 (N_4207,N_1484,N_195);
and U4208 (N_4208,N_1533,N_403);
nor U4209 (N_4209,N_2175,N_911);
and U4210 (N_4210,N_1709,N_2035);
and U4211 (N_4211,N_622,N_2184);
nand U4212 (N_4212,N_1808,N_2361);
xor U4213 (N_4213,N_2063,N_823);
nor U4214 (N_4214,N_324,N_987);
or U4215 (N_4215,N_1319,N_330);
xor U4216 (N_4216,N_935,N_1403);
xor U4217 (N_4217,N_1015,N_1146);
nor U4218 (N_4218,N_2028,N_565);
xnor U4219 (N_4219,N_1769,N_1604);
or U4220 (N_4220,N_1286,N_42);
or U4221 (N_4221,N_672,N_527);
or U4222 (N_4222,N_1180,N_2406);
xor U4223 (N_4223,N_2013,N_444);
and U4224 (N_4224,N_2151,N_477);
xor U4225 (N_4225,N_197,N_1331);
or U4226 (N_4226,N_1911,N_2015);
nand U4227 (N_4227,N_841,N_902);
xnor U4228 (N_4228,N_2365,N_2494);
xor U4229 (N_4229,N_271,N_2158);
nand U4230 (N_4230,N_1762,N_1550);
nor U4231 (N_4231,N_1129,N_954);
xor U4232 (N_4232,N_669,N_1732);
nor U4233 (N_4233,N_36,N_969);
nor U4234 (N_4234,N_540,N_1537);
nor U4235 (N_4235,N_236,N_1292);
xor U4236 (N_4236,N_2350,N_984);
or U4237 (N_4237,N_1689,N_2302);
nor U4238 (N_4238,N_1812,N_2181);
xor U4239 (N_4239,N_172,N_1525);
nor U4240 (N_4240,N_1160,N_342);
nor U4241 (N_4241,N_450,N_306);
xnor U4242 (N_4242,N_514,N_424);
nand U4243 (N_4243,N_1795,N_1652);
nor U4244 (N_4244,N_2178,N_394);
nor U4245 (N_4245,N_791,N_66);
or U4246 (N_4246,N_170,N_2494);
or U4247 (N_4247,N_2352,N_1370);
or U4248 (N_4248,N_345,N_188);
nor U4249 (N_4249,N_1831,N_946);
nor U4250 (N_4250,N_1788,N_1561);
and U4251 (N_4251,N_1134,N_2324);
nor U4252 (N_4252,N_1714,N_2360);
xor U4253 (N_4253,N_828,N_915);
nor U4254 (N_4254,N_311,N_265);
or U4255 (N_4255,N_1668,N_1759);
or U4256 (N_4256,N_2033,N_632);
and U4257 (N_4257,N_1169,N_1151);
xnor U4258 (N_4258,N_1637,N_1555);
xnor U4259 (N_4259,N_2237,N_613);
nor U4260 (N_4260,N_524,N_614);
and U4261 (N_4261,N_1791,N_773);
and U4262 (N_4262,N_1889,N_783);
xor U4263 (N_4263,N_1626,N_1694);
and U4264 (N_4264,N_1167,N_1207);
xor U4265 (N_4265,N_1787,N_747);
or U4266 (N_4266,N_648,N_555);
or U4267 (N_4267,N_918,N_2374);
nor U4268 (N_4268,N_1041,N_1244);
xor U4269 (N_4269,N_481,N_2329);
nand U4270 (N_4270,N_1650,N_1906);
nor U4271 (N_4271,N_988,N_1165);
or U4272 (N_4272,N_900,N_1353);
or U4273 (N_4273,N_1808,N_2039);
or U4274 (N_4274,N_792,N_1253);
nor U4275 (N_4275,N_150,N_78);
nand U4276 (N_4276,N_862,N_2417);
xnor U4277 (N_4277,N_2124,N_1219);
or U4278 (N_4278,N_2447,N_293);
nand U4279 (N_4279,N_1872,N_1263);
xor U4280 (N_4280,N_1950,N_822);
nand U4281 (N_4281,N_514,N_1178);
or U4282 (N_4282,N_2236,N_831);
or U4283 (N_4283,N_2095,N_751);
xnor U4284 (N_4284,N_1854,N_1813);
and U4285 (N_4285,N_858,N_29);
or U4286 (N_4286,N_1915,N_641);
and U4287 (N_4287,N_236,N_1686);
xnor U4288 (N_4288,N_1112,N_1586);
nor U4289 (N_4289,N_667,N_1679);
or U4290 (N_4290,N_1152,N_2174);
nor U4291 (N_4291,N_1319,N_1285);
nand U4292 (N_4292,N_1784,N_609);
or U4293 (N_4293,N_764,N_448);
nor U4294 (N_4294,N_1695,N_1976);
and U4295 (N_4295,N_2361,N_884);
xor U4296 (N_4296,N_583,N_2390);
or U4297 (N_4297,N_68,N_1483);
and U4298 (N_4298,N_1494,N_2169);
and U4299 (N_4299,N_1838,N_567);
and U4300 (N_4300,N_828,N_93);
nor U4301 (N_4301,N_578,N_1306);
nand U4302 (N_4302,N_46,N_1875);
and U4303 (N_4303,N_2479,N_2272);
or U4304 (N_4304,N_1678,N_1927);
xnor U4305 (N_4305,N_120,N_2031);
nand U4306 (N_4306,N_1528,N_850);
or U4307 (N_4307,N_326,N_2259);
nor U4308 (N_4308,N_514,N_2435);
or U4309 (N_4309,N_2495,N_1660);
xor U4310 (N_4310,N_1312,N_166);
nor U4311 (N_4311,N_761,N_1574);
nand U4312 (N_4312,N_735,N_840);
or U4313 (N_4313,N_508,N_1733);
nand U4314 (N_4314,N_447,N_2354);
nand U4315 (N_4315,N_547,N_575);
or U4316 (N_4316,N_620,N_1440);
and U4317 (N_4317,N_2223,N_2053);
nor U4318 (N_4318,N_1057,N_263);
xor U4319 (N_4319,N_1378,N_212);
or U4320 (N_4320,N_62,N_1223);
nor U4321 (N_4321,N_1865,N_2197);
or U4322 (N_4322,N_795,N_1969);
and U4323 (N_4323,N_1002,N_466);
or U4324 (N_4324,N_2350,N_1104);
and U4325 (N_4325,N_1761,N_292);
and U4326 (N_4326,N_1569,N_1821);
xnor U4327 (N_4327,N_2183,N_268);
nand U4328 (N_4328,N_1822,N_869);
xnor U4329 (N_4329,N_2434,N_1301);
xor U4330 (N_4330,N_1081,N_2352);
and U4331 (N_4331,N_964,N_1243);
and U4332 (N_4332,N_1507,N_764);
xnor U4333 (N_4333,N_923,N_1829);
nor U4334 (N_4334,N_2380,N_470);
and U4335 (N_4335,N_2065,N_618);
and U4336 (N_4336,N_158,N_1949);
and U4337 (N_4337,N_881,N_63);
or U4338 (N_4338,N_1596,N_2173);
nand U4339 (N_4339,N_1208,N_2128);
and U4340 (N_4340,N_679,N_2168);
and U4341 (N_4341,N_1883,N_773);
xnor U4342 (N_4342,N_1108,N_414);
nor U4343 (N_4343,N_1892,N_1120);
nand U4344 (N_4344,N_501,N_393);
and U4345 (N_4345,N_2066,N_232);
nor U4346 (N_4346,N_998,N_1664);
nand U4347 (N_4347,N_1717,N_2162);
or U4348 (N_4348,N_1448,N_848);
nand U4349 (N_4349,N_1444,N_428);
and U4350 (N_4350,N_710,N_97);
and U4351 (N_4351,N_2257,N_1988);
nand U4352 (N_4352,N_202,N_2021);
or U4353 (N_4353,N_143,N_1611);
xor U4354 (N_4354,N_1623,N_2270);
xor U4355 (N_4355,N_815,N_892);
xnor U4356 (N_4356,N_2347,N_748);
and U4357 (N_4357,N_90,N_1218);
nand U4358 (N_4358,N_1384,N_260);
xnor U4359 (N_4359,N_244,N_249);
or U4360 (N_4360,N_192,N_493);
xnor U4361 (N_4361,N_1275,N_2425);
or U4362 (N_4362,N_1590,N_215);
or U4363 (N_4363,N_1216,N_1920);
xnor U4364 (N_4364,N_1920,N_899);
nand U4365 (N_4365,N_1873,N_726);
xnor U4366 (N_4366,N_16,N_2270);
nand U4367 (N_4367,N_2212,N_930);
nand U4368 (N_4368,N_2462,N_552);
and U4369 (N_4369,N_206,N_515);
nand U4370 (N_4370,N_2457,N_1395);
and U4371 (N_4371,N_992,N_755);
xnor U4372 (N_4372,N_1798,N_1511);
and U4373 (N_4373,N_1371,N_857);
and U4374 (N_4374,N_2421,N_2227);
and U4375 (N_4375,N_1640,N_2498);
xor U4376 (N_4376,N_544,N_2147);
and U4377 (N_4377,N_253,N_1656);
xor U4378 (N_4378,N_281,N_1378);
or U4379 (N_4379,N_713,N_1931);
or U4380 (N_4380,N_1290,N_1713);
nor U4381 (N_4381,N_627,N_1074);
or U4382 (N_4382,N_17,N_468);
xor U4383 (N_4383,N_2349,N_591);
and U4384 (N_4384,N_147,N_1565);
xor U4385 (N_4385,N_343,N_821);
nand U4386 (N_4386,N_2280,N_1455);
nor U4387 (N_4387,N_2263,N_263);
nand U4388 (N_4388,N_1912,N_707);
or U4389 (N_4389,N_1240,N_797);
or U4390 (N_4390,N_1298,N_1865);
and U4391 (N_4391,N_1081,N_278);
or U4392 (N_4392,N_470,N_239);
nand U4393 (N_4393,N_1919,N_1572);
nand U4394 (N_4394,N_1803,N_966);
xnor U4395 (N_4395,N_2306,N_263);
or U4396 (N_4396,N_676,N_1240);
and U4397 (N_4397,N_1794,N_1156);
and U4398 (N_4398,N_1804,N_1450);
and U4399 (N_4399,N_445,N_466);
xor U4400 (N_4400,N_63,N_2235);
xnor U4401 (N_4401,N_216,N_716);
or U4402 (N_4402,N_1145,N_897);
nor U4403 (N_4403,N_1853,N_1390);
and U4404 (N_4404,N_1923,N_2465);
and U4405 (N_4405,N_281,N_1583);
nand U4406 (N_4406,N_2477,N_544);
nor U4407 (N_4407,N_1207,N_885);
or U4408 (N_4408,N_951,N_1236);
nand U4409 (N_4409,N_933,N_173);
nor U4410 (N_4410,N_251,N_1719);
and U4411 (N_4411,N_1526,N_1641);
and U4412 (N_4412,N_2031,N_1486);
and U4413 (N_4413,N_2460,N_2075);
or U4414 (N_4414,N_377,N_1863);
xor U4415 (N_4415,N_1104,N_1727);
or U4416 (N_4416,N_1254,N_596);
xor U4417 (N_4417,N_2314,N_1526);
xor U4418 (N_4418,N_1533,N_1367);
nor U4419 (N_4419,N_2123,N_1816);
xnor U4420 (N_4420,N_856,N_1642);
and U4421 (N_4421,N_1150,N_2385);
xnor U4422 (N_4422,N_1855,N_1705);
nor U4423 (N_4423,N_899,N_1314);
or U4424 (N_4424,N_1290,N_1197);
and U4425 (N_4425,N_1566,N_1458);
nor U4426 (N_4426,N_1422,N_2141);
nand U4427 (N_4427,N_321,N_1640);
nand U4428 (N_4428,N_100,N_931);
xnor U4429 (N_4429,N_800,N_2317);
nand U4430 (N_4430,N_819,N_578);
and U4431 (N_4431,N_2058,N_533);
xnor U4432 (N_4432,N_1823,N_755);
xnor U4433 (N_4433,N_1726,N_2310);
nand U4434 (N_4434,N_1891,N_700);
or U4435 (N_4435,N_2387,N_340);
nor U4436 (N_4436,N_143,N_1986);
xor U4437 (N_4437,N_629,N_517);
nand U4438 (N_4438,N_1963,N_1203);
nor U4439 (N_4439,N_751,N_1469);
nand U4440 (N_4440,N_1431,N_295);
nor U4441 (N_4441,N_1587,N_1955);
or U4442 (N_4442,N_2448,N_2348);
nand U4443 (N_4443,N_839,N_738);
or U4444 (N_4444,N_194,N_325);
nor U4445 (N_4445,N_886,N_1083);
nor U4446 (N_4446,N_68,N_1980);
xnor U4447 (N_4447,N_765,N_804);
nand U4448 (N_4448,N_182,N_705);
nand U4449 (N_4449,N_882,N_2044);
xnor U4450 (N_4450,N_2043,N_142);
nor U4451 (N_4451,N_1650,N_945);
nand U4452 (N_4452,N_2247,N_31);
or U4453 (N_4453,N_602,N_2253);
xor U4454 (N_4454,N_1859,N_132);
and U4455 (N_4455,N_907,N_761);
and U4456 (N_4456,N_20,N_2079);
and U4457 (N_4457,N_2455,N_471);
xnor U4458 (N_4458,N_102,N_87);
xnor U4459 (N_4459,N_1764,N_1814);
and U4460 (N_4460,N_1131,N_1567);
xnor U4461 (N_4461,N_1613,N_157);
xor U4462 (N_4462,N_1913,N_2162);
or U4463 (N_4463,N_1777,N_2084);
nor U4464 (N_4464,N_1078,N_1060);
and U4465 (N_4465,N_1052,N_89);
and U4466 (N_4466,N_573,N_42);
nor U4467 (N_4467,N_1461,N_250);
and U4468 (N_4468,N_710,N_1786);
and U4469 (N_4469,N_1288,N_582);
and U4470 (N_4470,N_1928,N_680);
nor U4471 (N_4471,N_1923,N_1839);
xor U4472 (N_4472,N_1257,N_2348);
xor U4473 (N_4473,N_1633,N_1594);
or U4474 (N_4474,N_2196,N_1440);
nor U4475 (N_4475,N_296,N_1829);
or U4476 (N_4476,N_701,N_953);
xnor U4477 (N_4477,N_178,N_2430);
nand U4478 (N_4478,N_53,N_2380);
nor U4479 (N_4479,N_375,N_361);
xor U4480 (N_4480,N_2026,N_2272);
nand U4481 (N_4481,N_1678,N_859);
and U4482 (N_4482,N_507,N_106);
nor U4483 (N_4483,N_1483,N_826);
nor U4484 (N_4484,N_249,N_2258);
or U4485 (N_4485,N_945,N_1744);
xor U4486 (N_4486,N_139,N_1299);
or U4487 (N_4487,N_604,N_461);
nor U4488 (N_4488,N_1362,N_2356);
nor U4489 (N_4489,N_1204,N_518);
nand U4490 (N_4490,N_1548,N_1518);
nand U4491 (N_4491,N_691,N_2428);
xnor U4492 (N_4492,N_1221,N_642);
or U4493 (N_4493,N_990,N_667);
nor U4494 (N_4494,N_900,N_961);
nand U4495 (N_4495,N_1741,N_1427);
xnor U4496 (N_4496,N_1723,N_2294);
or U4497 (N_4497,N_1445,N_1921);
nor U4498 (N_4498,N_538,N_1427);
nand U4499 (N_4499,N_1387,N_1988);
xnor U4500 (N_4500,N_954,N_1965);
nand U4501 (N_4501,N_1229,N_1127);
nor U4502 (N_4502,N_1437,N_1084);
nor U4503 (N_4503,N_1722,N_1255);
and U4504 (N_4504,N_1608,N_1314);
xnor U4505 (N_4505,N_955,N_340);
nor U4506 (N_4506,N_2068,N_447);
nand U4507 (N_4507,N_38,N_267);
nor U4508 (N_4508,N_1098,N_1819);
xnor U4509 (N_4509,N_1057,N_1865);
xnor U4510 (N_4510,N_1275,N_1683);
nor U4511 (N_4511,N_1329,N_1326);
or U4512 (N_4512,N_2201,N_2187);
nand U4513 (N_4513,N_744,N_1885);
or U4514 (N_4514,N_427,N_2475);
or U4515 (N_4515,N_548,N_1104);
and U4516 (N_4516,N_2068,N_894);
or U4517 (N_4517,N_430,N_1036);
or U4518 (N_4518,N_1560,N_46);
xor U4519 (N_4519,N_746,N_270);
xnor U4520 (N_4520,N_43,N_1474);
or U4521 (N_4521,N_503,N_828);
and U4522 (N_4522,N_1512,N_2255);
nand U4523 (N_4523,N_208,N_588);
and U4524 (N_4524,N_1352,N_1755);
or U4525 (N_4525,N_1348,N_1671);
nand U4526 (N_4526,N_315,N_1570);
nand U4527 (N_4527,N_1739,N_601);
and U4528 (N_4528,N_1180,N_808);
or U4529 (N_4529,N_383,N_528);
xnor U4530 (N_4530,N_1140,N_478);
nand U4531 (N_4531,N_56,N_2443);
xnor U4532 (N_4532,N_1779,N_718);
nor U4533 (N_4533,N_1604,N_1438);
nor U4534 (N_4534,N_345,N_1828);
or U4535 (N_4535,N_350,N_253);
nor U4536 (N_4536,N_1563,N_1754);
or U4537 (N_4537,N_1286,N_2414);
xnor U4538 (N_4538,N_1780,N_109);
and U4539 (N_4539,N_212,N_81);
nand U4540 (N_4540,N_2153,N_2336);
or U4541 (N_4541,N_1916,N_339);
xor U4542 (N_4542,N_1739,N_1479);
nor U4543 (N_4543,N_125,N_121);
or U4544 (N_4544,N_157,N_1121);
xor U4545 (N_4545,N_1941,N_702);
nand U4546 (N_4546,N_532,N_2071);
and U4547 (N_4547,N_1951,N_464);
nand U4548 (N_4548,N_1739,N_1107);
nor U4549 (N_4549,N_1176,N_825);
and U4550 (N_4550,N_1031,N_1084);
nor U4551 (N_4551,N_1174,N_2057);
xor U4552 (N_4552,N_1030,N_1762);
and U4553 (N_4553,N_1557,N_244);
nand U4554 (N_4554,N_2445,N_1032);
and U4555 (N_4555,N_480,N_1683);
xnor U4556 (N_4556,N_610,N_2318);
nand U4557 (N_4557,N_2278,N_1731);
or U4558 (N_4558,N_1418,N_2480);
nand U4559 (N_4559,N_2471,N_556);
xnor U4560 (N_4560,N_1597,N_2098);
xor U4561 (N_4561,N_377,N_1225);
and U4562 (N_4562,N_2160,N_72);
xor U4563 (N_4563,N_1891,N_2436);
and U4564 (N_4564,N_995,N_1011);
nor U4565 (N_4565,N_2108,N_314);
and U4566 (N_4566,N_2487,N_1227);
or U4567 (N_4567,N_701,N_2155);
nor U4568 (N_4568,N_1822,N_1636);
nor U4569 (N_4569,N_2057,N_1986);
nor U4570 (N_4570,N_1647,N_1797);
nand U4571 (N_4571,N_486,N_1454);
or U4572 (N_4572,N_1727,N_236);
nor U4573 (N_4573,N_740,N_2261);
and U4574 (N_4574,N_1597,N_2263);
nor U4575 (N_4575,N_1690,N_1386);
or U4576 (N_4576,N_2322,N_360);
or U4577 (N_4577,N_2468,N_1139);
xor U4578 (N_4578,N_1157,N_182);
nand U4579 (N_4579,N_2499,N_342);
xnor U4580 (N_4580,N_1673,N_2287);
xnor U4581 (N_4581,N_359,N_1164);
nor U4582 (N_4582,N_1285,N_69);
and U4583 (N_4583,N_448,N_464);
xnor U4584 (N_4584,N_625,N_189);
nor U4585 (N_4585,N_1828,N_2477);
nor U4586 (N_4586,N_94,N_416);
and U4587 (N_4587,N_952,N_2383);
or U4588 (N_4588,N_756,N_1952);
nor U4589 (N_4589,N_2041,N_985);
xnor U4590 (N_4590,N_1376,N_994);
nor U4591 (N_4591,N_1898,N_2141);
xor U4592 (N_4592,N_754,N_1203);
or U4593 (N_4593,N_2280,N_2380);
nor U4594 (N_4594,N_680,N_2097);
and U4595 (N_4595,N_2114,N_2313);
and U4596 (N_4596,N_674,N_262);
and U4597 (N_4597,N_614,N_1789);
nand U4598 (N_4598,N_52,N_1973);
nand U4599 (N_4599,N_224,N_239);
and U4600 (N_4600,N_1343,N_116);
nor U4601 (N_4601,N_721,N_2043);
and U4602 (N_4602,N_1333,N_1537);
and U4603 (N_4603,N_1664,N_157);
nor U4604 (N_4604,N_425,N_1089);
xor U4605 (N_4605,N_2293,N_1118);
and U4606 (N_4606,N_1368,N_285);
nand U4607 (N_4607,N_2403,N_1968);
and U4608 (N_4608,N_0,N_1107);
nand U4609 (N_4609,N_1221,N_1157);
xor U4610 (N_4610,N_1205,N_771);
nand U4611 (N_4611,N_2349,N_969);
xor U4612 (N_4612,N_1642,N_830);
and U4613 (N_4613,N_794,N_1356);
or U4614 (N_4614,N_635,N_444);
xnor U4615 (N_4615,N_1183,N_1286);
and U4616 (N_4616,N_495,N_407);
and U4617 (N_4617,N_1628,N_2485);
nand U4618 (N_4618,N_1805,N_1303);
nand U4619 (N_4619,N_1708,N_2440);
and U4620 (N_4620,N_1486,N_455);
or U4621 (N_4621,N_157,N_1637);
nor U4622 (N_4622,N_1776,N_553);
xnor U4623 (N_4623,N_1553,N_1220);
and U4624 (N_4624,N_1520,N_446);
and U4625 (N_4625,N_415,N_2096);
or U4626 (N_4626,N_457,N_775);
and U4627 (N_4627,N_906,N_1362);
or U4628 (N_4628,N_1933,N_583);
nor U4629 (N_4629,N_2437,N_2019);
and U4630 (N_4630,N_2407,N_1541);
nand U4631 (N_4631,N_883,N_1012);
nor U4632 (N_4632,N_840,N_244);
and U4633 (N_4633,N_1831,N_454);
xnor U4634 (N_4634,N_1148,N_922);
nand U4635 (N_4635,N_2255,N_1868);
nand U4636 (N_4636,N_1,N_1679);
and U4637 (N_4637,N_1265,N_2182);
xnor U4638 (N_4638,N_1823,N_689);
or U4639 (N_4639,N_658,N_1506);
nor U4640 (N_4640,N_1529,N_211);
nor U4641 (N_4641,N_1839,N_2153);
and U4642 (N_4642,N_312,N_1742);
nor U4643 (N_4643,N_983,N_1681);
nor U4644 (N_4644,N_850,N_2405);
nor U4645 (N_4645,N_539,N_1532);
nor U4646 (N_4646,N_576,N_2496);
and U4647 (N_4647,N_1391,N_367);
and U4648 (N_4648,N_1668,N_1673);
nor U4649 (N_4649,N_1122,N_1161);
nor U4650 (N_4650,N_1149,N_1781);
and U4651 (N_4651,N_2085,N_1553);
and U4652 (N_4652,N_1971,N_1224);
or U4653 (N_4653,N_311,N_233);
nand U4654 (N_4654,N_1234,N_1376);
and U4655 (N_4655,N_2096,N_2070);
and U4656 (N_4656,N_228,N_2353);
and U4657 (N_4657,N_598,N_814);
nor U4658 (N_4658,N_1040,N_1961);
or U4659 (N_4659,N_1182,N_2381);
xor U4660 (N_4660,N_896,N_229);
and U4661 (N_4661,N_1431,N_1257);
or U4662 (N_4662,N_713,N_1150);
nand U4663 (N_4663,N_1652,N_2170);
and U4664 (N_4664,N_81,N_2341);
nand U4665 (N_4665,N_274,N_2256);
xor U4666 (N_4666,N_1178,N_630);
nand U4667 (N_4667,N_1885,N_1396);
nand U4668 (N_4668,N_1631,N_909);
nor U4669 (N_4669,N_767,N_2029);
nor U4670 (N_4670,N_1630,N_176);
xor U4671 (N_4671,N_2052,N_1409);
nand U4672 (N_4672,N_1614,N_243);
nor U4673 (N_4673,N_2188,N_594);
nand U4674 (N_4674,N_951,N_637);
and U4675 (N_4675,N_1557,N_862);
nor U4676 (N_4676,N_1297,N_448);
nand U4677 (N_4677,N_1621,N_2355);
nor U4678 (N_4678,N_2160,N_1496);
or U4679 (N_4679,N_682,N_1323);
or U4680 (N_4680,N_2082,N_1150);
nor U4681 (N_4681,N_295,N_2213);
and U4682 (N_4682,N_2414,N_1921);
or U4683 (N_4683,N_1652,N_1406);
nor U4684 (N_4684,N_962,N_956);
nand U4685 (N_4685,N_1608,N_121);
or U4686 (N_4686,N_890,N_1102);
or U4687 (N_4687,N_1312,N_2049);
or U4688 (N_4688,N_1758,N_259);
nand U4689 (N_4689,N_7,N_947);
and U4690 (N_4690,N_2093,N_2223);
xor U4691 (N_4691,N_1102,N_808);
nand U4692 (N_4692,N_2230,N_636);
and U4693 (N_4693,N_755,N_428);
and U4694 (N_4694,N_1081,N_1209);
nor U4695 (N_4695,N_2134,N_2227);
xor U4696 (N_4696,N_1457,N_910);
nor U4697 (N_4697,N_192,N_2189);
nor U4698 (N_4698,N_96,N_805);
or U4699 (N_4699,N_1007,N_2307);
nand U4700 (N_4700,N_141,N_1013);
xor U4701 (N_4701,N_2058,N_2093);
nor U4702 (N_4702,N_1550,N_883);
xnor U4703 (N_4703,N_2023,N_1924);
or U4704 (N_4704,N_1105,N_1015);
nand U4705 (N_4705,N_1047,N_163);
and U4706 (N_4706,N_671,N_281);
and U4707 (N_4707,N_1105,N_305);
and U4708 (N_4708,N_2158,N_343);
and U4709 (N_4709,N_1162,N_543);
nand U4710 (N_4710,N_1030,N_1219);
and U4711 (N_4711,N_804,N_1177);
xnor U4712 (N_4712,N_1474,N_1740);
xnor U4713 (N_4713,N_63,N_843);
nand U4714 (N_4714,N_974,N_791);
or U4715 (N_4715,N_1228,N_2400);
xnor U4716 (N_4716,N_237,N_1495);
xnor U4717 (N_4717,N_1482,N_9);
and U4718 (N_4718,N_2218,N_324);
nor U4719 (N_4719,N_1931,N_416);
and U4720 (N_4720,N_153,N_1410);
nand U4721 (N_4721,N_1796,N_35);
nor U4722 (N_4722,N_673,N_2379);
and U4723 (N_4723,N_2272,N_533);
and U4724 (N_4724,N_803,N_429);
or U4725 (N_4725,N_54,N_906);
and U4726 (N_4726,N_204,N_42);
xor U4727 (N_4727,N_2327,N_998);
or U4728 (N_4728,N_1048,N_1906);
and U4729 (N_4729,N_1399,N_944);
nand U4730 (N_4730,N_1963,N_1311);
xnor U4731 (N_4731,N_820,N_1876);
or U4732 (N_4732,N_649,N_2369);
and U4733 (N_4733,N_1791,N_537);
or U4734 (N_4734,N_346,N_1809);
and U4735 (N_4735,N_713,N_2162);
xor U4736 (N_4736,N_1268,N_527);
and U4737 (N_4737,N_2482,N_1290);
nor U4738 (N_4738,N_551,N_254);
xor U4739 (N_4739,N_763,N_861);
and U4740 (N_4740,N_191,N_1175);
nor U4741 (N_4741,N_844,N_1448);
xor U4742 (N_4742,N_2209,N_2354);
xor U4743 (N_4743,N_1935,N_92);
and U4744 (N_4744,N_1971,N_1393);
nand U4745 (N_4745,N_1449,N_2245);
nor U4746 (N_4746,N_1632,N_764);
nor U4747 (N_4747,N_895,N_1484);
and U4748 (N_4748,N_735,N_170);
xor U4749 (N_4749,N_2185,N_1169);
and U4750 (N_4750,N_680,N_253);
nor U4751 (N_4751,N_363,N_1926);
xnor U4752 (N_4752,N_124,N_1957);
nor U4753 (N_4753,N_1302,N_1274);
nand U4754 (N_4754,N_2471,N_2243);
or U4755 (N_4755,N_2137,N_327);
or U4756 (N_4756,N_2150,N_2163);
nor U4757 (N_4757,N_18,N_1639);
xor U4758 (N_4758,N_714,N_1574);
and U4759 (N_4759,N_1332,N_2240);
nand U4760 (N_4760,N_1470,N_2032);
and U4761 (N_4761,N_1871,N_316);
xnor U4762 (N_4762,N_685,N_1193);
or U4763 (N_4763,N_1499,N_1789);
and U4764 (N_4764,N_172,N_690);
nor U4765 (N_4765,N_2126,N_651);
and U4766 (N_4766,N_2276,N_175);
or U4767 (N_4767,N_1752,N_1861);
xnor U4768 (N_4768,N_247,N_766);
and U4769 (N_4769,N_619,N_2344);
or U4770 (N_4770,N_2260,N_584);
nor U4771 (N_4771,N_114,N_304);
nor U4772 (N_4772,N_1417,N_1713);
and U4773 (N_4773,N_2282,N_1869);
or U4774 (N_4774,N_199,N_2117);
and U4775 (N_4775,N_329,N_2354);
or U4776 (N_4776,N_1490,N_2161);
xor U4777 (N_4777,N_810,N_539);
nand U4778 (N_4778,N_1382,N_2448);
or U4779 (N_4779,N_426,N_1578);
or U4780 (N_4780,N_1083,N_291);
xnor U4781 (N_4781,N_2390,N_260);
xor U4782 (N_4782,N_856,N_1456);
xnor U4783 (N_4783,N_1050,N_2026);
and U4784 (N_4784,N_2051,N_1915);
xnor U4785 (N_4785,N_2065,N_2007);
or U4786 (N_4786,N_1872,N_2445);
nand U4787 (N_4787,N_2372,N_763);
nor U4788 (N_4788,N_923,N_1417);
or U4789 (N_4789,N_1786,N_1835);
nand U4790 (N_4790,N_475,N_415);
and U4791 (N_4791,N_570,N_1924);
and U4792 (N_4792,N_617,N_1106);
or U4793 (N_4793,N_2278,N_3);
xnor U4794 (N_4794,N_179,N_2013);
and U4795 (N_4795,N_1548,N_1629);
or U4796 (N_4796,N_1695,N_1925);
nand U4797 (N_4797,N_337,N_1333);
nor U4798 (N_4798,N_1495,N_286);
xnor U4799 (N_4799,N_556,N_2054);
xor U4800 (N_4800,N_2397,N_282);
nor U4801 (N_4801,N_282,N_403);
or U4802 (N_4802,N_1983,N_439);
and U4803 (N_4803,N_1388,N_480);
or U4804 (N_4804,N_1532,N_671);
or U4805 (N_4805,N_75,N_2340);
nand U4806 (N_4806,N_1501,N_415);
nand U4807 (N_4807,N_805,N_441);
or U4808 (N_4808,N_1904,N_1597);
nand U4809 (N_4809,N_576,N_76);
or U4810 (N_4810,N_805,N_484);
xnor U4811 (N_4811,N_102,N_903);
nand U4812 (N_4812,N_1607,N_389);
or U4813 (N_4813,N_1253,N_71);
and U4814 (N_4814,N_752,N_1623);
and U4815 (N_4815,N_1935,N_476);
and U4816 (N_4816,N_942,N_812);
and U4817 (N_4817,N_770,N_1830);
nand U4818 (N_4818,N_445,N_1208);
xor U4819 (N_4819,N_305,N_1280);
nand U4820 (N_4820,N_89,N_22);
nor U4821 (N_4821,N_1822,N_80);
nor U4822 (N_4822,N_1394,N_1312);
and U4823 (N_4823,N_1986,N_204);
or U4824 (N_4824,N_2274,N_134);
nand U4825 (N_4825,N_1653,N_685);
nor U4826 (N_4826,N_1334,N_1505);
nor U4827 (N_4827,N_1835,N_1918);
nor U4828 (N_4828,N_378,N_2210);
nor U4829 (N_4829,N_730,N_662);
nand U4830 (N_4830,N_1225,N_2164);
nor U4831 (N_4831,N_745,N_644);
and U4832 (N_4832,N_2251,N_528);
nand U4833 (N_4833,N_1035,N_1589);
nand U4834 (N_4834,N_2447,N_370);
xnor U4835 (N_4835,N_125,N_1945);
nor U4836 (N_4836,N_1672,N_2213);
and U4837 (N_4837,N_1689,N_1882);
nand U4838 (N_4838,N_1242,N_1398);
or U4839 (N_4839,N_1557,N_1275);
and U4840 (N_4840,N_312,N_502);
nor U4841 (N_4841,N_1601,N_2283);
nand U4842 (N_4842,N_2170,N_2347);
nor U4843 (N_4843,N_1099,N_535);
nand U4844 (N_4844,N_1378,N_1646);
or U4845 (N_4845,N_470,N_1014);
nor U4846 (N_4846,N_117,N_2449);
xnor U4847 (N_4847,N_1807,N_1213);
or U4848 (N_4848,N_1781,N_941);
and U4849 (N_4849,N_434,N_575);
xnor U4850 (N_4850,N_2333,N_354);
nand U4851 (N_4851,N_2341,N_732);
nand U4852 (N_4852,N_1869,N_2120);
nor U4853 (N_4853,N_1918,N_357);
xnor U4854 (N_4854,N_788,N_421);
nor U4855 (N_4855,N_1449,N_800);
or U4856 (N_4856,N_1732,N_2034);
or U4857 (N_4857,N_1842,N_2386);
nor U4858 (N_4858,N_482,N_244);
and U4859 (N_4859,N_1357,N_2454);
or U4860 (N_4860,N_306,N_604);
nor U4861 (N_4861,N_16,N_273);
or U4862 (N_4862,N_1322,N_2109);
nand U4863 (N_4863,N_1524,N_1327);
and U4864 (N_4864,N_1876,N_1727);
and U4865 (N_4865,N_1686,N_773);
xor U4866 (N_4866,N_189,N_2319);
nor U4867 (N_4867,N_969,N_627);
xnor U4868 (N_4868,N_76,N_463);
nand U4869 (N_4869,N_139,N_1022);
nor U4870 (N_4870,N_966,N_1500);
xnor U4871 (N_4871,N_297,N_1587);
and U4872 (N_4872,N_683,N_231);
nor U4873 (N_4873,N_1639,N_1080);
and U4874 (N_4874,N_302,N_451);
nor U4875 (N_4875,N_1300,N_2213);
xnor U4876 (N_4876,N_1498,N_673);
or U4877 (N_4877,N_914,N_932);
xor U4878 (N_4878,N_2417,N_303);
xnor U4879 (N_4879,N_2313,N_383);
nor U4880 (N_4880,N_814,N_1437);
and U4881 (N_4881,N_1409,N_1549);
nand U4882 (N_4882,N_2492,N_2155);
and U4883 (N_4883,N_853,N_1365);
nand U4884 (N_4884,N_2437,N_135);
xnor U4885 (N_4885,N_600,N_1069);
nand U4886 (N_4886,N_1345,N_573);
or U4887 (N_4887,N_54,N_110);
or U4888 (N_4888,N_1187,N_183);
and U4889 (N_4889,N_2446,N_1365);
nor U4890 (N_4890,N_156,N_909);
xnor U4891 (N_4891,N_1268,N_429);
nand U4892 (N_4892,N_2208,N_930);
xor U4893 (N_4893,N_2437,N_2410);
nand U4894 (N_4894,N_2031,N_2481);
nand U4895 (N_4895,N_1815,N_1934);
xor U4896 (N_4896,N_2261,N_1953);
nor U4897 (N_4897,N_2355,N_201);
xnor U4898 (N_4898,N_1058,N_129);
xnor U4899 (N_4899,N_855,N_1230);
xor U4900 (N_4900,N_512,N_1148);
nand U4901 (N_4901,N_727,N_1092);
nor U4902 (N_4902,N_2094,N_2497);
and U4903 (N_4903,N_702,N_587);
xor U4904 (N_4904,N_1555,N_1493);
nand U4905 (N_4905,N_383,N_1181);
nand U4906 (N_4906,N_1664,N_1545);
nand U4907 (N_4907,N_1502,N_690);
nand U4908 (N_4908,N_287,N_576);
or U4909 (N_4909,N_322,N_2284);
nand U4910 (N_4910,N_323,N_784);
or U4911 (N_4911,N_1917,N_629);
or U4912 (N_4912,N_938,N_1795);
or U4913 (N_4913,N_1836,N_1712);
and U4914 (N_4914,N_1993,N_1466);
nor U4915 (N_4915,N_783,N_1083);
or U4916 (N_4916,N_1382,N_657);
and U4917 (N_4917,N_544,N_2334);
nand U4918 (N_4918,N_1506,N_138);
and U4919 (N_4919,N_1839,N_2088);
nor U4920 (N_4920,N_91,N_1929);
and U4921 (N_4921,N_563,N_89);
and U4922 (N_4922,N_143,N_770);
xor U4923 (N_4923,N_2412,N_2402);
or U4924 (N_4924,N_2084,N_719);
and U4925 (N_4925,N_1544,N_919);
or U4926 (N_4926,N_567,N_139);
nor U4927 (N_4927,N_1525,N_529);
and U4928 (N_4928,N_687,N_558);
or U4929 (N_4929,N_1343,N_784);
xnor U4930 (N_4930,N_1573,N_905);
or U4931 (N_4931,N_106,N_447);
or U4932 (N_4932,N_795,N_284);
nor U4933 (N_4933,N_610,N_157);
nor U4934 (N_4934,N_1338,N_1278);
and U4935 (N_4935,N_639,N_101);
nor U4936 (N_4936,N_784,N_286);
nand U4937 (N_4937,N_316,N_1350);
or U4938 (N_4938,N_275,N_2465);
nand U4939 (N_4939,N_264,N_1817);
nor U4940 (N_4940,N_135,N_1433);
nand U4941 (N_4941,N_60,N_1430);
nor U4942 (N_4942,N_450,N_1602);
and U4943 (N_4943,N_503,N_2432);
or U4944 (N_4944,N_840,N_799);
and U4945 (N_4945,N_1397,N_1066);
and U4946 (N_4946,N_2244,N_238);
or U4947 (N_4947,N_658,N_1415);
nand U4948 (N_4948,N_13,N_1411);
or U4949 (N_4949,N_1906,N_1333);
and U4950 (N_4950,N_2128,N_1329);
xnor U4951 (N_4951,N_114,N_534);
xor U4952 (N_4952,N_191,N_2055);
nand U4953 (N_4953,N_2185,N_2334);
nand U4954 (N_4954,N_1074,N_603);
nand U4955 (N_4955,N_930,N_975);
nand U4956 (N_4956,N_477,N_1279);
or U4957 (N_4957,N_2073,N_1486);
nand U4958 (N_4958,N_441,N_2460);
or U4959 (N_4959,N_528,N_2097);
nand U4960 (N_4960,N_859,N_641);
nor U4961 (N_4961,N_1764,N_2107);
nor U4962 (N_4962,N_2032,N_1326);
and U4963 (N_4963,N_578,N_454);
and U4964 (N_4964,N_1385,N_2393);
nand U4965 (N_4965,N_10,N_666);
and U4966 (N_4966,N_212,N_242);
or U4967 (N_4967,N_2138,N_241);
and U4968 (N_4968,N_2028,N_758);
xor U4969 (N_4969,N_1304,N_64);
nor U4970 (N_4970,N_2141,N_2378);
nor U4971 (N_4971,N_109,N_278);
xnor U4972 (N_4972,N_1510,N_788);
or U4973 (N_4973,N_2327,N_702);
xor U4974 (N_4974,N_452,N_182);
nand U4975 (N_4975,N_184,N_1839);
nor U4976 (N_4976,N_1803,N_1593);
or U4977 (N_4977,N_2,N_83);
or U4978 (N_4978,N_1861,N_1108);
and U4979 (N_4979,N_986,N_1106);
and U4980 (N_4980,N_660,N_84);
and U4981 (N_4981,N_509,N_617);
nor U4982 (N_4982,N_1063,N_612);
nand U4983 (N_4983,N_220,N_2213);
and U4984 (N_4984,N_2106,N_1583);
nand U4985 (N_4985,N_342,N_816);
nand U4986 (N_4986,N_2426,N_1849);
xnor U4987 (N_4987,N_1549,N_2286);
xnor U4988 (N_4988,N_434,N_1196);
nor U4989 (N_4989,N_477,N_2214);
and U4990 (N_4990,N_1483,N_1978);
or U4991 (N_4991,N_368,N_1206);
or U4992 (N_4992,N_1121,N_1638);
or U4993 (N_4993,N_1907,N_1408);
and U4994 (N_4994,N_2056,N_24);
and U4995 (N_4995,N_1273,N_2486);
nor U4996 (N_4996,N_741,N_517);
nor U4997 (N_4997,N_571,N_1011);
nor U4998 (N_4998,N_1551,N_2130);
nor U4999 (N_4999,N_1350,N_399);
xnor U5000 (N_5000,N_3981,N_4738);
nand U5001 (N_5001,N_3712,N_4016);
nand U5002 (N_5002,N_4229,N_4062);
or U5003 (N_5003,N_4419,N_3409);
nand U5004 (N_5004,N_2989,N_2506);
and U5005 (N_5005,N_4575,N_2845);
and U5006 (N_5006,N_4339,N_3542);
or U5007 (N_5007,N_4493,N_2945);
xor U5008 (N_5008,N_3722,N_3579);
or U5009 (N_5009,N_2515,N_4314);
and U5010 (N_5010,N_3753,N_2511);
xnor U5011 (N_5011,N_2628,N_2541);
or U5012 (N_5012,N_3291,N_2790);
xnor U5013 (N_5013,N_3425,N_3136);
xor U5014 (N_5014,N_2668,N_2882);
and U5015 (N_5015,N_2600,N_3193);
and U5016 (N_5016,N_2608,N_4191);
nor U5017 (N_5017,N_3661,N_3419);
and U5018 (N_5018,N_2656,N_3704);
nor U5019 (N_5019,N_2974,N_2630);
nand U5020 (N_5020,N_3870,N_4410);
nand U5021 (N_5021,N_3139,N_4904);
xor U5022 (N_5022,N_4031,N_3792);
nand U5023 (N_5023,N_3846,N_2926);
or U5024 (N_5024,N_4330,N_4392);
nor U5025 (N_5025,N_3490,N_3669);
or U5026 (N_5026,N_4847,N_4642);
nor U5027 (N_5027,N_3241,N_4375);
and U5028 (N_5028,N_3698,N_3924);
xnor U5029 (N_5029,N_2864,N_3342);
nor U5030 (N_5030,N_2946,N_2761);
nand U5031 (N_5031,N_4781,N_3585);
and U5032 (N_5032,N_3956,N_3536);
nor U5033 (N_5033,N_3236,N_2723);
nor U5034 (N_5034,N_3875,N_4487);
or U5035 (N_5035,N_3338,N_4131);
nand U5036 (N_5036,N_3955,N_3134);
nand U5037 (N_5037,N_3246,N_4301);
nand U5038 (N_5038,N_4013,N_4849);
nor U5039 (N_5039,N_3828,N_4261);
nor U5040 (N_5040,N_3449,N_3781);
nand U5041 (N_5041,N_3610,N_3808);
nand U5042 (N_5042,N_3160,N_3842);
nor U5043 (N_5043,N_2748,N_4030);
and U5044 (N_5044,N_4736,N_4910);
xnor U5045 (N_5045,N_4961,N_3263);
and U5046 (N_5046,N_3595,N_3575);
xor U5047 (N_5047,N_4058,N_2907);
nand U5048 (N_5048,N_3421,N_2805);
xnor U5049 (N_5049,N_3228,N_3582);
or U5050 (N_5050,N_4464,N_4799);
or U5051 (N_5051,N_2922,N_3878);
xor U5052 (N_5052,N_4675,N_3937);
and U5053 (N_5053,N_4621,N_2510);
xnor U5054 (N_5054,N_3057,N_4071);
nand U5055 (N_5055,N_3731,N_4587);
nand U5056 (N_5056,N_3564,N_2942);
nand U5057 (N_5057,N_3777,N_2767);
or U5058 (N_5058,N_4530,N_4443);
or U5059 (N_5059,N_3049,N_3133);
nor U5060 (N_5060,N_4853,N_4566);
nand U5061 (N_5061,N_3566,N_3560);
or U5062 (N_5062,N_2521,N_3090);
nor U5063 (N_5063,N_2919,N_3527);
or U5064 (N_5064,N_3507,N_3337);
nor U5065 (N_5065,N_4121,N_3882);
xnor U5066 (N_5066,N_4038,N_4551);
nor U5067 (N_5067,N_3772,N_3004);
xor U5068 (N_5068,N_3561,N_4693);
nor U5069 (N_5069,N_4457,N_4043);
or U5070 (N_5070,N_2673,N_3910);
nand U5071 (N_5071,N_4879,N_2858);
and U5072 (N_5072,N_3457,N_4559);
nand U5073 (N_5073,N_4913,N_2635);
or U5074 (N_5074,N_4873,N_4814);
nor U5075 (N_5075,N_3300,N_2804);
nor U5076 (N_5076,N_4204,N_4816);
nor U5077 (N_5077,N_4912,N_3369);
or U5078 (N_5078,N_3167,N_3638);
nand U5079 (N_5079,N_4571,N_3165);
xnor U5080 (N_5080,N_2976,N_4743);
and U5081 (N_5081,N_3353,N_3535);
nand U5082 (N_5082,N_3720,N_4715);
xor U5083 (N_5083,N_2969,N_2718);
xnor U5084 (N_5084,N_3015,N_3306);
nor U5085 (N_5085,N_3968,N_3410);
or U5086 (N_5086,N_3809,N_2717);
nor U5087 (N_5087,N_2513,N_3696);
xnor U5088 (N_5088,N_4285,N_2815);
xor U5089 (N_5089,N_4854,N_4288);
nor U5090 (N_5090,N_3444,N_4094);
and U5091 (N_5091,N_4304,N_3050);
nand U5092 (N_5092,N_4033,N_4984);
nand U5093 (N_5093,N_4472,N_3584);
xor U5094 (N_5094,N_4390,N_4459);
and U5095 (N_5095,N_3554,N_4309);
xor U5096 (N_5096,N_2712,N_4821);
nand U5097 (N_5097,N_3824,N_4686);
and U5098 (N_5098,N_4117,N_3628);
and U5099 (N_5099,N_3740,N_3303);
and U5100 (N_5100,N_3904,N_3774);
nand U5101 (N_5101,N_4277,N_4284);
nor U5102 (N_5102,N_2705,N_2849);
nand U5103 (N_5103,N_4810,N_4783);
xnor U5104 (N_5104,N_3395,N_4207);
xor U5105 (N_5105,N_3516,N_3547);
xnor U5106 (N_5106,N_3790,N_3392);
nor U5107 (N_5107,N_3270,N_3546);
xnor U5108 (N_5108,N_4046,N_3975);
xor U5109 (N_5109,N_4964,N_3298);
and U5110 (N_5110,N_3838,N_3806);
nor U5111 (N_5111,N_4612,N_4735);
and U5112 (N_5112,N_4084,N_4108);
and U5113 (N_5113,N_3744,N_4265);
nand U5114 (N_5114,N_2986,N_4927);
xnor U5115 (N_5115,N_2597,N_4272);
nor U5116 (N_5116,N_3636,N_3769);
and U5117 (N_5117,N_3428,N_4504);
or U5118 (N_5118,N_4196,N_4300);
xor U5119 (N_5119,N_4943,N_2592);
and U5120 (N_5120,N_3803,N_2870);
or U5121 (N_5121,N_3733,N_3592);
nand U5122 (N_5122,N_4906,N_2915);
or U5123 (N_5123,N_2566,N_3570);
or U5124 (N_5124,N_2885,N_3430);
xor U5125 (N_5125,N_4998,N_4403);
nand U5126 (N_5126,N_4951,N_3715);
xor U5127 (N_5127,N_3323,N_2822);
nor U5128 (N_5128,N_3426,N_3970);
nand U5129 (N_5129,N_4919,N_4548);
and U5130 (N_5130,N_3301,N_4510);
or U5131 (N_5131,N_4340,N_4660);
and U5132 (N_5132,N_3003,N_2619);
and U5133 (N_5133,N_3620,N_4159);
and U5134 (N_5134,N_3094,N_2990);
and U5135 (N_5135,N_4690,N_2602);
nand U5136 (N_5136,N_2734,N_4492);
nor U5137 (N_5137,N_4531,N_4422);
nor U5138 (N_5138,N_3710,N_2832);
nor U5139 (N_5139,N_4994,N_3484);
nor U5140 (N_5140,N_3158,N_3309);
and U5141 (N_5141,N_4862,N_2618);
xnor U5142 (N_5142,N_3260,N_2724);
and U5143 (N_5143,N_2562,N_3477);
or U5144 (N_5144,N_3416,N_4005);
or U5145 (N_5145,N_3209,N_3544);
or U5146 (N_5146,N_2979,N_3630);
and U5147 (N_5147,N_3349,N_4240);
nand U5148 (N_5148,N_4652,N_2752);
nand U5149 (N_5149,N_3952,N_4673);
nor U5150 (N_5150,N_4553,N_3601);
and U5151 (N_5151,N_3384,N_3683);
xnor U5152 (N_5152,N_4537,N_3156);
xnor U5153 (N_5153,N_2873,N_4750);
nand U5154 (N_5154,N_3130,N_3782);
or U5155 (N_5155,N_4971,N_4795);
or U5156 (N_5156,N_4831,N_3773);
nor U5157 (N_5157,N_3692,N_4331);
nor U5158 (N_5158,N_3014,N_4682);
or U5159 (N_5159,N_4593,N_2689);
nor U5160 (N_5160,N_2538,N_3599);
nand U5161 (N_5161,N_2936,N_4028);
or U5162 (N_5162,N_3044,N_3859);
and U5163 (N_5163,N_3713,N_4896);
and U5164 (N_5164,N_4133,N_2637);
xnor U5165 (N_5165,N_2737,N_3922);
xor U5166 (N_5166,N_4125,N_4397);
or U5167 (N_5167,N_4678,N_4112);
or U5168 (N_5168,N_4075,N_3695);
and U5169 (N_5169,N_2728,N_4498);
nand U5170 (N_5170,N_2794,N_4624);
xor U5171 (N_5171,N_3650,N_3286);
nand U5172 (N_5172,N_3857,N_4096);
nand U5173 (N_5173,N_2739,N_4177);
nand U5174 (N_5174,N_3245,N_3572);
or U5175 (N_5175,N_4655,N_3491);
nand U5176 (N_5176,N_4221,N_2660);
xnor U5177 (N_5177,N_4476,N_4730);
and U5178 (N_5178,N_2977,N_4485);
or U5179 (N_5179,N_3063,N_4577);
nor U5180 (N_5180,N_2740,N_3760);
nand U5181 (N_5181,N_2777,N_3187);
nand U5182 (N_5182,N_2759,N_3198);
nand U5183 (N_5183,N_4244,N_4313);
nor U5184 (N_5184,N_3819,N_3267);
and U5185 (N_5185,N_4921,N_3674);
or U5186 (N_5186,N_2590,N_4641);
nand U5187 (N_5187,N_4440,N_3997);
nand U5188 (N_5188,N_4562,N_2782);
and U5189 (N_5189,N_4463,N_4496);
or U5190 (N_5190,N_3205,N_2824);
nand U5191 (N_5191,N_3771,N_4305);
and U5192 (N_5192,N_4555,N_4480);
xor U5193 (N_5193,N_3532,N_4507);
nor U5194 (N_5194,N_3213,N_3990);
xor U5195 (N_5195,N_2738,N_3438);
xnor U5196 (N_5196,N_3707,N_3874);
nor U5197 (N_5197,N_3103,N_2935);
nand U5198 (N_5198,N_4742,N_3569);
xor U5199 (N_5199,N_3604,N_4585);
xnor U5200 (N_5200,N_4518,N_2779);
nand U5201 (N_5201,N_2693,N_4725);
xor U5202 (N_5202,N_3919,N_3664);
or U5203 (N_5203,N_3195,N_3675);
xnor U5204 (N_5204,N_2726,N_3653);
nand U5205 (N_5205,N_3957,N_3625);
nor U5206 (N_5206,N_3702,N_4249);
or U5207 (N_5207,N_4460,N_4850);
nand U5208 (N_5208,N_3708,N_3087);
nand U5209 (N_5209,N_4638,N_3497);
nor U5210 (N_5210,N_4271,N_2651);
xor U5211 (N_5211,N_3178,N_2902);
and U5212 (N_5212,N_2653,N_3266);
nand U5213 (N_5213,N_3853,N_3040);
nand U5214 (N_5214,N_4384,N_4701);
nand U5215 (N_5215,N_3468,N_3903);
xnor U5216 (N_5216,N_4465,N_3998);
nand U5217 (N_5217,N_2925,N_3471);
nor U5218 (N_5218,N_4428,N_2576);
and U5219 (N_5219,N_4570,N_4825);
xor U5220 (N_5220,N_4635,N_4944);
and U5221 (N_5221,N_3995,N_2793);
nor U5222 (N_5222,N_4000,N_4892);
nor U5223 (N_5223,N_3615,N_4081);
and U5224 (N_5224,N_4461,N_2943);
or U5225 (N_5225,N_3255,N_3510);
and U5226 (N_5226,N_4645,N_3999);
and U5227 (N_5227,N_3609,N_4891);
nand U5228 (N_5228,N_4223,N_3437);
or U5229 (N_5229,N_4274,N_4389);
nand U5230 (N_5230,N_4120,N_3310);
and U5231 (N_5231,N_4070,N_3032);
and U5232 (N_5232,N_2580,N_4431);
and U5233 (N_5233,N_3487,N_4595);
nand U5234 (N_5234,N_3574,N_2677);
nor U5235 (N_5235,N_3668,N_4748);
xor U5236 (N_5236,N_2509,N_4357);
nand U5237 (N_5237,N_3519,N_3069);
and U5238 (N_5238,N_4294,N_3233);
or U5239 (N_5239,N_3109,N_4224);
xnor U5240 (N_5240,N_4753,N_4909);
nand U5241 (N_5241,N_4206,N_3751);
nand U5242 (N_5242,N_3594,N_4486);
or U5243 (N_5243,N_3839,N_3046);
and U5244 (N_5244,N_3617,N_4728);
or U5245 (N_5245,N_4606,N_3450);
or U5246 (N_5246,N_3357,N_3591);
and U5247 (N_5247,N_3184,N_4015);
nand U5248 (N_5248,N_4266,N_4889);
nor U5249 (N_5249,N_3831,N_4158);
and U5250 (N_5250,N_4657,N_4004);
nand U5251 (N_5251,N_2964,N_4747);
xnor U5252 (N_5252,N_2847,N_3505);
nor U5253 (N_5253,N_4296,N_4306);
xnor U5254 (N_5254,N_2931,N_4996);
nand U5255 (N_5255,N_3935,N_3587);
and U5256 (N_5256,N_3833,N_4572);
nor U5257 (N_5257,N_3755,N_2980);
and U5258 (N_5258,N_3917,N_3432);
and U5259 (N_5259,N_3898,N_2833);
nand U5260 (N_5260,N_4356,N_4733);
or U5261 (N_5261,N_4199,N_2534);
nand U5262 (N_5262,N_3711,N_3688);
xnor U5263 (N_5263,N_2856,N_2801);
nand U5264 (N_5264,N_2621,N_4669);
and U5265 (N_5265,N_4448,N_2899);
xnor U5266 (N_5266,N_4222,N_3548);
and U5267 (N_5267,N_3538,N_3622);
or U5268 (N_5268,N_3647,N_3322);
nand U5269 (N_5269,N_2987,N_3210);
xor U5270 (N_5270,N_3912,N_2780);
nand U5271 (N_5271,N_4063,N_4823);
nor U5272 (N_5272,N_4517,N_4111);
xor U5273 (N_5273,N_3316,N_4582);
or U5274 (N_5274,N_3443,N_2883);
and U5275 (N_5275,N_3026,N_3915);
nor U5276 (N_5276,N_4774,N_4937);
nand U5277 (N_5277,N_3374,N_3693);
nand U5278 (N_5278,N_4218,N_4395);
and U5279 (N_5279,N_4547,N_3199);
xor U5280 (N_5280,N_4034,N_2788);
and U5281 (N_5281,N_3092,N_4438);
and U5282 (N_5282,N_4543,N_4036);
and U5283 (N_5283,N_3941,N_4771);
and U5284 (N_5284,N_2679,N_2898);
nor U5285 (N_5285,N_4534,N_3231);
or U5286 (N_5286,N_4414,N_4110);
nor U5287 (N_5287,N_3562,N_3146);
nor U5288 (N_5288,N_3216,N_4706);
or U5289 (N_5289,N_3754,N_4037);
xor U5290 (N_5290,N_4415,N_3775);
or U5291 (N_5291,N_4664,N_2877);
xor U5292 (N_5292,N_2839,N_4077);
nand U5293 (N_5293,N_4691,N_3151);
xor U5294 (N_5294,N_2881,N_4456);
xnor U5295 (N_5295,N_2722,N_3634);
and U5296 (N_5296,N_3344,N_3835);
or U5297 (N_5297,N_3041,N_3967);
nand U5298 (N_5298,N_2851,N_4405);
and U5299 (N_5299,N_4132,N_3393);
nor U5300 (N_5300,N_2760,N_2720);
and U5301 (N_5301,N_3404,N_4977);
or U5302 (N_5302,N_4928,N_3964);
nand U5303 (N_5303,N_4830,N_2762);
xnor U5304 (N_5304,N_2690,N_3480);
or U5305 (N_5305,N_4208,N_4985);
and U5306 (N_5306,N_2518,N_3802);
xnor U5307 (N_5307,N_3479,N_3991);
nor U5308 (N_5308,N_3992,N_4180);
or U5309 (N_5309,N_3515,N_2692);
xnor U5310 (N_5310,N_4088,N_3745);
nand U5311 (N_5311,N_4175,N_4716);
xor U5312 (N_5312,N_3402,N_3537);
xor U5313 (N_5313,N_2905,N_4039);
and U5314 (N_5314,N_2984,N_3363);
and U5315 (N_5315,N_3261,N_4417);
and U5316 (N_5316,N_3182,N_3873);
nor U5317 (N_5317,N_3372,N_3377);
xnor U5318 (N_5318,N_3943,N_4454);
nand U5319 (N_5319,N_4689,N_4292);
nor U5320 (N_5320,N_3927,N_2579);
xor U5321 (N_5321,N_3157,N_2848);
xnor U5322 (N_5322,N_4763,N_3208);
xor U5323 (N_5323,N_3958,N_4470);
xor U5324 (N_5324,N_4491,N_2559);
or U5325 (N_5325,N_2774,N_3563);
nand U5326 (N_5326,N_4329,N_2671);
nand U5327 (N_5327,N_4882,N_4109);
xnor U5328 (N_5328,N_4902,N_2582);
nand U5329 (N_5329,N_4250,N_3528);
or U5330 (N_5330,N_3971,N_4972);
nand U5331 (N_5331,N_4090,N_3124);
xor U5332 (N_5332,N_4720,N_2581);
or U5333 (N_5333,N_2798,N_4710);
xnor U5334 (N_5334,N_3820,N_3848);
nor U5335 (N_5335,N_2912,N_3851);
or U5336 (N_5336,N_3027,N_3463);
nand U5337 (N_5337,N_4091,N_2983);
and U5338 (N_5338,N_4851,N_4966);
xor U5339 (N_5339,N_2972,N_4508);
nor U5340 (N_5340,N_3053,N_4608);
or U5341 (N_5341,N_2997,N_3078);
or U5342 (N_5342,N_3834,N_2859);
xor U5343 (N_5343,N_3644,N_4903);
and U5344 (N_5344,N_3929,N_3779);
or U5345 (N_5345,N_3950,N_2638);
and U5346 (N_5346,N_3511,N_4561);
nand U5347 (N_5347,N_3916,N_4552);
or U5348 (N_5348,N_2505,N_2868);
and U5349 (N_5349,N_2574,N_3043);
and U5350 (N_5350,N_4366,N_4938);
nand U5351 (N_5351,N_4233,N_2751);
and U5352 (N_5352,N_3811,N_3945);
and U5353 (N_5353,N_4793,N_3214);
xnor U5354 (N_5354,N_3522,N_4367);
and U5355 (N_5355,N_3140,N_4458);
nor U5356 (N_5356,N_4796,N_3401);
nand U5357 (N_5357,N_4270,N_3765);
and U5358 (N_5358,N_3341,N_4886);
or U5359 (N_5359,N_3890,N_2799);
and U5360 (N_5360,N_3398,N_3451);
or U5361 (N_5361,N_2778,N_2520);
nor U5362 (N_5362,N_4149,N_4806);
and U5363 (N_5363,N_3361,N_3176);
and U5364 (N_5364,N_4800,N_2604);
and U5365 (N_5365,N_3007,N_3969);
and U5366 (N_5366,N_4045,N_2627);
or U5367 (N_5367,N_3531,N_3055);
and U5368 (N_5368,N_4859,N_4176);
xor U5369 (N_5369,N_4168,N_4979);
xnor U5370 (N_5370,N_3656,N_2958);
nor U5371 (N_5371,N_3680,N_4187);
nand U5372 (N_5372,N_4169,N_4598);
xor U5373 (N_5373,N_4687,N_4446);
nor U5374 (N_5374,N_3297,N_4614);
or U5375 (N_5375,N_3362,N_3099);
nand U5376 (N_5376,N_4542,N_2664);
nand U5377 (N_5377,N_4437,N_3258);
nor U5378 (N_5378,N_4729,N_3495);
xnor U5379 (N_5379,N_4128,N_4105);
nor U5380 (N_5380,N_4613,N_4786);
or U5381 (N_5381,N_4358,N_3716);
or U5382 (N_5382,N_4768,N_4711);
or U5383 (N_5383,N_3060,N_4140);
or U5384 (N_5384,N_2896,N_3520);
nand U5385 (N_5385,N_3223,N_4897);
xor U5386 (N_5386,N_4703,N_3045);
and U5387 (N_5387,N_3568,N_4416);
nand U5388 (N_5388,N_3496,N_4599);
and U5389 (N_5389,N_2878,N_3639);
and U5390 (N_5390,N_3222,N_3248);
or U5391 (N_5391,N_4662,N_4989);
or U5392 (N_5392,N_3960,N_4827);
nand U5393 (N_5393,N_3058,N_3276);
and U5394 (N_5394,N_3836,N_4836);
nor U5395 (N_5395,N_2901,N_4113);
nor U5396 (N_5396,N_4580,N_4129);
nand U5397 (N_5397,N_3197,N_4161);
nand U5398 (N_5398,N_4373,N_3289);
nand U5399 (N_5399,N_2991,N_2634);
nand U5400 (N_5400,N_4153,N_4391);
nand U5401 (N_5401,N_3414,N_3741);
or U5402 (N_5402,N_3893,N_4079);
and U5403 (N_5403,N_3739,N_2860);
xor U5404 (N_5404,N_2750,N_4318);
nor U5405 (N_5405,N_4987,N_3581);
and U5406 (N_5406,N_2818,N_2800);
nor U5407 (N_5407,N_3861,N_4393);
and U5408 (N_5408,N_3280,N_4259);
nor U5409 (N_5409,N_3162,N_4195);
xnor U5410 (N_5410,N_3714,N_4086);
nor U5411 (N_5411,N_4205,N_4003);
or U5412 (N_5412,N_4104,N_3204);
nand U5413 (N_5413,N_4731,N_3934);
and U5414 (N_5414,N_4727,N_4649);
or U5415 (N_5415,N_3881,N_3793);
or U5416 (N_5416,N_3949,N_4407);
and U5417 (N_5417,N_4967,N_4674);
xor U5418 (N_5418,N_4281,N_4138);
or U5419 (N_5419,N_4290,N_2644);
or U5420 (N_5420,N_3756,N_4170);
and U5421 (N_5421,N_4190,N_2701);
xnor U5422 (N_5422,N_3805,N_3234);
nor U5423 (N_5423,N_3307,N_4424);
nand U5424 (N_5424,N_3963,N_3655);
or U5425 (N_5425,N_3841,N_4435);
xnor U5426 (N_5426,N_3264,N_3186);
and U5427 (N_5427,N_3701,N_3606);
xor U5428 (N_5428,N_3493,N_3191);
nor U5429 (N_5429,N_4345,N_4950);
or U5430 (N_5430,N_3024,N_3849);
xnor U5431 (N_5431,N_3105,N_4087);
xnor U5432 (N_5432,N_3097,N_3106);
or U5433 (N_5433,N_4383,N_4505);
nand U5434 (N_5434,N_4146,N_3005);
xor U5435 (N_5435,N_2786,N_2616);
and U5436 (N_5436,N_3645,N_4893);
xor U5437 (N_5437,N_2956,N_2813);
and U5438 (N_5438,N_2944,N_4917);
nor U5439 (N_5439,N_4965,N_4442);
nand U5440 (N_5440,N_3886,N_3629);
nand U5441 (N_5441,N_2783,N_4436);
nor U5442 (N_5442,N_3220,N_4430);
xor U5443 (N_5443,N_4372,N_3230);
xor U5444 (N_5444,N_3555,N_3034);
or U5445 (N_5445,N_4022,N_4238);
xnor U5446 (N_5446,N_2894,N_4760);
and U5447 (N_5447,N_3102,N_3888);
and U5448 (N_5448,N_4709,N_3798);
xor U5449 (N_5449,N_3689,N_3390);
xnor U5450 (N_5450,N_3476,N_2715);
or U5451 (N_5451,N_2703,N_2613);
and U5452 (N_5452,N_4325,N_4455);
nor U5453 (N_5453,N_2807,N_3840);
nor U5454 (N_5454,N_2625,N_3954);
nor U5455 (N_5455,N_4402,N_4722);
or U5456 (N_5456,N_2552,N_4885);
and U5457 (N_5457,N_2999,N_4394);
nor U5458 (N_5458,N_3403,N_2917);
xor U5459 (N_5459,N_3219,N_4447);
and U5460 (N_5460,N_4425,N_3501);
and U5461 (N_5461,N_3518,N_4083);
and U5462 (N_5462,N_4804,N_4544);
xnor U5463 (N_5463,N_4767,N_2975);
nor U5464 (N_5464,N_3483,N_2587);
nand U5465 (N_5465,N_3351,N_3619);
nor U5466 (N_5466,N_4032,N_3441);
xor U5467 (N_5467,N_2516,N_2961);
nand U5468 (N_5468,N_4590,N_3940);
and U5469 (N_5469,N_4202,N_4230);
xnor U5470 (N_5470,N_3116,N_4256);
nand U5471 (N_5471,N_2729,N_3282);
nand U5472 (N_5472,N_2871,N_4907);
or U5473 (N_5473,N_4883,N_4920);
and U5474 (N_5474,N_3965,N_4002);
xor U5475 (N_5475,N_2570,N_3082);
xor U5476 (N_5476,N_3120,N_2594);
and U5477 (N_5477,N_2685,N_2672);
and U5478 (N_5478,N_4302,N_2826);
nand U5479 (N_5479,N_4656,N_4429);
or U5480 (N_5480,N_2829,N_4962);
and U5481 (N_5481,N_2887,N_4563);
nand U5482 (N_5482,N_3523,N_4363);
and U5483 (N_5483,N_4021,N_3679);
nor U5484 (N_5484,N_2655,N_2578);
nand U5485 (N_5485,N_4952,N_3659);
or U5486 (N_5486,N_3749,N_4007);
nand U5487 (N_5487,N_3667,N_4124);
xnor U5488 (N_5488,N_2642,N_3098);
nor U5489 (N_5489,N_3244,N_2749);
and U5490 (N_5490,N_4953,N_2988);
xnor U5491 (N_5491,N_3217,N_3897);
and U5492 (N_5492,N_2806,N_4260);
or U5493 (N_5493,N_4788,N_4672);
xor U5494 (N_5494,N_4792,N_3726);
and U5495 (N_5495,N_4881,N_4523);
or U5496 (N_5496,N_4494,N_2517);
nand U5497 (N_5497,N_4106,N_4201);
or U5498 (N_5498,N_4637,N_3492);
and U5499 (N_5499,N_3918,N_4065);
xor U5500 (N_5500,N_3311,N_3172);
xnor U5501 (N_5501,N_4975,N_4568);
and U5502 (N_5502,N_3478,N_2755);
nor U5503 (N_5503,N_4864,N_4677);
nand U5504 (N_5504,N_3901,N_3465);
nor U5505 (N_5505,N_3030,N_4970);
and U5506 (N_5506,N_3348,N_3961);
and U5507 (N_5507,N_2527,N_3239);
nor U5508 (N_5508,N_3226,N_3464);
or U5509 (N_5509,N_3776,N_3281);
and U5510 (N_5510,N_2657,N_3150);
xor U5511 (N_5511,N_3852,N_4157);
xnor U5512 (N_5512,N_3227,N_4018);
or U5513 (N_5513,N_3613,N_3972);
nor U5514 (N_5514,N_4665,N_4412);
xnor U5515 (N_5515,N_3304,N_4969);
xor U5516 (N_5516,N_2768,N_3259);
or U5517 (N_5517,N_2665,N_4719);
nand U5518 (N_5518,N_3183,N_3907);
xor U5519 (N_5519,N_3686,N_4216);
xor U5520 (N_5520,N_2891,N_2558);
nor U5521 (N_5521,N_4164,N_4012);
nor U5522 (N_5522,N_4670,N_2929);
nand U5523 (N_5523,N_3800,N_3326);
nand U5524 (N_5524,N_4348,N_3292);
or U5525 (N_5525,N_3405,N_4751);
xor U5526 (N_5526,N_2812,N_3481);
xnor U5527 (N_5527,N_4119,N_3734);
and U5528 (N_5528,N_3743,N_2640);
xnor U5529 (N_5529,N_4232,N_3365);
xor U5530 (N_5530,N_4809,N_4858);
and U5531 (N_5531,N_3580,N_2772);
nand U5532 (N_5532,N_4326,N_3672);
xor U5533 (N_5533,N_4116,N_4107);
nand U5534 (N_5534,N_4514,N_2756);
nor U5535 (N_5535,N_2924,N_3237);
or U5536 (N_5536,N_4775,N_3747);
nand U5537 (N_5537,N_4209,N_3394);
nand U5538 (N_5538,N_2609,N_3458);
and U5539 (N_5539,N_3166,N_4048);
nand U5540 (N_5540,N_4878,N_4546);
or U5541 (N_5541,N_4114,N_4840);
xnor U5542 (N_5542,N_2889,N_4601);
nor U5543 (N_5543,N_3062,N_4179);
and U5544 (N_5544,N_3330,N_4102);
xnor U5545 (N_5545,N_3042,N_4797);
nor U5546 (N_5546,N_4099,N_3845);
or U5547 (N_5547,N_3083,N_3525);
nor U5548 (N_5548,N_3869,N_3545);
nand U5549 (N_5549,N_3461,N_3114);
xor U5550 (N_5550,N_3383,N_4968);
and U5551 (N_5551,N_3285,N_3164);
nand U5552 (N_5552,N_4596,N_3913);
or U5553 (N_5553,N_3931,N_3272);
xnor U5554 (N_5554,N_4811,N_2809);
or U5555 (N_5555,N_3211,N_3814);
nand U5556 (N_5556,N_3470,N_4359);
nand U5557 (N_5557,N_2624,N_4680);
nand U5558 (N_5558,N_3169,N_2699);
xnor U5559 (N_5559,N_2884,N_3308);
and U5560 (N_5560,N_2707,N_3822);
or U5561 (N_5561,N_4923,N_3036);
or U5562 (N_5562,N_4887,N_2593);
and U5563 (N_5563,N_4721,N_2632);
xor U5564 (N_5564,N_3179,N_3902);
nor U5565 (N_5565,N_3827,N_3571);
and U5566 (N_5566,N_2810,N_3294);
nor U5567 (N_5567,N_4855,N_4757);
or U5568 (N_5568,N_2631,N_3761);
nor U5569 (N_5569,N_3657,N_2904);
or U5570 (N_5570,N_2547,N_3433);
nor U5571 (N_5571,N_3682,N_3611);
xor U5572 (N_5572,N_4741,N_2575);
and U5573 (N_5573,N_4298,N_3061);
or U5574 (N_5574,N_2796,N_2840);
xor U5575 (N_5575,N_2612,N_3690);
or U5576 (N_5576,N_2954,N_2838);
and U5577 (N_5577,N_3436,N_3000);
nand U5578 (N_5578,N_3144,N_3728);
nand U5579 (N_5579,N_4871,N_3725);
xor U5580 (N_5580,N_3445,N_3334);
xnor U5581 (N_5581,N_4185,N_4654);
and U5582 (N_5582,N_2537,N_4616);
nand U5583 (N_5583,N_4061,N_2758);
nand U5584 (N_5584,N_3795,N_3295);
and U5585 (N_5585,N_3723,N_3462);
nor U5586 (N_5586,N_2569,N_4789);
or U5587 (N_5587,N_4626,N_2539);
xnor U5588 (N_5588,N_4640,N_3442);
xnor U5589 (N_5589,N_2819,N_4080);
nand U5590 (N_5590,N_4336,N_4629);
xor U5591 (N_5591,N_4276,N_3152);
xnor U5592 (N_5592,N_3335,N_4976);
nor U5593 (N_5593,N_4374,N_4163);
nor U5594 (N_5594,N_4773,N_3503);
nor U5595 (N_5595,N_3324,N_2754);
nor U5596 (N_5596,N_4648,N_4068);
or U5597 (N_5597,N_2507,N_4700);
and U5598 (N_5598,N_4600,N_4311);
nor U5599 (N_5599,N_3534,N_3328);
or U5600 (N_5600,N_4867,N_4186);
or U5601 (N_5601,N_3126,N_4432);
nor U5602 (N_5602,N_4142,N_4581);
nand U5603 (N_5603,N_3813,N_3506);
or U5604 (N_5604,N_3906,N_3332);
xnor U5605 (N_5605,N_4625,N_3770);
xor U5606 (N_5606,N_3215,N_4019);
nor U5607 (N_5607,N_2560,N_4604);
nor U5608 (N_5608,N_4139,N_4268);
xor U5609 (N_5609,N_3268,N_4527);
nand U5610 (N_5610,N_3212,N_2773);
xor U5611 (N_5611,N_3885,N_3706);
nor U5612 (N_5612,N_2586,N_4752);
xor U5613 (N_5613,N_3283,N_3257);
or U5614 (N_5614,N_4386,N_3113);
xor U5615 (N_5615,N_4631,N_4802);
and U5616 (N_5616,N_4866,N_4127);
nor U5617 (N_5617,N_4258,N_4467);
or U5618 (N_5618,N_4264,N_3320);
nand U5619 (N_5619,N_3064,N_2681);
and U5620 (N_5620,N_2564,N_4085);
or U5621 (N_5621,N_4556,N_2725);
or U5622 (N_5622,N_2704,N_4666);
nor U5623 (N_5623,N_3346,N_3380);
nor U5624 (N_5624,N_4790,N_2525);
nand U5625 (N_5625,N_3551,N_3512);
or U5626 (N_5626,N_2797,N_2545);
nor U5627 (N_5627,N_4449,N_4759);
xnor U5628 (N_5628,N_4991,N_3333);
nor U5629 (N_5629,N_3588,N_2649);
nand U5630 (N_5630,N_4076,N_4597);
nor U5631 (N_5631,N_4838,N_3499);
nor U5632 (N_5632,N_3517,N_2551);
and U5633 (N_5633,N_2792,N_3021);
nor U5634 (N_5634,N_3705,N_3086);
nand U5635 (N_5635,N_3871,N_4451);
nand U5636 (N_5636,N_3118,N_2503);
or U5637 (N_5637,N_2605,N_4622);
nor U5638 (N_5638,N_4155,N_2504);
and U5639 (N_5639,N_4650,N_3758);
xnor U5640 (N_5640,N_4842,N_4942);
nor U5641 (N_5641,N_4573,N_3123);
or U5642 (N_5642,N_4780,N_4567);
or U5643 (N_5643,N_4468,N_4289);
nand U5644 (N_5644,N_3558,N_3161);
xor U5645 (N_5645,N_4538,N_4647);
xnor U5646 (N_5646,N_4844,N_2735);
or U5647 (N_5647,N_2874,N_3020);
nor U5648 (N_5648,N_2963,N_3096);
or U5649 (N_5649,N_3001,N_3068);
nand U5650 (N_5650,N_3111,N_4794);
xor U5651 (N_5651,N_2731,N_4837);
or U5652 (N_5652,N_4073,N_3033);
nor U5653 (N_5653,N_3694,N_2855);
nor U5654 (N_5654,N_2787,N_3091);
or U5655 (N_5655,N_4141,N_3553);
and U5656 (N_5656,N_4500,N_2764);
or U5657 (N_5657,N_4764,N_3766);
nor U5658 (N_5658,N_2937,N_4226);
nand U5659 (N_5659,N_4343,N_3951);
or U5660 (N_5660,N_2981,N_4933);
xnor U5661 (N_5661,N_4001,N_3142);
xnor U5662 (N_5662,N_4634,N_2854);
xnor U5663 (N_5663,N_2795,N_4247);
xor U5664 (N_5664,N_4122,N_4930);
nand U5665 (N_5665,N_4253,N_2775);
and U5666 (N_5666,N_3100,N_3104);
or U5667 (N_5667,N_2875,N_2763);
and U5668 (N_5668,N_3648,N_3596);
or U5669 (N_5669,N_2953,N_4526);
nor U5670 (N_5670,N_2876,N_2647);
or U5671 (N_5671,N_2633,N_4685);
or U5672 (N_5672,N_2682,N_4615);
or U5673 (N_5673,N_2747,N_3985);
or U5674 (N_5674,N_2960,N_2702);
nor U5675 (N_5675,N_4215,N_2680);
nand U5676 (N_5676,N_2554,N_3953);
xnor U5677 (N_5677,N_4100,N_2622);
nor U5678 (N_5678,N_4949,N_4815);
nor U5679 (N_5679,N_3149,N_3494);
nor U5680 (N_5680,N_3029,N_4589);
and U5681 (N_5681,N_3597,N_2951);
nand U5682 (N_5682,N_3079,N_2666);
and U5683 (N_5683,N_2522,N_3305);
or U5684 (N_5684,N_4385,N_3115);
or U5685 (N_5685,N_4605,N_3598);
or U5686 (N_5686,N_3107,N_4973);
and U5687 (N_5687,N_4278,N_3738);
nor U5688 (N_5688,N_2916,N_4696);
and U5689 (N_5689,N_2675,N_4704);
and U5690 (N_5690,N_4095,N_4623);
nor U5691 (N_5691,N_4017,N_4377);
nor U5692 (N_5692,N_3290,N_3977);
nand U5693 (N_5693,N_2837,N_4694);
nor U5694 (N_5694,N_2949,N_2836);
nand U5695 (N_5695,N_3948,N_4583);
nor U5696 (N_5696,N_4287,N_4263);
nand U5697 (N_5697,N_4777,N_3420);
and U5698 (N_5698,N_2880,N_2918);
and U5699 (N_5699,N_4052,N_3660);
nor U5700 (N_5700,N_4093,N_3540);
nor U5701 (N_5701,N_4619,N_4684);
xor U5702 (N_5702,N_4916,N_2670);
or U5703 (N_5703,N_2746,N_4522);
nand U5704 (N_5704,N_4813,N_2928);
xor U5705 (N_5705,N_3093,N_4705);
xor U5706 (N_5706,N_3837,N_3240);
and U5707 (N_5707,N_3252,N_3624);
nor U5708 (N_5708,N_4594,N_3067);
nor U5709 (N_5709,N_4932,N_3128);
and U5710 (N_5710,N_3767,N_4286);
and U5711 (N_5711,N_3048,N_4776);
xnor U5712 (N_5712,N_2663,N_3336);
nand U5713 (N_5713,N_4341,N_4115);
nand U5714 (N_5714,N_4734,N_3786);
and U5715 (N_5715,N_4495,N_2711);
or U5716 (N_5716,N_2636,N_3329);
and U5717 (N_5717,N_4565,N_4756);
and U5718 (N_5718,N_4832,N_2903);
xor U5719 (N_5719,N_3249,N_4828);
nor U5720 (N_5720,N_3590,N_3752);
xor U5721 (N_5721,N_2553,N_3411);
nand U5722 (N_5722,N_4915,N_2742);
or U5723 (N_5723,N_4165,N_2959);
and U5724 (N_5724,N_3631,N_3883);
nor U5725 (N_5725,N_3762,N_3018);
or U5726 (N_5726,N_3262,N_4148);
and U5727 (N_5727,N_3360,N_3973);
nand U5728 (N_5728,N_3699,N_2914);
or U5729 (N_5729,N_2890,N_3147);
nand U5730 (N_5730,N_4779,N_3340);
and U5731 (N_5731,N_4698,N_3318);
xnor U5732 (N_5732,N_4639,N_2921);
or U5733 (N_5733,N_3466,N_3832);
xnor U5734 (N_5734,N_4512,N_4008);
and U5735 (N_5735,N_4303,N_3550);
and U5736 (N_5736,N_4231,N_3391);
nand U5737 (N_5737,N_3880,N_4399);
xnor U5738 (N_5738,N_3987,N_2900);
nand U5739 (N_5739,N_3976,N_2523);
nand U5740 (N_5740,N_2650,N_4877);
xnor U5741 (N_5741,N_2957,N_3651);
nor U5742 (N_5742,N_3108,N_4929);
xor U5743 (N_5743,N_2568,N_3889);
or U5744 (N_5744,N_4519,N_4466);
xnor U5745 (N_5745,N_2733,N_2641);
xor U5746 (N_5746,N_2629,N_2591);
xnor U5747 (N_5747,N_3768,N_3287);
or U5748 (N_5748,N_4319,N_4181);
or U5749 (N_5749,N_2606,N_2817);
or U5750 (N_5750,N_3242,N_4400);
nand U5751 (N_5751,N_2583,N_3131);
or U5752 (N_5752,N_3993,N_3921);
xnor U5753 (N_5753,N_4211,N_4027);
nand U5754 (N_5754,N_4255,N_4267);
or U5755 (N_5755,N_4520,N_4826);
nor U5756 (N_5756,N_3469,N_2842);
or U5757 (N_5757,N_4557,N_4843);
xor U5758 (N_5758,N_4239,N_4957);
nand U5759 (N_5759,N_4484,N_3879);
nand U5760 (N_5760,N_4307,N_4327);
and U5761 (N_5761,N_4820,N_4769);
or U5762 (N_5762,N_3895,N_3173);
and U5763 (N_5763,N_4579,N_3011);
xnor U5764 (N_5764,N_3177,N_4934);
or U5765 (N_5765,N_3314,N_4354);
and U5766 (N_5766,N_4118,N_3207);
xor U5767 (N_5767,N_4041,N_3847);
nor U5768 (N_5768,N_3962,N_3830);
or U5769 (N_5769,N_2982,N_4997);
nor U5770 (N_5770,N_3135,N_3905);
and U5771 (N_5771,N_3844,N_3891);
xnor U5772 (N_5772,N_4280,N_3868);
and U5773 (N_5773,N_3541,N_4676);
and U5774 (N_5774,N_3729,N_4418);
or U5775 (N_5775,N_3475,N_2865);
or U5776 (N_5776,N_3382,N_4860);
or U5777 (N_5777,N_4754,N_4761);
nand U5778 (N_5778,N_4633,N_4452);
xor U5779 (N_5779,N_3339,N_3663);
and U5780 (N_5780,N_3138,N_4217);
xor U5781 (N_5781,N_2567,N_2695);
xnor U5782 (N_5782,N_3980,N_2684);
nand U5783 (N_5783,N_2676,N_3623);
or U5784 (N_5784,N_4603,N_3132);
and U5785 (N_5785,N_3939,N_3778);
nor U5786 (N_5786,N_3618,N_4396);
and U5787 (N_5787,N_4166,N_3129);
or U5788 (N_5788,N_3153,N_3452);
nor U5789 (N_5789,N_4010,N_4055);
nand U5790 (N_5790,N_4413,N_2993);
and U5791 (N_5791,N_4035,N_3603);
or U5792 (N_5792,N_4845,N_3256);
nand U5793 (N_5793,N_4026,N_3467);
nand U5794 (N_5794,N_4986,N_4474);
and U5795 (N_5795,N_3171,N_3225);
nor U5796 (N_5796,N_3559,N_3073);
and U5797 (N_5797,N_3070,N_4834);
and U5798 (N_5798,N_4338,N_3180);
nor U5799 (N_5799,N_3796,N_3238);
and U5800 (N_5800,N_4053,N_3854);
nand U5801 (N_5801,N_3110,N_3567);
or U5802 (N_5802,N_3407,N_2708);
or U5803 (N_5803,N_4421,N_3996);
nor U5804 (N_5804,N_4056,N_4011);
or U5805 (N_5805,N_4316,N_4980);
nand U5806 (N_5806,N_4958,N_2844);
xnor U5807 (N_5807,N_3850,N_4857);
or U5808 (N_5808,N_4241,N_3066);
nor U5809 (N_5809,N_3685,N_3385);
nand U5810 (N_5810,N_3431,N_4020);
nor U5811 (N_5811,N_2879,N_4679);
and U5812 (N_5812,N_4369,N_4192);
or U5813 (N_5813,N_3424,N_3439);
or U5814 (N_5814,N_4692,N_4558);
and U5815 (N_5815,N_3218,N_4954);
or U5816 (N_5816,N_4269,N_3359);
and U5817 (N_5817,N_3277,N_3253);
and U5818 (N_5818,N_3396,N_4360);
xor U5819 (N_5819,N_4805,N_4925);
xor U5820 (N_5820,N_4444,N_4632);
xor U5821 (N_5821,N_3137,N_4453);
nor U5822 (N_5822,N_3717,N_4074);
nand U5823 (N_5823,N_4434,N_2923);
and U5824 (N_5824,N_4151,N_4560);
and U5825 (N_5825,N_4990,N_3275);
nor U5826 (N_5826,N_4525,N_2706);
nand U5827 (N_5827,N_4332,N_3633);
xor U5828 (N_5828,N_2646,N_2714);
and U5829 (N_5829,N_4824,N_4047);
or U5830 (N_5830,N_3543,N_3418);
nor U5831 (N_5831,N_4550,N_3509);
nor U5832 (N_5832,N_2816,N_3039);
and U5833 (N_5833,N_4376,N_2577);
nand U5834 (N_5834,N_2697,N_4040);
nand U5835 (N_5835,N_3578,N_3221);
and U5836 (N_5836,N_3319,N_4337);
nand U5837 (N_5837,N_4541,N_3006);
or U5838 (N_5838,N_3533,N_4900);
and U5839 (N_5839,N_3938,N_2526);
and U5840 (N_5840,N_3288,N_3159);
nand U5841 (N_5841,N_4257,N_4433);
and U5842 (N_5842,N_3676,N_4335);
nor U5843 (N_5843,N_4993,N_4636);
xor U5844 (N_5844,N_3154,N_2930);
xnor U5845 (N_5845,N_3920,N_4940);
nand U5846 (N_5846,N_4228,N_3373);
xnor U5847 (N_5847,N_2713,N_4315);
or U5848 (N_5848,N_3936,N_4297);
and U5849 (N_5849,N_2659,N_2556);
or U5850 (N_5850,N_3388,N_3665);
xor U5851 (N_5851,N_2834,N_4248);
and U5852 (N_5852,N_4098,N_4688);
nor U5853 (N_5853,N_4251,N_4895);
or U5854 (N_5854,N_2617,N_2691);
xor U5855 (N_5855,N_4869,N_2543);
and U5856 (N_5856,N_3989,N_4511);
or U5857 (N_5857,N_4941,N_3978);
or U5858 (N_5858,N_4668,N_4643);
or U5859 (N_5859,N_2531,N_4852);
nand U5860 (N_5860,N_4661,N_4482);
or U5861 (N_5861,N_4762,N_4863);
and U5862 (N_5862,N_4060,N_3194);
or U5863 (N_5863,N_2830,N_3056);
xor U5864 (N_5864,N_3703,N_3299);
nand U5865 (N_5865,N_4194,N_3605);
xor U5866 (N_5866,N_2615,N_3247);
and U5867 (N_5867,N_3387,N_2585);
xor U5868 (N_5868,N_3155,N_4441);
and U5869 (N_5869,N_2540,N_4382);
and U5870 (N_5870,N_3823,N_4245);
xnor U5871 (N_5871,N_4723,N_4064);
nand U5872 (N_5872,N_3188,N_3678);
or U5873 (N_5873,N_4072,N_4798);
nand U5874 (N_5874,N_3556,N_4948);
and U5875 (N_5875,N_3023,N_4988);
or U5876 (N_5876,N_2850,N_4861);
and U5877 (N_5877,N_2710,N_4092);
nand U5878 (N_5878,N_3456,N_2978);
nor U5879 (N_5879,N_3417,N_4931);
nand U5880 (N_5880,N_3101,N_3911);
nor U5881 (N_5881,N_3892,N_3274);
xor U5882 (N_5882,N_4712,N_4908);
or U5883 (N_5883,N_2512,N_4981);
nor U5884 (N_5884,N_4355,N_4535);
or U5885 (N_5885,N_4312,N_4150);
and U5886 (N_5886,N_3974,N_4956);
and U5887 (N_5887,N_3794,N_4381);
xor U5888 (N_5888,N_2828,N_3926);
nor U5889 (N_5889,N_4137,N_4644);
and U5890 (N_5890,N_2920,N_4707);
or U5891 (N_5891,N_4714,N_4293);
nand U5892 (N_5892,N_2611,N_4982);
and U5893 (N_5893,N_2588,N_2992);
and U5894 (N_5894,N_4663,N_3736);
and U5895 (N_5895,N_4183,N_3313);
nand U5896 (N_5896,N_4726,N_3865);
nand U5897 (N_5897,N_4884,N_4936);
or U5898 (N_5898,N_3984,N_4778);
xnor U5899 (N_5899,N_3652,N_2536);
and U5900 (N_5900,N_3010,N_3413);
xnor U5901 (N_5901,N_3923,N_3742);
or U5902 (N_5902,N_2781,N_3816);
xor U5903 (N_5903,N_4054,N_4992);
nor U5904 (N_5904,N_3826,N_4529);
xor U5905 (N_5905,N_3866,N_2645);
nor U5906 (N_5906,N_4708,N_4351);
or U5907 (N_5907,N_2598,N_3666);
nand U5908 (N_5908,N_4846,N_4740);
or U5909 (N_5909,N_2757,N_3031);
and U5910 (N_5910,N_4380,N_3489);
or U5911 (N_5911,N_4333,N_2743);
xor U5912 (N_5912,N_4101,N_3942);
or U5913 (N_5913,N_4344,N_3658);
xor U5914 (N_5914,N_4234,N_4123);
and U5915 (N_5915,N_2791,N_2906);
and U5916 (N_5916,N_3909,N_4746);
nor U5917 (N_5917,N_3145,N_3641);
nor U5918 (N_5918,N_3757,N_4145);
or U5919 (N_5919,N_2895,N_3125);
xor U5920 (N_5920,N_4126,N_4219);
and U5921 (N_5921,N_4134,N_2573);
xnor U5922 (N_5922,N_3621,N_4999);
nand U5923 (N_5923,N_4197,N_4803);
nor U5924 (N_5924,N_4049,N_3812);
and U5925 (N_5925,N_4947,N_4724);
xor U5926 (N_5926,N_3019,N_4483);
xnor U5927 (N_5927,N_4945,N_3175);
xnor U5928 (N_5928,N_3932,N_4236);
nor U5929 (N_5929,N_3899,N_4770);
and U5930 (N_5930,N_3141,N_4143);
nand U5931 (N_5931,N_3459,N_3784);
nor U5932 (N_5932,N_2719,N_4899);
or U5933 (N_5933,N_4515,N_3293);
nor U5934 (N_5934,N_3988,N_2620);
or U5935 (N_5935,N_3576,N_2909);
or U5936 (N_5936,N_3072,N_4097);
nand U5937 (N_5937,N_4620,N_3504);
and U5938 (N_5938,N_4423,N_4588);
nand U5939 (N_5939,N_2995,N_3858);
nor U5940 (N_5940,N_3317,N_2603);
nand U5941 (N_5941,N_4282,N_3780);
or U5942 (N_5942,N_3979,N_4462);
nand U5943 (N_5943,N_3399,N_3640);
or U5944 (N_5944,N_3529,N_4044);
xnor U5945 (N_5945,N_2678,N_3877);
or U5946 (N_5946,N_4235,N_3265);
xor U5947 (N_5947,N_3654,N_4029);
xor U5948 (N_5948,N_2688,N_2610);
xor U5949 (N_5949,N_4513,N_4875);
nand U5950 (N_5950,N_3119,N_2709);
xor U5951 (N_5951,N_3345,N_4960);
nor U5952 (N_5952,N_3825,N_3017);
nand U5953 (N_5953,N_3121,N_2571);
nand U5954 (N_5954,N_2857,N_3783);
nand U5955 (N_5955,N_4254,N_4320);
or U5956 (N_5956,N_4162,N_2908);
or U5957 (N_5957,N_3224,N_4184);
and U5958 (N_5958,N_3229,N_4901);
or U5959 (N_5959,N_4025,N_4532);
nand U5960 (N_5960,N_3085,N_4388);
or U5961 (N_5961,N_3447,N_4554);
nand U5962 (N_5962,N_4242,N_2528);
xor U5963 (N_5963,N_4488,N_3700);
and U5964 (N_5964,N_4744,N_2546);
or U5965 (N_5965,N_3415,N_2643);
xor U5966 (N_5966,N_4227,N_3908);
nor U5967 (N_5967,N_3054,N_2841);
nand U5968 (N_5968,N_2595,N_3352);
nor U5969 (N_5969,N_4628,N_3810);
or U5970 (N_5970,N_4006,N_3691);
or U5971 (N_5971,N_2862,N_4497);
or U5972 (N_5972,N_3192,N_4506);
and U5973 (N_5973,N_3200,N_3080);
xor U5974 (N_5974,N_2674,N_4352);
or U5975 (N_5975,N_4856,N_3632);
xor U5976 (N_5976,N_2753,N_4935);
xor U5977 (N_5977,N_3347,N_3315);
and U5978 (N_5978,N_4819,N_4347);
or U5979 (N_5979,N_2911,N_2892);
and U5980 (N_5980,N_3946,N_3502);
or U5981 (N_5981,N_2686,N_3381);
nor U5982 (N_5982,N_2934,N_4469);
nor U5983 (N_5983,N_3804,N_3508);
xor U5984 (N_5984,N_4974,N_3148);
and U5985 (N_5985,N_4749,N_2765);
and U5986 (N_5986,N_3013,N_4671);
or U5987 (N_5987,N_2741,N_3206);
or U5988 (N_5988,N_3170,N_3807);
nor U5989 (N_5989,N_2652,N_4252);
xor U5990 (N_5990,N_3982,N_4182);
and U5991 (N_5991,N_2808,N_2811);
and U5992 (N_5992,N_2561,N_2965);
nor U5993 (N_5993,N_3269,N_4914);
and U5994 (N_5994,N_4310,N_3860);
xor U5995 (N_5995,N_4755,N_3627);
nor U5996 (N_5996,N_2544,N_3763);
or U5997 (N_5997,N_3746,N_4651);
nand U5998 (N_5998,N_3112,N_4658);
xnor U5999 (N_5999,N_3038,N_2548);
xor U6000 (N_6000,N_3434,N_2607);
nor U6001 (N_6001,N_3930,N_3608);
nor U6002 (N_6002,N_4398,N_4225);
and U6003 (N_6003,N_4509,N_4346);
nand U6004 (N_6004,N_4955,N_4160);
and U6005 (N_6005,N_4342,N_4591);
and U6006 (N_6006,N_3163,N_3358);
nor U6007 (N_6007,N_3412,N_3801);
or U6008 (N_6008,N_4308,N_3284);
and U6009 (N_6009,N_4772,N_3350);
nand U6010 (N_6010,N_2966,N_4739);
nor U6011 (N_6011,N_4172,N_3077);
nor U6012 (N_6012,N_3549,N_4611);
xor U6013 (N_6013,N_3250,N_2500);
nor U6014 (N_6014,N_3485,N_4578);
xor U6015 (N_6015,N_2985,N_2967);
and U6016 (N_6016,N_4350,N_2938);
xor U6017 (N_6017,N_2614,N_3379);
nor U6018 (N_6018,N_3455,N_3375);
nor U6019 (N_6019,N_4198,N_2872);
and U6020 (N_6020,N_2599,N_2654);
and U6021 (N_6021,N_3189,N_2863);
nor U6022 (N_6022,N_3008,N_2955);
and U6023 (N_6023,N_3829,N_4321);
xnor U6024 (N_6024,N_4023,N_3429);
and U6025 (N_6025,N_4528,N_4371);
nor U6026 (N_6026,N_3232,N_2998);
or U6027 (N_6027,N_4702,N_4220);
or U6028 (N_6028,N_4894,N_3602);
nand U6029 (N_6029,N_3190,N_3966);
nand U6030 (N_6030,N_3697,N_4411);
xnor U6031 (N_6031,N_4713,N_4057);
and U6032 (N_6032,N_3201,N_3626);
and U6033 (N_6033,N_4478,N_3370);
xor U6034 (N_6034,N_4370,N_3122);
nand U6035 (N_6035,N_3724,N_4243);
or U6036 (N_6036,N_3422,N_3681);
xnor U6037 (N_6037,N_3427,N_2769);
nor U6038 (N_6038,N_3514,N_3867);
nor U6039 (N_6039,N_3589,N_3472);
nand U6040 (N_6040,N_4584,N_4089);
and U6041 (N_6041,N_3074,N_4681);
nor U6042 (N_6042,N_3732,N_3440);
and U6043 (N_6043,N_4905,N_2555);
and U6044 (N_6044,N_4174,N_3435);
nor U6045 (N_6045,N_4766,N_2947);
and U6046 (N_6046,N_4328,N_4808);
or U6047 (N_6047,N_4521,N_3321);
nand U6048 (N_6048,N_4059,N_2683);
nand U6049 (N_6049,N_4876,N_4890);
or U6050 (N_6050,N_3799,N_3454);
xnor U6051 (N_6051,N_4214,N_2910);
nor U6052 (N_6052,N_2941,N_3354);
nor U6053 (N_6053,N_3423,N_4490);
and U6054 (N_6054,N_4978,N_2721);
nor U6055 (N_6055,N_3855,N_3168);
or U6056 (N_6056,N_2831,N_2897);
or U6057 (N_6057,N_2869,N_3028);
xnor U6058 (N_6058,N_3181,N_3719);
or U6059 (N_6059,N_4924,N_3642);
xnor U6060 (N_6060,N_4322,N_3460);
nor U6061 (N_6061,N_3887,N_3051);
xnor U6062 (N_6062,N_3959,N_3366);
nor U6063 (N_6063,N_4983,N_4536);
nand U6064 (N_6064,N_4295,N_3737);
or U6065 (N_6065,N_3271,N_4592);
nand U6066 (N_6066,N_4717,N_2893);
xnor U6067 (N_6067,N_3047,N_3876);
nand U6068 (N_6068,N_4317,N_3894);
and U6069 (N_6069,N_4785,N_3662);
nor U6070 (N_6070,N_4502,N_2535);
xnor U6071 (N_6071,N_2950,N_2820);
xor U6072 (N_6072,N_4503,N_2861);
and U6073 (N_6073,N_2886,N_3649);
and U6074 (N_6074,N_4564,N_3368);
xnor U6075 (N_6075,N_2565,N_2589);
nor U6076 (N_6076,N_3088,N_2927);
and U6077 (N_6077,N_4880,N_4479);
or U6078 (N_6078,N_4167,N_3355);
nand U6079 (N_6079,N_4152,N_3815);
nand U6080 (N_6080,N_4607,N_4787);
or U6081 (N_6081,N_2530,N_3474);
xnor U6082 (N_6082,N_4050,N_3254);
or U6083 (N_6083,N_3488,N_3513);
nand U6084 (N_6084,N_3900,N_3862);
xnor U6085 (N_6085,N_3037,N_2532);
xnor U6086 (N_6086,N_2501,N_3718);
xor U6087 (N_6087,N_3637,N_3202);
and U6088 (N_6088,N_2994,N_4299);
and U6089 (N_6089,N_4212,N_3185);
and U6090 (N_6090,N_3671,N_4409);
nor U6091 (N_6091,N_4833,N_4014);
or U6092 (N_6092,N_4874,N_4870);
or U6093 (N_6093,N_2821,N_4630);
or U6094 (N_6094,N_4237,N_4144);
xor U6095 (N_6095,N_4667,N_4533);
or U6096 (N_6096,N_3302,N_4203);
and U6097 (N_6097,N_2557,N_4586);
nand U6098 (N_6098,N_2843,N_3884);
or U6099 (N_6099,N_4445,N_4501);
and U6100 (N_6100,N_3552,N_3400);
nor U6101 (N_6101,N_3448,N_3797);
and U6102 (N_6102,N_4364,N_4812);
nor U6103 (N_6103,N_3684,N_4213);
and U6104 (N_6104,N_3677,N_2939);
or U6105 (N_6105,N_3872,N_3364);
and U6106 (N_6106,N_2789,N_3084);
xor U6107 (N_6107,N_2508,N_4627);
or U6108 (N_6108,N_3748,N_3089);
nor U6109 (N_6109,N_4427,N_3539);
nor U6110 (N_6110,N_4995,N_3817);
nor U6111 (N_6111,N_3530,N_4353);
nand U6112 (N_6112,N_4042,N_4922);
xnor U6113 (N_6113,N_2744,N_4732);
nand U6114 (N_6114,N_3586,N_3143);
and U6115 (N_6115,N_4807,N_4189);
nor U6116 (N_6116,N_4378,N_2563);
xnor U6117 (N_6117,N_2502,N_4481);
nor U6118 (N_6118,N_2696,N_2933);
nand U6119 (N_6119,N_4200,N_4009);
xnor U6120 (N_6120,N_4697,N_4193);
or U6121 (N_6121,N_3673,N_3012);
nor U6122 (N_6122,N_3583,N_4024);
nor U6123 (N_6123,N_4273,N_3709);
or U6124 (N_6124,N_4130,N_3095);
xor U6125 (N_6125,N_4574,N_2550);
and U6126 (N_6126,N_4066,N_4471);
xnor U6127 (N_6127,N_4765,N_3312);
xnor U6128 (N_6128,N_4489,N_4659);
or U6129 (N_6129,N_3983,N_3389);
and U6130 (N_6130,N_3278,N_4618);
or U6131 (N_6131,N_2667,N_4368);
nand U6132 (N_6132,N_4387,N_4758);
nand U6133 (N_6133,N_4822,N_4334);
and U6134 (N_6134,N_2533,N_2519);
or U6135 (N_6135,N_2745,N_3273);
nor U6136 (N_6136,N_3009,N_3607);
xor U6137 (N_6137,N_2700,N_3573);
or U6138 (N_6138,N_2776,N_4171);
nand U6139 (N_6139,N_3526,N_2770);
nor U6140 (N_6140,N_3016,N_3343);
and U6141 (N_6141,N_2866,N_4362);
nand U6142 (N_6142,N_4610,N_4549);
nor U6143 (N_6143,N_4745,N_3482);
or U6144 (N_6144,N_4911,N_4835);
or U6145 (N_6145,N_4868,N_4067);
nor U6146 (N_6146,N_4576,N_3331);
and U6147 (N_6147,N_3670,N_3059);
or U6148 (N_6148,N_3863,N_3127);
xor U6149 (N_6149,N_4737,N_3453);
or U6150 (N_6150,N_2962,N_2948);
nand U6151 (N_6151,N_3557,N_4324);
nor U6152 (N_6152,N_2932,N_4361);
nand U6153 (N_6153,N_3635,N_3643);
xor U6154 (N_6154,N_4888,N_3203);
nor U6155 (N_6155,N_4946,N_2542);
xor U6156 (N_6156,N_4683,N_4173);
or U6157 (N_6157,N_3486,N_4404);
or U6158 (N_6158,N_3174,N_2716);
nor U6159 (N_6159,N_4718,N_2529);
xnor U6160 (N_6160,N_2524,N_4898);
nand U6161 (N_6161,N_3896,N_3788);
and U6162 (N_6162,N_2784,N_4365);
xnor U6163 (N_6163,N_4408,N_2514);
nand U6164 (N_6164,N_3727,N_2694);
nor U6165 (N_6165,N_4473,N_4939);
or U6166 (N_6166,N_4602,N_3052);
or U6167 (N_6167,N_3081,N_3994);
and U6168 (N_6168,N_3327,N_3750);
nand U6169 (N_6169,N_4401,N_4262);
or U6170 (N_6170,N_2771,N_3818);
or U6171 (N_6171,N_2639,N_3371);
and U6172 (N_6172,N_4069,N_3500);
xor U6173 (N_6173,N_2825,N_3986);
nor U6174 (N_6174,N_3614,N_3789);
or U6175 (N_6175,N_4784,N_3616);
nor U6176 (N_6176,N_3759,N_3646);
nor U6177 (N_6177,N_4188,N_3196);
or U6178 (N_6178,N_2732,N_4829);
and U6179 (N_6179,N_3065,N_4545);
and U6180 (N_6180,N_2736,N_2648);
nor U6181 (N_6181,N_2669,N_2852);
xnor U6182 (N_6182,N_2952,N_2823);
nand U6183 (N_6183,N_3524,N_4135);
nor U6184 (N_6184,N_2996,N_2601);
and U6185 (N_6185,N_3730,N_3406);
nor U6186 (N_6186,N_3076,N_3821);
nor U6187 (N_6187,N_2698,N_3864);
or U6188 (N_6188,N_4279,N_2572);
and U6189 (N_6189,N_4609,N_4420);
nand U6190 (N_6190,N_3843,N_4918);
nand U6191 (N_6191,N_3914,N_4210);
or U6192 (N_6192,N_3612,N_4695);
and U6193 (N_6193,N_3025,N_2867);
and U6194 (N_6194,N_2803,N_4817);
and U6195 (N_6195,N_4963,N_3376);
xor U6196 (N_6196,N_3397,N_4275);
xor U6197 (N_6197,N_3785,N_2973);
nand U6198 (N_6198,N_3386,N_2827);
or U6199 (N_6199,N_4499,N_3764);
xor U6200 (N_6200,N_2549,N_4818);
or U6201 (N_6201,N_3022,N_2913);
xnor U6202 (N_6202,N_2970,N_2971);
nor U6203 (N_6203,N_4406,N_3117);
and U6204 (N_6204,N_2727,N_4699);
or U6205 (N_6205,N_4439,N_2835);
nor U6206 (N_6206,N_3356,N_4791);
nor U6207 (N_6207,N_3279,N_4156);
nand U6208 (N_6208,N_4782,N_3243);
or U6209 (N_6209,N_2888,N_3944);
nor U6210 (N_6210,N_4147,N_2814);
nor U6211 (N_6211,N_4178,N_4154);
xnor U6212 (N_6212,N_4246,N_4569);
and U6213 (N_6213,N_2661,N_4283);
nor U6214 (N_6214,N_3928,N_3075);
nand U6215 (N_6215,N_4291,N_4865);
nor U6216 (N_6216,N_3947,N_2662);
xor U6217 (N_6217,N_4426,N_3593);
nor U6218 (N_6218,N_4379,N_4103);
and U6219 (N_6219,N_3446,N_4540);
nand U6220 (N_6220,N_2626,N_4524);
or U6221 (N_6221,N_3521,N_4653);
xor U6222 (N_6222,N_4646,N_2846);
or U6223 (N_6223,N_3787,N_2687);
xnor U6224 (N_6224,N_3296,N_2596);
nor U6225 (N_6225,N_2940,N_4839);
nand U6226 (N_6226,N_3071,N_2584);
xnor U6227 (N_6227,N_3473,N_3925);
nand U6228 (N_6228,N_4841,N_2766);
or U6229 (N_6229,N_3721,N_3378);
xnor U6230 (N_6230,N_4477,N_2658);
nor U6231 (N_6231,N_3035,N_4078);
nand U6232 (N_6232,N_2853,N_3565);
nor U6233 (N_6233,N_3002,N_4051);
xnor U6234 (N_6234,N_3498,N_4617);
nand U6235 (N_6235,N_4801,N_3933);
and U6236 (N_6236,N_2785,N_4475);
xnor U6237 (N_6237,N_3600,N_3408);
nor U6238 (N_6238,N_4872,N_4349);
or U6239 (N_6239,N_4959,N_3325);
nand U6240 (N_6240,N_2802,N_2730);
nor U6241 (N_6241,N_4136,N_3791);
or U6242 (N_6242,N_4323,N_3735);
nand U6243 (N_6243,N_4516,N_2623);
and U6244 (N_6244,N_4539,N_3235);
and U6245 (N_6245,N_4450,N_3367);
nor U6246 (N_6246,N_3251,N_2968);
and U6247 (N_6247,N_3687,N_4926);
and U6248 (N_6248,N_4848,N_3856);
xnor U6249 (N_6249,N_3577,N_4082);
nand U6250 (N_6250,N_4099,N_2884);
xnor U6251 (N_6251,N_4641,N_3322);
nand U6252 (N_6252,N_4598,N_4725);
and U6253 (N_6253,N_4155,N_4823);
and U6254 (N_6254,N_4533,N_3397);
or U6255 (N_6255,N_2502,N_2992);
or U6256 (N_6256,N_2513,N_2996);
and U6257 (N_6257,N_4187,N_2813);
or U6258 (N_6258,N_3376,N_3748);
and U6259 (N_6259,N_3174,N_4376);
nand U6260 (N_6260,N_3725,N_3830);
nor U6261 (N_6261,N_4034,N_3913);
or U6262 (N_6262,N_3433,N_4135);
and U6263 (N_6263,N_3004,N_2802);
nand U6264 (N_6264,N_3649,N_4027);
and U6265 (N_6265,N_2669,N_4414);
or U6266 (N_6266,N_3655,N_2876);
xor U6267 (N_6267,N_3116,N_3582);
nand U6268 (N_6268,N_2622,N_4999);
xor U6269 (N_6269,N_4530,N_3183);
xor U6270 (N_6270,N_3618,N_3264);
nor U6271 (N_6271,N_3061,N_3979);
nor U6272 (N_6272,N_3891,N_3131);
and U6273 (N_6273,N_4456,N_2639);
nand U6274 (N_6274,N_3655,N_2962);
and U6275 (N_6275,N_2705,N_3155);
xnor U6276 (N_6276,N_4366,N_3537);
nand U6277 (N_6277,N_2683,N_4564);
and U6278 (N_6278,N_3043,N_3544);
nor U6279 (N_6279,N_3084,N_4955);
xor U6280 (N_6280,N_3452,N_4099);
nor U6281 (N_6281,N_4383,N_4775);
nor U6282 (N_6282,N_2949,N_4217);
nor U6283 (N_6283,N_4084,N_4792);
nor U6284 (N_6284,N_3594,N_3858);
or U6285 (N_6285,N_3245,N_3547);
nand U6286 (N_6286,N_2710,N_3410);
xor U6287 (N_6287,N_2881,N_2756);
and U6288 (N_6288,N_3365,N_2781);
and U6289 (N_6289,N_4338,N_4987);
xnor U6290 (N_6290,N_4919,N_4840);
xnor U6291 (N_6291,N_4453,N_4072);
nor U6292 (N_6292,N_3118,N_4875);
nor U6293 (N_6293,N_4116,N_3617);
nand U6294 (N_6294,N_4830,N_4217);
and U6295 (N_6295,N_2857,N_3232);
or U6296 (N_6296,N_4732,N_4879);
and U6297 (N_6297,N_4654,N_3908);
nor U6298 (N_6298,N_3391,N_2707);
nand U6299 (N_6299,N_3362,N_4041);
or U6300 (N_6300,N_4834,N_4073);
and U6301 (N_6301,N_4363,N_4214);
and U6302 (N_6302,N_4195,N_3184);
nor U6303 (N_6303,N_4480,N_4684);
and U6304 (N_6304,N_3084,N_3812);
nor U6305 (N_6305,N_4714,N_3856);
or U6306 (N_6306,N_3518,N_3397);
or U6307 (N_6307,N_3303,N_3498);
nor U6308 (N_6308,N_3077,N_3337);
xnor U6309 (N_6309,N_4596,N_2538);
and U6310 (N_6310,N_4453,N_3036);
nand U6311 (N_6311,N_3390,N_4806);
xor U6312 (N_6312,N_2792,N_2832);
nor U6313 (N_6313,N_3476,N_4683);
or U6314 (N_6314,N_2565,N_4919);
or U6315 (N_6315,N_3662,N_4344);
nor U6316 (N_6316,N_2630,N_2750);
and U6317 (N_6317,N_4334,N_3566);
nor U6318 (N_6318,N_2545,N_2749);
nor U6319 (N_6319,N_4620,N_4923);
nand U6320 (N_6320,N_3786,N_3858);
and U6321 (N_6321,N_4680,N_3950);
nor U6322 (N_6322,N_4722,N_4053);
xor U6323 (N_6323,N_4098,N_3231);
nand U6324 (N_6324,N_3360,N_2684);
xor U6325 (N_6325,N_3438,N_3890);
nor U6326 (N_6326,N_4021,N_3002);
nor U6327 (N_6327,N_3548,N_3522);
xor U6328 (N_6328,N_4272,N_3210);
and U6329 (N_6329,N_4343,N_3501);
or U6330 (N_6330,N_3736,N_3105);
xor U6331 (N_6331,N_3706,N_3630);
or U6332 (N_6332,N_3638,N_3980);
nor U6333 (N_6333,N_2837,N_2676);
or U6334 (N_6334,N_3550,N_3981);
nor U6335 (N_6335,N_2845,N_4508);
nand U6336 (N_6336,N_3357,N_4008);
nor U6337 (N_6337,N_3648,N_4616);
and U6338 (N_6338,N_4896,N_4581);
or U6339 (N_6339,N_4865,N_3010);
nand U6340 (N_6340,N_4274,N_2619);
nand U6341 (N_6341,N_4091,N_2545);
or U6342 (N_6342,N_3776,N_3651);
and U6343 (N_6343,N_4632,N_4117);
or U6344 (N_6344,N_2881,N_3940);
and U6345 (N_6345,N_4446,N_4787);
or U6346 (N_6346,N_2586,N_2794);
or U6347 (N_6347,N_3943,N_3212);
nor U6348 (N_6348,N_4715,N_3457);
and U6349 (N_6349,N_3793,N_3691);
or U6350 (N_6350,N_3537,N_2891);
nand U6351 (N_6351,N_2571,N_4230);
xor U6352 (N_6352,N_4195,N_4833);
nor U6353 (N_6353,N_2971,N_2533);
nor U6354 (N_6354,N_2666,N_4441);
nor U6355 (N_6355,N_2525,N_4712);
xnor U6356 (N_6356,N_3452,N_2836);
nand U6357 (N_6357,N_4069,N_3023);
or U6358 (N_6358,N_3966,N_2538);
nor U6359 (N_6359,N_3794,N_3230);
nor U6360 (N_6360,N_4019,N_4620);
nor U6361 (N_6361,N_4431,N_2691);
nor U6362 (N_6362,N_4558,N_3409);
xnor U6363 (N_6363,N_4373,N_4407);
xor U6364 (N_6364,N_2939,N_3724);
nor U6365 (N_6365,N_4691,N_4314);
or U6366 (N_6366,N_3033,N_2519);
or U6367 (N_6367,N_2790,N_4664);
or U6368 (N_6368,N_3528,N_4323);
nand U6369 (N_6369,N_3820,N_3145);
xnor U6370 (N_6370,N_3281,N_4018);
xnor U6371 (N_6371,N_4541,N_2545);
nor U6372 (N_6372,N_2737,N_2887);
or U6373 (N_6373,N_4924,N_3524);
nand U6374 (N_6374,N_4557,N_4660);
nand U6375 (N_6375,N_3334,N_4853);
or U6376 (N_6376,N_3427,N_4782);
nor U6377 (N_6377,N_4009,N_4084);
or U6378 (N_6378,N_4787,N_3292);
nor U6379 (N_6379,N_2596,N_3239);
and U6380 (N_6380,N_4016,N_2755);
nor U6381 (N_6381,N_3881,N_2600);
and U6382 (N_6382,N_4021,N_3375);
and U6383 (N_6383,N_4432,N_3961);
nand U6384 (N_6384,N_3390,N_2984);
xor U6385 (N_6385,N_4870,N_4216);
nor U6386 (N_6386,N_4854,N_4608);
xnor U6387 (N_6387,N_3864,N_2811);
xor U6388 (N_6388,N_4615,N_3315);
xor U6389 (N_6389,N_2624,N_3975);
nor U6390 (N_6390,N_4087,N_3963);
or U6391 (N_6391,N_4326,N_3691);
nor U6392 (N_6392,N_4705,N_4915);
xor U6393 (N_6393,N_3093,N_2615);
xnor U6394 (N_6394,N_4876,N_4485);
or U6395 (N_6395,N_2601,N_3266);
nor U6396 (N_6396,N_4616,N_2711);
xor U6397 (N_6397,N_3705,N_2935);
and U6398 (N_6398,N_3544,N_3000);
or U6399 (N_6399,N_2705,N_3214);
nor U6400 (N_6400,N_4483,N_4830);
or U6401 (N_6401,N_4382,N_3808);
nand U6402 (N_6402,N_2974,N_3982);
nand U6403 (N_6403,N_2729,N_4002);
or U6404 (N_6404,N_3265,N_4789);
xor U6405 (N_6405,N_3273,N_3935);
and U6406 (N_6406,N_4784,N_4415);
xnor U6407 (N_6407,N_4751,N_4288);
or U6408 (N_6408,N_3494,N_4308);
and U6409 (N_6409,N_2725,N_4204);
or U6410 (N_6410,N_3706,N_4084);
and U6411 (N_6411,N_2518,N_4266);
nand U6412 (N_6412,N_4956,N_4376);
and U6413 (N_6413,N_4294,N_3384);
xnor U6414 (N_6414,N_2935,N_3678);
nand U6415 (N_6415,N_3012,N_4228);
nand U6416 (N_6416,N_3925,N_3892);
and U6417 (N_6417,N_4509,N_2613);
nor U6418 (N_6418,N_3760,N_2838);
xnor U6419 (N_6419,N_2962,N_3229);
xnor U6420 (N_6420,N_4194,N_3328);
and U6421 (N_6421,N_3664,N_4651);
nand U6422 (N_6422,N_4640,N_2508);
and U6423 (N_6423,N_3977,N_2839);
and U6424 (N_6424,N_4291,N_3867);
nand U6425 (N_6425,N_2734,N_3965);
or U6426 (N_6426,N_4760,N_3740);
nand U6427 (N_6427,N_4081,N_2508);
or U6428 (N_6428,N_3633,N_4806);
nand U6429 (N_6429,N_3079,N_4205);
or U6430 (N_6430,N_3418,N_4854);
nand U6431 (N_6431,N_3268,N_4841);
nor U6432 (N_6432,N_3151,N_4371);
or U6433 (N_6433,N_4805,N_4904);
or U6434 (N_6434,N_4890,N_3959);
xor U6435 (N_6435,N_2993,N_2637);
xor U6436 (N_6436,N_4414,N_3993);
xnor U6437 (N_6437,N_2933,N_3197);
nand U6438 (N_6438,N_4771,N_2844);
nor U6439 (N_6439,N_3684,N_3752);
nand U6440 (N_6440,N_3994,N_4405);
xor U6441 (N_6441,N_4266,N_3607);
nand U6442 (N_6442,N_4972,N_3714);
or U6443 (N_6443,N_3682,N_3918);
nand U6444 (N_6444,N_3299,N_4121);
nor U6445 (N_6445,N_4472,N_3048);
nor U6446 (N_6446,N_3277,N_4048);
nor U6447 (N_6447,N_3486,N_3550);
or U6448 (N_6448,N_4508,N_4220);
or U6449 (N_6449,N_2801,N_4252);
or U6450 (N_6450,N_3410,N_4393);
nand U6451 (N_6451,N_4370,N_2989);
xor U6452 (N_6452,N_2906,N_3859);
nand U6453 (N_6453,N_4879,N_2955);
xor U6454 (N_6454,N_4312,N_2866);
xnor U6455 (N_6455,N_2674,N_2614);
nand U6456 (N_6456,N_3873,N_2798);
xnor U6457 (N_6457,N_3144,N_2800);
and U6458 (N_6458,N_4271,N_3182);
nand U6459 (N_6459,N_3802,N_4656);
and U6460 (N_6460,N_2732,N_4048);
and U6461 (N_6461,N_3296,N_4091);
or U6462 (N_6462,N_3500,N_4666);
or U6463 (N_6463,N_2574,N_4571);
nor U6464 (N_6464,N_2884,N_3522);
or U6465 (N_6465,N_4340,N_4868);
or U6466 (N_6466,N_3245,N_2876);
nor U6467 (N_6467,N_3909,N_4430);
or U6468 (N_6468,N_4982,N_4985);
nor U6469 (N_6469,N_3094,N_2503);
nor U6470 (N_6470,N_3381,N_2880);
nor U6471 (N_6471,N_2515,N_4482);
nand U6472 (N_6472,N_4753,N_3961);
nand U6473 (N_6473,N_4144,N_4793);
nand U6474 (N_6474,N_3836,N_3392);
or U6475 (N_6475,N_4537,N_2619);
nor U6476 (N_6476,N_3289,N_4027);
or U6477 (N_6477,N_3445,N_4809);
or U6478 (N_6478,N_3305,N_2847);
and U6479 (N_6479,N_3579,N_3950);
nor U6480 (N_6480,N_2831,N_3818);
or U6481 (N_6481,N_4234,N_3142);
nor U6482 (N_6482,N_3700,N_3797);
xor U6483 (N_6483,N_3861,N_3179);
nand U6484 (N_6484,N_4280,N_4858);
or U6485 (N_6485,N_4767,N_3661);
nand U6486 (N_6486,N_4275,N_3510);
and U6487 (N_6487,N_4190,N_3383);
xnor U6488 (N_6488,N_2973,N_3581);
and U6489 (N_6489,N_3716,N_3709);
nand U6490 (N_6490,N_2781,N_2993);
nand U6491 (N_6491,N_3504,N_2727);
nand U6492 (N_6492,N_4113,N_2513);
xor U6493 (N_6493,N_4040,N_3815);
and U6494 (N_6494,N_3913,N_3729);
or U6495 (N_6495,N_4886,N_2591);
or U6496 (N_6496,N_3979,N_2515);
xor U6497 (N_6497,N_3720,N_2751);
or U6498 (N_6498,N_2547,N_4097);
and U6499 (N_6499,N_2597,N_4633);
nor U6500 (N_6500,N_3505,N_3068);
and U6501 (N_6501,N_2536,N_4819);
and U6502 (N_6502,N_3562,N_4183);
and U6503 (N_6503,N_3895,N_4424);
or U6504 (N_6504,N_3080,N_3216);
and U6505 (N_6505,N_2791,N_4624);
xor U6506 (N_6506,N_3697,N_4575);
xor U6507 (N_6507,N_4572,N_3175);
nand U6508 (N_6508,N_4364,N_3963);
and U6509 (N_6509,N_3574,N_4138);
or U6510 (N_6510,N_4663,N_4700);
nor U6511 (N_6511,N_4977,N_2966);
xor U6512 (N_6512,N_4071,N_3350);
and U6513 (N_6513,N_3906,N_3891);
nand U6514 (N_6514,N_2611,N_4272);
and U6515 (N_6515,N_3818,N_2750);
nor U6516 (N_6516,N_3545,N_4636);
and U6517 (N_6517,N_2870,N_3794);
nor U6518 (N_6518,N_4384,N_3553);
nor U6519 (N_6519,N_3320,N_3372);
xor U6520 (N_6520,N_3774,N_4580);
and U6521 (N_6521,N_4552,N_3475);
and U6522 (N_6522,N_2895,N_3840);
or U6523 (N_6523,N_4432,N_3680);
and U6524 (N_6524,N_3986,N_4249);
xor U6525 (N_6525,N_3581,N_4129);
or U6526 (N_6526,N_4178,N_4624);
xor U6527 (N_6527,N_2875,N_4702);
and U6528 (N_6528,N_3306,N_2659);
nand U6529 (N_6529,N_3480,N_4905);
or U6530 (N_6530,N_3957,N_3638);
nand U6531 (N_6531,N_3000,N_2898);
nor U6532 (N_6532,N_3492,N_3682);
nand U6533 (N_6533,N_3849,N_4749);
and U6534 (N_6534,N_3925,N_3751);
xor U6535 (N_6535,N_2763,N_4708);
nand U6536 (N_6536,N_2737,N_4840);
nor U6537 (N_6537,N_4595,N_3605);
and U6538 (N_6538,N_4848,N_2904);
nand U6539 (N_6539,N_4364,N_3930);
or U6540 (N_6540,N_3299,N_3059);
nand U6541 (N_6541,N_2599,N_3324);
or U6542 (N_6542,N_3759,N_3383);
or U6543 (N_6543,N_3304,N_4998);
nor U6544 (N_6544,N_4402,N_3445);
and U6545 (N_6545,N_4874,N_4324);
nor U6546 (N_6546,N_3911,N_3620);
and U6547 (N_6547,N_4983,N_4395);
nand U6548 (N_6548,N_3838,N_4805);
or U6549 (N_6549,N_4051,N_3289);
and U6550 (N_6550,N_3591,N_2869);
or U6551 (N_6551,N_3541,N_3272);
nor U6552 (N_6552,N_4001,N_3309);
nand U6553 (N_6553,N_4273,N_3901);
nor U6554 (N_6554,N_2981,N_4223);
nor U6555 (N_6555,N_2601,N_3689);
nor U6556 (N_6556,N_4923,N_4485);
or U6557 (N_6557,N_4778,N_3506);
xor U6558 (N_6558,N_3634,N_3258);
xor U6559 (N_6559,N_2802,N_4733);
and U6560 (N_6560,N_4229,N_3763);
or U6561 (N_6561,N_3403,N_4752);
or U6562 (N_6562,N_4227,N_2637);
xor U6563 (N_6563,N_2743,N_4369);
nor U6564 (N_6564,N_3195,N_3209);
xor U6565 (N_6565,N_2643,N_4377);
nor U6566 (N_6566,N_4110,N_2544);
xnor U6567 (N_6567,N_4383,N_4536);
xor U6568 (N_6568,N_3733,N_3734);
and U6569 (N_6569,N_3991,N_4988);
nand U6570 (N_6570,N_3165,N_2885);
and U6571 (N_6571,N_3807,N_4254);
and U6572 (N_6572,N_4037,N_2701);
or U6573 (N_6573,N_4222,N_3950);
and U6574 (N_6574,N_3498,N_3295);
nand U6575 (N_6575,N_3827,N_3909);
xor U6576 (N_6576,N_3341,N_3454);
nor U6577 (N_6577,N_2806,N_3192);
or U6578 (N_6578,N_4487,N_4215);
xor U6579 (N_6579,N_3862,N_3608);
xor U6580 (N_6580,N_4263,N_4607);
xor U6581 (N_6581,N_2788,N_3769);
nor U6582 (N_6582,N_3837,N_4762);
and U6583 (N_6583,N_3343,N_2920);
and U6584 (N_6584,N_3232,N_3481);
or U6585 (N_6585,N_4595,N_2652);
nand U6586 (N_6586,N_3503,N_3554);
and U6587 (N_6587,N_3749,N_4948);
and U6588 (N_6588,N_3547,N_3170);
xnor U6589 (N_6589,N_2925,N_4863);
nor U6590 (N_6590,N_2542,N_3789);
or U6591 (N_6591,N_4948,N_4571);
and U6592 (N_6592,N_2733,N_2863);
or U6593 (N_6593,N_4729,N_4965);
nor U6594 (N_6594,N_4027,N_3242);
xnor U6595 (N_6595,N_4221,N_3034);
xor U6596 (N_6596,N_3542,N_3498);
nor U6597 (N_6597,N_3021,N_3003);
nand U6598 (N_6598,N_4341,N_4380);
xnor U6599 (N_6599,N_3112,N_2684);
nand U6600 (N_6600,N_4543,N_2734);
nand U6601 (N_6601,N_3409,N_2764);
nor U6602 (N_6602,N_2745,N_3685);
nor U6603 (N_6603,N_2693,N_2687);
nand U6604 (N_6604,N_4903,N_4148);
nand U6605 (N_6605,N_4778,N_4123);
nand U6606 (N_6606,N_4922,N_4431);
nor U6607 (N_6607,N_3525,N_2735);
and U6608 (N_6608,N_3658,N_4003);
and U6609 (N_6609,N_3411,N_3802);
nor U6610 (N_6610,N_4179,N_2875);
xnor U6611 (N_6611,N_3509,N_3227);
xor U6612 (N_6612,N_2643,N_3661);
or U6613 (N_6613,N_2709,N_3591);
xnor U6614 (N_6614,N_4078,N_3195);
nand U6615 (N_6615,N_3819,N_3683);
and U6616 (N_6616,N_3591,N_3799);
xnor U6617 (N_6617,N_3982,N_2887);
nand U6618 (N_6618,N_2914,N_2614);
and U6619 (N_6619,N_4741,N_3926);
or U6620 (N_6620,N_3652,N_4854);
nand U6621 (N_6621,N_3397,N_4263);
nor U6622 (N_6622,N_4872,N_4929);
nand U6623 (N_6623,N_4198,N_4451);
and U6624 (N_6624,N_3257,N_4268);
or U6625 (N_6625,N_2614,N_4541);
nor U6626 (N_6626,N_2614,N_3797);
nand U6627 (N_6627,N_4003,N_4130);
nand U6628 (N_6628,N_4364,N_2730);
and U6629 (N_6629,N_4426,N_4472);
nor U6630 (N_6630,N_2872,N_2574);
xor U6631 (N_6631,N_2500,N_4590);
and U6632 (N_6632,N_3189,N_3540);
nor U6633 (N_6633,N_4156,N_4280);
and U6634 (N_6634,N_3390,N_4512);
xnor U6635 (N_6635,N_3987,N_4962);
nor U6636 (N_6636,N_3646,N_4069);
or U6637 (N_6637,N_4419,N_3727);
or U6638 (N_6638,N_4363,N_2972);
and U6639 (N_6639,N_4347,N_4697);
nor U6640 (N_6640,N_4832,N_3093);
nand U6641 (N_6641,N_3807,N_4900);
xor U6642 (N_6642,N_4616,N_3917);
nand U6643 (N_6643,N_2802,N_3077);
and U6644 (N_6644,N_2563,N_4632);
and U6645 (N_6645,N_3089,N_4890);
nor U6646 (N_6646,N_4939,N_2983);
and U6647 (N_6647,N_2660,N_4469);
or U6648 (N_6648,N_4434,N_2573);
or U6649 (N_6649,N_3183,N_4789);
xor U6650 (N_6650,N_2599,N_2962);
xor U6651 (N_6651,N_4031,N_2800);
or U6652 (N_6652,N_3828,N_3023);
xnor U6653 (N_6653,N_3024,N_3279);
nor U6654 (N_6654,N_2904,N_2574);
xnor U6655 (N_6655,N_3083,N_4713);
and U6656 (N_6656,N_4284,N_2513);
and U6657 (N_6657,N_3187,N_2686);
and U6658 (N_6658,N_3596,N_2715);
nor U6659 (N_6659,N_4608,N_4571);
nand U6660 (N_6660,N_3090,N_4482);
or U6661 (N_6661,N_3356,N_3588);
nor U6662 (N_6662,N_4718,N_4070);
xor U6663 (N_6663,N_3874,N_4232);
nand U6664 (N_6664,N_3665,N_3386);
nand U6665 (N_6665,N_2797,N_2803);
xor U6666 (N_6666,N_3368,N_3208);
nand U6667 (N_6667,N_2612,N_3328);
nand U6668 (N_6668,N_3317,N_4207);
xor U6669 (N_6669,N_3480,N_3147);
and U6670 (N_6670,N_3973,N_2883);
or U6671 (N_6671,N_2917,N_3830);
and U6672 (N_6672,N_2995,N_3588);
nor U6673 (N_6673,N_3053,N_3710);
xor U6674 (N_6674,N_2973,N_3131);
and U6675 (N_6675,N_2970,N_4031);
nand U6676 (N_6676,N_3874,N_4526);
and U6677 (N_6677,N_3622,N_3707);
or U6678 (N_6678,N_3411,N_4196);
nor U6679 (N_6679,N_2953,N_4305);
nor U6680 (N_6680,N_4029,N_3554);
or U6681 (N_6681,N_3713,N_3146);
and U6682 (N_6682,N_4995,N_3642);
or U6683 (N_6683,N_2775,N_2638);
or U6684 (N_6684,N_3054,N_4914);
nand U6685 (N_6685,N_3489,N_3439);
or U6686 (N_6686,N_3808,N_3839);
xor U6687 (N_6687,N_2946,N_3711);
and U6688 (N_6688,N_2828,N_4447);
nand U6689 (N_6689,N_2787,N_2582);
or U6690 (N_6690,N_4440,N_3422);
nor U6691 (N_6691,N_3991,N_4147);
or U6692 (N_6692,N_2892,N_4805);
or U6693 (N_6693,N_4722,N_4898);
and U6694 (N_6694,N_4703,N_3341);
or U6695 (N_6695,N_4510,N_3346);
and U6696 (N_6696,N_2574,N_3566);
nor U6697 (N_6697,N_2992,N_4486);
nor U6698 (N_6698,N_3712,N_4796);
or U6699 (N_6699,N_4849,N_3513);
or U6700 (N_6700,N_3666,N_3425);
or U6701 (N_6701,N_4191,N_2796);
nor U6702 (N_6702,N_3188,N_3205);
xnor U6703 (N_6703,N_3084,N_4024);
nor U6704 (N_6704,N_2603,N_2976);
nand U6705 (N_6705,N_4372,N_2572);
xnor U6706 (N_6706,N_3484,N_2842);
or U6707 (N_6707,N_3810,N_2996);
and U6708 (N_6708,N_4896,N_4528);
nor U6709 (N_6709,N_4513,N_4903);
nand U6710 (N_6710,N_2827,N_4212);
nor U6711 (N_6711,N_4302,N_3845);
nor U6712 (N_6712,N_2543,N_3377);
or U6713 (N_6713,N_2649,N_4390);
or U6714 (N_6714,N_4943,N_3450);
and U6715 (N_6715,N_3614,N_4514);
and U6716 (N_6716,N_2762,N_2694);
nand U6717 (N_6717,N_4580,N_2661);
nand U6718 (N_6718,N_3648,N_3621);
or U6719 (N_6719,N_4134,N_3977);
xor U6720 (N_6720,N_2994,N_3004);
nand U6721 (N_6721,N_3128,N_2790);
and U6722 (N_6722,N_4217,N_4799);
xor U6723 (N_6723,N_3448,N_3429);
and U6724 (N_6724,N_3294,N_4083);
nand U6725 (N_6725,N_4447,N_2769);
nand U6726 (N_6726,N_4638,N_3064);
or U6727 (N_6727,N_3920,N_4684);
and U6728 (N_6728,N_2661,N_3477);
or U6729 (N_6729,N_3270,N_2503);
xor U6730 (N_6730,N_4541,N_2575);
nand U6731 (N_6731,N_4244,N_4085);
xnor U6732 (N_6732,N_3023,N_4796);
nand U6733 (N_6733,N_4650,N_2604);
xnor U6734 (N_6734,N_4272,N_3137);
nand U6735 (N_6735,N_2568,N_4973);
and U6736 (N_6736,N_4569,N_3298);
and U6737 (N_6737,N_4392,N_4448);
nand U6738 (N_6738,N_3401,N_2606);
or U6739 (N_6739,N_3526,N_4945);
or U6740 (N_6740,N_4944,N_2702);
xor U6741 (N_6741,N_4017,N_3685);
or U6742 (N_6742,N_3622,N_2964);
and U6743 (N_6743,N_2940,N_3354);
and U6744 (N_6744,N_4025,N_2799);
nor U6745 (N_6745,N_4203,N_4709);
and U6746 (N_6746,N_2663,N_2869);
nand U6747 (N_6747,N_3278,N_3092);
and U6748 (N_6748,N_4368,N_2706);
nor U6749 (N_6749,N_3844,N_3814);
nor U6750 (N_6750,N_2999,N_2566);
and U6751 (N_6751,N_4499,N_4228);
nand U6752 (N_6752,N_3494,N_2589);
xor U6753 (N_6753,N_4139,N_4342);
nand U6754 (N_6754,N_4552,N_2861);
xnor U6755 (N_6755,N_4409,N_3023);
nor U6756 (N_6756,N_3276,N_3144);
and U6757 (N_6757,N_2940,N_4983);
or U6758 (N_6758,N_3341,N_4491);
nand U6759 (N_6759,N_3930,N_3681);
nor U6760 (N_6760,N_4412,N_4555);
xnor U6761 (N_6761,N_3825,N_4097);
nor U6762 (N_6762,N_2924,N_4010);
nand U6763 (N_6763,N_4466,N_3094);
or U6764 (N_6764,N_2628,N_3431);
xor U6765 (N_6765,N_4994,N_3436);
nor U6766 (N_6766,N_3717,N_4739);
nand U6767 (N_6767,N_4907,N_3097);
or U6768 (N_6768,N_4913,N_4889);
xor U6769 (N_6769,N_4028,N_4910);
nand U6770 (N_6770,N_4079,N_4581);
nor U6771 (N_6771,N_2506,N_3329);
or U6772 (N_6772,N_4935,N_4311);
and U6773 (N_6773,N_4226,N_3573);
or U6774 (N_6774,N_3446,N_3050);
nor U6775 (N_6775,N_2694,N_2606);
and U6776 (N_6776,N_3840,N_3918);
xnor U6777 (N_6777,N_2856,N_3010);
nor U6778 (N_6778,N_2934,N_3526);
or U6779 (N_6779,N_3760,N_3700);
nor U6780 (N_6780,N_3046,N_4904);
nor U6781 (N_6781,N_3530,N_3893);
nor U6782 (N_6782,N_4482,N_3520);
or U6783 (N_6783,N_4932,N_2965);
or U6784 (N_6784,N_2967,N_4218);
and U6785 (N_6785,N_4587,N_3339);
nand U6786 (N_6786,N_3902,N_4590);
or U6787 (N_6787,N_3690,N_4504);
xnor U6788 (N_6788,N_3560,N_4129);
nor U6789 (N_6789,N_2610,N_3028);
or U6790 (N_6790,N_2947,N_2794);
or U6791 (N_6791,N_2536,N_3969);
xor U6792 (N_6792,N_4393,N_3700);
xnor U6793 (N_6793,N_3791,N_2765);
and U6794 (N_6794,N_3153,N_2760);
or U6795 (N_6795,N_2526,N_3168);
nand U6796 (N_6796,N_3598,N_2671);
and U6797 (N_6797,N_4762,N_4650);
nor U6798 (N_6798,N_4516,N_3536);
nand U6799 (N_6799,N_2947,N_3214);
and U6800 (N_6800,N_2572,N_4316);
or U6801 (N_6801,N_3463,N_4756);
or U6802 (N_6802,N_4015,N_4398);
and U6803 (N_6803,N_4130,N_2959);
and U6804 (N_6804,N_3992,N_4593);
xor U6805 (N_6805,N_3453,N_4619);
nand U6806 (N_6806,N_3187,N_3485);
xor U6807 (N_6807,N_4751,N_4863);
nor U6808 (N_6808,N_3202,N_4676);
and U6809 (N_6809,N_2637,N_4700);
and U6810 (N_6810,N_3109,N_2502);
and U6811 (N_6811,N_4479,N_3770);
nand U6812 (N_6812,N_4956,N_4611);
and U6813 (N_6813,N_2960,N_4698);
xnor U6814 (N_6814,N_4395,N_3432);
nor U6815 (N_6815,N_2543,N_4689);
xnor U6816 (N_6816,N_3845,N_2682);
and U6817 (N_6817,N_3062,N_3631);
nor U6818 (N_6818,N_4311,N_3739);
or U6819 (N_6819,N_3500,N_3531);
xor U6820 (N_6820,N_3295,N_3702);
nor U6821 (N_6821,N_4277,N_4617);
or U6822 (N_6822,N_3045,N_3709);
nor U6823 (N_6823,N_2954,N_3702);
nor U6824 (N_6824,N_4641,N_3930);
nand U6825 (N_6825,N_4847,N_4415);
xnor U6826 (N_6826,N_4926,N_4073);
nor U6827 (N_6827,N_3958,N_3408);
nand U6828 (N_6828,N_2858,N_3973);
or U6829 (N_6829,N_4004,N_4476);
nor U6830 (N_6830,N_3645,N_3582);
nor U6831 (N_6831,N_3364,N_4113);
nor U6832 (N_6832,N_3894,N_4281);
and U6833 (N_6833,N_4525,N_3075);
nand U6834 (N_6834,N_4216,N_4332);
nor U6835 (N_6835,N_2615,N_2952);
nor U6836 (N_6836,N_4382,N_3444);
and U6837 (N_6837,N_4755,N_4314);
or U6838 (N_6838,N_3894,N_4331);
nor U6839 (N_6839,N_3916,N_3413);
or U6840 (N_6840,N_4735,N_3613);
nand U6841 (N_6841,N_4904,N_4695);
and U6842 (N_6842,N_3262,N_4407);
or U6843 (N_6843,N_3220,N_3316);
nand U6844 (N_6844,N_3015,N_4602);
or U6845 (N_6845,N_3084,N_4460);
or U6846 (N_6846,N_2957,N_4762);
or U6847 (N_6847,N_4390,N_4148);
and U6848 (N_6848,N_3388,N_4061);
nand U6849 (N_6849,N_4322,N_2683);
nand U6850 (N_6850,N_4749,N_3858);
nor U6851 (N_6851,N_4252,N_2987);
nor U6852 (N_6852,N_4195,N_4603);
and U6853 (N_6853,N_4987,N_4774);
nand U6854 (N_6854,N_4115,N_4625);
and U6855 (N_6855,N_4428,N_3106);
xor U6856 (N_6856,N_3307,N_2584);
xnor U6857 (N_6857,N_3609,N_3303);
nor U6858 (N_6858,N_4562,N_3426);
and U6859 (N_6859,N_3643,N_3785);
nand U6860 (N_6860,N_4594,N_3371);
and U6861 (N_6861,N_4492,N_3364);
nand U6862 (N_6862,N_4438,N_4803);
or U6863 (N_6863,N_4011,N_2656);
or U6864 (N_6864,N_4236,N_3077);
and U6865 (N_6865,N_4008,N_2746);
nand U6866 (N_6866,N_3116,N_2840);
and U6867 (N_6867,N_3657,N_4144);
and U6868 (N_6868,N_4459,N_3549);
and U6869 (N_6869,N_3209,N_3529);
nand U6870 (N_6870,N_2628,N_3491);
xor U6871 (N_6871,N_2993,N_3189);
and U6872 (N_6872,N_3800,N_3227);
xnor U6873 (N_6873,N_3576,N_4230);
and U6874 (N_6874,N_3199,N_4367);
or U6875 (N_6875,N_2684,N_2963);
and U6876 (N_6876,N_2659,N_2781);
or U6877 (N_6877,N_4101,N_2870);
nor U6878 (N_6878,N_3683,N_2556);
nor U6879 (N_6879,N_4788,N_3624);
and U6880 (N_6880,N_4201,N_3976);
and U6881 (N_6881,N_4444,N_3650);
nor U6882 (N_6882,N_2826,N_4257);
nor U6883 (N_6883,N_3982,N_3364);
or U6884 (N_6884,N_2985,N_4676);
or U6885 (N_6885,N_4861,N_4256);
nor U6886 (N_6886,N_4408,N_3346);
xor U6887 (N_6887,N_2825,N_2645);
nand U6888 (N_6888,N_2642,N_3601);
or U6889 (N_6889,N_4497,N_4992);
nand U6890 (N_6890,N_4614,N_4635);
nor U6891 (N_6891,N_4385,N_4833);
xor U6892 (N_6892,N_3703,N_3794);
xor U6893 (N_6893,N_4486,N_3758);
or U6894 (N_6894,N_3409,N_2843);
or U6895 (N_6895,N_4194,N_2605);
and U6896 (N_6896,N_4924,N_4899);
nand U6897 (N_6897,N_4495,N_3902);
and U6898 (N_6898,N_4133,N_4817);
or U6899 (N_6899,N_4566,N_4637);
xor U6900 (N_6900,N_4044,N_2863);
or U6901 (N_6901,N_3244,N_3319);
xnor U6902 (N_6902,N_3387,N_2974);
nor U6903 (N_6903,N_2533,N_2727);
and U6904 (N_6904,N_4477,N_2634);
or U6905 (N_6905,N_2918,N_4439);
xnor U6906 (N_6906,N_3771,N_3440);
and U6907 (N_6907,N_2538,N_4386);
nand U6908 (N_6908,N_2772,N_4977);
xor U6909 (N_6909,N_4669,N_2527);
or U6910 (N_6910,N_2638,N_3880);
xnor U6911 (N_6911,N_2867,N_4885);
and U6912 (N_6912,N_3488,N_2840);
nand U6913 (N_6913,N_3501,N_3869);
and U6914 (N_6914,N_3160,N_3155);
or U6915 (N_6915,N_2859,N_4735);
and U6916 (N_6916,N_4698,N_3009);
nand U6917 (N_6917,N_4460,N_3876);
or U6918 (N_6918,N_4167,N_2716);
nor U6919 (N_6919,N_2868,N_4551);
xnor U6920 (N_6920,N_4478,N_4245);
nor U6921 (N_6921,N_3345,N_3017);
and U6922 (N_6922,N_4553,N_2521);
nor U6923 (N_6923,N_3720,N_3844);
xnor U6924 (N_6924,N_2573,N_2920);
and U6925 (N_6925,N_4136,N_3462);
and U6926 (N_6926,N_4857,N_4243);
nand U6927 (N_6927,N_4073,N_3052);
xor U6928 (N_6928,N_3318,N_3919);
and U6929 (N_6929,N_2588,N_4055);
or U6930 (N_6930,N_3482,N_4251);
nand U6931 (N_6931,N_4851,N_3706);
nor U6932 (N_6932,N_3563,N_2942);
or U6933 (N_6933,N_2730,N_3836);
xnor U6934 (N_6934,N_4042,N_4553);
nor U6935 (N_6935,N_4980,N_3571);
nor U6936 (N_6936,N_4120,N_4371);
and U6937 (N_6937,N_3951,N_4838);
or U6938 (N_6938,N_3622,N_4676);
or U6939 (N_6939,N_3965,N_3919);
xor U6940 (N_6940,N_3523,N_4855);
nand U6941 (N_6941,N_4395,N_3652);
and U6942 (N_6942,N_3049,N_4219);
nand U6943 (N_6943,N_4678,N_3008);
xnor U6944 (N_6944,N_4448,N_3068);
xnor U6945 (N_6945,N_4678,N_2949);
nor U6946 (N_6946,N_2733,N_4354);
or U6947 (N_6947,N_3406,N_3089);
nand U6948 (N_6948,N_3857,N_4652);
nor U6949 (N_6949,N_4299,N_4736);
xnor U6950 (N_6950,N_3472,N_3905);
nor U6951 (N_6951,N_2536,N_2925);
xor U6952 (N_6952,N_4929,N_2872);
and U6953 (N_6953,N_4630,N_3536);
or U6954 (N_6954,N_4836,N_4416);
xnor U6955 (N_6955,N_3933,N_3453);
xor U6956 (N_6956,N_3648,N_3585);
and U6957 (N_6957,N_3261,N_3660);
nand U6958 (N_6958,N_3831,N_2668);
nand U6959 (N_6959,N_4042,N_4283);
and U6960 (N_6960,N_3035,N_4372);
and U6961 (N_6961,N_3276,N_2907);
and U6962 (N_6962,N_4247,N_4743);
nand U6963 (N_6963,N_4330,N_2766);
nor U6964 (N_6964,N_4050,N_2641);
and U6965 (N_6965,N_4186,N_4338);
xnor U6966 (N_6966,N_2886,N_2747);
and U6967 (N_6967,N_4203,N_4651);
nand U6968 (N_6968,N_2732,N_3226);
nor U6969 (N_6969,N_4734,N_3929);
xor U6970 (N_6970,N_4083,N_4285);
or U6971 (N_6971,N_3013,N_4715);
nor U6972 (N_6972,N_4706,N_3093);
and U6973 (N_6973,N_3630,N_3820);
nor U6974 (N_6974,N_4402,N_4599);
xor U6975 (N_6975,N_3221,N_2989);
nor U6976 (N_6976,N_3512,N_4037);
and U6977 (N_6977,N_3513,N_3378);
nand U6978 (N_6978,N_4120,N_4775);
nand U6979 (N_6979,N_2584,N_2667);
xnor U6980 (N_6980,N_4308,N_3484);
or U6981 (N_6981,N_4971,N_4726);
xnor U6982 (N_6982,N_4960,N_3234);
xnor U6983 (N_6983,N_3757,N_3506);
nand U6984 (N_6984,N_4795,N_4391);
and U6985 (N_6985,N_4238,N_3857);
nor U6986 (N_6986,N_3020,N_3812);
xnor U6987 (N_6987,N_2615,N_4354);
nand U6988 (N_6988,N_2509,N_4874);
nand U6989 (N_6989,N_3163,N_4814);
or U6990 (N_6990,N_4662,N_4804);
nand U6991 (N_6991,N_2774,N_2632);
or U6992 (N_6992,N_2523,N_2913);
or U6993 (N_6993,N_4984,N_3459);
xnor U6994 (N_6994,N_3627,N_4626);
xnor U6995 (N_6995,N_3236,N_4122);
xor U6996 (N_6996,N_3456,N_4018);
or U6997 (N_6997,N_4357,N_4602);
and U6998 (N_6998,N_4660,N_3090);
nor U6999 (N_6999,N_3929,N_4619);
and U7000 (N_7000,N_2918,N_4846);
nor U7001 (N_7001,N_2958,N_4082);
xnor U7002 (N_7002,N_3998,N_4380);
xnor U7003 (N_7003,N_3210,N_3551);
xor U7004 (N_7004,N_4530,N_2708);
and U7005 (N_7005,N_4742,N_4400);
nand U7006 (N_7006,N_3908,N_2928);
nand U7007 (N_7007,N_4686,N_2583);
or U7008 (N_7008,N_3009,N_4753);
and U7009 (N_7009,N_3574,N_3297);
nor U7010 (N_7010,N_2893,N_2703);
or U7011 (N_7011,N_3347,N_4854);
nor U7012 (N_7012,N_4537,N_2837);
nor U7013 (N_7013,N_2680,N_4516);
nor U7014 (N_7014,N_3918,N_3620);
or U7015 (N_7015,N_3915,N_4850);
or U7016 (N_7016,N_3321,N_4037);
and U7017 (N_7017,N_2828,N_2654);
xor U7018 (N_7018,N_3059,N_4126);
and U7019 (N_7019,N_4572,N_3644);
or U7020 (N_7020,N_3476,N_2993);
or U7021 (N_7021,N_3459,N_4993);
or U7022 (N_7022,N_4668,N_4642);
nor U7023 (N_7023,N_2852,N_2744);
nand U7024 (N_7024,N_4700,N_3004);
xnor U7025 (N_7025,N_3002,N_4200);
nor U7026 (N_7026,N_4475,N_3009);
or U7027 (N_7027,N_3995,N_3700);
and U7028 (N_7028,N_3512,N_3244);
xnor U7029 (N_7029,N_3015,N_4469);
nand U7030 (N_7030,N_4460,N_4505);
nor U7031 (N_7031,N_2839,N_2582);
nand U7032 (N_7032,N_4039,N_2797);
nor U7033 (N_7033,N_3956,N_3742);
nand U7034 (N_7034,N_3273,N_4053);
xnor U7035 (N_7035,N_3146,N_2674);
xor U7036 (N_7036,N_4641,N_4076);
and U7037 (N_7037,N_4402,N_4775);
or U7038 (N_7038,N_4490,N_2961);
nand U7039 (N_7039,N_4325,N_3915);
nor U7040 (N_7040,N_2729,N_3863);
and U7041 (N_7041,N_3907,N_3379);
nor U7042 (N_7042,N_3325,N_3995);
xor U7043 (N_7043,N_4834,N_4534);
nor U7044 (N_7044,N_4678,N_3704);
and U7045 (N_7045,N_4570,N_3194);
or U7046 (N_7046,N_4412,N_4561);
or U7047 (N_7047,N_2942,N_3862);
xor U7048 (N_7048,N_2704,N_4987);
and U7049 (N_7049,N_2753,N_4650);
or U7050 (N_7050,N_2648,N_4174);
nor U7051 (N_7051,N_3692,N_2917);
or U7052 (N_7052,N_3496,N_3208);
nand U7053 (N_7053,N_2704,N_2777);
nand U7054 (N_7054,N_4847,N_3627);
or U7055 (N_7055,N_4394,N_4538);
xnor U7056 (N_7056,N_4180,N_3417);
and U7057 (N_7057,N_3557,N_3606);
or U7058 (N_7058,N_4952,N_4671);
nand U7059 (N_7059,N_2592,N_2883);
xor U7060 (N_7060,N_4889,N_2697);
xor U7061 (N_7061,N_3392,N_2809);
and U7062 (N_7062,N_4139,N_3599);
xnor U7063 (N_7063,N_3474,N_3642);
nand U7064 (N_7064,N_3858,N_3807);
and U7065 (N_7065,N_2514,N_2770);
and U7066 (N_7066,N_3009,N_3344);
xnor U7067 (N_7067,N_2798,N_4190);
nand U7068 (N_7068,N_3211,N_4474);
nand U7069 (N_7069,N_4032,N_3936);
and U7070 (N_7070,N_3964,N_3473);
nor U7071 (N_7071,N_3125,N_2889);
nand U7072 (N_7072,N_4002,N_3860);
and U7073 (N_7073,N_4701,N_3532);
xnor U7074 (N_7074,N_3340,N_4840);
xnor U7075 (N_7075,N_3480,N_2722);
or U7076 (N_7076,N_3211,N_3212);
and U7077 (N_7077,N_3307,N_3278);
xor U7078 (N_7078,N_4049,N_4980);
xnor U7079 (N_7079,N_3026,N_4638);
xor U7080 (N_7080,N_2749,N_4638);
xor U7081 (N_7081,N_4691,N_4999);
or U7082 (N_7082,N_2756,N_4033);
or U7083 (N_7083,N_2544,N_2533);
nand U7084 (N_7084,N_3237,N_3305);
nor U7085 (N_7085,N_4191,N_4796);
and U7086 (N_7086,N_2636,N_2712);
nor U7087 (N_7087,N_3815,N_3656);
and U7088 (N_7088,N_4388,N_4851);
and U7089 (N_7089,N_3556,N_3798);
and U7090 (N_7090,N_4281,N_4990);
nor U7091 (N_7091,N_4005,N_3305);
and U7092 (N_7092,N_3435,N_3062);
and U7093 (N_7093,N_2529,N_4539);
and U7094 (N_7094,N_3842,N_3996);
nor U7095 (N_7095,N_3183,N_4717);
and U7096 (N_7096,N_3656,N_3576);
nor U7097 (N_7097,N_3209,N_4313);
xnor U7098 (N_7098,N_3803,N_4180);
xor U7099 (N_7099,N_3806,N_2718);
xor U7100 (N_7100,N_4614,N_4546);
xnor U7101 (N_7101,N_2984,N_4542);
or U7102 (N_7102,N_4525,N_2817);
nor U7103 (N_7103,N_4557,N_4585);
nor U7104 (N_7104,N_3965,N_2972);
or U7105 (N_7105,N_3556,N_2992);
and U7106 (N_7106,N_2510,N_4706);
and U7107 (N_7107,N_3645,N_3338);
nand U7108 (N_7108,N_4724,N_3444);
and U7109 (N_7109,N_3624,N_4318);
and U7110 (N_7110,N_4884,N_4946);
or U7111 (N_7111,N_3656,N_3548);
nor U7112 (N_7112,N_3038,N_3126);
nor U7113 (N_7113,N_4438,N_4329);
xnor U7114 (N_7114,N_4882,N_4692);
and U7115 (N_7115,N_3124,N_3756);
or U7116 (N_7116,N_3349,N_3191);
nand U7117 (N_7117,N_3694,N_4443);
or U7118 (N_7118,N_2943,N_3796);
or U7119 (N_7119,N_4487,N_4087);
nand U7120 (N_7120,N_3292,N_3488);
xnor U7121 (N_7121,N_3486,N_3423);
nand U7122 (N_7122,N_4535,N_4625);
xnor U7123 (N_7123,N_4773,N_4691);
or U7124 (N_7124,N_4223,N_4120);
nand U7125 (N_7125,N_4811,N_3434);
nand U7126 (N_7126,N_2755,N_4548);
or U7127 (N_7127,N_4332,N_3581);
and U7128 (N_7128,N_2595,N_4718);
nor U7129 (N_7129,N_4534,N_3468);
xnor U7130 (N_7130,N_3592,N_2564);
xnor U7131 (N_7131,N_3532,N_4733);
nor U7132 (N_7132,N_3628,N_3807);
nand U7133 (N_7133,N_3967,N_2531);
nand U7134 (N_7134,N_2536,N_4864);
nand U7135 (N_7135,N_4277,N_2970);
and U7136 (N_7136,N_4257,N_2987);
xor U7137 (N_7137,N_3062,N_2742);
and U7138 (N_7138,N_4542,N_3794);
or U7139 (N_7139,N_3846,N_4133);
xnor U7140 (N_7140,N_4501,N_4419);
nand U7141 (N_7141,N_2958,N_2565);
or U7142 (N_7142,N_3369,N_3057);
nand U7143 (N_7143,N_3396,N_4518);
nand U7144 (N_7144,N_4220,N_3772);
nand U7145 (N_7145,N_2917,N_3064);
xnor U7146 (N_7146,N_4083,N_3651);
xnor U7147 (N_7147,N_3614,N_4776);
xnor U7148 (N_7148,N_2723,N_4879);
nand U7149 (N_7149,N_4851,N_4784);
nand U7150 (N_7150,N_3291,N_2640);
nor U7151 (N_7151,N_4408,N_4696);
or U7152 (N_7152,N_2813,N_3735);
xnor U7153 (N_7153,N_4886,N_2754);
xor U7154 (N_7154,N_3296,N_3435);
nand U7155 (N_7155,N_3227,N_3215);
xor U7156 (N_7156,N_3614,N_4448);
nor U7157 (N_7157,N_3622,N_3017);
xor U7158 (N_7158,N_4724,N_3720);
nand U7159 (N_7159,N_3003,N_3121);
nand U7160 (N_7160,N_4790,N_4956);
or U7161 (N_7161,N_3999,N_4191);
xnor U7162 (N_7162,N_2980,N_4864);
nor U7163 (N_7163,N_3523,N_2765);
or U7164 (N_7164,N_3039,N_4082);
and U7165 (N_7165,N_3467,N_4914);
nor U7166 (N_7166,N_2777,N_3849);
nor U7167 (N_7167,N_4987,N_3395);
and U7168 (N_7168,N_3979,N_4916);
or U7169 (N_7169,N_3124,N_3551);
xor U7170 (N_7170,N_3954,N_4687);
xor U7171 (N_7171,N_3229,N_4085);
nor U7172 (N_7172,N_3443,N_2828);
xnor U7173 (N_7173,N_2963,N_4229);
nor U7174 (N_7174,N_2598,N_3802);
or U7175 (N_7175,N_2829,N_4236);
nand U7176 (N_7176,N_4381,N_2587);
nor U7177 (N_7177,N_3414,N_3948);
and U7178 (N_7178,N_3258,N_2587);
and U7179 (N_7179,N_3210,N_3683);
or U7180 (N_7180,N_4265,N_4198);
and U7181 (N_7181,N_2839,N_3175);
xor U7182 (N_7182,N_2774,N_3570);
nand U7183 (N_7183,N_4947,N_3804);
nand U7184 (N_7184,N_4770,N_2761);
nor U7185 (N_7185,N_4321,N_4009);
nand U7186 (N_7186,N_4419,N_2786);
and U7187 (N_7187,N_2575,N_2926);
xnor U7188 (N_7188,N_2781,N_4426);
xor U7189 (N_7189,N_2799,N_3387);
and U7190 (N_7190,N_4395,N_4711);
and U7191 (N_7191,N_3692,N_3751);
or U7192 (N_7192,N_4140,N_3168);
xor U7193 (N_7193,N_4494,N_4754);
xor U7194 (N_7194,N_3930,N_4070);
and U7195 (N_7195,N_3418,N_3613);
nand U7196 (N_7196,N_4934,N_4594);
and U7197 (N_7197,N_4125,N_2585);
nand U7198 (N_7198,N_2839,N_3359);
nor U7199 (N_7199,N_4479,N_2832);
and U7200 (N_7200,N_2981,N_3680);
nand U7201 (N_7201,N_3279,N_3984);
or U7202 (N_7202,N_3306,N_4745);
xnor U7203 (N_7203,N_2891,N_4408);
or U7204 (N_7204,N_2574,N_3815);
and U7205 (N_7205,N_3420,N_4148);
nor U7206 (N_7206,N_4571,N_4278);
nand U7207 (N_7207,N_4505,N_3459);
xnor U7208 (N_7208,N_4899,N_4654);
or U7209 (N_7209,N_2684,N_2568);
xor U7210 (N_7210,N_3276,N_3999);
nor U7211 (N_7211,N_4069,N_4438);
and U7212 (N_7212,N_2945,N_3466);
nor U7213 (N_7213,N_4462,N_3328);
xnor U7214 (N_7214,N_4271,N_3818);
nor U7215 (N_7215,N_4218,N_3198);
nor U7216 (N_7216,N_2559,N_2961);
xnor U7217 (N_7217,N_4668,N_3511);
or U7218 (N_7218,N_3352,N_4005);
nor U7219 (N_7219,N_4287,N_3904);
or U7220 (N_7220,N_4695,N_4275);
nand U7221 (N_7221,N_3651,N_4285);
xnor U7222 (N_7222,N_2772,N_4575);
xnor U7223 (N_7223,N_3879,N_3763);
nand U7224 (N_7224,N_3951,N_3647);
xnor U7225 (N_7225,N_4873,N_3867);
and U7226 (N_7226,N_4648,N_3150);
or U7227 (N_7227,N_4824,N_3472);
xnor U7228 (N_7228,N_3432,N_2965);
or U7229 (N_7229,N_3271,N_2918);
nand U7230 (N_7230,N_3645,N_3157);
xor U7231 (N_7231,N_3277,N_4866);
or U7232 (N_7232,N_3957,N_4713);
nand U7233 (N_7233,N_4521,N_4996);
xor U7234 (N_7234,N_3056,N_4743);
or U7235 (N_7235,N_3652,N_4713);
or U7236 (N_7236,N_4644,N_4194);
and U7237 (N_7237,N_4770,N_2954);
nor U7238 (N_7238,N_2630,N_2705);
or U7239 (N_7239,N_2529,N_3566);
nor U7240 (N_7240,N_2612,N_4332);
or U7241 (N_7241,N_4989,N_2631);
and U7242 (N_7242,N_4524,N_4027);
and U7243 (N_7243,N_2692,N_2571);
xnor U7244 (N_7244,N_4640,N_2897);
nor U7245 (N_7245,N_3399,N_4374);
or U7246 (N_7246,N_4685,N_4721);
or U7247 (N_7247,N_2866,N_2907);
or U7248 (N_7248,N_3792,N_4848);
or U7249 (N_7249,N_3632,N_3312);
nand U7250 (N_7250,N_2679,N_4085);
and U7251 (N_7251,N_2794,N_3143);
and U7252 (N_7252,N_4904,N_3504);
xnor U7253 (N_7253,N_4215,N_3878);
xor U7254 (N_7254,N_4803,N_4048);
and U7255 (N_7255,N_2555,N_4295);
xor U7256 (N_7256,N_2905,N_4097);
and U7257 (N_7257,N_4981,N_3084);
and U7258 (N_7258,N_3965,N_3910);
xor U7259 (N_7259,N_4349,N_3623);
nand U7260 (N_7260,N_3959,N_3851);
nand U7261 (N_7261,N_2859,N_3020);
nor U7262 (N_7262,N_4260,N_4992);
xor U7263 (N_7263,N_3515,N_3363);
and U7264 (N_7264,N_4424,N_3387);
or U7265 (N_7265,N_2985,N_3733);
nand U7266 (N_7266,N_2757,N_3858);
nor U7267 (N_7267,N_4891,N_4270);
or U7268 (N_7268,N_3570,N_3133);
nor U7269 (N_7269,N_2847,N_2955);
or U7270 (N_7270,N_2711,N_3892);
nor U7271 (N_7271,N_4986,N_3805);
xor U7272 (N_7272,N_3681,N_4483);
or U7273 (N_7273,N_4302,N_3035);
and U7274 (N_7274,N_3967,N_3554);
or U7275 (N_7275,N_4141,N_4559);
xnor U7276 (N_7276,N_3514,N_4736);
xor U7277 (N_7277,N_3399,N_3239);
or U7278 (N_7278,N_4016,N_3374);
and U7279 (N_7279,N_2566,N_3775);
and U7280 (N_7280,N_4990,N_2863);
xor U7281 (N_7281,N_4727,N_4896);
nor U7282 (N_7282,N_4707,N_3397);
or U7283 (N_7283,N_3096,N_3840);
xor U7284 (N_7284,N_3084,N_2705);
and U7285 (N_7285,N_4429,N_4669);
and U7286 (N_7286,N_2821,N_3318);
xnor U7287 (N_7287,N_4907,N_3172);
xnor U7288 (N_7288,N_2648,N_2727);
or U7289 (N_7289,N_2884,N_3150);
nor U7290 (N_7290,N_4986,N_2591);
and U7291 (N_7291,N_4760,N_3325);
nor U7292 (N_7292,N_4371,N_4438);
nand U7293 (N_7293,N_3861,N_4056);
nor U7294 (N_7294,N_2935,N_2655);
and U7295 (N_7295,N_2709,N_4666);
nand U7296 (N_7296,N_3552,N_4436);
nor U7297 (N_7297,N_4201,N_3459);
nor U7298 (N_7298,N_4579,N_4667);
nand U7299 (N_7299,N_3194,N_3191);
and U7300 (N_7300,N_2820,N_3373);
or U7301 (N_7301,N_4910,N_3891);
and U7302 (N_7302,N_3380,N_3385);
nand U7303 (N_7303,N_3546,N_4304);
nor U7304 (N_7304,N_4327,N_4917);
nor U7305 (N_7305,N_4290,N_3861);
or U7306 (N_7306,N_2603,N_3302);
and U7307 (N_7307,N_4014,N_2991);
nor U7308 (N_7308,N_3017,N_4584);
and U7309 (N_7309,N_2808,N_4396);
xnor U7310 (N_7310,N_4295,N_4238);
nor U7311 (N_7311,N_3016,N_4654);
nor U7312 (N_7312,N_4705,N_2639);
and U7313 (N_7313,N_3995,N_3238);
nand U7314 (N_7314,N_4444,N_2544);
xor U7315 (N_7315,N_3299,N_4851);
or U7316 (N_7316,N_3704,N_2643);
or U7317 (N_7317,N_4405,N_4600);
and U7318 (N_7318,N_3175,N_4432);
nand U7319 (N_7319,N_4239,N_4480);
and U7320 (N_7320,N_4024,N_2965);
xor U7321 (N_7321,N_3152,N_2874);
nand U7322 (N_7322,N_3820,N_4719);
xnor U7323 (N_7323,N_4846,N_4321);
nor U7324 (N_7324,N_3862,N_4369);
and U7325 (N_7325,N_2500,N_4404);
nor U7326 (N_7326,N_3204,N_3706);
xor U7327 (N_7327,N_2717,N_3538);
and U7328 (N_7328,N_2707,N_3177);
or U7329 (N_7329,N_3618,N_4883);
xnor U7330 (N_7330,N_4842,N_3091);
xor U7331 (N_7331,N_3165,N_3817);
xnor U7332 (N_7332,N_4691,N_2608);
nor U7333 (N_7333,N_3183,N_2954);
nor U7334 (N_7334,N_4678,N_4957);
nor U7335 (N_7335,N_3861,N_4431);
and U7336 (N_7336,N_3551,N_4578);
xor U7337 (N_7337,N_4932,N_3814);
xnor U7338 (N_7338,N_3835,N_4185);
and U7339 (N_7339,N_3564,N_2690);
and U7340 (N_7340,N_3795,N_4792);
or U7341 (N_7341,N_3103,N_3311);
nor U7342 (N_7342,N_4059,N_4404);
xor U7343 (N_7343,N_4264,N_3831);
xor U7344 (N_7344,N_3511,N_4008);
xor U7345 (N_7345,N_2941,N_2780);
or U7346 (N_7346,N_4175,N_3183);
xor U7347 (N_7347,N_4270,N_2862);
and U7348 (N_7348,N_4855,N_3454);
and U7349 (N_7349,N_4885,N_4496);
nand U7350 (N_7350,N_4941,N_4432);
nor U7351 (N_7351,N_3672,N_4895);
nand U7352 (N_7352,N_4832,N_4249);
or U7353 (N_7353,N_3679,N_2719);
nand U7354 (N_7354,N_3562,N_2937);
or U7355 (N_7355,N_3543,N_4938);
xor U7356 (N_7356,N_3686,N_2794);
nand U7357 (N_7357,N_4790,N_3015);
nor U7358 (N_7358,N_4030,N_2632);
nand U7359 (N_7359,N_2873,N_3129);
and U7360 (N_7360,N_4323,N_4812);
or U7361 (N_7361,N_3181,N_4338);
and U7362 (N_7362,N_3903,N_2543);
nand U7363 (N_7363,N_4831,N_4622);
and U7364 (N_7364,N_3296,N_2846);
and U7365 (N_7365,N_4690,N_3398);
nand U7366 (N_7366,N_4071,N_2890);
or U7367 (N_7367,N_3542,N_3893);
nand U7368 (N_7368,N_2736,N_2718);
nand U7369 (N_7369,N_4164,N_3040);
or U7370 (N_7370,N_3552,N_4100);
xnor U7371 (N_7371,N_3090,N_4014);
nor U7372 (N_7372,N_2904,N_4353);
or U7373 (N_7373,N_3265,N_4248);
nor U7374 (N_7374,N_4977,N_2508);
xor U7375 (N_7375,N_3291,N_4491);
or U7376 (N_7376,N_4056,N_4288);
nor U7377 (N_7377,N_3579,N_4550);
nor U7378 (N_7378,N_3314,N_3156);
nor U7379 (N_7379,N_3321,N_4335);
or U7380 (N_7380,N_3045,N_3407);
xor U7381 (N_7381,N_4438,N_3909);
and U7382 (N_7382,N_4247,N_3669);
and U7383 (N_7383,N_4999,N_3035);
or U7384 (N_7384,N_4158,N_3741);
nor U7385 (N_7385,N_2762,N_4415);
and U7386 (N_7386,N_2817,N_3537);
nor U7387 (N_7387,N_3005,N_4304);
and U7388 (N_7388,N_3139,N_4999);
nor U7389 (N_7389,N_3328,N_4017);
nor U7390 (N_7390,N_4346,N_3442);
or U7391 (N_7391,N_2714,N_2583);
and U7392 (N_7392,N_4488,N_3219);
nor U7393 (N_7393,N_2678,N_3874);
xnor U7394 (N_7394,N_4418,N_3896);
and U7395 (N_7395,N_3456,N_3952);
nand U7396 (N_7396,N_2864,N_4541);
or U7397 (N_7397,N_3112,N_3151);
nor U7398 (N_7398,N_4959,N_4903);
nor U7399 (N_7399,N_2636,N_2801);
or U7400 (N_7400,N_4874,N_2964);
nand U7401 (N_7401,N_3730,N_3492);
nor U7402 (N_7402,N_3973,N_3972);
nand U7403 (N_7403,N_4513,N_3601);
xor U7404 (N_7404,N_4191,N_4523);
and U7405 (N_7405,N_4453,N_4370);
and U7406 (N_7406,N_4312,N_4392);
xnor U7407 (N_7407,N_4429,N_3478);
nor U7408 (N_7408,N_4132,N_3399);
xnor U7409 (N_7409,N_2968,N_3335);
xor U7410 (N_7410,N_2617,N_4914);
nor U7411 (N_7411,N_2804,N_2560);
and U7412 (N_7412,N_4354,N_4286);
xor U7413 (N_7413,N_2851,N_3433);
xor U7414 (N_7414,N_3367,N_2638);
xor U7415 (N_7415,N_3104,N_3469);
and U7416 (N_7416,N_3044,N_4564);
and U7417 (N_7417,N_4048,N_3832);
xnor U7418 (N_7418,N_3712,N_4786);
nand U7419 (N_7419,N_3847,N_4241);
nand U7420 (N_7420,N_4048,N_3907);
and U7421 (N_7421,N_4207,N_4473);
nor U7422 (N_7422,N_3176,N_3359);
or U7423 (N_7423,N_3985,N_4892);
nand U7424 (N_7424,N_2740,N_3094);
nand U7425 (N_7425,N_2607,N_4073);
nand U7426 (N_7426,N_3665,N_2537);
nor U7427 (N_7427,N_4162,N_2759);
xor U7428 (N_7428,N_3445,N_4038);
nand U7429 (N_7429,N_4993,N_4438);
nand U7430 (N_7430,N_4204,N_3536);
nand U7431 (N_7431,N_2774,N_2824);
nor U7432 (N_7432,N_4950,N_3588);
nor U7433 (N_7433,N_4383,N_3755);
or U7434 (N_7434,N_3063,N_3306);
or U7435 (N_7435,N_4971,N_3087);
nor U7436 (N_7436,N_3375,N_3045);
nor U7437 (N_7437,N_3090,N_4909);
and U7438 (N_7438,N_3312,N_3259);
and U7439 (N_7439,N_3515,N_3512);
nand U7440 (N_7440,N_4415,N_4759);
or U7441 (N_7441,N_3012,N_2625);
or U7442 (N_7442,N_3504,N_3081);
nand U7443 (N_7443,N_3182,N_4161);
or U7444 (N_7444,N_2620,N_3268);
nor U7445 (N_7445,N_3554,N_4816);
nand U7446 (N_7446,N_3677,N_4593);
or U7447 (N_7447,N_3372,N_3680);
nand U7448 (N_7448,N_2838,N_3074);
nor U7449 (N_7449,N_3314,N_4517);
or U7450 (N_7450,N_4023,N_3780);
nand U7451 (N_7451,N_4567,N_4795);
nand U7452 (N_7452,N_2834,N_4740);
nand U7453 (N_7453,N_3322,N_3827);
or U7454 (N_7454,N_4149,N_4843);
or U7455 (N_7455,N_3514,N_4195);
xnor U7456 (N_7456,N_4605,N_4405);
xor U7457 (N_7457,N_3877,N_4308);
nand U7458 (N_7458,N_3398,N_3210);
xnor U7459 (N_7459,N_4334,N_2700);
nand U7460 (N_7460,N_4925,N_3774);
xnor U7461 (N_7461,N_3507,N_3613);
nor U7462 (N_7462,N_4557,N_3312);
or U7463 (N_7463,N_4519,N_4246);
or U7464 (N_7464,N_2773,N_4370);
xnor U7465 (N_7465,N_2621,N_2522);
or U7466 (N_7466,N_4207,N_4140);
nand U7467 (N_7467,N_2747,N_3486);
nand U7468 (N_7468,N_4044,N_3153);
and U7469 (N_7469,N_4206,N_4689);
nand U7470 (N_7470,N_3144,N_2914);
nor U7471 (N_7471,N_4283,N_2879);
nor U7472 (N_7472,N_4381,N_4256);
xnor U7473 (N_7473,N_4060,N_4556);
nor U7474 (N_7474,N_2782,N_2703);
or U7475 (N_7475,N_3550,N_3985);
nand U7476 (N_7476,N_3211,N_4715);
nand U7477 (N_7477,N_4440,N_3600);
and U7478 (N_7478,N_2988,N_3919);
and U7479 (N_7479,N_3248,N_4987);
nand U7480 (N_7480,N_4432,N_3219);
and U7481 (N_7481,N_4612,N_4094);
or U7482 (N_7482,N_2918,N_2893);
xor U7483 (N_7483,N_3338,N_3032);
xnor U7484 (N_7484,N_3710,N_3651);
or U7485 (N_7485,N_4979,N_4467);
nor U7486 (N_7486,N_4563,N_3926);
nand U7487 (N_7487,N_3502,N_4507);
xor U7488 (N_7488,N_3230,N_4578);
nor U7489 (N_7489,N_3800,N_4413);
and U7490 (N_7490,N_4806,N_3268);
xor U7491 (N_7491,N_4261,N_3545);
or U7492 (N_7492,N_3170,N_3113);
or U7493 (N_7493,N_4135,N_3799);
nor U7494 (N_7494,N_4791,N_3739);
nor U7495 (N_7495,N_3358,N_3720);
nor U7496 (N_7496,N_4512,N_3769);
xnor U7497 (N_7497,N_4801,N_3383);
nand U7498 (N_7498,N_4969,N_3195);
and U7499 (N_7499,N_3291,N_3480);
and U7500 (N_7500,N_6251,N_7254);
nand U7501 (N_7501,N_5562,N_6956);
xnor U7502 (N_7502,N_5292,N_5654);
xor U7503 (N_7503,N_6871,N_6283);
nand U7504 (N_7504,N_5201,N_7119);
or U7505 (N_7505,N_7324,N_6490);
or U7506 (N_7506,N_5071,N_6985);
nand U7507 (N_7507,N_5150,N_6700);
and U7508 (N_7508,N_6659,N_6785);
nand U7509 (N_7509,N_7124,N_7084);
and U7510 (N_7510,N_6334,N_6476);
and U7511 (N_7511,N_7306,N_6284);
nand U7512 (N_7512,N_5543,N_5314);
nor U7513 (N_7513,N_5323,N_6382);
nor U7514 (N_7514,N_6606,N_5386);
or U7515 (N_7515,N_6524,N_5009);
and U7516 (N_7516,N_6523,N_5101);
or U7517 (N_7517,N_7095,N_5550);
nand U7518 (N_7518,N_6376,N_6215);
and U7519 (N_7519,N_7260,N_5085);
nand U7520 (N_7520,N_6591,N_7135);
nand U7521 (N_7521,N_5630,N_6001);
nor U7522 (N_7522,N_5560,N_6618);
nand U7523 (N_7523,N_5271,N_5304);
nor U7524 (N_7524,N_6620,N_6444);
or U7525 (N_7525,N_6602,N_5779);
nor U7526 (N_7526,N_5083,N_5475);
nor U7527 (N_7527,N_5269,N_5261);
or U7528 (N_7528,N_6677,N_7116);
nand U7529 (N_7529,N_6290,N_6086);
nor U7530 (N_7530,N_6635,N_7224);
nand U7531 (N_7531,N_6790,N_7017);
nor U7532 (N_7532,N_6625,N_5169);
nand U7533 (N_7533,N_7444,N_6170);
xor U7534 (N_7534,N_6321,N_6247);
and U7535 (N_7535,N_6336,N_7406);
nand U7536 (N_7536,N_6847,N_5871);
nor U7537 (N_7537,N_7189,N_7193);
nor U7538 (N_7538,N_5116,N_6157);
nor U7539 (N_7539,N_7377,N_7239);
and U7540 (N_7540,N_5882,N_6129);
and U7541 (N_7541,N_6220,N_6672);
nand U7542 (N_7542,N_5927,N_6471);
or U7543 (N_7543,N_5581,N_6031);
or U7544 (N_7544,N_6718,N_6588);
nor U7545 (N_7545,N_7191,N_5675);
nand U7546 (N_7546,N_7318,N_6802);
nand U7547 (N_7547,N_7482,N_6356);
and U7548 (N_7548,N_5748,N_7280);
and U7549 (N_7549,N_5342,N_6036);
or U7550 (N_7550,N_6680,N_6813);
nand U7551 (N_7551,N_6204,N_7255);
xnor U7552 (N_7552,N_7344,N_6128);
nand U7553 (N_7553,N_5322,N_7088);
xor U7554 (N_7554,N_7127,N_5552);
xnor U7555 (N_7555,N_7024,N_7461);
or U7556 (N_7556,N_6948,N_5032);
nand U7557 (N_7557,N_7131,N_5426);
and U7558 (N_7558,N_7345,N_5419);
and U7559 (N_7559,N_7400,N_6879);
nor U7560 (N_7560,N_6379,N_5457);
xor U7561 (N_7561,N_5258,N_5872);
and U7562 (N_7562,N_5088,N_6416);
nor U7563 (N_7563,N_6433,N_6870);
or U7564 (N_7564,N_5113,N_6933);
nand U7565 (N_7565,N_5362,N_7258);
and U7566 (N_7566,N_7082,N_7073);
and U7567 (N_7567,N_5856,N_6069);
nand U7568 (N_7568,N_7252,N_5579);
nor U7569 (N_7569,N_6598,N_7081);
nand U7570 (N_7570,N_5337,N_6093);
or U7571 (N_7571,N_7101,N_6633);
nor U7572 (N_7572,N_5517,N_5735);
or U7573 (N_7573,N_7064,N_6551);
nand U7574 (N_7574,N_5483,N_5055);
nor U7575 (N_7575,N_5284,N_5863);
or U7576 (N_7576,N_5325,N_6242);
and U7577 (N_7577,N_6200,N_5809);
or U7578 (N_7578,N_5092,N_7021);
nor U7579 (N_7579,N_6322,N_5665);
nand U7580 (N_7580,N_5217,N_6395);
and U7581 (N_7581,N_7360,N_5107);
and U7582 (N_7582,N_6011,N_6465);
nand U7583 (N_7583,N_6244,N_5839);
and U7584 (N_7584,N_5200,N_5246);
or U7585 (N_7585,N_5173,N_5143);
xor U7586 (N_7586,N_5868,N_6714);
nor U7587 (N_7587,N_5612,N_6197);
and U7588 (N_7588,N_6507,N_7106);
and U7589 (N_7589,N_5710,N_6827);
xor U7590 (N_7590,N_6347,N_5082);
xnor U7591 (N_7591,N_5448,N_5525);
nor U7592 (N_7592,N_6818,N_7477);
nor U7593 (N_7593,N_6357,N_6181);
or U7594 (N_7594,N_6768,N_7375);
nor U7595 (N_7595,N_6090,N_6609);
xnor U7596 (N_7596,N_7464,N_6561);
nand U7597 (N_7597,N_6019,N_7041);
and U7598 (N_7598,N_6469,N_5336);
or U7599 (N_7599,N_6358,N_5123);
nand U7600 (N_7600,N_6300,N_5230);
xor U7601 (N_7601,N_5673,N_5696);
xor U7602 (N_7602,N_5681,N_6450);
or U7603 (N_7603,N_6628,N_5077);
and U7604 (N_7604,N_5764,N_7034);
and U7605 (N_7605,N_5952,N_6994);
nor U7606 (N_7606,N_6041,N_6341);
xor U7607 (N_7607,N_6579,N_6339);
xnor U7608 (N_7608,N_6727,N_5390);
or U7609 (N_7609,N_6509,N_7039);
nand U7610 (N_7610,N_5918,N_7335);
nor U7611 (N_7611,N_7297,N_5470);
nand U7612 (N_7612,N_5734,N_5504);
nand U7613 (N_7613,N_5389,N_5851);
or U7614 (N_7614,N_7353,N_5841);
and U7615 (N_7615,N_5454,N_7080);
xnor U7616 (N_7616,N_5218,N_5741);
xnor U7617 (N_7617,N_5210,N_5640);
or U7618 (N_7618,N_6717,N_5164);
nor U7619 (N_7619,N_5094,N_6151);
nand U7620 (N_7620,N_6073,N_6571);
nor U7621 (N_7621,N_5294,N_7310);
xor U7622 (N_7622,N_5253,N_6867);
xnor U7623 (N_7623,N_6688,N_7069);
nor U7624 (N_7624,N_5761,N_5063);
xnor U7625 (N_7625,N_7229,N_6210);
or U7626 (N_7626,N_7428,N_6886);
nand U7627 (N_7627,N_5720,N_5155);
or U7628 (N_7628,N_5996,N_6246);
or U7629 (N_7629,N_7150,N_5418);
or U7630 (N_7630,N_5511,N_6730);
nand U7631 (N_7631,N_5984,N_5926);
nor U7632 (N_7632,N_5723,N_6682);
nor U7633 (N_7633,N_6616,N_6089);
xor U7634 (N_7634,N_6981,N_7126);
nand U7635 (N_7635,N_5182,N_6820);
and U7636 (N_7636,N_7234,N_5793);
nand U7637 (N_7637,N_6212,N_6259);
nor U7638 (N_7638,N_5042,N_5908);
nor U7639 (N_7639,N_6175,N_7295);
xor U7640 (N_7640,N_6281,N_6350);
or U7641 (N_7641,N_5633,N_7491);
and U7642 (N_7642,N_6883,N_6935);
xor U7643 (N_7643,N_6161,N_7371);
and U7644 (N_7644,N_6008,N_7376);
nand U7645 (N_7645,N_5848,N_6735);
or U7646 (N_7646,N_5672,N_7359);
xor U7647 (N_7647,N_5332,N_5003);
xnor U7648 (N_7648,N_7312,N_7032);
xnor U7649 (N_7649,N_6160,N_5249);
and U7650 (N_7650,N_5351,N_6120);
xor U7651 (N_7651,N_6065,N_6458);
xnor U7652 (N_7652,N_5354,N_6522);
or U7653 (N_7653,N_5225,N_5731);
nor U7654 (N_7654,N_7313,N_5034);
and U7655 (N_7655,N_7432,N_6410);
or U7656 (N_7656,N_5031,N_5431);
xnor U7657 (N_7657,N_6594,N_6343);
and U7658 (N_7658,N_6431,N_5541);
nand U7659 (N_7659,N_6520,N_7165);
nand U7660 (N_7660,N_7108,N_5580);
nand U7661 (N_7661,N_5870,N_5276);
xnor U7662 (N_7662,N_7175,N_5730);
nand U7663 (N_7663,N_6257,N_7060);
nor U7664 (N_7664,N_7070,N_5494);
and U7665 (N_7665,N_6307,N_7144);
xnor U7666 (N_7666,N_6627,N_6393);
and U7667 (N_7667,N_5570,N_7153);
or U7668 (N_7668,N_5174,N_6155);
xnor U7669 (N_7669,N_6560,N_5728);
xnor U7670 (N_7670,N_5035,N_6918);
and U7671 (N_7671,N_6117,N_7217);
xor U7672 (N_7672,N_6459,N_5188);
nor U7673 (N_7673,N_7004,N_7431);
or U7674 (N_7674,N_5762,N_6023);
nand U7675 (N_7675,N_6369,N_5435);
and U7676 (N_7676,N_5537,N_5137);
nor U7677 (N_7677,N_5666,N_6474);
nor U7678 (N_7678,N_5472,N_5905);
nor U7679 (N_7679,N_7192,N_6374);
or U7680 (N_7680,N_5698,N_5566);
nor U7681 (N_7681,N_5833,N_5505);
and U7682 (N_7682,N_5287,N_7307);
and U7683 (N_7683,N_6861,N_5030);
nand U7684 (N_7684,N_5774,N_6952);
nand U7685 (N_7685,N_5760,N_6044);
xnor U7686 (N_7686,N_5007,N_5649);
and U7687 (N_7687,N_6549,N_5135);
or U7688 (N_7688,N_7209,N_7057);
xor U7689 (N_7689,N_7350,N_6998);
and U7690 (N_7690,N_6171,N_6015);
nor U7691 (N_7691,N_5677,N_6983);
xor U7692 (N_7692,N_6608,N_6694);
nand U7693 (N_7693,N_6368,N_5939);
nor U7694 (N_7694,N_5595,N_5587);
xor U7695 (N_7695,N_6185,N_5670);
or U7696 (N_7696,N_5460,N_6791);
nor U7697 (N_7697,N_7040,N_7485);
nor U7698 (N_7698,N_7045,N_5985);
and U7699 (N_7699,N_5692,N_5133);
and U7700 (N_7700,N_5788,N_6763);
nor U7701 (N_7701,N_5158,N_6890);
xnor U7702 (N_7702,N_6586,N_5746);
and U7703 (N_7703,N_5096,N_7365);
or U7704 (N_7704,N_5616,N_6097);
nor U7705 (N_7705,N_6527,N_7190);
and U7706 (N_7706,N_7397,N_5706);
and U7707 (N_7707,N_6853,N_5958);
xnor U7708 (N_7708,N_5020,N_6081);
nand U7709 (N_7709,N_6399,N_5015);
xnor U7710 (N_7710,N_5852,N_6414);
nor U7711 (N_7711,N_6723,N_6868);
or U7712 (N_7712,N_5441,N_7141);
nand U7713 (N_7713,N_6613,N_5726);
xor U7714 (N_7714,N_5103,N_6519);
nand U7715 (N_7715,N_5471,N_6619);
nor U7716 (N_7716,N_6958,N_6388);
xnor U7717 (N_7717,N_6597,N_5530);
and U7718 (N_7718,N_5513,N_6139);
or U7719 (N_7719,N_6378,N_6596);
nand U7720 (N_7720,N_6119,N_6199);
xor U7721 (N_7721,N_7343,N_7257);
nor U7722 (N_7722,N_5213,N_7455);
xor U7723 (N_7723,N_6773,N_6759);
xor U7724 (N_7724,N_6141,N_6367);
xor U7725 (N_7725,N_5816,N_5738);
xor U7726 (N_7726,N_6530,N_7183);
and U7727 (N_7727,N_5144,N_7314);
nor U7728 (N_7728,N_5518,N_5241);
xnor U7729 (N_7729,N_5553,N_7302);
nor U7730 (N_7730,N_7471,N_5674);
xor U7731 (N_7731,N_7061,N_6434);
nor U7732 (N_7732,N_6074,N_5348);
or U7733 (N_7733,N_6990,N_5857);
or U7734 (N_7734,N_7227,N_6850);
nand U7735 (N_7735,N_7188,N_6102);
nor U7736 (N_7736,N_7405,N_6999);
nor U7737 (N_7737,N_6728,N_5736);
or U7738 (N_7738,N_5008,N_5819);
nor U7739 (N_7739,N_5648,N_5501);
xor U7740 (N_7740,N_7319,N_5924);
or U7741 (N_7741,N_6372,N_5281);
xor U7742 (N_7742,N_7468,N_5093);
nor U7743 (N_7743,N_5005,N_6748);
and U7744 (N_7744,N_5199,N_5944);
xor U7745 (N_7745,N_6296,N_5421);
and U7746 (N_7746,N_5686,N_6572);
xnor U7747 (N_7747,N_7240,N_7483);
and U7748 (N_7748,N_7075,N_7074);
nor U7749 (N_7749,N_6068,N_5676);
and U7750 (N_7750,N_7441,N_6510);
or U7751 (N_7751,N_6054,N_5974);
and U7752 (N_7752,N_7391,N_6463);
nor U7753 (N_7753,N_7404,N_6454);
and U7754 (N_7754,N_5953,N_7055);
nand U7755 (N_7755,N_5802,N_6130);
or U7756 (N_7756,N_6188,N_5423);
or U7757 (N_7757,N_7332,N_5668);
xnor U7758 (N_7758,N_5242,N_6592);
and U7759 (N_7759,N_7091,N_5345);
nor U7760 (N_7760,N_7129,N_6814);
or U7761 (N_7761,N_7293,N_6088);
nor U7762 (N_7762,N_7437,N_6266);
or U7763 (N_7763,N_5138,N_5862);
nor U7764 (N_7764,N_6462,N_7166);
nand U7765 (N_7765,N_5998,N_5955);
nor U7766 (N_7766,N_7452,N_6299);
and U7767 (N_7767,N_7311,N_5338);
nand U7768 (N_7768,N_6685,N_6754);
xor U7769 (N_7769,N_6042,N_6764);
or U7770 (N_7770,N_6062,N_5558);
xor U7771 (N_7771,N_5492,N_5982);
nand U7772 (N_7772,N_6538,N_6309);
and U7773 (N_7773,N_7351,N_6180);
nor U7774 (N_7774,N_5346,N_5983);
nand U7775 (N_7775,N_7076,N_7194);
and U7776 (N_7776,N_5778,N_7361);
nor U7777 (N_7777,N_5388,N_6902);
nand U7778 (N_7778,N_6734,N_6699);
and U7779 (N_7779,N_7147,N_7220);
and U7780 (N_7780,N_6061,N_5374);
and U7781 (N_7781,N_7120,N_6294);
or U7782 (N_7782,N_5873,N_6430);
nor U7783 (N_7783,N_6722,N_7243);
and U7784 (N_7784,N_5263,N_6788);
xor U7785 (N_7785,N_7364,N_5885);
xor U7786 (N_7786,N_6912,N_6456);
and U7787 (N_7787,N_5075,N_6110);
or U7788 (N_7788,N_7270,N_7264);
nor U7789 (N_7789,N_6240,N_6529);
or U7790 (N_7790,N_6265,N_5383);
nand U7791 (N_7791,N_6169,N_6154);
nand U7792 (N_7792,N_6192,N_5540);
nor U7793 (N_7793,N_6516,N_6252);
xor U7794 (N_7794,N_6955,N_6532);
xnor U7795 (N_7795,N_6479,N_6052);
nand U7796 (N_7796,N_5160,N_5806);
or U7797 (N_7797,N_6605,N_6131);
xnor U7798 (N_7798,N_6420,N_5946);
or U7799 (N_7799,N_6359,N_7230);
xor U7800 (N_7800,N_7445,N_7176);
nor U7801 (N_7801,N_6673,N_6118);
and U7802 (N_7802,N_5514,N_5745);
nand U7803 (N_7803,N_6238,N_5073);
and U7804 (N_7804,N_6231,N_7203);
nand U7805 (N_7805,N_6652,N_5744);
nand U7806 (N_7806,N_5527,N_7473);
xnor U7807 (N_7807,N_5299,N_6977);
and U7808 (N_7808,N_5010,N_6540);
xor U7809 (N_7809,N_7372,N_5267);
nand U7810 (N_7810,N_5500,N_5789);
or U7811 (N_7811,N_7366,N_5151);
xor U7812 (N_7812,N_5070,N_7138);
nor U7813 (N_7813,N_7218,N_6492);
xnor U7814 (N_7814,N_5963,N_6817);
and U7815 (N_7815,N_6397,N_5175);
nand U7816 (N_7816,N_5215,N_7370);
nor U7817 (N_7817,N_7182,N_6770);
nand U7818 (N_7818,N_5878,N_5936);
nor U7819 (N_7819,N_7448,N_6274);
and U7820 (N_7820,N_6101,N_7459);
or U7821 (N_7821,N_5100,N_6582);
and U7822 (N_7822,N_6288,N_7003);
nor U7823 (N_7823,N_7015,N_6761);
xnor U7824 (N_7824,N_5165,N_7282);
and U7825 (N_7825,N_6396,N_7490);
xor U7826 (N_7826,N_6317,N_6403);
nand U7827 (N_7827,N_7300,N_6846);
or U7828 (N_7828,N_6037,N_6924);
or U7829 (N_7829,N_7179,N_5154);
nand U7830 (N_7830,N_6711,N_6352);
nor U7831 (N_7831,N_6829,N_5987);
nand U7832 (N_7832,N_6013,N_5995);
nand U7833 (N_7833,N_7454,N_5221);
or U7834 (N_7834,N_5080,N_5349);
and U7835 (N_7835,N_5198,N_6387);
or U7836 (N_7836,N_6795,N_7164);
nor U7837 (N_7837,N_5922,N_6230);
and U7838 (N_7838,N_5324,N_7296);
nor U7839 (N_7839,N_5752,N_7232);
nor U7840 (N_7840,N_5656,N_7102);
and U7841 (N_7841,N_6452,N_6812);
or U7842 (N_7842,N_5397,N_5523);
and U7843 (N_7843,N_5476,N_5392);
and U7844 (N_7844,N_5934,N_7121);
or U7845 (N_7845,N_6320,N_6664);
nor U7846 (N_7846,N_5273,N_5443);
xor U7847 (N_7847,N_6781,N_5468);
and U7848 (N_7848,N_6866,N_6894);
nand U7849 (N_7849,N_5171,N_7130);
or U7850 (N_7850,N_7425,N_5810);
nand U7851 (N_7851,N_6132,N_7309);
and U7852 (N_7852,N_5787,N_6159);
nor U7853 (N_7853,N_5438,N_6934);
nor U7854 (N_7854,N_5847,N_5727);
nand U7855 (N_7855,N_5949,N_6544);
nor U7856 (N_7856,N_7422,N_5380);
nor U7857 (N_7857,N_6440,N_5347);
nor U7858 (N_7858,N_5220,N_7291);
and U7859 (N_7859,N_5621,N_5758);
xor U7860 (N_7860,N_6639,N_5311);
and U7861 (N_7861,N_7388,N_6280);
or U7862 (N_7862,N_6852,N_6679);
xnor U7863 (N_7863,N_6737,N_6856);
nand U7864 (N_7864,N_6874,N_6205);
nand U7865 (N_7865,N_6144,N_6292);
xnor U7866 (N_7866,N_5965,N_5339);
and U7867 (N_7867,N_7159,N_6769);
nand U7868 (N_7868,N_5854,N_6655);
nand U7869 (N_7869,N_5194,N_6908);
xor U7870 (N_7870,N_6354,N_6615);
xor U7871 (N_7871,N_6111,N_5486);
xnor U7872 (N_7872,N_5428,N_5573);
xnor U7873 (N_7873,N_6897,N_6899);
or U7874 (N_7874,N_6276,N_7418);
nor U7875 (N_7875,N_5202,N_6941);
nand U7876 (N_7876,N_7167,N_5935);
or U7877 (N_7877,N_7408,N_6056);
or U7878 (N_7878,N_5289,N_5663);
and U7879 (N_7879,N_7204,N_6642);
nand U7880 (N_7880,N_5288,N_6206);
and U7881 (N_7881,N_5685,N_5972);
and U7882 (N_7882,N_5180,N_7334);
or U7883 (N_7883,N_5260,N_6303);
nand U7884 (N_7884,N_5529,N_6910);
xor U7885 (N_7885,N_5781,N_6211);
and U7886 (N_7886,N_7356,N_6464);
xnor U7887 (N_7887,N_6701,N_6049);
and U7888 (N_7888,N_6145,N_6876);
and U7889 (N_7889,N_7256,N_5130);
nor U7890 (N_7890,N_7137,N_5193);
xnor U7891 (N_7891,N_6491,N_6822);
or U7892 (N_7892,N_5639,N_7488);
xnor U7893 (N_7893,N_5684,N_6992);
or U7894 (N_7894,N_6423,N_5427);
nand U7895 (N_7895,N_5398,N_5312);
and U7896 (N_7896,N_6961,N_7093);
or U7897 (N_7897,N_6928,N_5941);
xnor U7898 (N_7898,N_5384,N_5821);
and U7899 (N_7899,N_6810,N_5757);
or U7900 (N_7900,N_6564,N_5124);
xor U7901 (N_7901,N_5994,N_7265);
nand U7902 (N_7902,N_5526,N_5317);
and U7903 (N_7903,N_6649,N_5588);
nand U7904 (N_7904,N_5464,N_6498);
nand U7905 (N_7905,N_6483,N_7494);
nor U7906 (N_7906,N_6381,N_6715);
nor U7907 (N_7907,N_5724,N_6162);
xor U7908 (N_7908,N_6239,N_5843);
nor U7909 (N_7909,N_7052,N_6228);
nand U7910 (N_7910,N_6548,N_6721);
and U7911 (N_7911,N_5027,N_6756);
xor U7912 (N_7912,N_5229,N_5742);
nand U7913 (N_7913,N_6712,N_6392);
or U7914 (N_7914,N_6126,N_6332);
or U7915 (N_7915,N_5866,N_5382);
or U7916 (N_7916,N_6653,N_7429);
xor U7917 (N_7917,N_5831,N_7434);
and U7918 (N_7918,N_5282,N_6531);
or U7919 (N_7919,N_5330,N_7417);
and U7920 (N_7920,N_6318,N_5458);
nand U7921 (N_7921,N_7273,N_5571);
and U7922 (N_7922,N_6766,N_6346);
nor U7923 (N_7923,N_5480,N_7235);
or U7924 (N_7924,N_6344,N_6760);
nor U7925 (N_7925,N_7215,N_5968);
and U7926 (N_7926,N_6047,N_5232);
nand U7927 (N_7927,N_5086,N_6789);
or U7928 (N_7928,N_7259,N_6574);
and U7929 (N_7929,N_6226,N_6408);
xnor U7930 (N_7930,N_5000,N_6092);
nand U7931 (N_7931,N_6805,N_5799);
or U7932 (N_7932,N_6143,N_6777);
nor U7933 (N_7933,N_5148,N_5061);
nor U7934 (N_7934,N_6966,N_6447);
nand U7935 (N_7935,N_6187,N_5106);
and U7936 (N_7936,N_6738,N_6893);
or U7937 (N_7937,N_5978,N_6741);
xnor U7938 (N_7938,N_6308,N_5114);
and U7939 (N_7939,N_5224,N_6502);
xnor U7940 (N_7940,N_6708,N_6786);
and U7941 (N_7941,N_5084,N_5433);
and U7942 (N_7942,N_6799,N_5642);
or U7943 (N_7943,N_5628,N_5899);
and U7944 (N_7944,N_6815,N_7089);
or U7945 (N_7945,N_6293,N_7247);
xnor U7946 (N_7946,N_6198,N_5813);
nor U7947 (N_7947,N_5016,N_5247);
xnor U7948 (N_7948,N_6070,N_5928);
xor U7949 (N_7949,N_6124,N_6064);
nand U7950 (N_7950,N_6646,N_6569);
xor U7951 (N_7951,N_5274,N_7451);
nor U7952 (N_7952,N_6437,N_6631);
nand U7953 (N_7953,N_5313,N_6455);
and U7954 (N_7954,N_5373,N_5531);
nor U7955 (N_7955,N_5358,N_6179);
or U7956 (N_7956,N_5547,N_6427);
nor U7957 (N_7957,N_6168,N_5381);
or U7958 (N_7958,N_6807,N_6604);
nand U7959 (N_7959,N_6072,N_5679);
xor U7960 (N_7960,N_6050,N_6315);
or U7961 (N_7961,N_5490,N_7236);
xor U7962 (N_7962,N_6243,N_7357);
or U7963 (N_7963,N_5569,N_5259);
nand U7964 (N_7964,N_6740,N_6059);
or U7965 (N_7965,N_6800,N_6190);
nand U7966 (N_7966,N_5655,N_5617);
xor U7967 (N_7967,N_6978,N_5244);
xnor U7968 (N_7968,N_5750,N_6377);
nor U7969 (N_7969,N_5894,N_6643);
xor U7970 (N_7970,N_6589,N_6636);
or U7971 (N_7971,N_5089,N_7008);
xor U7972 (N_7972,N_5765,N_6443);
nor U7973 (N_7973,N_7284,N_7413);
and U7974 (N_7974,N_6645,N_6150);
and U7975 (N_7975,N_6552,N_6954);
or U7976 (N_7976,N_7379,N_5228);
nor U7977 (N_7977,N_5658,N_5950);
nand U7978 (N_7978,N_5783,N_5461);
xnor U7979 (N_7979,N_5522,N_6406);
nor U7980 (N_7980,N_6385,N_6104);
and U7981 (N_7981,N_6929,N_5700);
nand U7982 (N_7982,N_5129,N_6135);
and U7983 (N_7983,N_6327,N_5515);
or U7984 (N_7984,N_7207,N_7068);
nor U7985 (N_7985,N_6271,N_5499);
xor U7986 (N_7986,N_6779,N_6468);
nor U7987 (N_7987,N_5262,N_5119);
nand U7988 (N_7988,N_7022,N_6067);
and U7989 (N_7989,N_7440,N_6896);
or U7990 (N_7990,N_7027,N_7113);
nor U7991 (N_7991,N_6140,N_6980);
nor U7992 (N_7992,N_6512,N_5858);
nand U7993 (N_7993,N_5167,N_6648);
or U7994 (N_7994,N_5601,N_5545);
and U7995 (N_7995,N_6796,N_6967);
and U7996 (N_7996,N_6888,N_7132);
or U7997 (N_7997,N_5754,N_5917);
xor U7998 (N_7998,N_5297,N_5662);
and U7999 (N_7999,N_6287,N_6845);
nor U8000 (N_8000,N_5377,N_6422);
or U8001 (N_8001,N_5801,N_6710);
and U8002 (N_8002,N_5364,N_6996);
xor U8003 (N_8003,N_5590,N_5405);
xor U8004 (N_8004,N_6862,N_7325);
nor U8005 (N_8005,N_6250,N_7005);
nand U8006 (N_8006,N_5062,N_6881);
xor U8007 (N_8007,N_6503,N_7030);
nand U8008 (N_8008,N_5869,N_6725);
xnor U8009 (N_8009,N_5737,N_6138);
or U8010 (N_8010,N_6331,N_6457);
or U8011 (N_8011,N_7415,N_6745);
nand U8012 (N_8012,N_5659,N_7154);
xnor U8013 (N_8013,N_7096,N_6706);
xor U8014 (N_8014,N_6546,N_7480);
xnor U8015 (N_8015,N_7383,N_7267);
and U8016 (N_8016,N_5713,N_7042);
xor U8017 (N_8017,N_6445,N_5118);
nand U8018 (N_8018,N_7056,N_5127);
or U8019 (N_8019,N_7160,N_7063);
or U8020 (N_8020,N_6661,N_5308);
xor U8021 (N_8021,N_6323,N_6937);
xnor U8022 (N_8022,N_6662,N_7079);
and U8023 (N_8023,N_5614,N_6094);
or U8024 (N_8024,N_7245,N_6500);
nor U8025 (N_8025,N_5278,N_7281);
xor U8026 (N_8026,N_6329,N_6451);
or U8027 (N_8027,N_6484,N_6114);
nand U8028 (N_8028,N_5842,N_6448);
nand U8029 (N_8029,N_5076,N_6148);
nor U8030 (N_8030,N_6057,N_5520);
xor U8031 (N_8031,N_7143,N_5691);
and U8032 (N_8032,N_6217,N_5178);
xor U8033 (N_8033,N_5265,N_6480);
nor U8034 (N_8034,N_5102,N_7072);
nor U8035 (N_8035,N_6914,N_5768);
or U8036 (N_8036,N_6555,N_5533);
or U8037 (N_8037,N_7497,N_5333);
or U8038 (N_8038,N_6325,N_6577);
or U8039 (N_8039,N_6165,N_6963);
nand U8040 (N_8040,N_5067,N_6634);
nor U8041 (N_8041,N_6384,N_6732);
or U8042 (N_8042,N_6536,N_6953);
xnor U8043 (N_8043,N_6166,N_5524);
xnor U8044 (N_8044,N_5999,N_5855);
xor U8045 (N_8045,N_7155,N_5371);
nor U8046 (N_8046,N_5290,N_7331);
nor U8047 (N_8047,N_6203,N_5185);
nor U8048 (N_8048,N_5181,N_7195);
nand U8049 (N_8049,N_5785,N_5992);
nand U8050 (N_8050,N_6207,N_6473);
nand U8051 (N_8051,N_5367,N_5594);
or U8052 (N_8052,N_5065,N_5420);
xor U8053 (N_8053,N_5238,N_7048);
or U8054 (N_8054,N_7341,N_5850);
and U8055 (N_8055,N_7149,N_6747);
nand U8056 (N_8056,N_6731,N_5052);
and U8057 (N_8057,N_6167,N_7384);
and U8058 (N_8058,N_5867,N_5407);
nor U8059 (N_8059,N_6919,N_5945);
nor U8060 (N_8060,N_5404,N_6622);
or U8061 (N_8061,N_5931,N_5548);
nand U8062 (N_8062,N_7198,N_6957);
or U8063 (N_8063,N_6453,N_6663);
nor U8064 (N_8064,N_5179,N_6525);
and U8065 (N_8065,N_5702,N_6882);
nand U8066 (N_8066,N_6153,N_6578);
and U8067 (N_8067,N_6348,N_5183);
nor U8068 (N_8068,N_5660,N_5033);
or U8069 (N_8069,N_5823,N_5112);
and U8070 (N_8070,N_6736,N_6917);
or U8071 (N_8071,N_7067,N_6017);
xor U8072 (N_8072,N_5309,N_5141);
xor U8073 (N_8073,N_5449,N_6194);
or U8074 (N_8074,N_5399,N_7268);
and U8075 (N_8075,N_5719,N_6373);
nand U8076 (N_8076,N_6518,N_6146);
nand U8077 (N_8077,N_5361,N_6696);
nor U8078 (N_8078,N_6563,N_5874);
nor U8079 (N_8079,N_7094,N_6945);
nor U8080 (N_8080,N_6107,N_5487);
nand U8081 (N_8081,N_5159,N_6301);
xnor U8082 (N_8082,N_6782,N_6028);
and U8083 (N_8083,N_7304,N_7185);
nor U8084 (N_8084,N_5890,N_6671);
and U8085 (N_8085,N_7387,N_7274);
nand U8086 (N_8086,N_6439,N_7327);
or U8087 (N_8087,N_6164,N_6825);
nor U8088 (N_8088,N_5943,N_6380);
or U8089 (N_8089,N_5747,N_5604);
and U8090 (N_8090,N_5017,N_6261);
nand U8091 (N_8091,N_5266,N_6971);
nand U8092 (N_8092,N_7301,N_5385);
nand U8093 (N_8093,N_6219,N_5189);
xnor U8094 (N_8094,N_6824,N_5800);
nor U8095 (N_8095,N_6931,N_6657);
and U8096 (N_8096,N_5453,N_6900);
xnor U8097 (N_8097,N_5883,N_6232);
nand U8098 (N_8098,N_5714,N_5546);
nand U8099 (N_8099,N_6614,N_6505);
xor U8100 (N_8100,N_6920,N_6840);
or U8101 (N_8101,N_7180,N_7083);
and U8102 (N_8102,N_5919,N_6121);
xor U8103 (N_8103,N_6689,N_6803);
xnor U8104 (N_8104,N_5041,N_5519);
and U8105 (N_8105,N_6809,N_6302);
nor U8106 (N_8106,N_5416,N_7177);
nand U8107 (N_8107,N_7277,N_6202);
nor U8108 (N_8108,N_5425,N_7012);
xnor U8109 (N_8109,N_5913,N_6488);
and U8110 (N_8110,N_5990,N_7202);
nand U8111 (N_8111,N_7107,N_6547);
nor U8112 (N_8112,N_6418,N_7462);
and U8113 (N_8113,N_6461,N_5156);
or U8114 (N_8114,N_5310,N_6136);
nand U8115 (N_8115,N_6621,N_7037);
xnor U8116 (N_8116,N_6078,N_6310);
and U8117 (N_8117,N_7299,N_6035);
nand U8118 (N_8118,N_7054,N_5450);
and U8119 (N_8119,N_6103,N_5192);
and U8120 (N_8120,N_5319,N_5722);
and U8121 (N_8121,N_5328,N_5068);
nor U8122 (N_8122,N_6264,N_6972);
or U8123 (N_8123,N_5915,N_6066);
nor U8124 (N_8124,N_6641,N_5979);
or U8125 (N_8125,N_5301,N_7389);
nand U8126 (N_8126,N_5911,N_6386);
or U8127 (N_8127,N_5976,N_6316);
xor U8128 (N_8128,N_5286,N_7090);
or U8129 (N_8129,N_6864,N_6869);
and U8130 (N_8130,N_7077,N_5775);
or U8131 (N_8131,N_7380,N_6709);
and U8132 (N_8132,N_5997,N_5769);
nor U8133 (N_8133,N_5631,N_6364);
and U8134 (N_8134,N_5632,N_5623);
nor U8135 (N_8135,N_5794,N_7285);
xor U8136 (N_8136,N_6409,N_5251);
xnor U8137 (N_8137,N_6979,N_7340);
nor U8138 (N_8138,N_7251,N_6811);
or U8139 (N_8139,N_6003,N_7453);
or U8140 (N_8140,N_6757,N_6535);
or U8141 (N_8141,N_6637,N_5969);
nor U8142 (N_8142,N_5142,N_5610);
and U8143 (N_8143,N_7363,N_7421);
nor U8144 (N_8144,N_5341,N_5971);
and U8145 (N_8145,N_7495,N_5937);
and U8146 (N_8146,N_5066,N_5549);
and U8147 (N_8147,N_6030,N_7290);
nand U8148 (N_8148,N_5961,N_5759);
or U8149 (N_8149,N_5613,N_5396);
nor U8150 (N_8150,N_5393,N_6400);
or U8151 (N_8151,N_6580,N_5131);
xor U8152 (N_8152,N_5814,N_6865);
or U8153 (N_8153,N_5152,N_6305);
nor U8154 (N_8154,N_6877,N_6149);
or U8155 (N_8155,N_5898,N_6593);
and U8156 (N_8156,N_5844,N_6060);
xnor U8157 (N_8157,N_5805,N_6511);
nand U8158 (N_8158,N_7349,N_7122);
or U8159 (N_8159,N_5295,N_6964);
nor U8160 (N_8160,N_7470,N_6903);
and U8161 (N_8161,N_6987,N_7211);
and U8162 (N_8162,N_5484,N_7223);
nor U8163 (N_8163,N_7374,N_5442);
and U8164 (N_8164,N_6975,N_6022);
nor U8165 (N_8165,N_7049,N_6611);
nand U8166 (N_8166,N_6142,N_5766);
nor U8167 (N_8167,N_6177,N_5022);
xnor U8168 (N_8168,N_5140,N_6833);
nand U8169 (N_8169,N_6083,N_7146);
nand U8170 (N_8170,N_7336,N_6719);
and U8171 (N_8171,N_7033,N_6043);
nor U8172 (N_8172,N_7184,N_5277);
or U8173 (N_8173,N_5561,N_6319);
nor U8174 (N_8174,N_6984,N_6670);
or U8175 (N_8175,N_5584,N_5818);
xnor U8176 (N_8176,N_6201,N_5074);
xnor U8177 (N_8177,N_6733,N_5320);
xnor U8178 (N_8178,N_5593,N_5824);
xor U8179 (N_8179,N_5506,N_5884);
nand U8180 (N_8180,N_6134,N_7411);
nor U8181 (N_8181,N_6533,N_6255);
and U8182 (N_8182,N_6355,N_5059);
or U8183 (N_8183,N_5387,N_5410);
xnor U8184 (N_8184,N_7355,N_6746);
or U8185 (N_8185,N_7053,N_6435);
nand U8186 (N_8186,N_5028,N_5634);
xnor U8187 (N_8187,N_6394,N_5716);
nand U8188 (N_8188,N_6291,N_6233);
nor U8189 (N_8189,N_7424,N_7435);
nor U8190 (N_8190,N_5763,N_6550);
nor U8191 (N_8191,N_7222,N_7446);
nor U8192 (N_8192,N_5563,N_6806);
nor U8193 (N_8193,N_7469,N_6189);
nand U8194 (N_8194,N_5528,N_5248);
xnor U8195 (N_8195,N_5694,N_6046);
xor U8196 (N_8196,N_5697,N_5240);
or U8197 (N_8197,N_6940,N_6314);
nand U8198 (N_8198,N_6925,N_7020);
xor U8199 (N_8199,N_5196,N_5050);
nand U8200 (N_8200,N_6236,N_6109);
nor U8201 (N_8201,N_5647,N_5272);
xor U8202 (N_8202,N_7142,N_6724);
or U8203 (N_8203,N_5807,N_5556);
nand U8204 (N_8204,N_7219,N_5184);
or U8205 (N_8205,N_7499,N_5233);
nand U8206 (N_8206,N_5469,N_5053);
and U8207 (N_8207,N_5211,N_5018);
nor U8208 (N_8208,N_6947,N_7271);
and U8209 (N_8209,N_5892,N_5516);
and U8210 (N_8210,N_6105,N_5597);
xnor U8211 (N_8211,N_6687,N_6221);
or U8212 (N_8212,N_5845,N_7486);
or U8213 (N_8213,N_7029,N_5365);
nor U8214 (N_8214,N_6419,N_7023);
or U8215 (N_8215,N_5583,N_5564);
or U8216 (N_8216,N_6951,N_7476);
and U8217 (N_8217,N_6880,N_6742);
and U8218 (N_8218,N_6997,N_6024);
nand U8219 (N_8219,N_5717,N_5749);
or U8220 (N_8220,N_6916,N_7262);
or U8221 (N_8221,N_7298,N_5835);
and U8222 (N_8222,N_7316,N_6487);
and U8223 (N_8223,N_5575,N_6108);
nand U8224 (N_8224,N_6389,N_5413);
xor U8225 (N_8225,N_7221,N_7399);
xnor U8226 (N_8226,N_5740,N_5861);
or U8227 (N_8227,N_6581,N_7169);
or U8228 (N_8228,N_5832,N_7199);
xor U8229 (N_8229,N_6911,N_5417);
xnor U8230 (N_8230,N_7438,N_6630);
nor U8231 (N_8231,N_6324,N_6335);
or U8232 (N_8232,N_7342,N_7161);
or U8233 (N_8233,N_6923,N_5712);
nor U8234 (N_8234,N_6601,N_5255);
and U8235 (N_8235,N_6909,N_6675);
nand U8236 (N_8236,N_6429,N_7303);
nor U8237 (N_8237,N_6018,N_5914);
nand U8238 (N_8238,N_6904,N_7062);
and U8239 (N_8239,N_7329,N_6286);
or U8240 (N_8240,N_6055,N_6797);
nand U8241 (N_8241,N_7289,N_7019);
or U8242 (N_8242,N_6186,N_7288);
and U8243 (N_8243,N_5326,N_7046);
nor U8244 (N_8244,N_7481,N_5236);
nand U8245 (N_8245,N_7139,N_7463);
nor U8246 (N_8246,N_6794,N_6668);
nor U8247 (N_8247,N_6585,N_7287);
xnor U8248 (N_8248,N_7278,N_5923);
nand U8249 (N_8249,N_6176,N_7407);
and U8250 (N_8250,N_6021,N_5432);
nand U8251 (N_8251,N_7117,N_7458);
and U8252 (N_8252,N_6330,N_5859);
xor U8253 (N_8253,N_5970,N_6025);
xor U8254 (N_8254,N_6496,N_7443);
and U8255 (N_8255,N_5491,N_5400);
and U8256 (N_8256,N_6542,N_6277);
nor U8257 (N_8257,N_5002,N_5572);
and U8258 (N_8258,N_5452,N_6426);
or U8259 (N_8259,N_5991,N_6716);
xnor U8260 (N_8260,N_7460,N_6559);
or U8261 (N_8261,N_6472,N_5437);
nand U8262 (N_8262,N_6995,N_5368);
and U8263 (N_8263,N_5718,N_5353);
or U8264 (N_8264,N_5207,N_7231);
or U8265 (N_8265,N_6949,N_5609);
nand U8266 (N_8266,N_5576,N_6891);
and U8267 (N_8267,N_5864,N_6849);
or U8268 (N_8268,N_7128,N_5134);
nand U8269 (N_8269,N_7346,N_6541);
nand U8270 (N_8270,N_6854,N_7286);
and U8271 (N_8271,N_6349,N_5840);
nor U8272 (N_8272,N_7242,N_6943);
xor U8273 (N_8273,N_6944,N_6184);
or U8274 (N_8274,N_5836,N_6583);
and U8275 (N_8275,N_5128,N_6263);
and U8276 (N_8276,N_7416,N_5837);
nor U8277 (N_8277,N_5190,N_7279);
nor U8278 (N_8278,N_6428,N_7447);
and U8279 (N_8279,N_7315,N_5988);
nand U8280 (N_8280,N_5701,N_6986);
xor U8281 (N_8281,N_6702,N_6029);
xor U8282 (N_8282,N_5904,N_6587);
nand U8283 (N_8283,N_6793,N_6241);
or U8284 (N_8284,N_6223,N_6517);
or U8285 (N_8285,N_5036,N_6573);
xnor U8286 (N_8286,N_7333,N_5777);
nand U8287 (N_8287,N_5829,N_5257);
or U8288 (N_8288,N_5125,N_7171);
and U8289 (N_8289,N_6858,N_5705);
xor U8290 (N_8290,N_7233,N_6885);
or U8291 (N_8291,N_5669,N_6125);
or U8292 (N_8292,N_6258,N_7100);
nand U8293 (N_8293,N_5975,N_6798);
or U8294 (N_8294,N_5708,N_6402);
nor U8295 (N_8295,N_6304,N_5045);
or U8296 (N_8296,N_6855,N_5478);
nor U8297 (N_8297,N_5507,N_5796);
xor U8298 (N_8298,N_7237,N_5715);
nand U8299 (N_8299,N_6513,N_7394);
nor U8300 (N_8300,N_6638,N_5466);
nand U8301 (N_8301,N_5860,N_5268);
and U8302 (N_8302,N_5095,N_5977);
or U8303 (N_8303,N_6836,N_5098);
and U8304 (N_8304,N_6600,N_6629);
nor U8305 (N_8305,N_7133,N_5402);
nand U8306 (N_8306,N_7367,N_6697);
or U8307 (N_8307,N_7186,N_7044);
xor U8308 (N_8308,N_7347,N_5474);
nor U8309 (N_8309,N_5641,N_5372);
nor U8310 (N_8310,N_7283,N_5245);
nor U8311 (N_8311,N_5037,N_7014);
or U8312 (N_8312,N_6506,N_5815);
nand U8313 (N_8313,N_6640,N_7158);
and U8314 (N_8314,N_5895,N_6493);
xnor U8315 (N_8315,N_5582,N_5544);
xnor U8316 (N_8316,N_5542,N_6010);
xnor U8317 (N_8317,N_7071,N_6216);
xnor U8318 (N_8318,N_6819,N_6767);
xor U8319 (N_8319,N_6401,N_5252);
nand U8320 (N_8320,N_5149,N_6306);
and U8321 (N_8321,N_6844,N_7226);
and U8322 (N_8322,N_5600,N_6568);
and U8323 (N_8323,N_7426,N_6051);
nor U8324 (N_8324,N_6275,N_5429);
nand U8325 (N_8325,N_6993,N_5219);
or U8326 (N_8326,N_7410,N_7358);
or U8327 (N_8327,N_5555,N_7362);
nand U8328 (N_8328,N_5683,N_6834);
xor U8329 (N_8329,N_7378,N_6556);
nor U8330 (N_8330,N_5875,N_5574);
or U8331 (N_8331,N_5479,N_5004);
nor U8332 (N_8332,N_5162,N_5139);
nor U8333 (N_8333,N_6002,N_5485);
xor U8334 (N_8334,N_5456,N_7419);
xnor U8335 (N_8335,N_6566,N_7498);
xor U8336 (N_8336,N_5880,N_5462);
or U8337 (N_8337,N_6921,N_5006);
or U8338 (N_8338,N_6686,N_6256);
nand U8339 (N_8339,N_5916,N_5147);
xor U8340 (N_8340,N_5495,N_5038);
or U8341 (N_8341,N_7487,N_6539);
xor U8342 (N_8342,N_5090,N_5772);
nor U8343 (N_8343,N_5424,N_6780);
and U8344 (N_8344,N_5605,N_5729);
nor U8345 (N_8345,N_5414,N_5058);
or U8346 (N_8346,N_5315,N_5334);
and U8347 (N_8347,N_6053,N_5115);
nand U8348 (N_8348,N_5770,N_6099);
nand U8349 (N_8349,N_5619,N_6875);
nand U8350 (N_8350,N_5279,N_6654);
nand U8351 (N_8351,N_6494,N_6749);
nand U8352 (N_8352,N_5043,N_6595);
and U8353 (N_8353,N_6783,N_6938);
xor U8354 (N_8354,N_6489,N_5060);
or U8355 (N_8355,N_5316,N_6751);
nand U8356 (N_8356,N_5132,N_5707);
xor U8357 (N_8357,N_6370,N_5909);
nand U8358 (N_8358,N_6693,N_5191);
or U8359 (N_8359,N_5340,N_6224);
nor U8360 (N_8360,N_6270,N_7162);
or U8361 (N_8361,N_6851,N_6405);
nor U8362 (N_8362,N_7272,N_6326);
and U8363 (N_8363,N_5502,N_5108);
nor U8364 (N_8364,N_6020,N_5782);
nand U8365 (N_8365,N_6651,N_5888);
nor U8366 (N_8366,N_6801,N_6353);
nor U8367 (N_8367,N_7238,N_5512);
xor U8368 (N_8368,N_6843,N_6421);
or U8369 (N_8369,N_6739,N_5048);
xor U8370 (N_8370,N_7013,N_5305);
xor U8371 (N_8371,N_7112,N_6262);
or U8372 (N_8372,N_5329,N_7385);
nor U8373 (N_8373,N_6182,N_6475);
and U8374 (N_8374,N_6082,N_6599);
nor U8375 (N_8375,N_6080,N_5168);
nor U8376 (N_8376,N_7493,N_6222);
nand U8377 (N_8377,N_5026,N_5157);
nand U8378 (N_8378,N_7002,N_7086);
or U8379 (N_8379,N_5363,N_5493);
nor U8380 (N_8380,N_6758,N_5568);
xnor U8381 (N_8381,N_6158,N_7492);
nor U8382 (N_8382,N_6841,N_6009);
nand U8383 (N_8383,N_6006,N_5439);
nor U8384 (N_8384,N_6857,N_7205);
or U8385 (N_8385,N_5589,N_5645);
nor U8386 (N_8386,N_6227,N_6973);
xnor U8387 (N_8387,N_5830,N_6991);
xnor U8388 (N_8388,N_6084,N_7320);
nand U8389 (N_8389,N_7196,N_6163);
xnor U8390 (N_8390,N_7420,N_5817);
nor U8391 (N_8391,N_7038,N_7369);
nor U8392 (N_8392,N_6831,N_5001);
and U8393 (N_8393,N_6665,N_6860);
or U8394 (N_8394,N_7085,N_6338);
or U8395 (N_8395,N_5535,N_5902);
nand U8396 (N_8396,N_6750,N_5834);
nor U8397 (N_8397,N_7208,N_6534);
and U8398 (N_8398,N_7187,N_6026);
or U8399 (N_8399,N_6650,N_5331);
nor U8400 (N_8400,N_5488,N_5733);
nand U8401 (N_8401,N_6345,N_5293);
and U8402 (N_8402,N_5577,N_6575);
nand U8403 (N_8403,N_5693,N_6229);
or U8404 (N_8404,N_6942,N_6930);
and U8405 (N_8405,N_7148,N_7479);
xnor U8406 (N_8406,N_5234,N_7430);
and U8407 (N_8407,N_6989,N_6058);
nor U8408 (N_8408,N_5811,N_5667);
xnor U8409 (N_8409,N_5047,N_6774);
or U8410 (N_8410,N_5237,N_6778);
nand U8411 (N_8411,N_6837,N_6183);
nand U8412 (N_8412,N_7475,N_5951);
nand U8413 (N_8413,N_5767,N_5912);
nand U8414 (N_8414,N_6085,N_7178);
and U8415 (N_8415,N_7047,N_5622);
xor U8416 (N_8416,N_6122,N_5629);
and U8417 (N_8417,N_6039,N_6075);
xor U8418 (N_8418,N_6460,N_7382);
and U8419 (N_8419,N_5285,N_6040);
or U8420 (N_8420,N_5565,N_5153);
nor U8421 (N_8421,N_6683,N_6884);
or U8422 (N_8422,N_5369,N_6950);
or U8423 (N_8423,N_5509,N_7423);
nor U8424 (N_8424,N_5097,N_6842);
xor U8425 (N_8425,N_5921,N_6407);
and U8426 (N_8426,N_6442,N_5161);
nand U8427 (N_8427,N_7140,N_6932);
xnor U8428 (N_8428,N_6784,N_6100);
xor U8429 (N_8429,N_5534,N_6106);
or U8430 (N_8430,N_5620,N_6295);
xor U8431 (N_8431,N_6477,N_5624);
nor U8432 (N_8432,N_6333,N_5447);
xnor U8433 (N_8433,N_7172,N_6889);
and U8434 (N_8434,N_7134,N_6743);
nor U8435 (N_8435,N_5973,N_5296);
nand U8436 (N_8436,N_5360,N_6273);
xor U8437 (N_8437,N_5370,N_6045);
or U8438 (N_8438,N_5025,N_7249);
nand U8439 (N_8439,N_5881,N_5126);
nand U8440 (N_8440,N_6195,N_6839);
xor U8441 (N_8441,N_5643,N_6684);
xnor U8442 (N_8442,N_7496,N_7170);
or U8443 (N_8443,N_5352,N_6298);
nor U8444 (N_8444,N_7412,N_5021);
and U8445 (N_8445,N_7007,N_5962);
or U8446 (N_8446,N_5638,N_7103);
or U8447 (N_8447,N_6147,N_7092);
and U8448 (N_8448,N_5942,N_5664);
nand U8449 (N_8449,N_5503,N_5197);
xor U8450 (N_8450,N_5790,N_6366);
nand U8451 (N_8451,N_7214,N_6776);
xnor U8452 (N_8452,N_5680,N_5910);
or U8453 (N_8453,N_5344,N_6553);
nor U8454 (N_8454,N_5603,N_6253);
nor U8455 (N_8455,N_6391,N_6467);
nand U8456 (N_8456,N_5209,N_6248);
and U8457 (N_8457,N_7025,N_6375);
nor U8458 (N_8458,N_5012,N_5699);
and U8459 (N_8459,N_5467,N_5838);
or U8460 (N_8460,N_5376,N_6137);
nand U8461 (N_8461,N_5049,N_5206);
nor U8462 (N_8462,N_6570,N_5711);
or U8463 (N_8463,N_6174,N_5808);
nor U8464 (N_8464,N_7392,N_5145);
nand U8465 (N_8465,N_6436,N_5357);
xnor U8466 (N_8466,N_6360,N_5166);
or U8467 (N_8467,N_5163,N_6647);
or U8468 (N_8468,N_6832,N_5473);
nand U8469 (N_8469,N_5755,N_6034);
and U8470 (N_8470,N_6660,N_5203);
xor U8471 (N_8471,N_5117,N_5602);
xnor U8472 (N_8472,N_5599,N_5186);
or U8473 (N_8473,N_6969,N_5019);
or U8474 (N_8474,N_5786,N_5051);
nand U8475 (N_8475,N_6808,N_5521);
and U8476 (N_8476,N_5434,N_6267);
nor U8477 (N_8477,N_7099,N_6695);
or U8478 (N_8478,N_6116,N_6576);
xnor U8479 (N_8479,N_6590,N_6624);
nor U8480 (N_8480,N_5930,N_5901);
nand U8481 (N_8481,N_5321,N_7294);
nor U8482 (N_8482,N_6365,N_5827);
nor U8483 (N_8483,N_6269,N_6234);
or U8484 (N_8484,N_6237,N_6970);
nand U8485 (N_8485,N_5445,N_5356);
and U8486 (N_8486,N_5771,N_5459);
nor U8487 (N_8487,N_5721,N_6214);
nor U8488 (N_8488,N_7386,N_7354);
or U8489 (N_8489,N_5216,N_6565);
nor U8490 (N_8490,N_5412,N_6449);
nor U8491 (N_8491,N_5510,N_7317);
nor U8492 (N_8492,N_5212,N_6486);
and U8493 (N_8493,N_6762,N_5865);
and U8494 (N_8494,N_5064,N_5204);
xnor U8495 (N_8495,N_6173,N_7000);
and U8496 (N_8496,N_6612,N_5104);
or U8497 (N_8497,N_6526,N_7275);
and U8498 (N_8498,N_6960,N_7396);
or U8499 (N_8499,N_7036,N_6311);
and U8500 (N_8500,N_6744,N_5993);
nand U8501 (N_8501,N_7181,N_6249);
xnor U8502 (N_8502,N_6014,N_6497);
xnor U8503 (N_8503,N_5646,N_7105);
and U8504 (N_8504,N_5798,N_6415);
or U8505 (N_8505,N_5651,N_5343);
or U8506 (N_8506,N_5703,N_6417);
or U8507 (N_8507,N_5176,N_5239);
or U8508 (N_8508,N_5784,N_5214);
xnor U8509 (N_8509,N_6432,N_7401);
and U8510 (N_8510,N_6351,N_5948);
and U8511 (N_8511,N_5606,N_6959);
and U8512 (N_8512,N_7010,N_5989);
xor U8513 (N_8513,N_6328,N_6753);
xnor U8514 (N_8514,N_7212,N_6478);
nor U8515 (N_8515,N_5876,N_5690);
xnor U8516 (N_8516,N_5275,N_5256);
and U8517 (N_8517,N_5804,N_5897);
nor U8518 (N_8518,N_7436,N_6632);
or U8519 (N_8519,N_7261,N_6482);
xnor U8520 (N_8520,N_6729,N_6077);
nor U8521 (N_8521,N_6208,N_7409);
or U8522 (N_8522,N_7398,N_6048);
nand U8523 (N_8523,N_5732,N_5877);
and U8524 (N_8524,N_6016,N_5596);
and U8525 (N_8525,N_7466,N_7439);
or U8526 (N_8526,N_6412,N_5559);
or U8527 (N_8527,N_7228,N_5886);
or U8528 (N_8528,N_7206,N_5302);
and U8529 (N_8529,N_5925,N_6913);
nor U8530 (N_8530,N_5893,N_5298);
and U8531 (N_8531,N_6218,N_7031);
xor U8532 (N_8532,N_5072,N_5508);
or U8533 (N_8533,N_5250,N_5231);
and U8534 (N_8534,N_5920,N_7136);
and U8535 (N_8535,N_5079,N_5826);
nand U8536 (N_8536,N_5797,N_6156);
xor U8537 (N_8537,N_6004,N_6848);
nand U8538 (N_8538,N_5853,N_6113);
nor U8539 (N_8539,N_6644,N_5408);
nand U8540 (N_8540,N_6965,N_5430);
or U8541 (N_8541,N_7018,N_5496);
nor U8542 (N_8542,N_5688,N_5551);
xor U8543 (N_8543,N_5099,N_7197);
nand U8544 (N_8544,N_7145,N_5111);
xnor U8545 (N_8545,N_5300,N_5825);
xnor U8546 (N_8546,N_5446,N_7210);
xor U8547 (N_8547,N_7118,N_5753);
or U8548 (N_8548,N_7213,N_5465);
nand U8549 (N_8549,N_7403,N_6676);
and U8550 (N_8550,N_5172,N_6823);
and U8551 (N_8551,N_5105,N_7110);
nor U8552 (N_8552,N_7097,N_7266);
nor U8553 (N_8553,N_7115,N_6096);
and U8554 (N_8554,N_7414,N_6915);
nand U8555 (N_8555,N_6282,N_5280);
nor U8556 (N_8556,N_6926,N_5109);
and U8557 (N_8557,N_7200,N_5938);
and U8558 (N_8558,N_7337,N_5195);
or U8559 (N_8559,N_7393,N_5932);
nor U8560 (N_8560,N_7450,N_5954);
nand U8561 (N_8561,N_5704,N_6361);
nor U8562 (N_8562,N_7478,N_5375);
xor U8563 (N_8563,N_5792,N_5444);
xnor U8564 (N_8564,N_5498,N_5607);
and U8565 (N_8565,N_5415,N_7395);
nor U8566 (N_8566,N_7001,N_6667);
nor U8567 (N_8567,N_5751,N_6775);
and U8568 (N_8568,N_6623,N_6213);
and U8569 (N_8569,N_6962,N_6543);
nor U8570 (N_8570,N_7292,N_5057);
nand U8571 (N_8571,N_6584,N_6772);
and U8572 (N_8572,N_6038,N_6607);
or U8573 (N_8573,N_6830,N_6091);
xor U8574 (N_8574,N_6521,N_6390);
xor U8575 (N_8575,N_5539,N_6562);
or U8576 (N_8576,N_6071,N_7244);
and U8577 (N_8577,N_6537,N_7157);
and U8578 (N_8578,N_7368,N_6098);
or U8579 (N_8579,N_6289,N_7168);
xor U8580 (N_8580,N_5235,N_6703);
xnor U8581 (N_8581,N_7006,N_5611);
or U8582 (N_8582,N_6828,N_6470);
and U8583 (N_8583,N_6272,N_5170);
and U8584 (N_8584,N_5477,N_6698);
or U8585 (N_8585,N_7043,N_6872);
nand U8586 (N_8586,N_7201,N_7174);
and U8587 (N_8587,N_6898,N_5776);
or U8588 (N_8588,N_6260,N_5378);
xnor U8589 (N_8589,N_5091,N_6441);
or U8590 (N_8590,N_6095,N_7248);
xor U8591 (N_8591,N_5455,N_7163);
xor U8592 (N_8592,N_6705,N_5803);
xor U8593 (N_8593,N_5578,N_5682);
and U8594 (N_8594,N_7465,N_6079);
xor U8595 (N_8595,N_7026,N_7456);
xnor U8596 (N_8596,N_6545,N_6087);
nand U8597 (N_8597,N_7216,N_7328);
xnor U8598 (N_8598,N_7457,N_7339);
and U8599 (N_8599,N_6863,N_6254);
nand U8600 (N_8600,N_6936,N_6666);
xor U8601 (N_8601,N_5243,N_6127);
or U8602 (N_8602,N_6027,N_5966);
xnor U8603 (N_8603,N_6508,N_6678);
xor U8604 (N_8604,N_6285,N_5227);
or U8605 (N_8605,N_5743,N_6787);
xnor U8606 (N_8606,N_7058,N_5254);
nand U8607 (N_8607,N_7427,N_6152);
and U8608 (N_8608,N_5967,N_6063);
xnor U8609 (N_8609,N_7253,N_6826);
nand U8610 (N_8610,N_7276,N_6835);
xor U8611 (N_8611,N_7449,N_6501);
or U8612 (N_8612,N_6012,N_5395);
nor U8613 (N_8613,N_5947,N_5980);
nor U8614 (N_8614,N_6411,N_6804);
and U8615 (N_8615,N_6720,N_5013);
xor U8616 (N_8616,N_7152,N_5907);
and U8617 (N_8617,N_5046,N_5489);
nand U8618 (N_8618,N_5146,N_5403);
nor U8619 (N_8619,N_6755,N_6362);
and U8620 (N_8620,N_6906,N_5187);
nand U8621 (N_8621,N_7373,N_5964);
or U8622 (N_8622,N_5222,N_5591);
or U8623 (N_8623,N_7433,N_6398);
xor U8624 (N_8624,N_7011,N_6499);
xnor U8625 (N_8625,N_7246,N_6209);
xnor U8626 (N_8626,N_5887,N_5394);
and U8627 (N_8627,N_5307,N_5406);
xor U8628 (N_8628,N_6895,N_5391);
xor U8629 (N_8629,N_6225,N_5120);
or U8630 (N_8630,N_5773,N_5940);
xor U8631 (N_8631,N_5355,N_5933);
and U8632 (N_8632,N_5644,N_5585);
xnor U8633 (N_8633,N_7322,N_7225);
and U8634 (N_8634,N_5618,N_5291);
or U8635 (N_8635,N_6907,N_5029);
nand U8636 (N_8636,N_6446,N_6178);
and U8637 (N_8637,N_7390,N_5440);
or U8638 (N_8638,N_5078,N_5081);
nor U8639 (N_8639,N_7016,N_5401);
or U8640 (N_8640,N_6626,N_6438);
or U8641 (N_8641,N_5739,N_5586);
nor U8642 (N_8642,N_5678,N_6245);
nor U8643 (N_8643,N_5264,N_6485);
nand U8644 (N_8644,N_5812,N_5451);
nand U8645 (N_8645,N_6297,N_6892);
nor U8646 (N_8646,N_6704,N_7151);
and U8647 (N_8647,N_5554,N_5653);
xnor U8648 (N_8648,N_5687,N_7123);
and U8649 (N_8649,N_5327,N_5436);
nor U8650 (N_8650,N_7323,N_6669);
and U8651 (N_8651,N_6927,N_5023);
and U8652 (N_8652,N_7250,N_7352);
nand U8653 (N_8653,N_7305,N_6172);
nor U8654 (N_8654,N_5709,N_5671);
xor U8655 (N_8655,N_6859,N_5463);
xor U8656 (N_8656,N_5226,N_7484);
nand U8657 (N_8657,N_6674,N_6312);
xor U8658 (N_8658,N_6371,N_6752);
nand U8659 (N_8659,N_6838,N_5652);
xor U8660 (N_8660,N_5481,N_5205);
or U8661 (N_8661,N_6514,N_6974);
nand U8662 (N_8662,N_7442,N_5828);
and U8663 (N_8663,N_6976,N_5956);
nand U8664 (N_8664,N_6033,N_7087);
xnor U8665 (N_8665,N_5379,N_5635);
and U8666 (N_8666,N_7009,N_7059);
nand U8667 (N_8667,N_6515,N_7348);
nor U8668 (N_8668,N_5650,N_6191);
nand U8669 (N_8669,N_5122,N_5270);
or U8670 (N_8670,N_7263,N_6196);
nand U8671 (N_8671,N_5359,N_6425);
or U8672 (N_8672,N_6133,N_5615);
and U8673 (N_8673,N_5121,N_6342);
xnor U8674 (N_8674,N_7326,N_6424);
or U8675 (N_8675,N_5303,N_6413);
and U8676 (N_8676,N_6873,N_7402);
nand U8677 (N_8677,N_7173,N_6558);
nor U8678 (N_8678,N_5849,N_5725);
nor U8679 (N_8679,N_6939,N_5024);
nand U8680 (N_8680,N_6887,N_5557);
or U8681 (N_8681,N_5846,N_6363);
nand U8682 (N_8682,N_5538,N_5335);
nand U8683 (N_8683,N_6554,N_5087);
or U8684 (N_8684,N_6982,N_6495);
and U8685 (N_8685,N_5177,N_5136);
or U8686 (N_8686,N_5411,N_7125);
or U8687 (N_8687,N_5608,N_6340);
or U8688 (N_8688,N_5957,N_5906);
or U8689 (N_8689,N_6905,N_7109);
xor U8690 (N_8690,N_7051,N_6313);
or U8691 (N_8691,N_5657,N_6901);
xnor U8692 (N_8692,N_6404,N_6816);
nand U8693 (N_8693,N_6792,N_5822);
or U8694 (N_8694,N_5820,N_6617);
nor U8695 (N_8695,N_6988,N_6968);
nand U8696 (N_8696,N_6603,N_5366);
nand U8697 (N_8697,N_6383,N_6557);
nor U8698 (N_8698,N_5626,N_5011);
or U8699 (N_8699,N_6922,N_7111);
and U8700 (N_8700,N_6032,N_5409);
nand U8701 (N_8701,N_6278,N_6946);
xnor U8702 (N_8702,N_6765,N_5110);
or U8703 (N_8703,N_7066,N_7028);
xnor U8704 (N_8704,N_6235,N_6115);
nand U8705 (N_8705,N_6707,N_5306);
and U8706 (N_8706,N_7241,N_5592);
and U8707 (N_8707,N_6658,N_5959);
or U8708 (N_8708,N_5900,N_5661);
nor U8709 (N_8709,N_5689,N_5536);
nor U8710 (N_8710,N_5627,N_7381);
and U8711 (N_8711,N_6007,N_5780);
nor U8712 (N_8712,N_7321,N_5891);
or U8713 (N_8713,N_7078,N_6567);
or U8714 (N_8714,N_6112,N_7489);
or U8715 (N_8715,N_6076,N_5014);
and U8716 (N_8716,N_5756,N_6692);
xnor U8717 (N_8717,N_5318,N_5598);
xnor U8718 (N_8718,N_7467,N_6878);
and U8719 (N_8719,N_6771,N_5208);
nor U8720 (N_8720,N_6193,N_5637);
or U8721 (N_8721,N_5069,N_5889);
nor U8722 (N_8722,N_7156,N_5625);
and U8723 (N_8723,N_6821,N_7050);
xor U8724 (N_8724,N_7472,N_6337);
or U8725 (N_8725,N_5283,N_5040);
nor U8726 (N_8726,N_5795,N_5497);
xnor U8727 (N_8727,N_6504,N_7104);
nor U8728 (N_8728,N_6656,N_5695);
or U8729 (N_8729,N_6466,N_6681);
and U8730 (N_8730,N_6690,N_7065);
nor U8731 (N_8731,N_6005,N_7269);
xnor U8732 (N_8732,N_6691,N_5044);
nand U8733 (N_8733,N_5567,N_6610);
or U8734 (N_8734,N_7330,N_5903);
and U8735 (N_8735,N_5223,N_6268);
xnor U8736 (N_8736,N_7308,N_5981);
nor U8737 (N_8737,N_5039,N_6000);
xor U8738 (N_8738,N_5879,N_5929);
xor U8739 (N_8739,N_7035,N_7114);
xnor U8740 (N_8740,N_6123,N_7474);
or U8741 (N_8741,N_5986,N_5636);
xnor U8742 (N_8742,N_5896,N_5482);
or U8743 (N_8743,N_6481,N_7098);
or U8744 (N_8744,N_5056,N_6528);
or U8745 (N_8745,N_5350,N_5532);
nand U8746 (N_8746,N_6279,N_5960);
nand U8747 (N_8747,N_5422,N_5054);
xnor U8748 (N_8748,N_6726,N_6713);
nand U8749 (N_8749,N_7338,N_5791);
nand U8750 (N_8750,N_7030,N_6107);
and U8751 (N_8751,N_6494,N_6219);
or U8752 (N_8752,N_5721,N_5932);
xor U8753 (N_8753,N_5172,N_7382);
or U8754 (N_8754,N_5042,N_6843);
xor U8755 (N_8755,N_7146,N_7187);
and U8756 (N_8756,N_7333,N_5049);
xor U8757 (N_8757,N_5990,N_5976);
nand U8758 (N_8758,N_7443,N_6037);
and U8759 (N_8759,N_5215,N_7237);
and U8760 (N_8760,N_6769,N_7022);
nor U8761 (N_8761,N_6795,N_6327);
nand U8762 (N_8762,N_6231,N_6632);
nor U8763 (N_8763,N_6309,N_5176);
nand U8764 (N_8764,N_5726,N_6215);
or U8765 (N_8765,N_5783,N_5470);
or U8766 (N_8766,N_7285,N_5559);
nand U8767 (N_8767,N_6673,N_7200);
nor U8768 (N_8768,N_5430,N_6769);
and U8769 (N_8769,N_6280,N_6435);
xor U8770 (N_8770,N_5484,N_6201);
nand U8771 (N_8771,N_6267,N_5613);
xor U8772 (N_8772,N_5745,N_7014);
nor U8773 (N_8773,N_7159,N_6766);
and U8774 (N_8774,N_5716,N_6382);
nor U8775 (N_8775,N_6836,N_5281);
nand U8776 (N_8776,N_5712,N_6550);
or U8777 (N_8777,N_7426,N_6819);
xor U8778 (N_8778,N_6392,N_6140);
or U8779 (N_8779,N_6854,N_6531);
xor U8780 (N_8780,N_6763,N_6747);
xnor U8781 (N_8781,N_5004,N_6769);
nor U8782 (N_8782,N_7198,N_6653);
and U8783 (N_8783,N_7261,N_5314);
nor U8784 (N_8784,N_6671,N_5232);
nor U8785 (N_8785,N_6175,N_5737);
nand U8786 (N_8786,N_7235,N_5731);
nand U8787 (N_8787,N_5276,N_7333);
nand U8788 (N_8788,N_6224,N_5014);
and U8789 (N_8789,N_6342,N_6214);
and U8790 (N_8790,N_6185,N_6564);
and U8791 (N_8791,N_7274,N_6188);
nor U8792 (N_8792,N_7145,N_5755);
and U8793 (N_8793,N_5879,N_5990);
and U8794 (N_8794,N_5278,N_6237);
nand U8795 (N_8795,N_6586,N_6833);
nor U8796 (N_8796,N_6735,N_5227);
nand U8797 (N_8797,N_6942,N_5896);
or U8798 (N_8798,N_5703,N_6171);
and U8799 (N_8799,N_5900,N_6344);
xnor U8800 (N_8800,N_5813,N_7111);
and U8801 (N_8801,N_5069,N_5223);
nor U8802 (N_8802,N_7347,N_6152);
and U8803 (N_8803,N_5901,N_6995);
xor U8804 (N_8804,N_7487,N_5079);
and U8805 (N_8805,N_7051,N_5998);
nand U8806 (N_8806,N_6645,N_6881);
nor U8807 (N_8807,N_7106,N_5162);
nand U8808 (N_8808,N_7004,N_6591);
nand U8809 (N_8809,N_5249,N_6966);
nand U8810 (N_8810,N_5942,N_7240);
or U8811 (N_8811,N_5445,N_5848);
nor U8812 (N_8812,N_6304,N_7202);
and U8813 (N_8813,N_7005,N_6866);
and U8814 (N_8814,N_6412,N_5552);
nor U8815 (N_8815,N_6177,N_5938);
xnor U8816 (N_8816,N_5051,N_6527);
nor U8817 (N_8817,N_6877,N_6822);
nand U8818 (N_8818,N_7123,N_6157);
nand U8819 (N_8819,N_6103,N_6340);
or U8820 (N_8820,N_5407,N_7307);
nand U8821 (N_8821,N_6420,N_7153);
xor U8822 (N_8822,N_5979,N_6012);
nand U8823 (N_8823,N_7327,N_7272);
nor U8824 (N_8824,N_7279,N_6257);
or U8825 (N_8825,N_5081,N_7361);
or U8826 (N_8826,N_5129,N_7017);
or U8827 (N_8827,N_7287,N_5423);
and U8828 (N_8828,N_5160,N_6052);
and U8829 (N_8829,N_7055,N_5477);
or U8830 (N_8830,N_5423,N_7048);
nand U8831 (N_8831,N_7213,N_6392);
xnor U8832 (N_8832,N_6666,N_6403);
and U8833 (N_8833,N_5074,N_5016);
xnor U8834 (N_8834,N_5756,N_7002);
or U8835 (N_8835,N_7208,N_6452);
nor U8836 (N_8836,N_6307,N_6339);
or U8837 (N_8837,N_5366,N_6669);
xnor U8838 (N_8838,N_5694,N_5619);
and U8839 (N_8839,N_6461,N_6611);
or U8840 (N_8840,N_5694,N_5436);
or U8841 (N_8841,N_7458,N_5611);
or U8842 (N_8842,N_5794,N_6653);
xnor U8843 (N_8843,N_5194,N_5432);
or U8844 (N_8844,N_7350,N_5405);
nor U8845 (N_8845,N_7398,N_6882);
or U8846 (N_8846,N_6959,N_7167);
xnor U8847 (N_8847,N_6693,N_6301);
or U8848 (N_8848,N_5316,N_5877);
xor U8849 (N_8849,N_7333,N_7302);
nand U8850 (N_8850,N_5954,N_6551);
and U8851 (N_8851,N_5689,N_5187);
xnor U8852 (N_8852,N_7128,N_7124);
and U8853 (N_8853,N_6323,N_6370);
xor U8854 (N_8854,N_6062,N_5162);
nor U8855 (N_8855,N_5238,N_5865);
or U8856 (N_8856,N_5144,N_6322);
and U8857 (N_8857,N_7079,N_5716);
nor U8858 (N_8858,N_6924,N_5339);
or U8859 (N_8859,N_5526,N_5930);
nand U8860 (N_8860,N_5646,N_6551);
xor U8861 (N_8861,N_5146,N_5353);
and U8862 (N_8862,N_5727,N_7465);
or U8863 (N_8863,N_7069,N_7190);
xor U8864 (N_8864,N_7302,N_6585);
xor U8865 (N_8865,N_6186,N_6249);
nand U8866 (N_8866,N_5365,N_6474);
xor U8867 (N_8867,N_5579,N_6757);
nor U8868 (N_8868,N_5032,N_5158);
nor U8869 (N_8869,N_6606,N_7100);
nor U8870 (N_8870,N_7193,N_6882);
or U8871 (N_8871,N_5636,N_5386);
and U8872 (N_8872,N_6645,N_6232);
or U8873 (N_8873,N_7207,N_6339);
nand U8874 (N_8874,N_6467,N_5486);
and U8875 (N_8875,N_7289,N_5795);
nand U8876 (N_8876,N_5919,N_5128);
nand U8877 (N_8877,N_5388,N_6824);
nor U8878 (N_8878,N_7233,N_5687);
xnor U8879 (N_8879,N_7457,N_6947);
and U8880 (N_8880,N_6961,N_6725);
nor U8881 (N_8881,N_6493,N_7254);
and U8882 (N_8882,N_6913,N_5759);
and U8883 (N_8883,N_5456,N_6507);
xnor U8884 (N_8884,N_6059,N_6750);
or U8885 (N_8885,N_6561,N_5073);
nor U8886 (N_8886,N_7047,N_5663);
or U8887 (N_8887,N_6492,N_6248);
and U8888 (N_8888,N_6885,N_5236);
xnor U8889 (N_8889,N_6571,N_5432);
xnor U8890 (N_8890,N_5907,N_5932);
nor U8891 (N_8891,N_5637,N_6896);
xnor U8892 (N_8892,N_6685,N_7402);
and U8893 (N_8893,N_7315,N_6716);
nand U8894 (N_8894,N_5822,N_5750);
nor U8895 (N_8895,N_5084,N_6465);
nor U8896 (N_8896,N_5847,N_6511);
and U8897 (N_8897,N_6975,N_5495);
nand U8898 (N_8898,N_5699,N_6899);
nand U8899 (N_8899,N_5433,N_6709);
xnor U8900 (N_8900,N_6359,N_5084);
nand U8901 (N_8901,N_5111,N_7158);
nor U8902 (N_8902,N_6454,N_7366);
nor U8903 (N_8903,N_5867,N_5822);
nand U8904 (N_8904,N_5439,N_5084);
xor U8905 (N_8905,N_5669,N_5802);
and U8906 (N_8906,N_5799,N_5223);
xor U8907 (N_8907,N_7042,N_6444);
nand U8908 (N_8908,N_6535,N_6853);
or U8909 (N_8909,N_5516,N_5186);
nor U8910 (N_8910,N_7094,N_5529);
nand U8911 (N_8911,N_5256,N_5338);
nand U8912 (N_8912,N_5902,N_5883);
or U8913 (N_8913,N_5483,N_5977);
nor U8914 (N_8914,N_6535,N_5980);
and U8915 (N_8915,N_5895,N_5282);
and U8916 (N_8916,N_5308,N_5909);
nor U8917 (N_8917,N_5146,N_7020);
or U8918 (N_8918,N_5834,N_6898);
xnor U8919 (N_8919,N_7075,N_6156);
nand U8920 (N_8920,N_6245,N_5350);
and U8921 (N_8921,N_6025,N_6318);
and U8922 (N_8922,N_6288,N_7118);
nor U8923 (N_8923,N_6668,N_5077);
nand U8924 (N_8924,N_6150,N_5482);
and U8925 (N_8925,N_5436,N_5077);
xnor U8926 (N_8926,N_6252,N_7282);
nor U8927 (N_8927,N_5110,N_5550);
and U8928 (N_8928,N_7143,N_5004);
or U8929 (N_8929,N_5879,N_7241);
xor U8930 (N_8930,N_5679,N_5695);
nand U8931 (N_8931,N_5821,N_5990);
and U8932 (N_8932,N_5627,N_6203);
xnor U8933 (N_8933,N_6126,N_7477);
nand U8934 (N_8934,N_6057,N_5714);
xor U8935 (N_8935,N_5482,N_6483);
and U8936 (N_8936,N_5187,N_5557);
or U8937 (N_8937,N_5608,N_6325);
or U8938 (N_8938,N_5684,N_6954);
or U8939 (N_8939,N_6083,N_7278);
xnor U8940 (N_8940,N_5402,N_5859);
nor U8941 (N_8941,N_5721,N_5117);
or U8942 (N_8942,N_5036,N_6246);
xor U8943 (N_8943,N_6341,N_6061);
nand U8944 (N_8944,N_5265,N_6004);
and U8945 (N_8945,N_7098,N_6287);
nor U8946 (N_8946,N_6522,N_6194);
nor U8947 (N_8947,N_5955,N_6666);
nor U8948 (N_8948,N_6567,N_6707);
nor U8949 (N_8949,N_5963,N_5017);
nand U8950 (N_8950,N_6957,N_6622);
or U8951 (N_8951,N_6880,N_7004);
and U8952 (N_8952,N_6333,N_6968);
nor U8953 (N_8953,N_6200,N_5975);
xnor U8954 (N_8954,N_5614,N_5528);
and U8955 (N_8955,N_7136,N_6561);
or U8956 (N_8956,N_7135,N_5600);
nand U8957 (N_8957,N_6713,N_5173);
nand U8958 (N_8958,N_5386,N_5874);
xor U8959 (N_8959,N_6292,N_6406);
xnor U8960 (N_8960,N_5356,N_6476);
and U8961 (N_8961,N_5686,N_7479);
and U8962 (N_8962,N_7221,N_5480);
xnor U8963 (N_8963,N_5355,N_7092);
nor U8964 (N_8964,N_7349,N_7314);
nand U8965 (N_8965,N_6716,N_7497);
xnor U8966 (N_8966,N_5699,N_5161);
xnor U8967 (N_8967,N_5562,N_5872);
xor U8968 (N_8968,N_7413,N_7231);
xnor U8969 (N_8969,N_5648,N_6913);
xor U8970 (N_8970,N_6012,N_6032);
nand U8971 (N_8971,N_7010,N_5819);
or U8972 (N_8972,N_6543,N_6714);
or U8973 (N_8973,N_5933,N_6581);
nand U8974 (N_8974,N_6350,N_5397);
xor U8975 (N_8975,N_6084,N_6325);
xor U8976 (N_8976,N_6050,N_7362);
nand U8977 (N_8977,N_5054,N_5123);
nand U8978 (N_8978,N_6063,N_7035);
nor U8979 (N_8979,N_5364,N_5009);
and U8980 (N_8980,N_6258,N_6673);
nor U8981 (N_8981,N_6816,N_6208);
nor U8982 (N_8982,N_5450,N_6585);
or U8983 (N_8983,N_5524,N_6880);
or U8984 (N_8984,N_6561,N_6613);
nor U8985 (N_8985,N_6595,N_6856);
xnor U8986 (N_8986,N_6554,N_7416);
nand U8987 (N_8987,N_5817,N_5499);
nor U8988 (N_8988,N_5249,N_5576);
and U8989 (N_8989,N_5629,N_5519);
xor U8990 (N_8990,N_6625,N_7094);
or U8991 (N_8991,N_7049,N_6262);
nand U8992 (N_8992,N_6964,N_6624);
nand U8993 (N_8993,N_7052,N_7247);
nor U8994 (N_8994,N_7366,N_7243);
or U8995 (N_8995,N_6740,N_6974);
nor U8996 (N_8996,N_6498,N_5022);
xor U8997 (N_8997,N_7476,N_6775);
or U8998 (N_8998,N_5940,N_6792);
nor U8999 (N_8999,N_5166,N_5319);
nor U9000 (N_9000,N_5895,N_5644);
or U9001 (N_9001,N_5998,N_6349);
and U9002 (N_9002,N_5641,N_6859);
or U9003 (N_9003,N_7311,N_6350);
xor U9004 (N_9004,N_5302,N_5124);
and U9005 (N_9005,N_7128,N_7456);
xor U9006 (N_9006,N_5166,N_6086);
xnor U9007 (N_9007,N_7463,N_6282);
or U9008 (N_9008,N_7046,N_6945);
and U9009 (N_9009,N_5002,N_6488);
nor U9010 (N_9010,N_5290,N_6227);
and U9011 (N_9011,N_5205,N_5722);
nor U9012 (N_9012,N_5250,N_6006);
and U9013 (N_9013,N_6633,N_7061);
nand U9014 (N_9014,N_7091,N_6741);
and U9015 (N_9015,N_5039,N_7113);
nand U9016 (N_9016,N_5193,N_5161);
nor U9017 (N_9017,N_7258,N_5909);
nor U9018 (N_9018,N_7238,N_6831);
nor U9019 (N_9019,N_6576,N_7398);
nand U9020 (N_9020,N_7085,N_5402);
and U9021 (N_9021,N_6702,N_5771);
nand U9022 (N_9022,N_7115,N_6122);
nand U9023 (N_9023,N_7054,N_6585);
and U9024 (N_9024,N_5137,N_6826);
xor U9025 (N_9025,N_6640,N_5118);
nor U9026 (N_9026,N_5085,N_5953);
xor U9027 (N_9027,N_6118,N_5332);
nand U9028 (N_9028,N_6013,N_6843);
and U9029 (N_9029,N_6318,N_7188);
or U9030 (N_9030,N_6310,N_7178);
xor U9031 (N_9031,N_6038,N_6463);
xnor U9032 (N_9032,N_7467,N_6174);
nand U9033 (N_9033,N_5926,N_6178);
and U9034 (N_9034,N_6013,N_5914);
and U9035 (N_9035,N_6265,N_6719);
xor U9036 (N_9036,N_7478,N_7149);
or U9037 (N_9037,N_7073,N_6204);
and U9038 (N_9038,N_6485,N_6748);
or U9039 (N_9039,N_6194,N_7232);
or U9040 (N_9040,N_6576,N_5181);
nand U9041 (N_9041,N_5527,N_5399);
nor U9042 (N_9042,N_7294,N_5975);
and U9043 (N_9043,N_5539,N_6751);
and U9044 (N_9044,N_6065,N_7183);
xnor U9045 (N_9045,N_5695,N_5037);
and U9046 (N_9046,N_5694,N_6066);
nand U9047 (N_9047,N_5002,N_6282);
xor U9048 (N_9048,N_7367,N_5595);
nand U9049 (N_9049,N_5894,N_5248);
xnor U9050 (N_9050,N_5891,N_6582);
xor U9051 (N_9051,N_6045,N_5977);
nor U9052 (N_9052,N_5616,N_7212);
xnor U9053 (N_9053,N_7135,N_6028);
nand U9054 (N_9054,N_6559,N_5074);
or U9055 (N_9055,N_6949,N_5144);
nand U9056 (N_9056,N_6175,N_5587);
nor U9057 (N_9057,N_5909,N_6897);
or U9058 (N_9058,N_6026,N_6817);
nor U9059 (N_9059,N_6277,N_5484);
xor U9060 (N_9060,N_7392,N_5213);
nor U9061 (N_9061,N_7009,N_5764);
xor U9062 (N_9062,N_5975,N_6091);
nor U9063 (N_9063,N_5038,N_5787);
nor U9064 (N_9064,N_5970,N_5638);
nor U9065 (N_9065,N_5154,N_5800);
xor U9066 (N_9066,N_5753,N_7288);
and U9067 (N_9067,N_7436,N_6040);
nor U9068 (N_9068,N_5557,N_6340);
nor U9069 (N_9069,N_6116,N_6889);
xnor U9070 (N_9070,N_6951,N_6867);
and U9071 (N_9071,N_5950,N_5423);
and U9072 (N_9072,N_5658,N_5406);
or U9073 (N_9073,N_5206,N_5807);
or U9074 (N_9074,N_7048,N_5411);
nor U9075 (N_9075,N_5356,N_5076);
nand U9076 (N_9076,N_6727,N_5201);
or U9077 (N_9077,N_7313,N_7069);
nand U9078 (N_9078,N_6974,N_7162);
or U9079 (N_9079,N_5547,N_5000);
and U9080 (N_9080,N_6167,N_6007);
nor U9081 (N_9081,N_7169,N_5817);
xor U9082 (N_9082,N_6029,N_6975);
nand U9083 (N_9083,N_6573,N_5360);
and U9084 (N_9084,N_6133,N_7094);
or U9085 (N_9085,N_7005,N_5184);
nor U9086 (N_9086,N_5358,N_5141);
nor U9087 (N_9087,N_5961,N_6137);
nand U9088 (N_9088,N_6556,N_6585);
nor U9089 (N_9089,N_6073,N_6413);
nand U9090 (N_9090,N_5031,N_5033);
or U9091 (N_9091,N_6108,N_5571);
nand U9092 (N_9092,N_7261,N_5707);
nand U9093 (N_9093,N_6659,N_5596);
or U9094 (N_9094,N_7472,N_6386);
nor U9095 (N_9095,N_6786,N_6141);
xnor U9096 (N_9096,N_6238,N_5047);
xor U9097 (N_9097,N_6575,N_7445);
nand U9098 (N_9098,N_5230,N_6694);
xor U9099 (N_9099,N_6188,N_5163);
xnor U9100 (N_9100,N_5440,N_6585);
nor U9101 (N_9101,N_7021,N_5717);
or U9102 (N_9102,N_5373,N_5916);
or U9103 (N_9103,N_5708,N_6148);
xor U9104 (N_9104,N_5742,N_6333);
nor U9105 (N_9105,N_6398,N_5731);
xor U9106 (N_9106,N_7250,N_5738);
nor U9107 (N_9107,N_6963,N_6575);
or U9108 (N_9108,N_6737,N_6093);
and U9109 (N_9109,N_5643,N_5084);
or U9110 (N_9110,N_6738,N_6185);
nor U9111 (N_9111,N_6209,N_7080);
nand U9112 (N_9112,N_5314,N_5524);
and U9113 (N_9113,N_7496,N_5762);
or U9114 (N_9114,N_6663,N_6160);
xnor U9115 (N_9115,N_5888,N_7256);
nor U9116 (N_9116,N_7157,N_5385);
nand U9117 (N_9117,N_5698,N_5702);
nor U9118 (N_9118,N_6002,N_5076);
nand U9119 (N_9119,N_6751,N_5581);
nor U9120 (N_9120,N_5383,N_5359);
or U9121 (N_9121,N_5635,N_5362);
nor U9122 (N_9122,N_6248,N_5256);
or U9123 (N_9123,N_5543,N_6295);
xnor U9124 (N_9124,N_5341,N_5802);
and U9125 (N_9125,N_5068,N_5039);
xor U9126 (N_9126,N_5221,N_6840);
and U9127 (N_9127,N_5284,N_7268);
xnor U9128 (N_9128,N_6751,N_7001);
and U9129 (N_9129,N_7316,N_5206);
and U9130 (N_9130,N_5642,N_7045);
or U9131 (N_9131,N_7178,N_7036);
or U9132 (N_9132,N_6319,N_5668);
nor U9133 (N_9133,N_7186,N_6602);
xnor U9134 (N_9134,N_5730,N_6825);
nor U9135 (N_9135,N_7249,N_6597);
nand U9136 (N_9136,N_5919,N_6033);
and U9137 (N_9137,N_6502,N_6427);
xor U9138 (N_9138,N_7120,N_6691);
nand U9139 (N_9139,N_5483,N_5876);
or U9140 (N_9140,N_6280,N_5732);
nand U9141 (N_9141,N_6297,N_5414);
nor U9142 (N_9142,N_6705,N_5817);
or U9143 (N_9143,N_6855,N_6193);
xor U9144 (N_9144,N_5657,N_6210);
nor U9145 (N_9145,N_7265,N_6670);
nand U9146 (N_9146,N_5326,N_6896);
nand U9147 (N_9147,N_7493,N_5886);
xnor U9148 (N_9148,N_6318,N_5852);
xor U9149 (N_9149,N_6856,N_5052);
and U9150 (N_9150,N_5210,N_6230);
nor U9151 (N_9151,N_5500,N_5263);
and U9152 (N_9152,N_5370,N_7389);
or U9153 (N_9153,N_7077,N_5176);
and U9154 (N_9154,N_7385,N_5498);
xnor U9155 (N_9155,N_6485,N_7313);
and U9156 (N_9156,N_5002,N_5331);
and U9157 (N_9157,N_6889,N_7008);
nand U9158 (N_9158,N_7472,N_6588);
or U9159 (N_9159,N_6466,N_5619);
nand U9160 (N_9160,N_5783,N_7392);
xor U9161 (N_9161,N_5892,N_5505);
or U9162 (N_9162,N_5199,N_5608);
or U9163 (N_9163,N_6907,N_7367);
or U9164 (N_9164,N_6165,N_5836);
or U9165 (N_9165,N_6515,N_6087);
nand U9166 (N_9166,N_6005,N_6785);
nand U9167 (N_9167,N_6699,N_7318);
or U9168 (N_9168,N_5716,N_5620);
or U9169 (N_9169,N_6677,N_5941);
nor U9170 (N_9170,N_6742,N_6970);
and U9171 (N_9171,N_7373,N_5871);
nor U9172 (N_9172,N_5604,N_7378);
nor U9173 (N_9173,N_5510,N_5039);
nand U9174 (N_9174,N_6853,N_5196);
xnor U9175 (N_9175,N_7486,N_7058);
xor U9176 (N_9176,N_5091,N_5441);
and U9177 (N_9177,N_5382,N_7486);
nand U9178 (N_9178,N_5265,N_6243);
and U9179 (N_9179,N_6790,N_7485);
and U9180 (N_9180,N_5983,N_5112);
and U9181 (N_9181,N_5968,N_5660);
nor U9182 (N_9182,N_5112,N_6636);
and U9183 (N_9183,N_6277,N_5322);
nand U9184 (N_9184,N_7239,N_6590);
nor U9185 (N_9185,N_5526,N_6287);
and U9186 (N_9186,N_6089,N_5100);
nand U9187 (N_9187,N_5007,N_5718);
and U9188 (N_9188,N_5124,N_5710);
xnor U9189 (N_9189,N_7373,N_5013);
or U9190 (N_9190,N_6555,N_5851);
nor U9191 (N_9191,N_6432,N_7480);
nor U9192 (N_9192,N_6487,N_5122);
nand U9193 (N_9193,N_6432,N_7109);
xor U9194 (N_9194,N_5966,N_7253);
nand U9195 (N_9195,N_7104,N_5102);
xor U9196 (N_9196,N_5640,N_5294);
nand U9197 (N_9197,N_6245,N_7347);
or U9198 (N_9198,N_7023,N_6481);
and U9199 (N_9199,N_6576,N_5614);
xor U9200 (N_9200,N_5267,N_7327);
xor U9201 (N_9201,N_5656,N_6824);
nand U9202 (N_9202,N_5407,N_7200);
xor U9203 (N_9203,N_6415,N_5405);
or U9204 (N_9204,N_7030,N_6935);
and U9205 (N_9205,N_6044,N_5924);
nand U9206 (N_9206,N_6257,N_6598);
nor U9207 (N_9207,N_6292,N_5932);
and U9208 (N_9208,N_5915,N_5074);
or U9209 (N_9209,N_6497,N_5595);
nand U9210 (N_9210,N_7303,N_5626);
nor U9211 (N_9211,N_5900,N_5224);
or U9212 (N_9212,N_6262,N_6535);
nor U9213 (N_9213,N_7136,N_7255);
or U9214 (N_9214,N_5440,N_6915);
xor U9215 (N_9215,N_5481,N_6428);
nor U9216 (N_9216,N_5311,N_5477);
nor U9217 (N_9217,N_6699,N_7002);
nand U9218 (N_9218,N_7348,N_6800);
and U9219 (N_9219,N_7389,N_5609);
nand U9220 (N_9220,N_6677,N_7180);
and U9221 (N_9221,N_7050,N_6674);
xor U9222 (N_9222,N_6464,N_5584);
or U9223 (N_9223,N_7103,N_6368);
nor U9224 (N_9224,N_6426,N_5593);
xnor U9225 (N_9225,N_7353,N_6868);
nor U9226 (N_9226,N_6408,N_7190);
and U9227 (N_9227,N_5977,N_7339);
nor U9228 (N_9228,N_5372,N_5691);
xor U9229 (N_9229,N_5451,N_5393);
xor U9230 (N_9230,N_5387,N_6278);
nor U9231 (N_9231,N_6030,N_5828);
nand U9232 (N_9232,N_5779,N_5694);
or U9233 (N_9233,N_5541,N_6157);
or U9234 (N_9234,N_5261,N_5852);
xor U9235 (N_9235,N_6740,N_5536);
or U9236 (N_9236,N_5194,N_6782);
and U9237 (N_9237,N_6283,N_6960);
nor U9238 (N_9238,N_7463,N_5544);
and U9239 (N_9239,N_5122,N_6984);
nand U9240 (N_9240,N_5461,N_5113);
nor U9241 (N_9241,N_6819,N_5470);
and U9242 (N_9242,N_5007,N_6984);
nand U9243 (N_9243,N_6645,N_6478);
or U9244 (N_9244,N_7374,N_5040);
xnor U9245 (N_9245,N_5660,N_6288);
and U9246 (N_9246,N_6931,N_6817);
or U9247 (N_9247,N_6399,N_5456);
nand U9248 (N_9248,N_7407,N_6075);
and U9249 (N_9249,N_5288,N_5040);
xor U9250 (N_9250,N_5996,N_6732);
or U9251 (N_9251,N_6397,N_5967);
nor U9252 (N_9252,N_5597,N_6958);
or U9253 (N_9253,N_6164,N_5407);
nand U9254 (N_9254,N_6766,N_6519);
or U9255 (N_9255,N_6268,N_5275);
and U9256 (N_9256,N_7000,N_5372);
or U9257 (N_9257,N_6096,N_5361);
nand U9258 (N_9258,N_5581,N_7176);
xor U9259 (N_9259,N_6856,N_7490);
and U9260 (N_9260,N_5567,N_7009);
xor U9261 (N_9261,N_5350,N_5969);
nor U9262 (N_9262,N_6654,N_7167);
nor U9263 (N_9263,N_6985,N_5946);
xor U9264 (N_9264,N_7282,N_5709);
xnor U9265 (N_9265,N_6694,N_5684);
or U9266 (N_9266,N_5564,N_5241);
or U9267 (N_9267,N_5387,N_6486);
nand U9268 (N_9268,N_5464,N_5517);
xor U9269 (N_9269,N_6230,N_5830);
and U9270 (N_9270,N_7193,N_6025);
and U9271 (N_9271,N_7035,N_5582);
nand U9272 (N_9272,N_5829,N_5132);
xor U9273 (N_9273,N_7431,N_6275);
or U9274 (N_9274,N_5262,N_6971);
nand U9275 (N_9275,N_6807,N_5881);
or U9276 (N_9276,N_5767,N_7247);
and U9277 (N_9277,N_7159,N_5740);
or U9278 (N_9278,N_6344,N_7177);
nand U9279 (N_9279,N_5862,N_6384);
and U9280 (N_9280,N_5709,N_6155);
and U9281 (N_9281,N_6854,N_7267);
nand U9282 (N_9282,N_5332,N_6514);
and U9283 (N_9283,N_7217,N_5436);
or U9284 (N_9284,N_7461,N_6253);
xor U9285 (N_9285,N_7184,N_6895);
nor U9286 (N_9286,N_7351,N_5227);
nand U9287 (N_9287,N_5923,N_5716);
nor U9288 (N_9288,N_6013,N_6388);
xnor U9289 (N_9289,N_6661,N_6372);
xor U9290 (N_9290,N_7368,N_6790);
and U9291 (N_9291,N_5233,N_6972);
and U9292 (N_9292,N_5701,N_7310);
and U9293 (N_9293,N_6618,N_5703);
or U9294 (N_9294,N_5676,N_6402);
and U9295 (N_9295,N_6451,N_5916);
or U9296 (N_9296,N_7222,N_6362);
or U9297 (N_9297,N_5326,N_6085);
nor U9298 (N_9298,N_6412,N_6332);
nand U9299 (N_9299,N_5187,N_6281);
nor U9300 (N_9300,N_5211,N_5612);
nor U9301 (N_9301,N_6885,N_6302);
nand U9302 (N_9302,N_5448,N_5432);
xor U9303 (N_9303,N_7201,N_7158);
nor U9304 (N_9304,N_5421,N_7265);
nand U9305 (N_9305,N_5091,N_6267);
and U9306 (N_9306,N_7042,N_5526);
nand U9307 (N_9307,N_5022,N_5453);
nor U9308 (N_9308,N_6659,N_6821);
and U9309 (N_9309,N_7083,N_5638);
xnor U9310 (N_9310,N_6916,N_7038);
and U9311 (N_9311,N_5960,N_6059);
nand U9312 (N_9312,N_6426,N_7398);
xnor U9313 (N_9313,N_5464,N_5584);
and U9314 (N_9314,N_6688,N_6018);
nor U9315 (N_9315,N_6016,N_5917);
xnor U9316 (N_9316,N_6739,N_5146);
and U9317 (N_9317,N_6455,N_5790);
nor U9318 (N_9318,N_5720,N_6758);
xor U9319 (N_9319,N_5768,N_6145);
or U9320 (N_9320,N_6163,N_5567);
nand U9321 (N_9321,N_7386,N_6955);
and U9322 (N_9322,N_6802,N_5345);
nor U9323 (N_9323,N_5843,N_5387);
xnor U9324 (N_9324,N_5970,N_6213);
nand U9325 (N_9325,N_6517,N_7090);
nor U9326 (N_9326,N_6590,N_7096);
and U9327 (N_9327,N_7161,N_5286);
xnor U9328 (N_9328,N_5933,N_6057);
xnor U9329 (N_9329,N_6451,N_5906);
or U9330 (N_9330,N_5910,N_5988);
and U9331 (N_9331,N_6001,N_6893);
nor U9332 (N_9332,N_7439,N_7408);
and U9333 (N_9333,N_7292,N_5528);
and U9334 (N_9334,N_6495,N_6409);
or U9335 (N_9335,N_6875,N_6402);
xnor U9336 (N_9336,N_5527,N_7035);
xor U9337 (N_9337,N_6717,N_7130);
or U9338 (N_9338,N_6338,N_5581);
nor U9339 (N_9339,N_6938,N_5490);
or U9340 (N_9340,N_6965,N_7280);
or U9341 (N_9341,N_5293,N_6203);
nand U9342 (N_9342,N_6490,N_7188);
and U9343 (N_9343,N_7112,N_6236);
xor U9344 (N_9344,N_7024,N_6502);
and U9345 (N_9345,N_5408,N_7109);
or U9346 (N_9346,N_5247,N_6312);
nand U9347 (N_9347,N_5940,N_6941);
and U9348 (N_9348,N_5510,N_5145);
or U9349 (N_9349,N_5279,N_5989);
and U9350 (N_9350,N_6065,N_6209);
nand U9351 (N_9351,N_6003,N_6792);
and U9352 (N_9352,N_7020,N_5495);
or U9353 (N_9353,N_6262,N_6837);
and U9354 (N_9354,N_6994,N_6870);
nand U9355 (N_9355,N_5271,N_5839);
or U9356 (N_9356,N_5623,N_6522);
xor U9357 (N_9357,N_5685,N_6126);
and U9358 (N_9358,N_6520,N_5718);
xor U9359 (N_9359,N_6025,N_6666);
nand U9360 (N_9360,N_6835,N_6841);
or U9361 (N_9361,N_5411,N_5749);
nand U9362 (N_9362,N_5671,N_5455);
nor U9363 (N_9363,N_6193,N_5146);
nand U9364 (N_9364,N_5540,N_5961);
and U9365 (N_9365,N_5884,N_6535);
or U9366 (N_9366,N_6749,N_5369);
or U9367 (N_9367,N_6022,N_7411);
nand U9368 (N_9368,N_6161,N_6419);
nor U9369 (N_9369,N_5570,N_6509);
and U9370 (N_9370,N_5238,N_5041);
nor U9371 (N_9371,N_6855,N_5592);
or U9372 (N_9372,N_5157,N_6709);
nor U9373 (N_9373,N_6645,N_6797);
nor U9374 (N_9374,N_5729,N_5356);
or U9375 (N_9375,N_5264,N_6082);
or U9376 (N_9376,N_7258,N_6819);
nand U9377 (N_9377,N_5740,N_6322);
and U9378 (N_9378,N_6671,N_7479);
xnor U9379 (N_9379,N_7243,N_6966);
and U9380 (N_9380,N_7108,N_6491);
nor U9381 (N_9381,N_7306,N_6434);
nor U9382 (N_9382,N_6573,N_5278);
xnor U9383 (N_9383,N_5440,N_7010);
and U9384 (N_9384,N_6002,N_6785);
nor U9385 (N_9385,N_5239,N_6210);
nand U9386 (N_9386,N_5567,N_6838);
and U9387 (N_9387,N_6959,N_6372);
and U9388 (N_9388,N_5048,N_6724);
nand U9389 (N_9389,N_6871,N_5306);
nor U9390 (N_9390,N_6032,N_5479);
xor U9391 (N_9391,N_5470,N_6180);
nor U9392 (N_9392,N_6012,N_6558);
and U9393 (N_9393,N_7067,N_6624);
and U9394 (N_9394,N_7300,N_5491);
and U9395 (N_9395,N_5399,N_6355);
and U9396 (N_9396,N_5052,N_5965);
or U9397 (N_9397,N_5401,N_7139);
or U9398 (N_9398,N_6705,N_7174);
nor U9399 (N_9399,N_7172,N_6166);
nand U9400 (N_9400,N_6414,N_7495);
or U9401 (N_9401,N_5387,N_5422);
nand U9402 (N_9402,N_6800,N_6998);
xor U9403 (N_9403,N_7420,N_5169);
and U9404 (N_9404,N_6927,N_5557);
nor U9405 (N_9405,N_5605,N_5118);
nand U9406 (N_9406,N_6925,N_6546);
nand U9407 (N_9407,N_6646,N_7282);
nor U9408 (N_9408,N_7456,N_7378);
or U9409 (N_9409,N_5257,N_5825);
or U9410 (N_9410,N_6662,N_5923);
and U9411 (N_9411,N_6435,N_6134);
xor U9412 (N_9412,N_7486,N_6179);
or U9413 (N_9413,N_5518,N_6283);
and U9414 (N_9414,N_6230,N_6792);
nand U9415 (N_9415,N_6153,N_6477);
or U9416 (N_9416,N_6039,N_7414);
xnor U9417 (N_9417,N_6841,N_5533);
or U9418 (N_9418,N_5701,N_7449);
and U9419 (N_9419,N_5476,N_5685);
nand U9420 (N_9420,N_5459,N_6175);
nand U9421 (N_9421,N_7410,N_5520);
or U9422 (N_9422,N_6352,N_5401);
nand U9423 (N_9423,N_6003,N_5340);
and U9424 (N_9424,N_6897,N_6198);
and U9425 (N_9425,N_5380,N_5403);
nand U9426 (N_9426,N_5352,N_6705);
and U9427 (N_9427,N_7445,N_7355);
xnor U9428 (N_9428,N_6095,N_6953);
nor U9429 (N_9429,N_7208,N_5739);
nand U9430 (N_9430,N_6038,N_7485);
nand U9431 (N_9431,N_6681,N_6063);
xor U9432 (N_9432,N_5177,N_6237);
nor U9433 (N_9433,N_5831,N_6227);
and U9434 (N_9434,N_6087,N_5413);
nor U9435 (N_9435,N_5876,N_6410);
and U9436 (N_9436,N_5562,N_7170);
and U9437 (N_9437,N_7439,N_5798);
and U9438 (N_9438,N_7179,N_5861);
nand U9439 (N_9439,N_6913,N_7273);
or U9440 (N_9440,N_6547,N_5298);
xor U9441 (N_9441,N_5750,N_5891);
and U9442 (N_9442,N_6039,N_6576);
and U9443 (N_9443,N_7498,N_7426);
xor U9444 (N_9444,N_6215,N_5747);
nor U9445 (N_9445,N_5709,N_7334);
xnor U9446 (N_9446,N_7138,N_6436);
xnor U9447 (N_9447,N_5927,N_6412);
nand U9448 (N_9448,N_6230,N_5011);
nand U9449 (N_9449,N_7458,N_6780);
and U9450 (N_9450,N_5472,N_5807);
and U9451 (N_9451,N_7305,N_5362);
nor U9452 (N_9452,N_5513,N_6089);
xor U9453 (N_9453,N_7272,N_5168);
xor U9454 (N_9454,N_5794,N_5577);
nor U9455 (N_9455,N_5556,N_5266);
nand U9456 (N_9456,N_6504,N_5722);
and U9457 (N_9457,N_6082,N_7089);
or U9458 (N_9458,N_5732,N_6856);
nand U9459 (N_9459,N_5063,N_5314);
or U9460 (N_9460,N_6133,N_6853);
nor U9461 (N_9461,N_5408,N_6859);
and U9462 (N_9462,N_6790,N_7216);
nor U9463 (N_9463,N_5158,N_5483);
and U9464 (N_9464,N_6726,N_7246);
or U9465 (N_9465,N_6418,N_5112);
nand U9466 (N_9466,N_7362,N_7021);
nor U9467 (N_9467,N_6756,N_6087);
xnor U9468 (N_9468,N_5830,N_7467);
nand U9469 (N_9469,N_5927,N_6191);
or U9470 (N_9470,N_7171,N_6633);
xor U9471 (N_9471,N_5273,N_7287);
nand U9472 (N_9472,N_5321,N_6123);
nand U9473 (N_9473,N_6260,N_5689);
or U9474 (N_9474,N_6024,N_5944);
and U9475 (N_9475,N_5785,N_5612);
xnor U9476 (N_9476,N_5280,N_7052);
or U9477 (N_9477,N_7156,N_6968);
xor U9478 (N_9478,N_5213,N_6953);
nand U9479 (N_9479,N_5209,N_5478);
or U9480 (N_9480,N_5600,N_6513);
or U9481 (N_9481,N_6325,N_6029);
xnor U9482 (N_9482,N_6340,N_6630);
or U9483 (N_9483,N_6114,N_6708);
and U9484 (N_9484,N_5173,N_6095);
nor U9485 (N_9485,N_5953,N_5352);
and U9486 (N_9486,N_6235,N_7059);
or U9487 (N_9487,N_6019,N_5593);
and U9488 (N_9488,N_5977,N_7038);
or U9489 (N_9489,N_6535,N_6097);
and U9490 (N_9490,N_6057,N_5123);
nand U9491 (N_9491,N_5889,N_6116);
and U9492 (N_9492,N_5035,N_6325);
nand U9493 (N_9493,N_5078,N_7382);
xor U9494 (N_9494,N_6756,N_7427);
xor U9495 (N_9495,N_5351,N_6592);
nor U9496 (N_9496,N_5852,N_6549);
xor U9497 (N_9497,N_5262,N_6514);
nand U9498 (N_9498,N_7323,N_5661);
or U9499 (N_9499,N_6948,N_5108);
xnor U9500 (N_9500,N_6234,N_6519);
nor U9501 (N_9501,N_5409,N_6866);
nand U9502 (N_9502,N_7337,N_6346);
xor U9503 (N_9503,N_7064,N_7074);
nor U9504 (N_9504,N_6036,N_6832);
or U9505 (N_9505,N_6614,N_5871);
xor U9506 (N_9506,N_6991,N_6184);
nand U9507 (N_9507,N_7396,N_5427);
and U9508 (N_9508,N_5125,N_5262);
nand U9509 (N_9509,N_7161,N_6745);
xor U9510 (N_9510,N_5131,N_6839);
nor U9511 (N_9511,N_6150,N_6980);
nor U9512 (N_9512,N_6425,N_7258);
xnor U9513 (N_9513,N_5817,N_5533);
nand U9514 (N_9514,N_6807,N_5382);
nor U9515 (N_9515,N_5128,N_7182);
nor U9516 (N_9516,N_7081,N_6690);
and U9517 (N_9517,N_5608,N_5800);
nand U9518 (N_9518,N_6085,N_7291);
nor U9519 (N_9519,N_7209,N_6943);
nand U9520 (N_9520,N_7243,N_5049);
and U9521 (N_9521,N_6452,N_7317);
nand U9522 (N_9522,N_5883,N_6357);
or U9523 (N_9523,N_7087,N_5451);
nand U9524 (N_9524,N_6578,N_5259);
and U9525 (N_9525,N_5099,N_7172);
xor U9526 (N_9526,N_5512,N_6361);
or U9527 (N_9527,N_5483,N_7176);
or U9528 (N_9528,N_5519,N_6953);
nor U9529 (N_9529,N_5018,N_6120);
nor U9530 (N_9530,N_6673,N_6469);
nor U9531 (N_9531,N_5747,N_6164);
or U9532 (N_9532,N_6605,N_5761);
nor U9533 (N_9533,N_5906,N_6171);
or U9534 (N_9534,N_7464,N_7250);
nor U9535 (N_9535,N_6332,N_5578);
xnor U9536 (N_9536,N_6217,N_5648);
or U9537 (N_9537,N_7395,N_5834);
xor U9538 (N_9538,N_6588,N_5096);
and U9539 (N_9539,N_5307,N_5455);
and U9540 (N_9540,N_6964,N_6658);
and U9541 (N_9541,N_5153,N_6396);
nand U9542 (N_9542,N_6815,N_6598);
or U9543 (N_9543,N_5462,N_6997);
nor U9544 (N_9544,N_6430,N_6952);
or U9545 (N_9545,N_6774,N_7263);
nand U9546 (N_9546,N_7323,N_7022);
or U9547 (N_9547,N_5094,N_5272);
nand U9548 (N_9548,N_7240,N_5476);
or U9549 (N_9549,N_5412,N_7250);
or U9550 (N_9550,N_7232,N_5374);
xnor U9551 (N_9551,N_6939,N_7089);
nand U9552 (N_9552,N_6437,N_5317);
xor U9553 (N_9553,N_5656,N_6886);
xor U9554 (N_9554,N_5925,N_5227);
or U9555 (N_9555,N_5412,N_6175);
or U9556 (N_9556,N_5649,N_5181);
and U9557 (N_9557,N_7419,N_6162);
nor U9558 (N_9558,N_6547,N_5605);
or U9559 (N_9559,N_5011,N_5925);
nand U9560 (N_9560,N_7074,N_5350);
xnor U9561 (N_9561,N_6073,N_6461);
or U9562 (N_9562,N_6398,N_5765);
nand U9563 (N_9563,N_5738,N_5788);
nor U9564 (N_9564,N_5590,N_5548);
nor U9565 (N_9565,N_5271,N_5910);
xnor U9566 (N_9566,N_5092,N_5901);
and U9567 (N_9567,N_7309,N_7202);
or U9568 (N_9568,N_7155,N_5415);
nand U9569 (N_9569,N_5491,N_7135);
or U9570 (N_9570,N_7464,N_6038);
or U9571 (N_9571,N_6018,N_6917);
or U9572 (N_9572,N_5486,N_6353);
xnor U9573 (N_9573,N_7229,N_5390);
xor U9574 (N_9574,N_6148,N_7334);
or U9575 (N_9575,N_5362,N_5701);
xor U9576 (N_9576,N_6208,N_6785);
xor U9577 (N_9577,N_6983,N_6780);
xnor U9578 (N_9578,N_7165,N_5491);
or U9579 (N_9579,N_5350,N_7480);
xnor U9580 (N_9580,N_6020,N_7082);
xor U9581 (N_9581,N_5599,N_5983);
nand U9582 (N_9582,N_5312,N_6948);
or U9583 (N_9583,N_7416,N_6834);
or U9584 (N_9584,N_6759,N_6142);
xnor U9585 (N_9585,N_6292,N_6804);
xor U9586 (N_9586,N_5131,N_5478);
nand U9587 (N_9587,N_6833,N_5996);
xor U9588 (N_9588,N_6622,N_7342);
xor U9589 (N_9589,N_5058,N_6982);
or U9590 (N_9590,N_6019,N_6249);
nor U9591 (N_9591,N_7240,N_5123);
nor U9592 (N_9592,N_5169,N_6478);
and U9593 (N_9593,N_7172,N_7112);
nand U9594 (N_9594,N_7257,N_6899);
nand U9595 (N_9595,N_7424,N_5597);
nor U9596 (N_9596,N_6702,N_5145);
and U9597 (N_9597,N_6134,N_5843);
xnor U9598 (N_9598,N_6644,N_6478);
nand U9599 (N_9599,N_7113,N_6717);
nor U9600 (N_9600,N_5047,N_6116);
nand U9601 (N_9601,N_7109,N_5719);
nor U9602 (N_9602,N_6445,N_5352);
xor U9603 (N_9603,N_6122,N_5626);
and U9604 (N_9604,N_5553,N_6847);
or U9605 (N_9605,N_5360,N_5031);
nor U9606 (N_9606,N_6556,N_6590);
or U9607 (N_9607,N_5401,N_5953);
or U9608 (N_9608,N_5255,N_7325);
nor U9609 (N_9609,N_5506,N_6597);
nor U9610 (N_9610,N_6206,N_5770);
or U9611 (N_9611,N_5717,N_6047);
xor U9612 (N_9612,N_6001,N_6550);
nor U9613 (N_9613,N_7062,N_6115);
and U9614 (N_9614,N_6820,N_5339);
xnor U9615 (N_9615,N_5705,N_5628);
nand U9616 (N_9616,N_7313,N_6592);
and U9617 (N_9617,N_7311,N_7345);
nor U9618 (N_9618,N_6889,N_5847);
nand U9619 (N_9619,N_7158,N_5044);
or U9620 (N_9620,N_7277,N_6505);
nor U9621 (N_9621,N_5254,N_5263);
and U9622 (N_9622,N_7157,N_7401);
or U9623 (N_9623,N_6990,N_5204);
nor U9624 (N_9624,N_5131,N_5279);
xor U9625 (N_9625,N_5758,N_6879);
nor U9626 (N_9626,N_7313,N_5413);
nand U9627 (N_9627,N_6499,N_6621);
xor U9628 (N_9628,N_6824,N_5792);
and U9629 (N_9629,N_6349,N_5916);
or U9630 (N_9630,N_5844,N_5407);
and U9631 (N_9631,N_5180,N_7379);
and U9632 (N_9632,N_6752,N_7040);
nor U9633 (N_9633,N_5986,N_6219);
or U9634 (N_9634,N_6446,N_5032);
or U9635 (N_9635,N_6496,N_5454);
and U9636 (N_9636,N_5910,N_5673);
nand U9637 (N_9637,N_7315,N_6022);
nor U9638 (N_9638,N_7173,N_5328);
or U9639 (N_9639,N_7190,N_6240);
xnor U9640 (N_9640,N_5825,N_6943);
xnor U9641 (N_9641,N_6069,N_5990);
or U9642 (N_9642,N_7146,N_5804);
nor U9643 (N_9643,N_7493,N_6182);
nand U9644 (N_9644,N_5184,N_6112);
nor U9645 (N_9645,N_5845,N_5258);
xnor U9646 (N_9646,N_5129,N_5662);
or U9647 (N_9647,N_5145,N_6060);
and U9648 (N_9648,N_7070,N_7456);
xnor U9649 (N_9649,N_6644,N_6790);
or U9650 (N_9650,N_6917,N_6350);
xnor U9651 (N_9651,N_6415,N_6781);
or U9652 (N_9652,N_5730,N_7256);
nor U9653 (N_9653,N_7038,N_6016);
xnor U9654 (N_9654,N_6831,N_5978);
and U9655 (N_9655,N_6608,N_5327);
xnor U9656 (N_9656,N_5736,N_5570);
and U9657 (N_9657,N_6931,N_6210);
and U9658 (N_9658,N_6493,N_6828);
nor U9659 (N_9659,N_5878,N_5765);
nor U9660 (N_9660,N_5549,N_6471);
or U9661 (N_9661,N_6852,N_5393);
nor U9662 (N_9662,N_6786,N_6662);
xor U9663 (N_9663,N_5907,N_6774);
nor U9664 (N_9664,N_5754,N_6813);
and U9665 (N_9665,N_6958,N_5841);
xor U9666 (N_9666,N_6393,N_5025);
nor U9667 (N_9667,N_6535,N_5516);
xnor U9668 (N_9668,N_5814,N_7462);
xnor U9669 (N_9669,N_6329,N_6860);
nor U9670 (N_9670,N_7424,N_6891);
nand U9671 (N_9671,N_6732,N_5313);
and U9672 (N_9672,N_6135,N_7142);
nand U9673 (N_9673,N_6978,N_5291);
or U9674 (N_9674,N_5798,N_5979);
or U9675 (N_9675,N_6795,N_6819);
nand U9676 (N_9676,N_7158,N_5506);
and U9677 (N_9677,N_7011,N_6236);
nand U9678 (N_9678,N_5751,N_5503);
nand U9679 (N_9679,N_7382,N_6060);
and U9680 (N_9680,N_5669,N_6590);
nand U9681 (N_9681,N_6757,N_6664);
xnor U9682 (N_9682,N_6557,N_6193);
and U9683 (N_9683,N_7297,N_6768);
xor U9684 (N_9684,N_7145,N_5761);
or U9685 (N_9685,N_5467,N_5324);
nor U9686 (N_9686,N_5692,N_6560);
and U9687 (N_9687,N_7433,N_5222);
or U9688 (N_9688,N_6631,N_5097);
nor U9689 (N_9689,N_5929,N_5649);
or U9690 (N_9690,N_5435,N_5733);
nor U9691 (N_9691,N_5623,N_6961);
nand U9692 (N_9692,N_5288,N_5724);
nand U9693 (N_9693,N_5430,N_7348);
nor U9694 (N_9694,N_5020,N_6561);
or U9695 (N_9695,N_5583,N_6088);
nor U9696 (N_9696,N_6023,N_7302);
nor U9697 (N_9697,N_7407,N_6013);
xor U9698 (N_9698,N_6779,N_6572);
xnor U9699 (N_9699,N_5450,N_5967);
nand U9700 (N_9700,N_7207,N_5823);
and U9701 (N_9701,N_6815,N_6799);
xor U9702 (N_9702,N_5568,N_6203);
and U9703 (N_9703,N_5191,N_6736);
xnor U9704 (N_9704,N_5878,N_5641);
nor U9705 (N_9705,N_5998,N_5768);
xor U9706 (N_9706,N_6535,N_6738);
xnor U9707 (N_9707,N_7314,N_5542);
nand U9708 (N_9708,N_7141,N_7230);
nand U9709 (N_9709,N_5386,N_6300);
nand U9710 (N_9710,N_5666,N_5564);
nand U9711 (N_9711,N_7255,N_5011);
or U9712 (N_9712,N_7444,N_6958);
or U9713 (N_9713,N_6903,N_6294);
and U9714 (N_9714,N_7388,N_7251);
xor U9715 (N_9715,N_6263,N_5945);
nor U9716 (N_9716,N_5704,N_7279);
nor U9717 (N_9717,N_5291,N_7438);
or U9718 (N_9718,N_6971,N_6692);
nand U9719 (N_9719,N_7449,N_7317);
xnor U9720 (N_9720,N_6000,N_5731);
or U9721 (N_9721,N_6938,N_5635);
nor U9722 (N_9722,N_7381,N_6717);
and U9723 (N_9723,N_7454,N_7388);
and U9724 (N_9724,N_6597,N_5336);
xor U9725 (N_9725,N_6644,N_6632);
nor U9726 (N_9726,N_6392,N_6114);
or U9727 (N_9727,N_5797,N_6597);
and U9728 (N_9728,N_7282,N_5769);
and U9729 (N_9729,N_6411,N_5283);
xor U9730 (N_9730,N_7423,N_5656);
and U9731 (N_9731,N_6849,N_6648);
and U9732 (N_9732,N_5351,N_5824);
and U9733 (N_9733,N_5795,N_6077);
and U9734 (N_9734,N_6948,N_6005);
nand U9735 (N_9735,N_6557,N_5913);
and U9736 (N_9736,N_5635,N_6108);
nor U9737 (N_9737,N_5345,N_5111);
or U9738 (N_9738,N_6407,N_5172);
xor U9739 (N_9739,N_5660,N_5540);
and U9740 (N_9740,N_5063,N_5946);
nor U9741 (N_9741,N_6971,N_6873);
nor U9742 (N_9742,N_5385,N_6444);
nand U9743 (N_9743,N_6634,N_6885);
nand U9744 (N_9744,N_5860,N_6177);
and U9745 (N_9745,N_7489,N_7239);
nor U9746 (N_9746,N_6583,N_5194);
xnor U9747 (N_9747,N_6417,N_6117);
xor U9748 (N_9748,N_7220,N_7065);
nand U9749 (N_9749,N_5040,N_6789);
nor U9750 (N_9750,N_6071,N_6473);
nor U9751 (N_9751,N_6090,N_6486);
xor U9752 (N_9752,N_5862,N_7206);
nor U9753 (N_9753,N_5023,N_7473);
and U9754 (N_9754,N_6139,N_5418);
nor U9755 (N_9755,N_5901,N_5835);
or U9756 (N_9756,N_6719,N_7013);
nor U9757 (N_9757,N_5086,N_5776);
nand U9758 (N_9758,N_6161,N_5300);
and U9759 (N_9759,N_6025,N_6467);
nand U9760 (N_9760,N_5851,N_5148);
nor U9761 (N_9761,N_5160,N_5269);
nor U9762 (N_9762,N_5134,N_5293);
and U9763 (N_9763,N_5210,N_6383);
nor U9764 (N_9764,N_6675,N_6176);
xnor U9765 (N_9765,N_5139,N_6440);
or U9766 (N_9766,N_6078,N_7455);
or U9767 (N_9767,N_5320,N_7139);
or U9768 (N_9768,N_7122,N_7310);
and U9769 (N_9769,N_5291,N_5737);
nand U9770 (N_9770,N_6914,N_6306);
xor U9771 (N_9771,N_5518,N_7154);
or U9772 (N_9772,N_6632,N_6514);
nor U9773 (N_9773,N_5152,N_6837);
nor U9774 (N_9774,N_6944,N_7486);
nor U9775 (N_9775,N_7089,N_6846);
xnor U9776 (N_9776,N_6048,N_5762);
xor U9777 (N_9777,N_7397,N_6445);
xor U9778 (N_9778,N_6689,N_7212);
xnor U9779 (N_9779,N_7477,N_6858);
or U9780 (N_9780,N_6014,N_5403);
xor U9781 (N_9781,N_5485,N_6606);
xnor U9782 (N_9782,N_6087,N_5920);
and U9783 (N_9783,N_5123,N_5421);
or U9784 (N_9784,N_5220,N_7200);
nand U9785 (N_9785,N_5807,N_7143);
nand U9786 (N_9786,N_6973,N_7253);
xnor U9787 (N_9787,N_6978,N_5088);
nand U9788 (N_9788,N_5967,N_6501);
and U9789 (N_9789,N_5714,N_5534);
or U9790 (N_9790,N_5856,N_7122);
or U9791 (N_9791,N_7380,N_6227);
nand U9792 (N_9792,N_7318,N_6412);
and U9793 (N_9793,N_6705,N_7406);
nand U9794 (N_9794,N_6905,N_5383);
nand U9795 (N_9795,N_7022,N_7298);
nor U9796 (N_9796,N_5680,N_6920);
xnor U9797 (N_9797,N_5127,N_6333);
or U9798 (N_9798,N_5779,N_6294);
xor U9799 (N_9799,N_7335,N_5247);
nand U9800 (N_9800,N_7095,N_6404);
nand U9801 (N_9801,N_7375,N_6615);
nor U9802 (N_9802,N_6255,N_6150);
nand U9803 (N_9803,N_6338,N_5359);
or U9804 (N_9804,N_7411,N_6273);
and U9805 (N_9805,N_6113,N_7444);
xnor U9806 (N_9806,N_5678,N_5339);
and U9807 (N_9807,N_7036,N_5874);
or U9808 (N_9808,N_5763,N_5157);
and U9809 (N_9809,N_7416,N_5176);
or U9810 (N_9810,N_6683,N_6730);
or U9811 (N_9811,N_6000,N_5133);
xnor U9812 (N_9812,N_5418,N_5872);
nand U9813 (N_9813,N_5274,N_7431);
or U9814 (N_9814,N_5083,N_5334);
nor U9815 (N_9815,N_6832,N_7194);
or U9816 (N_9816,N_7259,N_7000);
nor U9817 (N_9817,N_6791,N_6237);
nor U9818 (N_9818,N_6152,N_5155);
xnor U9819 (N_9819,N_5093,N_6850);
or U9820 (N_9820,N_5192,N_7045);
nand U9821 (N_9821,N_6965,N_7033);
nor U9822 (N_9822,N_6751,N_7139);
nor U9823 (N_9823,N_7441,N_6740);
nor U9824 (N_9824,N_6195,N_7224);
or U9825 (N_9825,N_5267,N_6110);
nand U9826 (N_9826,N_7332,N_6664);
nand U9827 (N_9827,N_6492,N_6776);
nor U9828 (N_9828,N_7033,N_6018);
and U9829 (N_9829,N_5629,N_6557);
nor U9830 (N_9830,N_5052,N_7454);
or U9831 (N_9831,N_7316,N_6254);
and U9832 (N_9832,N_6574,N_7396);
nor U9833 (N_9833,N_6884,N_6883);
nand U9834 (N_9834,N_5035,N_6157);
and U9835 (N_9835,N_5561,N_6592);
nor U9836 (N_9836,N_5350,N_5054);
xor U9837 (N_9837,N_6157,N_5754);
or U9838 (N_9838,N_6950,N_7243);
nor U9839 (N_9839,N_6925,N_7211);
xnor U9840 (N_9840,N_6082,N_5550);
xnor U9841 (N_9841,N_6213,N_5710);
xnor U9842 (N_9842,N_5420,N_6090);
or U9843 (N_9843,N_5209,N_5281);
nor U9844 (N_9844,N_6940,N_7104);
xnor U9845 (N_9845,N_6686,N_6945);
xor U9846 (N_9846,N_5020,N_6008);
and U9847 (N_9847,N_7252,N_7384);
nor U9848 (N_9848,N_6871,N_5882);
and U9849 (N_9849,N_7077,N_5673);
and U9850 (N_9850,N_5954,N_5575);
and U9851 (N_9851,N_5389,N_6275);
xnor U9852 (N_9852,N_6981,N_6996);
or U9853 (N_9853,N_6384,N_6842);
nand U9854 (N_9854,N_6844,N_7239);
nand U9855 (N_9855,N_5751,N_5007);
nor U9856 (N_9856,N_7451,N_6017);
or U9857 (N_9857,N_7359,N_6378);
xnor U9858 (N_9858,N_6508,N_6435);
and U9859 (N_9859,N_6056,N_5306);
xor U9860 (N_9860,N_7265,N_5161);
xor U9861 (N_9861,N_5785,N_5959);
nand U9862 (N_9862,N_6595,N_5108);
nand U9863 (N_9863,N_6382,N_5506);
and U9864 (N_9864,N_6852,N_7492);
nand U9865 (N_9865,N_5774,N_6012);
xor U9866 (N_9866,N_6577,N_5265);
nand U9867 (N_9867,N_7061,N_6413);
or U9868 (N_9868,N_7366,N_5156);
or U9869 (N_9869,N_5516,N_6052);
xnor U9870 (N_9870,N_6708,N_5456);
xnor U9871 (N_9871,N_6931,N_7347);
nor U9872 (N_9872,N_7367,N_7482);
nor U9873 (N_9873,N_5850,N_6081);
or U9874 (N_9874,N_5564,N_5998);
nand U9875 (N_9875,N_5597,N_6729);
nand U9876 (N_9876,N_7043,N_7239);
nand U9877 (N_9877,N_6237,N_5257);
nand U9878 (N_9878,N_5496,N_6677);
nand U9879 (N_9879,N_6975,N_7344);
xnor U9880 (N_9880,N_5891,N_6337);
xnor U9881 (N_9881,N_6509,N_6300);
or U9882 (N_9882,N_7262,N_7485);
nor U9883 (N_9883,N_5488,N_6053);
nand U9884 (N_9884,N_5214,N_6590);
nand U9885 (N_9885,N_5902,N_5791);
nand U9886 (N_9886,N_6719,N_5885);
xor U9887 (N_9887,N_6469,N_7413);
or U9888 (N_9888,N_6359,N_5699);
xor U9889 (N_9889,N_7462,N_5942);
or U9890 (N_9890,N_6023,N_5071);
or U9891 (N_9891,N_5445,N_7286);
and U9892 (N_9892,N_5784,N_7038);
or U9893 (N_9893,N_6019,N_6910);
and U9894 (N_9894,N_5230,N_6417);
nand U9895 (N_9895,N_6519,N_5612);
and U9896 (N_9896,N_6349,N_6931);
xnor U9897 (N_9897,N_7114,N_5916);
and U9898 (N_9898,N_7159,N_5140);
or U9899 (N_9899,N_6318,N_6064);
or U9900 (N_9900,N_7146,N_6419);
xnor U9901 (N_9901,N_6211,N_5318);
nor U9902 (N_9902,N_5159,N_6293);
nor U9903 (N_9903,N_5640,N_6339);
xnor U9904 (N_9904,N_6324,N_7432);
nand U9905 (N_9905,N_6848,N_5840);
and U9906 (N_9906,N_6031,N_5273);
nand U9907 (N_9907,N_5751,N_5494);
and U9908 (N_9908,N_5000,N_6633);
or U9909 (N_9909,N_5862,N_5624);
nor U9910 (N_9910,N_6365,N_5841);
or U9911 (N_9911,N_5141,N_7410);
nand U9912 (N_9912,N_6732,N_5642);
nor U9913 (N_9913,N_6885,N_6689);
nand U9914 (N_9914,N_7009,N_5646);
or U9915 (N_9915,N_6627,N_6733);
and U9916 (N_9916,N_5540,N_7178);
nand U9917 (N_9917,N_6946,N_7460);
nor U9918 (N_9918,N_7414,N_6546);
nor U9919 (N_9919,N_5799,N_5791);
xnor U9920 (N_9920,N_5927,N_7221);
and U9921 (N_9921,N_6117,N_7357);
xor U9922 (N_9922,N_6705,N_6893);
and U9923 (N_9923,N_6836,N_6962);
and U9924 (N_9924,N_5439,N_6319);
xor U9925 (N_9925,N_6805,N_7367);
nand U9926 (N_9926,N_5176,N_6058);
and U9927 (N_9927,N_5419,N_7056);
or U9928 (N_9928,N_7100,N_7137);
and U9929 (N_9929,N_7123,N_7363);
and U9930 (N_9930,N_5971,N_6314);
xnor U9931 (N_9931,N_5769,N_6391);
xnor U9932 (N_9932,N_7370,N_7371);
nand U9933 (N_9933,N_7003,N_7239);
and U9934 (N_9934,N_5723,N_6568);
or U9935 (N_9935,N_7133,N_7287);
and U9936 (N_9936,N_7090,N_7129);
xor U9937 (N_9937,N_6179,N_6719);
and U9938 (N_9938,N_5346,N_6618);
and U9939 (N_9939,N_6681,N_6640);
nand U9940 (N_9940,N_5893,N_7031);
nand U9941 (N_9941,N_7474,N_6714);
nor U9942 (N_9942,N_5669,N_7117);
xor U9943 (N_9943,N_6816,N_7216);
nand U9944 (N_9944,N_6410,N_7112);
and U9945 (N_9945,N_6471,N_5075);
or U9946 (N_9946,N_5805,N_6303);
nor U9947 (N_9947,N_6906,N_6273);
or U9948 (N_9948,N_5365,N_6716);
xor U9949 (N_9949,N_6843,N_5694);
and U9950 (N_9950,N_6611,N_6208);
nand U9951 (N_9951,N_6517,N_7327);
xnor U9952 (N_9952,N_5586,N_6265);
nand U9953 (N_9953,N_5179,N_6980);
or U9954 (N_9954,N_6719,N_6661);
nor U9955 (N_9955,N_6983,N_6119);
and U9956 (N_9956,N_6033,N_5373);
nor U9957 (N_9957,N_6767,N_5784);
nor U9958 (N_9958,N_5121,N_6709);
or U9959 (N_9959,N_7187,N_6157);
and U9960 (N_9960,N_5757,N_7040);
nand U9961 (N_9961,N_6771,N_6246);
or U9962 (N_9962,N_5824,N_5151);
nor U9963 (N_9963,N_7076,N_5818);
or U9964 (N_9964,N_6072,N_6313);
or U9965 (N_9965,N_6222,N_7164);
xor U9966 (N_9966,N_6058,N_6967);
or U9967 (N_9967,N_6031,N_6670);
or U9968 (N_9968,N_6946,N_6209);
xor U9969 (N_9969,N_5541,N_6047);
xnor U9970 (N_9970,N_7038,N_7185);
xor U9971 (N_9971,N_6882,N_7324);
nand U9972 (N_9972,N_6106,N_5390);
xor U9973 (N_9973,N_7301,N_6771);
nand U9974 (N_9974,N_6637,N_7443);
nor U9975 (N_9975,N_7409,N_6281);
nand U9976 (N_9976,N_6167,N_5782);
nand U9977 (N_9977,N_5467,N_6347);
and U9978 (N_9978,N_5704,N_7103);
xnor U9979 (N_9979,N_6759,N_5311);
nor U9980 (N_9980,N_5849,N_6667);
nand U9981 (N_9981,N_6297,N_5632);
xnor U9982 (N_9982,N_7271,N_5171);
nand U9983 (N_9983,N_6482,N_6254);
and U9984 (N_9984,N_5839,N_5651);
nor U9985 (N_9985,N_6135,N_7339);
nand U9986 (N_9986,N_7489,N_7238);
nand U9987 (N_9987,N_6203,N_6702);
and U9988 (N_9988,N_5449,N_6543);
xnor U9989 (N_9989,N_5469,N_6732);
nand U9990 (N_9990,N_7413,N_7287);
nand U9991 (N_9991,N_7118,N_5749);
xor U9992 (N_9992,N_5673,N_6183);
or U9993 (N_9993,N_6962,N_5831);
or U9994 (N_9994,N_5989,N_5683);
nand U9995 (N_9995,N_6100,N_6617);
nor U9996 (N_9996,N_5546,N_7476);
or U9997 (N_9997,N_5339,N_5626);
nor U9998 (N_9998,N_6585,N_7473);
xor U9999 (N_9999,N_5062,N_5844);
and U10000 (N_10000,N_9871,N_7655);
nand U10001 (N_10001,N_8773,N_9600);
or U10002 (N_10002,N_9221,N_9073);
and U10003 (N_10003,N_9747,N_9301);
or U10004 (N_10004,N_9647,N_8678);
and U10005 (N_10005,N_8038,N_8606);
nand U10006 (N_10006,N_9344,N_9272);
nor U10007 (N_10007,N_9754,N_9827);
nand U10008 (N_10008,N_8858,N_7981);
nor U10009 (N_10009,N_8547,N_9205);
xnor U10010 (N_10010,N_8433,N_8629);
nor U10011 (N_10011,N_8745,N_9673);
or U10012 (N_10012,N_7987,N_7750);
nor U10013 (N_10013,N_7818,N_8125);
nor U10014 (N_10014,N_8541,N_7714);
xor U10015 (N_10015,N_9079,N_8870);
nand U10016 (N_10016,N_7680,N_7632);
nor U10017 (N_10017,N_9651,N_8388);
nand U10018 (N_10018,N_8073,N_9588);
nand U10019 (N_10019,N_9504,N_9749);
nor U10020 (N_10020,N_9609,N_8410);
or U10021 (N_10021,N_8015,N_8001);
or U10022 (N_10022,N_8810,N_9139);
or U10023 (N_10023,N_7914,N_9040);
xnor U10024 (N_10024,N_7940,N_9564);
nand U10025 (N_10025,N_9652,N_9523);
nand U10026 (N_10026,N_7924,N_8317);
or U10027 (N_10027,N_8123,N_8943);
nand U10028 (N_10028,N_8288,N_7595);
and U10029 (N_10029,N_9218,N_8998);
and U10030 (N_10030,N_7596,N_7722);
xor U10031 (N_10031,N_9349,N_9659);
nand U10032 (N_10032,N_9689,N_7705);
xor U10033 (N_10033,N_9922,N_9878);
or U10034 (N_10034,N_8596,N_7541);
or U10035 (N_10035,N_8489,N_9374);
xnor U10036 (N_10036,N_9741,N_8173);
xnor U10037 (N_10037,N_8681,N_9416);
or U10038 (N_10038,N_9787,N_8331);
nor U10039 (N_10039,N_9880,N_8270);
nor U10040 (N_10040,N_7540,N_9985);
or U10041 (N_10041,N_9126,N_9257);
and U10042 (N_10042,N_8281,N_9602);
nand U10043 (N_10043,N_8240,N_7549);
nor U10044 (N_10044,N_7839,N_9026);
or U10045 (N_10045,N_9593,N_8386);
nor U10046 (N_10046,N_9122,N_9382);
xor U10047 (N_10047,N_8222,N_9107);
and U10048 (N_10048,N_8689,N_9945);
and U10049 (N_10049,N_9797,N_7647);
nand U10050 (N_10050,N_8688,N_7737);
xor U10051 (N_10051,N_8712,N_8490);
xnor U10052 (N_10052,N_9840,N_7863);
or U10053 (N_10053,N_9315,N_8828);
or U10054 (N_10054,N_7523,N_8566);
nor U10055 (N_10055,N_9693,N_9502);
or U10056 (N_10056,N_8441,N_9406);
nand U10057 (N_10057,N_9043,N_8151);
nand U10058 (N_10058,N_9882,N_7889);
or U10059 (N_10059,N_9944,N_9543);
xnor U10060 (N_10060,N_8285,N_8319);
nand U10061 (N_10061,N_7600,N_7520);
or U10062 (N_10062,N_9032,N_8742);
nand U10063 (N_10063,N_7659,N_9118);
nand U10064 (N_10064,N_9428,N_9553);
and U10065 (N_10065,N_8508,N_9901);
or U10066 (N_10066,N_8289,N_8819);
nor U10067 (N_10067,N_9486,N_8776);
or U10068 (N_10068,N_7898,N_9756);
or U10069 (N_10069,N_8152,N_8396);
nor U10070 (N_10070,N_9595,N_8967);
and U10071 (N_10071,N_9070,N_8572);
and U10072 (N_10072,N_7920,N_9669);
or U10073 (N_10073,N_8296,N_9608);
or U10074 (N_10074,N_8725,N_9597);
and U10075 (N_10075,N_9303,N_8393);
nor U10076 (N_10076,N_9391,N_7525);
or U10077 (N_10077,N_7629,N_9851);
nor U10078 (N_10078,N_9239,N_8018);
xnor U10079 (N_10079,N_8461,N_8956);
and U10080 (N_10080,N_8932,N_9343);
xnor U10081 (N_10081,N_8590,N_9411);
or U10082 (N_10082,N_7663,N_8275);
or U10083 (N_10083,N_7562,N_9801);
and U10084 (N_10084,N_9852,N_8219);
or U10085 (N_10085,N_9816,N_8201);
or U10086 (N_10086,N_9215,N_8363);
nand U10087 (N_10087,N_9568,N_8183);
nor U10088 (N_10088,N_8320,N_9764);
nor U10089 (N_10089,N_8752,N_7650);
xor U10090 (N_10090,N_7518,N_7929);
or U10091 (N_10091,N_9183,N_7753);
or U10092 (N_10092,N_9578,N_8579);
and U10093 (N_10093,N_8595,N_9022);
xor U10094 (N_10094,N_7843,N_9772);
nand U10095 (N_10095,N_8326,N_8834);
and U10096 (N_10096,N_8782,N_9622);
or U10097 (N_10097,N_9630,N_9738);
nand U10098 (N_10098,N_9003,N_7618);
xnor U10099 (N_10099,N_8966,N_8225);
nand U10100 (N_10100,N_8592,N_9974);
xor U10101 (N_10101,N_8093,N_8087);
nand U10102 (N_10102,N_7891,N_9368);
nand U10103 (N_10103,N_9463,N_8497);
and U10104 (N_10104,N_9933,N_9113);
nor U10105 (N_10105,N_9238,N_7698);
or U10106 (N_10106,N_9867,N_8822);
or U10107 (N_10107,N_8677,N_8116);
nor U10108 (N_10108,N_8243,N_8069);
nor U10109 (N_10109,N_8658,N_9292);
or U10110 (N_10110,N_7997,N_8013);
nand U10111 (N_10111,N_8504,N_9781);
nor U10112 (N_10112,N_7746,N_7921);
and U10113 (N_10113,N_8733,N_7962);
or U10114 (N_10114,N_9488,N_8276);
nor U10115 (N_10115,N_9240,N_8696);
and U10116 (N_10116,N_8821,N_9033);
nor U10117 (N_10117,N_9063,N_8160);
xnor U10118 (N_10118,N_9972,N_9431);
and U10119 (N_10119,N_9132,N_8909);
nor U10120 (N_10120,N_8884,N_8652);
nand U10121 (N_10121,N_9761,N_7919);
xnor U10122 (N_10122,N_8163,N_8171);
and U10123 (N_10123,N_8165,N_9087);
or U10124 (N_10124,N_9295,N_8360);
nor U10125 (N_10125,N_8016,N_8362);
xor U10126 (N_10126,N_8423,N_8527);
nor U10127 (N_10127,N_8202,N_7604);
or U10128 (N_10128,N_7932,N_9655);
nor U10129 (N_10129,N_7884,N_8912);
xnor U10130 (N_10130,N_9685,N_8908);
and U10131 (N_10131,N_9104,N_8864);
nor U10132 (N_10132,N_7723,N_8984);
xnor U10133 (N_10133,N_7500,N_9581);
and U10134 (N_10134,N_7710,N_7986);
xor U10135 (N_10135,N_8898,N_7788);
nor U10136 (N_10136,N_7857,N_8398);
and U10137 (N_10137,N_9717,N_8237);
or U10138 (N_10138,N_8931,N_7909);
or U10139 (N_10139,N_9109,N_8506);
xor U10140 (N_10140,N_8211,N_9869);
nor U10141 (N_10141,N_9541,N_7777);
and U10142 (N_10142,N_9725,N_7996);
or U10143 (N_10143,N_8789,N_8722);
or U10144 (N_10144,N_8322,N_9101);
xnor U10145 (N_10145,N_8917,N_7826);
xnor U10146 (N_10146,N_7731,N_8985);
or U10147 (N_10147,N_8094,N_8124);
xor U10148 (N_10148,N_8012,N_8624);
nor U10149 (N_10149,N_7588,N_9610);
nand U10150 (N_10150,N_9847,N_9075);
and U10151 (N_10151,N_9672,N_9361);
or U10152 (N_10152,N_8389,N_8339);
xnor U10153 (N_10153,N_8394,N_8754);
and U10154 (N_10154,N_7984,N_8169);
nor U10155 (N_10155,N_7627,N_7881);
xor U10156 (N_10156,N_8346,N_8584);
nor U10157 (N_10157,N_8948,N_9373);
or U10158 (N_10158,N_7711,N_9779);
nor U10159 (N_10159,N_9188,N_9421);
nand U10160 (N_10160,N_7855,N_8006);
nor U10161 (N_10161,N_8993,N_7724);
and U10162 (N_10162,N_7886,N_9054);
nor U10163 (N_10163,N_8100,N_9489);
nor U10164 (N_10164,N_7539,N_8226);
nor U10165 (N_10165,N_8946,N_7639);
and U10166 (N_10166,N_8845,N_8418);
nor U10167 (N_10167,N_9106,N_8876);
and U10168 (N_10168,N_9895,N_9794);
or U10169 (N_10169,N_9220,N_9915);
or U10170 (N_10170,N_8888,N_9356);
and U10171 (N_10171,N_7972,N_9569);
xor U10172 (N_10172,N_7859,N_9558);
nor U10173 (N_10173,N_8848,N_9331);
and U10174 (N_10174,N_8758,N_8968);
or U10175 (N_10175,N_9358,N_9785);
and U10176 (N_10176,N_9511,N_9207);
nor U10177 (N_10177,N_9029,N_8859);
xnor U10178 (N_10178,N_8514,N_8809);
and U10179 (N_10179,N_9112,N_7586);
xnor U10180 (N_10180,N_9748,N_7736);
and U10181 (N_10181,N_7735,N_8347);
and U10182 (N_10182,N_8328,N_8559);
nand U10183 (N_10183,N_9923,N_8618);
or U10184 (N_10184,N_7558,N_9664);
or U10185 (N_10185,N_8426,N_8600);
xor U10186 (N_10186,N_7916,N_8885);
or U10187 (N_10187,N_9314,N_8891);
xor U10188 (N_10188,N_8445,N_8378);
nand U10189 (N_10189,N_9634,N_8267);
nor U10190 (N_10190,N_8768,N_9921);
nor U10191 (N_10191,N_8924,N_8313);
xor U10192 (N_10192,N_7566,N_9116);
or U10193 (N_10193,N_9500,N_9067);
and U10194 (N_10194,N_9582,N_9025);
or U10195 (N_10195,N_8027,N_7738);
xnor U10196 (N_10196,N_8042,N_9081);
nor U10197 (N_10197,N_8991,N_8464);
or U10198 (N_10198,N_8247,N_9963);
and U10199 (N_10199,N_8673,N_9249);
nand U10200 (N_10200,N_8692,N_7707);
xnor U10201 (N_10201,N_9348,N_8850);
nor U10202 (N_10202,N_9418,N_7960);
nand U10203 (N_10203,N_8741,N_9247);
or U10204 (N_10204,N_8196,N_8604);
and U10205 (N_10205,N_7715,N_8260);
and U10206 (N_10206,N_7630,N_9552);
nor U10207 (N_10207,N_8494,N_9204);
xnor U10208 (N_10208,N_9628,N_9235);
xor U10209 (N_10209,N_8772,N_9419);
nor U10210 (N_10210,N_8456,N_9508);
nor U10211 (N_10211,N_7955,N_7831);
nor U10212 (N_10212,N_9223,N_8206);
nand U10213 (N_10213,N_7694,N_9962);
nand U10214 (N_10214,N_9711,N_9913);
and U10215 (N_10215,N_9545,N_8990);
or U10216 (N_10216,N_8643,N_8665);
xnor U10217 (N_10217,N_9503,N_9147);
or U10218 (N_10218,N_9743,N_8997);
or U10219 (N_10219,N_7872,N_7875);
nand U10220 (N_10220,N_9364,N_8937);
and U10221 (N_10221,N_8976,N_8208);
xnor U10222 (N_10222,N_9309,N_9174);
nor U10223 (N_10223,N_8726,N_8952);
nor U10224 (N_10224,N_7508,N_8189);
nand U10225 (N_10225,N_9538,N_9679);
nand U10226 (N_10226,N_9594,N_8836);
nand U10227 (N_10227,N_8799,N_8186);
xnor U10228 (N_10228,N_7964,N_9667);
or U10229 (N_10229,N_7778,N_9253);
and U10230 (N_10230,N_8503,N_8448);
nand U10231 (N_10231,N_9185,N_7634);
or U10232 (N_10232,N_9484,N_8907);
nand U10233 (N_10233,N_8614,N_9380);
nor U10234 (N_10234,N_8539,N_9347);
or U10235 (N_10235,N_9413,N_9493);
or U10236 (N_10236,N_8184,N_8623);
or U10237 (N_10237,N_8298,N_9680);
xnor U10238 (N_10238,N_9156,N_8392);
and U10239 (N_10239,N_9120,N_7998);
xor U10240 (N_10240,N_9702,N_8251);
or U10241 (N_10241,N_7561,N_8528);
nand U10242 (N_10242,N_9810,N_7693);
and U10243 (N_10243,N_8594,N_9661);
xor U10244 (N_10244,N_8258,N_8483);
nor U10245 (N_10245,N_9002,N_8427);
xnor U10246 (N_10246,N_7868,N_9905);
or U10247 (N_10247,N_9920,N_8765);
or U10248 (N_10248,N_7880,N_7879);
and U10249 (N_10249,N_7907,N_9443);
or U10250 (N_10250,N_9030,N_7564);
nor U10251 (N_10251,N_8804,N_8699);
and U10252 (N_10252,N_9403,N_8355);
nand U10253 (N_10253,N_8996,N_9636);
xor U10254 (N_10254,N_8979,N_8080);
nand U10255 (N_10255,N_8283,N_8017);
xnor U10256 (N_10256,N_8304,N_7833);
nand U10257 (N_10257,N_7543,N_9793);
or U10258 (N_10258,N_8204,N_8477);
or U10259 (N_10259,N_9051,N_8540);
and U10260 (N_10260,N_9422,N_9395);
nor U10261 (N_10261,N_9698,N_9131);
nand U10262 (N_10262,N_8766,N_9294);
nor U10263 (N_10263,N_9142,N_9654);
xor U10264 (N_10264,N_7902,N_8405);
and U10265 (N_10265,N_9004,N_8972);
xnor U10266 (N_10266,N_7834,N_9585);
nor U10267 (N_10267,N_9626,N_7575);
nor U10268 (N_10268,N_8895,N_7672);
and U10269 (N_10269,N_9124,N_8861);
nand U10270 (N_10270,N_9455,N_9948);
xnor U10271 (N_10271,N_9213,N_8920);
nand U10272 (N_10272,N_9663,N_7524);
nor U10273 (N_10273,N_8089,N_9162);
nor U10274 (N_10274,N_9548,N_9408);
nand U10275 (N_10275,N_9320,N_8324);
nor U10276 (N_10276,N_9803,N_9496);
nor U10277 (N_10277,N_7503,N_9111);
nor U10278 (N_10278,N_9497,N_7887);
nand U10279 (N_10279,N_8312,N_9461);
nor U10280 (N_10280,N_7982,N_7592);
nand U10281 (N_10281,N_9219,N_7942);
and U10282 (N_10282,N_9724,N_8807);
or U10283 (N_10283,N_8144,N_7504);
nand U10284 (N_10284,N_8062,N_8071);
nand U10285 (N_10285,N_9889,N_8730);
and U10286 (N_10286,N_9179,N_8851);
xor U10287 (N_10287,N_8280,N_9532);
or U10288 (N_10288,N_9642,N_9352);
nor U10289 (N_10289,N_9099,N_9507);
or U10290 (N_10290,N_9912,N_9924);
nand U10291 (N_10291,N_8112,N_7699);
or U10292 (N_10292,N_8651,N_8367);
nand U10293 (N_10293,N_8532,N_9978);
or U10294 (N_10294,N_8295,N_9119);
xnor U10295 (N_10295,N_9960,N_8708);
xor U10296 (N_10296,N_9631,N_8941);
nand U10297 (N_10297,N_9955,N_7975);
nand U10298 (N_10298,N_9456,N_9163);
nor U10299 (N_10299,N_9445,N_9392);
and U10300 (N_10300,N_8359,N_7797);
nor U10301 (N_10301,N_7605,N_8079);
nor U10302 (N_10302,N_9557,N_7754);
nor U10303 (N_10303,N_8244,N_9580);
xnor U10304 (N_10304,N_8973,N_9362);
and U10305 (N_10305,N_8770,N_8628);
nor U10306 (N_10306,N_8669,N_9606);
nor U10307 (N_10307,N_9401,N_9259);
nor U10308 (N_10308,N_8193,N_7531);
nand U10309 (N_10309,N_7653,N_8823);
and U10310 (N_10310,N_8354,N_7802);
xor U10311 (N_10311,N_9533,N_7917);
nand U10312 (N_10312,N_7734,N_8117);
or U10313 (N_10313,N_8299,N_8019);
nor U10314 (N_10314,N_9467,N_9157);
nand U10315 (N_10315,N_8234,N_8390);
nand U10316 (N_10316,N_8223,N_8277);
xor U10317 (N_10317,N_7512,N_7821);
and U10318 (N_10318,N_8128,N_7517);
nand U10319 (N_10319,N_8710,N_7679);
nand U10320 (N_10320,N_8573,N_8182);
nand U10321 (N_10321,N_9399,N_8622);
or U10322 (N_10322,N_8660,N_9164);
nand U10323 (N_10323,N_7544,N_8009);
nor U10324 (N_10324,N_8101,N_8077);
or U10325 (N_10325,N_9313,N_8162);
nor U10326 (N_10326,N_8897,N_9397);
nand U10327 (N_10327,N_7757,N_8719);
xnor U10328 (N_10328,N_7676,N_9677);
xor U10329 (N_10329,N_8557,N_8523);
or U10330 (N_10330,N_7536,N_7684);
nor U10331 (N_10331,N_8102,N_8435);
nor U10332 (N_10332,N_9217,N_7692);
nand U10333 (N_10333,N_9078,N_9477);
or U10334 (N_10334,N_8357,N_8549);
xnor U10335 (N_10335,N_8440,N_8205);
xnor U10336 (N_10336,N_8522,N_9806);
xor U10337 (N_10337,N_7752,N_7871);
nor U10338 (N_10338,N_9214,N_8502);
nor U10339 (N_10339,N_9675,N_9263);
or U10340 (N_10340,N_8352,N_9114);
and U10341 (N_10341,N_7841,N_9285);
xor U10342 (N_10342,N_8602,N_9706);
or U10343 (N_10343,N_8130,N_7505);
and U10344 (N_10344,N_9243,N_9953);
xnor U10345 (N_10345,N_8238,N_9820);
and U10346 (N_10346,N_9539,N_9509);
or U10347 (N_10347,N_9760,N_8300);
and U10348 (N_10348,N_8122,N_7941);
and U10349 (N_10349,N_8228,N_8404);
nand U10350 (N_10350,N_8743,N_7905);
and U10351 (N_10351,N_7869,N_9514);
xor U10352 (N_10352,N_8350,N_9697);
nand U10353 (N_10353,N_8744,N_7611);
or U10354 (N_10354,N_8899,N_7874);
and U10355 (N_10355,N_9554,N_7696);
and U10356 (N_10356,N_8649,N_9482);
xnor U10357 (N_10357,N_8659,N_8625);
nand U10358 (N_10358,N_9704,N_8385);
xnor U10359 (N_10359,N_9023,N_7703);
and U10360 (N_10360,N_8338,N_7713);
nor U10361 (N_10361,N_8029,N_8365);
and U10362 (N_10362,N_7791,N_8034);
xnor U10363 (N_10363,N_7726,N_7851);
xnor U10364 (N_10364,N_8510,N_8425);
and U10365 (N_10365,N_9678,N_7645);
or U10366 (N_10366,N_8248,N_7999);
nand U10367 (N_10367,N_7966,N_9512);
and U10368 (N_10368,N_8983,N_9178);
nor U10369 (N_10369,N_8853,N_9956);
nand U10370 (N_10370,N_7521,N_8007);
xor U10371 (N_10371,N_9805,N_8466);
and U10372 (N_10372,N_8005,N_8060);
xnor U10373 (N_10373,N_9317,N_8509);
or U10374 (N_10374,N_7706,N_9809);
nor U10375 (N_10375,N_9042,N_8358);
nor U10376 (N_10376,N_9389,N_8814);
or U10377 (N_10377,N_8749,N_9616);
nand U10378 (N_10378,N_9316,N_9404);
nor U10379 (N_10379,N_7628,N_8512);
nand U10380 (N_10380,N_9121,N_8645);
nand U10381 (N_10381,N_7820,N_9020);
nor U10382 (N_10382,N_9175,N_9037);
nand U10383 (N_10383,N_8597,N_7601);
and U10384 (N_10384,N_9279,N_8798);
xor U10385 (N_10385,N_8747,N_9077);
xor U10386 (N_10386,N_8585,N_9006);
nand U10387 (N_10387,N_9570,N_8558);
nor U10388 (N_10388,N_9495,N_8098);
nand U10389 (N_10389,N_7944,N_8679);
xnor U10390 (N_10390,N_7812,N_9645);
nor U10391 (N_10391,N_8986,N_8561);
xor U10392 (N_10392,N_9357,N_9227);
nor U10393 (N_10393,N_8800,N_8786);
and U10394 (N_10394,N_9750,N_8316);
and U10395 (N_10395,N_9751,N_9981);
nor U10396 (N_10396,N_8762,N_8341);
and U10397 (N_10397,N_8090,N_8905);
xor U10398 (N_10398,N_9018,N_8458);
nor U10399 (N_10399,N_7864,N_8025);
nor U10400 (N_10400,N_9080,N_9321);
and U10401 (N_10401,N_8866,N_8524);
nor U10402 (N_10402,N_9877,N_8105);
and U10403 (N_10403,N_9815,N_9346);
xor U10404 (N_10404,N_9513,N_9879);
and U10405 (N_10405,N_9526,N_9470);
xnor U10406 (N_10406,N_8391,N_7641);
and U10407 (N_10407,N_9531,N_9264);
and U10408 (N_10408,N_9014,N_9886);
or U10409 (N_10409,N_8406,N_8369);
nor U10410 (N_10410,N_9910,N_9468);
or U10411 (N_10411,N_8261,N_8621);
or U10412 (N_10412,N_7923,N_9885);
nand U10413 (N_10413,N_7756,N_7948);
xnor U10414 (N_10414,N_8801,N_9351);
and U10415 (N_10415,N_9181,N_9900);
nor U10416 (N_10416,N_9907,N_9571);
nand U10417 (N_10417,N_8279,N_8545);
nor U10418 (N_10418,N_8777,N_8187);
nor U10419 (N_10419,N_8450,N_8701);
xnor U10420 (N_10420,N_8241,N_8307);
or U10421 (N_10421,N_7994,N_7938);
or U10422 (N_10422,N_8046,N_9719);
nor U10423 (N_10423,N_8879,N_9058);
and U10424 (N_10424,N_7903,N_7965);
nand U10425 (N_10425,N_8774,N_9377);
or U10426 (N_10426,N_9444,N_9336);
nor U10427 (N_10427,N_9757,N_9699);
xnor U10428 (N_10428,N_7652,N_9904);
nor U10429 (N_10429,N_9365,N_9031);
xor U10430 (N_10430,N_8608,N_8981);
nor U10431 (N_10431,N_7988,N_9641);
and U10432 (N_10432,N_8235,N_7732);
nand U10433 (N_10433,N_7983,N_8377);
or U10434 (N_10434,N_7958,N_8890);
nand U10435 (N_10435,N_8548,N_9036);
and U10436 (N_10436,N_8827,N_7571);
nor U10437 (N_10437,N_9433,N_9427);
and U10438 (N_10438,N_8886,N_9094);
and U10439 (N_10439,N_8321,N_8978);
or U10440 (N_10440,N_9123,N_7515);
and U10441 (N_10441,N_7893,N_8846);
or U10442 (N_10442,N_9278,N_8344);
xor U10443 (N_10443,N_7976,N_8936);
or U10444 (N_10444,N_7621,N_9231);
nor U10445 (N_10445,N_9472,N_8992);
xor U10446 (N_10446,N_9598,N_9055);
nand U10447 (N_10447,N_7691,N_9746);
and U10448 (N_10448,N_9200,N_9619);
and U10449 (N_10449,N_9478,N_9435);
or U10450 (N_10450,N_9372,N_7658);
and U10451 (N_10451,N_8308,N_8278);
nor U10452 (N_10452,N_9965,N_9767);
or U10453 (N_10453,N_9341,N_9858);
nand U10454 (N_10454,N_9085,N_8460);
nor U10455 (N_10455,N_8286,N_9402);
xnor U10456 (N_10456,N_8757,N_8644);
nand U10457 (N_10457,N_7720,N_9414);
nand U10458 (N_10458,N_8925,N_8428);
nand U10459 (N_10459,N_8065,N_7908);
and U10460 (N_10460,N_9583,N_8370);
or U10461 (N_10461,N_9605,N_9916);
nand U10462 (N_10462,N_7638,N_9190);
and U10463 (N_10463,N_8158,N_9536);
and U10464 (N_10464,N_9966,N_8264);
and U10465 (N_10465,N_8928,N_7814);
nor U10466 (N_10466,N_9485,N_9136);
nor U10467 (N_10467,N_9098,N_7950);
or U10468 (N_10468,N_8720,N_9745);
or U10469 (N_10469,N_8403,N_8697);
xor U10470 (N_10470,N_9975,N_8790);
nor U10471 (N_10471,N_9171,N_7827);
xor U10472 (N_10472,N_7502,N_8724);
xnor U10473 (N_10473,N_7766,N_8220);
nand U10474 (N_10474,N_7935,N_7928);
or U10475 (N_10475,N_7771,N_8753);
xor U10476 (N_10476,N_7795,N_7578);
nor U10477 (N_10477,N_7547,N_8654);
xor U10478 (N_10478,N_8942,N_7668);
nor U10479 (N_10479,N_8837,N_8672);
or U10480 (N_10480,N_9774,N_9198);
nor U10481 (N_10481,N_8256,N_8455);
or U10482 (N_10482,N_9941,N_7811);
or U10483 (N_10483,N_7816,N_8212);
xor U10484 (N_10484,N_8500,N_8104);
xnor U10485 (N_10485,N_7995,N_9244);
xor U10486 (N_10486,N_8233,N_8078);
nand U10487 (N_10487,N_8530,N_9836);
nor U10488 (N_10488,N_7642,N_9854);
nand U10489 (N_10489,N_8121,N_9499);
xnor U10490 (N_10490,N_8191,N_9782);
or U10491 (N_10491,N_8632,N_9562);
or U10492 (N_10492,N_8525,N_8434);
or U10493 (N_10493,N_9744,N_8430);
and U10494 (N_10494,N_8068,N_9596);
or U10495 (N_10495,N_8432,N_8167);
or U10496 (N_10496,N_8081,N_9450);
xor U10497 (N_10497,N_7612,N_8115);
xor U10498 (N_10498,N_9280,N_7763);
nor U10499 (N_10499,N_9384,N_9601);
nand U10500 (N_10500,N_8779,N_8271);
nor U10501 (N_10501,N_8422,N_9262);
or U10502 (N_10502,N_7662,N_7589);
nand U10503 (N_10503,N_8975,N_9130);
nor U10504 (N_10504,N_9892,N_9242);
xnor U10505 (N_10505,N_9225,N_8215);
xor U10506 (N_10506,N_8253,N_9935);
nor U10507 (N_10507,N_8763,N_9992);
nor U10508 (N_10508,N_8366,N_7644);
nand U10509 (N_10509,N_9252,N_9694);
xnor U10510 (N_10510,N_7729,N_7610);
or U10511 (N_10511,N_9049,N_7937);
nand U10512 (N_10512,N_8663,N_9909);
nand U10513 (N_10513,N_8473,N_8454);
or U10514 (N_10514,N_8929,N_9066);
nor U10515 (N_10515,N_9883,N_9074);
or U10516 (N_10516,N_8066,N_9771);
nor U10517 (N_10517,N_8647,N_9340);
or U10518 (N_10518,N_9224,N_8916);
nor U10519 (N_10519,N_9096,N_8199);
or U10520 (N_10520,N_8465,N_8791);
and U10521 (N_10521,N_9627,N_8265);
and U10522 (N_10522,N_9823,N_8227);
xnor U10523 (N_10523,N_9211,N_8601);
xnor U10524 (N_10524,N_7741,N_8671);
and U10525 (N_10525,N_8735,N_8302);
nor U10526 (N_10526,N_8578,N_8495);
xnor U10527 (N_10527,N_9818,N_7739);
nor U10528 (N_10528,N_9166,N_8259);
xnor U10529 (N_10529,N_9893,N_9060);
nand U10530 (N_10530,N_8805,N_8041);
xnor U10531 (N_10531,N_9481,N_8926);
xnor U10532 (N_10532,N_9759,N_8857);
and U10533 (N_10533,N_9453,N_9684);
and U10534 (N_10534,N_9083,N_7532);
nor U10535 (N_10535,N_9376,N_7507);
xor U10536 (N_10536,N_9015,N_9637);
xor U10537 (N_10537,N_8811,N_9592);
xnor U10538 (N_10538,N_7946,N_9674);
nor U10539 (N_10539,N_8813,N_9959);
or U10540 (N_10540,N_7620,N_9696);
nand U10541 (N_10541,N_7702,N_9928);
nor U10542 (N_10542,N_7514,N_8619);
nor U10543 (N_10543,N_7563,N_9091);
and U10544 (N_10544,N_9984,N_9890);
nor U10545 (N_10545,N_7603,N_9617);
or U10546 (N_10546,N_9970,N_8297);
and U10547 (N_10547,N_9202,N_9068);
xor U10548 (N_10548,N_8797,N_7697);
xnor U10549 (N_10549,N_8911,N_8408);
and U10550 (N_10550,N_8581,N_9286);
or U10551 (N_10551,N_7751,N_8734);
xor U10552 (N_10552,N_8210,N_9868);
nand U10553 (N_10553,N_8436,N_8412);
or U10554 (N_10554,N_9822,N_8070);
nor U10555 (N_10555,N_9804,N_9707);
nor U10556 (N_10556,N_7956,N_8372);
nand U10557 (N_10557,N_9172,N_8496);
or U10558 (N_10558,N_9375,N_9095);
nand U10559 (N_10559,N_7783,N_8411);
nand U10560 (N_10560,N_9260,N_9167);
nand U10561 (N_10561,N_9833,N_8076);
and U10562 (N_10562,N_9614,N_8882);
or U10563 (N_10563,N_8667,N_7992);
nand U10564 (N_10564,N_8159,N_8793);
and U10565 (N_10565,N_8775,N_8351);
nand U10566 (N_10566,N_8010,N_7542);
and U10567 (N_10567,N_8072,N_8867);
xnor U10568 (N_10568,N_9520,N_8064);
or U10569 (N_10569,N_8787,N_7718);
xor U10570 (N_10570,N_7643,N_8519);
or U10571 (N_10571,N_9097,N_9329);
and U10572 (N_10572,N_9476,N_9090);
nor U10573 (N_10573,N_9929,N_9491);
nor U10574 (N_10574,N_7598,N_8361);
or U10575 (N_10575,N_8231,N_8142);
nor U10576 (N_10576,N_9016,N_7636);
or U10577 (N_10577,N_9811,N_8035);
and U10578 (N_10578,N_7913,N_7892);
nand U10579 (N_10579,N_7623,N_8839);
or U10580 (N_10580,N_8429,N_9417);
nand U10581 (N_10581,N_7671,N_9480);
nor U10582 (N_10582,N_9576,N_9440);
nor U10583 (N_10583,N_8764,N_7538);
nor U10584 (N_10584,N_8551,N_8040);
nor U10585 (N_10585,N_8803,N_8249);
xnor U10586 (N_10586,N_9951,N_9407);
nor U10587 (N_10587,N_8097,N_8655);
nand U10588 (N_10588,N_8707,N_7704);
and U10589 (N_10589,N_9432,N_8008);
nand U10590 (N_10590,N_9199,N_8451);
or U10591 (N_10591,N_9337,N_8795);
or U10592 (N_10592,N_8333,N_9160);
nor U10593 (N_10593,N_7654,N_8164);
nand U10594 (N_10594,N_9950,N_8379);
nor U10595 (N_10595,N_9690,N_9150);
xnor U10596 (N_10596,N_8785,N_8301);
nor U10597 (N_10597,N_8816,N_8133);
and U10598 (N_10598,N_8310,N_9611);
nand U10599 (N_10599,N_9203,N_8371);
or U10600 (N_10600,N_9448,N_7953);
nor U10601 (N_10601,N_8021,N_8930);
and U10602 (N_10602,N_7910,N_8011);
and U10603 (N_10603,N_9250,N_8705);
nor U10604 (N_10604,N_9990,N_9986);
nand U10605 (N_10605,N_7534,N_9284);
xnor U10606 (N_10606,N_7583,N_9768);
nor U10607 (N_10607,N_8513,N_7573);
xor U10608 (N_10608,N_8444,N_8148);
and U10609 (N_10609,N_7877,N_7609);
nor U10610 (N_10610,N_7527,N_8095);
nor U10611 (N_10611,N_8702,N_9245);
xnor U10612 (N_10612,N_9729,N_9424);
xor U10613 (N_10613,N_9855,N_8170);
nand U10614 (N_10614,N_8751,N_8155);
and U10615 (N_10615,N_8686,N_8544);
or U10616 (N_10616,N_8447,N_8939);
xnor U10617 (N_10617,N_7667,N_8272);
or U10618 (N_10618,N_7683,N_7977);
xnor U10619 (N_10619,N_7931,N_8881);
and U10620 (N_10620,N_7943,N_7862);
or U10621 (N_10621,N_8844,N_9560);
and U10622 (N_10622,N_8588,N_9834);
nand U10623 (N_10623,N_9088,N_8918);
or U10624 (N_10624,N_9723,N_9127);
nand U10625 (N_10625,N_8282,N_9011);
and U10626 (N_10626,N_9731,N_8474);
nand U10627 (N_10627,N_8693,N_8437);
nor U10628 (N_10628,N_9379,N_8536);
and U10629 (N_10629,N_9938,N_9994);
nand U10630 (N_10630,N_9039,N_7570);
nor U10631 (N_10631,N_8047,N_9299);
nand U10632 (N_10632,N_9076,N_9035);
or U10633 (N_10633,N_9047,N_7614);
and U10634 (N_10634,N_8103,N_9210);
xnor U10635 (N_10635,N_8414,N_8521);
nand U10636 (N_10636,N_7989,N_8303);
nor U10637 (N_10637,N_9501,N_7730);
nand U10638 (N_10638,N_9038,N_7922);
xnor U10639 (N_10639,N_9550,N_8467);
xnor U10640 (N_10640,N_9932,N_9549);
nor U10641 (N_10641,N_8479,N_9814);
nor U10642 (N_10642,N_8778,N_7829);
nand U10643 (N_10643,N_9777,N_8889);
xnor U10644 (N_10644,N_9473,N_9911);
nor U10645 (N_10645,N_7824,N_8190);
and U10646 (N_10646,N_8865,N_9783);
nand U10647 (N_10647,N_9563,N_8598);
nand U10648 (N_10648,N_9808,N_9860);
nor U10649 (N_10649,N_8111,N_9736);
or U10650 (N_10650,N_8974,N_8874);
or U10651 (N_10651,N_8615,N_8533);
nor U10652 (N_10652,N_8309,N_7545);
xor U10653 (N_10653,N_9487,N_7954);
xnor U10654 (N_10654,N_8684,N_9233);
and U10655 (N_10655,N_8349,N_9000);
xor U10656 (N_10656,N_9367,N_8739);
nand U10657 (N_10657,N_7796,N_9360);
xor U10658 (N_10658,N_9590,N_8653);
and U10659 (N_10659,N_8482,N_7593);
nor U10660 (N_10660,N_8059,N_8817);
or U10661 (N_10661,N_9061,N_9439);
nand U10662 (N_10662,N_8737,N_8131);
xor U10663 (N_10663,N_8114,N_8893);
and U10664 (N_10664,N_7580,N_9490);
nand U10665 (N_10665,N_8784,N_8901);
xor U10666 (N_10666,N_7526,N_9269);
or U10667 (N_10667,N_8792,N_8988);
xnor U10668 (N_10668,N_9721,N_8092);
nand U10669 (N_10669,N_9780,N_9573);
and U10670 (N_10670,N_8746,N_9143);
or U10671 (N_10671,N_7674,N_8562);
xor U10672 (N_10672,N_8571,N_7535);
nand U10673 (N_10673,N_9134,N_8472);
nand U10674 (N_10674,N_9765,N_9438);
and U10675 (N_10675,N_9991,N_9149);
nor U10676 (N_10676,N_8449,N_9064);
nor U10677 (N_10677,N_8685,N_9686);
or U10678 (N_10678,N_9333,N_9682);
or U10679 (N_10679,N_8670,N_9282);
and U10680 (N_10680,N_9498,N_7742);
nand U10681 (N_10681,N_8383,N_9753);
nand U10682 (N_10682,N_9007,N_8195);
or U10683 (N_10683,N_8330,N_9383);
xnor U10684 (N_10684,N_8727,N_9492);
xnor U10685 (N_10685,N_8683,N_8736);
xnor U10686 (N_10686,N_9927,N_7633);
and U10687 (N_10687,N_8023,N_7894);
and U10688 (N_10688,N_9165,N_9145);
or U10689 (N_10689,N_9169,N_9624);
or U10690 (N_10690,N_9516,N_7585);
nor U10691 (N_10691,N_8568,N_8376);
and U10692 (N_10692,N_7830,N_9701);
and U10693 (N_10693,N_8630,N_7897);
or U10694 (N_10694,N_9668,N_8387);
xor U10695 (N_10695,N_8415,N_9366);
or U10696 (N_10696,N_9716,N_8587);
nand U10697 (N_10697,N_7767,N_9342);
nor U10698 (N_10698,N_9817,N_8830);
and U10699 (N_10699,N_9870,N_8994);
and U10700 (N_10700,N_9196,N_9325);
nor U10701 (N_10701,N_8904,N_8529);
or U10702 (N_10702,N_7823,N_7608);
xor U10703 (N_10703,N_8020,N_9005);
nand U10704 (N_10704,N_7838,N_8965);
xor U10705 (N_10705,N_9862,N_7568);
nand U10706 (N_10706,N_9515,N_8318);
nand U10707 (N_10707,N_8314,N_8055);
xnor U10708 (N_10708,N_8694,N_8825);
nor U10709 (N_10709,N_7776,N_7622);
nand U10710 (N_10710,N_8145,N_8954);
nand U10711 (N_10711,N_8620,N_7606);
nand U10712 (N_10712,N_8048,N_7785);
and U10713 (N_10713,N_8242,N_8407);
and U10714 (N_10714,N_9071,N_8960);
or U10715 (N_10715,N_9323,N_8342);
and U10716 (N_10716,N_7567,N_9228);
nor U10717 (N_10717,N_7690,N_9173);
nand U10718 (N_10718,N_8399,N_7688);
xnor U10719 (N_10719,N_9713,N_9201);
nand U10720 (N_10720,N_9287,N_7651);
xor U10721 (N_10721,N_8553,N_9649);
nand U10722 (N_10722,N_8031,N_9521);
nor U10723 (N_10723,N_7770,N_8675);
and U10724 (N_10724,N_9968,N_7613);
and U10725 (N_10725,N_8284,N_9261);
xnor U10726 (N_10726,N_9857,N_9758);
nand U10727 (N_10727,N_8709,N_9620);
and U10728 (N_10728,N_8721,N_9838);
nor U10729 (N_10729,N_7682,N_8197);
and U10730 (N_10730,N_8740,N_9853);
and U10731 (N_10731,N_9591,N_7509);
xnor U10732 (N_10732,N_8690,N_9676);
xor U10733 (N_10733,N_7768,N_8603);
and U10734 (N_10734,N_9599,N_7660);
or U10735 (N_10735,N_9584,N_9393);
nor U10736 (N_10736,N_8381,N_9052);
xor U10737 (N_10737,N_9300,N_9302);
or U10738 (N_10738,N_9623,N_8075);
nor U10739 (N_10739,N_9449,N_9381);
and U10740 (N_10740,N_9084,N_9979);
nand U10741 (N_10741,N_8229,N_8860);
or U10742 (N_10742,N_7717,N_9092);
or U10743 (N_10743,N_9934,N_9288);
nor U10744 (N_10744,N_7970,N_9873);
nand U10745 (N_10745,N_7860,N_8535);
nor U10746 (N_10746,N_9603,N_9115);
or U10747 (N_10747,N_8421,N_9138);
and U10748 (N_10748,N_7670,N_8695);
and U10749 (N_10749,N_9483,N_8232);
xnor U10750 (N_10750,N_8638,N_8656);
or U10751 (N_10751,N_8841,N_9462);
and U10752 (N_10752,N_8582,N_9812);
or U10753 (N_10753,N_9102,N_8153);
nand U10754 (N_10754,N_8480,N_8364);
nand U10755 (N_10755,N_8030,N_8401);
nor U10756 (N_10756,N_9338,N_8345);
or U10757 (N_10757,N_9266,N_8113);
or U10758 (N_10758,N_7743,N_9327);
or U10759 (N_10759,N_8878,N_9957);
or U10760 (N_10760,N_7845,N_9176);
and U10761 (N_10761,N_8910,N_7728);
and U10762 (N_10762,N_9671,N_9307);
and U10763 (N_10763,N_9028,N_9589);
or U10764 (N_10764,N_9265,N_9019);
xnor U10765 (N_10765,N_7837,N_8900);
or U10766 (N_10766,N_8294,N_9275);
and U10767 (N_10767,N_9825,N_9906);
and U10768 (N_10768,N_8137,N_7974);
and U10769 (N_10769,N_9001,N_9876);
and U10770 (N_10770,N_7579,N_9971);
xor U10771 (N_10771,N_9270,N_7708);
xnor U10772 (N_10772,N_9535,N_7656);
or U10773 (N_10773,N_7695,N_8054);
nor U10774 (N_10774,N_9423,N_8738);
or U10775 (N_10775,N_8168,N_7576);
xor U10776 (N_10776,N_9525,N_8612);
xnor U10777 (N_10777,N_8373,N_9931);
or U10778 (N_10778,N_7772,N_8591);
and U10779 (N_10779,N_9856,N_8488);
nand U10780 (N_10780,N_9875,N_8934);
or U10781 (N_10781,N_9662,N_7936);
and U10782 (N_10782,N_9012,N_8717);
xnor U10783 (N_10783,N_9140,N_8580);
or U10784 (N_10784,N_7828,N_7640);
or U10785 (N_10785,N_8446,N_8732);
nor U10786 (N_10786,N_8149,N_7719);
xnor U10787 (N_10787,N_8552,N_7817);
or U10788 (N_10788,N_8053,N_7721);
nor U10789 (N_10789,N_8374,N_8896);
nor U10790 (N_10790,N_9849,N_9577);
or U10791 (N_10791,N_8292,N_8914);
nand U10792 (N_10792,N_8963,N_9410);
nand U10793 (N_10793,N_9452,N_8877);
nor U10794 (N_10794,N_8863,N_8420);
and U10795 (N_10795,N_8218,N_7866);
nor U10796 (N_10796,N_8443,N_8050);
nand U10797 (N_10797,N_9304,N_8217);
or U10798 (N_10798,N_8818,N_8382);
xor U10799 (N_10799,N_8291,N_7528);
xor U10800 (N_10800,N_9194,N_8894);
xor U10801 (N_10801,N_8969,N_8485);
and U10802 (N_10802,N_9505,N_8439);
nor U10803 (N_10803,N_9778,N_9153);
or U10804 (N_10804,N_7804,N_8516);
or U10805 (N_10805,N_9232,N_8004);
and U10806 (N_10806,N_9297,N_9961);
nand U10807 (N_10807,N_8207,N_9246);
or U10808 (N_10808,N_9930,N_8849);
xnor U10809 (N_10809,N_8484,N_9987);
nand U10810 (N_10810,N_9355,N_7552);
or U10811 (N_10811,N_9918,N_7789);
nor U10812 (N_10812,N_8962,N_7786);
xnor U10813 (N_10813,N_9065,N_8254);
xnor U10814 (N_10814,N_8933,N_7895);
nor U10815 (N_10815,N_8783,N_7858);
and U10816 (N_10816,N_8213,N_7557);
nand U10817 (N_10817,N_7873,N_8674);
or U10818 (N_10818,N_7882,N_9692);
and U10819 (N_10819,N_9625,N_9795);
nor U10820 (N_10820,N_8982,N_9465);
nor U10821 (N_10821,N_8266,N_9788);
and U10822 (N_10822,N_7506,N_9008);
nor U10823 (N_10823,N_7899,N_8636);
nand U10824 (N_10824,N_7760,N_9050);
xor U10825 (N_10825,N_9949,N_8756);
nor U10826 (N_10826,N_8518,N_8118);
nand U10827 (N_10827,N_9056,N_7727);
nand U10828 (N_10828,N_8635,N_8634);
nor U10829 (N_10829,N_8486,N_7673);
xor U10830 (N_10830,N_8641,N_9353);
or U10831 (N_10831,N_7516,N_7890);
or U10832 (N_10832,N_9222,N_8067);
and U10833 (N_10833,N_9952,N_9865);
nand U10834 (N_10834,N_7669,N_8000);
nor U10835 (N_10835,N_7758,N_9914);
xor U10836 (N_10836,N_8820,N_9195);
and U10837 (N_10837,N_9648,N_9973);
xnor U10838 (N_10838,N_9844,N_9426);
nor U10839 (N_10839,N_9615,N_8611);
and U10840 (N_10840,N_9728,N_8862);
nor U10841 (N_10841,N_8091,N_7973);
and U10842 (N_10842,N_7689,N_8869);
or U10843 (N_10843,N_7784,N_8531);
and U10844 (N_10844,N_8088,N_8953);
nor U10845 (N_10845,N_9062,N_8613);
nand U10846 (N_10846,N_8269,N_8661);
nand U10847 (N_10847,N_9660,N_8174);
and U10848 (N_10848,N_8058,N_8129);
and U10849 (N_10849,N_8802,N_8397);
or U10850 (N_10850,N_9144,N_9556);
nand U10851 (N_10851,N_9540,N_8028);
xor U10852 (N_10852,N_9412,N_9363);
xnor U10853 (N_10853,N_8989,N_9574);
xnor U10854 (N_10854,N_7967,N_9330);
and U10855 (N_10855,N_8875,N_9789);
nor U10856 (N_10856,N_8833,N_8538);
nand U10857 (N_10857,N_8384,N_9983);
or U10858 (N_10858,N_9896,N_7876);
nor U10859 (N_10859,N_9197,N_7780);
and U10860 (N_10860,N_9369,N_7808);
nand U10861 (N_10861,N_8723,N_7712);
nor U10862 (N_10862,N_7513,N_9296);
xor U10863 (N_10863,N_8099,N_8824);
or U10864 (N_10864,N_8108,N_8156);
and U10865 (N_10865,N_8788,N_8662);
nor U10866 (N_10866,N_9273,N_8526);
nor U10867 (N_10867,N_8505,N_9133);
nor U10868 (N_10868,N_8838,N_8650);
nor U10869 (N_10869,N_9954,N_9718);
and U10870 (N_10870,N_9846,N_9209);
or U10871 (N_10871,N_7537,N_8332);
nor U10872 (N_10872,N_7906,N_8574);
nor U10873 (N_10873,N_8178,N_9755);
and U10874 (N_10874,N_7745,N_8453);
and U10875 (N_10875,N_8812,N_9283);
nand U10876 (N_10876,N_9378,N_7809);
nor U10877 (N_10877,N_9459,N_9193);
xor U10878 (N_10878,N_9848,N_7574);
xnor U10879 (N_10879,N_8325,N_7725);
xnor U10880 (N_10880,N_8599,N_8250);
and U10881 (N_10881,N_7749,N_9903);
nand U10882 (N_10882,N_8593,N_9180);
xnor U10883 (N_10883,N_8959,N_9575);
or U10884 (N_10884,N_8052,N_9864);
xor U10885 (N_10885,N_9587,N_9434);
xor U10886 (N_10886,N_8808,N_9710);
nor U10887 (N_10887,N_8700,N_9722);
and U10888 (N_10888,N_9613,N_7556);
nor U10889 (N_10889,N_8056,N_9874);
nor U10890 (N_10890,N_9936,N_7590);
and U10891 (N_10891,N_8609,N_7951);
and U10892 (N_10892,N_8380,N_8109);
xor U10893 (N_10893,N_9128,N_9995);
nand U10894 (N_10894,N_7551,N_9715);
nor U10895 (N_10895,N_8748,N_9048);
or U10896 (N_10896,N_7949,N_8475);
nand U10897 (N_10897,N_8534,N_8003);
and U10898 (N_10898,N_8586,N_7959);
nor U10899 (N_10899,N_8224,N_8245);
nor U10900 (N_10900,N_9943,N_9813);
or U10901 (N_10901,N_9212,N_9737);
xnor U10902 (N_10902,N_8039,N_8537);
and U10903 (N_10903,N_9632,N_9887);
xnor U10904 (N_10904,N_7616,N_9093);
nand U10905 (N_10905,N_7854,N_9475);
nand U10906 (N_10906,N_7501,N_8083);
nand U10907 (N_10907,N_9441,N_9335);
nor U10908 (N_10908,N_8515,N_7968);
and U10909 (N_10909,N_9542,N_9635);
xnor U10910 (N_10910,N_9045,N_8718);
nor U10911 (N_10911,N_9884,N_8074);
nor U10912 (N_10912,N_9471,N_8759);
and U10913 (N_10913,N_8147,N_7626);
xnor U10914 (N_10914,N_7666,N_7519);
nand U10915 (N_10915,N_8257,N_8402);
nor U10916 (N_10916,N_8637,N_9688);
or U10917 (N_10917,N_9277,N_9888);
xor U10918 (N_10918,N_9670,N_8995);
and U10919 (N_10919,N_9872,N_8476);
nand U10920 (N_10920,N_8487,N_8570);
nor U10921 (N_10921,N_8501,N_9639);
or U10922 (N_10922,N_8154,N_8348);
or U10923 (N_10923,N_9184,N_8424);
xnor U10924 (N_10924,N_8715,N_8471);
nand U10925 (N_10925,N_9437,N_8794);
nand U10926 (N_10926,N_8395,N_8082);
nand U10927 (N_10927,N_8329,N_9447);
nor U10928 (N_10928,N_9653,N_9226);
and U10929 (N_10929,N_8416,N_7985);
nand U10930 (N_10930,N_8273,N_8835);
xnor U10931 (N_10931,N_7861,N_9319);
nand U10932 (N_10932,N_8565,N_7748);
xnor U10933 (N_10933,N_9370,N_7806);
nand U10934 (N_10934,N_8413,N_9530);
nand U10935 (N_10935,N_8498,N_8438);
or U10936 (N_10936,N_8051,N_8546);
xor U10937 (N_10937,N_8305,N_9769);
nor U10938 (N_10938,N_9234,N_8511);
and U10939 (N_10939,N_8923,N_8713);
nor U10940 (N_10940,N_9565,N_8796);
and U10941 (N_10941,N_7607,N_8560);
nand U10942 (N_10942,N_7825,N_8014);
xor U10943 (N_10943,N_9996,N_9354);
and U10944 (N_10944,N_9831,N_9775);
nor U10945 (N_10945,N_9146,N_9824);
xnor U10946 (N_10946,N_9044,N_7835);
xnor U10947 (N_10947,N_8610,N_8086);
nand U10948 (N_10948,N_8036,N_7900);
nand U10949 (N_10949,N_8698,N_8648);
nand U10950 (N_10950,N_9776,N_8132);
nand U10951 (N_10951,N_9784,N_7555);
xnor U10952 (N_10952,N_9494,N_9216);
nand U10953 (N_10953,N_9863,N_7912);
xnor U10954 (N_10954,N_7646,N_8729);
and U10955 (N_10955,N_7800,N_9308);
xnor U10956 (N_10956,N_9604,N_8172);
and U10957 (N_10957,N_9248,N_7915);
or U10958 (N_10958,N_9830,N_9236);
nand U10959 (N_10959,N_8462,N_9638);
xnor U10960 (N_10960,N_8311,N_8955);
and U10961 (N_10961,N_8781,N_9189);
and U10962 (N_10962,N_9902,N_9845);
xnor U10963 (N_10963,N_9633,N_9976);
and U10964 (N_10964,N_9572,N_9141);
nor U10965 (N_10965,N_9524,N_7774);
nand U10966 (N_10966,N_9643,N_9733);
nor U10967 (N_10967,N_9691,N_9469);
or U10968 (N_10968,N_9135,N_7522);
nand U10969 (N_10969,N_7649,N_9409);
and U10970 (N_10970,N_9786,N_9894);
xnor U10971 (N_10971,N_9528,N_9155);
nand U10972 (N_10972,N_9708,N_8950);
and U10973 (N_10973,N_9618,N_9829);
or U10974 (N_10974,N_8555,N_7993);
or U10975 (N_10975,N_9229,N_9415);
nand U10976 (N_10976,N_8589,N_7657);
or U10977 (N_10977,N_7832,N_9843);
nor U10978 (N_10978,N_7569,N_9400);
nor U10979 (N_10979,N_9821,N_9559);
xor U10980 (N_10980,N_9255,N_9137);
nand U10981 (N_10981,N_8868,N_8293);
nand U10982 (N_10982,N_9807,N_9607);
nor U10983 (N_10983,N_9312,N_9522);
xnor U10984 (N_10984,N_8141,N_9740);
nand U10985 (N_10985,N_9850,N_9752);
or U10986 (N_10986,N_7803,N_7934);
xnor U10987 (N_10987,N_7963,N_8107);
xnor U10988 (N_10988,N_8268,N_8507);
or U10989 (N_10989,N_9186,N_7685);
and U10990 (N_10990,N_8287,N_8127);
nand U10991 (N_10991,N_9891,N_9683);
xor U10992 (N_10992,N_7847,N_7661);
nand U10993 (N_10993,N_8022,N_8666);
or U10994 (N_10994,N_9027,N_9739);
nor U10995 (N_10995,N_7602,N_9534);
or U10996 (N_10996,N_7952,N_8236);
or U10997 (N_10997,N_9734,N_8262);
and U10998 (N_10998,N_8057,N_9839);
nand U10999 (N_10999,N_8980,N_9866);
or U11000 (N_11000,N_7759,N_9289);
or U11001 (N_11001,N_8135,N_8126);
xor U11002 (N_11002,N_9946,N_8617);
nand U11003 (N_11003,N_8843,N_8871);
or U11004 (N_11004,N_8922,N_9182);
nor U11005 (N_11005,N_8564,N_9537);
and U11006 (N_11006,N_8964,N_8032);
nand U11007 (N_11007,N_8913,N_8542);
xor U11008 (N_11008,N_9646,N_9152);
or U11009 (N_11009,N_9980,N_8616);
xor U11010 (N_11010,N_8417,N_7530);
nor U11011 (N_11011,N_7686,N_9371);
nor U11012 (N_11012,N_7765,N_7591);
nand U11013 (N_11013,N_7553,N_9551);
nand U11014 (N_11014,N_9799,N_7793);
or U11015 (N_11015,N_8431,N_8583);
or U11016 (N_11016,N_9281,N_8353);
or U11017 (N_11017,N_8493,N_9964);
xnor U11018 (N_11018,N_8831,N_9398);
and U11019 (N_11019,N_7798,N_9658);
nand U11020 (N_11020,N_7546,N_8198);
xnor U11021 (N_11021,N_9835,N_9334);
and U11022 (N_11022,N_8633,N_7740);
nor U11023 (N_11023,N_7822,N_9908);
nor U11024 (N_11024,N_8750,N_7577);
xnor U11025 (N_11025,N_9271,N_9926);
nand U11026 (N_11026,N_8706,N_8940);
or U11027 (N_11027,N_7687,N_7635);
nor U11028 (N_11028,N_7597,N_8181);
nor U11029 (N_11029,N_8576,N_9919);
and U11030 (N_11030,N_7637,N_9105);
or U11031 (N_11031,N_9527,N_8569);
and U11032 (N_11032,N_9681,N_9518);
or U11033 (N_11033,N_9547,N_7584);
xnor U11034 (N_11034,N_7781,N_9208);
or U11035 (N_11035,N_8106,N_9969);
nor U11036 (N_11036,N_9013,N_8646);
and U11037 (N_11037,N_8657,N_9730);
nor U11038 (N_11038,N_7842,N_8987);
nand U11039 (N_11039,N_9192,N_8146);
or U11040 (N_11040,N_9695,N_7930);
nand U11041 (N_11041,N_7587,N_9089);
nor U11042 (N_11042,N_9267,N_8177);
nand U11043 (N_11043,N_7529,N_7755);
xnor U11044 (N_11044,N_8855,N_9274);
xor U11045 (N_11045,N_9712,N_9168);
or U11046 (N_11046,N_8463,N_7665);
nor U11047 (N_11047,N_8335,N_9305);
and U11048 (N_11048,N_7675,N_7991);
nor U11049 (N_11049,N_7807,N_9989);
nor U11050 (N_11050,N_7849,N_9621);
and U11051 (N_11051,N_8327,N_9687);
or U11052 (N_11052,N_7582,N_9258);
nand U11053 (N_11053,N_7790,N_9187);
or U11054 (N_11054,N_9072,N_9268);
and U11055 (N_11055,N_9766,N_9519);
nand U11056 (N_11056,N_8642,N_8915);
nand U11057 (N_11057,N_9206,N_8711);
nor U11058 (N_11058,N_9958,N_7810);
nand U11059 (N_11059,N_7594,N_9017);
nor U11060 (N_11060,N_8252,N_9332);
and U11061 (N_11061,N_8230,N_8577);
xor U11062 (N_11062,N_8192,N_9457);
and U11063 (N_11063,N_9629,N_9100);
nor U11064 (N_11064,N_8902,N_9709);
nand U11065 (N_11065,N_8550,N_8140);
or U11066 (N_11066,N_8044,N_9657);
nor U11067 (N_11067,N_9125,N_9290);
and U11068 (N_11068,N_7747,N_9254);
and U11069 (N_11069,N_8938,N_7813);
xnor U11070 (N_11070,N_9762,N_8143);
nor U11071 (N_11071,N_8239,N_8166);
xnor U11072 (N_11072,N_9727,N_7911);
nor U11073 (N_11073,N_9159,N_9881);
or U11074 (N_11074,N_9899,N_7978);
xnor U11075 (N_11075,N_9832,N_9790);
nor U11076 (N_11076,N_8492,N_8138);
or U11077 (N_11077,N_7961,N_9982);
nand U11078 (N_11078,N_8769,N_7969);
and U11079 (N_11079,N_7769,N_9720);
xnor U11080 (N_11080,N_9396,N_9714);
nor U11081 (N_11081,N_8903,N_8947);
and U11082 (N_11082,N_9024,N_9999);
or U11083 (N_11083,N_9276,N_8120);
nor U11084 (N_11084,N_9586,N_8520);
nand U11085 (N_11085,N_8203,N_9241);
xnor U11086 (N_11086,N_7581,N_7762);
and U11087 (N_11087,N_7933,N_9579);
nand U11088 (N_11088,N_9474,N_9010);
or U11089 (N_11089,N_8704,N_7701);
and U11090 (N_11090,N_7550,N_9666);
xor U11091 (N_11091,N_8134,N_9940);
or U11092 (N_11092,N_9897,N_8999);
or U11093 (N_11093,N_9773,N_7971);
nor U11094 (N_11094,N_7980,N_9566);
or U11095 (N_11095,N_7867,N_8263);
or U11096 (N_11096,N_9861,N_9069);
nor U11097 (N_11097,N_7787,N_8085);
and U11098 (N_11098,N_8150,N_7927);
xor U11099 (N_11099,N_9324,N_9436);
nand U11100 (N_11100,N_8951,N_9828);
nand U11101 (N_11101,N_8919,N_7709);
nor U11102 (N_11102,N_8832,N_7792);
nand U11103 (N_11103,N_9735,N_9117);
and U11104 (N_11104,N_8419,N_8563);
xnor U11105 (N_11105,N_9387,N_9510);
nor U11106 (N_11106,N_8343,N_9988);
xor U11107 (N_11107,N_8554,N_8337);
or U11108 (N_11108,N_9386,N_9977);
or U11109 (N_11109,N_9311,N_9705);
xnor U11110 (N_11110,N_9293,N_8906);
or U11111 (N_11111,N_9446,N_7619);
nor U11112 (N_11112,N_7888,N_8188);
nor U11113 (N_11113,N_7617,N_9394);
nor U11114 (N_11114,N_8806,N_9460);
nand U11115 (N_11115,N_9942,N_8605);
or U11116 (N_11116,N_8543,N_8002);
or U11117 (N_11117,N_9170,N_8400);
xnor U11118 (N_11118,N_8856,N_8961);
nand U11119 (N_11119,N_7979,N_9792);
nor U11120 (N_11120,N_9291,N_8627);
nand U11121 (N_11121,N_8336,N_9110);
xnor U11122 (N_11122,N_9151,N_9517);
nand U11123 (N_11123,N_7648,N_9700);
nor U11124 (N_11124,N_9644,N_8037);
nor U11125 (N_11125,N_8567,N_7844);
or U11126 (N_11126,N_8457,N_8927);
xor U11127 (N_11127,N_9326,N_8949);
nor U11128 (N_11128,N_7815,N_8872);
or U11129 (N_11129,N_8703,N_8200);
xnor U11130 (N_11130,N_7764,N_8687);
or U11131 (N_11131,N_9561,N_9059);
and U11132 (N_11132,N_8246,N_8176);
or U11133 (N_11133,N_9177,N_7716);
xnor U11134 (N_11134,N_8731,N_9612);
nand U11135 (N_11135,N_7559,N_9917);
or U11136 (N_11136,N_9842,N_9154);
and U11137 (N_11137,N_9800,N_8680);
nand U11138 (N_11138,N_9967,N_9742);
nand U11139 (N_11139,N_8935,N_9425);
and U11140 (N_11140,N_7761,N_8136);
nor U11141 (N_11141,N_8854,N_7848);
or U11142 (N_11142,N_9939,N_8556);
xor U11143 (N_11143,N_8852,N_7511);
xnor U11144 (N_11144,N_8045,N_8375);
or U11145 (N_11145,N_9947,N_8356);
xor U11146 (N_11146,N_7850,N_9298);
xnor U11147 (N_11147,N_7733,N_8043);
or U11148 (N_11148,N_7510,N_8771);
nor U11149 (N_11149,N_8829,N_8892);
or U11150 (N_11150,N_7773,N_9993);
or U11151 (N_11151,N_9148,N_8221);
or U11152 (N_11152,N_8255,N_8274);
or U11153 (N_11153,N_8306,N_9251);
nand U11154 (N_11154,N_7599,N_9420);
nor U11155 (N_11155,N_8957,N_9385);
and U11156 (N_11156,N_7554,N_8780);
nor U11157 (N_11157,N_8084,N_9791);
nand U11158 (N_11158,N_9256,N_8842);
nand U11159 (N_11159,N_9053,N_7883);
or U11160 (N_11160,N_7533,N_8315);
or U11161 (N_11161,N_9454,N_9429);
nor U11162 (N_11162,N_8691,N_9665);
or U11163 (N_11163,N_7904,N_8214);
and U11164 (N_11164,N_8945,N_9318);
and U11165 (N_11165,N_8883,N_8716);
and U11166 (N_11166,N_8873,N_8478);
xor U11167 (N_11167,N_9158,N_9103);
nor U11168 (N_11168,N_8815,N_8607);
or U11169 (N_11169,N_8290,N_7918);
nor U11170 (N_11170,N_8826,N_8139);
nor U11171 (N_11171,N_8323,N_8180);
or U11172 (N_11172,N_8761,N_9726);
nand U11173 (N_11173,N_8970,N_8179);
nor U11174 (N_11174,N_8682,N_7853);
nand U11175 (N_11175,N_8971,N_9230);
nor U11176 (N_11176,N_7878,N_9345);
and U11177 (N_11177,N_9826,N_9430);
or U11178 (N_11178,N_8631,N_9458);
or U11179 (N_11179,N_9819,N_7896);
nor U11180 (N_11180,N_9479,N_8161);
and U11181 (N_11181,N_9841,N_7631);
nand U11182 (N_11182,N_9770,N_8061);
nand U11183 (N_11183,N_8767,N_7548);
xnor U11184 (N_11184,N_8958,N_7572);
xnor U11185 (N_11185,N_8024,N_8714);
xor U11186 (N_11186,N_8216,N_9640);
and U11187 (N_11187,N_9129,N_7565);
and U11188 (N_11188,N_7805,N_7819);
nand U11189 (N_11189,N_7799,N_8676);
and U11190 (N_11190,N_9555,N_9388);
nand U11191 (N_11191,N_9306,N_7664);
xnor U11192 (N_11192,N_9451,N_9567);
xnor U11193 (N_11193,N_7700,N_9161);
xnor U11194 (N_11194,N_8640,N_9650);
nand U11195 (N_11195,N_8944,N_9339);
nor U11196 (N_11196,N_8491,N_8096);
xor U11197 (N_11197,N_9350,N_8977);
nor U11198 (N_11198,N_7870,N_7990);
xor U11199 (N_11199,N_9021,N_7856);
nor U11200 (N_11200,N_7782,N_9998);
and U11201 (N_11201,N_8517,N_9802);
or U11202 (N_11202,N_8499,N_7560);
and U11203 (N_11203,N_9925,N_9464);
nand U11204 (N_11204,N_8334,N_8033);
xor U11205 (N_11205,N_8847,N_9656);
and U11206 (N_11206,N_7947,N_8728);
nand U11207 (N_11207,N_9237,N_9796);
and U11208 (N_11208,N_9082,N_9322);
xnor U11209 (N_11209,N_7801,N_9859);
and U11210 (N_11210,N_8368,N_8840);
and U11211 (N_11211,N_7840,N_9763);
nor U11212 (N_11212,N_9009,N_9997);
or U11213 (N_11213,N_8442,N_7885);
nor U11214 (N_11214,N_9529,N_9506);
nor U11215 (N_11215,N_8470,N_7625);
and U11216 (N_11216,N_8110,N_8664);
nor U11217 (N_11217,N_9328,N_8887);
nor U11218 (N_11218,N_8481,N_8880);
and U11219 (N_11219,N_7925,N_8157);
nor U11220 (N_11220,N_8175,N_8049);
or U11221 (N_11221,N_8026,N_9057);
xnor U11222 (N_11222,N_8639,N_7775);
xor U11223 (N_11223,N_7926,N_8409);
or U11224 (N_11224,N_7901,N_8668);
nor U11225 (N_11225,N_9405,N_7779);
and U11226 (N_11226,N_7744,N_9041);
nor U11227 (N_11227,N_7794,N_8626);
nand U11228 (N_11228,N_9703,N_7677);
nand U11229 (N_11229,N_9390,N_9546);
or U11230 (N_11230,N_9937,N_9359);
xor U11231 (N_11231,N_7852,N_9046);
or U11232 (N_11232,N_8452,N_8185);
xnor U11233 (N_11233,N_9086,N_9798);
and U11234 (N_11234,N_8469,N_8755);
nand U11235 (N_11235,N_8459,N_9466);
nor U11236 (N_11236,N_8760,N_8575);
xnor U11237 (N_11237,N_8209,N_7836);
xnor U11238 (N_11238,N_7957,N_9898);
xor U11239 (N_11239,N_7846,N_9544);
xnor U11240 (N_11240,N_9310,N_8119);
or U11241 (N_11241,N_9108,N_8340);
nand U11242 (N_11242,N_7678,N_9034);
nand U11243 (N_11243,N_8194,N_8063);
or U11244 (N_11244,N_8921,N_7945);
or U11245 (N_11245,N_7624,N_9442);
nor U11246 (N_11246,N_9191,N_9837);
or U11247 (N_11247,N_9732,N_7865);
xor U11248 (N_11248,N_7939,N_7681);
or U11249 (N_11249,N_8468,N_7615);
and U11250 (N_11250,N_9447,N_8927);
nor U11251 (N_11251,N_9267,N_8635);
nor U11252 (N_11252,N_9121,N_7874);
nand U11253 (N_11253,N_7567,N_7732);
or U11254 (N_11254,N_9260,N_9148);
nor U11255 (N_11255,N_8782,N_8260);
nor U11256 (N_11256,N_9736,N_8249);
nor U11257 (N_11257,N_7980,N_9172);
or U11258 (N_11258,N_8391,N_8535);
xor U11259 (N_11259,N_8695,N_9288);
or U11260 (N_11260,N_9505,N_8261);
or U11261 (N_11261,N_8853,N_8405);
and U11262 (N_11262,N_7962,N_9105);
and U11263 (N_11263,N_8427,N_9125);
or U11264 (N_11264,N_8411,N_8739);
nor U11265 (N_11265,N_8956,N_8111);
and U11266 (N_11266,N_9412,N_8092);
xnor U11267 (N_11267,N_8674,N_9591);
and U11268 (N_11268,N_8798,N_8221);
nand U11269 (N_11269,N_7771,N_8699);
and U11270 (N_11270,N_8987,N_9838);
xnor U11271 (N_11271,N_7953,N_9735);
xnor U11272 (N_11272,N_9945,N_9487);
and U11273 (N_11273,N_8918,N_9743);
nor U11274 (N_11274,N_9840,N_9154);
xnor U11275 (N_11275,N_8839,N_8391);
nand U11276 (N_11276,N_7608,N_7840);
xor U11277 (N_11277,N_8352,N_8978);
xnor U11278 (N_11278,N_9628,N_8000);
xor U11279 (N_11279,N_9612,N_8168);
nor U11280 (N_11280,N_9876,N_8068);
or U11281 (N_11281,N_7689,N_7962);
or U11282 (N_11282,N_9292,N_9115);
nand U11283 (N_11283,N_8535,N_9198);
or U11284 (N_11284,N_9083,N_9934);
and U11285 (N_11285,N_7512,N_7838);
nor U11286 (N_11286,N_8725,N_9504);
or U11287 (N_11287,N_9250,N_7517);
nor U11288 (N_11288,N_9803,N_9644);
nand U11289 (N_11289,N_8766,N_8733);
nor U11290 (N_11290,N_8223,N_9883);
and U11291 (N_11291,N_8702,N_9525);
xor U11292 (N_11292,N_9317,N_7656);
nor U11293 (N_11293,N_9430,N_9905);
and U11294 (N_11294,N_9596,N_8303);
nand U11295 (N_11295,N_7713,N_7506);
or U11296 (N_11296,N_9314,N_8733);
or U11297 (N_11297,N_8728,N_7523);
nand U11298 (N_11298,N_8715,N_9581);
nor U11299 (N_11299,N_7534,N_9909);
nand U11300 (N_11300,N_7849,N_8983);
nand U11301 (N_11301,N_7848,N_9360);
and U11302 (N_11302,N_9088,N_8347);
nor U11303 (N_11303,N_8951,N_9733);
nand U11304 (N_11304,N_8465,N_9180);
xor U11305 (N_11305,N_9306,N_8773);
xnor U11306 (N_11306,N_9021,N_9440);
and U11307 (N_11307,N_9416,N_9429);
or U11308 (N_11308,N_8253,N_9082);
or U11309 (N_11309,N_7903,N_7677);
xnor U11310 (N_11310,N_8620,N_8528);
nand U11311 (N_11311,N_8210,N_8418);
nand U11312 (N_11312,N_8264,N_8842);
nor U11313 (N_11313,N_8884,N_7775);
and U11314 (N_11314,N_8803,N_9695);
nor U11315 (N_11315,N_8123,N_7838);
or U11316 (N_11316,N_8006,N_9856);
nor U11317 (N_11317,N_9550,N_9302);
nand U11318 (N_11318,N_8529,N_9283);
and U11319 (N_11319,N_9129,N_8609);
and U11320 (N_11320,N_8792,N_7516);
and U11321 (N_11321,N_8141,N_9485);
nor U11322 (N_11322,N_9538,N_9307);
or U11323 (N_11323,N_7741,N_9595);
xor U11324 (N_11324,N_8659,N_9813);
and U11325 (N_11325,N_8510,N_8000);
xor U11326 (N_11326,N_9292,N_9676);
nand U11327 (N_11327,N_8466,N_9529);
and U11328 (N_11328,N_8424,N_8163);
or U11329 (N_11329,N_7630,N_7585);
xor U11330 (N_11330,N_9660,N_9917);
nand U11331 (N_11331,N_9351,N_9483);
nor U11332 (N_11332,N_9813,N_9735);
nor U11333 (N_11333,N_8454,N_7702);
and U11334 (N_11334,N_7899,N_7559);
nor U11335 (N_11335,N_9393,N_7990);
nand U11336 (N_11336,N_8173,N_8186);
and U11337 (N_11337,N_8478,N_8487);
nor U11338 (N_11338,N_7732,N_9730);
nor U11339 (N_11339,N_8261,N_8473);
xor U11340 (N_11340,N_9691,N_8746);
xnor U11341 (N_11341,N_8367,N_8435);
nor U11342 (N_11342,N_8894,N_9996);
xor U11343 (N_11343,N_8573,N_9022);
or U11344 (N_11344,N_7894,N_7566);
nor U11345 (N_11345,N_8330,N_9443);
and U11346 (N_11346,N_7850,N_7786);
or U11347 (N_11347,N_9592,N_8944);
nor U11348 (N_11348,N_9398,N_7754);
or U11349 (N_11349,N_9623,N_9092);
or U11350 (N_11350,N_7691,N_9816);
or U11351 (N_11351,N_8355,N_8079);
and U11352 (N_11352,N_7605,N_9038);
and U11353 (N_11353,N_7758,N_8795);
xnor U11354 (N_11354,N_9432,N_7602);
and U11355 (N_11355,N_8987,N_8777);
and U11356 (N_11356,N_9498,N_8946);
nand U11357 (N_11357,N_8463,N_7792);
nand U11358 (N_11358,N_8759,N_9137);
or U11359 (N_11359,N_7694,N_9322);
nor U11360 (N_11360,N_9116,N_7516);
and U11361 (N_11361,N_7833,N_7776);
or U11362 (N_11362,N_9910,N_9092);
xor U11363 (N_11363,N_8728,N_9427);
nor U11364 (N_11364,N_9174,N_9684);
and U11365 (N_11365,N_7801,N_8748);
or U11366 (N_11366,N_7641,N_9736);
nor U11367 (N_11367,N_9984,N_7895);
and U11368 (N_11368,N_8051,N_9202);
and U11369 (N_11369,N_7713,N_9941);
and U11370 (N_11370,N_8144,N_9870);
and U11371 (N_11371,N_9984,N_9174);
nor U11372 (N_11372,N_9001,N_9986);
nand U11373 (N_11373,N_7574,N_7906);
nand U11374 (N_11374,N_7602,N_8996);
nand U11375 (N_11375,N_8096,N_9060);
nand U11376 (N_11376,N_9662,N_8561);
nor U11377 (N_11377,N_8937,N_8556);
and U11378 (N_11378,N_9475,N_9705);
nand U11379 (N_11379,N_9584,N_9719);
and U11380 (N_11380,N_7815,N_7978);
nand U11381 (N_11381,N_7513,N_9851);
nor U11382 (N_11382,N_7723,N_9418);
nor U11383 (N_11383,N_9304,N_9101);
or U11384 (N_11384,N_7608,N_7652);
nand U11385 (N_11385,N_9845,N_8929);
nand U11386 (N_11386,N_9123,N_9738);
xor U11387 (N_11387,N_9006,N_8824);
xor U11388 (N_11388,N_8836,N_8856);
xor U11389 (N_11389,N_7922,N_8104);
or U11390 (N_11390,N_9985,N_8593);
nand U11391 (N_11391,N_8328,N_9795);
nor U11392 (N_11392,N_8528,N_9080);
nor U11393 (N_11393,N_9169,N_9619);
nand U11394 (N_11394,N_8570,N_8691);
or U11395 (N_11395,N_7515,N_9072);
nor U11396 (N_11396,N_9661,N_7555);
and U11397 (N_11397,N_9652,N_8356);
xnor U11398 (N_11398,N_9325,N_9231);
xnor U11399 (N_11399,N_7973,N_8573);
xnor U11400 (N_11400,N_8249,N_9022);
nand U11401 (N_11401,N_9049,N_9948);
xnor U11402 (N_11402,N_7708,N_7602);
xor U11403 (N_11403,N_9716,N_9184);
xor U11404 (N_11404,N_9436,N_9808);
and U11405 (N_11405,N_8882,N_8872);
and U11406 (N_11406,N_7628,N_9177);
xnor U11407 (N_11407,N_8393,N_8217);
nand U11408 (N_11408,N_7926,N_8153);
nand U11409 (N_11409,N_9978,N_7572);
and U11410 (N_11410,N_8711,N_8382);
nand U11411 (N_11411,N_8465,N_9414);
and U11412 (N_11412,N_9382,N_8693);
nand U11413 (N_11413,N_9318,N_7740);
or U11414 (N_11414,N_8889,N_9838);
xor U11415 (N_11415,N_8790,N_8531);
nor U11416 (N_11416,N_8265,N_8651);
nand U11417 (N_11417,N_9016,N_9231);
xor U11418 (N_11418,N_8531,N_9975);
xnor U11419 (N_11419,N_7923,N_9294);
xor U11420 (N_11420,N_9281,N_8593);
xnor U11421 (N_11421,N_8719,N_8907);
or U11422 (N_11422,N_8272,N_9618);
and U11423 (N_11423,N_8155,N_9031);
nand U11424 (N_11424,N_7981,N_7761);
xor U11425 (N_11425,N_9628,N_9069);
xnor U11426 (N_11426,N_8595,N_8033);
or U11427 (N_11427,N_8968,N_9163);
or U11428 (N_11428,N_8097,N_8186);
or U11429 (N_11429,N_8032,N_9276);
nor U11430 (N_11430,N_9469,N_7867);
nand U11431 (N_11431,N_9357,N_9161);
xor U11432 (N_11432,N_9035,N_9022);
xor U11433 (N_11433,N_9827,N_9017);
or U11434 (N_11434,N_8936,N_9825);
or U11435 (N_11435,N_8909,N_9847);
and U11436 (N_11436,N_7862,N_7892);
nand U11437 (N_11437,N_8266,N_8806);
nor U11438 (N_11438,N_9663,N_8193);
nor U11439 (N_11439,N_9037,N_9709);
and U11440 (N_11440,N_8140,N_8215);
or U11441 (N_11441,N_9979,N_8264);
and U11442 (N_11442,N_9858,N_7612);
xnor U11443 (N_11443,N_9037,N_8237);
nor U11444 (N_11444,N_7678,N_9227);
nor U11445 (N_11445,N_9697,N_9578);
nor U11446 (N_11446,N_9646,N_8364);
xor U11447 (N_11447,N_8608,N_8670);
or U11448 (N_11448,N_8327,N_9006);
and U11449 (N_11449,N_9388,N_8694);
nand U11450 (N_11450,N_9139,N_7906);
and U11451 (N_11451,N_8901,N_8158);
nand U11452 (N_11452,N_9142,N_7711);
nand U11453 (N_11453,N_8443,N_7549);
or U11454 (N_11454,N_7807,N_8981);
xnor U11455 (N_11455,N_7945,N_9786);
xnor U11456 (N_11456,N_9579,N_8305);
nor U11457 (N_11457,N_9658,N_9844);
nand U11458 (N_11458,N_8572,N_8006);
and U11459 (N_11459,N_9580,N_8568);
and U11460 (N_11460,N_7942,N_9876);
and U11461 (N_11461,N_9434,N_8569);
or U11462 (N_11462,N_7734,N_8191);
nor U11463 (N_11463,N_7588,N_8751);
xor U11464 (N_11464,N_8417,N_9221);
nor U11465 (N_11465,N_7910,N_8602);
and U11466 (N_11466,N_8855,N_7818);
xnor U11467 (N_11467,N_8154,N_9841);
nor U11468 (N_11468,N_9027,N_8757);
xnor U11469 (N_11469,N_9928,N_9043);
nor U11470 (N_11470,N_7695,N_9708);
or U11471 (N_11471,N_7522,N_9264);
and U11472 (N_11472,N_8312,N_7846);
nand U11473 (N_11473,N_8654,N_7924);
nand U11474 (N_11474,N_7557,N_7672);
xor U11475 (N_11475,N_9066,N_7705);
and U11476 (N_11476,N_9905,N_9632);
or U11477 (N_11477,N_9967,N_7918);
and U11478 (N_11478,N_9403,N_9124);
nand U11479 (N_11479,N_9011,N_8549);
xor U11480 (N_11480,N_9574,N_8884);
and U11481 (N_11481,N_9316,N_8107);
and U11482 (N_11482,N_9179,N_7521);
nor U11483 (N_11483,N_7623,N_8914);
xnor U11484 (N_11484,N_9071,N_7854);
nor U11485 (N_11485,N_9749,N_9935);
nand U11486 (N_11486,N_8591,N_8458);
xor U11487 (N_11487,N_9237,N_8181);
nand U11488 (N_11488,N_9607,N_8622);
xor U11489 (N_11489,N_8597,N_8489);
xor U11490 (N_11490,N_8367,N_8222);
nand U11491 (N_11491,N_8653,N_7829);
and U11492 (N_11492,N_9269,N_8969);
xnor U11493 (N_11493,N_8201,N_7946);
or U11494 (N_11494,N_9735,N_9115);
nor U11495 (N_11495,N_9611,N_8282);
and U11496 (N_11496,N_8233,N_7744);
nand U11497 (N_11497,N_9402,N_8632);
nand U11498 (N_11498,N_8804,N_7735);
and U11499 (N_11499,N_8616,N_9202);
or U11500 (N_11500,N_7903,N_9749);
nor U11501 (N_11501,N_8217,N_8497);
nor U11502 (N_11502,N_7501,N_9542);
xor U11503 (N_11503,N_7571,N_8305);
nand U11504 (N_11504,N_8408,N_9186);
nor U11505 (N_11505,N_8397,N_8527);
and U11506 (N_11506,N_9915,N_7875);
xnor U11507 (N_11507,N_9153,N_9817);
or U11508 (N_11508,N_8537,N_9913);
and U11509 (N_11509,N_8258,N_8944);
and U11510 (N_11510,N_7671,N_9424);
nor U11511 (N_11511,N_9020,N_7976);
and U11512 (N_11512,N_8267,N_8895);
nor U11513 (N_11513,N_8915,N_8343);
or U11514 (N_11514,N_9663,N_9542);
nor U11515 (N_11515,N_8718,N_9460);
nand U11516 (N_11516,N_8767,N_8828);
nand U11517 (N_11517,N_9201,N_9569);
and U11518 (N_11518,N_8600,N_9062);
nand U11519 (N_11519,N_9435,N_9000);
xor U11520 (N_11520,N_8493,N_8572);
nand U11521 (N_11521,N_8576,N_9337);
or U11522 (N_11522,N_9416,N_9397);
and U11523 (N_11523,N_8898,N_8996);
and U11524 (N_11524,N_7867,N_9294);
xor U11525 (N_11525,N_9059,N_9660);
nand U11526 (N_11526,N_9167,N_7984);
nand U11527 (N_11527,N_8542,N_9453);
nor U11528 (N_11528,N_7693,N_8632);
xor U11529 (N_11529,N_9436,N_7684);
nand U11530 (N_11530,N_7574,N_9314);
and U11531 (N_11531,N_9248,N_7713);
or U11532 (N_11532,N_8762,N_7744);
and U11533 (N_11533,N_9825,N_9342);
and U11534 (N_11534,N_8129,N_8627);
or U11535 (N_11535,N_7685,N_9799);
xor U11536 (N_11536,N_8752,N_7661);
nand U11537 (N_11537,N_9713,N_8077);
nand U11538 (N_11538,N_8680,N_9279);
nand U11539 (N_11539,N_7510,N_8161);
or U11540 (N_11540,N_9965,N_9654);
xnor U11541 (N_11541,N_9806,N_9622);
or U11542 (N_11542,N_9589,N_9812);
and U11543 (N_11543,N_9365,N_8671);
and U11544 (N_11544,N_8801,N_8236);
nand U11545 (N_11545,N_9035,N_8547);
nand U11546 (N_11546,N_9998,N_9813);
and U11547 (N_11547,N_7727,N_8203);
nor U11548 (N_11548,N_7596,N_9647);
nor U11549 (N_11549,N_9741,N_8104);
or U11550 (N_11550,N_8725,N_8166);
and U11551 (N_11551,N_9493,N_9264);
and U11552 (N_11552,N_9126,N_8241);
and U11553 (N_11553,N_7731,N_8323);
and U11554 (N_11554,N_8792,N_8167);
nor U11555 (N_11555,N_8317,N_8577);
nand U11556 (N_11556,N_8709,N_8870);
nor U11557 (N_11557,N_9960,N_9567);
and U11558 (N_11558,N_9957,N_9338);
and U11559 (N_11559,N_8057,N_9743);
or U11560 (N_11560,N_9246,N_7542);
xor U11561 (N_11561,N_9002,N_9914);
and U11562 (N_11562,N_9861,N_8137);
or U11563 (N_11563,N_9116,N_8047);
nand U11564 (N_11564,N_8034,N_8110);
nor U11565 (N_11565,N_8021,N_9973);
nor U11566 (N_11566,N_9795,N_9244);
xor U11567 (N_11567,N_9579,N_8492);
nor U11568 (N_11568,N_9836,N_7861);
nor U11569 (N_11569,N_8214,N_8308);
or U11570 (N_11570,N_7719,N_9889);
or U11571 (N_11571,N_9366,N_8280);
nand U11572 (N_11572,N_8509,N_7677);
nor U11573 (N_11573,N_8499,N_7742);
and U11574 (N_11574,N_9366,N_8767);
nand U11575 (N_11575,N_9855,N_9512);
or U11576 (N_11576,N_9317,N_9740);
nor U11577 (N_11577,N_9375,N_7511);
or U11578 (N_11578,N_7529,N_9881);
nand U11579 (N_11579,N_8977,N_8758);
and U11580 (N_11580,N_7867,N_8514);
xor U11581 (N_11581,N_8412,N_8942);
nor U11582 (N_11582,N_9882,N_8458);
or U11583 (N_11583,N_9776,N_8655);
nand U11584 (N_11584,N_9115,N_9781);
nor U11585 (N_11585,N_9600,N_8291);
nand U11586 (N_11586,N_8269,N_8760);
or U11587 (N_11587,N_8288,N_8322);
nand U11588 (N_11588,N_9758,N_8922);
xnor U11589 (N_11589,N_8657,N_7957);
nor U11590 (N_11590,N_9189,N_9696);
nand U11591 (N_11591,N_7775,N_8435);
and U11592 (N_11592,N_8275,N_7798);
nand U11593 (N_11593,N_9720,N_9649);
or U11594 (N_11594,N_9284,N_9338);
and U11595 (N_11595,N_8252,N_8847);
or U11596 (N_11596,N_7594,N_9367);
or U11597 (N_11597,N_8530,N_9429);
xor U11598 (N_11598,N_7587,N_8012);
nand U11599 (N_11599,N_8611,N_7824);
or U11600 (N_11600,N_8573,N_7628);
nor U11601 (N_11601,N_7579,N_9219);
and U11602 (N_11602,N_8871,N_9683);
or U11603 (N_11603,N_8755,N_8738);
nand U11604 (N_11604,N_9724,N_8101);
xor U11605 (N_11605,N_8211,N_8594);
nand U11606 (N_11606,N_7697,N_8537);
or U11607 (N_11607,N_9158,N_7690);
xor U11608 (N_11608,N_9551,N_8579);
xor U11609 (N_11609,N_9029,N_9348);
nor U11610 (N_11610,N_8228,N_9429);
or U11611 (N_11611,N_7562,N_7754);
xor U11612 (N_11612,N_7526,N_8039);
nor U11613 (N_11613,N_9812,N_7625);
nand U11614 (N_11614,N_8465,N_8157);
and U11615 (N_11615,N_9191,N_7604);
and U11616 (N_11616,N_8027,N_8030);
nand U11617 (N_11617,N_8918,N_8753);
or U11618 (N_11618,N_8376,N_8751);
and U11619 (N_11619,N_7897,N_8586);
nor U11620 (N_11620,N_9185,N_7851);
or U11621 (N_11621,N_8228,N_9067);
and U11622 (N_11622,N_8116,N_8252);
nor U11623 (N_11623,N_9534,N_8467);
nor U11624 (N_11624,N_9413,N_7706);
or U11625 (N_11625,N_8343,N_9061);
and U11626 (N_11626,N_8903,N_8912);
nand U11627 (N_11627,N_8799,N_8887);
and U11628 (N_11628,N_9536,N_8306);
xor U11629 (N_11629,N_8874,N_8043);
xor U11630 (N_11630,N_9586,N_7510);
nor U11631 (N_11631,N_9617,N_7779);
or U11632 (N_11632,N_8988,N_9794);
xnor U11633 (N_11633,N_9129,N_9969);
and U11634 (N_11634,N_9308,N_7822);
and U11635 (N_11635,N_9913,N_7764);
and U11636 (N_11636,N_9096,N_9666);
nor U11637 (N_11637,N_8426,N_7582);
nand U11638 (N_11638,N_9887,N_7851);
nor U11639 (N_11639,N_8143,N_7697);
nor U11640 (N_11640,N_9035,N_8955);
nor U11641 (N_11641,N_8464,N_8923);
nand U11642 (N_11642,N_8751,N_8524);
and U11643 (N_11643,N_8625,N_7946);
or U11644 (N_11644,N_7531,N_9074);
and U11645 (N_11645,N_9407,N_8172);
nand U11646 (N_11646,N_8433,N_9007);
or U11647 (N_11647,N_7668,N_8598);
nor U11648 (N_11648,N_7769,N_8469);
xnor U11649 (N_11649,N_9639,N_9556);
nor U11650 (N_11650,N_9298,N_9419);
nor U11651 (N_11651,N_9985,N_9561);
xor U11652 (N_11652,N_8473,N_8281);
nand U11653 (N_11653,N_7511,N_8113);
nand U11654 (N_11654,N_8349,N_8709);
xnor U11655 (N_11655,N_8025,N_8522);
xnor U11656 (N_11656,N_9609,N_9670);
xor U11657 (N_11657,N_8997,N_9789);
nand U11658 (N_11658,N_8685,N_9870);
nand U11659 (N_11659,N_8782,N_9304);
or U11660 (N_11660,N_9679,N_8259);
or U11661 (N_11661,N_8923,N_8324);
nand U11662 (N_11662,N_8290,N_9990);
and U11663 (N_11663,N_9886,N_9436);
and U11664 (N_11664,N_9490,N_8406);
nor U11665 (N_11665,N_7966,N_8487);
or U11666 (N_11666,N_9395,N_9047);
nor U11667 (N_11667,N_9431,N_8923);
and U11668 (N_11668,N_8939,N_8993);
or U11669 (N_11669,N_8540,N_8842);
nand U11670 (N_11670,N_7977,N_8902);
nand U11671 (N_11671,N_8728,N_8193);
or U11672 (N_11672,N_8855,N_9031);
xor U11673 (N_11673,N_8417,N_7790);
nand U11674 (N_11674,N_8154,N_7663);
or U11675 (N_11675,N_8701,N_9465);
xor U11676 (N_11676,N_8914,N_9552);
and U11677 (N_11677,N_7584,N_7677);
or U11678 (N_11678,N_9670,N_7530);
or U11679 (N_11679,N_7721,N_9153);
or U11680 (N_11680,N_8253,N_8656);
xor U11681 (N_11681,N_8991,N_9622);
or U11682 (N_11682,N_9302,N_8896);
xor U11683 (N_11683,N_9482,N_9608);
nand U11684 (N_11684,N_8800,N_9939);
xnor U11685 (N_11685,N_8235,N_8271);
and U11686 (N_11686,N_7859,N_9470);
xor U11687 (N_11687,N_8582,N_8131);
or U11688 (N_11688,N_9848,N_8141);
nor U11689 (N_11689,N_8914,N_8408);
and U11690 (N_11690,N_8257,N_8681);
or U11691 (N_11691,N_8702,N_9084);
or U11692 (N_11692,N_9958,N_8176);
and U11693 (N_11693,N_8022,N_8534);
nor U11694 (N_11694,N_7677,N_8983);
and U11695 (N_11695,N_8494,N_9624);
xor U11696 (N_11696,N_8157,N_9782);
and U11697 (N_11697,N_9346,N_7648);
xor U11698 (N_11698,N_9264,N_8597);
xor U11699 (N_11699,N_8670,N_7749);
nand U11700 (N_11700,N_8891,N_9863);
nand U11701 (N_11701,N_7961,N_9419);
or U11702 (N_11702,N_9140,N_9724);
xor U11703 (N_11703,N_8045,N_7998);
or U11704 (N_11704,N_9028,N_9720);
nand U11705 (N_11705,N_9427,N_9265);
or U11706 (N_11706,N_8826,N_8565);
xnor U11707 (N_11707,N_8083,N_7965);
nor U11708 (N_11708,N_9822,N_9408);
xor U11709 (N_11709,N_9161,N_9282);
nor U11710 (N_11710,N_9203,N_8401);
or U11711 (N_11711,N_9856,N_8310);
and U11712 (N_11712,N_8979,N_8533);
or U11713 (N_11713,N_9569,N_8835);
and U11714 (N_11714,N_7656,N_7757);
xnor U11715 (N_11715,N_7512,N_8398);
or U11716 (N_11716,N_9866,N_9727);
nor U11717 (N_11717,N_9482,N_8301);
and U11718 (N_11718,N_9601,N_9095);
nand U11719 (N_11719,N_8419,N_9421);
and U11720 (N_11720,N_9921,N_8078);
nand U11721 (N_11721,N_8061,N_8057);
xor U11722 (N_11722,N_8522,N_7562);
and U11723 (N_11723,N_9216,N_8170);
nand U11724 (N_11724,N_8605,N_9324);
xor U11725 (N_11725,N_9407,N_7963);
and U11726 (N_11726,N_9694,N_7753);
xnor U11727 (N_11727,N_9381,N_8843);
nor U11728 (N_11728,N_9306,N_8183);
xor U11729 (N_11729,N_7979,N_9590);
nor U11730 (N_11730,N_9053,N_8540);
nand U11731 (N_11731,N_8132,N_9812);
or U11732 (N_11732,N_7969,N_8460);
and U11733 (N_11733,N_8729,N_9387);
xor U11734 (N_11734,N_8604,N_8730);
xor U11735 (N_11735,N_7575,N_9577);
and U11736 (N_11736,N_9863,N_8614);
nor U11737 (N_11737,N_9753,N_9497);
or U11738 (N_11738,N_8672,N_8813);
nand U11739 (N_11739,N_9223,N_9192);
xor U11740 (N_11740,N_8897,N_8333);
and U11741 (N_11741,N_8183,N_8895);
nor U11742 (N_11742,N_7943,N_8011);
xor U11743 (N_11743,N_7677,N_9932);
nand U11744 (N_11744,N_8016,N_8264);
or U11745 (N_11745,N_9035,N_8888);
nor U11746 (N_11746,N_9003,N_8144);
nor U11747 (N_11747,N_9761,N_8342);
nand U11748 (N_11748,N_7969,N_8858);
nor U11749 (N_11749,N_8946,N_9461);
and U11750 (N_11750,N_8119,N_8229);
and U11751 (N_11751,N_8732,N_7677);
and U11752 (N_11752,N_8095,N_7718);
and U11753 (N_11753,N_8405,N_9078);
or U11754 (N_11754,N_9398,N_9587);
and U11755 (N_11755,N_7794,N_7778);
nand U11756 (N_11756,N_9584,N_8429);
nand U11757 (N_11757,N_7620,N_7593);
or U11758 (N_11758,N_9814,N_8021);
nand U11759 (N_11759,N_7621,N_8889);
or U11760 (N_11760,N_8516,N_9595);
xnor U11761 (N_11761,N_8199,N_8116);
and U11762 (N_11762,N_8160,N_9910);
and U11763 (N_11763,N_8116,N_8823);
or U11764 (N_11764,N_8396,N_8155);
xor U11765 (N_11765,N_7660,N_9499);
or U11766 (N_11766,N_7898,N_7623);
nand U11767 (N_11767,N_7851,N_9547);
nor U11768 (N_11768,N_9841,N_7591);
nor U11769 (N_11769,N_8711,N_8202);
nor U11770 (N_11770,N_8725,N_9144);
and U11771 (N_11771,N_9446,N_9680);
xor U11772 (N_11772,N_7649,N_9917);
xnor U11773 (N_11773,N_8730,N_8757);
and U11774 (N_11774,N_8650,N_8229);
nor U11775 (N_11775,N_8151,N_7657);
and U11776 (N_11776,N_7742,N_9814);
and U11777 (N_11777,N_7805,N_8010);
nor U11778 (N_11778,N_9157,N_9505);
and U11779 (N_11779,N_7563,N_8970);
xnor U11780 (N_11780,N_7758,N_9647);
and U11781 (N_11781,N_9711,N_9338);
nand U11782 (N_11782,N_9186,N_7803);
xnor U11783 (N_11783,N_7606,N_9587);
xnor U11784 (N_11784,N_9609,N_8052);
xor U11785 (N_11785,N_9306,N_8767);
xnor U11786 (N_11786,N_7750,N_8826);
xor U11787 (N_11787,N_9263,N_8685);
and U11788 (N_11788,N_7868,N_8101);
and U11789 (N_11789,N_8120,N_8384);
xor U11790 (N_11790,N_8821,N_9197);
xnor U11791 (N_11791,N_8093,N_8930);
nand U11792 (N_11792,N_9057,N_9283);
nor U11793 (N_11793,N_7727,N_8378);
nand U11794 (N_11794,N_7534,N_8373);
and U11795 (N_11795,N_8671,N_8243);
xnor U11796 (N_11796,N_8012,N_9213);
xor U11797 (N_11797,N_8500,N_9110);
xor U11798 (N_11798,N_9385,N_8511);
nand U11799 (N_11799,N_8443,N_8045);
nand U11800 (N_11800,N_9658,N_8975);
nand U11801 (N_11801,N_9977,N_7868);
xor U11802 (N_11802,N_8794,N_7711);
or U11803 (N_11803,N_8139,N_8098);
and U11804 (N_11804,N_8130,N_9397);
xnor U11805 (N_11805,N_8499,N_8597);
and U11806 (N_11806,N_9014,N_9743);
and U11807 (N_11807,N_9979,N_9574);
nand U11808 (N_11808,N_8170,N_9503);
nor U11809 (N_11809,N_8356,N_9621);
or U11810 (N_11810,N_8016,N_9011);
and U11811 (N_11811,N_7949,N_8920);
nand U11812 (N_11812,N_7704,N_9750);
nand U11813 (N_11813,N_8254,N_9799);
nand U11814 (N_11814,N_8120,N_7571);
xor U11815 (N_11815,N_9385,N_7756);
xnor U11816 (N_11816,N_7801,N_7765);
or U11817 (N_11817,N_8143,N_9241);
and U11818 (N_11818,N_9117,N_7946);
xor U11819 (N_11819,N_8915,N_7595);
or U11820 (N_11820,N_9413,N_7974);
nor U11821 (N_11821,N_8876,N_9854);
or U11822 (N_11822,N_9729,N_8851);
nor U11823 (N_11823,N_9684,N_8316);
nor U11824 (N_11824,N_9615,N_8953);
xor U11825 (N_11825,N_8748,N_9823);
or U11826 (N_11826,N_9308,N_7775);
nor U11827 (N_11827,N_9164,N_8901);
or U11828 (N_11828,N_9479,N_8865);
and U11829 (N_11829,N_7910,N_7624);
or U11830 (N_11830,N_8103,N_9542);
nor U11831 (N_11831,N_7606,N_8088);
or U11832 (N_11832,N_7911,N_9186);
xor U11833 (N_11833,N_8720,N_9593);
nor U11834 (N_11834,N_9574,N_8247);
and U11835 (N_11835,N_7975,N_9761);
nor U11836 (N_11836,N_8462,N_9454);
nor U11837 (N_11837,N_9807,N_8756);
xor U11838 (N_11838,N_8103,N_7866);
and U11839 (N_11839,N_8023,N_9666);
or U11840 (N_11840,N_8979,N_9904);
and U11841 (N_11841,N_7608,N_7982);
nand U11842 (N_11842,N_8122,N_9500);
or U11843 (N_11843,N_8504,N_8665);
nand U11844 (N_11844,N_9030,N_9500);
nor U11845 (N_11845,N_7714,N_9380);
nand U11846 (N_11846,N_8646,N_9416);
xor U11847 (N_11847,N_8756,N_8701);
or U11848 (N_11848,N_8763,N_8585);
nand U11849 (N_11849,N_8868,N_9897);
xnor U11850 (N_11850,N_9961,N_7975);
xor U11851 (N_11851,N_9317,N_8579);
and U11852 (N_11852,N_8199,N_8935);
xnor U11853 (N_11853,N_9664,N_8471);
or U11854 (N_11854,N_9073,N_7760);
and U11855 (N_11855,N_7523,N_7963);
and U11856 (N_11856,N_8423,N_8146);
nand U11857 (N_11857,N_8784,N_9870);
xor U11858 (N_11858,N_9213,N_7515);
xnor U11859 (N_11859,N_8078,N_9233);
nand U11860 (N_11860,N_9885,N_7980);
nor U11861 (N_11861,N_7694,N_7813);
nand U11862 (N_11862,N_9647,N_9419);
and U11863 (N_11863,N_8677,N_9215);
nand U11864 (N_11864,N_8318,N_7889);
or U11865 (N_11865,N_9053,N_9324);
nor U11866 (N_11866,N_8079,N_7521);
and U11867 (N_11867,N_8290,N_9538);
or U11868 (N_11868,N_9195,N_9437);
nor U11869 (N_11869,N_9115,N_7948);
xor U11870 (N_11870,N_8682,N_7677);
or U11871 (N_11871,N_9025,N_7749);
nor U11872 (N_11872,N_9781,N_8103);
nor U11873 (N_11873,N_8693,N_9901);
or U11874 (N_11874,N_8565,N_9198);
nor U11875 (N_11875,N_9595,N_9095);
and U11876 (N_11876,N_9191,N_8758);
and U11877 (N_11877,N_8860,N_9553);
nor U11878 (N_11878,N_8086,N_9797);
xor U11879 (N_11879,N_8130,N_8837);
and U11880 (N_11880,N_9583,N_8228);
and U11881 (N_11881,N_9980,N_7899);
or U11882 (N_11882,N_9424,N_8258);
nor U11883 (N_11883,N_9219,N_7688);
nor U11884 (N_11884,N_7670,N_9178);
or U11885 (N_11885,N_9930,N_8907);
and U11886 (N_11886,N_8025,N_9624);
xnor U11887 (N_11887,N_9958,N_9363);
and U11888 (N_11888,N_8695,N_9521);
xnor U11889 (N_11889,N_9334,N_8941);
and U11890 (N_11890,N_8634,N_9426);
nand U11891 (N_11891,N_9143,N_7863);
nand U11892 (N_11892,N_9049,N_7994);
nor U11893 (N_11893,N_8236,N_8342);
nand U11894 (N_11894,N_9455,N_9359);
nand U11895 (N_11895,N_9068,N_9688);
xnor U11896 (N_11896,N_8479,N_9238);
nor U11897 (N_11897,N_9388,N_9272);
nor U11898 (N_11898,N_8812,N_9531);
or U11899 (N_11899,N_8589,N_9601);
or U11900 (N_11900,N_8704,N_8015);
or U11901 (N_11901,N_8495,N_9541);
and U11902 (N_11902,N_8544,N_8455);
nand U11903 (N_11903,N_9728,N_8296);
or U11904 (N_11904,N_8230,N_7968);
or U11905 (N_11905,N_8304,N_8909);
and U11906 (N_11906,N_9482,N_8975);
nand U11907 (N_11907,N_9303,N_9088);
and U11908 (N_11908,N_7807,N_9542);
nand U11909 (N_11909,N_8281,N_7713);
or U11910 (N_11910,N_9420,N_8352);
nand U11911 (N_11911,N_7764,N_9040);
nand U11912 (N_11912,N_8455,N_7509);
nand U11913 (N_11913,N_8346,N_8375);
nand U11914 (N_11914,N_8318,N_9655);
nand U11915 (N_11915,N_8209,N_7614);
or U11916 (N_11916,N_9031,N_9781);
xor U11917 (N_11917,N_9217,N_9377);
or U11918 (N_11918,N_8374,N_9109);
or U11919 (N_11919,N_9988,N_8140);
nand U11920 (N_11920,N_9283,N_8588);
xnor U11921 (N_11921,N_9868,N_9850);
and U11922 (N_11922,N_9668,N_9727);
xor U11923 (N_11923,N_8742,N_9660);
or U11924 (N_11924,N_8259,N_7865);
and U11925 (N_11925,N_8237,N_8587);
xor U11926 (N_11926,N_8153,N_9760);
nor U11927 (N_11927,N_8514,N_7572);
xor U11928 (N_11928,N_9705,N_9460);
xor U11929 (N_11929,N_7750,N_7722);
nand U11930 (N_11930,N_9942,N_8006);
nor U11931 (N_11931,N_9128,N_8788);
xor U11932 (N_11932,N_7533,N_7648);
and U11933 (N_11933,N_9637,N_8895);
or U11934 (N_11934,N_8859,N_7971);
nand U11935 (N_11935,N_9669,N_9869);
or U11936 (N_11936,N_8107,N_9772);
nor U11937 (N_11937,N_9143,N_7544);
or U11938 (N_11938,N_8697,N_9151);
and U11939 (N_11939,N_8362,N_9610);
nand U11940 (N_11940,N_8295,N_9439);
and U11941 (N_11941,N_7679,N_7916);
xnor U11942 (N_11942,N_8337,N_9253);
nor U11943 (N_11943,N_7569,N_9855);
or U11944 (N_11944,N_7980,N_7683);
xnor U11945 (N_11945,N_8865,N_8465);
xnor U11946 (N_11946,N_7587,N_8686);
or U11947 (N_11947,N_8140,N_8931);
or U11948 (N_11948,N_7816,N_8247);
nor U11949 (N_11949,N_9801,N_8832);
and U11950 (N_11950,N_7832,N_9050);
xnor U11951 (N_11951,N_8229,N_9375);
nor U11952 (N_11952,N_8655,N_9443);
or U11953 (N_11953,N_8930,N_9874);
and U11954 (N_11954,N_7731,N_7508);
or U11955 (N_11955,N_8994,N_8449);
nor U11956 (N_11956,N_8712,N_7842);
xor U11957 (N_11957,N_8120,N_7560);
xor U11958 (N_11958,N_9579,N_9244);
nand U11959 (N_11959,N_8595,N_8629);
nor U11960 (N_11960,N_7894,N_7514);
nand U11961 (N_11961,N_7707,N_9771);
and U11962 (N_11962,N_8265,N_7902);
xor U11963 (N_11963,N_7741,N_7600);
or U11964 (N_11964,N_7989,N_8089);
nor U11965 (N_11965,N_7813,N_7965);
and U11966 (N_11966,N_9644,N_7713);
or U11967 (N_11967,N_7506,N_9684);
xor U11968 (N_11968,N_8860,N_9136);
nor U11969 (N_11969,N_9008,N_7602);
or U11970 (N_11970,N_8499,N_9465);
and U11971 (N_11971,N_9914,N_7786);
or U11972 (N_11972,N_8549,N_9727);
or U11973 (N_11973,N_8703,N_9217);
nand U11974 (N_11974,N_9663,N_8104);
xor U11975 (N_11975,N_8738,N_9933);
nor U11976 (N_11976,N_8438,N_8511);
nand U11977 (N_11977,N_9939,N_9756);
nor U11978 (N_11978,N_8624,N_7735);
nor U11979 (N_11979,N_8895,N_7607);
or U11980 (N_11980,N_8439,N_9391);
xor U11981 (N_11981,N_9628,N_7695);
nor U11982 (N_11982,N_8597,N_9913);
or U11983 (N_11983,N_9471,N_9178);
xor U11984 (N_11984,N_8682,N_9356);
xor U11985 (N_11985,N_8077,N_8506);
xor U11986 (N_11986,N_8823,N_8848);
xor U11987 (N_11987,N_8135,N_9044);
xnor U11988 (N_11988,N_8389,N_8012);
nand U11989 (N_11989,N_7703,N_9338);
nor U11990 (N_11990,N_8185,N_8838);
or U11991 (N_11991,N_9358,N_9619);
or U11992 (N_11992,N_8415,N_8542);
or U11993 (N_11993,N_7839,N_8162);
or U11994 (N_11994,N_8340,N_8094);
nor U11995 (N_11995,N_9369,N_8645);
xor U11996 (N_11996,N_7735,N_9551);
nor U11997 (N_11997,N_7620,N_9805);
and U11998 (N_11998,N_8587,N_8618);
nor U11999 (N_11999,N_7954,N_8619);
or U12000 (N_12000,N_8074,N_8370);
nor U12001 (N_12001,N_9569,N_9872);
nor U12002 (N_12002,N_9278,N_8912);
nand U12003 (N_12003,N_7500,N_7940);
or U12004 (N_12004,N_9875,N_8374);
nand U12005 (N_12005,N_8677,N_9876);
and U12006 (N_12006,N_8464,N_7971);
nor U12007 (N_12007,N_8076,N_8199);
or U12008 (N_12008,N_8029,N_7731);
or U12009 (N_12009,N_9705,N_8277);
and U12010 (N_12010,N_7795,N_9120);
nand U12011 (N_12011,N_9691,N_9877);
nand U12012 (N_12012,N_8723,N_8224);
or U12013 (N_12013,N_7550,N_9578);
or U12014 (N_12014,N_7594,N_8376);
or U12015 (N_12015,N_9231,N_7704);
nor U12016 (N_12016,N_8717,N_8651);
or U12017 (N_12017,N_9934,N_9627);
or U12018 (N_12018,N_7949,N_9074);
and U12019 (N_12019,N_8059,N_8795);
xnor U12020 (N_12020,N_8845,N_8720);
nand U12021 (N_12021,N_8092,N_8363);
or U12022 (N_12022,N_9310,N_8427);
or U12023 (N_12023,N_9272,N_7863);
nand U12024 (N_12024,N_7912,N_7513);
nand U12025 (N_12025,N_9763,N_7888);
and U12026 (N_12026,N_8230,N_9745);
and U12027 (N_12027,N_9473,N_9408);
or U12028 (N_12028,N_7776,N_8885);
xor U12029 (N_12029,N_9567,N_7891);
and U12030 (N_12030,N_8326,N_7629);
nand U12031 (N_12031,N_9002,N_9128);
and U12032 (N_12032,N_8217,N_9870);
nand U12033 (N_12033,N_9385,N_8220);
nand U12034 (N_12034,N_8673,N_9936);
nand U12035 (N_12035,N_7783,N_9923);
and U12036 (N_12036,N_9786,N_7985);
or U12037 (N_12037,N_7773,N_9052);
or U12038 (N_12038,N_8863,N_8209);
and U12039 (N_12039,N_8058,N_7620);
xnor U12040 (N_12040,N_7819,N_7638);
and U12041 (N_12041,N_7728,N_8829);
nand U12042 (N_12042,N_8367,N_7843);
nor U12043 (N_12043,N_7732,N_7840);
xor U12044 (N_12044,N_8909,N_8029);
nor U12045 (N_12045,N_7839,N_8758);
nor U12046 (N_12046,N_8406,N_8967);
and U12047 (N_12047,N_8906,N_7874);
or U12048 (N_12048,N_7686,N_8471);
and U12049 (N_12049,N_9215,N_9159);
nor U12050 (N_12050,N_9190,N_9277);
nor U12051 (N_12051,N_8791,N_9944);
or U12052 (N_12052,N_7849,N_8239);
nand U12053 (N_12053,N_9123,N_9024);
nand U12054 (N_12054,N_7790,N_9204);
nor U12055 (N_12055,N_7772,N_8167);
xor U12056 (N_12056,N_9165,N_9042);
and U12057 (N_12057,N_9409,N_8070);
nor U12058 (N_12058,N_9089,N_7621);
and U12059 (N_12059,N_8092,N_9554);
xor U12060 (N_12060,N_9007,N_8157);
and U12061 (N_12061,N_7975,N_8529);
nor U12062 (N_12062,N_9095,N_8286);
or U12063 (N_12063,N_8353,N_9476);
nor U12064 (N_12064,N_9961,N_8721);
nor U12065 (N_12065,N_9989,N_9845);
xor U12066 (N_12066,N_9274,N_9798);
nor U12067 (N_12067,N_7955,N_8902);
nand U12068 (N_12068,N_8125,N_7510);
xor U12069 (N_12069,N_8936,N_9951);
and U12070 (N_12070,N_9577,N_8492);
xnor U12071 (N_12071,N_9610,N_8882);
nand U12072 (N_12072,N_9700,N_8312);
or U12073 (N_12073,N_9289,N_9993);
and U12074 (N_12074,N_9059,N_7715);
or U12075 (N_12075,N_8943,N_8415);
or U12076 (N_12076,N_8785,N_9044);
and U12077 (N_12077,N_8025,N_7655);
nor U12078 (N_12078,N_9528,N_9386);
and U12079 (N_12079,N_9811,N_9994);
or U12080 (N_12080,N_9467,N_9005);
nor U12081 (N_12081,N_8083,N_8893);
nor U12082 (N_12082,N_8920,N_9695);
nor U12083 (N_12083,N_9569,N_9792);
nor U12084 (N_12084,N_9806,N_7704);
nor U12085 (N_12085,N_9926,N_8314);
nand U12086 (N_12086,N_7518,N_7605);
and U12087 (N_12087,N_8507,N_9026);
nand U12088 (N_12088,N_7681,N_8585);
xnor U12089 (N_12089,N_8573,N_9857);
xor U12090 (N_12090,N_8104,N_9358);
or U12091 (N_12091,N_9239,N_8671);
nor U12092 (N_12092,N_7953,N_9624);
xor U12093 (N_12093,N_8253,N_7552);
nand U12094 (N_12094,N_8069,N_9483);
or U12095 (N_12095,N_8592,N_9749);
and U12096 (N_12096,N_9396,N_8127);
nor U12097 (N_12097,N_8347,N_9316);
or U12098 (N_12098,N_8984,N_9670);
or U12099 (N_12099,N_8894,N_9712);
nand U12100 (N_12100,N_9922,N_9583);
and U12101 (N_12101,N_7931,N_9991);
and U12102 (N_12102,N_8610,N_7629);
and U12103 (N_12103,N_9869,N_8940);
nand U12104 (N_12104,N_8319,N_8307);
and U12105 (N_12105,N_9604,N_8609);
or U12106 (N_12106,N_8586,N_7836);
xor U12107 (N_12107,N_8827,N_7792);
nand U12108 (N_12108,N_8652,N_8569);
or U12109 (N_12109,N_8029,N_9434);
nor U12110 (N_12110,N_8930,N_9098);
and U12111 (N_12111,N_7510,N_9696);
nand U12112 (N_12112,N_8955,N_8670);
xnor U12113 (N_12113,N_8878,N_8138);
and U12114 (N_12114,N_9438,N_8117);
nand U12115 (N_12115,N_9644,N_8588);
and U12116 (N_12116,N_7582,N_9737);
xor U12117 (N_12117,N_9482,N_8974);
or U12118 (N_12118,N_9430,N_8303);
and U12119 (N_12119,N_7736,N_9982);
xor U12120 (N_12120,N_9412,N_9825);
or U12121 (N_12121,N_8544,N_9958);
xor U12122 (N_12122,N_8695,N_9516);
or U12123 (N_12123,N_7523,N_8282);
xor U12124 (N_12124,N_9381,N_8080);
and U12125 (N_12125,N_7972,N_9937);
nand U12126 (N_12126,N_8875,N_9066);
and U12127 (N_12127,N_8208,N_9617);
nand U12128 (N_12128,N_9526,N_9723);
xor U12129 (N_12129,N_9314,N_9661);
and U12130 (N_12130,N_9648,N_7605);
nand U12131 (N_12131,N_8861,N_8153);
xor U12132 (N_12132,N_7744,N_8948);
xnor U12133 (N_12133,N_8765,N_7941);
nor U12134 (N_12134,N_7736,N_8510);
nand U12135 (N_12135,N_8288,N_7949);
xnor U12136 (N_12136,N_7647,N_8063);
nand U12137 (N_12137,N_9267,N_7641);
and U12138 (N_12138,N_8162,N_7581);
nor U12139 (N_12139,N_7853,N_7826);
xor U12140 (N_12140,N_8250,N_7914);
or U12141 (N_12141,N_8772,N_9709);
and U12142 (N_12142,N_7730,N_9403);
nor U12143 (N_12143,N_7616,N_8951);
nor U12144 (N_12144,N_9633,N_8576);
xor U12145 (N_12145,N_8854,N_9148);
xnor U12146 (N_12146,N_7595,N_9906);
nand U12147 (N_12147,N_8905,N_9590);
and U12148 (N_12148,N_7672,N_7520);
nand U12149 (N_12149,N_8188,N_9643);
and U12150 (N_12150,N_9978,N_9864);
and U12151 (N_12151,N_9069,N_9750);
and U12152 (N_12152,N_8847,N_9090);
xor U12153 (N_12153,N_8891,N_8971);
nand U12154 (N_12154,N_8989,N_7646);
nand U12155 (N_12155,N_9284,N_8537);
nand U12156 (N_12156,N_9008,N_7680);
nor U12157 (N_12157,N_7906,N_8428);
and U12158 (N_12158,N_8648,N_7513);
nand U12159 (N_12159,N_8391,N_8493);
and U12160 (N_12160,N_7682,N_8567);
nor U12161 (N_12161,N_8859,N_9390);
and U12162 (N_12162,N_8826,N_7547);
and U12163 (N_12163,N_8130,N_9349);
or U12164 (N_12164,N_9450,N_9274);
nor U12165 (N_12165,N_9645,N_8001);
nor U12166 (N_12166,N_9638,N_9832);
nor U12167 (N_12167,N_8934,N_7941);
nand U12168 (N_12168,N_9138,N_7763);
nor U12169 (N_12169,N_8445,N_9758);
and U12170 (N_12170,N_9345,N_8116);
nor U12171 (N_12171,N_8925,N_7755);
xor U12172 (N_12172,N_7750,N_8464);
nand U12173 (N_12173,N_8728,N_7903);
and U12174 (N_12174,N_8918,N_8557);
nand U12175 (N_12175,N_9213,N_7687);
xor U12176 (N_12176,N_9619,N_8576);
nand U12177 (N_12177,N_7852,N_8512);
and U12178 (N_12178,N_7777,N_8221);
xor U12179 (N_12179,N_7769,N_8204);
nand U12180 (N_12180,N_8077,N_8336);
and U12181 (N_12181,N_7975,N_9462);
nand U12182 (N_12182,N_8573,N_9754);
nor U12183 (N_12183,N_9413,N_7951);
or U12184 (N_12184,N_8143,N_8222);
xor U12185 (N_12185,N_7678,N_7640);
xor U12186 (N_12186,N_7979,N_7795);
nor U12187 (N_12187,N_9008,N_8160);
xnor U12188 (N_12188,N_7746,N_9541);
and U12189 (N_12189,N_9458,N_9323);
and U12190 (N_12190,N_7785,N_9583);
or U12191 (N_12191,N_9137,N_8388);
nor U12192 (N_12192,N_8571,N_9034);
nand U12193 (N_12193,N_7729,N_9625);
nor U12194 (N_12194,N_8874,N_7838);
xor U12195 (N_12195,N_9779,N_8225);
nand U12196 (N_12196,N_8402,N_8451);
xor U12197 (N_12197,N_7572,N_8649);
or U12198 (N_12198,N_9444,N_8662);
and U12199 (N_12199,N_8230,N_9043);
and U12200 (N_12200,N_9351,N_9156);
nand U12201 (N_12201,N_7785,N_9802);
xnor U12202 (N_12202,N_7531,N_7853);
xor U12203 (N_12203,N_9323,N_8310);
and U12204 (N_12204,N_8218,N_7637);
and U12205 (N_12205,N_9807,N_8302);
or U12206 (N_12206,N_7635,N_9127);
nand U12207 (N_12207,N_8352,N_9388);
and U12208 (N_12208,N_8529,N_9765);
and U12209 (N_12209,N_9489,N_8684);
nor U12210 (N_12210,N_8272,N_9312);
or U12211 (N_12211,N_8255,N_9055);
nor U12212 (N_12212,N_8946,N_8225);
nor U12213 (N_12213,N_8950,N_8462);
xnor U12214 (N_12214,N_9593,N_8880);
nor U12215 (N_12215,N_8051,N_7717);
nor U12216 (N_12216,N_7586,N_7825);
nand U12217 (N_12217,N_9944,N_8172);
xor U12218 (N_12218,N_7674,N_7946);
nor U12219 (N_12219,N_9086,N_9552);
xor U12220 (N_12220,N_9856,N_8906);
and U12221 (N_12221,N_9028,N_8018);
and U12222 (N_12222,N_9378,N_8529);
or U12223 (N_12223,N_9651,N_9712);
or U12224 (N_12224,N_8075,N_7559);
and U12225 (N_12225,N_8041,N_7522);
xor U12226 (N_12226,N_8776,N_9192);
xnor U12227 (N_12227,N_9020,N_8822);
or U12228 (N_12228,N_9463,N_9646);
nor U12229 (N_12229,N_9444,N_9517);
nor U12230 (N_12230,N_8905,N_7858);
or U12231 (N_12231,N_9793,N_9218);
or U12232 (N_12232,N_7695,N_8277);
and U12233 (N_12233,N_8659,N_8591);
nor U12234 (N_12234,N_7772,N_9899);
nor U12235 (N_12235,N_7721,N_8551);
or U12236 (N_12236,N_9150,N_7699);
nand U12237 (N_12237,N_8470,N_9811);
or U12238 (N_12238,N_9353,N_8577);
nor U12239 (N_12239,N_9791,N_8134);
nand U12240 (N_12240,N_8849,N_8243);
xor U12241 (N_12241,N_9459,N_9395);
nor U12242 (N_12242,N_8473,N_9053);
nand U12243 (N_12243,N_8566,N_9657);
xnor U12244 (N_12244,N_8792,N_7848);
xnor U12245 (N_12245,N_8526,N_7571);
or U12246 (N_12246,N_9312,N_8843);
nand U12247 (N_12247,N_7778,N_8109);
nand U12248 (N_12248,N_7734,N_9407);
or U12249 (N_12249,N_9262,N_9841);
nor U12250 (N_12250,N_8465,N_9676);
nand U12251 (N_12251,N_8477,N_7727);
xor U12252 (N_12252,N_9327,N_9282);
nor U12253 (N_12253,N_8503,N_8766);
and U12254 (N_12254,N_9315,N_9429);
nand U12255 (N_12255,N_8205,N_9459);
or U12256 (N_12256,N_9183,N_7547);
and U12257 (N_12257,N_7860,N_8994);
and U12258 (N_12258,N_8930,N_9126);
nor U12259 (N_12259,N_8249,N_8332);
nor U12260 (N_12260,N_9411,N_7664);
xnor U12261 (N_12261,N_8302,N_8619);
xor U12262 (N_12262,N_7743,N_9409);
nand U12263 (N_12263,N_7998,N_7738);
nor U12264 (N_12264,N_9018,N_8658);
xnor U12265 (N_12265,N_8847,N_9145);
and U12266 (N_12266,N_7857,N_9259);
nand U12267 (N_12267,N_8300,N_8843);
nand U12268 (N_12268,N_9718,N_9621);
nor U12269 (N_12269,N_7641,N_9951);
nor U12270 (N_12270,N_8931,N_8390);
or U12271 (N_12271,N_9298,N_7820);
and U12272 (N_12272,N_9275,N_8124);
and U12273 (N_12273,N_9442,N_7718);
nand U12274 (N_12274,N_7528,N_7867);
or U12275 (N_12275,N_7837,N_8593);
xnor U12276 (N_12276,N_9106,N_9537);
or U12277 (N_12277,N_8155,N_9554);
nand U12278 (N_12278,N_9847,N_9259);
nor U12279 (N_12279,N_8137,N_8533);
or U12280 (N_12280,N_8045,N_9798);
nand U12281 (N_12281,N_9800,N_7941);
nand U12282 (N_12282,N_7893,N_8055);
and U12283 (N_12283,N_8326,N_8548);
nor U12284 (N_12284,N_7988,N_7907);
nor U12285 (N_12285,N_9003,N_7635);
nand U12286 (N_12286,N_7622,N_8340);
nand U12287 (N_12287,N_9939,N_9139);
and U12288 (N_12288,N_8874,N_8223);
xnor U12289 (N_12289,N_7809,N_7841);
xor U12290 (N_12290,N_9139,N_7887);
and U12291 (N_12291,N_8366,N_9204);
nor U12292 (N_12292,N_9505,N_8318);
nand U12293 (N_12293,N_8691,N_7613);
nand U12294 (N_12294,N_8355,N_8551);
or U12295 (N_12295,N_8901,N_9203);
or U12296 (N_12296,N_8823,N_9396);
nand U12297 (N_12297,N_9276,N_9752);
and U12298 (N_12298,N_8291,N_9513);
nand U12299 (N_12299,N_8913,N_8544);
and U12300 (N_12300,N_8862,N_7814);
and U12301 (N_12301,N_9575,N_7862);
xor U12302 (N_12302,N_9644,N_7671);
nand U12303 (N_12303,N_9214,N_8608);
xor U12304 (N_12304,N_8720,N_8803);
xor U12305 (N_12305,N_9723,N_9156);
xnor U12306 (N_12306,N_7757,N_8433);
nand U12307 (N_12307,N_9128,N_9408);
or U12308 (N_12308,N_9438,N_8260);
nor U12309 (N_12309,N_9768,N_8311);
xor U12310 (N_12310,N_7687,N_7844);
or U12311 (N_12311,N_9706,N_9250);
and U12312 (N_12312,N_9596,N_8337);
or U12313 (N_12313,N_8023,N_9303);
nor U12314 (N_12314,N_9110,N_7954);
nor U12315 (N_12315,N_7636,N_7576);
and U12316 (N_12316,N_7870,N_8219);
nor U12317 (N_12317,N_9950,N_9480);
or U12318 (N_12318,N_8667,N_9891);
or U12319 (N_12319,N_8835,N_9865);
and U12320 (N_12320,N_8711,N_9021);
xnor U12321 (N_12321,N_7793,N_8016);
and U12322 (N_12322,N_8263,N_9426);
nand U12323 (N_12323,N_8897,N_9653);
nor U12324 (N_12324,N_8349,N_9924);
xor U12325 (N_12325,N_8142,N_7500);
nand U12326 (N_12326,N_8772,N_7778);
and U12327 (N_12327,N_8382,N_7833);
nand U12328 (N_12328,N_8200,N_7649);
xnor U12329 (N_12329,N_9189,N_7761);
or U12330 (N_12330,N_8416,N_9873);
xor U12331 (N_12331,N_9841,N_9404);
xor U12332 (N_12332,N_8129,N_8763);
or U12333 (N_12333,N_8041,N_9866);
and U12334 (N_12334,N_9268,N_9419);
and U12335 (N_12335,N_9607,N_8848);
xnor U12336 (N_12336,N_9006,N_9842);
or U12337 (N_12337,N_9093,N_9197);
and U12338 (N_12338,N_8560,N_8726);
xor U12339 (N_12339,N_9677,N_8626);
and U12340 (N_12340,N_9271,N_9028);
or U12341 (N_12341,N_7550,N_9822);
or U12342 (N_12342,N_9558,N_7694);
and U12343 (N_12343,N_7598,N_8341);
nand U12344 (N_12344,N_8154,N_8351);
and U12345 (N_12345,N_9699,N_9519);
nand U12346 (N_12346,N_7934,N_7887);
nor U12347 (N_12347,N_9789,N_9731);
and U12348 (N_12348,N_8864,N_9885);
or U12349 (N_12349,N_8646,N_7702);
and U12350 (N_12350,N_9576,N_9305);
nor U12351 (N_12351,N_9175,N_9452);
nand U12352 (N_12352,N_8302,N_9683);
nand U12353 (N_12353,N_8776,N_7577);
or U12354 (N_12354,N_9567,N_9169);
xor U12355 (N_12355,N_9633,N_9736);
nand U12356 (N_12356,N_9969,N_8634);
nand U12357 (N_12357,N_8176,N_8782);
and U12358 (N_12358,N_8468,N_8882);
nand U12359 (N_12359,N_9694,N_7654);
nor U12360 (N_12360,N_8811,N_8438);
nor U12361 (N_12361,N_9708,N_7613);
xor U12362 (N_12362,N_9115,N_8941);
nor U12363 (N_12363,N_9652,N_9510);
nand U12364 (N_12364,N_9644,N_8640);
nor U12365 (N_12365,N_8131,N_8231);
or U12366 (N_12366,N_8343,N_8932);
nand U12367 (N_12367,N_8977,N_7957);
nand U12368 (N_12368,N_9571,N_9252);
or U12369 (N_12369,N_9744,N_8636);
nand U12370 (N_12370,N_7805,N_8552);
xor U12371 (N_12371,N_7841,N_9847);
or U12372 (N_12372,N_8674,N_8696);
nor U12373 (N_12373,N_9245,N_8302);
nand U12374 (N_12374,N_8049,N_9182);
nand U12375 (N_12375,N_8421,N_9570);
and U12376 (N_12376,N_7967,N_7645);
nor U12377 (N_12377,N_9436,N_9006);
and U12378 (N_12378,N_8156,N_7767);
and U12379 (N_12379,N_9884,N_9778);
nor U12380 (N_12380,N_7922,N_8433);
nor U12381 (N_12381,N_8031,N_8576);
and U12382 (N_12382,N_7925,N_8250);
nand U12383 (N_12383,N_8117,N_9208);
nand U12384 (N_12384,N_8788,N_7505);
or U12385 (N_12385,N_8929,N_9020);
nand U12386 (N_12386,N_9287,N_9346);
and U12387 (N_12387,N_9009,N_7753);
or U12388 (N_12388,N_7807,N_9487);
xnor U12389 (N_12389,N_8094,N_9895);
xor U12390 (N_12390,N_9605,N_8753);
nor U12391 (N_12391,N_9551,N_8539);
nor U12392 (N_12392,N_8180,N_8030);
or U12393 (N_12393,N_8157,N_8785);
or U12394 (N_12394,N_8433,N_8987);
nor U12395 (N_12395,N_9261,N_9848);
nor U12396 (N_12396,N_8589,N_8377);
nor U12397 (N_12397,N_9385,N_9925);
xnor U12398 (N_12398,N_7946,N_8915);
and U12399 (N_12399,N_8033,N_8402);
nor U12400 (N_12400,N_9266,N_7770);
and U12401 (N_12401,N_8716,N_7573);
nor U12402 (N_12402,N_8618,N_8280);
nor U12403 (N_12403,N_8632,N_9463);
or U12404 (N_12404,N_9124,N_9793);
and U12405 (N_12405,N_9654,N_8492);
nand U12406 (N_12406,N_7596,N_9093);
or U12407 (N_12407,N_8825,N_7567);
nand U12408 (N_12408,N_9362,N_9185);
or U12409 (N_12409,N_9894,N_9802);
nand U12410 (N_12410,N_9813,N_8789);
and U12411 (N_12411,N_9255,N_7874);
nor U12412 (N_12412,N_7653,N_9612);
nand U12413 (N_12413,N_8348,N_9601);
xnor U12414 (N_12414,N_8672,N_8988);
nand U12415 (N_12415,N_8398,N_8295);
nand U12416 (N_12416,N_8400,N_7846);
xor U12417 (N_12417,N_8237,N_9616);
or U12418 (N_12418,N_7787,N_8533);
nand U12419 (N_12419,N_9551,N_9184);
nand U12420 (N_12420,N_7580,N_8208);
or U12421 (N_12421,N_9565,N_7775);
and U12422 (N_12422,N_8975,N_7553);
nand U12423 (N_12423,N_9878,N_7762);
xnor U12424 (N_12424,N_8975,N_8509);
xnor U12425 (N_12425,N_7509,N_9973);
xor U12426 (N_12426,N_8395,N_8687);
xor U12427 (N_12427,N_8347,N_9075);
xnor U12428 (N_12428,N_9867,N_9699);
and U12429 (N_12429,N_8688,N_9692);
or U12430 (N_12430,N_8827,N_9640);
xnor U12431 (N_12431,N_9200,N_9812);
nand U12432 (N_12432,N_8381,N_8351);
nor U12433 (N_12433,N_9596,N_9280);
nand U12434 (N_12434,N_8573,N_7941);
xor U12435 (N_12435,N_9297,N_9174);
nand U12436 (N_12436,N_8305,N_8941);
nand U12437 (N_12437,N_9782,N_9854);
nand U12438 (N_12438,N_7803,N_9344);
xnor U12439 (N_12439,N_8874,N_8508);
and U12440 (N_12440,N_9766,N_8198);
nor U12441 (N_12441,N_8744,N_8225);
nand U12442 (N_12442,N_9915,N_8847);
nand U12443 (N_12443,N_8637,N_8972);
xnor U12444 (N_12444,N_9194,N_9204);
or U12445 (N_12445,N_9005,N_8772);
or U12446 (N_12446,N_7571,N_9008);
nand U12447 (N_12447,N_8450,N_8383);
and U12448 (N_12448,N_9664,N_9596);
and U12449 (N_12449,N_8094,N_9848);
or U12450 (N_12450,N_8501,N_8742);
xor U12451 (N_12451,N_8262,N_9505);
or U12452 (N_12452,N_9238,N_9160);
and U12453 (N_12453,N_7843,N_8176);
xnor U12454 (N_12454,N_8018,N_8050);
nor U12455 (N_12455,N_8497,N_9724);
nor U12456 (N_12456,N_9378,N_8613);
xnor U12457 (N_12457,N_7871,N_8050);
nor U12458 (N_12458,N_7997,N_9811);
and U12459 (N_12459,N_9403,N_8041);
nand U12460 (N_12460,N_9754,N_9952);
nand U12461 (N_12461,N_9041,N_9779);
xor U12462 (N_12462,N_8894,N_8892);
or U12463 (N_12463,N_8385,N_8323);
nor U12464 (N_12464,N_9666,N_8432);
and U12465 (N_12465,N_9104,N_9381);
or U12466 (N_12466,N_9966,N_9917);
and U12467 (N_12467,N_9854,N_9655);
or U12468 (N_12468,N_9639,N_7828);
xor U12469 (N_12469,N_9150,N_7592);
and U12470 (N_12470,N_9449,N_8226);
nand U12471 (N_12471,N_8926,N_8735);
and U12472 (N_12472,N_9482,N_9947);
xnor U12473 (N_12473,N_8034,N_8180);
nand U12474 (N_12474,N_7848,N_9052);
xnor U12475 (N_12475,N_7775,N_9721);
or U12476 (N_12476,N_7736,N_9881);
xnor U12477 (N_12477,N_8243,N_9773);
xor U12478 (N_12478,N_9874,N_7739);
xor U12479 (N_12479,N_9868,N_8847);
nand U12480 (N_12480,N_8451,N_9796);
nand U12481 (N_12481,N_7841,N_9503);
nand U12482 (N_12482,N_7658,N_8840);
or U12483 (N_12483,N_8554,N_9489);
or U12484 (N_12484,N_9762,N_9575);
nand U12485 (N_12485,N_8508,N_8463);
xor U12486 (N_12486,N_8785,N_9782);
or U12487 (N_12487,N_8498,N_9290);
xnor U12488 (N_12488,N_9500,N_9290);
nor U12489 (N_12489,N_9235,N_8139);
xor U12490 (N_12490,N_9408,N_9383);
and U12491 (N_12491,N_8663,N_7811);
nand U12492 (N_12492,N_9065,N_8989);
xor U12493 (N_12493,N_8648,N_7536);
nor U12494 (N_12494,N_8361,N_9380);
nor U12495 (N_12495,N_7842,N_7732);
xnor U12496 (N_12496,N_7661,N_8171);
and U12497 (N_12497,N_9779,N_8944);
nor U12498 (N_12498,N_7506,N_8670);
nand U12499 (N_12499,N_9588,N_8348);
xnor U12500 (N_12500,N_12427,N_11624);
xnor U12501 (N_12501,N_11499,N_10657);
or U12502 (N_12502,N_10469,N_11974);
nand U12503 (N_12503,N_12495,N_11238);
or U12504 (N_12504,N_10609,N_12459);
and U12505 (N_12505,N_11159,N_10590);
nand U12506 (N_12506,N_11464,N_11224);
and U12507 (N_12507,N_12447,N_10567);
and U12508 (N_12508,N_11562,N_11750);
xor U12509 (N_12509,N_11380,N_10053);
xnor U12510 (N_12510,N_11665,N_10734);
xor U12511 (N_12511,N_11104,N_11094);
nor U12512 (N_12512,N_12349,N_10160);
xnor U12513 (N_12513,N_10763,N_10117);
or U12514 (N_12514,N_10833,N_10549);
and U12515 (N_12515,N_10244,N_12087);
and U12516 (N_12516,N_11424,N_11091);
nor U12517 (N_12517,N_11272,N_10937);
xnor U12518 (N_12518,N_11827,N_11821);
and U12519 (N_12519,N_10996,N_10111);
and U12520 (N_12520,N_12372,N_11412);
xor U12521 (N_12521,N_11641,N_10258);
nand U12522 (N_12522,N_12010,N_10843);
xnor U12523 (N_12523,N_10808,N_11218);
xnor U12524 (N_12524,N_11907,N_12211);
xnor U12525 (N_12525,N_11168,N_10642);
xor U12526 (N_12526,N_12364,N_10551);
or U12527 (N_12527,N_11889,N_12411);
or U12528 (N_12528,N_10685,N_10901);
nor U12529 (N_12529,N_11014,N_11186);
or U12530 (N_12530,N_12445,N_10182);
xnor U12531 (N_12531,N_12022,N_10449);
and U12532 (N_12532,N_11814,N_11400);
or U12533 (N_12533,N_11275,N_12353);
nand U12534 (N_12534,N_11637,N_11708);
or U12535 (N_12535,N_11900,N_10080);
nand U12536 (N_12536,N_10109,N_12057);
xor U12537 (N_12537,N_10806,N_10380);
nor U12538 (N_12538,N_10761,N_11269);
nor U12539 (N_12539,N_11385,N_10351);
or U12540 (N_12540,N_11735,N_10048);
or U12541 (N_12541,N_10968,N_10706);
nor U12542 (N_12542,N_12428,N_10526);
xnor U12543 (N_12543,N_11959,N_11375);
nand U12544 (N_12544,N_11683,N_11266);
nand U12545 (N_12545,N_11939,N_10035);
and U12546 (N_12546,N_11520,N_12272);
nor U12547 (N_12547,N_11219,N_11942);
nand U12548 (N_12548,N_10429,N_11663);
and U12549 (N_12549,N_12007,N_11132);
or U12550 (N_12550,N_10569,N_12258);
and U12551 (N_12551,N_11461,N_10520);
xnor U12552 (N_12552,N_10142,N_11930);
nand U12553 (N_12553,N_10457,N_12037);
xor U12554 (N_12554,N_11926,N_11246);
xnor U12555 (N_12555,N_11801,N_11475);
nor U12556 (N_12556,N_12336,N_10556);
xnor U12557 (N_12557,N_10592,N_10508);
nor U12558 (N_12558,N_12361,N_10804);
nor U12559 (N_12559,N_11027,N_10497);
and U12560 (N_12560,N_12152,N_11072);
nor U12561 (N_12561,N_11032,N_10991);
and U12562 (N_12562,N_11000,N_10897);
xnor U12563 (N_12563,N_12449,N_10702);
and U12564 (N_12564,N_10153,N_11722);
and U12565 (N_12565,N_11941,N_11728);
nand U12566 (N_12566,N_11998,N_10286);
and U12567 (N_12567,N_10411,N_11618);
nor U12568 (N_12568,N_11441,N_11182);
nor U12569 (N_12569,N_11241,N_12288);
or U12570 (N_12570,N_10493,N_12252);
nand U12571 (N_12571,N_11668,N_10326);
xor U12572 (N_12572,N_10980,N_10423);
or U12573 (N_12573,N_11096,N_10122);
or U12574 (N_12574,N_11395,N_10445);
nand U12575 (N_12575,N_11770,N_10077);
nand U12576 (N_12576,N_10369,N_11541);
xor U12577 (N_12577,N_11554,N_10249);
nand U12578 (N_12578,N_11732,N_11929);
nor U12579 (N_12579,N_11397,N_11011);
or U12580 (N_12580,N_11351,N_12292);
or U12581 (N_12581,N_12457,N_10951);
or U12582 (N_12582,N_11766,N_10613);
nand U12583 (N_12583,N_12480,N_10066);
nor U12584 (N_12584,N_12492,N_10263);
or U12585 (N_12585,N_10013,N_11048);
nor U12586 (N_12586,N_12233,N_12180);
or U12587 (N_12587,N_11629,N_10916);
and U12588 (N_12588,N_11830,N_11674);
and U12589 (N_12589,N_11713,N_11955);
nor U12590 (N_12590,N_12337,N_11632);
and U12591 (N_12591,N_12226,N_10585);
xor U12592 (N_12592,N_11374,N_10417);
nand U12593 (N_12593,N_12198,N_11928);
xor U12594 (N_12594,N_11281,N_10269);
nor U12595 (N_12595,N_11954,N_10056);
nor U12596 (N_12596,N_10938,N_11625);
xor U12597 (N_12597,N_12385,N_12170);
and U12598 (N_12598,N_10643,N_11856);
nand U12599 (N_12599,N_11913,N_10272);
xnor U12600 (N_12600,N_12270,N_10061);
nor U12601 (N_12601,N_11899,N_10076);
xor U12602 (N_12602,N_11515,N_10416);
nand U12603 (N_12603,N_12329,N_10754);
or U12604 (N_12604,N_11428,N_10479);
nor U12605 (N_12605,N_11612,N_10055);
or U12606 (N_12606,N_10157,N_11070);
xor U12607 (N_12607,N_11640,N_12316);
nor U12608 (N_12608,N_10426,N_11324);
xor U12609 (N_12609,N_12222,N_12267);
nand U12610 (N_12610,N_11059,N_12109);
nor U12611 (N_12611,N_10335,N_12467);
nand U12612 (N_12612,N_11411,N_11533);
xnor U12613 (N_12613,N_11106,N_11079);
and U12614 (N_12614,N_10633,N_11359);
and U12615 (N_12615,N_10752,N_11843);
nor U12616 (N_12616,N_11378,N_11114);
xnor U12617 (N_12617,N_12444,N_11084);
and U12618 (N_12618,N_11992,N_11600);
nor U12619 (N_12619,N_10791,N_10782);
or U12620 (N_12620,N_11905,N_11200);
xnor U12621 (N_12621,N_10972,N_11321);
xnor U12622 (N_12622,N_11245,N_11524);
nor U12623 (N_12623,N_10009,N_10820);
and U12624 (N_12624,N_10525,N_12308);
nor U12625 (N_12625,N_10383,N_11588);
nor U12626 (N_12626,N_11230,N_12038);
nor U12627 (N_12627,N_11042,N_10384);
nor U12628 (N_12628,N_11968,N_10583);
or U12629 (N_12629,N_10072,N_12432);
nor U12630 (N_12630,N_11152,N_11053);
and U12631 (N_12631,N_12391,N_10559);
or U12632 (N_12632,N_11675,N_12334);
nor U12633 (N_12633,N_10166,N_10612);
or U12634 (N_12634,N_10719,N_11308);
xor U12635 (N_12635,N_10807,N_12118);
nand U12636 (N_12636,N_10409,N_10862);
and U12637 (N_12637,N_10329,N_10623);
xor U12638 (N_12638,N_10145,N_10490);
and U12639 (N_12639,N_11251,N_11172);
and U12640 (N_12640,N_10994,N_11818);
nor U12641 (N_12641,N_10029,N_12499);
nand U12642 (N_12642,N_10043,N_12307);
nor U12643 (N_12643,N_11195,N_10577);
and U12644 (N_12644,N_10415,N_11613);
xor U12645 (N_12645,N_11088,N_12042);
or U12646 (N_12646,N_11769,N_11466);
nor U12647 (N_12647,N_11537,N_10582);
and U12648 (N_12648,N_11690,N_10016);
and U12649 (N_12649,N_10733,N_11216);
or U12650 (N_12650,N_12435,N_10505);
xor U12651 (N_12651,N_11903,N_12023);
nor U12652 (N_12652,N_10507,N_11639);
nor U12653 (N_12653,N_11416,N_11381);
nand U12654 (N_12654,N_11473,N_11006);
nor U12655 (N_12655,N_12327,N_11121);
nor U12656 (N_12656,N_12441,N_12205);
xor U12657 (N_12657,N_10163,N_11509);
and U12658 (N_12658,N_10535,N_11495);
xnor U12659 (N_12659,N_11952,N_11505);
and U12660 (N_12660,N_11825,N_10750);
or U12661 (N_12661,N_11883,N_10026);
nand U12662 (N_12662,N_10017,N_12303);
or U12663 (N_12663,N_12021,N_11366);
xor U12664 (N_12664,N_10971,N_11702);
nand U12665 (N_12665,N_11972,N_11760);
nor U12666 (N_12666,N_11575,N_11022);
nor U12667 (N_12667,N_11782,N_11243);
and U12668 (N_12668,N_11463,N_12130);
nor U12669 (N_12669,N_12423,N_10467);
and U12670 (N_12670,N_11966,N_12473);
or U12671 (N_12671,N_11166,N_12401);
and U12672 (N_12672,N_11623,N_12145);
and U12673 (N_12673,N_11310,N_12187);
or U12674 (N_12674,N_12373,N_10087);
nor U12675 (N_12675,N_10841,N_12297);
nor U12676 (N_12676,N_10516,N_12408);
nor U12677 (N_12677,N_11016,N_10599);
nand U12678 (N_12678,N_11797,N_11469);
or U12679 (N_12679,N_11858,N_10958);
and U12680 (N_12680,N_10755,N_11815);
or U12681 (N_12681,N_10579,N_11566);
or U12682 (N_12682,N_11868,N_11589);
xor U12683 (N_12683,N_12494,N_10581);
nand U12684 (N_12684,N_11286,N_11456);
nor U12685 (N_12685,N_12063,N_10736);
nor U12686 (N_12686,N_12490,N_10855);
nor U12687 (N_12687,N_11250,N_11044);
nand U12688 (N_12688,N_10290,N_10267);
or U12689 (N_12689,N_10014,N_10046);
nand U12690 (N_12690,N_12067,N_10760);
xnor U12691 (N_12691,N_12363,N_12069);
nand U12692 (N_12692,N_11633,N_11795);
nand U12693 (N_12693,N_12246,N_11871);
or U12694 (N_12694,N_11707,N_10941);
nand U12695 (N_12695,N_11301,N_10953);
nand U12696 (N_12696,N_11291,N_12485);
xor U12697 (N_12697,N_11130,N_12347);
nand U12698 (N_12698,N_12017,N_10187);
nand U12699 (N_12699,N_11470,N_12192);
and U12700 (N_12700,N_11787,N_11692);
nor U12701 (N_12701,N_10159,N_11817);
xnor U12702 (N_12702,N_10461,N_11339);
xor U12703 (N_12703,N_10596,N_11529);
xnor U12704 (N_12704,N_11488,N_10969);
or U12705 (N_12705,N_11978,N_11360);
and U12706 (N_12706,N_10717,N_12181);
nand U12707 (N_12707,N_11785,N_12281);
nand U12708 (N_12708,N_10407,N_12020);
and U12709 (N_12709,N_11323,N_11671);
or U12710 (N_12710,N_10798,N_12218);
and U12711 (N_12711,N_10375,N_11631);
nor U12712 (N_12712,N_10434,N_11676);
or U12713 (N_12713,N_11514,N_12279);
and U12714 (N_12714,N_10280,N_10718);
or U12715 (N_12715,N_11264,N_11962);
xor U12716 (N_12716,N_10175,N_11489);
nand U12717 (N_12717,N_11687,N_10898);
xnor U12718 (N_12718,N_12350,N_10176);
xnor U12719 (N_12719,N_12393,N_11727);
nor U12720 (N_12720,N_12050,N_10872);
nor U12721 (N_12721,N_11109,N_12210);
and U12722 (N_12722,N_10907,N_11240);
xnor U12723 (N_12723,N_11398,N_11806);
xnor U12724 (N_12724,N_11848,N_11384);
nor U12725 (N_12725,N_10195,N_10031);
xor U12726 (N_12726,N_11136,N_11571);
nand U12727 (N_12727,N_10611,N_12131);
and U12728 (N_12728,N_10406,N_12129);
and U12729 (N_12729,N_10876,N_10970);
nor U12730 (N_12730,N_10438,N_11560);
and U12731 (N_12731,N_12165,N_11666);
or U12732 (N_12732,N_12249,N_10494);
nor U12733 (N_12733,N_12462,N_10295);
nand U12734 (N_12734,N_10730,N_11531);
nor U12735 (N_12735,N_10805,N_12151);
nor U12736 (N_12736,N_11517,N_10923);
xnor U12737 (N_12737,N_11128,N_10977);
xnor U12738 (N_12738,N_11828,N_10487);
nand U12739 (N_12739,N_10931,N_10568);
and U12740 (N_12740,N_10044,N_10322);
or U12741 (N_12741,N_11309,N_11902);
or U12742 (N_12742,N_11145,N_11895);
nor U12743 (N_12743,N_10127,N_10037);
and U12744 (N_12744,N_11338,N_11574);
nand U12745 (N_12745,N_10709,N_11936);
and U12746 (N_12746,N_11890,N_10541);
or U12747 (N_12747,N_10388,N_11764);
and U12748 (N_12748,N_11578,N_11617);
nand U12749 (N_12749,N_11918,N_11596);
or U12750 (N_12750,N_10889,N_11957);
nand U12751 (N_12751,N_12225,N_10676);
nand U12752 (N_12752,N_10352,N_11607);
nand U12753 (N_12753,N_11300,N_11696);
or U12754 (N_12754,N_12477,N_11142);
nor U12755 (N_12755,N_11661,N_12139);
or U12756 (N_12756,N_12240,N_11544);
or U12757 (N_12757,N_10000,N_10155);
nor U12758 (N_12758,N_11755,N_12196);
nand U12759 (N_12759,N_10878,N_10981);
and U12760 (N_12760,N_12236,N_11893);
xor U12761 (N_12761,N_10238,N_11069);
nand U12762 (N_12762,N_10363,N_10962);
nor U12763 (N_12763,N_12434,N_10165);
or U12764 (N_12764,N_11345,N_12284);
nor U12765 (N_12765,N_11915,N_11382);
and U12766 (N_12766,N_10894,N_10131);
nor U12767 (N_12767,N_11174,N_11140);
nor U12768 (N_12768,N_12128,N_11584);
nand U12769 (N_12769,N_10892,N_10699);
xor U12770 (N_12770,N_12138,N_10631);
nand U12771 (N_12771,N_11294,N_11151);
xor U12772 (N_12772,N_10903,N_12250);
and U12773 (N_12773,N_10119,N_10832);
nor U12774 (N_12774,N_10687,N_12403);
xnor U12775 (N_12775,N_10584,N_11963);
and U12776 (N_12776,N_12355,N_10105);
or U12777 (N_12777,N_11803,N_10476);
nor U12778 (N_12778,N_12458,N_11812);
xnor U12779 (N_12779,N_12259,N_11144);
nor U12780 (N_12780,N_11552,N_11223);
and U12781 (N_12781,N_10049,N_11153);
nand U12782 (N_12782,N_11045,N_10501);
nor U12783 (N_12783,N_10557,N_12018);
xor U12784 (N_12784,N_11256,N_11860);
nand U12785 (N_12785,N_12464,N_12164);
nand U12786 (N_12786,N_11660,N_11759);
nand U12787 (N_12787,N_12224,N_11352);
or U12788 (N_12788,N_11282,N_11539);
xor U12789 (N_12789,N_11320,N_10391);
and U12790 (N_12790,N_10141,N_10517);
or U12791 (N_12791,N_12331,N_11302);
nand U12792 (N_12792,N_12471,N_11415);
or U12793 (N_12793,N_12387,N_11001);
nand U12794 (N_12794,N_12009,N_12352);
xnor U12795 (N_12795,N_12256,N_11154);
or U12796 (N_12796,N_11160,N_11709);
xor U12797 (N_12797,N_10513,N_10271);
or U12798 (N_12798,N_10108,N_12275);
and U12799 (N_12799,N_11158,N_11932);
nand U12800 (N_12800,N_10193,N_12304);
nand U12801 (N_12801,N_11569,N_10337);
and U12802 (N_12802,N_11725,N_12206);
and U12803 (N_12803,N_10431,N_10543);
or U12804 (N_12804,N_12371,N_10020);
xnor U12805 (N_12805,N_10462,N_10846);
and U12806 (N_12806,N_11831,N_10902);
and U12807 (N_12807,N_12463,N_10886);
or U12808 (N_12808,N_11744,N_12008);
xnor U12809 (N_12809,N_12289,N_11976);
xor U12810 (N_12810,N_10936,N_10877);
and U12811 (N_12811,N_11943,N_12024);
xor U12812 (N_12812,N_11211,N_12268);
xor U12813 (N_12813,N_10514,N_11947);
nand U12814 (N_12814,N_12419,N_10860);
and U12815 (N_12815,N_12443,N_10885);
nand U12816 (N_12816,N_11587,N_12147);
nor U12817 (N_12817,N_11861,N_11143);
xor U12818 (N_12818,N_11399,N_10226);
xor U12819 (N_12819,N_12003,N_11285);
and U12820 (N_12820,N_12141,N_12199);
nand U12821 (N_12821,N_10812,N_10181);
and U12822 (N_12822,N_11226,N_11228);
nand U12823 (N_12823,N_10089,N_10914);
nor U12824 (N_12824,N_10961,N_10795);
xor U12825 (N_12825,N_11191,N_10527);
nand U12826 (N_12826,N_10368,N_10632);
nor U12827 (N_12827,N_12340,N_10059);
and U12828 (N_12828,N_11206,N_11009);
xnor U12829 (N_12829,N_10118,N_11793);
xnor U12830 (N_12830,N_11118,N_11884);
nand U12831 (N_12831,N_10975,N_11171);
nand U12832 (N_12832,N_12412,N_10540);
and U12833 (N_12833,N_11066,N_10635);
nand U12834 (N_12834,N_10146,N_10616);
and U12835 (N_12835,N_10197,N_10819);
and U12836 (N_12836,N_11741,N_10148);
xnor U12837 (N_12837,N_10291,N_10453);
nand U12838 (N_12838,N_11227,N_10560);
nor U12839 (N_12839,N_11579,N_10742);
nor U12840 (N_12840,N_11842,N_10666);
nor U12841 (N_12841,N_10600,N_11894);
nor U12842 (N_12842,N_11789,N_11838);
nor U12843 (N_12843,N_10988,N_10485);
or U12844 (N_12844,N_11307,N_10854);
xnor U12845 (N_12845,N_12166,N_10521);
or U12846 (N_12846,N_11527,N_11317);
or U12847 (N_12847,N_10664,N_11185);
nor U12848 (N_12848,N_10716,N_10942);
or U12849 (N_12849,N_10587,N_10617);
nor U12850 (N_12850,N_11844,N_12001);
nand U12851 (N_12851,N_11414,N_12150);
xnor U12852 (N_12852,N_11492,N_11577);
xnor U12853 (N_12853,N_11512,N_10829);
xor U12854 (N_12854,N_11076,N_10315);
nor U12855 (N_12855,N_12048,N_12148);
or U12856 (N_12856,N_11874,N_11887);
nand U12857 (N_12857,N_11846,N_10670);
nor U12858 (N_12858,N_11064,N_10740);
and U12859 (N_12859,N_10356,N_10194);
xor U12860 (N_12860,N_12342,N_11327);
and U12861 (N_12861,N_10484,N_10308);
and U12862 (N_12862,N_10324,N_10661);
nor U12863 (N_12863,N_12169,N_11592);
nor U12864 (N_12864,N_10311,N_11901);
nor U12865 (N_12865,N_10850,N_10439);
nor U12866 (N_12866,N_11880,N_10221);
or U12867 (N_12867,N_11178,N_12266);
xnor U12868 (N_12868,N_10070,N_10094);
xnor U12869 (N_12869,N_10232,N_10104);
xor U12870 (N_12870,N_11126,N_12136);
nor U12871 (N_12871,N_11427,N_10361);
xor U12872 (N_12872,N_10724,N_10769);
xnor U12873 (N_12873,N_11925,N_11179);
nor U12874 (N_12874,N_11598,N_12497);
nand U12875 (N_12875,N_11602,N_10728);
and U12876 (N_12876,N_10690,N_10998);
nand U12877 (N_12877,N_11985,N_11036);
nor U12878 (N_12878,N_11404,N_10496);
nor U12879 (N_12879,N_10033,N_10034);
or U12880 (N_12880,N_10229,N_10727);
and U12881 (N_12881,N_12237,N_10400);
nand U12882 (N_12882,N_10475,N_11330);
nand U12883 (N_12883,N_10614,N_11038);
nand U12884 (N_12884,N_11839,N_10816);
or U12885 (N_12885,N_10838,N_11026);
or U12886 (N_12886,N_11102,N_11994);
nand U12887 (N_12887,N_10864,N_10714);
nor U12888 (N_12888,N_12276,N_10986);
nor U12889 (N_12889,N_11657,N_11477);
and U12890 (N_12890,N_11518,N_10373);
nand U12891 (N_12891,N_11372,N_10102);
xnor U12892 (N_12892,N_12120,N_11402);
nor U12893 (N_12893,N_12006,N_10649);
and U12894 (N_12894,N_11681,N_11288);
xor U12895 (N_12895,N_10510,N_10607);
nor U12896 (N_12896,N_10450,N_11325);
nand U12897 (N_12897,N_11650,N_12107);
nor U12898 (N_12898,N_11553,N_10054);
nand U12899 (N_12899,N_11855,N_11703);
nand U12900 (N_12900,N_12062,N_10663);
or U12901 (N_12901,N_10436,N_10684);
nand U12902 (N_12902,N_11762,N_10576);
nor U12903 (N_12903,N_10241,N_10564);
nand U12904 (N_12904,N_10116,N_11335);
and U12905 (N_12905,N_10533,N_10873);
and U12906 (N_12906,N_10506,N_10367);
xor U12907 (N_12907,N_12452,N_12498);
nor U12908 (N_12908,N_10477,N_12319);
nand U12909 (N_12909,N_12396,N_11207);
xor U12910 (N_12910,N_11736,N_10848);
xnor U12911 (N_12911,N_10353,N_11999);
xor U12912 (N_12912,N_11347,N_12468);
or U12913 (N_12913,N_11496,N_11263);
and U12914 (N_12914,N_12422,N_12066);
nand U12915 (N_12915,N_11919,N_11115);
nor U12916 (N_12916,N_10317,N_12114);
nor U12917 (N_12917,N_10949,N_10911);
nand U12918 (N_12918,N_10647,N_11538);
or U12919 (N_12919,N_12054,N_11802);
and U12920 (N_12920,N_11739,N_10783);
xor U12921 (N_12921,N_11433,N_10321);
nor U12922 (N_12922,N_11854,N_12168);
or U12923 (N_12923,N_11080,N_10561);
or U12924 (N_12924,N_11326,N_12213);
and U12925 (N_12925,N_10327,N_10636);
nor U12926 (N_12926,N_10174,N_10360);
or U12927 (N_12927,N_10206,N_11133);
or U12928 (N_12928,N_11387,N_10999);
and U12929 (N_12929,N_11396,N_11869);
xor U12930 (N_12930,N_10398,N_10235);
or U12931 (N_12931,N_11268,N_12032);
xnor U12932 (N_12932,N_10973,N_12309);
nand U12933 (N_12933,N_11807,N_11314);
xor U12934 (N_12934,N_12099,N_11244);
xor U12935 (N_12935,N_11593,N_10345);
and U12936 (N_12936,N_11670,N_10339);
xnor U12937 (N_12937,N_10817,N_11892);
nand U12938 (N_12938,N_10482,N_11811);
nand U12939 (N_12939,N_11742,N_11964);
nand U12940 (N_12940,N_11567,N_10430);
nor U12941 (N_12941,N_10788,N_11467);
xnor U12942 (N_12942,N_10680,N_11406);
or U12943 (N_12943,N_11849,N_10480);
nor U12944 (N_12944,N_10167,N_12162);
nor U12945 (N_12945,N_10265,N_10529);
and U12946 (N_12946,N_10084,N_11277);
and U12947 (N_12947,N_10987,N_11125);
or U12948 (N_12948,N_10976,N_10191);
nand U12949 (N_12949,N_10149,N_10256);
or U12950 (N_12950,N_10071,N_10320);
nor U12951 (N_12951,N_10947,N_11720);
nor U12952 (N_12952,N_11638,N_11063);
nand U12953 (N_12953,N_10741,N_10671);
xnor U12954 (N_12954,N_12178,N_10578);
nor U12955 (N_12955,N_11864,N_11311);
nor U12956 (N_12956,N_11318,N_12125);
nor U12957 (N_12957,N_11446,N_11788);
and U12958 (N_12958,N_11083,N_12366);
nor U12959 (N_12959,N_11111,N_12343);
xor U12960 (N_12960,N_11937,N_10691);
and U12961 (N_12961,N_10171,N_10250);
and U12962 (N_12962,N_12354,N_11479);
nor U12963 (N_12963,N_11459,N_11134);
or U12964 (N_12964,N_11209,N_11035);
and U12965 (N_12965,N_10503,N_11156);
and U12966 (N_12966,N_10648,N_12228);
nand U12967 (N_12967,N_10512,N_10261);
and U12968 (N_12968,N_11711,N_10114);
and U12969 (N_12969,N_10879,N_10654);
or U12970 (N_12970,N_12415,N_11995);
xor U12971 (N_12971,N_10757,N_12269);
or U12972 (N_12972,N_11570,N_11155);
nor U12973 (N_12973,N_11337,N_11581);
and U12974 (N_12974,N_11622,N_11551);
nor U12975 (N_12975,N_10784,N_11098);
xor U12976 (N_12976,N_10528,N_12474);
nor U12977 (N_12977,N_10917,N_10224);
xnor U12978 (N_12978,N_10301,N_12126);
or U12979 (N_12979,N_12101,N_11876);
and U12980 (N_12980,N_10097,N_11877);
or U12981 (N_12981,N_10922,N_10408);
or U12982 (N_12982,N_10726,N_12320);
nand U12983 (N_12983,N_12328,N_11095);
nor U12984 (N_12984,N_11239,N_11701);
nand U12985 (N_12985,N_11157,N_11262);
or U12986 (N_12986,N_12358,N_11214);
xor U12987 (N_12987,N_11576,N_12430);
and U12988 (N_12988,N_11405,N_11455);
and U12989 (N_12989,N_11977,N_12060);
nand U12990 (N_12990,N_10452,N_10722);
xor U12991 (N_12991,N_11113,N_11599);
nand U12992 (N_12992,N_11328,N_11525);
nand U12993 (N_12993,N_10939,N_10233);
xnor U12994 (N_12994,N_10347,N_12338);
or U12995 (N_12995,N_12472,N_12123);
nor U12996 (N_12996,N_10394,N_10900);
nor U12997 (N_12997,N_12056,N_10481);
or U12998 (N_12998,N_12231,N_10943);
nor U12999 (N_12999,N_11761,N_12247);
nor U13000 (N_13000,N_11659,N_11232);
or U13001 (N_13001,N_11845,N_10143);
and U13002 (N_13002,N_10615,N_11257);
xnor U13003 (N_13003,N_11355,N_10603);
xnor U13004 (N_13004,N_11047,N_10694);
xor U13005 (N_13005,N_10103,N_12466);
or U13006 (N_13006,N_11336,N_10777);
xnor U13007 (N_13007,N_11834,N_11279);
nor U13008 (N_13008,N_11090,N_11124);
xor U13009 (N_13009,N_11819,N_12344);
nand U13010 (N_13010,N_12191,N_10858);
and U13011 (N_13011,N_11689,N_10758);
nor U13012 (N_13012,N_11847,N_10336);
xor U13013 (N_13013,N_11117,N_10305);
and U13014 (N_13014,N_10796,N_11714);
and U13015 (N_13015,N_11829,N_11346);
and U13016 (N_13016,N_10285,N_10201);
or U13017 (N_13017,N_10523,N_10818);
and U13018 (N_13018,N_11700,N_10304);
nand U13019 (N_13019,N_10284,N_12073);
nand U13020 (N_13020,N_10729,N_12124);
nor U13021 (N_13021,N_10251,N_10209);
xor U13022 (N_13022,N_11984,N_11511);
nor U13023 (N_13023,N_11075,N_11667);
nand U13024 (N_13024,N_11103,N_10101);
nand U13025 (N_13025,N_12194,N_11127);
xor U13026 (N_13026,N_11559,N_10154);
nand U13027 (N_13027,N_10638,N_10751);
or U13028 (N_13028,N_10797,N_11192);
or U13029 (N_13029,N_10323,N_10124);
and U13030 (N_13030,N_10940,N_11835);
nand U13031 (N_13031,N_11630,N_10575);
xor U13032 (N_13032,N_10254,N_12386);
or U13033 (N_13033,N_11857,N_11749);
or U13034 (N_13034,N_11987,N_10342);
and U13035 (N_13035,N_10689,N_11163);
xnor U13036 (N_13036,N_10189,N_10027);
and U13037 (N_13037,N_10207,N_12360);
and U13038 (N_13038,N_11840,N_10925);
nand U13039 (N_13039,N_10082,N_12088);
nor U13040 (N_13040,N_10152,N_10723);
or U13041 (N_13041,N_11341,N_11046);
and U13042 (N_13042,N_10177,N_10828);
or U13043 (N_13043,N_11779,N_12221);
nand U13044 (N_13044,N_10421,N_12154);
xnor U13045 (N_13045,N_10554,N_10586);
or U13046 (N_13046,N_10288,N_10093);
nand U13047 (N_13047,N_10281,N_10773);
and U13048 (N_13048,N_11885,N_12195);
nand U13049 (N_13049,N_10202,N_11745);
xor U13050 (N_13050,N_12326,N_12405);
or U13051 (N_13051,N_10313,N_11501);
xor U13052 (N_13052,N_10010,N_10625);
nand U13053 (N_13053,N_11606,N_10025);
xnor U13054 (N_13054,N_10770,N_10793);
nor U13055 (N_13055,N_11685,N_12414);
xnor U13056 (N_13056,N_11924,N_12341);
and U13057 (N_13057,N_10966,N_12388);
nand U13058 (N_13058,N_12440,N_10110);
nor U13059 (N_13059,N_11349,N_10130);
nand U13060 (N_13060,N_10906,N_11472);
and U13061 (N_13061,N_10478,N_12286);
xor U13062 (N_13062,N_10606,N_10222);
xor U13063 (N_13063,N_11545,N_11361);
nor U13064 (N_13064,N_12175,N_11729);
and U13065 (N_13065,N_11777,N_11784);
and U13066 (N_13066,N_10859,N_12217);
nand U13067 (N_13067,N_11393,N_11089);
nor U13068 (N_13068,N_10282,N_11056);
nor U13069 (N_13069,N_11573,N_10963);
nor U13070 (N_13070,N_10933,N_10563);
nand U13071 (N_13071,N_10239,N_11916);
or U13072 (N_13072,N_10057,N_10882);
nand U13073 (N_13073,N_11099,N_12086);
or U13074 (N_13074,N_10144,N_10218);
nand U13075 (N_13075,N_10875,N_10753);
xnor U13076 (N_13076,N_11927,N_11733);
nor U13077 (N_13077,N_10880,N_10861);
nor U13078 (N_13078,N_10771,N_12325);
or U13079 (N_13079,N_12053,N_12059);
nand U13080 (N_13080,N_10619,N_11236);
or U13081 (N_13081,N_11493,N_12019);
and U13082 (N_13082,N_10168,N_11370);
or U13083 (N_13083,N_10137,N_12156);
nand U13084 (N_13084,N_10762,N_11447);
and U13085 (N_13085,N_11547,N_11261);
nor U13086 (N_13086,N_10799,N_10683);
and U13087 (N_13087,N_10835,N_12330);
nor U13088 (N_13088,N_11970,N_10532);
or U13089 (N_13089,N_11184,N_12431);
nand U13090 (N_13090,N_11710,N_11187);
xnor U13091 (N_13091,N_10451,N_12047);
nor U13092 (N_13092,N_10519,N_10735);
or U13093 (N_13093,N_10045,N_10573);
nor U13094 (N_13094,N_11054,N_11724);
nor U13095 (N_13095,N_11866,N_10822);
and U13096 (N_13096,N_11394,N_11267);
nand U13097 (N_13097,N_11148,N_11969);
and U13098 (N_13098,N_11392,N_11454);
xnor U13099 (N_13099,N_11023,N_10455);
nor U13100 (N_13100,N_10107,N_11176);
xnor U13101 (N_13101,N_10021,N_11716);
nand U13102 (N_13102,N_10932,N_11550);
nand U13103 (N_13103,N_12311,N_10213);
and U13104 (N_13104,N_10183,N_11058);
xor U13105 (N_13105,N_10161,N_12390);
and U13106 (N_13106,N_12305,N_11922);
nand U13107 (N_13107,N_11715,N_11853);
and U13108 (N_13108,N_11296,N_11458);
nor U13109 (N_13109,N_10934,N_10653);
nand U13110 (N_13110,N_10658,N_10464);
or U13111 (N_13111,N_10418,N_11933);
nor U13112 (N_13112,N_10064,N_10869);
nand U13113 (N_13113,N_11951,N_12476);
nor U13114 (N_13114,N_10673,N_10492);
or U13115 (N_13115,N_10589,N_11315);
or U13116 (N_13116,N_11658,N_11254);
and U13117 (N_13117,N_10065,N_10646);
and U13118 (N_13118,N_12241,N_10008);
and U13119 (N_13119,N_10092,N_10184);
xor U13120 (N_13120,N_11101,N_10705);
and U13121 (N_13121,N_12439,N_10299);
and U13122 (N_13122,N_11914,N_10095);
and U13123 (N_13123,N_10377,N_10626);
nor U13124 (N_13124,N_10789,N_10240);
and U13125 (N_13125,N_10359,N_12381);
or U13126 (N_13126,N_12190,N_10444);
xor U13127 (N_13127,N_11429,N_11146);
nand U13128 (N_13128,N_12014,N_12171);
and U13129 (N_13129,N_11037,N_10824);
nand U13130 (N_13130,N_11621,N_11500);
or U13131 (N_13131,N_10225,N_10410);
or U13132 (N_13132,N_10571,N_11012);
nand U13133 (N_13133,N_11440,N_12369);
nand U13134 (N_13134,N_11478,N_12376);
xor U13135 (N_13135,N_12287,N_10954);
xor U13136 (N_13136,N_12298,N_10538);
nand U13137 (N_13137,N_10135,N_12324);
xnor U13138 (N_13138,N_10696,N_10790);
and U13139 (N_13139,N_10597,N_11376);
nand U13140 (N_13140,N_11971,N_11137);
xnor U13141 (N_13141,N_12404,N_11813);
xnor U13142 (N_13142,N_10669,N_11609);
nor U13143 (N_13143,N_10083,N_11604);
or U13144 (N_13144,N_12093,N_11030);
or U13145 (N_13145,N_10136,N_11289);
nor U13146 (N_13146,N_12436,N_11595);
and U13147 (N_13147,N_11391,N_10036);
nand U13148 (N_13148,N_11758,N_10539);
nand U13149 (N_13149,N_11188,N_10196);
and U13150 (N_13150,N_12098,N_10682);
and U13151 (N_13151,N_10246,N_11331);
nor U13152 (N_13152,N_10839,N_12277);
nor U13153 (N_13153,N_10621,N_11862);
nand U13154 (N_13154,N_11530,N_10598);
and U13155 (N_13155,N_11734,N_12089);
and U13156 (N_13156,N_12179,N_12068);
xor U13157 (N_13157,N_12064,N_10248);
nor U13158 (N_13158,N_10314,N_10262);
and U13159 (N_13159,N_10547,N_10624);
and U13160 (N_13160,N_11614,N_12255);
xnor U13161 (N_13161,N_12112,N_12215);
xor U13162 (N_13162,N_10865,N_10959);
and U13163 (N_13163,N_11451,N_12159);
and U13164 (N_13164,N_11255,N_12478);
and U13165 (N_13165,N_11419,N_10787);
xnor U13166 (N_13166,N_12437,N_11794);
and U13167 (N_13167,N_12106,N_12167);
xor U13168 (N_13168,N_11837,N_11608);
nor U13169 (N_13169,N_10997,N_10836);
or U13170 (N_13170,N_10454,N_12134);
and U13171 (N_13171,N_11648,N_12397);
nand U13172 (N_13172,N_11975,N_12121);
xor U13173 (N_13173,N_11010,N_12482);
xnor U13174 (N_13174,N_11175,N_12248);
and U13175 (N_13175,N_11189,N_10173);
and U13176 (N_13176,N_10038,N_10545);
nor U13177 (N_13177,N_11804,N_10803);
nand U13178 (N_13178,N_12155,N_10810);
xor U13179 (N_13179,N_11757,N_10259);
nor U13180 (N_13180,N_10553,N_12481);
nand U13181 (N_13181,N_10420,N_11445);
or U13182 (N_13182,N_11119,N_11523);
xor U13183 (N_13183,N_11450,N_12058);
and U13184 (N_13184,N_10811,N_11695);
nand U13185 (N_13185,N_11350,N_10266);
nand U13186 (N_13186,N_10403,N_11235);
nand U13187 (N_13187,N_10318,N_12251);
nand U13188 (N_13188,N_10536,N_11850);
nand U13189 (N_13189,N_12016,N_12212);
or U13190 (N_13190,N_11342,N_10593);
and U13191 (N_13191,N_11698,N_10252);
and U13192 (N_13192,N_10381,N_10989);
or U13193 (N_13193,N_10018,N_10428);
nand U13194 (N_13194,N_10005,N_12046);
and U13195 (N_13195,N_12294,N_10983);
nand U13196 (N_13196,N_12132,N_11586);
or U13197 (N_13197,N_12382,N_11062);
nand U13198 (N_13198,N_11055,N_11150);
nor U13199 (N_13199,N_11443,N_11253);
xnor U13200 (N_13200,N_10069,N_12282);
xnor U13201 (N_13201,N_10910,N_12140);
nor U13202 (N_13202,N_10715,N_12378);
xnor U13203 (N_13203,N_10744,N_11180);
nor U13204 (N_13204,N_11147,N_10441);
and U13205 (N_13205,N_11222,N_10738);
and U13206 (N_13206,N_12072,N_11521);
nor U13207 (N_13207,N_10794,N_11278);
nand U13208 (N_13208,N_11334,N_10928);
nand U13209 (N_13209,N_12465,N_11923);
or U13210 (N_13210,N_11555,N_11677);
nand U13211 (N_13211,N_11270,N_11940);
xor U13212 (N_13212,N_11878,N_11365);
and U13213 (N_13213,N_12455,N_11580);
and U13214 (N_13214,N_11897,N_12094);
xnor U13215 (N_13215,N_12488,N_10891);
nand U13216 (N_13216,N_11221,N_10809);
and U13217 (N_13217,N_12185,N_12295);
and U13218 (N_13218,N_10214,N_11737);
or U13219 (N_13219,N_12127,N_10134);
and U13220 (N_13220,N_12223,N_10712);
nand U13221 (N_13221,N_10852,N_11386);
nor U13222 (N_13222,N_11563,N_11196);
or U13223 (N_13223,N_11796,N_10720);
and U13224 (N_13224,N_10594,N_12044);
nand U13225 (N_13225,N_10200,N_11616);
nand U13226 (N_13226,N_12301,N_11491);
and U13227 (N_13227,N_10483,N_11763);
nor U13228 (N_13228,N_11436,N_10007);
and U13229 (N_13229,N_12299,N_11653);
xnor U13230 (N_13230,N_10686,N_10277);
nand U13231 (N_13231,N_10550,N_10776);
or U13232 (N_13232,N_10424,N_10985);
or U13233 (N_13233,N_12027,N_10273);
nor U13234 (N_13234,N_11280,N_11662);
xnor U13235 (N_13235,N_10292,N_11549);
nor U13236 (N_13236,N_11215,N_12034);
nand U13237 (N_13237,N_12257,N_10466);
xnor U13238 (N_13238,N_11765,N_10674);
xor U13239 (N_13239,N_10815,N_10442);
and U13240 (N_13240,N_11162,N_10952);
xnor U13241 (N_13241,N_10075,N_10678);
or U13242 (N_13242,N_11627,N_11203);
and U13243 (N_13243,N_10219,N_12345);
or U13244 (N_13244,N_11043,N_10471);
nand U13245 (N_13245,N_11031,N_12029);
and U13246 (N_13246,N_10370,N_11513);
or U13247 (N_13247,N_10679,N_12158);
nor U13248 (N_13248,N_10074,N_12380);
nor U13249 (N_13249,N_12074,N_10060);
nand U13250 (N_13250,N_11771,N_10170);
xor U13251 (N_13251,N_10629,N_11204);
nor U13252 (N_13252,N_10307,N_11504);
and U13253 (N_13253,N_11212,N_11210);
and U13254 (N_13254,N_12253,N_11388);
nor U13255 (N_13255,N_12486,N_12456);
nand U13256 (N_13256,N_10672,N_11965);
and U13257 (N_13257,N_11833,N_10935);
or U13258 (N_13258,N_11073,N_11680);
xor U13259 (N_13259,N_10874,N_12004);
and U13260 (N_13260,N_12033,N_10950);
nand U13261 (N_13261,N_10402,N_11503);
nand U13262 (N_13262,N_10856,N_12031);
or U13263 (N_13263,N_10732,N_10399);
and U13264 (N_13264,N_11061,N_11906);
nor U13265 (N_13265,N_11556,N_11875);
xor U13266 (N_13266,N_10840,N_10644);
and U13267 (N_13267,N_10278,N_12296);
nand U13268 (N_13268,N_10708,N_11316);
nor U13269 (N_13269,N_11528,N_10552);
xnor U13270 (N_13270,N_11259,N_10309);
and U13271 (N_13271,N_10641,N_11823);
and U13272 (N_13272,N_10100,N_11421);
nand U13273 (N_13273,N_11486,N_10178);
or U13274 (N_13274,N_12271,N_12362);
and U13275 (N_13275,N_12417,N_12399);
nand U13276 (N_13276,N_10208,N_10058);
xnor U13277 (N_13277,N_10534,N_10303);
nor U13278 (N_13278,N_12406,N_11721);
xor U13279 (N_13279,N_10341,N_11422);
nand U13280 (N_13280,N_11799,N_11688);
or U13281 (N_13281,N_10325,N_10591);
and U13282 (N_13282,N_11699,N_11645);
or U13283 (N_13283,N_10169,N_11007);
or U13284 (N_13284,N_10460,N_10212);
xor U13285 (N_13285,N_11273,N_10404);
nand U13286 (N_13286,N_11247,N_11982);
or U13287 (N_13287,N_10667,N_10778);
and U13288 (N_13288,N_11497,N_12115);
or U13289 (N_13289,N_11886,N_12263);
xnor U13290 (N_13290,N_11967,N_10566);
or U13291 (N_13291,N_12077,N_11718);
nand U13292 (N_13292,N_11021,N_11067);
nand U13293 (N_13293,N_11561,N_10260);
and U13294 (N_13294,N_11836,N_12013);
and U13295 (N_13295,N_12487,N_11008);
nand U13296 (N_13296,N_11322,N_11672);
nor U13297 (N_13297,N_10050,N_11005);
and U13298 (N_13298,N_11202,N_11536);
or U13299 (N_13299,N_10365,N_12314);
or U13300 (N_13300,N_11449,N_12216);
nor U13301 (N_13301,N_11002,N_10502);
nor U13302 (N_13302,N_10524,N_12070);
nand U13303 (N_13303,N_10710,N_10389);
nand U13304 (N_13304,N_10982,N_10884);
nand U13305 (N_13305,N_10279,N_10293);
nand U13306 (N_13306,N_10096,N_10499);
nand U13307 (N_13307,N_10227,N_10470);
nor U13308 (N_13308,N_10842,N_10665);
nor U13309 (N_13309,N_10588,N_10945);
or U13310 (N_13310,N_10199,N_11407);
nand U13311 (N_13311,N_11498,N_10944);
or U13312 (N_13312,N_11234,N_12264);
xor U13313 (N_13313,N_10486,N_11909);
or U13314 (N_13314,N_11437,N_10179);
and U13315 (N_13315,N_10927,N_10870);
and U13316 (N_13316,N_11851,N_10446);
or U13317 (N_13317,N_11293,N_12339);
nand U13318 (N_13318,N_11983,N_11237);
and U13319 (N_13319,N_12280,N_11481);
nand U13320 (N_13320,N_10405,N_12078);
or U13321 (N_13321,N_10542,N_11583);
or U13322 (N_13322,N_10747,N_11810);
or U13323 (N_13323,N_11024,N_11958);
nand U13324 (N_13324,N_10800,N_10126);
or U13325 (N_13325,N_10162,N_10711);
nand U13326 (N_13326,N_11986,N_12015);
xnor U13327 (N_13327,N_10395,N_10264);
nor U13328 (N_13328,N_12161,N_10888);
nor U13329 (N_13329,N_12451,N_10253);
nor U13330 (N_13330,N_11462,N_10041);
nor U13331 (N_13331,N_11442,N_10548);
or U13332 (N_13332,N_10652,N_12394);
nand U13333 (N_13333,N_10139,N_11938);
nor U13334 (N_13334,N_10780,N_10090);
nand U13335 (N_13335,N_11543,N_11664);
or U13336 (N_13336,N_10604,N_11430);
and U13337 (N_13337,N_11208,N_10422);
xor U13338 (N_13338,N_10223,N_10188);
nand U13339 (N_13339,N_12243,N_12189);
nand U13340 (N_13340,N_11712,N_10129);
xor U13341 (N_13341,N_11390,N_12035);
or U13342 (N_13342,N_11367,N_10677);
nand U13343 (N_13343,N_12103,N_11057);
nand U13344 (N_13344,N_11774,N_10024);
nand U13345 (N_13345,N_10147,N_10427);
xor U13346 (N_13346,N_10330,N_10433);
nand U13347 (N_13347,N_12000,N_11615);
xnor U13348 (N_13348,N_12418,N_12096);
nand U13349 (N_13349,N_12144,N_11678);
xnor U13350 (N_13350,N_11494,N_12300);
or U13351 (N_13351,N_12095,N_11824);
nor U13352 (N_13352,N_11950,N_10759);
and U13353 (N_13353,N_11704,N_10456);
or U13354 (N_13354,N_10472,N_12119);
or U13355 (N_13355,N_10371,N_12454);
or U13356 (N_13356,N_11805,N_11120);
xor U13357 (N_13357,N_10247,N_11468);
xnor U13358 (N_13358,N_11049,N_10332);
xnor U13359 (N_13359,N_11465,N_12475);
or U13360 (N_13360,N_11747,N_11258);
nor U13361 (N_13361,N_11242,N_11644);
and U13362 (N_13362,N_12383,N_10302);
and U13363 (N_13363,N_11679,N_11767);
xnor U13364 (N_13364,N_12079,N_10693);
xnor U13365 (N_13365,N_11646,N_10993);
or U13366 (N_13366,N_12395,N_11197);
or U13367 (N_13367,N_11274,N_11642);
or U13368 (N_13368,N_11333,N_11997);
nand U13369 (N_13369,N_10385,N_11693);
nor U13370 (N_13370,N_11135,N_12235);
nand U13371 (N_13371,N_12025,N_10562);
and U13372 (N_13372,N_11358,N_11694);
and U13373 (N_13373,N_10745,N_12416);
xor U13374 (N_13374,N_11859,N_10319);
nor U13375 (N_13375,N_10028,N_11565);
nor U13376 (N_13376,N_10237,N_11652);
or U13377 (N_13377,N_10121,N_11389);
nand U13378 (N_13378,N_12091,N_10704);
nand U13379 (N_13379,N_11798,N_12318);
xor U13380 (N_13380,N_10681,N_10544);
xor U13381 (N_13381,N_10918,N_11480);
or U13382 (N_13382,N_10511,N_11781);
nor U13383 (N_13383,N_10489,N_11655);
xor U13384 (N_13384,N_11508,N_11979);
or U13385 (N_13385,N_12496,N_11110);
or U13386 (N_13386,N_12293,N_11564);
and U13387 (N_13387,N_11773,N_12332);
or U13388 (N_13388,N_10637,N_12377);
nor U13389 (N_13389,N_12108,N_10749);
and U13390 (N_13390,N_10992,N_11364);
nor U13391 (N_13391,N_12039,N_10287);
or U13392 (N_13392,N_10650,N_10830);
nand U13393 (N_13393,N_11752,N_10965);
and U13394 (N_13394,N_11904,N_11033);
xnor U13395 (N_13395,N_11434,N_10956);
nand U13396 (N_13396,N_10814,N_11684);
xnor U13397 (N_13397,N_11649,N_10032);
or U13398 (N_13398,N_10651,N_11077);
and U13399 (N_13399,N_12110,N_11299);
xor U13400 (N_13400,N_12232,N_10192);
xnor U13401 (N_13401,N_10984,N_12245);
or U13402 (N_13402,N_10270,N_12450);
nor U13403 (N_13403,N_10042,N_10115);
and U13404 (N_13404,N_11431,N_10565);
or U13405 (N_13405,N_11585,N_12193);
nand U13406 (N_13406,N_11557,N_10608);
nor U13407 (N_13407,N_12163,N_11423);
or U13408 (N_13408,N_10412,N_11357);
or U13409 (N_13409,N_10863,N_10459);
nand U13410 (N_13410,N_11123,N_12200);
nor U13411 (N_13411,N_10350,N_10158);
or U13412 (N_13412,N_12315,N_10236);
and U13413 (N_13413,N_10707,N_12479);
or U13414 (N_13414,N_10306,N_10378);
or U13415 (N_13415,N_11377,N_10926);
xor U13416 (N_13416,N_12238,N_10376);
and U13417 (N_13417,N_11295,N_11457);
nand U13418 (N_13418,N_11425,N_11074);
nand U13419 (N_13419,N_11792,N_11888);
nor U13420 (N_13420,N_11444,N_11990);
xnor U13421 (N_13421,N_10002,N_11603);
nor U13422 (N_13422,N_10276,N_10298);
or U13423 (N_13423,N_10138,N_10853);
nand U13424 (N_13424,N_11383,N_11013);
xnor U13425 (N_13425,N_11471,N_11682);
and U13426 (N_13426,N_10721,N_11808);
nor U13427 (N_13427,N_10343,N_10955);
xor U13428 (N_13428,N_10210,N_12283);
or U13429 (N_13429,N_11460,N_10458);
and U13430 (N_13430,N_12075,N_10255);
nand U13431 (N_13431,N_10834,N_10495);
or U13432 (N_13432,N_12262,N_11004);
and U13433 (N_13433,N_10346,N_11287);
nand U13434 (N_13434,N_12183,N_11438);
or U13435 (N_13435,N_11348,N_10328);
and U13436 (N_13436,N_10580,N_12274);
nand U13437 (N_13437,N_10172,N_10081);
xnor U13438 (N_13438,N_11107,N_10946);
xor U13439 (N_13439,N_11582,N_11164);
nand U13440 (N_13440,N_11626,N_12113);
or U13441 (N_13441,N_11017,N_11078);
nand U13442 (N_13442,N_11453,N_11343);
and U13443 (N_13443,N_11620,N_11643);
xnor U13444 (N_13444,N_11304,N_11988);
nand U13445 (N_13445,N_10504,N_11526);
nor U13446 (N_13446,N_11917,N_10821);
nand U13447 (N_13447,N_11717,N_11780);
and U13448 (N_13448,N_10156,N_10245);
and U13449 (N_13449,N_12208,N_11371);
and U13450 (N_13450,N_11432,N_12085);
xnor U13451 (N_13451,N_10372,N_12402);
xor U13452 (N_13452,N_11822,N_10448);
and U13453 (N_13453,N_10474,N_10920);
or U13454 (N_13454,N_11312,N_10443);
nor U13455 (N_13455,N_10465,N_11401);
or U13456 (N_13456,N_11740,N_11673);
nor U13457 (N_13457,N_11476,N_10713);
nand U13458 (N_13458,N_12321,N_10618);
xor U13459 (N_13459,N_11948,N_10823);
xnor U13460 (N_13460,N_11019,N_12219);
nand U13461 (N_13461,N_12278,N_12061);
nor U13462 (N_13462,N_11165,N_10413);
and U13463 (N_13463,N_10164,N_10801);
nand U13464 (N_13464,N_10743,N_10150);
and U13465 (N_13465,N_11116,N_11949);
nand U13466 (N_13466,N_10331,N_10392);
xnor U13467 (N_13467,N_10775,N_10358);
nor U13468 (N_13468,N_11534,N_12111);
or U13469 (N_13469,N_11050,N_11097);
xor U13470 (N_13470,N_11791,N_11149);
nor U13471 (N_13471,N_11935,N_10078);
xor U13472 (N_13472,N_10622,N_10688);
xor U13473 (N_13473,N_11139,N_12333);
or U13474 (N_13474,N_11532,N_12448);
or U13475 (N_13475,N_10257,N_12375);
or U13476 (N_13476,N_11340,N_10558);
or U13477 (N_13477,N_11956,N_12491);
nand U13478 (N_13478,N_12469,N_10572);
xnor U13479 (N_13479,N_11568,N_10390);
or U13480 (N_13480,N_11991,N_12433);
nor U13481 (N_13481,N_11863,N_10703);
and U13482 (N_13482,N_10366,N_11034);
or U13483 (N_13483,N_10022,N_10509);
or U13484 (N_13484,N_11973,N_11635);
xor U13485 (N_13485,N_10242,N_10498);
nand U13486 (N_13486,N_12142,N_10948);
nand U13487 (N_13487,N_12229,N_11051);
nor U13488 (N_13488,N_10957,N_10079);
nor U13489 (N_13489,N_12160,N_10871);
and U13490 (N_13490,N_12172,N_11015);
xor U13491 (N_13491,N_11920,N_11490);
nor U13492 (N_13492,N_11507,N_12174);
xor U13493 (N_13493,N_12188,N_11233);
and U13494 (N_13494,N_10893,N_12365);
nand U13495 (N_13495,N_11946,N_10700);
xor U13496 (N_13496,N_10030,N_10349);
xnor U13497 (N_13497,N_11768,N_10283);
and U13498 (N_13498,N_10052,N_11068);
nor U13499 (N_13499,N_12370,N_11298);
nand U13500 (N_13500,N_11252,N_11778);
nand U13501 (N_13501,N_12357,N_11260);
xor U13502 (N_13502,N_11953,N_10185);
xor U13503 (N_13503,N_12429,N_12157);
xor U13504 (N_13504,N_12065,N_11516);
nor U13505 (N_13505,N_12100,N_11413);
nand U13506 (N_13506,N_10530,N_10905);
nand U13507 (N_13507,N_12026,N_10845);
nor U13508 (N_13508,N_11591,N_10921);
nand U13509 (N_13509,N_12227,N_11292);
and U13510 (N_13510,N_10003,N_12470);
or U13511 (N_13511,N_11535,N_12105);
xnor U13512 (N_13512,N_11167,N_11220);
and U13513 (N_13513,N_12389,N_12104);
nand U13514 (N_13514,N_10468,N_10039);
nor U13515 (N_13515,N_10019,N_12197);
and U13516 (N_13516,N_11870,N_11020);
and U13517 (N_13517,N_10610,N_11485);
nor U13518 (N_13518,N_11249,N_12002);
nand U13519 (N_13519,N_10354,N_10967);
and U13520 (N_13520,N_11572,N_10006);
xnor U13521 (N_13521,N_10697,N_10570);
xnor U13522 (N_13522,N_10979,N_10602);
and U13523 (N_13523,N_11297,N_10725);
xor U13524 (N_13524,N_11912,N_11706);
or U13525 (N_13525,N_11654,N_11173);
and U13526 (N_13526,N_12203,N_11052);
nand U13527 (N_13527,N_10203,N_11082);
and U13528 (N_13528,N_12204,N_11439);
and U13529 (N_13529,N_10929,N_10357);
xnor U13530 (N_13530,N_12051,N_10779);
nor U13531 (N_13531,N_10675,N_11379);
nor U13532 (N_13532,N_10362,N_12323);
nor U13533 (N_13533,N_11908,N_10639);
nand U13534 (N_13534,N_11122,N_12489);
nor U13535 (N_13535,N_10868,N_10447);
nand U13536 (N_13536,N_10766,N_11041);
xnor U13537 (N_13537,N_11981,N_12421);
and U13538 (N_13538,N_11369,N_11131);
nor U13539 (N_13539,N_11435,N_12214);
nand U13540 (N_13540,N_11290,N_10887);
xnor U13541 (N_13541,N_10851,N_10132);
nor U13542 (N_13542,N_10300,N_10692);
xnor U13543 (N_13543,N_11590,N_10746);
or U13544 (N_13544,N_11756,N_11746);
and U13545 (N_13545,N_12116,N_11989);
xnor U13546 (N_13546,N_11558,N_10231);
nor U13547 (N_13547,N_10120,N_11426);
xor U13548 (N_13548,N_12239,N_12076);
or U13549 (N_13549,N_11993,N_10731);
xor U13550 (N_13550,N_12379,N_11738);
nand U13551 (N_13551,N_10106,N_10063);
nor U13552 (N_13552,N_10627,N_10881);
or U13553 (N_13553,N_12071,N_11138);
or U13554 (N_13554,N_10023,N_12410);
or U13555 (N_13555,N_10866,N_11487);
nand U13556 (N_13556,N_11306,N_12483);
or U13557 (N_13557,N_12092,N_10964);
nor U13558 (N_13558,N_10217,N_10500);
xnor U13559 (N_13559,N_11931,N_10531);
xor U13560 (N_13560,N_11181,N_11283);
and U13561 (N_13561,N_11783,N_10001);
nand U13562 (N_13562,N_12202,N_11161);
xnor U13563 (N_13563,N_11100,N_11040);
nand U13564 (N_13564,N_10211,N_11980);
and U13565 (N_13565,N_11417,N_11108);
or U13566 (N_13566,N_11628,N_11093);
or U13567 (N_13567,N_11448,N_12460);
or U13568 (N_13568,N_12493,N_11362);
xnor U13569 (N_13569,N_10140,N_11597);
nor U13570 (N_13570,N_10113,N_11723);
nor U13571 (N_13571,N_10190,N_12052);
and U13572 (N_13572,N_11753,N_10216);
xor U13573 (N_13573,N_11354,N_11697);
or U13574 (N_13574,N_10774,N_11669);
and U13575 (N_13575,N_12122,N_12149);
xor U13576 (N_13576,N_10628,N_10813);
xor U13577 (N_13577,N_11826,N_11611);
nor U13578 (N_13578,N_10091,N_11820);
nand U13579 (N_13579,N_11081,N_10294);
and U13580 (N_13580,N_12082,N_11754);
nand U13581 (N_13581,N_10086,N_12097);
or U13582 (N_13582,N_12398,N_10978);
nand U13583 (N_13583,N_10355,N_11420);
and U13584 (N_13584,N_10180,N_12356);
and U13585 (N_13585,N_10737,N_11408);
nor U13586 (N_13586,N_12143,N_11071);
and U13587 (N_13587,N_12348,N_10792);
nand U13588 (N_13588,N_10268,N_11944);
or U13589 (N_13589,N_12012,N_11483);
xor U13590 (N_13590,N_11329,N_11522);
or U13591 (N_13591,N_12368,N_11775);
nor U13592 (N_13592,N_10924,N_11229);
xnor U13593 (N_13593,N_10414,N_10274);
or U13594 (N_13594,N_10895,N_12177);
nand U13595 (N_13595,N_11686,N_10437);
nor U13596 (N_13596,N_10297,N_12234);
nand U13597 (N_13597,N_11647,N_11540);
nand U13598 (N_13598,N_10068,N_12055);
nand U13599 (N_13599,N_10827,N_12302);
nand U13600 (N_13600,N_12322,N_11619);
nor U13601 (N_13601,N_11403,N_11170);
nor U13602 (N_13602,N_11961,N_10768);
nor U13603 (N_13603,N_10098,N_10640);
or U13604 (N_13604,N_12392,N_10133);
or U13605 (N_13605,N_10004,N_12133);
or U13606 (N_13606,N_10913,N_11039);
nand U13607 (N_13607,N_12080,N_10919);
or U13608 (N_13608,N_10128,N_10364);
and U13609 (N_13609,N_11911,N_12201);
nand U13610 (N_13610,N_11790,N_12137);
and U13611 (N_13611,N_12285,N_10837);
and U13612 (N_13612,N_10425,N_11519);
nand U13613 (N_13613,N_10085,N_11891);
or U13614 (N_13614,N_10435,N_12359);
nor U13615 (N_13615,N_10396,N_11800);
xnor U13616 (N_13616,N_12453,N_10662);
nand U13617 (N_13617,N_10786,N_11201);
or U13618 (N_13618,N_10634,N_11169);
nor U13619 (N_13619,N_10695,N_10344);
xnor U13620 (N_13620,N_10310,N_11852);
and U13621 (N_13621,N_11353,N_11177);
nand U13622 (N_13622,N_11865,N_10432);
and U13623 (N_13623,N_10522,N_11373);
or U13624 (N_13624,N_12384,N_12409);
and U13625 (N_13625,N_10015,N_12242);
or U13626 (N_13626,N_12117,N_12244);
xor U13627 (N_13627,N_10204,N_12424);
nor U13628 (N_13628,N_11205,N_10088);
nor U13629 (N_13629,N_12273,N_12005);
xnor U13630 (N_13630,N_10215,N_11719);
xnor U13631 (N_13631,N_12040,N_11601);
xnor U13632 (N_13632,N_11231,N_10831);
nor U13633 (N_13633,N_11225,N_12306);
nor U13634 (N_13634,N_10333,N_10960);
nor U13635 (N_13635,N_11996,N_10334);
nand U13636 (N_13636,N_12413,N_10764);
nor U13637 (N_13637,N_11313,N_11748);
xnor U13638 (N_13638,N_10047,N_11248);
xnor U13639 (N_13639,N_10748,N_11129);
nor U13640 (N_13640,N_11910,N_12317);
nand U13641 (N_13641,N_10781,N_10574);
and U13642 (N_13642,N_10668,N_12207);
nor U13643 (N_13643,N_11356,N_11634);
xnor U13644 (N_13644,N_11506,N_10825);
and U13645 (N_13645,N_11199,N_10340);
and U13646 (N_13646,N_11656,N_11284);
nor U13647 (N_13647,N_10387,N_11691);
or U13648 (N_13648,N_11881,N_11065);
nor U13649 (N_13649,N_11198,N_11213);
nor U13650 (N_13650,N_12313,N_11085);
nor U13651 (N_13651,N_11867,N_11743);
or U13652 (N_13652,N_10228,N_10915);
and U13653 (N_13653,N_12184,N_11872);
nand U13654 (N_13654,N_12081,N_12102);
nand U13655 (N_13655,N_11651,N_10012);
and U13656 (N_13656,N_10990,N_10826);
nand U13657 (N_13657,N_12400,N_12367);
xor U13658 (N_13658,N_12041,N_11344);
nor U13659 (N_13659,N_12290,N_11772);
xnor U13660 (N_13660,N_10756,N_12186);
nor U13661 (N_13661,N_10125,N_11305);
or U13662 (N_13662,N_12442,N_11882);
nor U13663 (N_13663,N_11368,N_10051);
nor U13664 (N_13664,N_10198,N_12182);
xnor U13665 (N_13665,N_12426,N_11921);
or U13666 (N_13666,N_10151,N_10338);
nand U13667 (N_13667,N_10659,N_10440);
and U13668 (N_13668,N_11751,N_10515);
and U13669 (N_13669,N_10620,N_12425);
and U13670 (N_13670,N_12030,N_11474);
and U13671 (N_13671,N_10847,N_10348);
and U13672 (N_13672,N_12084,N_11482);
nor U13673 (N_13673,N_12261,N_11832);
xor U13674 (N_13674,N_11217,N_11484);
nand U13675 (N_13675,N_11776,N_10067);
nand U13676 (N_13676,N_10660,N_10518);
nor U13677 (N_13677,N_12461,N_11896);
nand U13678 (N_13678,N_10463,N_10230);
xor U13679 (N_13679,N_11960,N_11276);
nand U13680 (N_13680,N_11594,N_11731);
xnor U13681 (N_13681,N_11873,N_11636);
nor U13682 (N_13682,N_11786,N_12209);
nor U13683 (N_13683,N_11086,N_12028);
nand U13684 (N_13684,N_10896,N_10645);
nand U13685 (N_13685,N_10857,N_11025);
nand U13686 (N_13686,N_10767,N_10701);
nand U13687 (N_13687,N_11319,N_10656);
nand U13688 (N_13688,N_12291,N_11028);
or U13689 (N_13689,N_10491,N_10630);
and U13690 (N_13690,N_10123,N_10555);
and U13691 (N_13691,N_11809,N_10379);
nor U13692 (N_13692,N_12049,N_11945);
nor U13693 (N_13693,N_10912,N_10537);
or U13694 (N_13694,N_12446,N_10099);
nor U13695 (N_13695,N_12135,N_10765);
nor U13696 (N_13696,N_10802,N_10867);
nand U13697 (N_13697,N_10289,N_12173);
and U13698 (N_13698,N_11141,N_11003);
xnor U13699 (N_13699,N_11546,N_12346);
nor U13700 (N_13700,N_11363,N_10112);
nor U13701 (N_13701,N_11816,N_12083);
nor U13702 (N_13702,N_11730,N_12153);
nand U13703 (N_13703,N_10655,N_12036);
xor U13704 (N_13704,N_10234,N_10397);
nand U13705 (N_13705,N_12335,N_11060);
nor U13706 (N_13706,N_11271,N_11029);
nor U13707 (N_13707,N_10601,N_11898);
and U13708 (N_13708,N_12260,N_11605);
nand U13709 (N_13709,N_12374,N_10899);
and U13710 (N_13710,N_10883,N_11879);
xor U13711 (N_13711,N_11610,N_11193);
and U13712 (N_13712,N_11303,N_12220);
and U13713 (N_13713,N_10401,N_10849);
nand U13714 (N_13714,N_10488,N_11018);
nand U13715 (N_13715,N_10312,N_10995);
and U13716 (N_13716,N_10904,N_10844);
xnor U13717 (N_13717,N_10909,N_12484);
xnor U13718 (N_13718,N_12407,N_10040);
xnor U13719 (N_13719,N_10316,N_12420);
or U13720 (N_13720,N_10698,N_10595);
xor U13721 (N_13721,N_11332,N_12045);
nand U13722 (N_13722,N_11183,N_11105);
nor U13723 (N_13723,N_10205,N_12351);
and U13724 (N_13724,N_11092,N_12312);
or U13725 (N_13725,N_10186,N_10890);
and U13726 (N_13726,N_12176,N_12146);
xnor U13727 (N_13727,N_10393,N_11705);
nand U13728 (N_13728,N_10073,N_10908);
nor U13729 (N_13729,N_11190,N_11409);
or U13730 (N_13730,N_12310,N_12043);
and U13731 (N_13731,N_10382,N_10220);
nand U13732 (N_13732,N_10419,N_11542);
nor U13733 (N_13733,N_11726,N_11502);
nor U13734 (N_13734,N_10473,N_12011);
and U13735 (N_13735,N_10275,N_11265);
xnor U13736 (N_13736,N_10374,N_10772);
nor U13737 (N_13737,N_12438,N_11510);
or U13738 (N_13738,N_10296,N_10974);
or U13739 (N_13739,N_11410,N_12254);
or U13740 (N_13740,N_11934,N_10930);
nand U13741 (N_13741,N_10062,N_10011);
or U13742 (N_13742,N_10785,N_11548);
and U13743 (N_13743,N_11841,N_11418);
and U13744 (N_13744,N_12265,N_10386);
and U13745 (N_13745,N_11112,N_10739);
xnor U13746 (N_13746,N_12230,N_10605);
xor U13747 (N_13747,N_12090,N_11194);
xnor U13748 (N_13748,N_11087,N_10546);
and U13749 (N_13749,N_11452,N_10243);
or U13750 (N_13750,N_10778,N_10910);
nand U13751 (N_13751,N_11201,N_11039);
xor U13752 (N_13752,N_11304,N_12233);
or U13753 (N_13753,N_12352,N_10544);
xor U13754 (N_13754,N_11428,N_12260);
nor U13755 (N_13755,N_10336,N_10964);
nor U13756 (N_13756,N_10761,N_10936);
or U13757 (N_13757,N_11128,N_11732);
nand U13758 (N_13758,N_12012,N_11686);
and U13759 (N_13759,N_10528,N_12302);
and U13760 (N_13760,N_11794,N_11330);
and U13761 (N_13761,N_10764,N_11419);
nor U13762 (N_13762,N_11549,N_11172);
nand U13763 (N_13763,N_10566,N_11026);
or U13764 (N_13764,N_11440,N_10140);
xnor U13765 (N_13765,N_10114,N_11966);
xor U13766 (N_13766,N_10435,N_10964);
nor U13767 (N_13767,N_10006,N_10579);
xor U13768 (N_13768,N_10295,N_10700);
and U13769 (N_13769,N_11247,N_10454);
xnor U13770 (N_13770,N_11992,N_12198);
nor U13771 (N_13771,N_10140,N_11536);
and U13772 (N_13772,N_11474,N_10746);
or U13773 (N_13773,N_10492,N_12357);
or U13774 (N_13774,N_12182,N_10117);
or U13775 (N_13775,N_10616,N_10006);
and U13776 (N_13776,N_10172,N_12289);
xor U13777 (N_13777,N_11990,N_10156);
xnor U13778 (N_13778,N_10516,N_10252);
nor U13779 (N_13779,N_10556,N_11581);
xnor U13780 (N_13780,N_12226,N_12188);
nor U13781 (N_13781,N_11495,N_10173);
and U13782 (N_13782,N_10945,N_12138);
nor U13783 (N_13783,N_11354,N_11331);
and U13784 (N_13784,N_11034,N_10288);
and U13785 (N_13785,N_11639,N_11610);
and U13786 (N_13786,N_11248,N_10820);
and U13787 (N_13787,N_10141,N_12107);
and U13788 (N_13788,N_10392,N_12090);
or U13789 (N_13789,N_11503,N_10289);
nor U13790 (N_13790,N_10730,N_12148);
nand U13791 (N_13791,N_10536,N_10273);
xnor U13792 (N_13792,N_12317,N_11143);
or U13793 (N_13793,N_12070,N_11553);
or U13794 (N_13794,N_12493,N_11798);
or U13795 (N_13795,N_12373,N_10461);
nor U13796 (N_13796,N_11021,N_10510);
or U13797 (N_13797,N_11421,N_10756);
nand U13798 (N_13798,N_11935,N_12272);
xor U13799 (N_13799,N_11762,N_11493);
nor U13800 (N_13800,N_11306,N_12084);
xor U13801 (N_13801,N_12106,N_11988);
xor U13802 (N_13802,N_10796,N_10322);
or U13803 (N_13803,N_11704,N_10557);
and U13804 (N_13804,N_10763,N_11401);
or U13805 (N_13805,N_11519,N_11075);
or U13806 (N_13806,N_11310,N_10069);
nand U13807 (N_13807,N_11096,N_12268);
nor U13808 (N_13808,N_11499,N_11552);
or U13809 (N_13809,N_10103,N_11594);
or U13810 (N_13810,N_10973,N_10077);
and U13811 (N_13811,N_11830,N_11954);
and U13812 (N_13812,N_10044,N_10947);
xor U13813 (N_13813,N_11212,N_10467);
nor U13814 (N_13814,N_10221,N_12227);
xnor U13815 (N_13815,N_11631,N_11629);
and U13816 (N_13816,N_11772,N_11166);
nand U13817 (N_13817,N_11132,N_12139);
or U13818 (N_13818,N_12033,N_11466);
or U13819 (N_13819,N_12414,N_10116);
or U13820 (N_13820,N_10235,N_12387);
nor U13821 (N_13821,N_12010,N_11162);
xor U13822 (N_13822,N_10030,N_10769);
nor U13823 (N_13823,N_10337,N_10827);
nand U13824 (N_13824,N_10903,N_10371);
xnor U13825 (N_13825,N_11368,N_12243);
and U13826 (N_13826,N_10006,N_11935);
nor U13827 (N_13827,N_11915,N_10241);
xor U13828 (N_13828,N_12187,N_10298);
xor U13829 (N_13829,N_12273,N_10753);
nand U13830 (N_13830,N_10031,N_11132);
and U13831 (N_13831,N_10562,N_11380);
nor U13832 (N_13832,N_11812,N_11100);
and U13833 (N_13833,N_11601,N_10898);
or U13834 (N_13834,N_12092,N_11398);
xor U13835 (N_13835,N_10166,N_10616);
xnor U13836 (N_13836,N_11052,N_10903);
and U13837 (N_13837,N_11905,N_10247);
and U13838 (N_13838,N_10326,N_11001);
and U13839 (N_13839,N_11219,N_11627);
and U13840 (N_13840,N_11658,N_11445);
nor U13841 (N_13841,N_12087,N_11441);
xnor U13842 (N_13842,N_11169,N_12296);
or U13843 (N_13843,N_12076,N_10329);
xor U13844 (N_13844,N_10143,N_12142);
nand U13845 (N_13845,N_11307,N_10090);
nor U13846 (N_13846,N_12425,N_10355);
nand U13847 (N_13847,N_11159,N_10401);
and U13848 (N_13848,N_10345,N_11411);
nor U13849 (N_13849,N_12344,N_10837);
or U13850 (N_13850,N_10687,N_11451);
nand U13851 (N_13851,N_10274,N_11031);
nand U13852 (N_13852,N_11708,N_11849);
xor U13853 (N_13853,N_12470,N_11579);
xor U13854 (N_13854,N_10894,N_10450);
nor U13855 (N_13855,N_11469,N_10798);
xnor U13856 (N_13856,N_11914,N_11704);
nor U13857 (N_13857,N_11131,N_10783);
or U13858 (N_13858,N_11764,N_10153);
xor U13859 (N_13859,N_10142,N_11650);
xor U13860 (N_13860,N_10245,N_12084);
nor U13861 (N_13861,N_12406,N_10902);
xnor U13862 (N_13862,N_11951,N_12336);
xor U13863 (N_13863,N_12451,N_12213);
xnor U13864 (N_13864,N_11704,N_10227);
or U13865 (N_13865,N_10434,N_11637);
nand U13866 (N_13866,N_10060,N_12206);
and U13867 (N_13867,N_10503,N_12088);
or U13868 (N_13868,N_11132,N_10369);
xnor U13869 (N_13869,N_12205,N_12169);
nor U13870 (N_13870,N_10122,N_10974);
nor U13871 (N_13871,N_12048,N_10466);
nand U13872 (N_13872,N_11745,N_10191);
nor U13873 (N_13873,N_10774,N_10622);
nand U13874 (N_13874,N_11505,N_10755);
nand U13875 (N_13875,N_11299,N_11075);
nor U13876 (N_13876,N_11512,N_12131);
nor U13877 (N_13877,N_11329,N_10708);
or U13878 (N_13878,N_10917,N_10247);
or U13879 (N_13879,N_10210,N_10778);
nand U13880 (N_13880,N_11837,N_12192);
xor U13881 (N_13881,N_11202,N_11410);
nand U13882 (N_13882,N_12206,N_11183);
nand U13883 (N_13883,N_10086,N_11402);
nor U13884 (N_13884,N_12399,N_11188);
or U13885 (N_13885,N_10924,N_11737);
or U13886 (N_13886,N_12478,N_12431);
xor U13887 (N_13887,N_10671,N_11024);
or U13888 (N_13888,N_10784,N_10269);
and U13889 (N_13889,N_10479,N_11980);
xnor U13890 (N_13890,N_10773,N_11683);
or U13891 (N_13891,N_11602,N_11925);
nor U13892 (N_13892,N_10736,N_12238);
nand U13893 (N_13893,N_10315,N_11064);
xnor U13894 (N_13894,N_11122,N_11247);
xnor U13895 (N_13895,N_12277,N_11033);
or U13896 (N_13896,N_10051,N_10547);
or U13897 (N_13897,N_12163,N_11610);
or U13898 (N_13898,N_11066,N_10487);
nand U13899 (N_13899,N_11582,N_11620);
and U13900 (N_13900,N_10824,N_11508);
or U13901 (N_13901,N_10805,N_11231);
xnor U13902 (N_13902,N_11752,N_11075);
nand U13903 (N_13903,N_10373,N_11438);
nor U13904 (N_13904,N_11803,N_11954);
and U13905 (N_13905,N_11345,N_11480);
or U13906 (N_13906,N_12250,N_10607);
nor U13907 (N_13907,N_10211,N_10086);
nor U13908 (N_13908,N_10902,N_10989);
or U13909 (N_13909,N_12201,N_10297);
nor U13910 (N_13910,N_10593,N_10580);
or U13911 (N_13911,N_12105,N_11105);
xor U13912 (N_13912,N_11611,N_10874);
and U13913 (N_13913,N_11036,N_10595);
xor U13914 (N_13914,N_10794,N_11640);
or U13915 (N_13915,N_12097,N_11170);
and U13916 (N_13916,N_10829,N_10950);
or U13917 (N_13917,N_11088,N_10377);
or U13918 (N_13918,N_10801,N_11630);
or U13919 (N_13919,N_10424,N_11947);
or U13920 (N_13920,N_10352,N_10621);
or U13921 (N_13921,N_10456,N_10065);
nor U13922 (N_13922,N_12068,N_12008);
nand U13923 (N_13923,N_11127,N_11456);
nand U13924 (N_13924,N_10864,N_12332);
and U13925 (N_13925,N_10172,N_10238);
nor U13926 (N_13926,N_11904,N_11548);
nand U13927 (N_13927,N_10993,N_12064);
nor U13928 (N_13928,N_11352,N_10844);
nor U13929 (N_13929,N_12475,N_11735);
xor U13930 (N_13930,N_12132,N_10567);
nand U13931 (N_13931,N_11735,N_12232);
and U13932 (N_13932,N_12470,N_11217);
nor U13933 (N_13933,N_12290,N_11131);
and U13934 (N_13934,N_10597,N_10326);
or U13935 (N_13935,N_10389,N_12113);
nand U13936 (N_13936,N_10822,N_11865);
nand U13937 (N_13937,N_10306,N_11954);
xnor U13938 (N_13938,N_11508,N_12055);
nor U13939 (N_13939,N_10800,N_10064);
and U13940 (N_13940,N_10761,N_10418);
and U13941 (N_13941,N_10924,N_10608);
xor U13942 (N_13942,N_10745,N_10954);
and U13943 (N_13943,N_12041,N_11399);
or U13944 (N_13944,N_11652,N_11412);
and U13945 (N_13945,N_11297,N_11160);
nand U13946 (N_13946,N_11442,N_12462);
and U13947 (N_13947,N_11209,N_11372);
nand U13948 (N_13948,N_10499,N_12177);
nand U13949 (N_13949,N_10616,N_10129);
and U13950 (N_13950,N_12039,N_10175);
or U13951 (N_13951,N_11040,N_10049);
nor U13952 (N_13952,N_11412,N_11363);
or U13953 (N_13953,N_10152,N_10337);
xor U13954 (N_13954,N_11401,N_12297);
xnor U13955 (N_13955,N_10564,N_10842);
nor U13956 (N_13956,N_11396,N_11671);
or U13957 (N_13957,N_11444,N_10123);
xor U13958 (N_13958,N_12169,N_12167);
and U13959 (N_13959,N_11486,N_10470);
and U13960 (N_13960,N_10964,N_11946);
or U13961 (N_13961,N_12280,N_12284);
nor U13962 (N_13962,N_10397,N_11413);
or U13963 (N_13963,N_11699,N_10095);
or U13964 (N_13964,N_11293,N_11590);
or U13965 (N_13965,N_11035,N_11015);
nor U13966 (N_13966,N_11952,N_11332);
nor U13967 (N_13967,N_10844,N_10527);
nand U13968 (N_13968,N_11208,N_11144);
and U13969 (N_13969,N_11450,N_11350);
xor U13970 (N_13970,N_11949,N_11115);
and U13971 (N_13971,N_10943,N_12489);
and U13972 (N_13972,N_10110,N_10235);
nor U13973 (N_13973,N_12368,N_11102);
nor U13974 (N_13974,N_12134,N_10514);
nand U13975 (N_13975,N_10938,N_11039);
and U13976 (N_13976,N_11608,N_12156);
nor U13977 (N_13977,N_10531,N_10343);
xnor U13978 (N_13978,N_12098,N_10834);
nor U13979 (N_13979,N_11140,N_12420);
or U13980 (N_13980,N_11317,N_11237);
xor U13981 (N_13981,N_10653,N_11313);
and U13982 (N_13982,N_10835,N_11052);
xor U13983 (N_13983,N_10654,N_12489);
nor U13984 (N_13984,N_10127,N_11695);
and U13985 (N_13985,N_11273,N_11828);
nand U13986 (N_13986,N_11714,N_12052);
or U13987 (N_13987,N_10162,N_10533);
or U13988 (N_13988,N_10063,N_12127);
xnor U13989 (N_13989,N_11654,N_10461);
nand U13990 (N_13990,N_11448,N_11850);
nand U13991 (N_13991,N_10071,N_10596);
and U13992 (N_13992,N_11561,N_10271);
nand U13993 (N_13993,N_10336,N_10638);
or U13994 (N_13994,N_11951,N_10852);
nand U13995 (N_13995,N_10238,N_11673);
xor U13996 (N_13996,N_10155,N_10458);
or U13997 (N_13997,N_10635,N_11430);
or U13998 (N_13998,N_11802,N_10623);
xnor U13999 (N_13999,N_12180,N_11097);
or U14000 (N_14000,N_11738,N_11794);
and U14001 (N_14001,N_11777,N_11587);
or U14002 (N_14002,N_10171,N_11697);
nand U14003 (N_14003,N_11417,N_11166);
nor U14004 (N_14004,N_12373,N_11195);
or U14005 (N_14005,N_11839,N_11118);
and U14006 (N_14006,N_12363,N_10876);
or U14007 (N_14007,N_12166,N_11163);
nor U14008 (N_14008,N_12356,N_10593);
and U14009 (N_14009,N_10934,N_12126);
and U14010 (N_14010,N_10653,N_10930);
nor U14011 (N_14011,N_12263,N_11975);
or U14012 (N_14012,N_11179,N_12091);
nor U14013 (N_14013,N_12257,N_11912);
and U14014 (N_14014,N_11172,N_10183);
or U14015 (N_14015,N_11238,N_10990);
nand U14016 (N_14016,N_12200,N_11200);
and U14017 (N_14017,N_11214,N_12443);
and U14018 (N_14018,N_12359,N_11811);
or U14019 (N_14019,N_11594,N_10034);
nand U14020 (N_14020,N_10939,N_11628);
and U14021 (N_14021,N_12211,N_10774);
or U14022 (N_14022,N_12031,N_10488);
xor U14023 (N_14023,N_11615,N_12299);
nand U14024 (N_14024,N_10651,N_11130);
or U14025 (N_14025,N_10336,N_10912);
nor U14026 (N_14026,N_10687,N_11669);
xnor U14027 (N_14027,N_11293,N_12198);
and U14028 (N_14028,N_11758,N_10754);
xnor U14029 (N_14029,N_10170,N_12141);
or U14030 (N_14030,N_10236,N_12425);
and U14031 (N_14031,N_10195,N_12092);
and U14032 (N_14032,N_10068,N_12361);
nand U14033 (N_14033,N_12257,N_11333);
or U14034 (N_14034,N_12353,N_10354);
and U14035 (N_14035,N_12428,N_11984);
nor U14036 (N_14036,N_10536,N_10668);
nand U14037 (N_14037,N_12273,N_10439);
or U14038 (N_14038,N_10785,N_11120);
or U14039 (N_14039,N_10453,N_11392);
xnor U14040 (N_14040,N_11161,N_10358);
xor U14041 (N_14041,N_12298,N_11895);
nand U14042 (N_14042,N_12074,N_11001);
and U14043 (N_14043,N_10398,N_10407);
xor U14044 (N_14044,N_10033,N_11559);
nor U14045 (N_14045,N_11073,N_11421);
and U14046 (N_14046,N_11362,N_11696);
or U14047 (N_14047,N_11341,N_10945);
nand U14048 (N_14048,N_11080,N_12119);
nor U14049 (N_14049,N_11074,N_10189);
and U14050 (N_14050,N_10319,N_11204);
and U14051 (N_14051,N_10624,N_11576);
and U14052 (N_14052,N_10770,N_11780);
and U14053 (N_14053,N_11949,N_10092);
nor U14054 (N_14054,N_10539,N_11746);
xor U14055 (N_14055,N_11168,N_11023);
nand U14056 (N_14056,N_11599,N_11528);
nand U14057 (N_14057,N_12006,N_10479);
nor U14058 (N_14058,N_11018,N_11407);
or U14059 (N_14059,N_10371,N_12444);
and U14060 (N_14060,N_12076,N_10035);
xor U14061 (N_14061,N_11085,N_12303);
nand U14062 (N_14062,N_12430,N_12254);
and U14063 (N_14063,N_10543,N_11713);
xnor U14064 (N_14064,N_11898,N_12042);
nor U14065 (N_14065,N_11049,N_10199);
nand U14066 (N_14066,N_11266,N_10853);
or U14067 (N_14067,N_11107,N_11401);
and U14068 (N_14068,N_11194,N_12380);
or U14069 (N_14069,N_12083,N_12169);
nand U14070 (N_14070,N_10182,N_11283);
or U14071 (N_14071,N_10585,N_11350);
and U14072 (N_14072,N_10270,N_10741);
or U14073 (N_14073,N_11078,N_11946);
and U14074 (N_14074,N_11794,N_11374);
xor U14075 (N_14075,N_11580,N_11337);
xor U14076 (N_14076,N_11823,N_10616);
nand U14077 (N_14077,N_11929,N_10222);
or U14078 (N_14078,N_12146,N_12224);
xnor U14079 (N_14079,N_11933,N_11812);
and U14080 (N_14080,N_10521,N_11256);
nor U14081 (N_14081,N_11887,N_12259);
xor U14082 (N_14082,N_10025,N_12414);
or U14083 (N_14083,N_10466,N_12380);
and U14084 (N_14084,N_10648,N_10357);
nor U14085 (N_14085,N_11957,N_10041);
and U14086 (N_14086,N_11321,N_10096);
and U14087 (N_14087,N_10236,N_12423);
nand U14088 (N_14088,N_11920,N_11985);
nor U14089 (N_14089,N_12296,N_11381);
nand U14090 (N_14090,N_12155,N_11939);
or U14091 (N_14091,N_11786,N_10459);
nand U14092 (N_14092,N_10985,N_12067);
nor U14093 (N_14093,N_12446,N_10974);
and U14094 (N_14094,N_10578,N_11318);
nand U14095 (N_14095,N_11668,N_11005);
nor U14096 (N_14096,N_11632,N_10957);
nand U14097 (N_14097,N_10764,N_10268);
or U14098 (N_14098,N_11545,N_10199);
nor U14099 (N_14099,N_12070,N_12450);
nor U14100 (N_14100,N_11099,N_11464);
nand U14101 (N_14101,N_10636,N_10072);
xor U14102 (N_14102,N_11628,N_10051);
xnor U14103 (N_14103,N_11065,N_11352);
or U14104 (N_14104,N_12263,N_10200);
or U14105 (N_14105,N_11045,N_12364);
nand U14106 (N_14106,N_10357,N_11846);
nor U14107 (N_14107,N_11840,N_11625);
nor U14108 (N_14108,N_10700,N_10610);
nor U14109 (N_14109,N_12308,N_12341);
nand U14110 (N_14110,N_10719,N_10338);
nor U14111 (N_14111,N_11012,N_12171);
xor U14112 (N_14112,N_10092,N_12136);
and U14113 (N_14113,N_11124,N_10198);
and U14114 (N_14114,N_11047,N_11388);
and U14115 (N_14115,N_11663,N_10650);
nand U14116 (N_14116,N_11819,N_11690);
and U14117 (N_14117,N_11938,N_11547);
xnor U14118 (N_14118,N_10937,N_11763);
nor U14119 (N_14119,N_11088,N_10164);
and U14120 (N_14120,N_12410,N_10303);
xnor U14121 (N_14121,N_10899,N_11874);
nand U14122 (N_14122,N_10122,N_11959);
xnor U14123 (N_14123,N_11871,N_10571);
or U14124 (N_14124,N_11528,N_10406);
nand U14125 (N_14125,N_11833,N_11109);
nand U14126 (N_14126,N_12470,N_11154);
and U14127 (N_14127,N_12141,N_12319);
and U14128 (N_14128,N_11095,N_11958);
nand U14129 (N_14129,N_11032,N_11524);
and U14130 (N_14130,N_10125,N_11851);
nand U14131 (N_14131,N_11121,N_12078);
or U14132 (N_14132,N_11812,N_11486);
xor U14133 (N_14133,N_10150,N_11958);
or U14134 (N_14134,N_11117,N_12086);
or U14135 (N_14135,N_11877,N_10358);
nand U14136 (N_14136,N_10170,N_11672);
xnor U14137 (N_14137,N_12078,N_11180);
and U14138 (N_14138,N_10641,N_10625);
and U14139 (N_14139,N_10710,N_12002);
and U14140 (N_14140,N_10458,N_10225);
nand U14141 (N_14141,N_10909,N_10976);
or U14142 (N_14142,N_11313,N_12132);
nand U14143 (N_14143,N_12434,N_12042);
nand U14144 (N_14144,N_10664,N_11055);
nor U14145 (N_14145,N_11662,N_11725);
nand U14146 (N_14146,N_10086,N_10162);
nor U14147 (N_14147,N_11023,N_11312);
xnor U14148 (N_14148,N_12066,N_11277);
nor U14149 (N_14149,N_11407,N_12233);
xor U14150 (N_14150,N_10896,N_12397);
nor U14151 (N_14151,N_10719,N_11816);
or U14152 (N_14152,N_11327,N_12381);
nor U14153 (N_14153,N_12149,N_11007);
nand U14154 (N_14154,N_10944,N_10642);
xnor U14155 (N_14155,N_10284,N_11690);
nand U14156 (N_14156,N_10622,N_12333);
nor U14157 (N_14157,N_11115,N_12273);
xnor U14158 (N_14158,N_11327,N_10148);
or U14159 (N_14159,N_11462,N_10853);
or U14160 (N_14160,N_10530,N_12447);
nand U14161 (N_14161,N_10519,N_10398);
and U14162 (N_14162,N_12436,N_10945);
xnor U14163 (N_14163,N_10212,N_11769);
or U14164 (N_14164,N_10129,N_10749);
xor U14165 (N_14165,N_12467,N_10351);
xnor U14166 (N_14166,N_10926,N_12067);
nor U14167 (N_14167,N_10593,N_12498);
and U14168 (N_14168,N_11606,N_12267);
xnor U14169 (N_14169,N_11563,N_12117);
nand U14170 (N_14170,N_12419,N_11930);
xor U14171 (N_14171,N_10506,N_10285);
nand U14172 (N_14172,N_10170,N_11935);
nor U14173 (N_14173,N_10254,N_10122);
and U14174 (N_14174,N_10033,N_10630);
nor U14175 (N_14175,N_11253,N_11753);
and U14176 (N_14176,N_10836,N_10421);
nand U14177 (N_14177,N_12368,N_10810);
nor U14178 (N_14178,N_11334,N_12459);
xnor U14179 (N_14179,N_11003,N_10298);
nand U14180 (N_14180,N_11076,N_12154);
or U14181 (N_14181,N_11480,N_10260);
nand U14182 (N_14182,N_10448,N_12361);
nor U14183 (N_14183,N_11576,N_10564);
xor U14184 (N_14184,N_12230,N_12085);
and U14185 (N_14185,N_11271,N_11907);
nand U14186 (N_14186,N_11853,N_12151);
nand U14187 (N_14187,N_11022,N_10445);
nand U14188 (N_14188,N_12110,N_10530);
or U14189 (N_14189,N_12240,N_10310);
xnor U14190 (N_14190,N_10373,N_11342);
nor U14191 (N_14191,N_11234,N_11570);
xnor U14192 (N_14192,N_10014,N_10675);
nor U14193 (N_14193,N_10370,N_10588);
or U14194 (N_14194,N_10640,N_10824);
or U14195 (N_14195,N_10165,N_11232);
xor U14196 (N_14196,N_11775,N_10386);
or U14197 (N_14197,N_11843,N_10123);
or U14198 (N_14198,N_10001,N_10366);
and U14199 (N_14199,N_11834,N_11012);
or U14200 (N_14200,N_10231,N_11650);
or U14201 (N_14201,N_11876,N_11377);
and U14202 (N_14202,N_11435,N_11841);
nor U14203 (N_14203,N_10200,N_12355);
and U14204 (N_14204,N_12279,N_12034);
nand U14205 (N_14205,N_10487,N_10239);
nor U14206 (N_14206,N_10264,N_10568);
or U14207 (N_14207,N_10373,N_11633);
nand U14208 (N_14208,N_10922,N_10750);
nor U14209 (N_14209,N_11590,N_10268);
xnor U14210 (N_14210,N_10411,N_11906);
nand U14211 (N_14211,N_11203,N_12135);
nand U14212 (N_14212,N_12075,N_12241);
nor U14213 (N_14213,N_10836,N_10088);
nor U14214 (N_14214,N_12014,N_11719);
and U14215 (N_14215,N_12165,N_11009);
or U14216 (N_14216,N_10436,N_10372);
xnor U14217 (N_14217,N_11754,N_11189);
or U14218 (N_14218,N_11788,N_12231);
xnor U14219 (N_14219,N_11482,N_10817);
or U14220 (N_14220,N_10529,N_10047);
or U14221 (N_14221,N_10942,N_11115);
or U14222 (N_14222,N_11149,N_10824);
xor U14223 (N_14223,N_10712,N_12493);
nor U14224 (N_14224,N_11473,N_12346);
xor U14225 (N_14225,N_11054,N_10810);
nor U14226 (N_14226,N_12317,N_12491);
and U14227 (N_14227,N_12037,N_11242);
nor U14228 (N_14228,N_12370,N_11487);
or U14229 (N_14229,N_10652,N_11734);
nor U14230 (N_14230,N_12299,N_11741);
nor U14231 (N_14231,N_11093,N_12046);
nor U14232 (N_14232,N_11521,N_11845);
or U14233 (N_14233,N_10064,N_12256);
nand U14234 (N_14234,N_11580,N_10735);
nor U14235 (N_14235,N_11733,N_12127);
and U14236 (N_14236,N_10422,N_11977);
xor U14237 (N_14237,N_12161,N_12448);
and U14238 (N_14238,N_10927,N_10215);
nand U14239 (N_14239,N_10542,N_10129);
nand U14240 (N_14240,N_10958,N_11437);
and U14241 (N_14241,N_11173,N_11361);
and U14242 (N_14242,N_10168,N_10081);
nor U14243 (N_14243,N_11225,N_11217);
nor U14244 (N_14244,N_11237,N_11232);
xnor U14245 (N_14245,N_10890,N_11868);
or U14246 (N_14246,N_10800,N_12103);
xor U14247 (N_14247,N_11550,N_11847);
nor U14248 (N_14248,N_11734,N_11990);
or U14249 (N_14249,N_11540,N_11566);
and U14250 (N_14250,N_12043,N_11091);
xor U14251 (N_14251,N_12192,N_11994);
nor U14252 (N_14252,N_11324,N_11512);
or U14253 (N_14253,N_10541,N_11961);
xor U14254 (N_14254,N_11136,N_12342);
or U14255 (N_14255,N_10633,N_12098);
xor U14256 (N_14256,N_11077,N_12082);
nand U14257 (N_14257,N_11764,N_10040);
and U14258 (N_14258,N_12142,N_10475);
nand U14259 (N_14259,N_11553,N_11402);
or U14260 (N_14260,N_12455,N_12150);
xnor U14261 (N_14261,N_11693,N_12488);
xor U14262 (N_14262,N_11085,N_12463);
nor U14263 (N_14263,N_11304,N_10427);
nor U14264 (N_14264,N_11103,N_12366);
nand U14265 (N_14265,N_10101,N_11222);
nor U14266 (N_14266,N_10345,N_11014);
xnor U14267 (N_14267,N_10383,N_11016);
nand U14268 (N_14268,N_12031,N_10358);
nor U14269 (N_14269,N_11064,N_11019);
nor U14270 (N_14270,N_10999,N_12316);
nand U14271 (N_14271,N_11676,N_12268);
or U14272 (N_14272,N_11258,N_10535);
and U14273 (N_14273,N_11626,N_11758);
xor U14274 (N_14274,N_11914,N_10428);
and U14275 (N_14275,N_11552,N_11163);
xnor U14276 (N_14276,N_12037,N_10316);
or U14277 (N_14277,N_10882,N_11098);
and U14278 (N_14278,N_11092,N_10105);
nand U14279 (N_14279,N_10500,N_11841);
or U14280 (N_14280,N_12199,N_10456);
and U14281 (N_14281,N_10315,N_12462);
or U14282 (N_14282,N_12258,N_12367);
and U14283 (N_14283,N_10007,N_12114);
nor U14284 (N_14284,N_11465,N_11148);
and U14285 (N_14285,N_10921,N_12446);
and U14286 (N_14286,N_12470,N_11826);
xor U14287 (N_14287,N_10746,N_11535);
nand U14288 (N_14288,N_10016,N_11281);
xnor U14289 (N_14289,N_12010,N_11824);
and U14290 (N_14290,N_12225,N_10030);
nand U14291 (N_14291,N_12197,N_10049);
xnor U14292 (N_14292,N_11156,N_10971);
nand U14293 (N_14293,N_11713,N_10675);
nor U14294 (N_14294,N_12428,N_11017);
or U14295 (N_14295,N_10768,N_12442);
or U14296 (N_14296,N_10673,N_12312);
nor U14297 (N_14297,N_10956,N_11258);
and U14298 (N_14298,N_11662,N_12140);
xnor U14299 (N_14299,N_10453,N_11655);
xnor U14300 (N_14300,N_11088,N_10235);
and U14301 (N_14301,N_11621,N_10931);
nor U14302 (N_14302,N_10736,N_12350);
and U14303 (N_14303,N_10285,N_11352);
or U14304 (N_14304,N_10766,N_10658);
xor U14305 (N_14305,N_10497,N_11010);
xor U14306 (N_14306,N_10107,N_10424);
or U14307 (N_14307,N_10264,N_12000);
nand U14308 (N_14308,N_12391,N_11046);
or U14309 (N_14309,N_10562,N_10707);
and U14310 (N_14310,N_11019,N_10708);
nand U14311 (N_14311,N_11424,N_12009);
and U14312 (N_14312,N_12373,N_10081);
nand U14313 (N_14313,N_11253,N_11387);
nand U14314 (N_14314,N_10168,N_10945);
nor U14315 (N_14315,N_12425,N_11500);
nand U14316 (N_14316,N_11123,N_12080);
or U14317 (N_14317,N_11821,N_12461);
or U14318 (N_14318,N_11804,N_11619);
nor U14319 (N_14319,N_10980,N_10013);
or U14320 (N_14320,N_10699,N_12375);
xnor U14321 (N_14321,N_10003,N_10999);
nor U14322 (N_14322,N_10034,N_10355);
nor U14323 (N_14323,N_10779,N_10540);
xor U14324 (N_14324,N_10229,N_10297);
or U14325 (N_14325,N_12413,N_10849);
or U14326 (N_14326,N_11535,N_11678);
or U14327 (N_14327,N_12319,N_10043);
nor U14328 (N_14328,N_10921,N_10200);
or U14329 (N_14329,N_10622,N_11388);
xnor U14330 (N_14330,N_10648,N_11880);
nand U14331 (N_14331,N_10882,N_12319);
nor U14332 (N_14332,N_10335,N_10290);
nand U14333 (N_14333,N_10828,N_11588);
xor U14334 (N_14334,N_11412,N_10557);
xor U14335 (N_14335,N_12255,N_10705);
xnor U14336 (N_14336,N_11636,N_10786);
nand U14337 (N_14337,N_10836,N_11622);
or U14338 (N_14338,N_11809,N_10290);
and U14339 (N_14339,N_10644,N_11363);
and U14340 (N_14340,N_11539,N_11876);
and U14341 (N_14341,N_10606,N_12393);
or U14342 (N_14342,N_10761,N_10616);
and U14343 (N_14343,N_10908,N_12266);
and U14344 (N_14344,N_11319,N_12109);
nand U14345 (N_14345,N_10311,N_11163);
nor U14346 (N_14346,N_10210,N_11105);
or U14347 (N_14347,N_11694,N_10368);
and U14348 (N_14348,N_11354,N_10270);
nand U14349 (N_14349,N_10990,N_10794);
nor U14350 (N_14350,N_12259,N_11417);
nand U14351 (N_14351,N_11332,N_11045);
nor U14352 (N_14352,N_10694,N_12038);
xnor U14353 (N_14353,N_10956,N_11809);
nand U14354 (N_14354,N_10627,N_10377);
and U14355 (N_14355,N_10514,N_10257);
xor U14356 (N_14356,N_12324,N_11050);
xnor U14357 (N_14357,N_10700,N_12321);
or U14358 (N_14358,N_10023,N_10687);
nand U14359 (N_14359,N_10769,N_10313);
xnor U14360 (N_14360,N_11772,N_10039);
or U14361 (N_14361,N_11033,N_12227);
xor U14362 (N_14362,N_10952,N_10097);
and U14363 (N_14363,N_11151,N_10992);
nand U14364 (N_14364,N_12374,N_10206);
xor U14365 (N_14365,N_11658,N_10579);
nor U14366 (N_14366,N_10786,N_10710);
or U14367 (N_14367,N_11672,N_10374);
nor U14368 (N_14368,N_12194,N_12433);
nand U14369 (N_14369,N_10272,N_11508);
or U14370 (N_14370,N_11142,N_11494);
nor U14371 (N_14371,N_11051,N_11688);
xnor U14372 (N_14372,N_11220,N_10925);
or U14373 (N_14373,N_10043,N_10099);
and U14374 (N_14374,N_11815,N_11076);
or U14375 (N_14375,N_11488,N_10436);
or U14376 (N_14376,N_12182,N_12391);
nand U14377 (N_14377,N_11963,N_11800);
or U14378 (N_14378,N_10204,N_10462);
or U14379 (N_14379,N_11650,N_11115);
nand U14380 (N_14380,N_11310,N_10307);
and U14381 (N_14381,N_12098,N_11745);
nand U14382 (N_14382,N_11320,N_12083);
and U14383 (N_14383,N_12493,N_12475);
nand U14384 (N_14384,N_11083,N_10332);
nand U14385 (N_14385,N_11745,N_10882);
xnor U14386 (N_14386,N_11716,N_12002);
nand U14387 (N_14387,N_12372,N_10166);
or U14388 (N_14388,N_10381,N_11115);
nor U14389 (N_14389,N_12483,N_11288);
and U14390 (N_14390,N_10575,N_11531);
xor U14391 (N_14391,N_11932,N_10999);
nor U14392 (N_14392,N_10758,N_11228);
xnor U14393 (N_14393,N_11297,N_11608);
and U14394 (N_14394,N_12138,N_10085);
nor U14395 (N_14395,N_12000,N_11320);
xor U14396 (N_14396,N_11454,N_11705);
nor U14397 (N_14397,N_10143,N_11884);
and U14398 (N_14398,N_12012,N_11518);
nand U14399 (N_14399,N_10759,N_12213);
and U14400 (N_14400,N_11282,N_11760);
nor U14401 (N_14401,N_11423,N_10741);
and U14402 (N_14402,N_11777,N_10983);
xnor U14403 (N_14403,N_10366,N_10281);
or U14404 (N_14404,N_10237,N_10372);
xor U14405 (N_14405,N_10261,N_11940);
xor U14406 (N_14406,N_10768,N_10140);
or U14407 (N_14407,N_11928,N_10789);
nor U14408 (N_14408,N_11973,N_12440);
or U14409 (N_14409,N_12044,N_11954);
nor U14410 (N_14410,N_11488,N_12489);
or U14411 (N_14411,N_10266,N_10811);
and U14412 (N_14412,N_10530,N_11225);
and U14413 (N_14413,N_11392,N_12076);
or U14414 (N_14414,N_12494,N_11365);
nor U14415 (N_14415,N_11701,N_12078);
and U14416 (N_14416,N_12343,N_11657);
nand U14417 (N_14417,N_10777,N_10056);
and U14418 (N_14418,N_11227,N_10994);
or U14419 (N_14419,N_12402,N_10866);
and U14420 (N_14420,N_11664,N_10330);
nor U14421 (N_14421,N_11989,N_10400);
or U14422 (N_14422,N_10702,N_11676);
or U14423 (N_14423,N_11210,N_10624);
xor U14424 (N_14424,N_11993,N_12155);
and U14425 (N_14425,N_11637,N_11184);
nor U14426 (N_14426,N_12310,N_10853);
nor U14427 (N_14427,N_11100,N_11217);
or U14428 (N_14428,N_10336,N_11038);
or U14429 (N_14429,N_10283,N_11224);
nand U14430 (N_14430,N_12072,N_12027);
nand U14431 (N_14431,N_10797,N_11294);
or U14432 (N_14432,N_11624,N_10251);
xnor U14433 (N_14433,N_10748,N_10120);
xnor U14434 (N_14434,N_12387,N_10189);
or U14435 (N_14435,N_10528,N_10597);
nor U14436 (N_14436,N_12216,N_11258);
or U14437 (N_14437,N_11225,N_12292);
nand U14438 (N_14438,N_11937,N_10163);
and U14439 (N_14439,N_11204,N_10698);
or U14440 (N_14440,N_11610,N_11969);
nand U14441 (N_14441,N_10177,N_11390);
or U14442 (N_14442,N_12467,N_12328);
nand U14443 (N_14443,N_12249,N_11655);
or U14444 (N_14444,N_10434,N_10893);
and U14445 (N_14445,N_11094,N_10056);
nand U14446 (N_14446,N_11770,N_10490);
nand U14447 (N_14447,N_10711,N_10654);
nand U14448 (N_14448,N_12038,N_10743);
nand U14449 (N_14449,N_12126,N_11591);
and U14450 (N_14450,N_11809,N_11639);
nand U14451 (N_14451,N_10698,N_12025);
nand U14452 (N_14452,N_11967,N_12128);
and U14453 (N_14453,N_11300,N_10101);
nand U14454 (N_14454,N_11883,N_11054);
xor U14455 (N_14455,N_10679,N_12474);
nor U14456 (N_14456,N_11943,N_10141);
nand U14457 (N_14457,N_11917,N_11066);
and U14458 (N_14458,N_11852,N_11028);
nor U14459 (N_14459,N_10527,N_11670);
xor U14460 (N_14460,N_12055,N_11292);
xnor U14461 (N_14461,N_11670,N_11528);
and U14462 (N_14462,N_12489,N_10949);
or U14463 (N_14463,N_11475,N_12251);
nor U14464 (N_14464,N_11436,N_10024);
xor U14465 (N_14465,N_12038,N_11506);
and U14466 (N_14466,N_11574,N_10048);
xnor U14467 (N_14467,N_11159,N_10691);
and U14468 (N_14468,N_11272,N_10795);
nor U14469 (N_14469,N_10672,N_12289);
nand U14470 (N_14470,N_11937,N_10020);
xor U14471 (N_14471,N_10706,N_10644);
and U14472 (N_14472,N_11669,N_11984);
nand U14473 (N_14473,N_10096,N_11332);
nand U14474 (N_14474,N_10321,N_11960);
or U14475 (N_14475,N_11080,N_10059);
and U14476 (N_14476,N_11374,N_10690);
xnor U14477 (N_14477,N_11617,N_11064);
xor U14478 (N_14478,N_11944,N_12007);
xnor U14479 (N_14479,N_10845,N_11176);
and U14480 (N_14480,N_10442,N_10672);
and U14481 (N_14481,N_11698,N_11989);
xor U14482 (N_14482,N_11750,N_10026);
nor U14483 (N_14483,N_12341,N_10898);
xnor U14484 (N_14484,N_11981,N_11682);
nand U14485 (N_14485,N_10103,N_11925);
xnor U14486 (N_14486,N_11176,N_10818);
nand U14487 (N_14487,N_10637,N_10536);
nor U14488 (N_14488,N_11300,N_11200);
and U14489 (N_14489,N_11985,N_10507);
nand U14490 (N_14490,N_11770,N_11931);
and U14491 (N_14491,N_11313,N_10746);
xor U14492 (N_14492,N_10410,N_10060);
nand U14493 (N_14493,N_11001,N_12409);
nand U14494 (N_14494,N_10778,N_10006);
xnor U14495 (N_14495,N_11534,N_10609);
xnor U14496 (N_14496,N_10398,N_11978);
xor U14497 (N_14497,N_11864,N_12035);
and U14498 (N_14498,N_12492,N_10053);
or U14499 (N_14499,N_10082,N_10168);
xor U14500 (N_14500,N_11426,N_10608);
nand U14501 (N_14501,N_11661,N_10116);
or U14502 (N_14502,N_10903,N_12329);
nand U14503 (N_14503,N_10220,N_11089);
or U14504 (N_14504,N_11499,N_12488);
nor U14505 (N_14505,N_12482,N_11978);
xor U14506 (N_14506,N_10610,N_10878);
nor U14507 (N_14507,N_12014,N_11000);
nand U14508 (N_14508,N_10056,N_12207);
and U14509 (N_14509,N_10405,N_10764);
and U14510 (N_14510,N_11988,N_10384);
nor U14511 (N_14511,N_12301,N_11235);
nand U14512 (N_14512,N_11751,N_11443);
or U14513 (N_14513,N_10827,N_11885);
nand U14514 (N_14514,N_12492,N_11552);
nand U14515 (N_14515,N_11670,N_11674);
xnor U14516 (N_14516,N_12467,N_11272);
or U14517 (N_14517,N_10785,N_11512);
or U14518 (N_14518,N_10033,N_11683);
or U14519 (N_14519,N_10434,N_11152);
or U14520 (N_14520,N_11361,N_11972);
xor U14521 (N_14521,N_10156,N_11373);
nor U14522 (N_14522,N_12143,N_10600);
nand U14523 (N_14523,N_10457,N_12056);
xor U14524 (N_14524,N_11640,N_11443);
nor U14525 (N_14525,N_11516,N_10172);
nor U14526 (N_14526,N_11353,N_12405);
and U14527 (N_14527,N_11707,N_11717);
or U14528 (N_14528,N_10017,N_10851);
or U14529 (N_14529,N_11039,N_10310);
nand U14530 (N_14530,N_11180,N_10424);
and U14531 (N_14531,N_11099,N_10566);
and U14532 (N_14532,N_10070,N_11270);
nand U14533 (N_14533,N_10139,N_11902);
and U14534 (N_14534,N_11912,N_11396);
nand U14535 (N_14535,N_10973,N_10075);
nand U14536 (N_14536,N_10681,N_11704);
xor U14537 (N_14537,N_10120,N_11513);
xor U14538 (N_14538,N_10414,N_11608);
xnor U14539 (N_14539,N_11201,N_11395);
nand U14540 (N_14540,N_11972,N_10378);
and U14541 (N_14541,N_10871,N_10272);
xor U14542 (N_14542,N_10996,N_11617);
xnor U14543 (N_14543,N_10046,N_10135);
and U14544 (N_14544,N_11379,N_11629);
xor U14545 (N_14545,N_12131,N_10638);
nor U14546 (N_14546,N_10225,N_11663);
or U14547 (N_14547,N_10027,N_10965);
nand U14548 (N_14548,N_10373,N_11900);
and U14549 (N_14549,N_10651,N_11602);
nor U14550 (N_14550,N_12147,N_12356);
and U14551 (N_14551,N_10126,N_10330);
and U14552 (N_14552,N_12449,N_11061);
xor U14553 (N_14553,N_11418,N_11372);
xor U14554 (N_14554,N_10371,N_10280);
xor U14555 (N_14555,N_12083,N_11998);
nor U14556 (N_14556,N_10462,N_12157);
nor U14557 (N_14557,N_10587,N_10479);
and U14558 (N_14558,N_10326,N_11551);
nand U14559 (N_14559,N_12150,N_10353);
xnor U14560 (N_14560,N_11076,N_10801);
and U14561 (N_14561,N_10359,N_11884);
nand U14562 (N_14562,N_10347,N_12374);
and U14563 (N_14563,N_12041,N_11902);
nand U14564 (N_14564,N_11205,N_12434);
nand U14565 (N_14565,N_11755,N_11279);
xor U14566 (N_14566,N_10000,N_12406);
nand U14567 (N_14567,N_10614,N_11479);
and U14568 (N_14568,N_10579,N_10186);
nor U14569 (N_14569,N_11616,N_12019);
nor U14570 (N_14570,N_10536,N_10582);
or U14571 (N_14571,N_11973,N_12095);
and U14572 (N_14572,N_10156,N_11717);
nand U14573 (N_14573,N_10187,N_11229);
and U14574 (N_14574,N_11511,N_10950);
or U14575 (N_14575,N_11289,N_10041);
nor U14576 (N_14576,N_12394,N_10850);
nor U14577 (N_14577,N_12491,N_10936);
and U14578 (N_14578,N_10963,N_11406);
nor U14579 (N_14579,N_11391,N_11857);
and U14580 (N_14580,N_11719,N_10013);
nor U14581 (N_14581,N_12015,N_12271);
nand U14582 (N_14582,N_10838,N_10168);
and U14583 (N_14583,N_11418,N_12280);
and U14584 (N_14584,N_12421,N_10099);
and U14585 (N_14585,N_12312,N_11029);
nor U14586 (N_14586,N_10734,N_10435);
nor U14587 (N_14587,N_11490,N_11670);
and U14588 (N_14588,N_10112,N_11999);
nor U14589 (N_14589,N_12085,N_11874);
xor U14590 (N_14590,N_11898,N_12283);
or U14591 (N_14591,N_10254,N_10117);
or U14592 (N_14592,N_10883,N_11178);
or U14593 (N_14593,N_10885,N_10124);
nor U14594 (N_14594,N_12222,N_10448);
xor U14595 (N_14595,N_11095,N_10123);
nor U14596 (N_14596,N_11823,N_11569);
or U14597 (N_14597,N_10848,N_12114);
nand U14598 (N_14598,N_11673,N_11839);
and U14599 (N_14599,N_12001,N_10051);
nor U14600 (N_14600,N_10209,N_11321);
xnor U14601 (N_14601,N_10234,N_11314);
nand U14602 (N_14602,N_12042,N_10718);
nor U14603 (N_14603,N_11963,N_11582);
xnor U14604 (N_14604,N_11711,N_10149);
xnor U14605 (N_14605,N_10986,N_11087);
xor U14606 (N_14606,N_10155,N_12245);
and U14607 (N_14607,N_11816,N_12193);
or U14608 (N_14608,N_10123,N_11573);
or U14609 (N_14609,N_10811,N_11558);
or U14610 (N_14610,N_10167,N_11834);
and U14611 (N_14611,N_10588,N_11906);
xnor U14612 (N_14612,N_11995,N_11616);
nand U14613 (N_14613,N_12295,N_10272);
xnor U14614 (N_14614,N_11269,N_12372);
nand U14615 (N_14615,N_10569,N_10410);
xor U14616 (N_14616,N_10115,N_11822);
or U14617 (N_14617,N_10812,N_10850);
nor U14618 (N_14618,N_11290,N_12261);
and U14619 (N_14619,N_11490,N_11639);
xnor U14620 (N_14620,N_10548,N_10497);
and U14621 (N_14621,N_10878,N_10505);
or U14622 (N_14622,N_11887,N_12303);
or U14623 (N_14623,N_10389,N_10199);
xnor U14624 (N_14624,N_10126,N_12237);
and U14625 (N_14625,N_10237,N_11849);
and U14626 (N_14626,N_10264,N_11842);
nor U14627 (N_14627,N_10921,N_10301);
and U14628 (N_14628,N_12381,N_11887);
nand U14629 (N_14629,N_10983,N_10108);
xor U14630 (N_14630,N_10507,N_10754);
nand U14631 (N_14631,N_10585,N_12017);
nand U14632 (N_14632,N_10895,N_11295);
nand U14633 (N_14633,N_10197,N_10922);
nor U14634 (N_14634,N_12194,N_12493);
or U14635 (N_14635,N_10994,N_10852);
or U14636 (N_14636,N_10256,N_12174);
or U14637 (N_14637,N_10126,N_11594);
or U14638 (N_14638,N_11918,N_12414);
nor U14639 (N_14639,N_11474,N_10846);
or U14640 (N_14640,N_11213,N_10600);
nand U14641 (N_14641,N_10457,N_11401);
and U14642 (N_14642,N_10093,N_10396);
or U14643 (N_14643,N_11637,N_10913);
nor U14644 (N_14644,N_10947,N_11768);
nand U14645 (N_14645,N_10830,N_10845);
and U14646 (N_14646,N_12402,N_10851);
and U14647 (N_14647,N_12402,N_10114);
and U14648 (N_14648,N_10908,N_12127);
nand U14649 (N_14649,N_11643,N_10838);
xor U14650 (N_14650,N_12121,N_11791);
nor U14651 (N_14651,N_10560,N_12092);
xnor U14652 (N_14652,N_12201,N_11181);
nand U14653 (N_14653,N_10918,N_12363);
xor U14654 (N_14654,N_10847,N_10433);
nand U14655 (N_14655,N_11452,N_11830);
nand U14656 (N_14656,N_10512,N_10753);
nand U14657 (N_14657,N_12122,N_10212);
or U14658 (N_14658,N_10343,N_12122);
xnor U14659 (N_14659,N_11225,N_11621);
nand U14660 (N_14660,N_10946,N_12472);
nand U14661 (N_14661,N_10616,N_11988);
xor U14662 (N_14662,N_12495,N_10094);
or U14663 (N_14663,N_10988,N_10174);
nor U14664 (N_14664,N_10945,N_10225);
nor U14665 (N_14665,N_10497,N_11002);
nand U14666 (N_14666,N_10343,N_10988);
nor U14667 (N_14667,N_11711,N_11898);
and U14668 (N_14668,N_10181,N_12195);
or U14669 (N_14669,N_12054,N_11027);
xnor U14670 (N_14670,N_11155,N_10539);
and U14671 (N_14671,N_10605,N_10583);
and U14672 (N_14672,N_11835,N_11157);
xnor U14673 (N_14673,N_10986,N_10452);
nor U14674 (N_14674,N_11196,N_11003);
or U14675 (N_14675,N_12203,N_10587);
and U14676 (N_14676,N_11905,N_11902);
xnor U14677 (N_14677,N_11973,N_11478);
or U14678 (N_14678,N_11289,N_10185);
xor U14679 (N_14679,N_10742,N_12228);
nor U14680 (N_14680,N_12431,N_11728);
and U14681 (N_14681,N_11419,N_11739);
nor U14682 (N_14682,N_10245,N_10223);
nand U14683 (N_14683,N_10176,N_11044);
nand U14684 (N_14684,N_10434,N_12252);
nor U14685 (N_14685,N_11741,N_10050);
and U14686 (N_14686,N_11260,N_12457);
and U14687 (N_14687,N_11369,N_11365);
and U14688 (N_14688,N_11772,N_11859);
and U14689 (N_14689,N_11224,N_11323);
or U14690 (N_14690,N_11299,N_11116);
nand U14691 (N_14691,N_10467,N_12398);
nor U14692 (N_14692,N_12208,N_11320);
and U14693 (N_14693,N_12050,N_10663);
nor U14694 (N_14694,N_11354,N_10881);
or U14695 (N_14695,N_11155,N_10153);
and U14696 (N_14696,N_11207,N_10982);
and U14697 (N_14697,N_12472,N_10829);
nor U14698 (N_14698,N_12204,N_10105);
and U14699 (N_14699,N_12456,N_10294);
xor U14700 (N_14700,N_10017,N_11287);
and U14701 (N_14701,N_10746,N_10487);
xnor U14702 (N_14702,N_10265,N_10797);
xnor U14703 (N_14703,N_12023,N_12109);
xor U14704 (N_14704,N_10936,N_11015);
and U14705 (N_14705,N_11437,N_11866);
nor U14706 (N_14706,N_12160,N_10507);
xor U14707 (N_14707,N_10315,N_11129);
nor U14708 (N_14708,N_10760,N_12136);
and U14709 (N_14709,N_10712,N_10240);
and U14710 (N_14710,N_12469,N_11061);
xor U14711 (N_14711,N_11895,N_10496);
and U14712 (N_14712,N_10732,N_10000);
and U14713 (N_14713,N_11419,N_10768);
nand U14714 (N_14714,N_11864,N_11299);
xor U14715 (N_14715,N_12056,N_11200);
nand U14716 (N_14716,N_10553,N_10713);
or U14717 (N_14717,N_12365,N_11408);
xor U14718 (N_14718,N_10495,N_10820);
nand U14719 (N_14719,N_10060,N_10696);
nand U14720 (N_14720,N_12125,N_10036);
and U14721 (N_14721,N_11695,N_11497);
and U14722 (N_14722,N_12345,N_12408);
xor U14723 (N_14723,N_11260,N_11925);
or U14724 (N_14724,N_11942,N_10590);
or U14725 (N_14725,N_12104,N_10070);
or U14726 (N_14726,N_10024,N_11488);
xor U14727 (N_14727,N_11825,N_12078);
xor U14728 (N_14728,N_11537,N_10469);
nand U14729 (N_14729,N_10842,N_11630);
nand U14730 (N_14730,N_11970,N_11811);
xnor U14731 (N_14731,N_12308,N_12449);
or U14732 (N_14732,N_10965,N_11129);
nor U14733 (N_14733,N_11271,N_10252);
or U14734 (N_14734,N_11654,N_12419);
nand U14735 (N_14735,N_11616,N_10978);
xor U14736 (N_14736,N_10346,N_10288);
nor U14737 (N_14737,N_12169,N_10417);
and U14738 (N_14738,N_10854,N_10160);
and U14739 (N_14739,N_12187,N_12448);
xor U14740 (N_14740,N_10106,N_10338);
nor U14741 (N_14741,N_10757,N_11853);
or U14742 (N_14742,N_11765,N_12463);
and U14743 (N_14743,N_12348,N_10331);
and U14744 (N_14744,N_12081,N_10055);
nand U14745 (N_14745,N_11728,N_11186);
xnor U14746 (N_14746,N_10836,N_10665);
and U14747 (N_14747,N_10759,N_12337);
or U14748 (N_14748,N_10553,N_11427);
nand U14749 (N_14749,N_11494,N_10338);
nor U14750 (N_14750,N_11276,N_10661);
nor U14751 (N_14751,N_12158,N_11656);
nor U14752 (N_14752,N_10781,N_11864);
nor U14753 (N_14753,N_10411,N_10142);
or U14754 (N_14754,N_10209,N_11546);
and U14755 (N_14755,N_10296,N_11577);
xor U14756 (N_14756,N_11808,N_11443);
nor U14757 (N_14757,N_10772,N_10120);
and U14758 (N_14758,N_11060,N_10173);
nor U14759 (N_14759,N_11461,N_10240);
or U14760 (N_14760,N_10820,N_12287);
nand U14761 (N_14761,N_11224,N_11594);
or U14762 (N_14762,N_11711,N_12360);
and U14763 (N_14763,N_12462,N_10675);
nand U14764 (N_14764,N_12212,N_10824);
nand U14765 (N_14765,N_11825,N_12145);
and U14766 (N_14766,N_11554,N_11194);
nand U14767 (N_14767,N_10367,N_10557);
or U14768 (N_14768,N_11524,N_11128);
xnor U14769 (N_14769,N_12334,N_10574);
or U14770 (N_14770,N_11563,N_10164);
xnor U14771 (N_14771,N_12482,N_10785);
and U14772 (N_14772,N_10473,N_11113);
or U14773 (N_14773,N_10582,N_11735);
xnor U14774 (N_14774,N_11589,N_10720);
and U14775 (N_14775,N_10021,N_10958);
and U14776 (N_14776,N_11411,N_11271);
nand U14777 (N_14777,N_10540,N_10767);
or U14778 (N_14778,N_10678,N_10587);
or U14779 (N_14779,N_10815,N_10356);
nor U14780 (N_14780,N_12013,N_10259);
or U14781 (N_14781,N_11272,N_11608);
and U14782 (N_14782,N_11711,N_10647);
or U14783 (N_14783,N_11686,N_11687);
or U14784 (N_14784,N_10915,N_12309);
xor U14785 (N_14785,N_11776,N_10326);
and U14786 (N_14786,N_11146,N_11170);
and U14787 (N_14787,N_11210,N_12418);
nor U14788 (N_14788,N_10471,N_11886);
and U14789 (N_14789,N_11426,N_12149);
and U14790 (N_14790,N_10720,N_10830);
nor U14791 (N_14791,N_11188,N_10277);
and U14792 (N_14792,N_12051,N_10415);
and U14793 (N_14793,N_10238,N_12135);
and U14794 (N_14794,N_11783,N_10804);
and U14795 (N_14795,N_10735,N_12296);
or U14796 (N_14796,N_10274,N_12072);
nor U14797 (N_14797,N_12007,N_10261);
and U14798 (N_14798,N_11251,N_12284);
nand U14799 (N_14799,N_10422,N_10085);
and U14800 (N_14800,N_11473,N_12125);
and U14801 (N_14801,N_12204,N_10911);
or U14802 (N_14802,N_11299,N_11322);
nor U14803 (N_14803,N_11542,N_10154);
nand U14804 (N_14804,N_12209,N_11804);
xor U14805 (N_14805,N_11457,N_12462);
and U14806 (N_14806,N_11520,N_11277);
and U14807 (N_14807,N_10320,N_10799);
or U14808 (N_14808,N_11230,N_11086);
nor U14809 (N_14809,N_10131,N_10583);
nand U14810 (N_14810,N_11614,N_12142);
and U14811 (N_14811,N_10696,N_11581);
or U14812 (N_14812,N_12340,N_10553);
or U14813 (N_14813,N_11207,N_10351);
nand U14814 (N_14814,N_10845,N_12101);
xnor U14815 (N_14815,N_11438,N_10745);
and U14816 (N_14816,N_10735,N_12293);
or U14817 (N_14817,N_12241,N_10521);
xor U14818 (N_14818,N_10156,N_10520);
and U14819 (N_14819,N_12345,N_11156);
nor U14820 (N_14820,N_11949,N_10793);
xor U14821 (N_14821,N_10413,N_11696);
or U14822 (N_14822,N_12360,N_10448);
nor U14823 (N_14823,N_10357,N_12349);
and U14824 (N_14824,N_12193,N_10841);
and U14825 (N_14825,N_11020,N_12237);
xnor U14826 (N_14826,N_12072,N_12257);
or U14827 (N_14827,N_11242,N_12004);
or U14828 (N_14828,N_12092,N_10332);
nand U14829 (N_14829,N_12355,N_10471);
nor U14830 (N_14830,N_11445,N_11157);
xnor U14831 (N_14831,N_12464,N_10457);
and U14832 (N_14832,N_11229,N_11669);
nor U14833 (N_14833,N_12304,N_10304);
and U14834 (N_14834,N_10165,N_10055);
nor U14835 (N_14835,N_11616,N_10374);
xor U14836 (N_14836,N_12109,N_11600);
and U14837 (N_14837,N_11371,N_11492);
and U14838 (N_14838,N_12186,N_11546);
or U14839 (N_14839,N_11900,N_10605);
or U14840 (N_14840,N_11010,N_11846);
xnor U14841 (N_14841,N_11186,N_10139);
and U14842 (N_14842,N_11320,N_11583);
xor U14843 (N_14843,N_12160,N_10406);
or U14844 (N_14844,N_10072,N_11989);
nand U14845 (N_14845,N_10063,N_10292);
nor U14846 (N_14846,N_12458,N_10565);
nor U14847 (N_14847,N_11024,N_12305);
nand U14848 (N_14848,N_11660,N_11164);
and U14849 (N_14849,N_10089,N_11712);
nor U14850 (N_14850,N_11310,N_10044);
and U14851 (N_14851,N_12067,N_12404);
xnor U14852 (N_14852,N_10561,N_11179);
xor U14853 (N_14853,N_10549,N_11879);
nor U14854 (N_14854,N_11691,N_10263);
nand U14855 (N_14855,N_11084,N_12011);
nor U14856 (N_14856,N_11996,N_10907);
nor U14857 (N_14857,N_10323,N_10789);
nand U14858 (N_14858,N_11989,N_11975);
and U14859 (N_14859,N_10914,N_11698);
xnor U14860 (N_14860,N_11228,N_11511);
xor U14861 (N_14861,N_10801,N_10805);
xor U14862 (N_14862,N_11961,N_12064);
and U14863 (N_14863,N_11862,N_11144);
and U14864 (N_14864,N_11500,N_10988);
and U14865 (N_14865,N_10673,N_10093);
xnor U14866 (N_14866,N_10931,N_11728);
xnor U14867 (N_14867,N_11856,N_10525);
xnor U14868 (N_14868,N_10861,N_10901);
xor U14869 (N_14869,N_12279,N_11263);
nand U14870 (N_14870,N_12272,N_12124);
or U14871 (N_14871,N_11057,N_10243);
xor U14872 (N_14872,N_10492,N_11744);
or U14873 (N_14873,N_11800,N_12336);
nand U14874 (N_14874,N_11349,N_10255);
and U14875 (N_14875,N_11438,N_10915);
or U14876 (N_14876,N_12222,N_11470);
nor U14877 (N_14877,N_10532,N_11498);
nor U14878 (N_14878,N_10121,N_10507);
nand U14879 (N_14879,N_12305,N_10777);
nor U14880 (N_14880,N_12083,N_12018);
nand U14881 (N_14881,N_10736,N_10066);
and U14882 (N_14882,N_10646,N_11345);
nor U14883 (N_14883,N_12344,N_12322);
and U14884 (N_14884,N_10565,N_10029);
and U14885 (N_14885,N_10701,N_11967);
and U14886 (N_14886,N_10505,N_10921);
xnor U14887 (N_14887,N_10225,N_10098);
nor U14888 (N_14888,N_10985,N_10429);
or U14889 (N_14889,N_11840,N_10993);
or U14890 (N_14890,N_10017,N_12216);
or U14891 (N_14891,N_10453,N_11292);
or U14892 (N_14892,N_10154,N_11714);
xnor U14893 (N_14893,N_11206,N_11126);
and U14894 (N_14894,N_11900,N_11603);
xnor U14895 (N_14895,N_11472,N_11180);
nor U14896 (N_14896,N_11354,N_11056);
nor U14897 (N_14897,N_11892,N_11085);
or U14898 (N_14898,N_12236,N_10001);
or U14899 (N_14899,N_10298,N_12180);
or U14900 (N_14900,N_11893,N_12448);
nor U14901 (N_14901,N_10750,N_11888);
nor U14902 (N_14902,N_11210,N_10413);
nor U14903 (N_14903,N_10637,N_11493);
xnor U14904 (N_14904,N_12409,N_11704);
or U14905 (N_14905,N_11992,N_10651);
xor U14906 (N_14906,N_10268,N_10522);
or U14907 (N_14907,N_12470,N_12367);
xnor U14908 (N_14908,N_11790,N_12376);
and U14909 (N_14909,N_10876,N_11438);
nand U14910 (N_14910,N_12154,N_10536);
nor U14911 (N_14911,N_10533,N_11895);
nor U14912 (N_14912,N_11763,N_11734);
xor U14913 (N_14913,N_11289,N_10206);
nor U14914 (N_14914,N_12144,N_12053);
xor U14915 (N_14915,N_11411,N_11701);
nand U14916 (N_14916,N_12193,N_10006);
nor U14917 (N_14917,N_10221,N_11985);
and U14918 (N_14918,N_10738,N_10338);
or U14919 (N_14919,N_12160,N_10736);
or U14920 (N_14920,N_10764,N_11667);
nand U14921 (N_14921,N_12459,N_12073);
nand U14922 (N_14922,N_10738,N_11929);
nor U14923 (N_14923,N_12310,N_10850);
nor U14924 (N_14924,N_10465,N_11196);
or U14925 (N_14925,N_10879,N_11595);
xnor U14926 (N_14926,N_12109,N_11555);
nor U14927 (N_14927,N_12328,N_12461);
and U14928 (N_14928,N_11510,N_10996);
xnor U14929 (N_14929,N_12459,N_11482);
nand U14930 (N_14930,N_11307,N_10389);
and U14931 (N_14931,N_10205,N_11981);
and U14932 (N_14932,N_10731,N_12285);
nand U14933 (N_14933,N_10150,N_12056);
or U14934 (N_14934,N_10129,N_10250);
or U14935 (N_14935,N_10614,N_10757);
nand U14936 (N_14936,N_11665,N_11245);
or U14937 (N_14937,N_11636,N_11198);
nand U14938 (N_14938,N_10691,N_10761);
nand U14939 (N_14939,N_10676,N_12046);
or U14940 (N_14940,N_11585,N_10658);
or U14941 (N_14941,N_10618,N_11963);
nand U14942 (N_14942,N_10872,N_12412);
or U14943 (N_14943,N_11250,N_12173);
nand U14944 (N_14944,N_10687,N_10581);
xor U14945 (N_14945,N_12279,N_11294);
and U14946 (N_14946,N_11805,N_10228);
nand U14947 (N_14947,N_10557,N_12468);
nor U14948 (N_14948,N_10700,N_11762);
nand U14949 (N_14949,N_11299,N_12243);
nand U14950 (N_14950,N_12091,N_10123);
and U14951 (N_14951,N_11638,N_11427);
or U14952 (N_14952,N_12486,N_11037);
nor U14953 (N_14953,N_11762,N_11698);
nor U14954 (N_14954,N_11195,N_11143);
or U14955 (N_14955,N_10410,N_10093);
and U14956 (N_14956,N_11004,N_10966);
nand U14957 (N_14957,N_11626,N_10120);
and U14958 (N_14958,N_12155,N_10118);
nand U14959 (N_14959,N_12012,N_12169);
and U14960 (N_14960,N_10483,N_11105);
nor U14961 (N_14961,N_12412,N_11783);
and U14962 (N_14962,N_11546,N_11988);
nand U14963 (N_14963,N_11950,N_12076);
or U14964 (N_14964,N_10182,N_10622);
xnor U14965 (N_14965,N_10094,N_12408);
nand U14966 (N_14966,N_12203,N_12414);
nor U14967 (N_14967,N_10670,N_10712);
and U14968 (N_14968,N_10927,N_12363);
nand U14969 (N_14969,N_10948,N_10546);
or U14970 (N_14970,N_12348,N_11300);
or U14971 (N_14971,N_10597,N_10753);
and U14972 (N_14972,N_12120,N_10679);
nor U14973 (N_14973,N_12149,N_11052);
xor U14974 (N_14974,N_10075,N_10905);
nor U14975 (N_14975,N_11336,N_10383);
nand U14976 (N_14976,N_10884,N_11378);
nand U14977 (N_14977,N_11840,N_11100);
nand U14978 (N_14978,N_10944,N_12011);
or U14979 (N_14979,N_10223,N_10149);
or U14980 (N_14980,N_12475,N_12364);
or U14981 (N_14981,N_12104,N_10105);
and U14982 (N_14982,N_11919,N_10296);
nor U14983 (N_14983,N_12156,N_12245);
or U14984 (N_14984,N_11547,N_11084);
nand U14985 (N_14985,N_11449,N_10002);
and U14986 (N_14986,N_10737,N_10391);
or U14987 (N_14987,N_11067,N_10958);
and U14988 (N_14988,N_12144,N_12010);
and U14989 (N_14989,N_10982,N_10148);
and U14990 (N_14990,N_12104,N_10737);
and U14991 (N_14991,N_11893,N_11550);
and U14992 (N_14992,N_11721,N_12342);
or U14993 (N_14993,N_12491,N_10893);
xnor U14994 (N_14994,N_10048,N_10278);
nand U14995 (N_14995,N_10992,N_11658);
and U14996 (N_14996,N_11722,N_11226);
and U14997 (N_14997,N_10351,N_10734);
and U14998 (N_14998,N_11956,N_10611);
nor U14999 (N_14999,N_12161,N_11685);
xnor U15000 (N_15000,N_13021,N_12586);
xor U15001 (N_15001,N_12857,N_12853);
nor U15002 (N_15002,N_14900,N_14304);
nor U15003 (N_15003,N_13091,N_13040);
nand U15004 (N_15004,N_13259,N_13568);
nand U15005 (N_15005,N_12817,N_13075);
nand U15006 (N_15006,N_12641,N_14416);
nor U15007 (N_15007,N_13024,N_14614);
nor U15008 (N_15008,N_13474,N_13762);
nor U15009 (N_15009,N_14366,N_14895);
and U15010 (N_15010,N_12511,N_13839);
nand U15011 (N_15011,N_12854,N_13123);
and U15012 (N_15012,N_13368,N_13353);
or U15013 (N_15013,N_14111,N_13890);
nand U15014 (N_15014,N_14270,N_13529);
and U15015 (N_15015,N_12660,N_13711);
xnor U15016 (N_15016,N_14972,N_13946);
xnor U15017 (N_15017,N_12856,N_13071);
nand U15018 (N_15018,N_12985,N_13935);
or U15019 (N_15019,N_13563,N_13057);
nor U15020 (N_15020,N_14051,N_13692);
nor U15021 (N_15021,N_13210,N_12613);
or U15022 (N_15022,N_14915,N_14894);
nand U15023 (N_15023,N_13352,N_14163);
xnor U15024 (N_15024,N_12737,N_14365);
xnor U15025 (N_15025,N_12756,N_14743);
or U15026 (N_15026,N_14092,N_13241);
nor U15027 (N_15027,N_14642,N_14695);
nor U15028 (N_15028,N_12674,N_13208);
xnor U15029 (N_15029,N_13826,N_13332);
xor U15030 (N_15030,N_13077,N_14734);
nor U15031 (N_15031,N_12678,N_12934);
nand U15032 (N_15032,N_12848,N_14218);
nand U15033 (N_15033,N_13911,N_14951);
nand U15034 (N_15034,N_13429,N_13171);
and U15035 (N_15035,N_13666,N_13899);
and U15036 (N_15036,N_14841,N_14648);
xor U15037 (N_15037,N_14262,N_13672);
nand U15038 (N_15038,N_14344,N_12640);
nand U15039 (N_15039,N_14714,N_14637);
and U15040 (N_15040,N_13402,N_12813);
or U15041 (N_15041,N_13074,N_13199);
nand U15042 (N_15042,N_13416,N_12529);
nand U15043 (N_15043,N_13372,N_12734);
nor U15044 (N_15044,N_14122,N_14280);
xor U15045 (N_15045,N_13482,N_13141);
and U15046 (N_15046,N_13460,N_14861);
nor U15047 (N_15047,N_14465,N_13824);
or U15048 (N_15048,N_12928,N_13318);
or U15049 (N_15049,N_13113,N_12929);
and U15050 (N_15050,N_12900,N_14212);
and U15051 (N_15051,N_13876,N_13580);
nor U15052 (N_15052,N_14526,N_12587);
nor U15053 (N_15053,N_13884,N_12581);
nor U15054 (N_15054,N_13090,N_12534);
nor U15055 (N_15055,N_14959,N_13206);
xor U15056 (N_15056,N_13599,N_14474);
nor U15057 (N_15057,N_13971,N_14472);
xnor U15058 (N_15058,N_14460,N_14878);
nor U15059 (N_15059,N_12805,N_13847);
nor U15060 (N_15060,N_12606,N_14077);
and U15061 (N_15061,N_14965,N_13183);
nor U15062 (N_15062,N_14192,N_14947);
xor U15063 (N_15063,N_14118,N_13357);
and U15064 (N_15064,N_13817,N_12912);
nor U15065 (N_15065,N_14055,N_14574);
nor U15066 (N_15066,N_13850,N_12924);
nor U15067 (N_15067,N_14740,N_13565);
nor U15068 (N_15068,N_13926,N_12758);
nor U15069 (N_15069,N_13735,N_14473);
nand U15070 (N_15070,N_12607,N_13653);
xnor U15071 (N_15071,N_13302,N_14263);
or U15072 (N_15072,N_13697,N_12712);
and U15073 (N_15073,N_12576,N_13301);
and U15074 (N_15074,N_13542,N_14483);
nand U15075 (N_15075,N_14679,N_13182);
xnor U15076 (N_15076,N_12878,N_12903);
or U15077 (N_15077,N_14957,N_14249);
and U15078 (N_15078,N_14333,N_12776);
and U15079 (N_15079,N_14004,N_14626);
and U15080 (N_15080,N_12802,N_14613);
and U15081 (N_15081,N_13006,N_14384);
xnor U15082 (N_15082,N_13651,N_14834);
and U15083 (N_15083,N_12648,N_13225);
and U15084 (N_15084,N_14401,N_13828);
xnor U15085 (N_15085,N_13224,N_13039);
nor U15086 (N_15086,N_13745,N_12974);
xor U15087 (N_15087,N_14730,N_13415);
nand U15088 (N_15088,N_14064,N_14583);
xnor U15089 (N_15089,N_12514,N_14228);
and U15090 (N_15090,N_14949,N_12620);
nor U15091 (N_15091,N_13596,N_12738);
xor U15092 (N_15092,N_13195,N_12736);
nor U15093 (N_15093,N_14508,N_14499);
and U15094 (N_15094,N_14133,N_14315);
xnor U15095 (N_15095,N_14413,N_13325);
or U15096 (N_15096,N_14265,N_12575);
nor U15097 (N_15097,N_14721,N_12894);
and U15098 (N_15098,N_14071,N_13881);
and U15099 (N_15099,N_14143,N_14034);
nor U15100 (N_15100,N_12713,N_13139);
or U15101 (N_15101,N_14288,N_14966);
nor U15102 (N_15102,N_13275,N_13780);
and U15103 (N_15103,N_13009,N_13766);
nor U15104 (N_15104,N_12793,N_13300);
and U15105 (N_15105,N_12763,N_13079);
or U15106 (N_15106,N_14693,N_14551);
nor U15107 (N_15107,N_14036,N_14833);
xor U15108 (N_15108,N_13437,N_12692);
or U15109 (N_15109,N_12783,N_14053);
or U15110 (N_15110,N_13231,N_13988);
or U15111 (N_15111,N_14439,N_12968);
xnor U15112 (N_15112,N_12787,N_14813);
nor U15113 (N_15113,N_13457,N_13747);
xor U15114 (N_15114,N_14598,N_14516);
xnor U15115 (N_15115,N_14805,N_13701);
nand U15116 (N_15116,N_12739,N_14845);
or U15117 (N_15117,N_14941,N_13055);
xor U15118 (N_15118,N_13291,N_13716);
and U15119 (N_15119,N_13041,N_14742);
nor U15120 (N_15120,N_13158,N_13549);
and U15121 (N_15121,N_14561,N_14292);
xnor U15122 (N_15122,N_13084,N_13710);
nand U15123 (N_15123,N_14425,N_14119);
nor U15124 (N_15124,N_13990,N_12530);
nor U15125 (N_15125,N_13401,N_12862);
or U15126 (N_15126,N_14308,N_14183);
or U15127 (N_15127,N_13648,N_13669);
or U15128 (N_15128,N_13865,N_12623);
nor U15129 (N_15129,N_13829,N_14698);
and U15130 (N_15130,N_14625,N_13103);
nand U15131 (N_15131,N_13362,N_13782);
nand U15132 (N_15132,N_14647,N_14584);
and U15133 (N_15133,N_14736,N_13894);
nand U15134 (N_15134,N_14496,N_14847);
or U15135 (N_15135,N_13956,N_14312);
and U15136 (N_15136,N_14872,N_12922);
and U15137 (N_15137,N_12957,N_12765);
nor U15138 (N_15138,N_13518,N_12730);
nor U15139 (N_15139,N_14198,N_12936);
nand U15140 (N_15140,N_13223,N_12914);
xnor U15141 (N_15141,N_14411,N_14552);
nand U15142 (N_15142,N_14083,N_13625);
or U15143 (N_15143,N_14402,N_12784);
and U15144 (N_15144,N_14671,N_14398);
nand U15145 (N_15145,N_13133,N_12927);
nor U15146 (N_15146,N_14152,N_13134);
or U15147 (N_15147,N_14891,N_12653);
and U15148 (N_15148,N_12506,N_13752);
xor U15149 (N_15149,N_13661,N_13382);
xor U15150 (N_15150,N_14432,N_14633);
nand U15151 (N_15151,N_14569,N_13554);
nand U15152 (N_15152,N_14171,N_14624);
and U15153 (N_15153,N_13665,N_13121);
nand U15154 (N_15154,N_13366,N_13067);
and U15155 (N_15155,N_12554,N_13720);
nor U15156 (N_15156,N_14423,N_14141);
nor U15157 (N_15157,N_14830,N_14375);
nor U15158 (N_15158,N_14520,N_13179);
nor U15159 (N_15159,N_13010,N_12639);
nor U15160 (N_15160,N_13583,N_12879);
xnor U15161 (N_15161,N_13546,N_14147);
and U15162 (N_15162,N_14126,N_13045);
nor U15163 (N_15163,N_14391,N_14291);
nand U15164 (N_15164,N_12532,N_13938);
nand U15165 (N_15165,N_12883,N_14911);
nand U15166 (N_15166,N_13432,N_14854);
nand U15167 (N_15167,N_13900,N_13691);
xor U15168 (N_15168,N_14128,N_12896);
or U15169 (N_15169,N_13390,N_12901);
nor U15170 (N_15170,N_13703,N_12637);
and U15171 (N_15171,N_12790,N_13029);
xor U15172 (N_15172,N_12944,N_14724);
nor U15173 (N_15173,N_14204,N_14576);
nor U15174 (N_15174,N_13386,N_13512);
xnor U15175 (N_15175,N_13879,N_13683);
nor U15176 (N_15176,N_13977,N_12995);
nor U15177 (N_15177,N_12709,N_13414);
and U15178 (N_15178,N_14210,N_13144);
or U15179 (N_15179,N_13165,N_13778);
nor U15180 (N_15180,N_14880,N_14162);
and U15181 (N_15181,N_13324,N_14142);
and U15182 (N_15182,N_12518,N_12565);
nand U15183 (N_15183,N_13030,N_14705);
nor U15184 (N_15184,N_12832,N_14362);
or U15185 (N_15185,N_13874,N_12838);
nand U15186 (N_15186,N_12899,N_14889);
and U15187 (N_15187,N_13545,N_13910);
nand U15188 (N_15188,N_12797,N_13586);
nand U15189 (N_15189,N_13145,N_12815);
nand U15190 (N_15190,N_12583,N_13532);
and U15191 (N_15191,N_14357,N_14992);
or U15192 (N_15192,N_14011,N_13557);
xor U15193 (N_15193,N_12723,N_14239);
nor U15194 (N_15194,N_14961,N_14999);
or U15195 (N_15195,N_13376,N_14471);
xor U15196 (N_15196,N_12604,N_13724);
or U15197 (N_15197,N_13870,N_12542);
or U15198 (N_15198,N_14794,N_13060);
nand U15199 (N_15199,N_14101,N_14106);
xor U15200 (N_15200,N_13394,N_14898);
or U15201 (N_15201,N_13571,N_13983);
xnor U15202 (N_15202,N_14843,N_14136);
and U15203 (N_15203,N_13775,N_14420);
xnor U15204 (N_15204,N_12963,N_13348);
and U15205 (N_15205,N_13633,N_13269);
and U15206 (N_15206,N_13449,N_13825);
or U15207 (N_15207,N_14103,N_14490);
nor U15208 (N_15208,N_13528,N_13837);
nand U15209 (N_15209,N_14683,N_14342);
nor U15210 (N_15210,N_13685,N_12543);
and U15211 (N_15211,N_13163,N_13732);
or U15212 (N_15212,N_14793,N_14699);
xor U15213 (N_15213,N_14719,N_14568);
or U15214 (N_15214,N_13730,N_14546);
and U15215 (N_15215,N_13388,N_14597);
or U15216 (N_15216,N_12906,N_13008);
and U15217 (N_15217,N_12726,N_14912);
nand U15218 (N_15218,N_14829,N_12778);
nand U15219 (N_15219,N_14823,N_13805);
xnor U15220 (N_15220,N_12722,N_13963);
nor U15221 (N_15221,N_13205,N_12917);
xnor U15222 (N_15222,N_14761,N_14662);
nor U15223 (N_15223,N_14305,N_12522);
nor U15224 (N_15224,N_13230,N_12907);
and U15225 (N_15225,N_13581,N_14766);
nand U15226 (N_15226,N_14603,N_14984);
nor U15227 (N_15227,N_14974,N_13750);
or U15228 (N_15228,N_14573,N_14187);
and U15229 (N_15229,N_12842,N_12701);
and U15230 (N_15230,N_14217,N_14336);
nor U15231 (N_15231,N_12958,N_14500);
and U15232 (N_15232,N_13834,N_13883);
xnor U15233 (N_15233,N_13383,N_14430);
nor U15234 (N_15234,N_12803,N_13843);
xnor U15235 (N_15235,N_14368,N_13806);
nor U15236 (N_15236,N_13342,N_14802);
or U15237 (N_15237,N_14628,N_13792);
xnor U15238 (N_15238,N_13168,N_13438);
nand U15239 (N_15239,N_14453,N_14021);
or U15240 (N_15240,N_12754,N_12889);
or U15241 (N_15241,N_14075,N_14247);
and U15242 (N_15242,N_12557,N_12560);
xor U15243 (N_15243,N_13840,N_14787);
nand U15244 (N_15244,N_12809,N_12845);
nand U15245 (N_15245,N_12685,N_13475);
and U15246 (N_15246,N_14246,N_14224);
nor U15247 (N_15247,N_14673,N_14195);
and U15248 (N_15248,N_12810,N_12647);
and U15249 (N_15249,N_14986,N_13048);
nor U15250 (N_15250,N_13212,N_12750);
nand U15251 (N_15251,N_13795,N_13652);
nor U15252 (N_15252,N_13235,N_13251);
xor U15253 (N_15253,N_14243,N_12682);
or U15254 (N_15254,N_12992,N_14388);
and U15255 (N_15255,N_14219,N_12686);
xor U15256 (N_15256,N_14556,N_14924);
xnor U15257 (N_15257,N_13303,N_12512);
or U15258 (N_15258,N_13214,N_14820);
nand U15259 (N_15259,N_14358,N_12749);
nor U15260 (N_15260,N_14919,N_14539);
and U15261 (N_15261,N_12932,N_13909);
and U15262 (N_15262,N_14571,N_12996);
xor U15263 (N_15263,N_12638,N_14073);
nand U15264 (N_15264,N_13934,N_14089);
and U15265 (N_15265,N_13455,N_13481);
nand U15266 (N_15266,N_14170,N_14370);
nor U15267 (N_15267,N_14562,N_12962);
xnor U15268 (N_15268,N_14528,N_12930);
nor U15269 (N_15269,N_13587,N_14776);
nor U15270 (N_15270,N_13738,N_14596);
nor U15271 (N_15271,N_14522,N_13072);
xor U15272 (N_15272,N_14079,N_14138);
and U15273 (N_15273,N_13517,N_14922);
or U15274 (N_15274,N_14713,N_13062);
or U15275 (N_15275,N_14864,N_14789);
nor U15276 (N_15276,N_13051,N_12649);
xnor U15277 (N_15277,N_14723,N_12866);
nand U15278 (N_15278,N_14942,N_14524);
and U15279 (N_15279,N_14301,N_13255);
xor U15280 (N_15280,N_13679,N_12579);
nor U15281 (N_15281,N_13328,N_14014);
and U15282 (N_15282,N_14026,N_12524);
and U15283 (N_15283,N_12875,N_13410);
xor U15284 (N_15284,N_13688,N_12696);
or U15285 (N_15285,N_13391,N_14165);
nor U15286 (N_15286,N_13660,N_14888);
and U15287 (N_15287,N_12855,N_14298);
nand U15288 (N_15288,N_13564,N_14995);
nor U15289 (N_15289,N_13480,N_14355);
and U15290 (N_15290,N_13823,N_13112);
xnor U15291 (N_15291,N_13734,N_14221);
and U15292 (N_15292,N_14241,N_12547);
xor U15293 (N_15293,N_14454,N_14801);
nor U15294 (N_15294,N_13603,N_14550);
nor U15295 (N_15295,N_13418,N_12510);
xnor U15296 (N_15296,N_13190,N_14741);
and U15297 (N_15297,N_14871,N_13490);
and U15298 (N_15298,N_13634,N_13459);
or U15299 (N_15299,N_14293,N_13802);
nor U15300 (N_15300,N_14792,N_14746);
xnor U15301 (N_15301,N_13717,N_13960);
or U15302 (N_15302,N_14545,N_14067);
nand U15303 (N_15303,N_13516,N_14168);
nor U15304 (N_15304,N_12688,N_14720);
nand U15305 (N_15305,N_14709,N_13308);
and U15306 (N_15306,N_14360,N_14710);
nor U15307 (N_15307,N_13708,N_14314);
nor U15308 (N_15308,N_14166,N_13638);
xnor U15309 (N_15309,N_13358,N_14252);
or U15310 (N_15310,N_13036,N_13411);
and U15311 (N_15311,N_12973,N_14988);
nor U15312 (N_15312,N_14767,N_13769);
nand U15313 (N_15313,N_14824,N_12675);
and U15314 (N_15314,N_14727,N_14859);
or U15315 (N_15315,N_13536,N_14918);
xnor U15316 (N_15316,N_14969,N_14117);
nor U15317 (N_15317,N_12905,N_14604);
xor U15318 (N_15318,N_13948,N_14404);
and U15319 (N_15319,N_13495,N_13675);
xor U15320 (N_15320,N_14784,N_14846);
nor U15321 (N_15321,N_14797,N_13019);
or U15322 (N_15322,N_13381,N_14890);
xnor U15323 (N_15323,N_13064,N_14739);
or U15324 (N_15324,N_13450,N_14428);
nand U15325 (N_15325,N_12634,N_14444);
and U15326 (N_15326,N_14809,N_13867);
or U15327 (N_15327,N_13526,N_13790);
and U15328 (N_15328,N_14121,N_13155);
or U15329 (N_15329,N_13256,N_13065);
or U15330 (N_15330,N_12741,N_13849);
nand U15331 (N_15331,N_13632,N_14635);
and U15332 (N_15332,N_14674,N_14334);
nor U15333 (N_15333,N_14735,N_14097);
and U15334 (N_15334,N_12567,N_14094);
nand U15335 (N_15335,N_13310,N_14786);
xnor U15336 (N_15336,N_12652,N_14160);
and U15337 (N_15337,N_14385,N_12646);
or U15338 (N_15338,N_14790,N_14663);
nor U15339 (N_15339,N_14948,N_14692);
nand U15340 (N_15340,N_13556,N_13830);
or U15341 (N_15341,N_13872,N_14634);
xnor U15342 (N_15342,N_14237,N_14901);
and U15343 (N_15343,N_14356,N_14191);
nand U15344 (N_15344,N_13476,N_13346);
nor U15345 (N_15345,N_13351,N_12695);
nor U15346 (N_15346,N_13500,N_13271);
xnor U15347 (N_15347,N_13667,N_13326);
or U15348 (N_15348,N_13470,N_14885);
and U15349 (N_15349,N_14837,N_14655);
and U15350 (N_15350,N_13969,N_14715);
xor U15351 (N_15351,N_12588,N_12538);
or U15352 (N_15352,N_13317,N_14641);
nand U15353 (N_15353,N_13550,N_12733);
nand U15354 (N_15354,N_14675,N_13932);
and U15355 (N_15355,N_13644,N_14234);
nor U15356 (N_15356,N_13868,N_13781);
or U15357 (N_15357,N_13746,N_13279);
and U15358 (N_15358,N_14232,N_12782);
xnor U15359 (N_15359,N_14436,N_14282);
nand U15360 (N_15360,N_14478,N_14681);
nor U15361 (N_15361,N_13033,N_13469);
nand U15362 (N_15362,N_13365,N_14669);
nand U15363 (N_15363,N_13807,N_14575);
and U15364 (N_15364,N_12779,N_14441);
and U15365 (N_15365,N_13201,N_13777);
and U15366 (N_15366,N_14883,N_14586);
or U15367 (N_15367,N_13125,N_12556);
nand U15368 (N_15368,N_12720,N_12852);
or U15369 (N_15369,N_13726,N_14914);
or U15370 (N_15370,N_12667,N_14866);
nor U15371 (N_15371,N_14803,N_14652);
and U15372 (N_15372,N_14560,N_12847);
xnor U15373 (N_15373,N_14410,N_13811);
xnor U15374 (N_15374,N_13026,N_14137);
or U15375 (N_15375,N_13392,N_13579);
nand U15376 (N_15376,N_13215,N_13111);
nand U15377 (N_15377,N_13582,N_13178);
xnor U15378 (N_15378,N_13860,N_13164);
xnor U15379 (N_15379,N_12550,N_12707);
and U15380 (N_15380,N_13612,N_12622);
nand U15381 (N_15381,N_13642,N_13445);
or U15382 (N_15382,N_14701,N_13323);
nand U15383 (N_15383,N_14572,N_14194);
nor U15384 (N_15384,N_14733,N_14704);
nor U15385 (N_15385,N_12888,N_12627);
nor U15386 (N_15386,N_12743,N_14372);
xnor U15387 (N_15387,N_14124,N_12745);
and U15388 (N_15388,N_14456,N_14328);
and U15389 (N_15389,N_13135,N_13740);
or U15390 (N_15390,N_13227,N_12504);
or U15391 (N_15391,N_14618,N_13770);
nor U15392 (N_15392,N_13345,N_13032);
nor U15393 (N_15393,N_13374,N_13265);
or U15394 (N_15394,N_13187,N_13809);
and U15395 (N_15395,N_13037,N_14341);
and U15396 (N_15396,N_14003,N_12697);
xor U15397 (N_15397,N_13405,N_12535);
and U15398 (N_15398,N_14236,N_13439);
and U15399 (N_15399,N_13728,N_13754);
nand U15400 (N_15400,N_12614,N_12540);
xnor U15401 (N_15401,N_13142,N_14134);
nand U15402 (N_15402,N_13501,N_13011);
and U15403 (N_15403,N_12561,N_13204);
xnor U15404 (N_15404,N_12700,N_14527);
nor U15405 (N_15405,N_14485,N_14050);
and U15406 (N_15406,N_14035,N_13160);
and U15407 (N_15407,N_13785,N_13764);
or U15408 (N_15408,N_13589,N_13943);
nor U15409 (N_15409,N_14033,N_13192);
and U15410 (N_15410,N_13404,N_14159);
nor U15411 (N_15411,N_14184,N_12811);
nor U15412 (N_15412,N_13798,N_14340);
xor U15413 (N_15413,N_13330,N_14795);
and U15414 (N_15414,N_13000,N_12822);
or U15415 (N_15415,N_14838,N_12578);
nor U15416 (N_15416,N_14081,N_12689);
xor U15417 (N_15417,N_13656,N_14181);
nor U15418 (N_15418,N_14040,N_12501);
or U15419 (N_15419,N_14349,N_12771);
or U15420 (N_15420,N_13184,N_14352);
xor U15421 (N_15421,N_12960,N_13491);
or U15422 (N_15422,N_14361,N_14608);
or U15423 (N_15423,N_12869,N_14629);
and U15424 (N_15424,N_14131,N_14935);
and U15425 (N_15425,N_13737,N_14758);
xnor U15426 (N_15426,N_12618,N_14459);
and U15427 (N_15427,N_13087,N_14798);
and U15428 (N_15428,N_14072,N_14065);
or U15429 (N_15429,N_13624,N_13797);
xor U15430 (N_15430,N_14707,N_14728);
and U15431 (N_15431,N_13851,N_13757);
nor U15432 (N_15432,N_13061,N_13560);
nor U15433 (N_15433,N_12877,N_13788);
and U15434 (N_15434,N_12943,N_13170);
or U15435 (N_15435,N_14354,N_14172);
nand U15436 (N_15436,N_13869,N_13947);
nor U15437 (N_15437,N_13114,N_13425);
or U15438 (N_15438,N_14863,N_13494);
nand U15439 (N_15439,N_14238,N_13319);
nor U15440 (N_15440,N_14156,N_14418);
and U15441 (N_15441,N_13329,N_14009);
and U15442 (N_15442,N_13502,N_13393);
nor U15443 (N_15443,N_13497,N_14382);
and U15444 (N_15444,N_12595,N_14022);
nor U15445 (N_15445,N_14320,N_14585);
xnor U15446 (N_15446,N_14543,N_13083);
or U15447 (N_15447,N_13349,N_14250);
and U15448 (N_15448,N_14373,N_13217);
or U15449 (N_15449,N_14811,N_14182);
and U15450 (N_15450,N_14645,N_14825);
nand U15451 (N_15451,N_13743,N_14529);
or U15452 (N_15452,N_13298,N_14831);
or U15453 (N_15453,N_13982,N_14929);
nor U15454 (N_15454,N_13246,N_14203);
or U15455 (N_15455,N_12863,N_12572);
xor U15456 (N_15456,N_14690,N_14667);
nand U15457 (N_15457,N_14994,N_14495);
and U15458 (N_15458,N_13094,N_13548);
xor U15459 (N_15459,N_13191,N_12961);
nand U15460 (N_15460,N_13631,N_13668);
nand U15461 (N_15461,N_14466,N_12629);
nor U15462 (N_15462,N_13397,N_13422);
and U15463 (N_15463,N_14916,N_14819);
nand U15464 (N_15464,N_14330,N_12661);
or U15465 (N_15465,N_12824,N_13306);
nand U15466 (N_15466,N_12904,N_13361);
and U15467 (N_15467,N_14744,N_14627);
nand U15468 (N_15468,N_13428,N_14477);
and U15469 (N_15469,N_13095,N_13248);
xnor U15470 (N_15470,N_12564,N_14599);
nand U15471 (N_15471,N_13974,N_13477);
nor U15472 (N_15472,N_12525,N_13796);
xor U15473 (N_15473,N_13493,N_13994);
or U15474 (N_15474,N_12999,N_13233);
and U15475 (N_15475,N_14818,N_13772);
xor U15476 (N_15476,N_14945,N_14504);
or U15477 (N_15477,N_12761,N_13435);
or U15478 (N_15478,N_12570,N_12990);
xor U15479 (N_15479,N_14016,N_13143);
xnor U15480 (N_15480,N_14174,N_13132);
or U15481 (N_15481,N_12791,N_14415);
nand U15482 (N_15482,N_13857,N_12600);
nor U15483 (N_15483,N_14407,N_14879);
xnor U15484 (N_15484,N_14509,N_14567);
nor U15485 (N_15485,N_13373,N_13588);
or U15486 (N_15486,N_12502,N_13186);
xor U15487 (N_15487,N_14983,N_14093);
nor U15488 (N_15488,N_14844,N_12585);
nor U15489 (N_15489,N_14541,N_12757);
or U15490 (N_15490,N_14056,N_14000);
nand U15491 (N_15491,N_12704,N_14505);
and U15492 (N_15492,N_13846,N_13263);
and U15493 (N_15493,N_12965,N_14595);
or U15494 (N_15494,N_12898,N_13098);
or U15495 (N_15495,N_14881,N_14343);
xnor U15496 (N_15496,N_13050,N_14849);
or U15497 (N_15497,N_13022,N_14737);
or U15498 (N_15498,N_13028,N_14353);
nor U15499 (N_15499,N_14756,N_13447);
xor U15500 (N_15500,N_14445,N_14109);
or U15501 (N_15501,N_13942,N_13140);
nor U15502 (N_15502,N_13268,N_13174);
nand U15503 (N_15503,N_14007,N_12979);
xor U15504 (N_15504,N_14222,N_13069);
xnor U15505 (N_15505,N_14037,N_13654);
nor U15506 (N_15506,N_13852,N_14917);
xnor U15507 (N_15507,N_14462,N_14082);
nand U15508 (N_15508,N_12887,N_12939);
or U15509 (N_15509,N_13896,N_13842);
xnor U15510 (N_15510,N_14013,N_14799);
nand U15511 (N_15511,N_13610,N_14964);
xor U15512 (N_15512,N_13012,N_14113);
and U15513 (N_15513,N_13014,N_13479);
or U15514 (N_15514,N_12799,N_14893);
and U15515 (N_15515,N_14680,N_13451);
nor U15516 (N_15516,N_14621,N_14158);
or U15517 (N_15517,N_14302,N_13068);
and U15518 (N_15518,N_13955,N_14976);
xor U15519 (N_15519,N_13901,N_13923);
nand U15520 (N_15520,N_14610,N_13995);
nor U15521 (N_15521,N_12975,N_13194);
and U15522 (N_15522,N_14449,N_13446);
nand U15523 (N_15523,N_12735,N_13487);
and U15524 (N_15524,N_13765,N_13907);
or U15525 (N_15525,N_14279,N_14745);
xor U15526 (N_15526,N_12827,N_12507);
nand U15527 (N_15527,N_14877,N_14380);
nand U15528 (N_15528,N_13262,N_13761);
xor U15529 (N_15529,N_14763,N_14087);
and U15530 (N_15530,N_13294,N_13862);
xor U15531 (N_15531,N_12989,N_13698);
nand U15532 (N_15532,N_14294,N_12794);
xnor U15533 (N_15533,N_13334,N_14271);
nor U15534 (N_15534,N_12633,N_14409);
nand U15535 (N_15535,N_14010,N_13931);
or U15536 (N_15536,N_14587,N_13944);
and U15537 (N_15537,N_12873,N_13573);
xor U15538 (N_15538,N_14507,N_14902);
xnor U15539 (N_15539,N_12706,N_12621);
nand U15540 (N_15540,N_14731,N_14486);
or U15541 (N_15541,N_14835,N_14856);
nand U15542 (N_15542,N_14175,N_13906);
nand U15543 (N_15543,N_14677,N_13838);
or U15544 (N_15544,N_13277,N_13104);
or U15545 (N_15545,N_13154,N_13292);
and U15546 (N_15546,N_13025,N_14078);
or U15547 (N_15547,N_12603,N_14268);
nand U15548 (N_15548,N_14654,N_13222);
nand U15549 (N_15549,N_13590,N_13289);
xor U15550 (N_15550,N_13617,N_13034);
xnor U15551 (N_15551,N_14150,N_13288);
nand U15552 (N_15552,N_13722,N_13871);
nand U15553 (N_15553,N_12785,N_14909);
nand U15554 (N_15554,N_13063,N_13454);
xor U15555 (N_15555,N_13727,N_13917);
or U15556 (N_15556,N_12828,N_13370);
nor U15557 (N_15557,N_13767,N_12573);
xnor U15558 (N_15558,N_14908,N_13736);
and U15559 (N_15559,N_13835,N_12643);
xnor U15560 (N_15560,N_14685,N_14297);
nor U15561 (N_15561,N_13385,N_13998);
nor U15562 (N_15562,N_14286,N_14682);
or U15563 (N_15563,N_14855,N_12755);
or U15564 (N_15564,N_13086,N_13167);
nand U15565 (N_15565,N_13137,N_14242);
xnor U15566 (N_15566,N_14289,N_13774);
xor U15567 (N_15567,N_14201,N_13902);
xor U15568 (N_15568,N_13359,N_13677);
and U15569 (N_15569,N_12569,N_13013);
or U15570 (N_15570,N_12945,N_14632);
xnor U15571 (N_15571,N_13254,N_13209);
xnor U15572 (N_15572,N_14266,N_14132);
nor U15573 (N_15573,N_13478,N_14812);
and U15574 (N_15574,N_13066,N_13929);
or U15575 (N_15575,N_14594,N_13569);
xnor U15576 (N_15576,N_13885,N_14532);
or U15577 (N_15577,N_14392,N_13898);
xnor U15578 (N_15578,N_13522,N_14157);
and U15579 (N_15579,N_14503,N_13696);
and U15580 (N_15580,N_14639,N_14980);
and U15581 (N_15581,N_14419,N_14920);
nor U15582 (N_15582,N_14395,N_14070);
xor U15583 (N_15583,N_13379,N_13196);
xor U15584 (N_15584,N_13097,N_13047);
and U15585 (N_15585,N_14538,N_13059);
xor U15586 (N_15586,N_13702,N_14069);
and U15587 (N_15587,N_13641,N_14451);
and U15588 (N_15588,N_14827,N_14497);
nand U15589 (N_15589,N_14455,N_13198);
xnor U15590 (N_15590,N_14619,N_13007);
xor U15591 (N_15591,N_14311,N_13316);
xnor U15592 (N_15592,N_13693,N_13472);
or U15593 (N_15593,N_12568,N_14110);
nor U15594 (N_15594,N_14295,N_14853);
or U15595 (N_15595,N_13577,N_14190);
or U15596 (N_15596,N_14042,N_14753);
or U15597 (N_15597,N_13887,N_14140);
nand U15598 (N_15598,N_13753,N_12775);
nor U15599 (N_15599,N_13150,N_12931);
or U15600 (N_15600,N_13530,N_14778);
nand U15601 (N_15601,N_14227,N_14934);
and U15602 (N_15602,N_13367,N_13783);
or U15603 (N_15603,N_14440,N_14264);
and U15604 (N_15604,N_12994,N_14927);
nand U15605 (N_15605,N_14697,N_13813);
and U15606 (N_15606,N_12610,N_14781);
xor U15607 (N_15607,N_13681,N_14359);
nand U15608 (N_15608,N_14638,N_12670);
and U15609 (N_15609,N_13819,N_14005);
nor U15610 (N_15610,N_13848,N_12959);
and U15611 (N_15611,N_14332,N_14207);
and U15612 (N_15612,N_14257,N_13629);
or U15613 (N_15613,N_13489,N_14732);
nand U15614 (N_15614,N_13620,N_13339);
and U15615 (N_15615,N_14167,N_14696);
xor U15616 (N_15616,N_14002,N_13670);
or U15617 (N_15617,N_12672,N_14422);
xnor U15618 (N_15618,N_13311,N_14678);
nand U15619 (N_15619,N_13314,N_13207);
or U15620 (N_15620,N_12951,N_12976);
xor U15621 (N_15621,N_12562,N_13290);
and U15622 (N_15622,N_13682,N_13771);
nor U15623 (N_15623,N_13636,N_13122);
xor U15624 (N_15624,N_13115,N_13453);
or U15625 (N_15625,N_13733,N_14897);
xor U15626 (N_15626,N_14031,N_13739);
nor U15627 (N_15627,N_13966,N_13985);
and U15628 (N_15628,N_12897,N_12744);
nand U15629 (N_15629,N_13044,N_14606);
and U15630 (N_15630,N_13338,N_13552);
or U15631 (N_15631,N_14408,N_14046);
nand U15632 (N_15632,N_12582,N_14501);
nor U15633 (N_15633,N_12800,N_14565);
nand U15634 (N_15634,N_12978,N_14276);
and U15635 (N_15635,N_14684,N_12839);
nand U15636 (N_15636,N_14400,N_14102);
and U15637 (N_15637,N_13915,N_12972);
nor U15638 (N_15638,N_14600,N_13360);
and U15639 (N_15639,N_14179,N_12657);
nor U15640 (N_15640,N_12865,N_13551);
nor U15641 (N_15641,N_14383,N_13964);
or U15642 (N_15642,N_14043,N_13193);
or U15643 (N_15643,N_13570,N_13488);
nor U15644 (N_15644,N_12705,N_14750);
nand U15645 (N_15645,N_13157,N_14326);
or U15646 (N_15646,N_12804,N_14852);
xnor U15647 (N_15647,N_13464,N_14044);
or U15648 (N_15648,N_13341,N_14953);
nand U15649 (N_15649,N_14389,N_12611);
xnor U15650 (N_15650,N_14154,N_13002);
and U15651 (N_15651,N_13177,N_14839);
nor U15652 (N_15652,N_14985,N_14665);
nand U15653 (N_15653,N_13156,N_13120);
nand U15654 (N_15654,N_13356,N_12777);
xnor U15655 (N_15655,N_13020,N_12694);
and U15656 (N_15656,N_13704,N_12703);
nand U15657 (N_15657,N_14135,N_13803);
or U15658 (N_15658,N_13804,N_12806);
nand U15659 (N_15659,N_14273,N_12768);
and U15660 (N_15660,N_14582,N_14765);
xor U15661 (N_15661,N_12858,N_14782);
or U15662 (N_15662,N_12505,N_14689);
and U15663 (N_15663,N_12690,N_13908);
nor U15664 (N_15664,N_14115,N_14832);
nor U15665 (N_15665,N_14518,N_14609);
and U15666 (N_15666,N_14602,N_13169);
or U15667 (N_15667,N_14099,N_13864);
or U15668 (N_15668,N_13043,N_13371);
or U15669 (N_15669,N_13575,N_14622);
nand U15670 (N_15670,N_12955,N_12859);
xnor U15671 (N_15671,N_13604,N_14189);
xor U15672 (N_15672,N_13784,N_13786);
or U15673 (N_15673,N_12599,N_14202);
xor U15674 (N_15674,N_14272,N_14973);
nor U15675 (N_15675,N_13646,N_13327);
nand U15676 (N_15676,N_13893,N_14048);
and U15677 (N_15677,N_13389,N_14952);
xor U15678 (N_15678,N_13426,N_13678);
nand U15679 (N_15679,N_12624,N_14636);
nand U15680 (N_15680,N_12753,N_13615);
or U15681 (N_15681,N_14318,N_12503);
or U15682 (N_15682,N_12580,N_14519);
nor U15683 (N_15683,N_14484,N_14962);
or U15684 (N_15684,N_12981,N_13949);
and U15685 (N_15685,N_12593,N_12954);
nand U15686 (N_15686,N_12528,N_12772);
and U15687 (N_15687,N_13801,N_14275);
nor U15688 (N_15688,N_14762,N_12876);
and U15689 (N_15689,N_13891,N_12515);
nor U15690 (N_15690,N_13240,N_14876);
xnor U15691 (N_15691,N_13742,N_13886);
xor U15692 (N_15692,N_13607,N_14788);
or U15693 (N_15693,N_12868,N_14085);
nand U15694 (N_15694,N_13286,N_14722);
and U15695 (N_15695,N_13831,N_12792);
or U15696 (N_15696,N_12764,N_14084);
nand U15697 (N_15697,N_14105,N_12964);
nor U15698 (N_15698,N_14299,N_14796);
nor U15699 (N_15699,N_14397,N_13967);
and U15700 (N_15700,N_14656,N_14329);
nand U15701 (N_15701,N_13705,N_12710);
and U15702 (N_15702,N_13505,N_14027);
or U15703 (N_15703,N_14188,N_12601);
nor U15704 (N_15704,N_13856,N_13627);
xnor U15705 (N_15705,N_13082,N_14536);
nor U15706 (N_15706,N_14930,N_13015);
nor U15707 (N_15707,N_13544,N_13004);
and U15708 (N_15708,N_12748,N_13566);
or U15709 (N_15709,N_13562,N_13431);
xor U15710 (N_15710,N_14772,N_14339);
nor U15711 (N_15711,N_13380,N_13543);
nand U15712 (N_15712,N_14593,N_14590);
nor U15713 (N_15713,N_13689,N_14650);
or U15714 (N_15714,N_14012,N_13073);
nor U15715 (N_15715,N_14506,N_13510);
nor U15716 (N_15716,N_13524,N_12508);
nor U15717 (N_15717,N_13553,N_13448);
xnor U15718 (N_15718,N_13593,N_12691);
xor U15719 (N_15719,N_14489,N_13108);
and U15720 (N_15720,N_12807,N_13855);
and U15721 (N_15721,N_13748,N_14620);
or U15722 (N_15722,N_13398,N_14955);
nand U15723 (N_15723,N_14946,N_13833);
xnor U15724 (N_15724,N_13052,N_13313);
or U15725 (N_15725,N_14414,N_14531);
and U15726 (N_15726,N_13088,N_14660);
xnor U15727 (N_15727,N_14278,N_12969);
xnor U15728 (N_15728,N_13647,N_13109);
or U15729 (N_15729,N_12841,N_13611);
nor U15730 (N_15730,N_12500,N_14738);
nand U15731 (N_15731,N_13723,N_13239);
nor U15732 (N_15732,N_12752,N_13247);
nand U15733 (N_15733,N_13309,N_14394);
nor U15734 (N_15734,N_14542,N_12926);
nor U15735 (N_15735,N_14350,N_14517);
or U15736 (N_15736,N_13639,N_12921);
nand U15737 (N_15737,N_14899,N_12589);
and U15738 (N_15738,N_13699,N_13396);
xnor U15739 (N_15739,N_14549,N_12814);
nor U15740 (N_15740,N_13594,N_14615);
and U15741 (N_15741,N_14860,N_12919);
xor U15742 (N_15742,N_13503,N_12592);
nor U15743 (N_15743,N_13226,N_14749);
and U15744 (N_15744,N_14164,N_13337);
nor U15745 (N_15745,N_13515,N_12642);
xnor U15746 (N_15746,N_14672,N_14393);
nor U15747 (N_15747,N_13185,N_14448);
or U15748 (N_15748,N_13499,N_12654);
or U15749 (N_15749,N_13130,N_13147);
and U15750 (N_15750,N_12615,N_14646);
nand U15751 (N_15751,N_14525,N_14932);
nor U15752 (N_15752,N_12673,N_12993);
nand U15753 (N_15753,N_14963,N_13597);
or U15754 (N_15754,N_13211,N_13321);
or U15755 (N_15755,N_13853,N_13649);
or U15756 (N_15756,N_12544,N_13744);
xnor U15757 (N_15757,N_13602,N_13430);
nor U15758 (N_15758,N_13245,N_14261);
and U15759 (N_15759,N_14868,N_14579);
nand U15760 (N_15760,N_14978,N_13913);
nand U15761 (N_15761,N_14989,N_13725);
nor U15762 (N_15762,N_13866,N_14338);
xor U15763 (N_15763,N_12555,N_14323);
xnor U15764 (N_15764,N_12892,N_14925);
or U15765 (N_15765,N_14944,N_13662);
nand U15766 (N_15766,N_13315,N_14480);
nand U15767 (N_15767,N_14417,N_14706);
xor U15768 (N_15768,N_13875,N_13166);
or U15769 (N_15769,N_14426,N_14269);
nor U15770 (N_15770,N_13078,N_13729);
and U15771 (N_15771,N_12984,N_14547);
nand U15772 (N_15772,N_13151,N_12594);
nor U15773 (N_15773,N_14403,N_13939);
and U15774 (N_15774,N_13295,N_14535);
and U15775 (N_15775,N_13335,N_14018);
and U15776 (N_15776,N_14324,N_12655);
or U15777 (N_15777,N_12751,N_14231);
xor U15778 (N_15778,N_13252,N_14666);
xnor U15779 (N_15779,N_14566,N_13975);
nand U15780 (N_15780,N_14127,N_13640);
nor U15781 (N_15781,N_13585,N_14283);
nor U15782 (N_15782,N_13751,N_14810);
and U15783 (N_15783,N_14346,N_13873);
nor U15784 (N_15784,N_12521,N_12840);
nand U15785 (N_15785,N_14437,N_13281);
or U15786 (N_15786,N_13107,N_12881);
or U15787 (N_15787,N_13375,N_12902);
nor U15788 (N_15788,N_12849,N_13547);
nand U15789 (N_15789,N_14708,N_12526);
xor U15790 (N_15790,N_12983,N_14253);
nor U15791 (N_15791,N_13650,N_14510);
and U15792 (N_15792,N_13759,N_14379);
nand U15793 (N_15793,N_13001,N_14570);
or U15794 (N_15794,N_14309,N_13897);
or U15795 (N_15795,N_14169,N_13659);
nor U15796 (N_15796,N_13331,N_14664);
and U15797 (N_15797,N_12911,N_12509);
and U15798 (N_15798,N_12727,N_13463);
and U15799 (N_15799,N_12666,N_13674);
nor U15800 (N_15800,N_14039,N_14651);
nand U15801 (N_15801,N_14998,N_14494);
xor U15802 (N_15802,N_12988,N_12886);
nand U15803 (N_15803,N_14442,N_13458);
nor U15804 (N_15804,N_14225,N_12684);
nand U15805 (N_15805,N_13053,N_14661);
xor U15806 (N_15806,N_14653,N_13096);
or U15807 (N_15807,N_13820,N_13320);
and U15808 (N_15808,N_13953,N_13676);
xnor U15809 (N_15809,N_13854,N_13136);
nor U15810 (N_15810,N_13486,N_13093);
nor U15811 (N_15811,N_12831,N_13408);
or U15812 (N_15812,N_13621,N_14718);
xor U15813 (N_15813,N_13567,N_14821);
or U15814 (N_15814,N_14668,N_14213);
nor U15815 (N_15815,N_12882,N_13080);
and U15816 (N_15816,N_13799,N_12786);
xnor U15817 (N_15817,N_14882,N_14095);
or U15818 (N_15818,N_14145,N_13814);
and U15819 (N_15819,N_12759,N_14631);
nand U15820 (N_15820,N_14367,N_13236);
nor U15821 (N_15821,N_14726,N_14589);
and U15822 (N_15822,N_13118,N_12728);
xor U15823 (N_15823,N_12773,N_12837);
nand U15824 (N_15824,N_13049,N_13755);
and U15825 (N_15825,N_13272,N_14024);
nor U15826 (N_15826,N_14644,N_14267);
nand U15827 (N_15827,N_14049,N_13219);
xor U15828 (N_15828,N_13818,N_12874);
or U15829 (N_15829,N_14230,N_13102);
nor U15830 (N_15830,N_13344,N_12789);
xor U15831 (N_15831,N_13081,N_13962);
xor U15832 (N_15832,N_13616,N_14054);
or U15833 (N_15833,N_14327,N_13282);
nand U15834 (N_15834,N_14091,N_13863);
nor U15835 (N_15835,N_14139,N_14245);
or U15836 (N_15836,N_13712,N_14857);
or U15837 (N_15837,N_12539,N_12942);
or U15838 (N_15838,N_13260,N_13101);
or U15839 (N_15839,N_14967,N_14285);
nor U15840 (N_15840,N_12812,N_12651);
or U15841 (N_15841,N_13152,N_13110);
and U15842 (N_15842,N_14406,N_13076);
nor U15843 (N_15843,N_12867,N_14104);
nor U15844 (N_15844,N_12551,N_12788);
nor U15845 (N_15845,N_13986,N_13442);
nor U15846 (N_15846,N_12533,N_12818);
xor U15847 (N_15847,N_14061,N_13521);
nor U15848 (N_15848,N_13541,N_14216);
xnor U15849 (N_15849,N_13249,N_13238);
xor U15850 (N_15850,N_12762,N_13419);
xor U15851 (N_15851,N_12658,N_13250);
nand U15852 (N_15852,N_12915,N_13417);
nand U15853 (N_15853,N_13197,N_14319);
nand U15854 (N_15854,N_14098,N_12766);
and U15855 (N_15855,N_14173,N_13138);
nand U15856 (N_15856,N_13299,N_13574);
or U15857 (N_15857,N_13343,N_13354);
or U15858 (N_15858,N_12531,N_12645);
xnor U15859 (N_15859,N_12909,N_12520);
and U15860 (N_15860,N_14226,N_13919);
and U15861 (N_15861,N_13280,N_13623);
xor U15862 (N_15862,N_14248,N_12884);
xnor U15863 (N_15863,N_13606,N_14256);
or U15864 (N_15864,N_12851,N_13999);
and U15865 (N_15865,N_13003,N_13131);
nand U15866 (N_15866,N_12850,N_14347);
xor U15867 (N_15867,N_14533,N_14421);
and U15868 (N_15868,N_13484,N_14059);
xnor U15869 (N_15869,N_13922,N_14300);
nor U15870 (N_15870,N_14178,N_14433);
or U15871 (N_15871,N_14153,N_14928);
xor U15872 (N_15872,N_13129,N_14875);
nor U15873 (N_15873,N_14498,N_13468);
or U15874 (N_15874,N_14939,N_14450);
xor U15875 (N_15875,N_14468,N_14557);
xor U15876 (N_15876,N_13117,N_14559);
xnor U15877 (N_15877,N_12659,N_13128);
or U15878 (N_15878,N_14757,N_14514);
nor U15879 (N_15879,N_13858,N_14612);
or U15880 (N_15880,N_13456,N_13601);
nand U15881 (N_15881,N_12552,N_12671);
and U15882 (N_15882,N_13462,N_14970);
nor U15883 (N_15883,N_12724,N_12997);
xnor U15884 (N_15884,N_12774,N_13808);
nor U15885 (N_15885,N_13105,N_13664);
or U15886 (N_15886,N_12681,N_12864);
xnor U15887 (N_15887,N_13461,N_12541);
nand U15888 (N_15888,N_14146,N_13687);
nor U15889 (N_15889,N_13626,N_12747);
and U15890 (N_15890,N_12796,N_14493);
xor U15891 (N_15891,N_13903,N_14251);
nor U15892 (N_15892,N_13161,N_12725);
xnor U15893 (N_15893,N_14659,N_14008);
or U15894 (N_15894,N_14025,N_13492);
or U15895 (N_15895,N_14716,N_12767);
nand U15896 (N_15896,N_12861,N_12947);
or U15897 (N_15897,N_14960,N_14933);
nor U15898 (N_15898,N_14185,N_13645);
nor U15899 (N_15899,N_12933,N_14544);
nand U15900 (N_15900,N_14783,N_14771);
or U15901 (N_15901,N_14047,N_14700);
nand U15902 (N_15902,N_13523,N_12602);
nand U15903 (N_15903,N_12920,N_12967);
and U15904 (N_15904,N_14405,N_14826);
or U15905 (N_15905,N_14816,N_13188);
nand U15906 (N_15906,N_13673,N_13914);
or U15907 (N_15907,N_14284,N_14020);
or U15908 (N_15908,N_13832,N_13972);
or U15909 (N_15909,N_14817,N_13941);
or U15910 (N_15910,N_12716,N_13619);
and U15911 (N_15911,N_14607,N_12836);
nor U15912 (N_15912,N_13928,N_14446);
nand U15913 (N_15913,N_13598,N_14096);
xor U15914 (N_15914,N_13421,N_13527);
xor U15915 (N_15915,N_13878,N_14006);
or U15916 (N_15916,N_12980,N_14755);
and U15917 (N_15917,N_14381,N_13038);
xnor U15918 (N_15918,N_13749,N_13534);
or U15919 (N_15919,N_14769,N_13810);
and U15920 (N_15920,N_13537,N_13369);
or U15921 (N_15921,N_13159,N_14068);
xnor U15922 (N_15922,N_14862,N_12699);
or U15923 (N_15923,N_14979,N_14427);
nand U15924 (N_15924,N_12662,N_13950);
or U15925 (N_15925,N_13794,N_14435);
nand U15926 (N_15926,N_13148,N_14197);
and U15927 (N_15927,N_14828,N_12880);
or U15928 (N_15928,N_12517,N_13924);
or U15929 (N_15929,N_14903,N_13403);
or U15930 (N_15930,N_14438,N_14206);
or U15931 (N_15931,N_14371,N_13471);
xnor U15932 (N_15932,N_13042,N_13296);
nor U15933 (N_15933,N_13816,N_14151);
xnor U15934 (N_15934,N_12656,N_13525);
xor U15935 (N_15935,N_13387,N_14307);
nor U15936 (N_15936,N_14592,N_12935);
and U15937 (N_15937,N_13508,N_13787);
and U15938 (N_15938,N_13173,N_13216);
or U15939 (N_15939,N_14694,N_14676);
and U15940 (N_15940,N_13930,N_14937);
nor U15941 (N_15941,N_13731,N_13609);
and U15942 (N_15942,N_12714,N_13466);
xor U15943 (N_15943,N_13409,N_14971);
xnor U15944 (N_15944,N_13538,N_13558);
or U15945 (N_15945,N_13465,N_14591);
nor U15946 (N_15946,N_13336,N_14467);
nand U15947 (N_15947,N_13089,N_12663);
nor U15948 (N_15948,N_14931,N_14977);
or U15949 (N_15949,N_12632,N_12574);
nor U15950 (N_15950,N_13700,N_12970);
and U15951 (N_15951,N_14475,N_13741);
xnor U15952 (N_15952,N_14555,N_13836);
and U15953 (N_15953,N_13056,N_13017);
and U15954 (N_15954,N_14896,N_14842);
xor U15955 (N_15955,N_14534,N_13779);
nand U15956 (N_15956,N_12826,N_12740);
nor U15957 (N_15957,N_14814,N_13980);
or U15958 (N_15958,N_14431,N_14848);
nand U15959 (N_15959,N_14161,N_12721);
nand U15960 (N_15960,N_14725,N_13441);
xnor U15961 (N_15961,N_13618,N_13507);
or U15962 (N_15962,N_14112,N_14815);
xor U15963 (N_15963,N_12708,N_13513);
or U15964 (N_15964,N_13984,N_14956);
or U15965 (N_15965,N_13485,N_12746);
xnor U15966 (N_15966,N_12636,N_13509);
nand U15967 (N_15967,N_14205,N_14523);
xnor U15968 (N_15968,N_13116,N_13531);
nand U15969 (N_15969,N_12553,N_13827);
or U15970 (N_15970,N_13242,N_13822);
and U15971 (N_15971,N_12549,N_14791);
or U15972 (N_15972,N_14649,N_14840);
xnor U15973 (N_15973,N_14255,N_13153);
nor U15974 (N_15974,N_12890,N_13377);
nor U15975 (N_15975,N_12571,N_13916);
xor U15976 (N_15976,N_14982,N_13278);
xor U15977 (N_15977,N_14884,N_13576);
nand U15978 (N_15978,N_14996,N_13364);
nor U15979 (N_15979,N_12584,N_14390);
or U15980 (N_15980,N_13180,N_14443);
nor U15981 (N_15981,N_13092,N_12835);
or U15982 (N_15982,N_14479,N_12558);
and U15983 (N_15983,N_13126,N_14214);
nor U15984 (N_15984,N_13584,N_13951);
xor U15985 (N_15985,N_14850,N_14521);
or U15986 (N_15986,N_12537,N_13937);
or U15987 (N_15987,N_14345,N_13232);
nand U15988 (N_15988,N_14429,N_12729);
or U15989 (N_15989,N_14074,N_13952);
nand U15990 (N_15990,N_12546,N_14476);
nand U15991 (N_15991,N_13220,N_12605);
nor U15992 (N_15992,N_14808,N_14657);
nor U15993 (N_15993,N_13498,N_13812);
nor U15994 (N_15994,N_12948,N_13005);
xor U15995 (N_15995,N_14144,N_12987);
nor U15996 (N_15996,N_12664,N_14325);
nand U15997 (N_15997,N_13229,N_14259);
nand U15998 (N_15998,N_12952,N_13655);
nand U15999 (N_15999,N_13877,N_13763);
or U16000 (N_16000,N_13106,N_14457);
xnor U16001 (N_16001,N_13473,N_13940);
and U16002 (N_16002,N_14463,N_14611);
xnor U16003 (N_16003,N_14363,N_14374);
or U16004 (N_16004,N_14975,N_14260);
nand U16005 (N_16005,N_14041,N_14936);
and U16006 (N_16006,N_14196,N_13927);
and U16007 (N_16007,N_13162,N_14123);
nor U16008 (N_16008,N_14088,N_14910);
xnor U16009 (N_16009,N_12770,N_14155);
nor U16010 (N_16010,N_14116,N_12844);
or U16011 (N_16011,N_13895,N_12698);
or U16012 (N_16012,N_14887,N_13407);
nor U16013 (N_16013,N_12871,N_12635);
nor U16014 (N_16014,N_13202,N_14066);
nor U16015 (N_16015,N_14554,N_13958);
xnor U16016 (N_16016,N_14886,N_13707);
nand U16017 (N_16017,N_13483,N_14296);
nand U16018 (N_16018,N_14223,N_13452);
xnor U16019 (N_16019,N_14254,N_13533);
or U16020 (N_16020,N_14424,N_13307);
nand U16021 (N_16021,N_14687,N_13613);
xnor U16022 (N_16022,N_14376,N_13970);
nor U16023 (N_16023,N_13413,N_13189);
xnor U16024 (N_16024,N_14943,N_12563);
and U16025 (N_16025,N_12918,N_14215);
nor U16026 (N_16026,N_12619,N_14488);
or U16027 (N_16027,N_13719,N_14804);
or U16028 (N_16028,N_12949,N_13221);
nor U16029 (N_16029,N_13172,N_14461);
nor U16030 (N_16030,N_14208,N_12825);
xnor U16031 (N_16031,N_14114,N_12950);
nand U16032 (N_16032,N_12625,N_14001);
nor U16033 (N_16033,N_13355,N_14938);
xor U16034 (N_16034,N_13882,N_13099);
and U16035 (N_16035,N_14277,N_14564);
nand U16036 (N_16036,N_13535,N_12617);
or U16037 (N_16037,N_14090,N_13384);
xor U16038 (N_16038,N_14062,N_14588);
nand U16039 (N_16039,N_14748,N_14369);
nor U16040 (N_16040,N_12925,N_14806);
or U16041 (N_16041,N_14702,N_13572);
or U16042 (N_16042,N_13243,N_12781);
xor U16043 (N_16043,N_12680,N_13959);
or U16044 (N_16044,N_14211,N_14530);
or U16045 (N_16045,N_14869,N_12513);
and U16046 (N_16046,N_14540,N_14108);
or U16047 (N_16047,N_12908,N_13423);
or U16048 (N_16048,N_12910,N_14511);
xnor U16049 (N_16049,N_12891,N_13514);
nand U16050 (N_16050,N_14873,N_13578);
xnor U16051 (N_16051,N_12953,N_13312);
nand U16052 (N_16052,N_14038,N_13695);
or U16053 (N_16053,N_13680,N_13228);
xnor U16054 (N_16054,N_13844,N_12711);
xor U16055 (N_16055,N_13146,N_14670);
or U16056 (N_16056,N_14399,N_14658);
xor U16057 (N_16057,N_14537,N_14987);
and U16058 (N_16058,N_13976,N_12966);
nand U16059 (N_16059,N_13264,N_14515);
and U16060 (N_16060,N_14310,N_14623);
nand U16061 (N_16061,N_14774,N_13347);
or U16062 (N_16062,N_14149,N_12516);
nand U16063 (N_16063,N_14563,N_14032);
nand U16064 (N_16064,N_12693,N_13023);
or U16065 (N_16065,N_13176,N_13433);
nor U16066 (N_16066,N_14630,N_13506);
or U16067 (N_16067,N_14076,N_14913);
or U16068 (N_16068,N_13561,N_12577);
nand U16069 (N_16069,N_12846,N_12742);
xor U16070 (N_16070,N_12536,N_14865);
xor U16071 (N_16071,N_14030,N_12937);
and U16072 (N_16072,N_14274,N_13511);
nor U16073 (N_16073,N_12843,N_13996);
nor U16074 (N_16074,N_14258,N_12977);
xor U16075 (N_16075,N_13234,N_12870);
or U16076 (N_16076,N_14686,N_13981);
nor U16077 (N_16077,N_12616,N_14997);
and U16078 (N_16078,N_14120,N_14364);
nand U16079 (N_16079,N_14502,N_13504);
nor U16080 (N_16080,N_13758,N_13768);
nand U16081 (N_16081,N_13436,N_13237);
nor U16082 (N_16082,N_13637,N_14822);
nand U16083 (N_16083,N_14447,N_13889);
nor U16084 (N_16084,N_13175,N_13904);
nand U16085 (N_16085,N_13119,N_13709);
and U16086 (N_16086,N_13760,N_14316);
or U16087 (N_16087,N_14335,N_14858);
nor U16088 (N_16088,N_13519,N_13287);
nor U16089 (N_16089,N_14950,N_13715);
or U16090 (N_16090,N_13018,N_14751);
and U16091 (N_16091,N_13622,N_14923);
nand U16092 (N_16092,N_13841,N_13181);
nor U16093 (N_16093,N_14785,N_13845);
or U16094 (N_16094,N_13605,N_12715);
or U16095 (N_16095,N_14244,N_12590);
nand U16096 (N_16096,N_13444,N_13035);
and U16097 (N_16097,N_14921,N_14240);
or U16098 (N_16098,N_13244,N_12598);
nor U16099 (N_16099,N_12872,N_12609);
xor U16100 (N_16100,N_14052,N_14209);
and U16101 (N_16101,N_13663,N_13671);
xor U16102 (N_16102,N_14229,N_13993);
and U16103 (N_16103,N_14717,N_14492);
or U16104 (N_16104,N_12719,N_14045);
xnor U16105 (N_16105,N_14235,N_13085);
or U16106 (N_16106,N_12677,N_12683);
or U16107 (N_16107,N_13694,N_14452);
nand U16108 (N_16108,N_12718,N_12991);
xor U16109 (N_16109,N_12717,N_13016);
nand U16110 (N_16110,N_14331,N_14558);
nor U16111 (N_16111,N_12860,N_12769);
nor U16112 (N_16112,N_14412,N_14601);
or U16113 (N_16113,N_13058,N_14867);
xnor U16114 (N_16114,N_14015,N_12687);
nor U16115 (N_16115,N_13333,N_12612);
xnor U16116 (N_16116,N_14780,N_12527);
and U16117 (N_16117,N_14290,N_13070);
and U16118 (N_16118,N_13559,N_13149);
or U16119 (N_16119,N_14306,N_13789);
or U16120 (N_16120,N_13297,N_13200);
nor U16121 (N_16121,N_14464,N_13261);
or U16122 (N_16122,N_14086,N_14640);
xor U16123 (N_16123,N_13267,N_13635);
nand U16124 (N_16124,N_12548,N_12566);
nor U16125 (N_16125,N_14851,N_12830);
nand U16126 (N_16126,N_12596,N_13630);
nand U16127 (N_16127,N_13933,N_14779);
xor U16128 (N_16128,N_14712,N_12834);
and U16129 (N_16129,N_13684,N_14643);
nand U16130 (N_16130,N_13713,N_12676);
or U16131 (N_16131,N_13945,N_14029);
or U16132 (N_16132,N_14954,N_13539);
nand U16133 (N_16133,N_14752,N_14512);
or U16134 (N_16134,N_12946,N_14617);
nand U16135 (N_16135,N_14605,N_13821);
nand U16136 (N_16136,N_13399,N_14378);
or U16137 (N_16137,N_14434,N_13284);
nand U16138 (N_16138,N_14487,N_14616);
and U16139 (N_16139,N_14019,N_13054);
or U16140 (N_16140,N_13027,N_13718);
nor U16141 (N_16141,N_14470,N_14023);
nor U16142 (N_16142,N_13614,N_14107);
and U16143 (N_16143,N_12608,N_14481);
and U16144 (N_16144,N_14125,N_12591);
nor U16145 (N_16145,N_13706,N_13363);
and U16146 (N_16146,N_14513,N_13957);
xor U16147 (N_16147,N_12630,N_13608);
or U16148 (N_16148,N_13257,N_13434);
and U16149 (N_16149,N_12956,N_12816);
or U16150 (N_16150,N_14892,N_12669);
xnor U16151 (N_16151,N_12940,N_13888);
and U16152 (N_16152,N_12801,N_12732);
nor U16153 (N_16153,N_14990,N_12833);
nand U16154 (N_16154,N_14177,N_13815);
nand U16155 (N_16155,N_13773,N_13520);
xnor U16156 (N_16156,N_12523,N_14129);
xor U16157 (N_16157,N_13540,N_13987);
nor U16158 (N_16158,N_12893,N_13793);
nor U16159 (N_16159,N_13378,N_14396);
nor U16160 (N_16160,N_14968,N_13968);
or U16161 (N_16161,N_12559,N_14580);
and U16162 (N_16162,N_14176,N_13880);
nor U16163 (N_16163,N_12798,N_14491);
nand U16164 (N_16164,N_13979,N_13555);
xor U16165 (N_16165,N_12631,N_13412);
and U16166 (N_16166,N_13467,N_13686);
and U16167 (N_16167,N_13400,N_14870);
nor U16168 (N_16168,N_13600,N_12780);
or U16169 (N_16169,N_12829,N_13270);
or U16170 (N_16170,N_14458,N_13274);
and U16171 (N_16171,N_13643,N_14321);
nor U16172 (N_16172,N_14993,N_13658);
and U16173 (N_16173,N_14729,N_14577);
or U16174 (N_16174,N_14377,N_14193);
nor U16175 (N_16175,N_14199,N_13420);
and U16176 (N_16176,N_13213,N_12731);
xnor U16177 (N_16177,N_13427,N_13496);
or U16178 (N_16178,N_14703,N_12519);
nand U16179 (N_16179,N_13322,N_14317);
and U16180 (N_16180,N_13276,N_13721);
nand U16181 (N_16181,N_13591,N_12795);
or U16182 (N_16182,N_14348,N_12679);
nor U16183 (N_16183,N_13925,N_14080);
or U16184 (N_16184,N_14836,N_12819);
and U16185 (N_16185,N_13690,N_13218);
nor U16186 (N_16186,N_13440,N_12941);
and U16187 (N_16187,N_14760,N_13100);
nor U16188 (N_16188,N_12895,N_12702);
xor U16189 (N_16189,N_12998,N_14058);
xor U16190 (N_16190,N_14180,N_14351);
xnor U16191 (N_16191,N_13628,N_14017);
xor U16192 (N_16192,N_12665,N_14773);
and U16193 (N_16193,N_13921,N_12668);
nand U16194 (N_16194,N_14233,N_12916);
nand U16195 (N_16195,N_14991,N_14981);
xnor U16196 (N_16196,N_12823,N_14688);
nor U16197 (N_16197,N_14482,N_14130);
xor U16198 (N_16198,N_14907,N_14303);
xor U16199 (N_16199,N_14337,N_13592);
nor U16200 (N_16200,N_14754,N_14581);
nor U16201 (N_16201,N_13203,N_13714);
or U16202 (N_16202,N_14148,N_14759);
xnor U16203 (N_16203,N_14287,N_13936);
nor U16204 (N_16204,N_14281,N_13127);
xor U16205 (N_16205,N_14186,N_14313);
and U16206 (N_16206,N_13657,N_14906);
and U16207 (N_16207,N_13892,N_14905);
and U16208 (N_16208,N_13350,N_13266);
and U16209 (N_16209,N_14800,N_13031);
xor U16210 (N_16210,N_14387,N_14057);
and U16211 (N_16211,N_13124,N_13283);
xnor U16212 (N_16212,N_14200,N_13595);
nor U16213 (N_16213,N_13989,N_12808);
nand U16214 (N_16214,N_14028,N_12982);
and U16215 (N_16215,N_14553,N_14958);
and U16216 (N_16216,N_12938,N_13954);
nand U16217 (N_16217,N_13258,N_14711);
nor U16218 (N_16218,N_14386,N_14060);
nor U16219 (N_16219,N_14063,N_14691);
or U16220 (N_16220,N_12986,N_14578);
nand U16221 (N_16221,N_13800,N_13965);
xnor U16222 (N_16222,N_14469,N_14100);
or U16223 (N_16223,N_14764,N_14768);
nor U16224 (N_16224,N_13912,N_13756);
and U16225 (N_16225,N_13424,N_13406);
or U16226 (N_16226,N_12628,N_13920);
xor U16227 (N_16227,N_14775,N_12760);
nor U16228 (N_16228,N_12650,N_13791);
xor U16229 (N_16229,N_14770,N_13978);
xor U16230 (N_16230,N_12597,N_12885);
or U16231 (N_16231,N_13859,N_12820);
and U16232 (N_16232,N_13861,N_13905);
xnor U16233 (N_16233,N_14322,N_12923);
nor U16234 (N_16234,N_13918,N_12971);
or U16235 (N_16235,N_13293,N_13991);
nand U16236 (N_16236,N_13340,N_14220);
nand U16237 (N_16237,N_14747,N_14926);
xnor U16238 (N_16238,N_13776,N_13046);
and U16239 (N_16239,N_13253,N_12626);
xor U16240 (N_16240,N_13273,N_14940);
nor U16241 (N_16241,N_13304,N_12821);
nor U16242 (N_16242,N_13285,N_13997);
nand U16243 (N_16243,N_14777,N_13992);
nand U16244 (N_16244,N_14874,N_12545);
and U16245 (N_16245,N_12913,N_13443);
and U16246 (N_16246,N_12644,N_13395);
or U16247 (N_16247,N_13305,N_13961);
or U16248 (N_16248,N_13973,N_14904);
or U16249 (N_16249,N_14807,N_14548);
xor U16250 (N_16250,N_14263,N_14822);
xnor U16251 (N_16251,N_13003,N_14824);
or U16252 (N_16252,N_13689,N_14182);
nor U16253 (N_16253,N_14273,N_12872);
nand U16254 (N_16254,N_14477,N_12826);
nand U16255 (N_16255,N_13994,N_14310);
xnor U16256 (N_16256,N_13850,N_13523);
or U16257 (N_16257,N_14297,N_13502);
or U16258 (N_16258,N_13687,N_12948);
nor U16259 (N_16259,N_13637,N_13963);
and U16260 (N_16260,N_14720,N_13168);
nand U16261 (N_16261,N_12908,N_12886);
nor U16262 (N_16262,N_12883,N_13950);
xor U16263 (N_16263,N_12941,N_12907);
and U16264 (N_16264,N_14380,N_13236);
nor U16265 (N_16265,N_14488,N_13508);
xnor U16266 (N_16266,N_13149,N_13332);
and U16267 (N_16267,N_14239,N_13137);
and U16268 (N_16268,N_12703,N_13090);
or U16269 (N_16269,N_13472,N_13947);
or U16270 (N_16270,N_13575,N_13010);
nor U16271 (N_16271,N_13599,N_13785);
or U16272 (N_16272,N_13610,N_14708);
and U16273 (N_16273,N_14957,N_14012);
nand U16274 (N_16274,N_14550,N_13047);
nor U16275 (N_16275,N_14027,N_13762);
or U16276 (N_16276,N_12832,N_14961);
nand U16277 (N_16277,N_13645,N_14865);
xor U16278 (N_16278,N_13236,N_13673);
or U16279 (N_16279,N_14991,N_14136);
nand U16280 (N_16280,N_14664,N_13159);
nand U16281 (N_16281,N_13501,N_13379);
nor U16282 (N_16282,N_12756,N_13148);
xnor U16283 (N_16283,N_12905,N_14958);
xnor U16284 (N_16284,N_14750,N_13960);
xor U16285 (N_16285,N_14170,N_14748);
and U16286 (N_16286,N_14857,N_14742);
or U16287 (N_16287,N_14638,N_14999);
nor U16288 (N_16288,N_14954,N_12786);
xnor U16289 (N_16289,N_12561,N_13602);
and U16290 (N_16290,N_14111,N_13411);
nor U16291 (N_16291,N_13972,N_12629);
nand U16292 (N_16292,N_12974,N_14246);
nand U16293 (N_16293,N_13549,N_14067);
nand U16294 (N_16294,N_12825,N_14088);
xor U16295 (N_16295,N_13597,N_13024);
nand U16296 (N_16296,N_14987,N_14686);
nor U16297 (N_16297,N_14755,N_12838);
nor U16298 (N_16298,N_13281,N_14076);
nor U16299 (N_16299,N_13931,N_14807);
xor U16300 (N_16300,N_14318,N_12683);
or U16301 (N_16301,N_14779,N_12804);
and U16302 (N_16302,N_13298,N_14474);
nor U16303 (N_16303,N_13815,N_14596);
or U16304 (N_16304,N_14052,N_14592);
xor U16305 (N_16305,N_14982,N_12627);
xnor U16306 (N_16306,N_12988,N_13629);
nor U16307 (N_16307,N_12597,N_13805);
nand U16308 (N_16308,N_14850,N_13408);
and U16309 (N_16309,N_13323,N_12912);
xor U16310 (N_16310,N_13222,N_14916);
xnor U16311 (N_16311,N_12831,N_13995);
or U16312 (N_16312,N_13217,N_12520);
xnor U16313 (N_16313,N_13295,N_13030);
nor U16314 (N_16314,N_13083,N_13757);
or U16315 (N_16315,N_12586,N_14301);
and U16316 (N_16316,N_14050,N_14449);
and U16317 (N_16317,N_13823,N_14477);
xnor U16318 (N_16318,N_12907,N_12790);
or U16319 (N_16319,N_13428,N_13638);
or U16320 (N_16320,N_14236,N_13317);
nor U16321 (N_16321,N_12629,N_14414);
nand U16322 (N_16322,N_13612,N_14295);
xor U16323 (N_16323,N_14719,N_13435);
nand U16324 (N_16324,N_14068,N_13448);
and U16325 (N_16325,N_14729,N_14557);
and U16326 (N_16326,N_14623,N_13296);
nor U16327 (N_16327,N_14549,N_14657);
xnor U16328 (N_16328,N_13331,N_13679);
xnor U16329 (N_16329,N_13755,N_13051);
nand U16330 (N_16330,N_14284,N_14272);
nand U16331 (N_16331,N_13003,N_13090);
and U16332 (N_16332,N_13528,N_13479);
nand U16333 (N_16333,N_14122,N_13502);
nor U16334 (N_16334,N_14415,N_14249);
nand U16335 (N_16335,N_14482,N_13434);
xor U16336 (N_16336,N_14213,N_12678);
xnor U16337 (N_16337,N_12564,N_14805);
nand U16338 (N_16338,N_14723,N_13104);
and U16339 (N_16339,N_12566,N_14544);
nand U16340 (N_16340,N_12615,N_13121);
or U16341 (N_16341,N_14995,N_14357);
nand U16342 (N_16342,N_14133,N_14158);
xnor U16343 (N_16343,N_13521,N_12779);
nand U16344 (N_16344,N_14403,N_14593);
or U16345 (N_16345,N_13656,N_13652);
or U16346 (N_16346,N_14379,N_14905);
xor U16347 (N_16347,N_12649,N_12885);
or U16348 (N_16348,N_13082,N_14286);
and U16349 (N_16349,N_14853,N_14728);
and U16350 (N_16350,N_13143,N_14075);
or U16351 (N_16351,N_14840,N_13771);
and U16352 (N_16352,N_13040,N_13834);
or U16353 (N_16353,N_14543,N_12905);
nand U16354 (N_16354,N_13027,N_14613);
xor U16355 (N_16355,N_14328,N_13758);
and U16356 (N_16356,N_13538,N_13178);
and U16357 (N_16357,N_14293,N_13150);
nand U16358 (N_16358,N_14635,N_14086);
nor U16359 (N_16359,N_14521,N_14517);
nand U16360 (N_16360,N_13859,N_14164);
and U16361 (N_16361,N_12798,N_14647);
xor U16362 (N_16362,N_13333,N_14562);
and U16363 (N_16363,N_12545,N_12912);
or U16364 (N_16364,N_13286,N_12806);
and U16365 (N_16365,N_13274,N_13935);
nand U16366 (N_16366,N_13141,N_14901);
nand U16367 (N_16367,N_12525,N_14598);
nand U16368 (N_16368,N_13927,N_14437);
xor U16369 (N_16369,N_13267,N_14546);
or U16370 (N_16370,N_14930,N_13211);
or U16371 (N_16371,N_13832,N_12523);
or U16372 (N_16372,N_12561,N_12740);
xnor U16373 (N_16373,N_14059,N_13642);
nor U16374 (N_16374,N_12794,N_12782);
nand U16375 (N_16375,N_13337,N_14591);
nor U16376 (N_16376,N_14744,N_13768);
nor U16377 (N_16377,N_14736,N_14323);
nor U16378 (N_16378,N_12532,N_13988);
nor U16379 (N_16379,N_14718,N_14149);
nand U16380 (N_16380,N_14967,N_14384);
nand U16381 (N_16381,N_14229,N_14206);
or U16382 (N_16382,N_12633,N_14948);
nand U16383 (N_16383,N_12979,N_12828);
or U16384 (N_16384,N_14155,N_13665);
and U16385 (N_16385,N_14481,N_13626);
and U16386 (N_16386,N_14599,N_14914);
xnor U16387 (N_16387,N_13829,N_12759);
xor U16388 (N_16388,N_13416,N_14678);
nor U16389 (N_16389,N_14614,N_13179);
and U16390 (N_16390,N_13853,N_14932);
nand U16391 (N_16391,N_13678,N_12745);
nand U16392 (N_16392,N_13255,N_14195);
or U16393 (N_16393,N_12534,N_12721);
nor U16394 (N_16394,N_14214,N_14854);
nand U16395 (N_16395,N_12973,N_12903);
xor U16396 (N_16396,N_14557,N_12931);
nand U16397 (N_16397,N_14181,N_13005);
or U16398 (N_16398,N_12676,N_14965);
and U16399 (N_16399,N_13718,N_13468);
and U16400 (N_16400,N_12699,N_13168);
xor U16401 (N_16401,N_14506,N_14537);
nand U16402 (N_16402,N_14046,N_14527);
or U16403 (N_16403,N_12779,N_13490);
nand U16404 (N_16404,N_13692,N_13640);
xor U16405 (N_16405,N_13327,N_14709);
or U16406 (N_16406,N_13970,N_12890);
or U16407 (N_16407,N_14552,N_14439);
and U16408 (N_16408,N_13204,N_13241);
or U16409 (N_16409,N_13031,N_13200);
or U16410 (N_16410,N_13578,N_12822);
nand U16411 (N_16411,N_13462,N_12806);
and U16412 (N_16412,N_14681,N_14760);
nand U16413 (N_16413,N_13802,N_14493);
nor U16414 (N_16414,N_13638,N_13677);
and U16415 (N_16415,N_12941,N_14998);
or U16416 (N_16416,N_14303,N_13077);
nor U16417 (N_16417,N_13299,N_13200);
or U16418 (N_16418,N_12662,N_13492);
xnor U16419 (N_16419,N_14070,N_14660);
and U16420 (N_16420,N_14921,N_14919);
xnor U16421 (N_16421,N_14331,N_14313);
nor U16422 (N_16422,N_13647,N_14053);
xor U16423 (N_16423,N_12813,N_12548);
nand U16424 (N_16424,N_13416,N_14454);
and U16425 (N_16425,N_14453,N_14732);
or U16426 (N_16426,N_12513,N_13193);
nor U16427 (N_16427,N_14747,N_14470);
xnor U16428 (N_16428,N_14738,N_12700);
xor U16429 (N_16429,N_14336,N_12569);
xnor U16430 (N_16430,N_13349,N_13746);
and U16431 (N_16431,N_14119,N_14348);
and U16432 (N_16432,N_14221,N_14714);
nand U16433 (N_16433,N_13540,N_13819);
nand U16434 (N_16434,N_12944,N_14115);
nor U16435 (N_16435,N_13993,N_14682);
nand U16436 (N_16436,N_14450,N_14363);
or U16437 (N_16437,N_13757,N_13291);
and U16438 (N_16438,N_14363,N_12852);
xor U16439 (N_16439,N_14879,N_14504);
or U16440 (N_16440,N_14016,N_13683);
nor U16441 (N_16441,N_13738,N_13019);
or U16442 (N_16442,N_14166,N_14027);
xor U16443 (N_16443,N_14357,N_14185);
xor U16444 (N_16444,N_13594,N_14255);
and U16445 (N_16445,N_12649,N_13831);
nor U16446 (N_16446,N_12564,N_13841);
or U16447 (N_16447,N_12628,N_13258);
nand U16448 (N_16448,N_13164,N_13159);
or U16449 (N_16449,N_14956,N_14101);
nor U16450 (N_16450,N_13059,N_12909);
xnor U16451 (N_16451,N_12688,N_12912);
and U16452 (N_16452,N_14866,N_14055);
xor U16453 (N_16453,N_13322,N_14731);
nand U16454 (N_16454,N_14031,N_13551);
and U16455 (N_16455,N_14218,N_13099);
and U16456 (N_16456,N_12580,N_13872);
or U16457 (N_16457,N_14613,N_14107);
nor U16458 (N_16458,N_13210,N_14141);
and U16459 (N_16459,N_13834,N_12962);
xnor U16460 (N_16460,N_12876,N_13003);
nor U16461 (N_16461,N_13011,N_13512);
xor U16462 (N_16462,N_14852,N_14950);
or U16463 (N_16463,N_13218,N_12787);
or U16464 (N_16464,N_14528,N_13537);
nor U16465 (N_16465,N_14620,N_12784);
and U16466 (N_16466,N_13480,N_13774);
xnor U16467 (N_16467,N_14421,N_14474);
or U16468 (N_16468,N_12553,N_13404);
and U16469 (N_16469,N_13840,N_14739);
nand U16470 (N_16470,N_14614,N_14172);
xor U16471 (N_16471,N_13165,N_13640);
or U16472 (N_16472,N_14189,N_13570);
xor U16473 (N_16473,N_12578,N_13803);
xnor U16474 (N_16474,N_14487,N_14511);
nor U16475 (N_16475,N_14319,N_14369);
nand U16476 (N_16476,N_12654,N_13339);
nand U16477 (N_16477,N_12531,N_14829);
nand U16478 (N_16478,N_12973,N_13082);
xnor U16479 (N_16479,N_14324,N_13793);
nand U16480 (N_16480,N_14831,N_14534);
or U16481 (N_16481,N_13207,N_13568);
nand U16482 (N_16482,N_14813,N_13170);
or U16483 (N_16483,N_14889,N_12853);
xnor U16484 (N_16484,N_14430,N_14978);
and U16485 (N_16485,N_12725,N_12590);
or U16486 (N_16486,N_14513,N_14450);
xnor U16487 (N_16487,N_14946,N_13393);
and U16488 (N_16488,N_14715,N_12757);
nor U16489 (N_16489,N_14748,N_14630);
nor U16490 (N_16490,N_14877,N_12926);
nor U16491 (N_16491,N_13595,N_12571);
and U16492 (N_16492,N_14306,N_14512);
and U16493 (N_16493,N_14906,N_12547);
or U16494 (N_16494,N_13507,N_12961);
nor U16495 (N_16495,N_13804,N_14622);
nor U16496 (N_16496,N_14116,N_14249);
nand U16497 (N_16497,N_14060,N_12577);
nand U16498 (N_16498,N_13645,N_13447);
nor U16499 (N_16499,N_12643,N_13349);
nand U16500 (N_16500,N_14351,N_13705);
nor U16501 (N_16501,N_12668,N_13501);
or U16502 (N_16502,N_14038,N_14132);
or U16503 (N_16503,N_12766,N_13973);
or U16504 (N_16504,N_13302,N_14032);
or U16505 (N_16505,N_13980,N_13866);
nand U16506 (N_16506,N_14021,N_14662);
xor U16507 (N_16507,N_13551,N_14989);
and U16508 (N_16508,N_12698,N_12637);
xnor U16509 (N_16509,N_14574,N_13355);
xor U16510 (N_16510,N_14894,N_14121);
nand U16511 (N_16511,N_12564,N_12727);
and U16512 (N_16512,N_14132,N_13591);
and U16513 (N_16513,N_13308,N_13963);
nor U16514 (N_16514,N_12669,N_13631);
nor U16515 (N_16515,N_12538,N_14321);
and U16516 (N_16516,N_13070,N_14486);
or U16517 (N_16517,N_14310,N_12933);
or U16518 (N_16518,N_13162,N_13211);
and U16519 (N_16519,N_14298,N_13253);
or U16520 (N_16520,N_14569,N_14189);
nand U16521 (N_16521,N_14628,N_12942);
or U16522 (N_16522,N_13964,N_13396);
or U16523 (N_16523,N_14365,N_13778);
or U16524 (N_16524,N_14635,N_13929);
nand U16525 (N_16525,N_12628,N_14816);
nand U16526 (N_16526,N_14693,N_14823);
nor U16527 (N_16527,N_13264,N_13185);
nand U16528 (N_16528,N_12647,N_14389);
and U16529 (N_16529,N_14883,N_14207);
xor U16530 (N_16530,N_12928,N_13652);
nor U16531 (N_16531,N_14190,N_14656);
and U16532 (N_16532,N_14446,N_13903);
or U16533 (N_16533,N_13630,N_12671);
xnor U16534 (N_16534,N_12725,N_13486);
nand U16535 (N_16535,N_13147,N_12979);
xor U16536 (N_16536,N_12748,N_12945);
xor U16537 (N_16537,N_13427,N_13686);
nor U16538 (N_16538,N_14866,N_13942);
or U16539 (N_16539,N_13431,N_14360);
nor U16540 (N_16540,N_13799,N_14260);
nand U16541 (N_16541,N_13712,N_14372);
xor U16542 (N_16542,N_12941,N_14986);
nand U16543 (N_16543,N_14278,N_13179);
nor U16544 (N_16544,N_13620,N_14086);
or U16545 (N_16545,N_14114,N_13863);
nor U16546 (N_16546,N_14939,N_12932);
xor U16547 (N_16547,N_13585,N_13812);
nor U16548 (N_16548,N_14071,N_13632);
nand U16549 (N_16549,N_14276,N_13122);
xor U16550 (N_16550,N_12757,N_14772);
nand U16551 (N_16551,N_12606,N_12943);
and U16552 (N_16552,N_13458,N_13552);
nand U16553 (N_16553,N_13907,N_13836);
or U16554 (N_16554,N_14477,N_14184);
or U16555 (N_16555,N_14755,N_14813);
nor U16556 (N_16556,N_14777,N_13887);
nand U16557 (N_16557,N_13519,N_13964);
and U16558 (N_16558,N_14178,N_13277);
and U16559 (N_16559,N_14525,N_13988);
nand U16560 (N_16560,N_12545,N_14413);
and U16561 (N_16561,N_14893,N_13477);
and U16562 (N_16562,N_13063,N_12864);
or U16563 (N_16563,N_14683,N_14160);
nand U16564 (N_16564,N_14416,N_12900);
or U16565 (N_16565,N_14388,N_12978);
nor U16566 (N_16566,N_14770,N_13149);
nand U16567 (N_16567,N_14635,N_14169);
nor U16568 (N_16568,N_14130,N_13182);
and U16569 (N_16569,N_14290,N_14266);
nor U16570 (N_16570,N_13885,N_12730);
and U16571 (N_16571,N_13608,N_14703);
or U16572 (N_16572,N_13970,N_13003);
and U16573 (N_16573,N_13216,N_14902);
and U16574 (N_16574,N_12931,N_13525);
or U16575 (N_16575,N_13801,N_13674);
nand U16576 (N_16576,N_14414,N_13581);
nor U16577 (N_16577,N_14158,N_14775);
xnor U16578 (N_16578,N_13623,N_14335);
xnor U16579 (N_16579,N_14402,N_14048);
nor U16580 (N_16580,N_14109,N_14252);
xnor U16581 (N_16581,N_12530,N_14994);
nand U16582 (N_16582,N_13043,N_14318);
or U16583 (N_16583,N_13853,N_12796);
nor U16584 (N_16584,N_13293,N_13530);
and U16585 (N_16585,N_12964,N_12873);
and U16586 (N_16586,N_13072,N_14380);
nand U16587 (N_16587,N_14690,N_14502);
nor U16588 (N_16588,N_14862,N_14926);
xnor U16589 (N_16589,N_12952,N_13352);
nand U16590 (N_16590,N_13399,N_13203);
nor U16591 (N_16591,N_13268,N_13618);
or U16592 (N_16592,N_13141,N_12907);
nand U16593 (N_16593,N_13666,N_13210);
xor U16594 (N_16594,N_14962,N_14541);
nand U16595 (N_16595,N_12614,N_13941);
nor U16596 (N_16596,N_13586,N_13959);
and U16597 (N_16597,N_13790,N_14333);
nor U16598 (N_16598,N_14024,N_14469);
and U16599 (N_16599,N_12671,N_12575);
or U16600 (N_16600,N_12747,N_12743);
xor U16601 (N_16601,N_14084,N_13331);
nor U16602 (N_16602,N_14481,N_14528);
or U16603 (N_16603,N_12860,N_14570);
nand U16604 (N_16604,N_14558,N_13065);
xor U16605 (N_16605,N_13241,N_12979);
nor U16606 (N_16606,N_12842,N_14884);
nor U16607 (N_16607,N_14351,N_13525);
xnor U16608 (N_16608,N_13674,N_13046);
nand U16609 (N_16609,N_13709,N_14399);
nor U16610 (N_16610,N_12664,N_13466);
nor U16611 (N_16611,N_14566,N_13421);
and U16612 (N_16612,N_14331,N_14288);
nand U16613 (N_16613,N_14188,N_13191);
and U16614 (N_16614,N_13445,N_12676);
xor U16615 (N_16615,N_14695,N_14458);
nor U16616 (N_16616,N_12717,N_14809);
or U16617 (N_16617,N_12813,N_13014);
nor U16618 (N_16618,N_14557,N_14318);
or U16619 (N_16619,N_12776,N_14933);
and U16620 (N_16620,N_13589,N_12910);
xnor U16621 (N_16621,N_13039,N_13827);
and U16622 (N_16622,N_13816,N_13849);
xnor U16623 (N_16623,N_12674,N_13760);
nor U16624 (N_16624,N_13044,N_14533);
and U16625 (N_16625,N_13739,N_13493);
and U16626 (N_16626,N_14974,N_13971);
and U16627 (N_16627,N_14722,N_12788);
nand U16628 (N_16628,N_13759,N_13515);
or U16629 (N_16629,N_13546,N_13936);
or U16630 (N_16630,N_13393,N_13134);
xor U16631 (N_16631,N_13010,N_13424);
nor U16632 (N_16632,N_13808,N_12905);
nand U16633 (N_16633,N_12532,N_13563);
and U16634 (N_16634,N_14448,N_14498);
or U16635 (N_16635,N_14968,N_14631);
and U16636 (N_16636,N_14992,N_14379);
xor U16637 (N_16637,N_12881,N_14030);
xnor U16638 (N_16638,N_13410,N_13919);
nor U16639 (N_16639,N_13577,N_13110);
nor U16640 (N_16640,N_13548,N_13653);
nand U16641 (N_16641,N_12971,N_14110);
nand U16642 (N_16642,N_14602,N_14487);
and U16643 (N_16643,N_12750,N_13377);
xnor U16644 (N_16644,N_13435,N_13544);
or U16645 (N_16645,N_14913,N_14655);
and U16646 (N_16646,N_14452,N_14346);
and U16647 (N_16647,N_13875,N_14826);
nand U16648 (N_16648,N_13041,N_12936);
nand U16649 (N_16649,N_14108,N_14992);
nand U16650 (N_16650,N_13835,N_14483);
nor U16651 (N_16651,N_13019,N_13190);
nand U16652 (N_16652,N_13560,N_13827);
xnor U16653 (N_16653,N_13555,N_12553);
or U16654 (N_16654,N_13591,N_14631);
nor U16655 (N_16655,N_14361,N_12858);
and U16656 (N_16656,N_14075,N_14638);
nand U16657 (N_16657,N_13108,N_14055);
nand U16658 (N_16658,N_14361,N_13018);
nand U16659 (N_16659,N_13260,N_14908);
xnor U16660 (N_16660,N_14358,N_14588);
nor U16661 (N_16661,N_14078,N_13284);
nor U16662 (N_16662,N_13851,N_14826);
and U16663 (N_16663,N_13664,N_13269);
nor U16664 (N_16664,N_13917,N_13407);
and U16665 (N_16665,N_13221,N_14280);
or U16666 (N_16666,N_13696,N_14695);
nor U16667 (N_16667,N_13736,N_13851);
xnor U16668 (N_16668,N_14573,N_13362);
and U16669 (N_16669,N_13112,N_13347);
xnor U16670 (N_16670,N_13640,N_14058);
or U16671 (N_16671,N_14419,N_14325);
nand U16672 (N_16672,N_14092,N_12957);
and U16673 (N_16673,N_14177,N_13286);
xnor U16674 (N_16674,N_12609,N_12844);
or U16675 (N_16675,N_14796,N_14340);
nand U16676 (N_16676,N_12550,N_14231);
or U16677 (N_16677,N_14153,N_14579);
and U16678 (N_16678,N_14552,N_12999);
xnor U16679 (N_16679,N_14534,N_12573);
xnor U16680 (N_16680,N_14865,N_14912);
and U16681 (N_16681,N_13025,N_14363);
and U16682 (N_16682,N_13385,N_14521);
or U16683 (N_16683,N_14870,N_13538);
xor U16684 (N_16684,N_13623,N_13353);
nand U16685 (N_16685,N_12546,N_12719);
xor U16686 (N_16686,N_12853,N_12502);
and U16687 (N_16687,N_14517,N_12724);
xor U16688 (N_16688,N_14002,N_14944);
nand U16689 (N_16689,N_12962,N_14917);
xnor U16690 (N_16690,N_12989,N_14405);
nor U16691 (N_16691,N_13679,N_14980);
and U16692 (N_16692,N_13608,N_13506);
or U16693 (N_16693,N_14698,N_13251);
or U16694 (N_16694,N_14164,N_13055);
and U16695 (N_16695,N_13957,N_12933);
nor U16696 (N_16696,N_13065,N_12803);
nor U16697 (N_16697,N_12720,N_14916);
xor U16698 (N_16698,N_13777,N_13332);
and U16699 (N_16699,N_14337,N_13307);
nor U16700 (N_16700,N_12638,N_12629);
or U16701 (N_16701,N_13116,N_13550);
nor U16702 (N_16702,N_13700,N_14501);
xnor U16703 (N_16703,N_14075,N_14956);
and U16704 (N_16704,N_13162,N_13072);
nand U16705 (N_16705,N_12660,N_13779);
and U16706 (N_16706,N_13695,N_12935);
or U16707 (N_16707,N_12962,N_13182);
and U16708 (N_16708,N_13706,N_14570);
or U16709 (N_16709,N_14603,N_13999);
or U16710 (N_16710,N_13449,N_13398);
or U16711 (N_16711,N_12868,N_14659);
or U16712 (N_16712,N_13900,N_14814);
or U16713 (N_16713,N_13255,N_13539);
nand U16714 (N_16714,N_12863,N_14699);
and U16715 (N_16715,N_13082,N_13013);
nand U16716 (N_16716,N_14066,N_12504);
xnor U16717 (N_16717,N_12504,N_14722);
nor U16718 (N_16718,N_13828,N_13293);
and U16719 (N_16719,N_12754,N_14941);
nor U16720 (N_16720,N_12647,N_14321);
xnor U16721 (N_16721,N_12605,N_12563);
nor U16722 (N_16722,N_12606,N_13133);
xor U16723 (N_16723,N_14979,N_13615);
nor U16724 (N_16724,N_13702,N_12980);
xor U16725 (N_16725,N_13956,N_12914);
xnor U16726 (N_16726,N_13430,N_14742);
or U16727 (N_16727,N_13252,N_13262);
nand U16728 (N_16728,N_12809,N_12947);
nand U16729 (N_16729,N_14050,N_13501);
or U16730 (N_16730,N_13195,N_14372);
and U16731 (N_16731,N_13332,N_14729);
or U16732 (N_16732,N_12907,N_13615);
nand U16733 (N_16733,N_14243,N_12603);
nor U16734 (N_16734,N_13613,N_14026);
or U16735 (N_16735,N_12621,N_14191);
or U16736 (N_16736,N_13581,N_14610);
and U16737 (N_16737,N_13149,N_13656);
nand U16738 (N_16738,N_14093,N_12709);
xnor U16739 (N_16739,N_13857,N_14858);
and U16740 (N_16740,N_14111,N_13847);
and U16741 (N_16741,N_13965,N_14481);
xnor U16742 (N_16742,N_14083,N_13687);
and U16743 (N_16743,N_12785,N_12928);
xor U16744 (N_16744,N_13190,N_14234);
and U16745 (N_16745,N_12753,N_13929);
nand U16746 (N_16746,N_13786,N_13674);
and U16747 (N_16747,N_13713,N_14680);
nor U16748 (N_16748,N_13592,N_12896);
xor U16749 (N_16749,N_12625,N_14397);
and U16750 (N_16750,N_14790,N_13353);
or U16751 (N_16751,N_13641,N_14448);
xnor U16752 (N_16752,N_13332,N_14717);
nor U16753 (N_16753,N_13045,N_14174);
nand U16754 (N_16754,N_12603,N_12896);
nand U16755 (N_16755,N_12914,N_14673);
nand U16756 (N_16756,N_12937,N_14353);
xnor U16757 (N_16757,N_14337,N_13209);
and U16758 (N_16758,N_13950,N_13058);
xnor U16759 (N_16759,N_14513,N_13434);
xor U16760 (N_16760,N_13136,N_13141);
or U16761 (N_16761,N_12655,N_13019);
or U16762 (N_16762,N_14976,N_12646);
xnor U16763 (N_16763,N_13708,N_14496);
and U16764 (N_16764,N_13964,N_14294);
xor U16765 (N_16765,N_12576,N_12850);
nor U16766 (N_16766,N_13008,N_14541);
nor U16767 (N_16767,N_14715,N_12756);
xnor U16768 (N_16768,N_14612,N_13223);
nor U16769 (N_16769,N_12859,N_12514);
nor U16770 (N_16770,N_12891,N_14086);
xnor U16771 (N_16771,N_12912,N_12833);
nand U16772 (N_16772,N_13933,N_13392);
or U16773 (N_16773,N_13995,N_12744);
xor U16774 (N_16774,N_14957,N_13988);
or U16775 (N_16775,N_14250,N_13805);
xor U16776 (N_16776,N_13360,N_12841);
xnor U16777 (N_16777,N_13833,N_14758);
xor U16778 (N_16778,N_13928,N_12975);
nor U16779 (N_16779,N_12618,N_12774);
and U16780 (N_16780,N_14849,N_14878);
nand U16781 (N_16781,N_14951,N_13550);
nand U16782 (N_16782,N_14994,N_12848);
and U16783 (N_16783,N_14536,N_14732);
nand U16784 (N_16784,N_12810,N_14405);
or U16785 (N_16785,N_13820,N_13619);
xor U16786 (N_16786,N_13825,N_14047);
nor U16787 (N_16787,N_14451,N_14046);
and U16788 (N_16788,N_13738,N_14934);
or U16789 (N_16789,N_14778,N_14423);
xor U16790 (N_16790,N_14536,N_14349);
nand U16791 (N_16791,N_14206,N_13679);
nand U16792 (N_16792,N_14935,N_13403);
nor U16793 (N_16793,N_12879,N_13491);
xor U16794 (N_16794,N_14864,N_12759);
nand U16795 (N_16795,N_14831,N_14893);
or U16796 (N_16796,N_13287,N_12518);
xnor U16797 (N_16797,N_14923,N_14918);
xor U16798 (N_16798,N_14949,N_12856);
or U16799 (N_16799,N_12671,N_13100);
or U16800 (N_16800,N_13563,N_14790);
and U16801 (N_16801,N_12614,N_13841);
nand U16802 (N_16802,N_12747,N_13312);
nand U16803 (N_16803,N_13919,N_14046);
or U16804 (N_16804,N_13619,N_13325);
nor U16805 (N_16805,N_14302,N_14487);
nand U16806 (N_16806,N_14812,N_14021);
or U16807 (N_16807,N_12548,N_14643);
nand U16808 (N_16808,N_14142,N_14390);
and U16809 (N_16809,N_14983,N_14254);
or U16810 (N_16810,N_13255,N_14207);
xor U16811 (N_16811,N_13042,N_14347);
and U16812 (N_16812,N_12677,N_12987);
and U16813 (N_16813,N_14163,N_14475);
nor U16814 (N_16814,N_12613,N_14323);
nand U16815 (N_16815,N_13583,N_14039);
nor U16816 (N_16816,N_14651,N_14841);
nor U16817 (N_16817,N_14371,N_12502);
or U16818 (N_16818,N_14421,N_14025);
nor U16819 (N_16819,N_14587,N_12628);
xor U16820 (N_16820,N_14585,N_13948);
nor U16821 (N_16821,N_13280,N_13329);
nand U16822 (N_16822,N_12611,N_14757);
nand U16823 (N_16823,N_12908,N_12648);
xor U16824 (N_16824,N_13215,N_13709);
nand U16825 (N_16825,N_14651,N_12594);
or U16826 (N_16826,N_13952,N_13906);
or U16827 (N_16827,N_14977,N_13811);
nor U16828 (N_16828,N_14999,N_14460);
xor U16829 (N_16829,N_13810,N_13576);
or U16830 (N_16830,N_14012,N_13518);
nor U16831 (N_16831,N_12958,N_14249);
or U16832 (N_16832,N_13390,N_14225);
and U16833 (N_16833,N_14964,N_14354);
or U16834 (N_16834,N_14074,N_13702);
xnor U16835 (N_16835,N_13714,N_12923);
or U16836 (N_16836,N_13142,N_12918);
xor U16837 (N_16837,N_14510,N_13583);
nor U16838 (N_16838,N_13213,N_13736);
xor U16839 (N_16839,N_13395,N_14270);
or U16840 (N_16840,N_12915,N_12612);
or U16841 (N_16841,N_14873,N_14452);
and U16842 (N_16842,N_14047,N_14999);
xnor U16843 (N_16843,N_13978,N_13047);
or U16844 (N_16844,N_12966,N_14318);
and U16845 (N_16845,N_14146,N_12689);
and U16846 (N_16846,N_13165,N_14004);
xor U16847 (N_16847,N_12666,N_12888);
nor U16848 (N_16848,N_14404,N_12604);
nand U16849 (N_16849,N_13606,N_12953);
nand U16850 (N_16850,N_13150,N_14294);
or U16851 (N_16851,N_13001,N_14777);
or U16852 (N_16852,N_14572,N_14496);
nor U16853 (N_16853,N_13472,N_13747);
and U16854 (N_16854,N_14798,N_12984);
nand U16855 (N_16855,N_13056,N_13621);
and U16856 (N_16856,N_13329,N_13653);
nor U16857 (N_16857,N_13287,N_13611);
nand U16858 (N_16858,N_14872,N_14077);
and U16859 (N_16859,N_13316,N_13690);
nor U16860 (N_16860,N_12502,N_14430);
nor U16861 (N_16861,N_13341,N_13781);
xnor U16862 (N_16862,N_14815,N_13898);
nand U16863 (N_16863,N_14150,N_13709);
nand U16864 (N_16864,N_13625,N_12914);
nor U16865 (N_16865,N_14604,N_14981);
xnor U16866 (N_16866,N_12945,N_12923);
or U16867 (N_16867,N_14254,N_12717);
nor U16868 (N_16868,N_14420,N_13733);
xnor U16869 (N_16869,N_14490,N_14804);
nor U16870 (N_16870,N_13879,N_13538);
nor U16871 (N_16871,N_13110,N_13736);
and U16872 (N_16872,N_14923,N_14010);
nand U16873 (N_16873,N_13222,N_13924);
and U16874 (N_16874,N_13489,N_14246);
xnor U16875 (N_16875,N_14052,N_14500);
or U16876 (N_16876,N_14993,N_14361);
nand U16877 (N_16877,N_12726,N_13869);
nand U16878 (N_16878,N_13307,N_14651);
and U16879 (N_16879,N_12845,N_13079);
or U16880 (N_16880,N_14963,N_13158);
and U16881 (N_16881,N_14057,N_13745);
nor U16882 (N_16882,N_14360,N_13489);
and U16883 (N_16883,N_14849,N_14626);
nand U16884 (N_16884,N_14150,N_13695);
nor U16885 (N_16885,N_13028,N_13664);
xnor U16886 (N_16886,N_14095,N_12559);
xnor U16887 (N_16887,N_14985,N_13478);
nor U16888 (N_16888,N_14742,N_14326);
nor U16889 (N_16889,N_13001,N_13017);
or U16890 (N_16890,N_13660,N_14024);
nand U16891 (N_16891,N_14180,N_13325);
nand U16892 (N_16892,N_14786,N_14113);
and U16893 (N_16893,N_14370,N_13145);
or U16894 (N_16894,N_14085,N_13693);
nor U16895 (N_16895,N_13143,N_14507);
and U16896 (N_16896,N_13502,N_14159);
or U16897 (N_16897,N_14024,N_14332);
nand U16898 (N_16898,N_12902,N_13704);
xnor U16899 (N_16899,N_13232,N_13634);
and U16900 (N_16900,N_13227,N_14083);
xnor U16901 (N_16901,N_13248,N_14231);
xor U16902 (N_16902,N_13065,N_13434);
and U16903 (N_16903,N_14241,N_14136);
or U16904 (N_16904,N_14176,N_13057);
nand U16905 (N_16905,N_12837,N_13021);
xor U16906 (N_16906,N_14498,N_13456);
xor U16907 (N_16907,N_13079,N_12755);
nand U16908 (N_16908,N_13952,N_14810);
and U16909 (N_16909,N_12745,N_13925);
xnor U16910 (N_16910,N_12789,N_12939);
and U16911 (N_16911,N_13268,N_14717);
nor U16912 (N_16912,N_14867,N_14498);
nor U16913 (N_16913,N_13207,N_13310);
and U16914 (N_16914,N_14383,N_13630);
xnor U16915 (N_16915,N_14000,N_14975);
nand U16916 (N_16916,N_12761,N_12904);
or U16917 (N_16917,N_14942,N_13612);
nand U16918 (N_16918,N_13575,N_13663);
or U16919 (N_16919,N_14825,N_13005);
or U16920 (N_16920,N_13335,N_13118);
xnor U16921 (N_16921,N_14455,N_13932);
nor U16922 (N_16922,N_12531,N_14058);
and U16923 (N_16923,N_13813,N_12709);
nor U16924 (N_16924,N_12518,N_14997);
xnor U16925 (N_16925,N_14878,N_13853);
and U16926 (N_16926,N_13278,N_12741);
xnor U16927 (N_16927,N_13434,N_14247);
nor U16928 (N_16928,N_13099,N_14280);
xnor U16929 (N_16929,N_14214,N_13459);
xor U16930 (N_16930,N_13335,N_13695);
nand U16931 (N_16931,N_13451,N_13850);
nor U16932 (N_16932,N_14096,N_13077);
and U16933 (N_16933,N_13373,N_14784);
or U16934 (N_16934,N_12849,N_14695);
or U16935 (N_16935,N_13390,N_12997);
xnor U16936 (N_16936,N_13669,N_14619);
xnor U16937 (N_16937,N_14025,N_14513);
xor U16938 (N_16938,N_12500,N_14893);
and U16939 (N_16939,N_14786,N_14386);
nand U16940 (N_16940,N_13331,N_14032);
nand U16941 (N_16941,N_14123,N_13792);
xnor U16942 (N_16942,N_14811,N_14320);
xnor U16943 (N_16943,N_14656,N_13762);
and U16944 (N_16944,N_13303,N_12695);
and U16945 (N_16945,N_13127,N_13634);
nor U16946 (N_16946,N_13414,N_12995);
nor U16947 (N_16947,N_14909,N_14466);
and U16948 (N_16948,N_13929,N_12818);
xor U16949 (N_16949,N_13745,N_13540);
nor U16950 (N_16950,N_13094,N_14326);
xnor U16951 (N_16951,N_14384,N_12561);
and U16952 (N_16952,N_13155,N_13169);
and U16953 (N_16953,N_14745,N_12630);
and U16954 (N_16954,N_12664,N_13220);
nand U16955 (N_16955,N_14492,N_13445);
nor U16956 (N_16956,N_12919,N_14461);
or U16957 (N_16957,N_13286,N_14882);
nand U16958 (N_16958,N_12509,N_14161);
nor U16959 (N_16959,N_13426,N_12756);
and U16960 (N_16960,N_14884,N_14976);
and U16961 (N_16961,N_14684,N_13776);
nor U16962 (N_16962,N_14720,N_13439);
xor U16963 (N_16963,N_14345,N_13186);
and U16964 (N_16964,N_12674,N_14202);
nand U16965 (N_16965,N_12670,N_14609);
nand U16966 (N_16966,N_13371,N_12842);
nand U16967 (N_16967,N_13982,N_12592);
nor U16968 (N_16968,N_13514,N_14838);
nand U16969 (N_16969,N_13208,N_13466);
nand U16970 (N_16970,N_12992,N_14190);
and U16971 (N_16971,N_13487,N_13572);
nor U16972 (N_16972,N_13274,N_13677);
and U16973 (N_16973,N_14793,N_14556);
nand U16974 (N_16974,N_13074,N_14573);
or U16975 (N_16975,N_13184,N_14853);
nor U16976 (N_16976,N_13705,N_14130);
or U16977 (N_16977,N_14109,N_14236);
xor U16978 (N_16978,N_14554,N_14095);
and U16979 (N_16979,N_12750,N_14907);
or U16980 (N_16980,N_14062,N_14102);
nand U16981 (N_16981,N_12629,N_12869);
and U16982 (N_16982,N_14464,N_12683);
nand U16983 (N_16983,N_13747,N_12743);
nand U16984 (N_16984,N_14788,N_13004);
and U16985 (N_16985,N_12951,N_14483);
nand U16986 (N_16986,N_14112,N_14944);
and U16987 (N_16987,N_12684,N_14873);
or U16988 (N_16988,N_14335,N_14183);
nor U16989 (N_16989,N_12796,N_14169);
xor U16990 (N_16990,N_13323,N_14549);
or U16991 (N_16991,N_13432,N_12845);
nor U16992 (N_16992,N_14839,N_14901);
xnor U16993 (N_16993,N_14860,N_13503);
nor U16994 (N_16994,N_14204,N_14144);
nor U16995 (N_16995,N_13427,N_13158);
nor U16996 (N_16996,N_12645,N_14442);
xor U16997 (N_16997,N_13805,N_12950);
xnor U16998 (N_16998,N_14179,N_12889);
or U16999 (N_16999,N_12544,N_14586);
and U17000 (N_17000,N_13421,N_12864);
xnor U17001 (N_17001,N_13437,N_14809);
nor U17002 (N_17002,N_14722,N_14630);
and U17003 (N_17003,N_14730,N_13455);
nand U17004 (N_17004,N_14221,N_13689);
xnor U17005 (N_17005,N_12648,N_14907);
or U17006 (N_17006,N_14518,N_13885);
or U17007 (N_17007,N_14980,N_14442);
nand U17008 (N_17008,N_13482,N_12789);
nor U17009 (N_17009,N_14026,N_14138);
and U17010 (N_17010,N_14766,N_14560);
nand U17011 (N_17011,N_13133,N_14884);
nor U17012 (N_17012,N_14519,N_14959);
or U17013 (N_17013,N_13402,N_13472);
and U17014 (N_17014,N_14756,N_12940);
and U17015 (N_17015,N_13350,N_13562);
and U17016 (N_17016,N_12854,N_13601);
nor U17017 (N_17017,N_12561,N_14173);
or U17018 (N_17018,N_14986,N_12981);
or U17019 (N_17019,N_13719,N_13975);
and U17020 (N_17020,N_12867,N_14692);
nand U17021 (N_17021,N_14353,N_14418);
and U17022 (N_17022,N_12875,N_12513);
nand U17023 (N_17023,N_14069,N_13968);
nand U17024 (N_17024,N_13434,N_12852);
nand U17025 (N_17025,N_14069,N_13913);
and U17026 (N_17026,N_14174,N_12888);
nand U17027 (N_17027,N_14377,N_14807);
or U17028 (N_17028,N_13609,N_13097);
nor U17029 (N_17029,N_13253,N_12888);
nor U17030 (N_17030,N_13679,N_13542);
nand U17031 (N_17031,N_14722,N_13689);
and U17032 (N_17032,N_14686,N_12536);
nor U17033 (N_17033,N_12683,N_14905);
or U17034 (N_17034,N_14228,N_13780);
or U17035 (N_17035,N_12659,N_12963);
or U17036 (N_17036,N_14873,N_14343);
nand U17037 (N_17037,N_13348,N_13649);
nor U17038 (N_17038,N_14997,N_13356);
and U17039 (N_17039,N_13879,N_12883);
nand U17040 (N_17040,N_14448,N_14449);
nor U17041 (N_17041,N_14127,N_14130);
nand U17042 (N_17042,N_13427,N_13924);
xnor U17043 (N_17043,N_13765,N_12650);
and U17044 (N_17044,N_13799,N_13964);
nor U17045 (N_17045,N_13918,N_13044);
and U17046 (N_17046,N_14384,N_13542);
nor U17047 (N_17047,N_12797,N_14154);
nand U17048 (N_17048,N_14405,N_12697);
nand U17049 (N_17049,N_14875,N_13870);
and U17050 (N_17050,N_14504,N_14759);
nor U17051 (N_17051,N_12785,N_14406);
nor U17052 (N_17052,N_13729,N_12505);
nand U17053 (N_17053,N_14533,N_13722);
or U17054 (N_17054,N_14988,N_12836);
or U17055 (N_17055,N_14639,N_13044);
and U17056 (N_17056,N_13627,N_12702);
and U17057 (N_17057,N_13936,N_13659);
nand U17058 (N_17058,N_12567,N_12685);
xor U17059 (N_17059,N_13097,N_14909);
nand U17060 (N_17060,N_13496,N_14746);
nor U17061 (N_17061,N_14755,N_14908);
and U17062 (N_17062,N_14612,N_13831);
or U17063 (N_17063,N_13918,N_12627);
xnor U17064 (N_17064,N_12721,N_13924);
or U17065 (N_17065,N_14731,N_12840);
nor U17066 (N_17066,N_14506,N_13177);
nor U17067 (N_17067,N_13399,N_13110);
xnor U17068 (N_17068,N_13405,N_13721);
and U17069 (N_17069,N_14763,N_12928);
and U17070 (N_17070,N_12750,N_12748);
or U17071 (N_17071,N_13697,N_12547);
xor U17072 (N_17072,N_13171,N_12857);
xor U17073 (N_17073,N_14741,N_14523);
xnor U17074 (N_17074,N_13848,N_12985);
xor U17075 (N_17075,N_13455,N_14838);
nand U17076 (N_17076,N_12582,N_13517);
or U17077 (N_17077,N_14754,N_14775);
nand U17078 (N_17078,N_14103,N_13979);
nor U17079 (N_17079,N_13070,N_13683);
nand U17080 (N_17080,N_14813,N_12808);
and U17081 (N_17081,N_14529,N_13333);
nor U17082 (N_17082,N_13082,N_14548);
xnor U17083 (N_17083,N_12512,N_14878);
nand U17084 (N_17084,N_13105,N_13433);
and U17085 (N_17085,N_13750,N_13212);
and U17086 (N_17086,N_14217,N_14860);
and U17087 (N_17087,N_13514,N_13492);
and U17088 (N_17088,N_13738,N_13676);
xor U17089 (N_17089,N_14342,N_14560);
and U17090 (N_17090,N_14239,N_13652);
nor U17091 (N_17091,N_14108,N_12685);
or U17092 (N_17092,N_14823,N_14862);
or U17093 (N_17093,N_13751,N_13328);
and U17094 (N_17094,N_14406,N_14794);
nand U17095 (N_17095,N_14442,N_14527);
nor U17096 (N_17096,N_14689,N_13304);
xor U17097 (N_17097,N_14710,N_14805);
or U17098 (N_17098,N_13276,N_14163);
nand U17099 (N_17099,N_12651,N_14130);
and U17100 (N_17100,N_14782,N_14665);
or U17101 (N_17101,N_12908,N_13640);
xnor U17102 (N_17102,N_13564,N_14865);
nor U17103 (N_17103,N_14845,N_13676);
xor U17104 (N_17104,N_14562,N_13283);
nor U17105 (N_17105,N_13452,N_14027);
nand U17106 (N_17106,N_13284,N_12773);
or U17107 (N_17107,N_12834,N_14250);
xnor U17108 (N_17108,N_14270,N_12618);
nand U17109 (N_17109,N_12941,N_14192);
and U17110 (N_17110,N_13361,N_14062);
or U17111 (N_17111,N_14253,N_14767);
nand U17112 (N_17112,N_14124,N_14711);
or U17113 (N_17113,N_12641,N_14550);
and U17114 (N_17114,N_14099,N_13582);
nand U17115 (N_17115,N_12686,N_13286);
and U17116 (N_17116,N_13524,N_12677);
nand U17117 (N_17117,N_13914,N_14880);
and U17118 (N_17118,N_14972,N_14008);
nand U17119 (N_17119,N_13515,N_14799);
nor U17120 (N_17120,N_12645,N_12616);
and U17121 (N_17121,N_12840,N_13379);
nand U17122 (N_17122,N_12922,N_12789);
nor U17123 (N_17123,N_14255,N_12879);
nor U17124 (N_17124,N_13858,N_13568);
xor U17125 (N_17125,N_13429,N_14669);
nand U17126 (N_17126,N_13581,N_13163);
or U17127 (N_17127,N_14311,N_13858);
xor U17128 (N_17128,N_12912,N_13240);
nand U17129 (N_17129,N_13720,N_13697);
or U17130 (N_17130,N_14387,N_14783);
nor U17131 (N_17131,N_13338,N_14535);
nor U17132 (N_17132,N_13045,N_13976);
nand U17133 (N_17133,N_14555,N_12615);
nand U17134 (N_17134,N_14065,N_12741);
nor U17135 (N_17135,N_12599,N_13460);
and U17136 (N_17136,N_13472,N_12899);
nor U17137 (N_17137,N_13296,N_12588);
xor U17138 (N_17138,N_13725,N_14438);
or U17139 (N_17139,N_13321,N_12860);
xnor U17140 (N_17140,N_14778,N_13009);
nor U17141 (N_17141,N_13243,N_13285);
or U17142 (N_17142,N_14524,N_13052);
and U17143 (N_17143,N_13709,N_13856);
nor U17144 (N_17144,N_12754,N_14783);
or U17145 (N_17145,N_14836,N_14055);
xnor U17146 (N_17146,N_14299,N_13961);
and U17147 (N_17147,N_12850,N_13566);
nand U17148 (N_17148,N_13613,N_14488);
and U17149 (N_17149,N_13098,N_12769);
and U17150 (N_17150,N_14441,N_14120);
nand U17151 (N_17151,N_14487,N_13138);
nor U17152 (N_17152,N_14314,N_14978);
nand U17153 (N_17153,N_13599,N_14240);
and U17154 (N_17154,N_12585,N_13623);
nor U17155 (N_17155,N_14003,N_14784);
xor U17156 (N_17156,N_13812,N_12621);
nand U17157 (N_17157,N_14118,N_13418);
nand U17158 (N_17158,N_12515,N_13325);
nor U17159 (N_17159,N_12559,N_13474);
and U17160 (N_17160,N_14819,N_14091);
nand U17161 (N_17161,N_14863,N_12771);
or U17162 (N_17162,N_13272,N_14824);
nand U17163 (N_17163,N_13210,N_14135);
nand U17164 (N_17164,N_14631,N_13230);
xnor U17165 (N_17165,N_13659,N_13491);
and U17166 (N_17166,N_13990,N_14942);
nand U17167 (N_17167,N_14362,N_14849);
or U17168 (N_17168,N_13637,N_12816);
xnor U17169 (N_17169,N_13113,N_14460);
nand U17170 (N_17170,N_14385,N_13011);
and U17171 (N_17171,N_13814,N_13146);
or U17172 (N_17172,N_13643,N_13024);
and U17173 (N_17173,N_12689,N_12912);
xor U17174 (N_17174,N_13114,N_13390);
xnor U17175 (N_17175,N_14711,N_14350);
xor U17176 (N_17176,N_14439,N_13297);
nor U17177 (N_17177,N_14939,N_12589);
or U17178 (N_17178,N_12777,N_14895);
xor U17179 (N_17179,N_12735,N_14919);
or U17180 (N_17180,N_14262,N_13918);
xor U17181 (N_17181,N_14179,N_12570);
and U17182 (N_17182,N_14706,N_13973);
nor U17183 (N_17183,N_12581,N_13346);
nand U17184 (N_17184,N_14890,N_12929);
nand U17185 (N_17185,N_12525,N_13724);
nor U17186 (N_17186,N_13930,N_13779);
nand U17187 (N_17187,N_14907,N_13585);
and U17188 (N_17188,N_14651,N_14276);
or U17189 (N_17189,N_14412,N_14407);
and U17190 (N_17190,N_14525,N_14365);
xor U17191 (N_17191,N_13686,N_12946);
nor U17192 (N_17192,N_13826,N_14569);
and U17193 (N_17193,N_13721,N_13537);
and U17194 (N_17194,N_14363,N_13937);
and U17195 (N_17195,N_14350,N_13647);
xnor U17196 (N_17196,N_13476,N_13794);
or U17197 (N_17197,N_13592,N_12545);
xnor U17198 (N_17198,N_13267,N_13725);
xor U17199 (N_17199,N_12684,N_13953);
or U17200 (N_17200,N_13519,N_12591);
nor U17201 (N_17201,N_12691,N_13075);
or U17202 (N_17202,N_14853,N_12693);
and U17203 (N_17203,N_14580,N_13152);
nor U17204 (N_17204,N_12951,N_14981);
nor U17205 (N_17205,N_13414,N_14755);
xnor U17206 (N_17206,N_13032,N_14314);
and U17207 (N_17207,N_13333,N_12597);
xnor U17208 (N_17208,N_12574,N_12532);
xor U17209 (N_17209,N_14371,N_13225);
nand U17210 (N_17210,N_13021,N_14515);
nor U17211 (N_17211,N_12699,N_13083);
nand U17212 (N_17212,N_13725,N_14770);
or U17213 (N_17213,N_13069,N_13821);
and U17214 (N_17214,N_13100,N_13529);
or U17215 (N_17215,N_13750,N_13724);
nand U17216 (N_17216,N_14959,N_14832);
xnor U17217 (N_17217,N_12776,N_14971);
nand U17218 (N_17218,N_12986,N_14294);
nand U17219 (N_17219,N_14205,N_14688);
nand U17220 (N_17220,N_13302,N_14391);
nand U17221 (N_17221,N_14885,N_13391);
and U17222 (N_17222,N_13404,N_14708);
xnor U17223 (N_17223,N_12982,N_12770);
or U17224 (N_17224,N_12600,N_14044);
nand U17225 (N_17225,N_13548,N_14377);
nand U17226 (N_17226,N_12595,N_13227);
nor U17227 (N_17227,N_13301,N_13194);
or U17228 (N_17228,N_13987,N_13323);
nand U17229 (N_17229,N_13950,N_14277);
xor U17230 (N_17230,N_14726,N_14182);
xnor U17231 (N_17231,N_14270,N_13183);
and U17232 (N_17232,N_12880,N_13892);
and U17233 (N_17233,N_13720,N_12833);
and U17234 (N_17234,N_13808,N_13716);
xor U17235 (N_17235,N_12604,N_12981);
or U17236 (N_17236,N_14724,N_14771);
nor U17237 (N_17237,N_14882,N_13456);
and U17238 (N_17238,N_12925,N_13750);
or U17239 (N_17239,N_14531,N_13430);
or U17240 (N_17240,N_14767,N_14993);
nor U17241 (N_17241,N_14509,N_14324);
nand U17242 (N_17242,N_12879,N_14474);
or U17243 (N_17243,N_13313,N_13320);
and U17244 (N_17244,N_13930,N_14375);
xnor U17245 (N_17245,N_13020,N_13391);
or U17246 (N_17246,N_14422,N_13565);
nor U17247 (N_17247,N_13106,N_13663);
nor U17248 (N_17248,N_12683,N_12665);
xor U17249 (N_17249,N_14858,N_14819);
and U17250 (N_17250,N_14509,N_14304);
nor U17251 (N_17251,N_14401,N_13057);
nor U17252 (N_17252,N_14218,N_12789);
nand U17253 (N_17253,N_13746,N_12911);
and U17254 (N_17254,N_13368,N_13765);
xnor U17255 (N_17255,N_12681,N_14626);
nand U17256 (N_17256,N_13882,N_13848);
or U17257 (N_17257,N_14957,N_14408);
xor U17258 (N_17258,N_14875,N_13661);
and U17259 (N_17259,N_14944,N_13155);
xor U17260 (N_17260,N_13848,N_14579);
xor U17261 (N_17261,N_13672,N_14057);
and U17262 (N_17262,N_13335,N_12734);
or U17263 (N_17263,N_14619,N_12756);
and U17264 (N_17264,N_12846,N_13827);
xnor U17265 (N_17265,N_13248,N_13626);
nand U17266 (N_17266,N_13609,N_14829);
nand U17267 (N_17267,N_13635,N_14068);
nor U17268 (N_17268,N_12547,N_14658);
nor U17269 (N_17269,N_13633,N_13274);
or U17270 (N_17270,N_14784,N_14655);
nor U17271 (N_17271,N_13537,N_12918);
xnor U17272 (N_17272,N_13986,N_14422);
xnor U17273 (N_17273,N_12821,N_13991);
xor U17274 (N_17274,N_14416,N_13928);
or U17275 (N_17275,N_14460,N_13682);
xnor U17276 (N_17276,N_14615,N_14700);
nand U17277 (N_17277,N_12738,N_14767);
xnor U17278 (N_17278,N_13131,N_12706);
nand U17279 (N_17279,N_13574,N_13269);
nor U17280 (N_17280,N_13044,N_12987);
nor U17281 (N_17281,N_14718,N_12827);
nand U17282 (N_17282,N_12579,N_12854);
and U17283 (N_17283,N_12821,N_14088);
nand U17284 (N_17284,N_13206,N_13122);
nand U17285 (N_17285,N_14703,N_12812);
xnor U17286 (N_17286,N_14141,N_14394);
nand U17287 (N_17287,N_14294,N_13461);
nand U17288 (N_17288,N_13679,N_13636);
nor U17289 (N_17289,N_13418,N_13535);
or U17290 (N_17290,N_13103,N_13153);
or U17291 (N_17291,N_14690,N_14246);
or U17292 (N_17292,N_12948,N_13030);
xor U17293 (N_17293,N_13348,N_14873);
or U17294 (N_17294,N_14994,N_14497);
nor U17295 (N_17295,N_14492,N_14164);
nand U17296 (N_17296,N_12745,N_13011);
nor U17297 (N_17297,N_14986,N_13951);
and U17298 (N_17298,N_14930,N_12652);
xor U17299 (N_17299,N_14044,N_12650);
nor U17300 (N_17300,N_14861,N_14818);
and U17301 (N_17301,N_13435,N_14406);
xnor U17302 (N_17302,N_14189,N_14025);
or U17303 (N_17303,N_14267,N_13081);
or U17304 (N_17304,N_12823,N_14266);
nand U17305 (N_17305,N_13219,N_12924);
nand U17306 (N_17306,N_14295,N_13823);
nand U17307 (N_17307,N_14660,N_14112);
and U17308 (N_17308,N_13531,N_13194);
nand U17309 (N_17309,N_13796,N_14972);
xor U17310 (N_17310,N_13039,N_13268);
or U17311 (N_17311,N_13159,N_14546);
xor U17312 (N_17312,N_13057,N_14886);
xor U17313 (N_17313,N_14895,N_14821);
or U17314 (N_17314,N_13301,N_14939);
and U17315 (N_17315,N_12556,N_13974);
and U17316 (N_17316,N_13967,N_12694);
nor U17317 (N_17317,N_14868,N_12863);
and U17318 (N_17318,N_13847,N_14209);
or U17319 (N_17319,N_14290,N_14838);
xor U17320 (N_17320,N_13575,N_14997);
nor U17321 (N_17321,N_13344,N_12593);
or U17322 (N_17322,N_12649,N_13969);
xnor U17323 (N_17323,N_14614,N_13893);
nand U17324 (N_17324,N_12727,N_13620);
nand U17325 (N_17325,N_14485,N_13298);
or U17326 (N_17326,N_13416,N_13898);
nand U17327 (N_17327,N_14014,N_13590);
nand U17328 (N_17328,N_14895,N_13356);
and U17329 (N_17329,N_13807,N_12622);
xor U17330 (N_17330,N_12729,N_13426);
and U17331 (N_17331,N_13982,N_14367);
nand U17332 (N_17332,N_12698,N_14061);
nand U17333 (N_17333,N_14477,N_12754);
or U17334 (N_17334,N_14776,N_12552);
nand U17335 (N_17335,N_13757,N_12724);
nand U17336 (N_17336,N_13950,N_14905);
or U17337 (N_17337,N_14615,N_12809);
nand U17338 (N_17338,N_14080,N_14947);
nand U17339 (N_17339,N_13325,N_12575);
nor U17340 (N_17340,N_12768,N_12889);
xnor U17341 (N_17341,N_13058,N_13282);
or U17342 (N_17342,N_12586,N_12504);
or U17343 (N_17343,N_14693,N_12979);
xor U17344 (N_17344,N_13194,N_13701);
or U17345 (N_17345,N_12881,N_12649);
and U17346 (N_17346,N_13917,N_12594);
xnor U17347 (N_17347,N_13405,N_13902);
nor U17348 (N_17348,N_12826,N_13337);
and U17349 (N_17349,N_12892,N_13851);
nand U17350 (N_17350,N_12996,N_12904);
nor U17351 (N_17351,N_14373,N_12901);
xor U17352 (N_17352,N_14445,N_13545);
nand U17353 (N_17353,N_13452,N_14943);
nor U17354 (N_17354,N_12640,N_14121);
and U17355 (N_17355,N_14243,N_13731);
and U17356 (N_17356,N_14800,N_13564);
xor U17357 (N_17357,N_14960,N_14111);
and U17358 (N_17358,N_14300,N_13476);
and U17359 (N_17359,N_12974,N_13362);
xnor U17360 (N_17360,N_14129,N_12902);
xnor U17361 (N_17361,N_13203,N_13872);
xor U17362 (N_17362,N_13498,N_13542);
xor U17363 (N_17363,N_14146,N_13338);
nor U17364 (N_17364,N_13098,N_13363);
or U17365 (N_17365,N_13122,N_12775);
nand U17366 (N_17366,N_12580,N_13793);
or U17367 (N_17367,N_14008,N_13839);
nor U17368 (N_17368,N_14237,N_13042);
and U17369 (N_17369,N_12681,N_14671);
xor U17370 (N_17370,N_14721,N_14703);
and U17371 (N_17371,N_14078,N_14305);
or U17372 (N_17372,N_14851,N_12934);
xnor U17373 (N_17373,N_12733,N_14178);
or U17374 (N_17374,N_14066,N_12611);
nand U17375 (N_17375,N_13174,N_14478);
and U17376 (N_17376,N_14882,N_13550);
or U17377 (N_17377,N_14660,N_14584);
xnor U17378 (N_17378,N_14485,N_13706);
and U17379 (N_17379,N_13892,N_14484);
nand U17380 (N_17380,N_12729,N_12574);
xor U17381 (N_17381,N_12887,N_14181);
xor U17382 (N_17382,N_12872,N_13056);
nand U17383 (N_17383,N_13017,N_13673);
and U17384 (N_17384,N_14183,N_12664);
nor U17385 (N_17385,N_14620,N_13223);
nor U17386 (N_17386,N_14262,N_14460);
xor U17387 (N_17387,N_12958,N_14130);
nor U17388 (N_17388,N_14427,N_13952);
and U17389 (N_17389,N_14424,N_13016);
nor U17390 (N_17390,N_13241,N_13431);
xor U17391 (N_17391,N_14795,N_12912);
nor U17392 (N_17392,N_13279,N_14669);
nand U17393 (N_17393,N_13204,N_12829);
xnor U17394 (N_17394,N_12598,N_13863);
nor U17395 (N_17395,N_12548,N_12533);
nor U17396 (N_17396,N_14196,N_13862);
xnor U17397 (N_17397,N_14815,N_14810);
and U17398 (N_17398,N_13411,N_14847);
xnor U17399 (N_17399,N_13629,N_14215);
nand U17400 (N_17400,N_14651,N_13135);
nand U17401 (N_17401,N_13429,N_14364);
xnor U17402 (N_17402,N_12873,N_14541);
xor U17403 (N_17403,N_13023,N_13668);
and U17404 (N_17404,N_13870,N_14698);
nor U17405 (N_17405,N_13757,N_12793);
or U17406 (N_17406,N_13968,N_13347);
or U17407 (N_17407,N_12791,N_13494);
nor U17408 (N_17408,N_13521,N_14869);
xnor U17409 (N_17409,N_14665,N_13195);
and U17410 (N_17410,N_12912,N_12696);
nand U17411 (N_17411,N_13638,N_13277);
xnor U17412 (N_17412,N_13572,N_12759);
xor U17413 (N_17413,N_14815,N_12607);
or U17414 (N_17414,N_14051,N_14535);
nor U17415 (N_17415,N_12503,N_12841);
and U17416 (N_17416,N_13183,N_12810);
or U17417 (N_17417,N_14670,N_14384);
nand U17418 (N_17418,N_12672,N_14654);
nor U17419 (N_17419,N_14608,N_13770);
nand U17420 (N_17420,N_12755,N_13948);
and U17421 (N_17421,N_14358,N_13558);
nand U17422 (N_17422,N_12741,N_13345);
or U17423 (N_17423,N_13718,N_13513);
xor U17424 (N_17424,N_12930,N_14527);
xnor U17425 (N_17425,N_14119,N_13474);
nand U17426 (N_17426,N_13067,N_14205);
nor U17427 (N_17427,N_14636,N_14675);
nand U17428 (N_17428,N_14018,N_13087);
and U17429 (N_17429,N_13424,N_13226);
nand U17430 (N_17430,N_13163,N_13753);
or U17431 (N_17431,N_14383,N_14147);
or U17432 (N_17432,N_14219,N_13519);
xnor U17433 (N_17433,N_13168,N_14998);
xor U17434 (N_17434,N_13145,N_12676);
nand U17435 (N_17435,N_14282,N_13966);
and U17436 (N_17436,N_14005,N_14922);
nor U17437 (N_17437,N_14197,N_13836);
nor U17438 (N_17438,N_13252,N_13114);
nand U17439 (N_17439,N_14156,N_14478);
xnor U17440 (N_17440,N_13705,N_13114);
nand U17441 (N_17441,N_14426,N_12761);
xor U17442 (N_17442,N_13225,N_13855);
xnor U17443 (N_17443,N_12797,N_12693);
nand U17444 (N_17444,N_14359,N_14470);
and U17445 (N_17445,N_13119,N_14189);
nand U17446 (N_17446,N_13480,N_14123);
xnor U17447 (N_17447,N_13054,N_14361);
and U17448 (N_17448,N_12833,N_13703);
and U17449 (N_17449,N_12708,N_12897);
xor U17450 (N_17450,N_14073,N_13284);
and U17451 (N_17451,N_14920,N_13270);
and U17452 (N_17452,N_14773,N_13006);
nand U17453 (N_17453,N_14876,N_12720);
xor U17454 (N_17454,N_14330,N_14934);
nor U17455 (N_17455,N_13562,N_13248);
nor U17456 (N_17456,N_12934,N_13581);
and U17457 (N_17457,N_14040,N_13006);
nand U17458 (N_17458,N_13986,N_13822);
nor U17459 (N_17459,N_12576,N_12983);
nor U17460 (N_17460,N_14518,N_12540);
and U17461 (N_17461,N_13260,N_14396);
nor U17462 (N_17462,N_14681,N_13402);
nand U17463 (N_17463,N_13512,N_14274);
nand U17464 (N_17464,N_13300,N_14570);
nand U17465 (N_17465,N_13073,N_13171);
nor U17466 (N_17466,N_14771,N_12791);
or U17467 (N_17467,N_12921,N_13966);
and U17468 (N_17468,N_14846,N_12730);
nand U17469 (N_17469,N_13117,N_14794);
xnor U17470 (N_17470,N_14711,N_14310);
xor U17471 (N_17471,N_13358,N_13999);
or U17472 (N_17472,N_13060,N_13411);
xor U17473 (N_17473,N_12898,N_14996);
or U17474 (N_17474,N_12501,N_12739);
and U17475 (N_17475,N_13211,N_12776);
or U17476 (N_17476,N_13654,N_12556);
xnor U17477 (N_17477,N_13674,N_14102);
or U17478 (N_17478,N_13777,N_12880);
or U17479 (N_17479,N_14592,N_12775);
xor U17480 (N_17480,N_14879,N_13104);
and U17481 (N_17481,N_13883,N_12782);
and U17482 (N_17482,N_14094,N_12781);
nand U17483 (N_17483,N_14247,N_13519);
or U17484 (N_17484,N_13129,N_13141);
nand U17485 (N_17485,N_14334,N_14883);
and U17486 (N_17486,N_13940,N_12541);
nand U17487 (N_17487,N_12942,N_14479);
and U17488 (N_17488,N_13370,N_14285);
and U17489 (N_17489,N_13441,N_14188);
xnor U17490 (N_17490,N_12843,N_13446);
and U17491 (N_17491,N_14900,N_13926);
xor U17492 (N_17492,N_13127,N_13154);
xnor U17493 (N_17493,N_14643,N_12876);
and U17494 (N_17494,N_14519,N_14008);
nor U17495 (N_17495,N_12508,N_13816);
and U17496 (N_17496,N_13471,N_13755);
nor U17497 (N_17497,N_14024,N_14563);
nand U17498 (N_17498,N_13338,N_14555);
xor U17499 (N_17499,N_14199,N_13298);
xnor U17500 (N_17500,N_15812,N_15384);
xnor U17501 (N_17501,N_16814,N_15354);
or U17502 (N_17502,N_17132,N_16734);
or U17503 (N_17503,N_17473,N_17184);
nand U17504 (N_17504,N_16993,N_15853);
xnor U17505 (N_17505,N_16237,N_17433);
and U17506 (N_17506,N_17074,N_17030);
nand U17507 (N_17507,N_15945,N_17093);
or U17508 (N_17508,N_15326,N_16575);
or U17509 (N_17509,N_15901,N_15111);
nand U17510 (N_17510,N_17039,N_16870);
nor U17511 (N_17511,N_17259,N_16348);
nand U17512 (N_17512,N_15439,N_16883);
nor U17513 (N_17513,N_16083,N_15232);
xor U17514 (N_17514,N_17495,N_15217);
or U17515 (N_17515,N_17373,N_17091);
nand U17516 (N_17516,N_17250,N_15295);
or U17517 (N_17517,N_15026,N_15946);
nand U17518 (N_17518,N_17040,N_16319);
xnor U17519 (N_17519,N_15759,N_16470);
xor U17520 (N_17520,N_15712,N_16151);
or U17521 (N_17521,N_16094,N_15592);
xnor U17522 (N_17522,N_15995,N_16712);
nor U17523 (N_17523,N_16971,N_16843);
xnor U17524 (N_17524,N_16309,N_16748);
nor U17525 (N_17525,N_15125,N_16068);
nand U17526 (N_17526,N_16086,N_17018);
nand U17527 (N_17527,N_15392,N_15615);
xor U17528 (N_17528,N_16245,N_15211);
xnor U17529 (N_17529,N_15842,N_17222);
and U17530 (N_17530,N_15166,N_17151);
and U17531 (N_17531,N_17211,N_16585);
and U17532 (N_17532,N_16477,N_15618);
nand U17533 (N_17533,N_15802,N_17042);
or U17534 (N_17534,N_17029,N_17300);
nand U17535 (N_17535,N_15917,N_16879);
xnor U17536 (N_17536,N_16567,N_17261);
and U17537 (N_17537,N_17068,N_16703);
or U17538 (N_17538,N_16177,N_17244);
nand U17539 (N_17539,N_15892,N_17032);
and U17540 (N_17540,N_16028,N_15997);
nand U17541 (N_17541,N_16218,N_16176);
nor U17542 (N_17542,N_17427,N_17327);
or U17543 (N_17543,N_17139,N_15385);
nand U17544 (N_17544,N_15721,N_15330);
nor U17545 (N_17545,N_16987,N_17426);
nand U17546 (N_17546,N_15181,N_15985);
and U17547 (N_17547,N_16142,N_15776);
nand U17548 (N_17548,N_17106,N_17240);
nor U17549 (N_17549,N_15113,N_15305);
and U17550 (N_17550,N_15383,N_15374);
and U17551 (N_17551,N_16458,N_16440);
nor U17552 (N_17552,N_17306,N_15424);
nor U17553 (N_17553,N_16277,N_15839);
and U17554 (N_17554,N_15414,N_16615);
nand U17555 (N_17555,N_17437,N_17041);
or U17556 (N_17556,N_17435,N_16017);
or U17557 (N_17557,N_16728,N_16653);
xnor U17558 (N_17558,N_15240,N_16099);
xor U17559 (N_17559,N_15192,N_17078);
or U17560 (N_17560,N_16239,N_15662);
or U17561 (N_17561,N_15980,N_15971);
xor U17562 (N_17562,N_17263,N_16763);
or U17563 (N_17563,N_16483,N_15137);
and U17564 (N_17564,N_15926,N_15698);
or U17565 (N_17565,N_16494,N_16493);
nand U17566 (N_17566,N_15937,N_15527);
nor U17567 (N_17567,N_17090,N_17406);
nor U17568 (N_17568,N_16584,N_16383);
or U17569 (N_17569,N_16503,N_15203);
or U17570 (N_17570,N_16906,N_16947);
and U17571 (N_17571,N_15609,N_16121);
nor U17572 (N_17572,N_16327,N_15426);
nand U17573 (N_17573,N_16749,N_16699);
nand U17574 (N_17574,N_16621,N_15179);
nand U17575 (N_17575,N_16290,N_16112);
nand U17576 (N_17576,N_16652,N_16427);
nand U17577 (N_17577,N_16650,N_15018);
xor U17578 (N_17578,N_17123,N_15284);
or U17579 (N_17579,N_17297,N_15611);
and U17580 (N_17580,N_16235,N_16551);
nor U17581 (N_17581,N_16045,N_16469);
nand U17582 (N_17582,N_17095,N_17299);
and U17583 (N_17583,N_16217,N_16233);
nand U17584 (N_17584,N_17447,N_16449);
or U17585 (N_17585,N_15796,N_17432);
xor U17586 (N_17586,N_15331,N_15158);
and U17587 (N_17587,N_16945,N_15906);
xnor U17588 (N_17588,N_16223,N_15627);
or U17589 (N_17589,N_17363,N_16297);
xnor U17590 (N_17590,N_15785,N_15189);
or U17591 (N_17591,N_16027,N_15047);
or U17592 (N_17592,N_16617,N_15480);
nand U17593 (N_17593,N_17186,N_16507);
nand U17594 (N_17594,N_15274,N_17019);
or U17595 (N_17595,N_15630,N_16411);
xnor U17596 (N_17596,N_15228,N_17143);
or U17597 (N_17597,N_17197,N_15780);
or U17598 (N_17598,N_16171,N_16779);
xor U17599 (N_17599,N_16522,N_15220);
or U17600 (N_17600,N_16591,N_15795);
and U17601 (N_17601,N_15098,N_16974);
nor U17602 (N_17602,N_16042,N_15154);
or U17603 (N_17603,N_15883,N_15329);
and U17604 (N_17604,N_17469,N_16680);
nand U17605 (N_17605,N_16131,N_17136);
or U17606 (N_17606,N_17077,N_17146);
nor U17607 (N_17607,N_15935,N_15001);
xnor U17608 (N_17608,N_17434,N_15344);
and U17609 (N_17609,N_17452,N_16289);
nand U17610 (N_17610,N_15754,N_16733);
nor U17611 (N_17611,N_15578,N_15040);
nand U17612 (N_17612,N_16249,N_15248);
xnor U17613 (N_17613,N_16729,N_15895);
or U17614 (N_17614,N_17051,N_16273);
and U17615 (N_17615,N_16926,N_16847);
and U17616 (N_17616,N_15368,N_17203);
and U17617 (N_17617,N_15949,N_15381);
nor U17618 (N_17618,N_15606,N_16528);
and U17619 (N_17619,N_15719,N_16865);
or U17620 (N_17620,N_15782,N_15521);
nand U17621 (N_17621,N_17079,N_15043);
nor U17622 (N_17622,N_16769,N_15556);
or U17623 (N_17623,N_15416,N_17241);
nor U17624 (N_17624,N_15438,N_16101);
xor U17625 (N_17625,N_16828,N_15637);
xor U17626 (N_17626,N_16334,N_17446);
or U17627 (N_17627,N_15273,N_15826);
and U17628 (N_17628,N_15168,N_16124);
xnor U17629 (N_17629,N_16010,N_16534);
xnor U17630 (N_17630,N_15778,N_17122);
or U17631 (N_17631,N_15277,N_17451);
or U17632 (N_17632,N_17298,N_17168);
nor U17633 (N_17633,N_17423,N_17057);
xor U17634 (N_17634,N_16572,N_15535);
nand U17635 (N_17635,N_16946,N_16571);
and U17636 (N_17636,N_16921,N_17142);
nand U17637 (N_17637,N_15509,N_15770);
xnor U17638 (N_17638,N_17127,N_16495);
nor U17639 (N_17639,N_16446,N_15593);
nand U17640 (N_17640,N_15991,N_17471);
xor U17641 (N_17641,N_15049,N_17404);
xnor U17642 (N_17642,N_15089,N_15324);
xnor U17643 (N_17643,N_15436,N_15824);
and U17644 (N_17644,N_16633,N_15897);
and U17645 (N_17645,N_17158,N_16034);
and U17646 (N_17646,N_15886,N_16484);
and U17647 (N_17647,N_15144,N_15707);
or U17648 (N_17648,N_16878,N_17442);
or U17649 (N_17649,N_15038,N_15737);
or U17650 (N_17650,N_15756,N_16443);
or U17651 (N_17651,N_16614,N_16152);
xor U17652 (N_17652,N_16444,N_15687);
and U17653 (N_17653,N_16746,N_17171);
and U17654 (N_17654,N_15915,N_15666);
xnor U17655 (N_17655,N_17475,N_15835);
and U17656 (N_17656,N_15084,N_16800);
nand U17657 (N_17657,N_16658,N_15827);
and U17658 (N_17658,N_15085,N_16471);
and U17659 (N_17659,N_16691,N_15852);
nand U17660 (N_17660,N_17238,N_17135);
or U17661 (N_17661,N_16560,N_16335);
nand U17662 (N_17662,N_15380,N_16163);
nand U17663 (N_17663,N_15610,N_16819);
nor U17664 (N_17664,N_16358,N_17163);
nand U17665 (N_17665,N_17159,N_17118);
xnor U17666 (N_17666,N_15417,N_17008);
nor U17667 (N_17667,N_17431,N_16558);
or U17668 (N_17668,N_15287,N_16675);
or U17669 (N_17669,N_15878,N_15936);
and U17670 (N_17670,N_16808,N_16861);
or U17671 (N_17671,N_17192,N_16807);
xnor U17672 (N_17672,N_17459,N_17190);
or U17673 (N_17673,N_16721,N_15391);
nand U17674 (N_17674,N_17349,N_15619);
xor U17675 (N_17675,N_15280,N_16340);
nand U17676 (N_17676,N_15009,N_17418);
or U17677 (N_17677,N_16399,N_15227);
and U17678 (N_17678,N_15118,N_15742);
and U17679 (N_17679,N_17054,N_15027);
and U17680 (N_17680,N_15891,N_16356);
nand U17681 (N_17681,N_15499,N_15840);
nor U17682 (N_17682,N_15488,N_16917);
and U17683 (N_17683,N_15775,N_16530);
nor U17684 (N_17684,N_16950,N_15703);
or U17685 (N_17685,N_16908,N_15431);
and U17686 (N_17686,N_17398,N_15565);
nor U17687 (N_17687,N_15820,N_17063);
and U17688 (N_17688,N_15024,N_15131);
nor U17689 (N_17689,N_15761,N_15312);
xor U17690 (N_17690,N_15966,N_16566);
and U17691 (N_17691,N_15924,N_15120);
xnor U17692 (N_17692,N_16430,N_16887);
xnor U17693 (N_17693,N_17342,N_16873);
xnor U17694 (N_17694,N_16296,N_17174);
xor U17695 (N_17695,N_17048,N_15572);
or U17696 (N_17696,N_15221,N_17302);
and U17697 (N_17697,N_15710,N_16380);
nand U17698 (N_17698,N_17455,N_15612);
or U17699 (N_17699,N_15779,N_15147);
nor U17700 (N_17700,N_15752,N_16428);
nand U17701 (N_17701,N_16934,N_15903);
nor U17702 (N_17702,N_15806,N_16339);
xor U17703 (N_17703,N_16542,N_17392);
xnor U17704 (N_17704,N_15452,N_16820);
nand U17705 (N_17705,N_15404,N_16665);
nand U17706 (N_17706,N_15000,N_15358);
or U17707 (N_17707,N_17149,N_16106);
xor U17708 (N_17708,N_17361,N_15484);
and U17709 (N_17709,N_16753,N_16231);
nand U17710 (N_17710,N_17110,N_15641);
nand U17711 (N_17711,N_17286,N_15718);
or U17712 (N_17712,N_15366,N_15992);
or U17713 (N_17713,N_15941,N_16127);
and U17714 (N_17714,N_16541,N_16644);
and U17715 (N_17715,N_16715,N_15393);
or U17716 (N_17716,N_16359,N_15979);
and U17717 (N_17717,N_16088,N_16637);
or U17718 (N_17718,N_16225,N_17058);
or U17719 (N_17719,N_17323,N_15469);
nand U17720 (N_17720,N_15164,N_16855);
nor U17721 (N_17721,N_17120,N_15807);
nand U17722 (N_17722,N_15389,N_16561);
nor U17723 (N_17723,N_15573,N_15055);
xnor U17724 (N_17724,N_16352,N_16091);
nor U17725 (N_17725,N_16778,N_15832);
xnor U17726 (N_17726,N_16126,N_15957);
nor U17727 (N_17727,N_16016,N_17346);
xnor U17728 (N_17728,N_15021,N_15516);
nand U17729 (N_17729,N_16418,N_16139);
nand U17730 (N_17730,N_16582,N_15898);
nand U17731 (N_17731,N_15205,N_15256);
or U17732 (N_17732,N_15302,N_17488);
xnor U17733 (N_17733,N_15275,N_15545);
nand U17734 (N_17734,N_15073,N_15003);
xnor U17735 (N_17735,N_15628,N_16222);
or U17736 (N_17736,N_15281,N_16514);
nand U17737 (N_17737,N_16153,N_17417);
and U17738 (N_17738,N_17338,N_17028);
or U17739 (N_17739,N_15023,N_15540);
nand U17740 (N_17740,N_16043,N_16556);
and U17741 (N_17741,N_15307,N_17470);
nor U17742 (N_17742,N_16431,N_16351);
nor U17743 (N_17743,N_15559,N_15973);
xor U17744 (N_17744,N_15373,N_16811);
nor U17745 (N_17745,N_17276,N_16073);
xnor U17746 (N_17746,N_15760,N_15942);
nor U17747 (N_17747,N_16000,N_16674);
xor U17748 (N_17748,N_15011,N_16269);
or U17749 (N_17749,N_16312,N_16825);
nor U17750 (N_17750,N_15485,N_15223);
or U17751 (N_17751,N_15953,N_15555);
and U17752 (N_17752,N_17319,N_15048);
nor U17753 (N_17753,N_15542,N_17231);
xor U17754 (N_17754,N_16647,N_16997);
or U17755 (N_17755,N_15071,N_17484);
and U17756 (N_17756,N_15323,N_15660);
xnor U17757 (N_17757,N_15463,N_16246);
nor U17758 (N_17758,N_16679,N_16254);
or U17759 (N_17759,N_16710,N_16853);
and U17760 (N_17760,N_16620,N_17479);
xnor U17761 (N_17761,N_17026,N_15849);
xnor U17762 (N_17762,N_16859,N_15529);
xnor U17763 (N_17763,N_17109,N_16607);
nand U17764 (N_17764,N_15976,N_15216);
xnor U17765 (N_17765,N_15743,N_15286);
nand U17766 (N_17766,N_17287,N_17152);
nor U17767 (N_17767,N_15097,N_16708);
or U17768 (N_17768,N_16626,N_15146);
nor U17769 (N_17769,N_16041,N_15646);
nor U17770 (N_17770,N_15507,N_17121);
and U17771 (N_17771,N_16848,N_17111);
or U17772 (N_17772,N_15504,N_16550);
and U17773 (N_17773,N_16098,N_15151);
or U17774 (N_17774,N_17044,N_17157);
and U17775 (N_17775,N_15920,N_16146);
nand U17776 (N_17776,N_15190,N_16479);
or U17777 (N_17777,N_15303,N_16473);
nand U17778 (N_17778,N_17464,N_17137);
nor U17779 (N_17779,N_15290,N_16294);
xor U17780 (N_17780,N_16333,N_15601);
and U17781 (N_17781,N_16755,N_16581);
nand U17782 (N_17782,N_16284,N_16777);
or U17783 (N_17783,N_16386,N_15677);
nand U17784 (N_17784,N_15651,N_16285);
or U17785 (N_17785,N_17315,N_15236);
nand U17786 (N_17786,N_15183,N_16595);
or U17787 (N_17787,N_16688,N_15339);
nor U17788 (N_17788,N_16909,N_17007);
nor U17789 (N_17789,N_15254,N_16918);
xnor U17790 (N_17790,N_17397,N_17356);
and U17791 (N_17791,N_16698,N_16024);
xor U17792 (N_17792,N_15500,N_15433);
or U17793 (N_17793,N_16212,N_15667);
nor U17794 (N_17794,N_15828,N_17490);
xor U17795 (N_17795,N_15790,N_17410);
xnor U17796 (N_17796,N_15894,N_16019);
and U17797 (N_17797,N_15680,N_16070);
xnor U17798 (N_17798,N_15948,N_15947);
nor U17799 (N_17799,N_15270,N_15854);
and U17800 (N_17800,N_17049,N_15034);
or U17801 (N_17801,N_15092,N_16508);
xor U17802 (N_17802,N_16377,N_15345);
nor U17803 (N_17803,N_16221,N_16573);
and U17804 (N_17804,N_15296,N_16841);
or U17805 (N_17805,N_15258,N_16476);
and U17806 (N_17806,N_16895,N_15437);
or U17807 (N_17807,N_16743,N_17477);
xnor U17808 (N_17808,N_15640,N_15989);
xnor U17809 (N_17809,N_15411,N_16718);
or U17810 (N_17810,N_16268,N_16738);
nand U17811 (N_17811,N_17295,N_17370);
nand U17812 (N_17812,N_16834,N_15700);
nor U17813 (N_17813,N_15800,N_17036);
xnor U17814 (N_17814,N_16162,N_15874);
nor U17815 (N_17815,N_15467,N_15266);
or U17816 (N_17816,N_16166,N_16329);
and U17817 (N_17817,N_16774,N_15007);
xnor U17818 (N_17818,N_17009,N_15105);
and U17819 (N_17819,N_16320,N_16211);
or U17820 (N_17820,N_16536,N_17156);
nor U17821 (N_17821,N_15006,N_16929);
nor U17822 (N_17822,N_16107,N_17215);
or U17823 (N_17823,N_16662,N_16164);
nor U17824 (N_17824,N_17084,N_16057);
and U17825 (N_17825,N_15259,N_15633);
and U17826 (N_17826,N_16740,N_16750);
and U17827 (N_17827,N_15430,N_16447);
xnor U17828 (N_17828,N_17440,N_15461);
xnor U17829 (N_17829,N_15596,N_15624);
or U17830 (N_17830,N_15420,N_15999);
or U17831 (N_17831,N_16395,N_16668);
and U17832 (N_17832,N_16173,N_15191);
or U17833 (N_17833,N_15093,N_16021);
or U17834 (N_17834,N_15732,N_16578);
and U17835 (N_17835,N_15934,N_16685);
nand U17836 (N_17836,N_17177,N_17462);
nand U17837 (N_17837,N_15174,N_16316);
xor U17838 (N_17838,N_16622,N_16772);
nand U17839 (N_17839,N_16280,N_16817);
nand U17840 (N_17840,N_15621,N_15123);
and U17841 (N_17841,N_17129,N_15132);
or U17842 (N_17842,N_15528,N_16303);
nand U17843 (N_17843,N_16453,N_15696);
and U17844 (N_17844,N_15033,N_15929);
nand U17845 (N_17845,N_16697,N_15199);
xor U17846 (N_17846,N_15153,N_16999);
and U17847 (N_17847,N_17133,N_16160);
nor U17848 (N_17848,N_16323,N_15337);
nand U17849 (N_17849,N_17235,N_15673);
and U17850 (N_17850,N_17085,N_17329);
or U17851 (N_17851,N_15247,N_15402);
nor U17852 (N_17852,N_16326,N_17069);
nand U17853 (N_17853,N_16829,N_16346);
xnor U17854 (N_17854,N_16343,N_16006);
nand U17855 (N_17855,N_16973,N_16149);
or U17856 (N_17856,N_17020,N_16454);
xor U17857 (N_17857,N_16818,N_16511);
and U17858 (N_17858,N_15140,N_17000);
nand U17859 (N_17859,N_15019,N_16457);
or U17860 (N_17860,N_17246,N_15686);
and U17861 (N_17861,N_16948,N_16760);
nand U17862 (N_17862,N_15145,N_16365);
or U17863 (N_17863,N_15141,N_15731);
or U17864 (N_17864,N_15805,N_16336);
nor U17865 (N_17865,N_17234,N_17059);
and U17866 (N_17866,N_16036,N_16806);
xor U17867 (N_17867,N_17296,N_16201);
xnor U17868 (N_17868,N_16498,N_17180);
xnor U17869 (N_17869,N_16373,N_16310);
nand U17870 (N_17870,N_15133,N_15860);
nand U17871 (N_17871,N_16109,N_15714);
xor U17872 (N_17872,N_15473,N_15562);
nand U17873 (N_17873,N_17467,N_15347);
nor U17874 (N_17874,N_16695,N_16451);
nor U17875 (N_17875,N_17169,N_17201);
nor U17876 (N_17876,N_17113,N_16337);
nand U17877 (N_17877,N_15589,N_16396);
nor U17878 (N_17878,N_15341,N_15253);
and U17879 (N_17879,N_16604,N_15557);
or U17880 (N_17880,N_17175,N_16586);
nand U17881 (N_17881,N_15747,N_15445);
nand U17882 (N_17882,N_15520,N_16513);
and U17883 (N_17883,N_15993,N_16810);
or U17884 (N_17884,N_16338,N_15745);
nor U17885 (N_17885,N_15362,N_16900);
xnor U17886 (N_17886,N_16849,N_16158);
xor U17887 (N_17887,N_15727,N_17038);
nand U17888 (N_17888,N_15933,N_16824);
and U17889 (N_17889,N_17027,N_17311);
nor U17890 (N_17890,N_16893,N_15202);
and U17891 (N_17891,N_16884,N_16897);
xor U17892 (N_17892,N_15927,N_16216);
xor U17893 (N_17893,N_16429,N_16243);
xnor U17894 (N_17894,N_15306,N_15625);
xnor U17895 (N_17895,N_15872,N_15738);
xor U17896 (N_17896,N_17303,N_15208);
nor U17897 (N_17897,N_16058,N_17277);
nand U17898 (N_17898,N_15422,N_15334);
nor U17899 (N_17899,N_15665,N_15044);
nor U17900 (N_17900,N_15481,N_15057);
and U17901 (N_17901,N_16354,N_15536);
nand U17902 (N_17902,N_16240,N_15613);
and U17903 (N_17903,N_16672,N_16739);
nand U17904 (N_17904,N_17413,N_17428);
xnor U17905 (N_17905,N_15896,N_15799);
xnor U17906 (N_17906,N_15964,N_15702);
or U17907 (N_17907,N_16549,N_16433);
xnor U17908 (N_17908,N_16627,N_16191);
nor U17909 (N_17909,N_16767,N_17067);
and U17910 (N_17910,N_17396,N_15109);
or U17911 (N_17911,N_17262,N_17460);
xor U17912 (N_17912,N_16785,N_15343);
nand U17913 (N_17913,N_15161,N_15576);
or U17914 (N_17914,N_16899,N_16826);
nor U17915 (N_17915,N_17187,N_15127);
xor U17916 (N_17916,N_17412,N_16353);
nand U17917 (N_17917,N_17482,N_17249);
and U17918 (N_17918,N_17326,N_17284);
nor U17919 (N_17919,N_15209,N_16912);
nand U17920 (N_17920,N_17046,N_15939);
and U17921 (N_17921,N_17436,N_16179);
or U17922 (N_17922,N_17421,N_16678);
nand U17923 (N_17923,N_16417,N_15285);
nand U17924 (N_17924,N_15925,N_16078);
xor U17925 (N_17925,N_15005,N_16659);
nor U17926 (N_17926,N_15950,N_16448);
nand U17927 (N_17927,N_17448,N_15814);
or U17928 (N_17928,N_17202,N_15583);
nand U17929 (N_17929,N_16260,N_17390);
nor U17930 (N_17930,N_16461,N_16804);
nand U17931 (N_17931,N_15278,N_15553);
or U17932 (N_17932,N_15657,N_17489);
nand U17933 (N_17933,N_16293,N_17289);
xor U17934 (N_17934,N_17371,N_16535);
nor U17935 (N_17935,N_15194,N_16903);
nor U17936 (N_17936,N_15954,N_16060);
or U17937 (N_17937,N_15321,N_15602);
nand U17938 (N_17938,N_15333,N_15088);
nand U17939 (N_17939,N_15585,N_16998);
xor U17940 (N_17940,N_16361,N_16518);
nor U17941 (N_17941,N_16317,N_16564);
or U17942 (N_17942,N_16111,N_16989);
xnor U17943 (N_17943,N_15879,N_17154);
and U17944 (N_17944,N_16606,N_15547);
xnor U17945 (N_17945,N_15599,N_16264);
xor U17946 (N_17946,N_17260,N_15722);
nor U17947 (N_17947,N_15196,N_15479);
xnor U17948 (N_17948,N_16587,N_16251);
nor U17949 (N_17949,N_16932,N_16069);
nor U17950 (N_17950,N_15741,N_15716);
or U17951 (N_17951,N_16301,N_15983);
xnor U17952 (N_17952,N_15550,N_16437);
xor U17953 (N_17953,N_16412,N_15272);
nor U17954 (N_17954,N_15268,N_15900);
nor U17955 (N_17955,N_16363,N_16119);
xnor U17956 (N_17956,N_16113,N_16130);
and U17957 (N_17957,N_16725,N_16044);
xnor U17958 (N_17958,N_16464,N_15928);
xor U17959 (N_17959,N_15050,N_15068);
and U17960 (N_17960,N_15880,N_17013);
nand U17961 (N_17961,N_15245,N_15735);
and U17962 (N_17962,N_17394,N_16958);
nand U17963 (N_17963,N_17369,N_16491);
nor U17964 (N_17964,N_16156,N_17468);
nand U17965 (N_17965,N_16636,N_17140);
nand U17966 (N_17966,N_16018,N_16631);
xnor U17967 (N_17967,N_16543,N_16227);
nor U17968 (N_17968,N_17011,N_17131);
nor U17969 (N_17969,N_16482,N_15186);
and U17970 (N_17970,N_15525,N_16082);
or U17971 (N_17971,N_17003,N_16553);
or U17972 (N_17972,N_16362,N_15910);
xnor U17973 (N_17973,N_16816,N_16723);
and U17974 (N_17974,N_16924,N_16271);
nand U17975 (N_17975,N_17278,N_16474);
xnor U17976 (N_17976,N_16704,N_16207);
nor U17977 (N_17977,N_16988,N_16915);
or U17978 (N_17978,N_15902,N_16305);
and U17979 (N_17979,N_16015,N_15739);
xor U17980 (N_17980,N_15590,N_16379);
xor U17981 (N_17981,N_16262,N_17381);
nor U17982 (N_17982,N_15676,N_17247);
nand U17983 (N_17983,N_15315,N_15685);
nand U17984 (N_17984,N_17497,N_16991);
nor U17985 (N_17985,N_15923,N_15159);
xor U17986 (N_17986,N_16540,N_15864);
and U17987 (N_17987,N_16574,N_15283);
or U17988 (N_17988,N_15534,N_15115);
and U17989 (N_17989,N_16832,N_15847);
xor U17990 (N_17990,N_16904,N_17282);
and U17991 (N_17991,N_17336,N_15427);
nor U17992 (N_17992,N_16654,N_15212);
xnor U17993 (N_17993,N_17325,N_17348);
or U17994 (N_17994,N_15830,N_15863);
nand U17995 (N_17995,N_17116,N_17454);
nor U17996 (N_17996,N_16032,N_15455);
and U17997 (N_17997,N_17208,N_17395);
or U17998 (N_17998,N_15691,N_16224);
xor U17999 (N_17999,N_15108,N_16798);
and U18000 (N_18000,N_15442,N_15152);
nand U18001 (N_18001,N_16376,N_17274);
nor U18002 (N_18002,N_17257,N_15866);
xnor U18003 (N_18003,N_16257,N_15390);
and U18004 (N_18004,N_16707,N_15128);
and U18005 (N_18005,N_17310,N_16823);
or U18006 (N_18006,N_15981,N_15905);
xor U18007 (N_18007,N_15564,N_15042);
and U18008 (N_18008,N_16962,N_15031);
nand U18009 (N_18009,N_16406,N_16981);
or U18010 (N_18010,N_15193,N_16986);
nand U18011 (N_18011,N_16026,N_16079);
and U18012 (N_18012,N_16442,N_15204);
nor U18013 (N_18013,N_17387,N_16669);
nand U18014 (N_18014,N_16565,N_15631);
or U18015 (N_18015,N_16624,N_15423);
and U18016 (N_18016,N_16613,N_15963);
nor U18017 (N_18017,N_16882,N_15541);
or U18018 (N_18018,N_15600,N_16141);
nand U18019 (N_18019,N_15054,N_17141);
nand U18020 (N_18020,N_15100,N_15608);
or U18021 (N_18021,N_15282,N_16341);
xnor U18022 (N_18022,N_16521,N_15289);
and U18023 (N_18023,N_15669,N_16432);
nor U18024 (N_18024,N_17364,N_17493);
nand U18025 (N_18025,N_17258,N_16350);
or U18026 (N_18026,N_15299,N_16197);
xor U18027 (N_18027,N_16764,N_16463);
and U18028 (N_18028,N_15308,N_17367);
and U18029 (N_18029,N_15486,N_16939);
xnor U18030 (N_18030,N_16758,N_16439);
or U18031 (N_18031,N_15787,N_15080);
xor U18032 (N_18032,N_15620,N_16259);
or U18033 (N_18033,N_17214,N_15769);
nor U18034 (N_18034,N_17359,N_16372);
and U18035 (N_18035,N_15030,N_15235);
nand U18036 (N_18036,N_15091,N_16056);
xnor U18037 (N_18037,N_16067,N_15661);
nand U18038 (N_18038,N_15792,N_15538);
and U18039 (N_18039,N_16881,N_16593);
or U18040 (N_18040,N_15311,N_16649);
nor U18041 (N_18041,N_15882,N_15032);
xnor U18042 (N_18042,N_15457,N_15548);
and U18043 (N_18043,N_16964,N_16322);
nor U18044 (N_18044,N_15370,N_16398);
nand U18045 (N_18045,N_16189,N_16421);
and U18046 (N_18046,N_15503,N_15498);
or U18047 (N_18047,N_16072,N_15884);
nor U18048 (N_18048,N_16047,N_16786);
and U18049 (N_18049,N_15435,N_15052);
nor U18050 (N_18050,N_15859,N_16095);
xnor U18051 (N_18051,N_17166,N_16941);
or U18052 (N_18052,N_15587,N_15728);
and U18053 (N_18053,N_16896,N_17223);
nand U18054 (N_18054,N_16014,N_15875);
and U18055 (N_18055,N_17499,N_17366);
or U18056 (N_18056,N_16594,N_17466);
nor U18057 (N_18057,N_17309,N_16076);
nand U18058 (N_18058,N_15574,N_16300);
nand U18059 (N_18059,N_16771,N_15348);
xnor U18060 (N_18060,N_17178,N_16527);
and U18061 (N_18061,N_15288,N_16694);
nor U18062 (N_18062,N_17045,N_15246);
and U18063 (N_18063,N_16602,N_16074);
nand U18064 (N_18064,N_15119,N_15683);
or U18065 (N_18065,N_15398,N_15156);
xnor U18066 (N_18066,N_15231,N_15332);
nand U18067 (N_18067,N_17064,N_15143);
or U18068 (N_18068,N_16605,N_15351);
xnor U18069 (N_18069,N_15229,N_16890);
nand U18070 (N_18070,N_17001,N_17453);
xor U18071 (N_18071,N_16456,N_16726);
nand U18072 (N_18072,N_16963,N_17233);
nor U18073 (N_18073,N_17496,N_16858);
and U18074 (N_18074,N_16618,N_16496);
xor U18075 (N_18075,N_16258,N_15195);
and U18076 (N_18076,N_16184,N_15519);
xnor U18077 (N_18077,N_15506,N_16468);
and U18078 (N_18078,N_16759,N_16559);
nand U18079 (N_18079,N_16842,N_15346);
xor U18080 (N_18080,N_16520,N_15165);
and U18081 (N_18081,N_17155,N_15222);
and U18082 (N_18082,N_17424,N_15591);
xor U18083 (N_18083,N_15960,N_15581);
nor U18084 (N_18084,N_15889,N_16115);
nor U18085 (N_18085,N_17320,N_15453);
and U18086 (N_18086,N_16623,N_17419);
nor U18087 (N_18087,N_15579,N_16276);
and U18088 (N_18088,N_15206,N_15508);
and U18089 (N_18089,N_16836,N_17265);
nor U18090 (N_18090,N_16837,N_16690);
or U18091 (N_18091,N_16780,N_16253);
or U18092 (N_18092,N_15397,N_16390);
xnor U18093 (N_18093,N_15010,N_15352);
nand U18094 (N_18094,N_16434,N_16425);
nand U18095 (N_18095,N_15588,N_17445);
and U18096 (N_18096,N_15234,N_15013);
xnor U18097 (N_18097,N_16857,N_16366);
nor U18098 (N_18098,N_16794,N_16592);
xor U18099 (N_18099,N_16588,N_15635);
nand U18100 (N_18100,N_15409,N_17429);
and U18101 (N_18101,N_16270,N_17147);
nor U18102 (N_18102,N_15102,N_16775);
or U18103 (N_18103,N_15734,N_15566);
or U18104 (N_18104,N_15822,N_15793);
xnor U18105 (N_18105,N_17271,N_15642);
or U18106 (N_18106,N_17377,N_15766);
nand U18107 (N_18107,N_17486,N_16081);
xor U18108 (N_18108,N_16247,N_15497);
nand U18109 (N_18109,N_15036,N_15319);
xnor U18110 (N_18110,N_16874,N_17280);
xor U18111 (N_18111,N_16169,N_15784);
nor U18112 (N_18112,N_17096,N_15269);
or U18113 (N_18113,N_17266,N_16922);
nand U18114 (N_18114,N_16210,N_17034);
nand U18115 (N_18115,N_16689,N_17205);
nor U18116 (N_18116,N_15096,N_17088);
xor U18117 (N_18117,N_16325,N_15149);
nor U18118 (N_18118,N_15207,N_16938);
nand U18119 (N_18119,N_16291,N_15255);
nand U18120 (N_18120,N_15413,N_15064);
and U18121 (N_18121,N_15629,N_17405);
and U18122 (N_18122,N_15035,N_15974);
and U18123 (N_18123,N_17207,N_17070);
or U18124 (N_18124,N_15861,N_15363);
nor U18125 (N_18125,N_16255,N_17087);
or U18126 (N_18126,N_16940,N_17425);
or U18127 (N_18127,N_16388,N_17465);
xor U18128 (N_18128,N_17104,N_15359);
or U18129 (N_18129,N_15697,N_16409);
nor U18130 (N_18130,N_16190,N_16892);
nor U18131 (N_18131,N_16554,N_17102);
or U18132 (N_18132,N_16852,N_16480);
nand U18133 (N_18133,N_16875,N_15444);
and U18134 (N_18134,N_16700,N_15626);
xnor U18135 (N_18135,N_17402,N_16783);
and U18136 (N_18136,N_17461,N_16367);
and U18137 (N_18137,N_15532,N_15575);
xnor U18138 (N_18138,N_17360,N_17124);
xor U18139 (N_18139,N_15378,N_17199);
or U18140 (N_18140,N_16092,N_16754);
nor U18141 (N_18141,N_16732,N_15369);
and U18142 (N_18142,N_15705,N_16097);
xnor U18143 (N_18143,N_17403,N_15733);
nand U18144 (N_18144,N_15134,N_15309);
nor U18145 (N_18145,N_16500,N_17232);
xnor U18146 (N_18146,N_16129,N_15386);
nor U18147 (N_18147,N_16040,N_16486);
and U18148 (N_18148,N_15877,N_15659);
or U18149 (N_18149,N_15544,N_16332);
nand U18150 (N_18150,N_15846,N_15355);
nor U18151 (N_18151,N_15515,N_15768);
and U18152 (N_18152,N_15689,N_15713);
xor U18153 (N_18153,N_16701,N_15823);
and U18154 (N_18154,N_16845,N_17195);
nor U18155 (N_18155,N_16478,N_15099);
xor U18156 (N_18156,N_15400,N_17209);
nor U18157 (N_18157,N_15829,N_15294);
and U18158 (N_18158,N_15711,N_16185);
or U18159 (N_18159,N_15751,N_16061);
or U18160 (N_18160,N_17138,N_15142);
nor U18161 (N_18161,N_16570,N_16410);
or U18162 (N_18162,N_16928,N_16720);
nor U18163 (N_18163,N_17248,N_16944);
nand U18164 (N_18164,N_17082,N_15773);
xnor U18165 (N_18165,N_15060,N_17340);
nor U18166 (N_18166,N_15450,N_15616);
xnor U18167 (N_18167,N_15182,N_17357);
xor U18168 (N_18168,N_16002,N_17407);
nand U18169 (N_18169,N_16404,N_16187);
and U18170 (N_18170,N_16096,N_16472);
nor U18171 (N_18171,N_15720,N_17491);
xnor U18172 (N_18172,N_16756,N_15605);
xor U18173 (N_18173,N_16994,N_15172);
nor U18174 (N_18174,N_17376,N_15650);
nand U18175 (N_18175,N_15184,N_16175);
and U18176 (N_18176,N_17061,N_16791);
or U18177 (N_18177,N_15495,N_15265);
and U18178 (N_18178,N_16022,N_15396);
or U18179 (N_18179,N_15644,N_17279);
nor U18180 (N_18180,N_17441,N_16007);
xnor U18181 (N_18181,N_15395,N_16752);
and U18182 (N_18182,N_15675,N_16951);
or U18183 (N_18183,N_15490,N_17388);
xor U18184 (N_18184,N_17251,N_15876);
or U18185 (N_18185,N_15944,N_15938);
nand U18186 (N_18186,N_16306,N_17218);
and U18187 (N_18187,N_15213,N_15148);
xnor U18188 (N_18188,N_17374,N_16544);
nor U18189 (N_18189,N_16046,N_15401);
or U18190 (N_18190,N_15517,N_15746);
or U18191 (N_18191,N_15645,N_16328);
or U18192 (N_18192,N_15918,N_15104);
and U18193 (N_18193,N_17353,N_15474);
or U18194 (N_18194,N_15483,N_15449);
xor U18195 (N_18195,N_15462,N_15376);
xor U18196 (N_18196,N_16597,N_16170);
and U18197 (N_18197,N_15264,N_17333);
or U18198 (N_18198,N_15428,N_16781);
and U18199 (N_18199,N_15750,N_16717);
and U18200 (N_18200,N_16168,N_17162);
and U18201 (N_18201,N_16552,N_16275);
nor U18202 (N_18202,N_17358,N_17224);
nand U18203 (N_18203,N_17380,N_16274);
and U18204 (N_18204,N_17219,N_17227);
xor U18205 (N_18205,N_17411,N_16867);
xnor U18206 (N_18206,N_15167,N_16331);
nor U18207 (N_18207,N_15598,N_16512);
or U18208 (N_18208,N_16736,N_15051);
or U18209 (N_18209,N_15037,N_15238);
and U18210 (N_18210,N_17017,N_16318);
nand U18211 (N_18211,N_15244,N_15571);
xnor U18212 (N_18212,N_16369,N_15679);
xor U18213 (N_18213,N_15293,N_15717);
nand U18214 (N_18214,N_17288,N_16382);
and U18215 (N_18215,N_16295,N_17474);
nor U18216 (N_18216,N_17170,N_16713);
or U18217 (N_18217,N_15114,N_17185);
or U18218 (N_18218,N_16198,N_16250);
nand U18219 (N_18219,N_16742,N_15233);
nand U18220 (N_18220,N_16681,N_16868);
or U18221 (N_18221,N_15492,N_16568);
nor U18222 (N_18222,N_15798,N_17322);
xnor U18223 (N_18223,N_16423,N_16167);
xnor U18224 (N_18224,N_15634,N_15730);
nand U18225 (N_18225,N_16537,N_15399);
nor U18226 (N_18226,N_17150,N_15340);
xor U18227 (N_18227,N_15851,N_16499);
nand U18228 (N_18228,N_16182,N_15514);
nand U18229 (N_18229,N_15129,N_16134);
xor U18230 (N_18230,N_15959,N_16984);
xnor U18231 (N_18231,N_15304,N_16809);
nand U18232 (N_18232,N_16394,N_15017);
or U18233 (N_18233,N_16030,N_16706);
xnor U18234 (N_18234,N_15567,N_15025);
xnor U18235 (N_18235,N_15825,N_15867);
nor U18236 (N_18236,N_16911,N_15988);
and U18237 (N_18237,N_15982,N_15322);
and U18238 (N_18238,N_16995,N_15797);
nand U18239 (N_18239,N_16952,N_17379);
nand U18240 (N_18240,N_17268,N_16302);
and U18241 (N_18241,N_15459,N_15984);
or U18242 (N_18242,N_16265,N_17422);
nand U18243 (N_18243,N_15764,N_17444);
nand U18244 (N_18244,N_16196,N_15511);
and U18245 (N_18245,N_17378,N_17290);
nor U18246 (N_18246,N_16792,N_16776);
or U18247 (N_18247,N_17350,N_16370);
or U18248 (N_18248,N_15382,N_16525);
or U18249 (N_18249,N_15597,N_16504);
nor U18250 (N_18250,N_15725,N_15136);
or U18251 (N_18251,N_15187,N_17160);
nor U18252 (N_18252,N_15360,N_17006);
xor U18253 (N_18253,N_15412,N_16796);
and U18254 (N_18254,N_17115,N_15338);
nand U18255 (N_18255,N_17053,N_15173);
nor U18256 (N_18256,N_16682,N_16801);
nand U18257 (N_18257,N_16242,N_16577);
and U18258 (N_18258,N_17372,N_15978);
xor U18259 (N_18259,N_16719,N_16608);
nand U18260 (N_18260,N_16517,N_15914);
xor U18261 (N_18261,N_15301,N_17275);
nor U18262 (N_18262,N_15922,N_15607);
or U18263 (N_18263,N_15456,N_17443);
nor U18264 (N_18264,N_16093,N_15771);
xnor U18265 (N_18265,N_17339,N_16641);
nor U18266 (N_18266,N_15786,N_17409);
xnor U18267 (N_18267,N_16510,N_15834);
nand U18268 (N_18268,N_16833,N_16628);
nor U18269 (N_18269,N_16108,N_16634);
nor U18270 (N_18270,N_15029,N_16186);
xor U18271 (N_18271,N_16803,N_16632);
xnor U18272 (N_18272,N_15951,N_15850);
nor U18273 (N_18273,N_15524,N_15250);
nand U18274 (N_18274,N_16850,N_15090);
nand U18275 (N_18275,N_15464,N_15004);
nor U18276 (N_18276,N_17341,N_16208);
xor U18277 (N_18277,N_15967,N_15931);
nor U18278 (N_18278,N_17430,N_17213);
or U18279 (N_18279,N_16344,N_16103);
or U18280 (N_18280,N_15478,N_16117);
xor U18281 (N_18281,N_16120,N_16961);
and U18282 (N_18282,N_15817,N_15701);
nand U18283 (N_18283,N_15491,N_15350);
nand U18284 (N_18284,N_17456,N_16515);
or U18285 (N_18285,N_17283,N_15833);
or U18286 (N_18286,N_15361,N_16489);
nor U18287 (N_18287,N_16789,N_16100);
nand U18288 (N_18288,N_16831,N_16533);
xor U18289 (N_18289,N_15969,N_16220);
or U18290 (N_18290,N_15243,N_16601);
xor U18291 (N_18291,N_16384,N_16967);
nor U18292 (N_18292,N_16315,N_16886);
nor U18293 (N_18293,N_15155,N_15791);
or U18294 (N_18294,N_15975,N_16797);
or U18295 (N_18295,N_16228,N_16465);
nand U18296 (N_18296,N_16979,N_16914);
xnor U18297 (N_18297,N_15405,N_16630);
xnor U18298 (N_18298,N_17179,N_16646);
nor U18299 (N_18299,N_17483,N_16860);
xnor U18300 (N_18300,N_17130,N_17071);
or U18301 (N_18301,N_17086,N_17354);
xor U18302 (N_18302,N_16226,N_15261);
nand U18303 (N_18303,N_17216,N_16137);
xnor U18304 (N_18304,N_16660,N_16199);
xnor U18305 (N_18305,N_15074,N_15470);
nor U18306 (N_18306,N_16954,N_16894);
and U18307 (N_18307,N_16526,N_16123);
or U18308 (N_18308,N_16209,N_16716);
xnor U18309 (N_18309,N_16992,N_16747);
nand U18310 (N_18310,N_15921,N_17285);
nand U18311 (N_18311,N_15809,N_17052);
and U18312 (N_18312,N_16165,N_17344);
xor U18313 (N_18313,N_16125,N_16090);
and U18314 (N_18314,N_15990,N_16872);
xnor U18315 (N_18315,N_16144,N_16840);
nand U18316 (N_18316,N_15454,N_15570);
nand U18317 (N_18317,N_15838,N_16400);
xor U18318 (N_18318,N_15215,N_16539);
nand U18319 (N_18319,N_15909,N_16880);
nor U18320 (N_18320,N_15320,N_16898);
nand U18321 (N_18321,N_15056,N_16064);
nor U18322 (N_18322,N_15458,N_17230);
and U18323 (N_18323,N_16762,N_15075);
nor U18324 (N_18324,N_15582,N_16140);
nand U18325 (N_18325,N_15482,N_15487);
or U18326 (N_18326,N_16205,N_15318);
and U18327 (N_18327,N_16345,N_16230);
nand U18328 (N_18328,N_16286,N_17229);
and U18329 (N_18329,N_15095,N_15116);
and U18330 (N_18330,N_16378,N_16299);
nand U18331 (N_18331,N_15169,N_15045);
nor U18332 (N_18332,N_16138,N_15257);
nor U18333 (N_18333,N_16445,N_17337);
nor U18334 (N_18334,N_17145,N_17375);
xor U18335 (N_18335,N_16787,N_16625);
or U18336 (N_18336,N_16488,N_17128);
or U18337 (N_18337,N_15678,N_15740);
and U18338 (N_18338,N_16136,N_15059);
and U18339 (N_18339,N_17439,N_16692);
xnor U18340 (N_18340,N_16116,N_16600);
xor U18341 (N_18341,N_17416,N_16648);
and U18342 (N_18342,N_16714,N_15658);
nand U18343 (N_18343,N_16077,N_15623);
and U18344 (N_18344,N_15443,N_15671);
or U18345 (N_18345,N_16854,N_15692);
xor U18346 (N_18346,N_15058,N_16773);
xnor U18347 (N_18347,N_16349,N_15178);
and U18348 (N_18348,N_16693,N_15162);
nand U18349 (N_18349,N_17055,N_17225);
and U18350 (N_18350,N_16155,N_15531);
and U18351 (N_18351,N_16656,N_17031);
and U18352 (N_18352,N_15079,N_17005);
xnor U18353 (N_18353,N_16524,N_16048);
or U18354 (N_18354,N_15441,N_15690);
or U18355 (N_18355,N_16812,N_16066);
nor U18356 (N_18356,N_16039,N_15139);
and U18357 (N_18357,N_17316,N_16071);
and U18358 (N_18358,N_15082,N_15788);
nand U18359 (N_18359,N_16460,N_17272);
or U18360 (N_18360,N_15135,N_15239);
nand U18361 (N_18361,N_15663,N_15356);
nor U18362 (N_18362,N_15965,N_17384);
nand U18363 (N_18363,N_15406,N_16596);
or U18364 (N_18364,N_15241,N_16279);
nand U18365 (N_18365,N_15081,N_16402);
and U18366 (N_18366,N_16143,N_17002);
nor U18367 (N_18367,N_15408,N_17226);
and U18368 (N_18368,N_16381,N_15020);
xor U18369 (N_18369,N_15622,N_15069);
nand U18370 (N_18370,N_16815,N_15377);
xnor U18371 (N_18371,N_16970,N_17305);
and U18372 (N_18372,N_15899,N_15837);
xor U18373 (N_18373,N_17073,N_17210);
and U18374 (N_18374,N_15501,N_17033);
or U18375 (N_18375,N_15325,N_16502);
nor U18376 (N_18376,N_16104,N_15015);
and U18377 (N_18377,N_15836,N_16422);
nand U18378 (N_18378,N_17196,N_16705);
and U18379 (N_18379,N_15112,N_17035);
nor U18380 (N_18380,N_17253,N_16128);
or U18381 (N_18381,N_15753,N_16105);
nand U18382 (N_18382,N_15314,N_16174);
or U18383 (N_18383,N_17281,N_15577);
or U18384 (N_18384,N_15594,N_16059);
nand U18385 (N_18385,N_17012,N_15972);
nor U18386 (N_18386,N_15549,N_16557);
or U18387 (N_18387,N_17400,N_17457);
or U18388 (N_18388,N_16516,N_15419);
nand U18389 (N_18389,N_15086,N_17107);
nor U18390 (N_18390,N_17307,N_17294);
nor U18391 (N_18391,N_17144,N_16214);
and U18392 (N_18392,N_17352,N_15300);
nor U18393 (N_18393,N_15237,N_15157);
xor U18394 (N_18394,N_16619,N_16959);
and U18395 (N_18395,N_16925,N_15977);
and U18396 (N_18396,N_16065,N_15744);
xor U18397 (N_18397,N_16063,N_15407);
xnor U18398 (N_18398,N_16183,N_15563);
and U18399 (N_18399,N_17101,N_15349);
and U18400 (N_18400,N_16009,N_15881);
or U18401 (N_18401,N_16419,N_17221);
and U18402 (N_18402,N_17383,N_15956);
nand U18403 (N_18403,N_16266,N_16757);
xnor U18404 (N_18404,N_16523,N_15736);
nand U18405 (N_18405,N_17347,N_15072);
nand U18406 (N_18406,N_15758,N_16145);
or U18407 (N_18407,N_17117,N_16157);
and U18408 (N_18408,N_15958,N_16110);
xor U18409 (N_18409,N_15729,N_16569);
and U18410 (N_18410,N_16455,N_16953);
nor U18411 (N_18411,N_16889,N_16937);
xnor U18412 (N_18412,N_17254,N_15335);
and U18413 (N_18413,N_16393,N_16181);
nand U18414 (N_18414,N_15371,N_16407);
xor U18415 (N_18415,N_15388,N_15638);
and U18416 (N_18416,N_15772,N_16545);
nor U18417 (N_18417,N_16876,N_16206);
nor U18418 (N_18418,N_16085,N_16001);
and U18419 (N_18419,N_16416,N_16178);
nand U18420 (N_18420,N_16813,N_17365);
nand U18421 (N_18421,N_15150,N_15715);
and U18422 (N_18422,N_16531,N_15249);
nand U18423 (N_18423,N_16788,N_15094);
or U18424 (N_18424,N_16956,N_17220);
and U18425 (N_18425,N_15225,N_15460);
nor U18426 (N_18426,N_16133,N_16192);
and U18427 (N_18427,N_16696,N_16052);
or U18428 (N_18428,N_15694,N_16888);
or U18429 (N_18429,N_16610,N_16931);
nand U18430 (N_18430,N_16357,N_16683);
and U18431 (N_18431,N_16905,N_16936);
and U18432 (N_18432,N_16612,N_17328);
xor U18433 (N_18433,N_15062,N_15649);
or U18434 (N_18434,N_15087,N_17487);
xnor U18435 (N_18435,N_16248,N_15869);
nor U18436 (N_18436,N_17264,N_15214);
nand U18437 (N_18437,N_17389,N_16972);
and U18438 (N_18438,N_15176,N_15961);
and U18439 (N_18439,N_16761,N_16862);
nor U18440 (N_18440,N_15066,N_15317);
nand U18441 (N_18441,N_17391,N_17334);
or U18442 (N_18442,N_15130,N_15365);
or U18443 (N_18443,N_15940,N_15670);
and U18444 (N_18444,N_16856,N_15364);
nor U18445 (N_18445,N_15313,N_17014);
nand U18446 (N_18446,N_15681,N_16450);
or U18447 (N_18447,N_17269,N_17022);
nor U18448 (N_18448,N_16038,N_16670);
nor U18449 (N_18449,N_16835,N_15765);
or U18450 (N_18450,N_17023,N_15276);
and U18451 (N_18451,N_17172,N_17236);
nand U18452 (N_18452,N_15994,N_16546);
or U18453 (N_18453,N_15505,N_15682);
or U18454 (N_18454,N_16751,N_15636);
nor U18455 (N_18455,N_16003,N_16202);
nor U18456 (N_18456,N_15197,N_17243);
and U18457 (N_18457,N_16330,N_16148);
nand U18458 (N_18458,N_16053,N_16538);
nand U18459 (N_18459,N_16180,N_17415);
nand U18460 (N_18460,N_15171,N_16871);
xor U18461 (N_18461,N_15561,N_16639);
xor U18462 (N_18462,N_15674,N_16241);
xor U18463 (N_18463,N_16966,N_15904);
or U18464 (N_18464,N_17408,N_16204);
and U18465 (N_18465,N_15263,N_17239);
nand U18466 (N_18466,N_16008,N_16598);
nand U18467 (N_18467,N_17362,N_15353);
or U18468 (N_18468,N_15552,N_15873);
nand U18469 (N_18469,N_16532,N_16188);
and U18470 (N_18470,N_16438,N_17189);
and U18471 (N_18471,N_16282,N_17270);
or U18472 (N_18472,N_17228,N_16487);
nor U18473 (N_18473,N_16004,N_15569);
xor U18474 (N_18474,N_15200,N_16805);
and U18475 (N_18475,N_16244,N_16193);
nor U18476 (N_18476,N_15845,N_15617);
and U18477 (N_18477,N_16256,N_17076);
nand U18478 (N_18478,N_15821,N_15870);
nor U18479 (N_18479,N_16949,N_16267);
or U18480 (N_18480,N_16505,N_16342);
and U18481 (N_18481,N_15078,N_17385);
or U18482 (N_18482,N_17188,N_17217);
or U18483 (N_18483,N_16851,N_17485);
nor U18484 (N_18484,N_15810,N_15777);
xnor U18485 (N_18485,N_15117,N_15816);
and U18486 (N_18486,N_16368,N_15170);
nand U18487 (N_18487,N_16467,N_16555);
nor U18488 (N_18488,N_16147,N_16968);
xnor U18489 (N_18489,N_16459,N_15188);
nand U18490 (N_18490,N_15328,N_15425);
or U18491 (N_18491,N_15201,N_17103);
nor U18492 (N_18492,N_15865,N_16827);
nor U18493 (N_18493,N_17438,N_16150);
nor U18494 (N_18494,N_16580,N_17368);
and U18495 (N_18495,N_15526,N_16263);
or U18496 (N_18496,N_16347,N_17324);
nand U18497 (N_18497,N_16590,N_16252);
xnor U18498 (N_18498,N_16033,N_16281);
and U18499 (N_18499,N_16005,N_16314);
and U18500 (N_18500,N_16102,N_16229);
or U18501 (N_18501,N_16709,N_15210);
or U18502 (N_18502,N_15518,N_17165);
or U18503 (N_18503,N_17242,N_16219);
xor U18504 (N_18504,N_15831,N_15652);
or U18505 (N_18505,N_15041,N_15440);
or U18506 (N_18506,N_16307,N_16054);
nand U18507 (N_18507,N_16877,N_16547);
and U18508 (N_18508,N_15789,N_17193);
or U18509 (N_18509,N_16490,N_17015);
nor U18510 (N_18510,N_17083,N_15755);
nor U18511 (N_18511,N_15655,N_16509);
and U18512 (N_18512,N_15801,N_16737);
nor U18513 (N_18513,N_16635,N_15053);
xnor U18514 (N_18514,N_15039,N_16037);
or U18515 (N_18515,N_16089,N_15968);
and U18516 (N_18516,N_15911,N_16023);
or U18517 (N_18517,N_16324,N_15763);
and U18518 (N_18518,N_16935,N_15762);
and U18519 (N_18519,N_17126,N_15008);
and U18520 (N_18520,N_15919,N_17321);
xor U18521 (N_18521,N_16313,N_16677);
and U18522 (N_18522,N_16311,N_15654);
or U18523 (N_18523,N_17125,N_15014);
nand U18524 (N_18524,N_17112,N_16385);
xnor U18525 (N_18525,N_16200,N_16194);
nor U18526 (N_18526,N_17494,N_16839);
nand U18527 (N_18527,N_15468,N_17314);
nand U18528 (N_18528,N_16802,N_17492);
nor U18529 (N_18529,N_17089,N_17255);
or U18530 (N_18530,N_16114,N_17212);
xor U18531 (N_18531,N_16485,N_16519);
nand U18532 (N_18532,N_15291,N_17386);
nor U18533 (N_18533,N_15106,N_16965);
and U18534 (N_18534,N_17308,N_16838);
and U18535 (N_18535,N_15998,N_17037);
nor U18536 (N_18536,N_16664,N_17480);
and U18537 (N_18537,N_16684,N_16288);
and U18538 (N_18538,N_17382,N_15757);
xnor U18539 (N_18539,N_15783,N_16741);
and U18540 (N_18540,N_16927,N_15668);
and U18541 (N_18541,N_17267,N_15415);
xor U18542 (N_18542,N_15451,N_17134);
nor U18543 (N_18543,N_16492,N_16397);
or U18544 (N_18544,N_17393,N_15955);
nor U18545 (N_18545,N_16667,N_16920);
and U18546 (N_18546,N_16923,N_16885);
nor U18547 (N_18547,N_15580,N_16821);
xor U18548 (N_18548,N_15083,N_16506);
xnor U18549 (N_18549,N_15695,N_17047);
xnor U18550 (N_18550,N_16864,N_16308);
nor U18551 (N_18551,N_15708,N_16869);
nor U18552 (N_18552,N_16955,N_17335);
nand U18553 (N_18553,N_16292,N_16589);
or U18554 (N_18554,N_16977,N_16969);
or U18555 (N_18555,N_15124,N_15819);
nand U18556 (N_18556,N_15357,N_16651);
or U18557 (N_18557,N_16655,N_15603);
and U18558 (N_18558,N_16982,N_15063);
nand U18559 (N_18559,N_17450,N_16583);
xnor U18560 (N_18560,N_15558,N_15639);
and U18561 (N_18561,N_16236,N_15546);
nand U18562 (N_18562,N_16159,N_15434);
xor U18563 (N_18563,N_15533,N_16676);
nand U18564 (N_18564,N_15110,N_15046);
or U18565 (N_18565,N_17198,N_16943);
nor U18566 (N_18566,N_15175,N_16298);
xnor U18567 (N_18567,N_16599,N_15379);
and U18568 (N_18568,N_16087,N_16238);
nor U18569 (N_18569,N_16844,N_15070);
or U18570 (N_18570,N_16321,N_16983);
nand U18571 (N_18571,N_15781,N_15316);
nor U18572 (N_18572,N_15327,N_16563);
or U18573 (N_18573,N_16401,N_15890);
or U18574 (N_18574,N_15403,N_16930);
nand U18575 (N_18575,N_15672,N_17312);
xor U18576 (N_18576,N_16360,N_16795);
nor U18577 (N_18577,N_15475,N_17153);
or U18578 (N_18578,N_17245,N_15292);
nand U18579 (N_18579,N_16731,N_16616);
nand U18580 (N_18580,N_16901,N_16232);
or U18581 (N_18581,N_15163,N_17351);
xnor U18582 (N_18582,N_15367,N_16435);
nand U18583 (N_18583,N_17292,N_16661);
xnor U18584 (N_18584,N_16172,N_15543);
and U18585 (N_18585,N_15022,N_17458);
xnor U18586 (N_18586,N_17204,N_16735);
or U18587 (N_18587,N_15107,N_15871);
or U18588 (N_18588,N_16657,N_16426);
xnor U18589 (N_18589,N_15912,N_17463);
nand U18590 (N_18590,N_15512,N_16919);
xor U18591 (N_18591,N_15279,N_17081);
nand U18592 (N_18592,N_15996,N_16122);
nor U18593 (N_18593,N_16799,N_15855);
nand U18594 (N_18594,N_15523,N_16933);
nand U18595 (N_18595,N_15913,N_16375);
xnor U18596 (N_18596,N_16213,N_15930);
xnor U18597 (N_18597,N_16278,N_16916);
nor U18598 (N_18598,N_15723,N_16686);
and U18599 (N_18599,N_15267,N_15180);
nand U18600 (N_18600,N_17173,N_17472);
and U18601 (N_18601,N_17332,N_17313);
xor U18602 (N_18602,N_17481,N_16976);
nor U18603 (N_18603,N_17099,N_15643);
xor U18604 (N_18604,N_16405,N_16671);
and U18605 (N_18605,N_17066,N_16387);
or U18606 (N_18606,N_15952,N_17317);
and U18607 (N_18607,N_15342,N_16579);
xor U18608 (N_18608,N_15077,N_16902);
nor U18609 (N_18609,N_15076,N_17024);
xnor U18610 (N_18610,N_17200,N_16374);
or U18611 (N_18611,N_17167,N_15465);
nor U18612 (N_18612,N_16645,N_16666);
nand U18613 (N_18613,N_15522,N_15604);
xor U18614 (N_18614,N_17498,N_16793);
xor U18615 (N_18615,N_15862,N_15868);
xor U18616 (N_18616,N_15493,N_16629);
xnor U18617 (N_18617,N_16643,N_16050);
nand U18618 (N_18618,N_16745,N_17181);
nand U18619 (N_18619,N_17318,N_15653);
and U18620 (N_18620,N_15709,N_16203);
xnor U18621 (N_18621,N_17293,N_15887);
xor U18622 (N_18622,N_16975,N_16603);
nor U18623 (N_18623,N_15429,N_17021);
nor U18624 (N_18624,N_17164,N_17399);
nand U18625 (N_18625,N_17345,N_15813);
nor U18626 (N_18626,N_16013,N_16035);
xor U18627 (N_18627,N_16371,N_17075);
nor U18628 (N_18628,N_16084,N_17108);
xnor U18629 (N_18629,N_15466,N_15242);
xnor U18630 (N_18630,N_16985,N_15803);
and U18631 (N_18631,N_16768,N_16075);
xor U18632 (N_18632,N_16408,N_15496);
xor U18633 (N_18633,N_15394,N_16055);
nand U18634 (N_18634,N_17194,N_15177);
nor U18635 (N_18635,N_15560,N_16576);
nor U18636 (N_18636,N_15539,N_15185);
or U18637 (N_18637,N_15693,N_17098);
nand U18638 (N_18638,N_16392,N_15432);
or U18639 (N_18639,N_15688,N_16441);
xor U18640 (N_18640,N_16765,N_15804);
and U18641 (N_18641,N_15476,N_15595);
nand U18642 (N_18642,N_16770,N_15916);
or U18643 (N_18643,N_15856,N_16389);
and U18644 (N_18644,N_15198,N_15218);
nand U18645 (N_18645,N_17401,N_15012);
nor U18646 (N_18646,N_16466,N_17330);
xor U18647 (N_18647,N_17414,N_15684);
and U18648 (N_18648,N_16548,N_17420);
or U18649 (N_18649,N_16640,N_15943);
nand U18650 (N_18650,N_15664,N_16702);
or U18651 (N_18651,N_15028,N_16609);
or U18652 (N_18652,N_15808,N_15447);
nand U18653 (N_18653,N_16942,N_16403);
nor U18654 (N_18654,N_15586,N_15537);
xor U18655 (N_18655,N_15219,N_16031);
and U18656 (N_18656,N_15726,N_15067);
xnor U18657 (N_18657,N_15418,N_15848);
or U18658 (N_18658,N_15101,N_16907);
xor U18659 (N_18659,N_17478,N_16611);
nand U18660 (N_18660,N_15699,N_15061);
and U18661 (N_18661,N_16957,N_16863);
nand U18662 (N_18662,N_15126,N_15310);
nand U18663 (N_18663,N_17080,N_15648);
xnor U18664 (N_18664,N_15843,N_15632);
xor U18665 (N_18665,N_15794,N_17291);
nor U18666 (N_18666,N_16822,N_17191);
or U18667 (N_18667,N_15749,N_15647);
nand U18668 (N_18668,N_15986,N_15002);
nand U18669 (N_18669,N_15554,N_15962);
nor U18670 (N_18670,N_15568,N_15065);
nor U18671 (N_18671,N_15226,N_16663);
or U18672 (N_18672,N_15656,N_15489);
nand U18673 (N_18673,N_15502,N_15908);
xor U18674 (N_18674,N_15297,N_16529);
nand U18675 (N_18675,N_16215,N_16012);
or U18676 (N_18676,N_15774,N_17056);
xnor U18677 (N_18677,N_15841,N_17252);
or U18678 (N_18678,N_17273,N_15103);
nor U18679 (N_18679,N_16724,N_16990);
nor U18680 (N_18680,N_15375,N_17331);
nor U18681 (N_18681,N_17343,N_16272);
nand U18682 (N_18682,N_16980,N_15970);
xnor U18683 (N_18683,N_15410,N_16261);
xnor U18684 (N_18684,N_15298,N_17148);
and U18685 (N_18685,N_15421,N_16711);
nand U18686 (N_18686,N_15724,N_15138);
nor U18687 (N_18687,N_16025,N_16364);
nor U18688 (N_18688,N_16475,N_15907);
xnor U18689 (N_18689,N_16287,N_15706);
xnor U18690 (N_18690,N_15387,N_15016);
or U18691 (N_18691,N_17301,N_17025);
or U18692 (N_18692,N_16234,N_16687);
or U18693 (N_18693,N_17062,N_15471);
or U18694 (N_18694,N_15513,N_15160);
nand U18695 (N_18695,N_16497,N_15767);
or U18696 (N_18696,N_16830,N_16722);
xnor U18697 (N_18697,N_16730,N_16436);
and U18698 (N_18698,N_17004,N_15251);
xor U18699 (N_18699,N_15858,N_15614);
or U18700 (N_18700,N_17183,N_17206);
and U18701 (N_18701,N_15448,N_15336);
xnor U18702 (N_18702,N_17476,N_17355);
and U18703 (N_18703,N_15893,N_16727);
and U18704 (N_18704,N_15477,N_15811);
nand U18705 (N_18705,N_15472,N_17119);
or U18706 (N_18706,N_16562,N_17092);
or U18707 (N_18707,N_17256,N_15584);
nand U18708 (N_18708,N_16413,N_17114);
or U18709 (N_18709,N_16051,N_16996);
or U18710 (N_18710,N_15857,N_16910);
nor U18711 (N_18711,N_15494,N_17237);
nand U18712 (N_18712,N_15748,N_17105);
or U18713 (N_18713,N_16462,N_16029);
and U18714 (N_18714,N_17304,N_16135);
nor U18715 (N_18715,N_16132,N_16866);
nand U18716 (N_18716,N_15815,N_16481);
nand U18717 (N_18717,N_15987,N_16355);
or U18718 (N_18718,N_17016,N_16414);
xor U18719 (N_18719,N_15122,N_16011);
nand U18720 (N_18720,N_15510,N_15704);
xnor U18721 (N_18721,N_15818,N_16154);
xor U18722 (N_18722,N_17097,N_16420);
nor U18723 (N_18723,N_16784,N_15844);
nor U18724 (N_18724,N_16304,N_17043);
and U18725 (N_18725,N_15230,N_15932);
nand U18726 (N_18726,N_16195,N_17010);
and U18727 (N_18727,N_16391,N_16673);
and U18728 (N_18728,N_17072,N_17182);
or U18729 (N_18729,N_16452,N_17065);
or U18730 (N_18730,N_16118,N_15224);
nor U18731 (N_18731,N_16782,N_16638);
or U18732 (N_18732,N_16790,N_15372);
or U18733 (N_18733,N_16161,N_15446);
or U18734 (N_18734,N_16978,N_16960);
xnor U18735 (N_18735,N_17094,N_16080);
or U18736 (N_18736,N_16846,N_17176);
and U18737 (N_18737,N_16020,N_16766);
nor U18738 (N_18738,N_17449,N_16891);
or U18739 (N_18739,N_15885,N_17100);
and U18740 (N_18740,N_15530,N_15252);
xor U18741 (N_18741,N_15271,N_15262);
nor U18742 (N_18742,N_16501,N_15888);
nor U18743 (N_18743,N_16424,N_16913);
and U18744 (N_18744,N_16415,N_16062);
or U18745 (N_18745,N_17060,N_16642);
xnor U18746 (N_18746,N_16744,N_16049);
nor U18747 (N_18747,N_15121,N_17050);
nand U18748 (N_18748,N_15551,N_15260);
nand U18749 (N_18749,N_16283,N_17161);
nand U18750 (N_18750,N_15039,N_16593);
nand U18751 (N_18751,N_16852,N_16320);
or U18752 (N_18752,N_16623,N_15930);
and U18753 (N_18753,N_16655,N_16368);
nand U18754 (N_18754,N_16132,N_16649);
nor U18755 (N_18755,N_16351,N_16504);
nor U18756 (N_18756,N_16702,N_17100);
xnor U18757 (N_18757,N_16782,N_15441);
nor U18758 (N_18758,N_17461,N_16082);
xor U18759 (N_18759,N_16443,N_15395);
nor U18760 (N_18760,N_15233,N_15159);
nor U18761 (N_18761,N_15033,N_16254);
xnor U18762 (N_18762,N_15502,N_16200);
nand U18763 (N_18763,N_16728,N_16516);
nor U18764 (N_18764,N_15545,N_17125);
nor U18765 (N_18765,N_16403,N_15609);
or U18766 (N_18766,N_16645,N_15367);
or U18767 (N_18767,N_15209,N_17494);
xor U18768 (N_18768,N_17022,N_17079);
or U18769 (N_18769,N_17423,N_15261);
or U18770 (N_18770,N_15864,N_16589);
xor U18771 (N_18771,N_15401,N_17105);
xor U18772 (N_18772,N_15679,N_15575);
nor U18773 (N_18773,N_15706,N_17471);
nor U18774 (N_18774,N_16665,N_16936);
or U18775 (N_18775,N_16552,N_17179);
xnor U18776 (N_18776,N_15501,N_16956);
xor U18777 (N_18777,N_15196,N_15921);
nor U18778 (N_18778,N_15171,N_17213);
and U18779 (N_18779,N_15271,N_17426);
nand U18780 (N_18780,N_16936,N_16121);
xnor U18781 (N_18781,N_16961,N_15095);
nor U18782 (N_18782,N_17087,N_15454);
nor U18783 (N_18783,N_15183,N_16167);
nand U18784 (N_18784,N_17384,N_16439);
or U18785 (N_18785,N_15517,N_15545);
and U18786 (N_18786,N_16205,N_16123);
xor U18787 (N_18787,N_15569,N_15852);
xnor U18788 (N_18788,N_17106,N_15599);
and U18789 (N_18789,N_15800,N_16482);
nand U18790 (N_18790,N_16724,N_15624);
nand U18791 (N_18791,N_15625,N_16386);
and U18792 (N_18792,N_15005,N_16206);
and U18793 (N_18793,N_16178,N_15698);
xor U18794 (N_18794,N_15831,N_15835);
nor U18795 (N_18795,N_15111,N_15676);
nand U18796 (N_18796,N_15136,N_17297);
and U18797 (N_18797,N_16169,N_16238);
xor U18798 (N_18798,N_16677,N_17429);
and U18799 (N_18799,N_17244,N_17379);
xor U18800 (N_18800,N_16663,N_15874);
xor U18801 (N_18801,N_15111,N_16455);
xor U18802 (N_18802,N_16734,N_15341);
nand U18803 (N_18803,N_16619,N_16740);
or U18804 (N_18804,N_16283,N_15123);
nand U18805 (N_18805,N_16561,N_15189);
xnor U18806 (N_18806,N_16883,N_16148);
xnor U18807 (N_18807,N_16735,N_16754);
nand U18808 (N_18808,N_16252,N_15102);
nand U18809 (N_18809,N_15000,N_17142);
or U18810 (N_18810,N_16562,N_17400);
and U18811 (N_18811,N_15205,N_15335);
or U18812 (N_18812,N_16471,N_16881);
nand U18813 (N_18813,N_17091,N_16705);
or U18814 (N_18814,N_17284,N_16680);
xor U18815 (N_18815,N_17163,N_15813);
xor U18816 (N_18816,N_16326,N_16172);
nand U18817 (N_18817,N_17014,N_17495);
and U18818 (N_18818,N_17325,N_15283);
nand U18819 (N_18819,N_16538,N_17002);
and U18820 (N_18820,N_16959,N_15841);
xnor U18821 (N_18821,N_17093,N_15343);
or U18822 (N_18822,N_17496,N_16163);
nand U18823 (N_18823,N_16914,N_17098);
nor U18824 (N_18824,N_15584,N_17076);
xor U18825 (N_18825,N_17286,N_17325);
nor U18826 (N_18826,N_15686,N_15355);
or U18827 (N_18827,N_16012,N_16412);
or U18828 (N_18828,N_16506,N_16278);
xor U18829 (N_18829,N_16905,N_16256);
nor U18830 (N_18830,N_15102,N_17266);
and U18831 (N_18831,N_16726,N_15776);
and U18832 (N_18832,N_16396,N_16504);
nand U18833 (N_18833,N_16419,N_15451);
and U18834 (N_18834,N_16979,N_15927);
and U18835 (N_18835,N_16098,N_15917);
nor U18836 (N_18836,N_16895,N_15322);
and U18837 (N_18837,N_16451,N_15581);
nor U18838 (N_18838,N_16433,N_15293);
and U18839 (N_18839,N_16647,N_16289);
nand U18840 (N_18840,N_16367,N_15613);
xor U18841 (N_18841,N_16454,N_16827);
nand U18842 (N_18842,N_16431,N_16468);
nor U18843 (N_18843,N_15528,N_17265);
or U18844 (N_18844,N_15972,N_15268);
nand U18845 (N_18845,N_15846,N_16436);
nand U18846 (N_18846,N_16970,N_15177);
nand U18847 (N_18847,N_15719,N_15363);
nor U18848 (N_18848,N_15405,N_15579);
or U18849 (N_18849,N_17306,N_16445);
nor U18850 (N_18850,N_16219,N_15063);
or U18851 (N_18851,N_16402,N_15902);
or U18852 (N_18852,N_15176,N_16675);
xor U18853 (N_18853,N_16921,N_15019);
xnor U18854 (N_18854,N_15313,N_16885);
nor U18855 (N_18855,N_15470,N_15963);
nand U18856 (N_18856,N_16240,N_17386);
or U18857 (N_18857,N_17430,N_16107);
nand U18858 (N_18858,N_15824,N_15505);
xor U18859 (N_18859,N_16507,N_16298);
and U18860 (N_18860,N_15623,N_15553);
nand U18861 (N_18861,N_15289,N_16738);
xnor U18862 (N_18862,N_17011,N_15679);
nand U18863 (N_18863,N_16850,N_15024);
xor U18864 (N_18864,N_16205,N_17401);
and U18865 (N_18865,N_15008,N_15910);
xnor U18866 (N_18866,N_15366,N_15000);
or U18867 (N_18867,N_15542,N_15955);
nor U18868 (N_18868,N_16447,N_15529);
and U18869 (N_18869,N_17320,N_16078);
nand U18870 (N_18870,N_16032,N_15676);
nor U18871 (N_18871,N_16603,N_15700);
nor U18872 (N_18872,N_16882,N_15211);
xor U18873 (N_18873,N_15988,N_17339);
nor U18874 (N_18874,N_15901,N_16211);
nand U18875 (N_18875,N_16932,N_16615);
nand U18876 (N_18876,N_16204,N_16590);
xnor U18877 (N_18877,N_17014,N_17109);
xnor U18878 (N_18878,N_16120,N_16106);
nor U18879 (N_18879,N_15449,N_15444);
nand U18880 (N_18880,N_16240,N_16257);
nor U18881 (N_18881,N_16569,N_15114);
or U18882 (N_18882,N_17201,N_16929);
xor U18883 (N_18883,N_15679,N_16378);
nand U18884 (N_18884,N_17264,N_17383);
and U18885 (N_18885,N_15842,N_17475);
nor U18886 (N_18886,N_16844,N_17364);
nor U18887 (N_18887,N_15457,N_16723);
or U18888 (N_18888,N_16725,N_15367);
nand U18889 (N_18889,N_16897,N_16565);
and U18890 (N_18890,N_16821,N_15584);
and U18891 (N_18891,N_15694,N_16670);
nor U18892 (N_18892,N_17020,N_16526);
xnor U18893 (N_18893,N_17022,N_16462);
or U18894 (N_18894,N_16923,N_16755);
nor U18895 (N_18895,N_15757,N_15365);
xnor U18896 (N_18896,N_15934,N_17188);
or U18897 (N_18897,N_15387,N_16051);
or U18898 (N_18898,N_15570,N_16644);
xor U18899 (N_18899,N_16224,N_17382);
nor U18900 (N_18900,N_16981,N_16596);
or U18901 (N_18901,N_16655,N_16907);
nor U18902 (N_18902,N_15863,N_17368);
or U18903 (N_18903,N_16646,N_17259);
and U18904 (N_18904,N_17346,N_16831);
or U18905 (N_18905,N_16512,N_17429);
xnor U18906 (N_18906,N_15172,N_16768);
and U18907 (N_18907,N_15195,N_15877);
xnor U18908 (N_18908,N_16808,N_15761);
xor U18909 (N_18909,N_15237,N_16264);
nor U18910 (N_18910,N_15647,N_15209);
xnor U18911 (N_18911,N_15719,N_16380);
nor U18912 (N_18912,N_15385,N_15607);
nor U18913 (N_18913,N_16385,N_17290);
or U18914 (N_18914,N_16190,N_16931);
or U18915 (N_18915,N_16494,N_15337);
xor U18916 (N_18916,N_15631,N_15257);
or U18917 (N_18917,N_17188,N_16728);
or U18918 (N_18918,N_17212,N_15080);
and U18919 (N_18919,N_15230,N_16303);
or U18920 (N_18920,N_17087,N_16275);
nor U18921 (N_18921,N_16769,N_17015);
xnor U18922 (N_18922,N_15243,N_16329);
xnor U18923 (N_18923,N_17435,N_15463);
xnor U18924 (N_18924,N_17348,N_15636);
nand U18925 (N_18925,N_15863,N_17087);
and U18926 (N_18926,N_15465,N_16185);
xnor U18927 (N_18927,N_15235,N_15653);
and U18928 (N_18928,N_16912,N_15531);
nand U18929 (N_18929,N_15058,N_15318);
or U18930 (N_18930,N_16088,N_15970);
and U18931 (N_18931,N_16896,N_16129);
nand U18932 (N_18932,N_16931,N_15824);
and U18933 (N_18933,N_15520,N_16520);
nor U18934 (N_18934,N_16786,N_16526);
nand U18935 (N_18935,N_15711,N_15698);
or U18936 (N_18936,N_17415,N_15437);
or U18937 (N_18937,N_16188,N_15003);
xnor U18938 (N_18938,N_15071,N_17207);
nor U18939 (N_18939,N_16321,N_15725);
and U18940 (N_18940,N_16604,N_15398);
or U18941 (N_18941,N_16532,N_16468);
nor U18942 (N_18942,N_15797,N_15300);
xnor U18943 (N_18943,N_16595,N_17018);
and U18944 (N_18944,N_16599,N_17357);
xor U18945 (N_18945,N_15266,N_16330);
or U18946 (N_18946,N_16225,N_16988);
xor U18947 (N_18947,N_15436,N_16194);
and U18948 (N_18948,N_15186,N_15985);
nand U18949 (N_18949,N_15133,N_15576);
nor U18950 (N_18950,N_15861,N_17281);
xor U18951 (N_18951,N_16097,N_15181);
xor U18952 (N_18952,N_16152,N_15549);
and U18953 (N_18953,N_16342,N_17490);
and U18954 (N_18954,N_15413,N_17452);
nand U18955 (N_18955,N_16824,N_16430);
or U18956 (N_18956,N_15484,N_15613);
nor U18957 (N_18957,N_15249,N_16546);
xor U18958 (N_18958,N_16414,N_15902);
nand U18959 (N_18959,N_15380,N_17406);
and U18960 (N_18960,N_15850,N_16867);
nor U18961 (N_18961,N_15020,N_15978);
or U18962 (N_18962,N_16094,N_15779);
nand U18963 (N_18963,N_17149,N_17005);
nand U18964 (N_18964,N_16819,N_16271);
nand U18965 (N_18965,N_15532,N_17408);
nor U18966 (N_18966,N_17152,N_16457);
or U18967 (N_18967,N_16573,N_17476);
or U18968 (N_18968,N_17121,N_15644);
xor U18969 (N_18969,N_15693,N_17453);
nand U18970 (N_18970,N_16133,N_15441);
or U18971 (N_18971,N_16071,N_15896);
nor U18972 (N_18972,N_16954,N_17136);
nand U18973 (N_18973,N_15818,N_16234);
nand U18974 (N_18974,N_17006,N_16980);
nor U18975 (N_18975,N_15450,N_17478);
nand U18976 (N_18976,N_16073,N_16377);
nand U18977 (N_18977,N_15338,N_16383);
or U18978 (N_18978,N_16394,N_15583);
or U18979 (N_18979,N_16351,N_15304);
nand U18980 (N_18980,N_15169,N_15099);
xor U18981 (N_18981,N_15052,N_15280);
nand U18982 (N_18982,N_15793,N_16141);
nand U18983 (N_18983,N_16777,N_16458);
and U18984 (N_18984,N_16375,N_17109);
and U18985 (N_18985,N_16362,N_16783);
or U18986 (N_18986,N_16452,N_15145);
or U18987 (N_18987,N_17036,N_17130);
or U18988 (N_18988,N_17097,N_15844);
nand U18989 (N_18989,N_15650,N_16169);
or U18990 (N_18990,N_17446,N_17254);
xnor U18991 (N_18991,N_15606,N_17329);
nand U18992 (N_18992,N_15014,N_16103);
xnor U18993 (N_18993,N_16363,N_17343);
or U18994 (N_18994,N_16019,N_16575);
or U18995 (N_18995,N_16419,N_15413);
nand U18996 (N_18996,N_15357,N_16558);
and U18997 (N_18997,N_15808,N_15115);
xor U18998 (N_18998,N_16412,N_16280);
or U18999 (N_18999,N_15243,N_16473);
nand U19000 (N_19000,N_15947,N_15935);
nor U19001 (N_19001,N_15837,N_15242);
or U19002 (N_19002,N_16202,N_17029);
nand U19003 (N_19003,N_15072,N_15333);
xor U19004 (N_19004,N_16604,N_16639);
xnor U19005 (N_19005,N_15490,N_16223);
nand U19006 (N_19006,N_17272,N_16336);
and U19007 (N_19007,N_17445,N_15724);
nor U19008 (N_19008,N_15150,N_15246);
nor U19009 (N_19009,N_17460,N_16278);
nor U19010 (N_19010,N_17251,N_16166);
nand U19011 (N_19011,N_17491,N_16304);
and U19012 (N_19012,N_15425,N_16594);
nor U19013 (N_19013,N_16798,N_15781);
nor U19014 (N_19014,N_17223,N_17002);
or U19015 (N_19015,N_15922,N_16217);
nor U19016 (N_19016,N_16697,N_17060);
nor U19017 (N_19017,N_15346,N_15587);
nand U19018 (N_19018,N_16456,N_15392);
nand U19019 (N_19019,N_17166,N_16340);
nor U19020 (N_19020,N_15473,N_15812);
nor U19021 (N_19021,N_16235,N_16314);
nand U19022 (N_19022,N_17202,N_16199);
nand U19023 (N_19023,N_17362,N_15852);
or U19024 (N_19024,N_15899,N_15117);
nand U19025 (N_19025,N_16089,N_15516);
and U19026 (N_19026,N_17118,N_15250);
nor U19027 (N_19027,N_15061,N_17358);
or U19028 (N_19028,N_15938,N_16576);
nand U19029 (N_19029,N_15728,N_15394);
or U19030 (N_19030,N_16688,N_16247);
xor U19031 (N_19031,N_16813,N_15550);
nor U19032 (N_19032,N_16888,N_16691);
and U19033 (N_19033,N_16431,N_17235);
or U19034 (N_19034,N_16891,N_17335);
nor U19035 (N_19035,N_15427,N_15425);
nor U19036 (N_19036,N_16798,N_15990);
xnor U19037 (N_19037,N_15856,N_16312);
or U19038 (N_19038,N_16164,N_16525);
and U19039 (N_19039,N_16683,N_15655);
and U19040 (N_19040,N_17399,N_15982);
xor U19041 (N_19041,N_16558,N_15108);
or U19042 (N_19042,N_15330,N_15208);
and U19043 (N_19043,N_15411,N_15025);
xnor U19044 (N_19044,N_15997,N_17035);
and U19045 (N_19045,N_16522,N_16790);
xor U19046 (N_19046,N_15991,N_17293);
xnor U19047 (N_19047,N_15227,N_16478);
and U19048 (N_19048,N_15930,N_16319);
or U19049 (N_19049,N_15577,N_15142);
or U19050 (N_19050,N_16285,N_15310);
and U19051 (N_19051,N_17393,N_16292);
or U19052 (N_19052,N_15724,N_16159);
nor U19053 (N_19053,N_16567,N_15128);
nand U19054 (N_19054,N_15311,N_16267);
or U19055 (N_19055,N_16754,N_16783);
xnor U19056 (N_19056,N_16583,N_15105);
or U19057 (N_19057,N_17153,N_16244);
xnor U19058 (N_19058,N_16755,N_16004);
and U19059 (N_19059,N_16348,N_17225);
and U19060 (N_19060,N_15902,N_16077);
xnor U19061 (N_19061,N_16168,N_15669);
and U19062 (N_19062,N_15213,N_16594);
and U19063 (N_19063,N_15099,N_15725);
nor U19064 (N_19064,N_16320,N_16872);
nand U19065 (N_19065,N_16880,N_15867);
nand U19066 (N_19066,N_15431,N_15228);
and U19067 (N_19067,N_15396,N_15591);
and U19068 (N_19068,N_15234,N_15138);
xor U19069 (N_19069,N_16409,N_17209);
xor U19070 (N_19070,N_15352,N_16705);
or U19071 (N_19071,N_15313,N_17494);
and U19072 (N_19072,N_15865,N_17085);
or U19073 (N_19073,N_17464,N_15303);
or U19074 (N_19074,N_16743,N_15991);
or U19075 (N_19075,N_15271,N_15899);
nor U19076 (N_19076,N_17472,N_15540);
xor U19077 (N_19077,N_17004,N_15564);
nor U19078 (N_19078,N_15815,N_17303);
and U19079 (N_19079,N_17340,N_16662);
nand U19080 (N_19080,N_15300,N_15102);
xor U19081 (N_19081,N_17387,N_15721);
xor U19082 (N_19082,N_17206,N_15419);
nor U19083 (N_19083,N_16338,N_15545);
nor U19084 (N_19084,N_17180,N_16554);
or U19085 (N_19085,N_15830,N_16005);
or U19086 (N_19086,N_15816,N_17116);
nor U19087 (N_19087,N_15785,N_16433);
xor U19088 (N_19088,N_15146,N_15229);
or U19089 (N_19089,N_17193,N_17137);
or U19090 (N_19090,N_15674,N_15791);
xnor U19091 (N_19091,N_17431,N_15412);
xor U19092 (N_19092,N_17142,N_15399);
or U19093 (N_19093,N_16516,N_16854);
and U19094 (N_19094,N_15270,N_15823);
and U19095 (N_19095,N_15509,N_16466);
and U19096 (N_19096,N_16545,N_15025);
and U19097 (N_19097,N_15542,N_15715);
xor U19098 (N_19098,N_15038,N_17205);
and U19099 (N_19099,N_16001,N_17352);
nor U19100 (N_19100,N_15740,N_17243);
nand U19101 (N_19101,N_16756,N_15897);
nand U19102 (N_19102,N_17326,N_17348);
nor U19103 (N_19103,N_15582,N_17365);
or U19104 (N_19104,N_17317,N_15641);
or U19105 (N_19105,N_17175,N_16272);
xor U19106 (N_19106,N_17484,N_15684);
and U19107 (N_19107,N_17190,N_15470);
nor U19108 (N_19108,N_15016,N_16501);
nand U19109 (N_19109,N_16728,N_17325);
xnor U19110 (N_19110,N_16682,N_17047);
nand U19111 (N_19111,N_15153,N_17139);
xnor U19112 (N_19112,N_17480,N_16621);
and U19113 (N_19113,N_16370,N_16179);
nand U19114 (N_19114,N_17194,N_16682);
nand U19115 (N_19115,N_16834,N_17349);
nor U19116 (N_19116,N_17120,N_16707);
nand U19117 (N_19117,N_16246,N_15995);
nand U19118 (N_19118,N_17140,N_17260);
nor U19119 (N_19119,N_16147,N_15850);
and U19120 (N_19120,N_17299,N_15547);
nand U19121 (N_19121,N_15443,N_16804);
and U19122 (N_19122,N_16116,N_15837);
and U19123 (N_19123,N_15064,N_16978);
xnor U19124 (N_19124,N_15971,N_16148);
and U19125 (N_19125,N_16078,N_17031);
xnor U19126 (N_19126,N_16866,N_16114);
nand U19127 (N_19127,N_16450,N_15601);
xnor U19128 (N_19128,N_16261,N_16320);
nand U19129 (N_19129,N_17116,N_17251);
or U19130 (N_19130,N_16692,N_16380);
and U19131 (N_19131,N_16316,N_17170);
nand U19132 (N_19132,N_15294,N_16595);
nor U19133 (N_19133,N_15702,N_17069);
xnor U19134 (N_19134,N_15255,N_15399);
xor U19135 (N_19135,N_15472,N_15223);
and U19136 (N_19136,N_15553,N_17129);
xnor U19137 (N_19137,N_16995,N_16400);
nor U19138 (N_19138,N_15132,N_17346);
nor U19139 (N_19139,N_17128,N_16314);
and U19140 (N_19140,N_16528,N_16675);
nand U19141 (N_19141,N_15968,N_16257);
or U19142 (N_19142,N_15945,N_15995);
nor U19143 (N_19143,N_17376,N_15944);
nor U19144 (N_19144,N_15344,N_17499);
xnor U19145 (N_19145,N_15113,N_15562);
nand U19146 (N_19146,N_16280,N_17188);
nor U19147 (N_19147,N_17157,N_15986);
nand U19148 (N_19148,N_15747,N_16290);
xnor U19149 (N_19149,N_17187,N_16299);
nor U19150 (N_19150,N_15744,N_16021);
xnor U19151 (N_19151,N_17222,N_15505);
nand U19152 (N_19152,N_16916,N_16976);
nor U19153 (N_19153,N_16430,N_15847);
nor U19154 (N_19154,N_16736,N_15119);
nor U19155 (N_19155,N_15191,N_16186);
xor U19156 (N_19156,N_16382,N_15563);
or U19157 (N_19157,N_15934,N_15388);
nand U19158 (N_19158,N_15629,N_15636);
and U19159 (N_19159,N_16206,N_17374);
nor U19160 (N_19160,N_16416,N_16506);
xnor U19161 (N_19161,N_17273,N_16215);
xnor U19162 (N_19162,N_16440,N_16729);
nor U19163 (N_19163,N_16222,N_15743);
nand U19164 (N_19164,N_16124,N_15399);
nor U19165 (N_19165,N_15494,N_16769);
nand U19166 (N_19166,N_16403,N_17169);
xnor U19167 (N_19167,N_15253,N_15182);
nand U19168 (N_19168,N_16179,N_15986);
xnor U19169 (N_19169,N_15001,N_15158);
or U19170 (N_19170,N_16337,N_16425);
nand U19171 (N_19171,N_17373,N_16813);
and U19172 (N_19172,N_15832,N_15485);
nand U19173 (N_19173,N_15420,N_15948);
and U19174 (N_19174,N_16716,N_16036);
nand U19175 (N_19175,N_15622,N_17060);
nor U19176 (N_19176,N_16098,N_17370);
and U19177 (N_19177,N_15227,N_15213);
or U19178 (N_19178,N_17006,N_15844);
nand U19179 (N_19179,N_16321,N_15882);
nor U19180 (N_19180,N_15139,N_16062);
and U19181 (N_19181,N_16626,N_16956);
xnor U19182 (N_19182,N_15243,N_15758);
and U19183 (N_19183,N_17486,N_15680);
xor U19184 (N_19184,N_15380,N_16174);
nor U19185 (N_19185,N_16087,N_16612);
nand U19186 (N_19186,N_15406,N_16173);
and U19187 (N_19187,N_17153,N_17300);
nand U19188 (N_19188,N_15919,N_16021);
xnor U19189 (N_19189,N_16362,N_16740);
xor U19190 (N_19190,N_16092,N_16707);
nand U19191 (N_19191,N_17133,N_17491);
xor U19192 (N_19192,N_15874,N_15006);
nor U19193 (N_19193,N_15215,N_15674);
and U19194 (N_19194,N_15902,N_17411);
nor U19195 (N_19195,N_16604,N_17054);
nor U19196 (N_19196,N_15357,N_17473);
nand U19197 (N_19197,N_15045,N_16669);
nand U19198 (N_19198,N_16730,N_17483);
and U19199 (N_19199,N_15483,N_16079);
and U19200 (N_19200,N_16861,N_16475);
nand U19201 (N_19201,N_17356,N_15784);
or U19202 (N_19202,N_17202,N_16327);
and U19203 (N_19203,N_15618,N_16622);
or U19204 (N_19204,N_16790,N_16377);
nor U19205 (N_19205,N_16245,N_15622);
or U19206 (N_19206,N_15165,N_16409);
nand U19207 (N_19207,N_15136,N_17225);
or U19208 (N_19208,N_15021,N_16889);
nor U19209 (N_19209,N_16904,N_16217);
and U19210 (N_19210,N_15765,N_16454);
nand U19211 (N_19211,N_15533,N_16397);
or U19212 (N_19212,N_16606,N_15927);
nand U19213 (N_19213,N_16217,N_16292);
and U19214 (N_19214,N_16871,N_17115);
or U19215 (N_19215,N_15771,N_16667);
and U19216 (N_19216,N_16717,N_17439);
nand U19217 (N_19217,N_15136,N_15979);
xor U19218 (N_19218,N_15753,N_15848);
or U19219 (N_19219,N_15505,N_15095);
xnor U19220 (N_19220,N_16473,N_15763);
xor U19221 (N_19221,N_15757,N_15235);
or U19222 (N_19222,N_16667,N_17184);
nand U19223 (N_19223,N_15314,N_15482);
nand U19224 (N_19224,N_15714,N_16689);
xnor U19225 (N_19225,N_15482,N_15412);
xor U19226 (N_19226,N_17260,N_16228);
xor U19227 (N_19227,N_15508,N_17085);
nand U19228 (N_19228,N_16442,N_16982);
and U19229 (N_19229,N_15563,N_15630);
nand U19230 (N_19230,N_17149,N_16633);
xnor U19231 (N_19231,N_15976,N_16753);
and U19232 (N_19232,N_16954,N_16885);
nor U19233 (N_19233,N_16650,N_16646);
nor U19234 (N_19234,N_16298,N_15152);
xnor U19235 (N_19235,N_16651,N_15868);
xor U19236 (N_19236,N_17193,N_15565);
xnor U19237 (N_19237,N_15605,N_16061);
or U19238 (N_19238,N_17386,N_17220);
or U19239 (N_19239,N_17065,N_17028);
or U19240 (N_19240,N_16305,N_17253);
nor U19241 (N_19241,N_15317,N_16238);
xnor U19242 (N_19242,N_16212,N_16732);
nor U19243 (N_19243,N_16884,N_17220);
nand U19244 (N_19244,N_16769,N_16612);
and U19245 (N_19245,N_16139,N_16966);
or U19246 (N_19246,N_16579,N_16672);
nor U19247 (N_19247,N_15421,N_16845);
nor U19248 (N_19248,N_16833,N_16806);
nor U19249 (N_19249,N_15818,N_17224);
and U19250 (N_19250,N_15770,N_15687);
and U19251 (N_19251,N_15213,N_15432);
and U19252 (N_19252,N_15418,N_16817);
and U19253 (N_19253,N_17100,N_16386);
or U19254 (N_19254,N_15596,N_16218);
nand U19255 (N_19255,N_16362,N_16424);
nor U19256 (N_19256,N_15734,N_16868);
xnor U19257 (N_19257,N_16790,N_15805);
or U19258 (N_19258,N_15180,N_16666);
nor U19259 (N_19259,N_16828,N_16356);
xor U19260 (N_19260,N_16229,N_16540);
and U19261 (N_19261,N_15377,N_16644);
or U19262 (N_19262,N_15283,N_15859);
and U19263 (N_19263,N_15774,N_15453);
nor U19264 (N_19264,N_16194,N_15961);
and U19265 (N_19265,N_17386,N_17029);
nand U19266 (N_19266,N_16085,N_16650);
and U19267 (N_19267,N_16878,N_16369);
xnor U19268 (N_19268,N_16770,N_17385);
and U19269 (N_19269,N_15766,N_15439);
nand U19270 (N_19270,N_16261,N_15948);
and U19271 (N_19271,N_15880,N_16186);
or U19272 (N_19272,N_17088,N_17156);
nand U19273 (N_19273,N_16609,N_15125);
or U19274 (N_19274,N_17099,N_16555);
nor U19275 (N_19275,N_15941,N_16452);
or U19276 (N_19276,N_16804,N_15161);
nand U19277 (N_19277,N_17046,N_15623);
and U19278 (N_19278,N_15103,N_15754);
or U19279 (N_19279,N_16705,N_15911);
or U19280 (N_19280,N_16520,N_15458);
xor U19281 (N_19281,N_15646,N_15300);
or U19282 (N_19282,N_16769,N_16186);
xnor U19283 (N_19283,N_17404,N_15053);
nor U19284 (N_19284,N_16705,N_15591);
nor U19285 (N_19285,N_16090,N_15276);
xnor U19286 (N_19286,N_16967,N_15310);
nor U19287 (N_19287,N_15005,N_15090);
xnor U19288 (N_19288,N_15971,N_16196);
xor U19289 (N_19289,N_15545,N_15157);
and U19290 (N_19290,N_15276,N_16609);
and U19291 (N_19291,N_16990,N_17203);
nor U19292 (N_19292,N_16914,N_17467);
nand U19293 (N_19293,N_16729,N_16185);
nor U19294 (N_19294,N_17245,N_16787);
and U19295 (N_19295,N_15057,N_16222);
or U19296 (N_19296,N_15355,N_17451);
nor U19297 (N_19297,N_17217,N_15991);
nor U19298 (N_19298,N_16450,N_15695);
or U19299 (N_19299,N_15043,N_15725);
nor U19300 (N_19300,N_16534,N_16063);
nor U19301 (N_19301,N_17054,N_15477);
and U19302 (N_19302,N_16357,N_16011);
or U19303 (N_19303,N_15191,N_15725);
nand U19304 (N_19304,N_15415,N_17326);
xnor U19305 (N_19305,N_16872,N_15949);
and U19306 (N_19306,N_15727,N_16481);
nor U19307 (N_19307,N_16303,N_16630);
nand U19308 (N_19308,N_16794,N_16627);
nand U19309 (N_19309,N_15741,N_16914);
or U19310 (N_19310,N_17065,N_17097);
nor U19311 (N_19311,N_15213,N_15971);
or U19312 (N_19312,N_15094,N_15249);
nor U19313 (N_19313,N_16327,N_16117);
or U19314 (N_19314,N_15123,N_16320);
and U19315 (N_19315,N_16741,N_16250);
or U19316 (N_19316,N_16305,N_17167);
or U19317 (N_19317,N_16546,N_16661);
or U19318 (N_19318,N_15095,N_15408);
nand U19319 (N_19319,N_15187,N_16173);
or U19320 (N_19320,N_16205,N_16126);
xnor U19321 (N_19321,N_15255,N_16501);
and U19322 (N_19322,N_16867,N_15679);
nor U19323 (N_19323,N_16174,N_15227);
or U19324 (N_19324,N_17067,N_16650);
nor U19325 (N_19325,N_17226,N_17445);
xor U19326 (N_19326,N_16915,N_15023);
nand U19327 (N_19327,N_16399,N_17131);
or U19328 (N_19328,N_16176,N_16936);
and U19329 (N_19329,N_17497,N_16112);
xnor U19330 (N_19330,N_15175,N_16555);
or U19331 (N_19331,N_16891,N_17135);
or U19332 (N_19332,N_16465,N_15448);
nor U19333 (N_19333,N_17362,N_17327);
nor U19334 (N_19334,N_16560,N_16534);
xnor U19335 (N_19335,N_15633,N_17272);
and U19336 (N_19336,N_16190,N_15826);
xnor U19337 (N_19337,N_17423,N_17456);
nor U19338 (N_19338,N_16968,N_15613);
nand U19339 (N_19339,N_17344,N_17380);
xor U19340 (N_19340,N_16145,N_15536);
and U19341 (N_19341,N_15255,N_15982);
xor U19342 (N_19342,N_15943,N_15586);
nor U19343 (N_19343,N_16905,N_15896);
nand U19344 (N_19344,N_15682,N_17249);
xnor U19345 (N_19345,N_15045,N_16529);
and U19346 (N_19346,N_15565,N_15794);
xor U19347 (N_19347,N_17071,N_16627);
nor U19348 (N_19348,N_16394,N_15838);
nor U19349 (N_19349,N_15525,N_15081);
and U19350 (N_19350,N_15785,N_16828);
nand U19351 (N_19351,N_15483,N_15234);
and U19352 (N_19352,N_16443,N_16147);
and U19353 (N_19353,N_16863,N_15877);
and U19354 (N_19354,N_16207,N_16578);
or U19355 (N_19355,N_17071,N_17261);
and U19356 (N_19356,N_15573,N_15424);
nor U19357 (N_19357,N_16796,N_16141);
and U19358 (N_19358,N_16347,N_15577);
nand U19359 (N_19359,N_16323,N_15926);
nand U19360 (N_19360,N_16876,N_15834);
xnor U19361 (N_19361,N_15432,N_16148);
and U19362 (N_19362,N_17132,N_16077);
xor U19363 (N_19363,N_16202,N_17433);
xnor U19364 (N_19364,N_16743,N_16657);
xor U19365 (N_19365,N_16166,N_15668);
nor U19366 (N_19366,N_16248,N_17069);
and U19367 (N_19367,N_17491,N_16022);
and U19368 (N_19368,N_16281,N_16780);
nand U19369 (N_19369,N_17122,N_16407);
or U19370 (N_19370,N_16289,N_15450);
and U19371 (N_19371,N_17423,N_16696);
or U19372 (N_19372,N_15025,N_17427);
nor U19373 (N_19373,N_15342,N_16324);
nand U19374 (N_19374,N_16886,N_15061);
or U19375 (N_19375,N_17143,N_15379);
and U19376 (N_19376,N_15969,N_17201);
nand U19377 (N_19377,N_17261,N_16182);
nor U19378 (N_19378,N_16304,N_15868);
and U19379 (N_19379,N_16910,N_16293);
xor U19380 (N_19380,N_16679,N_16735);
or U19381 (N_19381,N_15365,N_17022);
xnor U19382 (N_19382,N_16499,N_17438);
nor U19383 (N_19383,N_17024,N_16939);
nor U19384 (N_19384,N_16619,N_16054);
nand U19385 (N_19385,N_16320,N_16599);
or U19386 (N_19386,N_16086,N_16810);
nand U19387 (N_19387,N_15574,N_17059);
or U19388 (N_19388,N_15205,N_16817);
or U19389 (N_19389,N_15871,N_16486);
or U19390 (N_19390,N_15251,N_15870);
nor U19391 (N_19391,N_17304,N_17079);
nand U19392 (N_19392,N_16598,N_16528);
nor U19393 (N_19393,N_16205,N_16949);
xor U19394 (N_19394,N_15036,N_16503);
nor U19395 (N_19395,N_17485,N_15531);
and U19396 (N_19396,N_16890,N_15440);
and U19397 (N_19397,N_16358,N_16024);
nand U19398 (N_19398,N_16830,N_16649);
and U19399 (N_19399,N_16967,N_15619);
and U19400 (N_19400,N_16449,N_16304);
or U19401 (N_19401,N_15031,N_16415);
and U19402 (N_19402,N_17213,N_15036);
or U19403 (N_19403,N_15306,N_16256);
and U19404 (N_19404,N_15768,N_15710);
or U19405 (N_19405,N_15965,N_15412);
nand U19406 (N_19406,N_16361,N_16047);
nand U19407 (N_19407,N_15279,N_15458);
nand U19408 (N_19408,N_17270,N_16419);
nor U19409 (N_19409,N_15286,N_16351);
nand U19410 (N_19410,N_15928,N_16125);
and U19411 (N_19411,N_16218,N_15500);
xor U19412 (N_19412,N_16305,N_16153);
nor U19413 (N_19413,N_16872,N_15363);
xor U19414 (N_19414,N_16951,N_17285);
xnor U19415 (N_19415,N_15533,N_16517);
and U19416 (N_19416,N_16338,N_15744);
xor U19417 (N_19417,N_17240,N_15900);
or U19418 (N_19418,N_16597,N_15235);
nand U19419 (N_19419,N_17034,N_16355);
or U19420 (N_19420,N_17060,N_17116);
and U19421 (N_19421,N_16907,N_15880);
nand U19422 (N_19422,N_17435,N_16181);
xor U19423 (N_19423,N_17382,N_16822);
or U19424 (N_19424,N_17101,N_17462);
xnor U19425 (N_19425,N_16104,N_16937);
xor U19426 (N_19426,N_15986,N_17287);
and U19427 (N_19427,N_15455,N_16469);
and U19428 (N_19428,N_16578,N_15624);
or U19429 (N_19429,N_16933,N_16875);
xor U19430 (N_19430,N_15453,N_15458);
nand U19431 (N_19431,N_15933,N_16643);
and U19432 (N_19432,N_16379,N_17465);
or U19433 (N_19433,N_16999,N_15964);
nor U19434 (N_19434,N_15466,N_16152);
nand U19435 (N_19435,N_15347,N_15390);
nor U19436 (N_19436,N_17238,N_15563);
nor U19437 (N_19437,N_16333,N_15253);
and U19438 (N_19438,N_15482,N_16111);
nor U19439 (N_19439,N_15291,N_16115);
nor U19440 (N_19440,N_16496,N_16177);
and U19441 (N_19441,N_17011,N_16070);
nand U19442 (N_19442,N_15382,N_15144);
nand U19443 (N_19443,N_16009,N_17309);
nand U19444 (N_19444,N_15384,N_16479);
or U19445 (N_19445,N_15985,N_16992);
xnor U19446 (N_19446,N_17147,N_15434);
or U19447 (N_19447,N_17113,N_16156);
or U19448 (N_19448,N_16392,N_15215);
and U19449 (N_19449,N_16262,N_17228);
and U19450 (N_19450,N_15586,N_16233);
or U19451 (N_19451,N_15370,N_15684);
nor U19452 (N_19452,N_16453,N_15071);
nor U19453 (N_19453,N_15230,N_15939);
and U19454 (N_19454,N_15813,N_15320);
nand U19455 (N_19455,N_16845,N_15271);
or U19456 (N_19456,N_16311,N_16537);
or U19457 (N_19457,N_16414,N_16010);
nand U19458 (N_19458,N_15472,N_16394);
or U19459 (N_19459,N_15983,N_16285);
xnor U19460 (N_19460,N_17404,N_15164);
or U19461 (N_19461,N_16453,N_15368);
xor U19462 (N_19462,N_15203,N_16211);
nor U19463 (N_19463,N_16770,N_16835);
and U19464 (N_19464,N_17286,N_16826);
and U19465 (N_19465,N_15127,N_16889);
xor U19466 (N_19466,N_17035,N_17200);
or U19467 (N_19467,N_15934,N_15413);
and U19468 (N_19468,N_15350,N_16365);
or U19469 (N_19469,N_17044,N_16200);
nand U19470 (N_19470,N_15198,N_17392);
and U19471 (N_19471,N_16047,N_15182);
xnor U19472 (N_19472,N_15023,N_16446);
and U19473 (N_19473,N_16385,N_16504);
or U19474 (N_19474,N_17049,N_15671);
or U19475 (N_19475,N_16872,N_16352);
xor U19476 (N_19476,N_15779,N_15328);
xor U19477 (N_19477,N_15898,N_17381);
or U19478 (N_19478,N_15046,N_16753);
xor U19479 (N_19479,N_16942,N_16642);
or U19480 (N_19480,N_15025,N_16441);
xor U19481 (N_19481,N_15651,N_16196);
or U19482 (N_19482,N_16975,N_17146);
nand U19483 (N_19483,N_15298,N_16768);
or U19484 (N_19484,N_17041,N_17241);
and U19485 (N_19485,N_15482,N_17085);
nand U19486 (N_19486,N_15013,N_16824);
or U19487 (N_19487,N_15047,N_16849);
and U19488 (N_19488,N_17086,N_16533);
nand U19489 (N_19489,N_16258,N_15601);
xor U19490 (N_19490,N_15757,N_17094);
xor U19491 (N_19491,N_15164,N_15842);
nor U19492 (N_19492,N_17062,N_16397);
nor U19493 (N_19493,N_16135,N_16396);
and U19494 (N_19494,N_16480,N_15652);
or U19495 (N_19495,N_16154,N_15783);
nand U19496 (N_19496,N_16975,N_15423);
and U19497 (N_19497,N_16778,N_16751);
xor U19498 (N_19498,N_16380,N_17098);
or U19499 (N_19499,N_16228,N_15608);
or U19500 (N_19500,N_15827,N_15534);
and U19501 (N_19501,N_16932,N_16732);
nor U19502 (N_19502,N_17134,N_15032);
xnor U19503 (N_19503,N_16163,N_16411);
xor U19504 (N_19504,N_16675,N_15928);
nand U19505 (N_19505,N_15258,N_16367);
or U19506 (N_19506,N_17200,N_15411);
nand U19507 (N_19507,N_17002,N_17322);
nor U19508 (N_19508,N_16635,N_15856);
or U19509 (N_19509,N_16900,N_17298);
or U19510 (N_19510,N_15515,N_16826);
nor U19511 (N_19511,N_15020,N_17080);
nand U19512 (N_19512,N_17479,N_15620);
xnor U19513 (N_19513,N_16049,N_16025);
nor U19514 (N_19514,N_15028,N_17071);
nor U19515 (N_19515,N_15174,N_16671);
nand U19516 (N_19516,N_17001,N_17280);
nor U19517 (N_19517,N_17126,N_15133);
nor U19518 (N_19518,N_16399,N_16330);
and U19519 (N_19519,N_16698,N_16105);
or U19520 (N_19520,N_16280,N_16335);
or U19521 (N_19521,N_17167,N_15935);
or U19522 (N_19522,N_15273,N_17480);
nand U19523 (N_19523,N_15423,N_16982);
or U19524 (N_19524,N_15992,N_16155);
nand U19525 (N_19525,N_15101,N_15505);
or U19526 (N_19526,N_17154,N_16031);
or U19527 (N_19527,N_16735,N_16412);
nand U19528 (N_19528,N_16288,N_15004);
nand U19529 (N_19529,N_15877,N_15597);
or U19530 (N_19530,N_16404,N_17145);
nor U19531 (N_19531,N_17467,N_17292);
nor U19532 (N_19532,N_17163,N_16834);
nor U19533 (N_19533,N_15082,N_16965);
or U19534 (N_19534,N_17151,N_17363);
nand U19535 (N_19535,N_15472,N_17242);
or U19536 (N_19536,N_16941,N_16399);
or U19537 (N_19537,N_15650,N_16513);
nand U19538 (N_19538,N_16583,N_15876);
xnor U19539 (N_19539,N_17085,N_15039);
or U19540 (N_19540,N_15595,N_17418);
or U19541 (N_19541,N_16967,N_15693);
or U19542 (N_19542,N_16164,N_15314);
or U19543 (N_19543,N_15614,N_16287);
and U19544 (N_19544,N_15756,N_17113);
and U19545 (N_19545,N_15806,N_15273);
and U19546 (N_19546,N_16093,N_15393);
and U19547 (N_19547,N_15044,N_16502);
and U19548 (N_19548,N_16947,N_17285);
or U19549 (N_19549,N_15316,N_17451);
and U19550 (N_19550,N_15856,N_16319);
nand U19551 (N_19551,N_15776,N_15232);
and U19552 (N_19552,N_15244,N_17296);
xor U19553 (N_19553,N_16548,N_17241);
nand U19554 (N_19554,N_16898,N_15481);
and U19555 (N_19555,N_17316,N_15998);
or U19556 (N_19556,N_15598,N_17457);
nand U19557 (N_19557,N_16743,N_16721);
or U19558 (N_19558,N_15801,N_15962);
xnor U19559 (N_19559,N_17179,N_15311);
nor U19560 (N_19560,N_16741,N_17005);
and U19561 (N_19561,N_17122,N_15889);
nor U19562 (N_19562,N_16578,N_17054);
xor U19563 (N_19563,N_16303,N_16629);
nand U19564 (N_19564,N_16809,N_15014);
and U19565 (N_19565,N_15204,N_16336);
nand U19566 (N_19566,N_15658,N_17419);
nor U19567 (N_19567,N_17490,N_15361);
nand U19568 (N_19568,N_16651,N_17463);
and U19569 (N_19569,N_17059,N_15263);
xor U19570 (N_19570,N_15359,N_17441);
xor U19571 (N_19571,N_15930,N_16166);
nand U19572 (N_19572,N_16834,N_16326);
xor U19573 (N_19573,N_15970,N_16142);
and U19574 (N_19574,N_16600,N_16768);
and U19575 (N_19575,N_17181,N_15475);
or U19576 (N_19576,N_17098,N_16826);
xor U19577 (N_19577,N_15943,N_16261);
or U19578 (N_19578,N_15527,N_16375);
nor U19579 (N_19579,N_15491,N_15479);
nand U19580 (N_19580,N_16570,N_16789);
or U19581 (N_19581,N_16209,N_16461);
and U19582 (N_19582,N_15716,N_16992);
or U19583 (N_19583,N_15352,N_15710);
nand U19584 (N_19584,N_15249,N_16308);
nand U19585 (N_19585,N_16385,N_15567);
or U19586 (N_19586,N_17189,N_16120);
xnor U19587 (N_19587,N_15545,N_15723);
nand U19588 (N_19588,N_15038,N_17447);
nor U19589 (N_19589,N_16949,N_15089);
or U19590 (N_19590,N_15296,N_17399);
and U19591 (N_19591,N_16615,N_17310);
nand U19592 (N_19592,N_15299,N_16025);
nor U19593 (N_19593,N_15591,N_15141);
and U19594 (N_19594,N_15214,N_15532);
and U19595 (N_19595,N_15682,N_15886);
and U19596 (N_19596,N_17031,N_15655);
or U19597 (N_19597,N_16870,N_16927);
nand U19598 (N_19598,N_15443,N_16828);
and U19599 (N_19599,N_17007,N_17095);
nand U19600 (N_19600,N_16619,N_16666);
nand U19601 (N_19601,N_15378,N_15686);
nor U19602 (N_19602,N_16401,N_17305);
xnor U19603 (N_19603,N_15932,N_15268);
and U19604 (N_19604,N_17143,N_15040);
nor U19605 (N_19605,N_16521,N_15485);
xnor U19606 (N_19606,N_16674,N_16201);
xnor U19607 (N_19607,N_15179,N_15973);
nor U19608 (N_19608,N_15103,N_17208);
and U19609 (N_19609,N_17145,N_15801);
xor U19610 (N_19610,N_16525,N_15597);
xor U19611 (N_19611,N_16868,N_15348);
and U19612 (N_19612,N_16628,N_15787);
or U19613 (N_19613,N_15775,N_16568);
nand U19614 (N_19614,N_17296,N_15674);
nand U19615 (N_19615,N_16990,N_15937);
or U19616 (N_19616,N_15033,N_17082);
or U19617 (N_19617,N_17481,N_16013);
or U19618 (N_19618,N_15054,N_16933);
and U19619 (N_19619,N_16766,N_17167);
and U19620 (N_19620,N_16233,N_16205);
or U19621 (N_19621,N_15089,N_16146);
or U19622 (N_19622,N_15024,N_16673);
or U19623 (N_19623,N_17161,N_17427);
or U19624 (N_19624,N_16823,N_17003);
and U19625 (N_19625,N_15256,N_17283);
or U19626 (N_19626,N_15735,N_17327);
nor U19627 (N_19627,N_15901,N_16473);
or U19628 (N_19628,N_15056,N_15769);
or U19629 (N_19629,N_15249,N_16010);
or U19630 (N_19630,N_16290,N_16933);
or U19631 (N_19631,N_15900,N_16827);
nor U19632 (N_19632,N_17254,N_16432);
nor U19633 (N_19633,N_15724,N_15259);
xor U19634 (N_19634,N_15129,N_15922);
or U19635 (N_19635,N_15718,N_17059);
or U19636 (N_19636,N_15735,N_15849);
or U19637 (N_19637,N_15929,N_16899);
nor U19638 (N_19638,N_15883,N_17497);
and U19639 (N_19639,N_15497,N_15964);
nand U19640 (N_19640,N_15635,N_16241);
xnor U19641 (N_19641,N_15436,N_15597);
or U19642 (N_19642,N_15597,N_15424);
or U19643 (N_19643,N_16500,N_15220);
xnor U19644 (N_19644,N_15098,N_17401);
nand U19645 (N_19645,N_15874,N_15064);
nor U19646 (N_19646,N_15416,N_16309);
xnor U19647 (N_19647,N_15192,N_17370);
xnor U19648 (N_19648,N_16814,N_15003);
nand U19649 (N_19649,N_15656,N_17132);
and U19650 (N_19650,N_16756,N_17435);
or U19651 (N_19651,N_15265,N_15405);
xnor U19652 (N_19652,N_15659,N_16216);
nor U19653 (N_19653,N_16044,N_15046);
xnor U19654 (N_19654,N_16412,N_16602);
xnor U19655 (N_19655,N_17406,N_16791);
or U19656 (N_19656,N_15960,N_15616);
nor U19657 (N_19657,N_17304,N_15958);
xnor U19658 (N_19658,N_15474,N_15890);
and U19659 (N_19659,N_16571,N_15744);
nor U19660 (N_19660,N_16009,N_16305);
nor U19661 (N_19661,N_16214,N_15681);
nor U19662 (N_19662,N_17237,N_16802);
nand U19663 (N_19663,N_16660,N_15620);
nand U19664 (N_19664,N_17050,N_17186);
xor U19665 (N_19665,N_17287,N_15653);
nor U19666 (N_19666,N_16899,N_16095);
nor U19667 (N_19667,N_15050,N_17068);
nor U19668 (N_19668,N_16808,N_15915);
and U19669 (N_19669,N_17436,N_16097);
nor U19670 (N_19670,N_15830,N_16930);
nor U19671 (N_19671,N_16115,N_16816);
xnor U19672 (N_19672,N_15375,N_15667);
xor U19673 (N_19673,N_15199,N_16351);
or U19674 (N_19674,N_16871,N_16321);
nor U19675 (N_19675,N_16958,N_15614);
and U19676 (N_19676,N_16754,N_16232);
and U19677 (N_19677,N_16565,N_16315);
nand U19678 (N_19678,N_16749,N_17046);
nor U19679 (N_19679,N_16635,N_15083);
nand U19680 (N_19680,N_17332,N_16375);
nand U19681 (N_19681,N_15974,N_15412);
nor U19682 (N_19682,N_16317,N_16559);
and U19683 (N_19683,N_17457,N_16784);
nand U19684 (N_19684,N_15818,N_17274);
nor U19685 (N_19685,N_15409,N_15056);
and U19686 (N_19686,N_15106,N_15749);
nor U19687 (N_19687,N_16739,N_16132);
and U19688 (N_19688,N_16801,N_15943);
xnor U19689 (N_19689,N_16786,N_16565);
nand U19690 (N_19690,N_16849,N_15109);
nor U19691 (N_19691,N_17163,N_16600);
xor U19692 (N_19692,N_15228,N_16794);
xnor U19693 (N_19693,N_17201,N_15650);
xnor U19694 (N_19694,N_16048,N_17486);
or U19695 (N_19695,N_17095,N_16704);
and U19696 (N_19696,N_15023,N_16219);
and U19697 (N_19697,N_16575,N_16656);
xor U19698 (N_19698,N_16448,N_16561);
nor U19699 (N_19699,N_17400,N_15959);
and U19700 (N_19700,N_15091,N_16283);
or U19701 (N_19701,N_16319,N_15719);
or U19702 (N_19702,N_16514,N_17334);
nor U19703 (N_19703,N_17290,N_15988);
and U19704 (N_19704,N_15373,N_16373);
nor U19705 (N_19705,N_17218,N_15898);
or U19706 (N_19706,N_15770,N_16791);
nor U19707 (N_19707,N_17375,N_16427);
nand U19708 (N_19708,N_15780,N_17389);
nor U19709 (N_19709,N_16837,N_15970);
or U19710 (N_19710,N_16610,N_16567);
and U19711 (N_19711,N_15684,N_16684);
or U19712 (N_19712,N_16745,N_16411);
and U19713 (N_19713,N_15519,N_15932);
nor U19714 (N_19714,N_15990,N_15725);
nand U19715 (N_19715,N_16332,N_16187);
or U19716 (N_19716,N_16280,N_16314);
and U19717 (N_19717,N_15158,N_16906);
xor U19718 (N_19718,N_17000,N_15165);
nand U19719 (N_19719,N_16752,N_16029);
nor U19720 (N_19720,N_16164,N_16260);
nand U19721 (N_19721,N_16384,N_15084);
nand U19722 (N_19722,N_15646,N_15909);
and U19723 (N_19723,N_17181,N_15056);
nor U19724 (N_19724,N_15792,N_17498);
nand U19725 (N_19725,N_15750,N_15590);
or U19726 (N_19726,N_15013,N_15511);
or U19727 (N_19727,N_17464,N_16257);
or U19728 (N_19728,N_16052,N_15176);
nand U19729 (N_19729,N_16915,N_16215);
nor U19730 (N_19730,N_15806,N_17143);
or U19731 (N_19731,N_15959,N_16359);
and U19732 (N_19732,N_16146,N_15431);
or U19733 (N_19733,N_16026,N_16945);
nand U19734 (N_19734,N_16913,N_16395);
or U19735 (N_19735,N_15954,N_16816);
xnor U19736 (N_19736,N_16398,N_15013);
and U19737 (N_19737,N_15658,N_15780);
and U19738 (N_19738,N_15993,N_15244);
or U19739 (N_19739,N_15657,N_15186);
nor U19740 (N_19740,N_16266,N_15137);
and U19741 (N_19741,N_16982,N_17451);
and U19742 (N_19742,N_16756,N_15052);
and U19743 (N_19743,N_15382,N_15772);
nor U19744 (N_19744,N_15272,N_16967);
nor U19745 (N_19745,N_16472,N_16996);
or U19746 (N_19746,N_15705,N_16141);
nand U19747 (N_19747,N_17385,N_15842);
and U19748 (N_19748,N_15973,N_17402);
and U19749 (N_19749,N_17335,N_17414);
xor U19750 (N_19750,N_15892,N_15336);
xnor U19751 (N_19751,N_17367,N_15251);
nor U19752 (N_19752,N_16725,N_15754);
nor U19753 (N_19753,N_16007,N_15292);
nand U19754 (N_19754,N_17023,N_15408);
or U19755 (N_19755,N_15325,N_15649);
or U19756 (N_19756,N_16480,N_15678);
nor U19757 (N_19757,N_17078,N_15926);
nor U19758 (N_19758,N_16113,N_16623);
or U19759 (N_19759,N_15904,N_16241);
nor U19760 (N_19760,N_16638,N_16524);
and U19761 (N_19761,N_16608,N_16997);
xnor U19762 (N_19762,N_16725,N_15251);
nor U19763 (N_19763,N_16204,N_17281);
nand U19764 (N_19764,N_16786,N_16740);
and U19765 (N_19765,N_15190,N_16630);
or U19766 (N_19766,N_17085,N_16045);
and U19767 (N_19767,N_15654,N_15872);
or U19768 (N_19768,N_17491,N_17048);
nand U19769 (N_19769,N_15874,N_16107);
nor U19770 (N_19770,N_16355,N_16176);
xnor U19771 (N_19771,N_15720,N_16072);
nand U19772 (N_19772,N_15030,N_17219);
or U19773 (N_19773,N_17405,N_16941);
nand U19774 (N_19774,N_17074,N_15598);
or U19775 (N_19775,N_15306,N_15928);
and U19776 (N_19776,N_15023,N_16401);
nor U19777 (N_19777,N_15411,N_17228);
nor U19778 (N_19778,N_16730,N_17316);
nor U19779 (N_19779,N_16480,N_16629);
nand U19780 (N_19780,N_15293,N_16467);
nor U19781 (N_19781,N_16531,N_16471);
or U19782 (N_19782,N_17389,N_15597);
and U19783 (N_19783,N_16671,N_15745);
and U19784 (N_19784,N_16210,N_16072);
and U19785 (N_19785,N_17414,N_15832);
nand U19786 (N_19786,N_16124,N_17314);
xnor U19787 (N_19787,N_15511,N_15018);
nand U19788 (N_19788,N_17059,N_15236);
or U19789 (N_19789,N_16417,N_16630);
and U19790 (N_19790,N_15111,N_15073);
or U19791 (N_19791,N_16370,N_16951);
nand U19792 (N_19792,N_16673,N_15071);
and U19793 (N_19793,N_16393,N_15853);
and U19794 (N_19794,N_15483,N_17094);
or U19795 (N_19795,N_15542,N_15697);
nor U19796 (N_19796,N_15517,N_16226);
nand U19797 (N_19797,N_16264,N_16168);
xnor U19798 (N_19798,N_15498,N_15367);
xor U19799 (N_19799,N_15351,N_16611);
xor U19800 (N_19800,N_16528,N_17382);
nand U19801 (N_19801,N_16176,N_17232);
or U19802 (N_19802,N_15113,N_15556);
nand U19803 (N_19803,N_15780,N_16383);
or U19804 (N_19804,N_16972,N_16916);
or U19805 (N_19805,N_16565,N_15613);
xnor U19806 (N_19806,N_17228,N_16255);
and U19807 (N_19807,N_15080,N_15878);
and U19808 (N_19808,N_17433,N_16557);
xnor U19809 (N_19809,N_16427,N_16889);
nor U19810 (N_19810,N_15811,N_17120);
nand U19811 (N_19811,N_16859,N_16213);
nand U19812 (N_19812,N_15772,N_16998);
nand U19813 (N_19813,N_16995,N_16218);
nor U19814 (N_19814,N_15317,N_15852);
nor U19815 (N_19815,N_17269,N_17293);
or U19816 (N_19816,N_16518,N_17201);
xor U19817 (N_19817,N_17175,N_15011);
nand U19818 (N_19818,N_15470,N_16111);
nor U19819 (N_19819,N_16413,N_15204);
nand U19820 (N_19820,N_17135,N_16655);
and U19821 (N_19821,N_16686,N_16268);
and U19822 (N_19822,N_15672,N_16013);
and U19823 (N_19823,N_15052,N_15008);
nor U19824 (N_19824,N_16229,N_16552);
xor U19825 (N_19825,N_15159,N_16656);
nor U19826 (N_19826,N_15911,N_15938);
nor U19827 (N_19827,N_17172,N_15746);
nand U19828 (N_19828,N_15530,N_15406);
nor U19829 (N_19829,N_16514,N_15723);
and U19830 (N_19830,N_15986,N_16999);
and U19831 (N_19831,N_17309,N_15551);
nand U19832 (N_19832,N_15483,N_16709);
or U19833 (N_19833,N_17136,N_15218);
nand U19834 (N_19834,N_17166,N_15071);
xnor U19835 (N_19835,N_16632,N_17001);
and U19836 (N_19836,N_15657,N_16513);
nor U19837 (N_19837,N_16704,N_16994);
and U19838 (N_19838,N_15466,N_15984);
nand U19839 (N_19839,N_17499,N_16298);
xnor U19840 (N_19840,N_16427,N_17443);
xnor U19841 (N_19841,N_17390,N_15932);
nand U19842 (N_19842,N_15342,N_15006);
and U19843 (N_19843,N_15482,N_16438);
or U19844 (N_19844,N_16189,N_15453);
xnor U19845 (N_19845,N_16678,N_16106);
xnor U19846 (N_19846,N_15683,N_15337);
xnor U19847 (N_19847,N_15707,N_15666);
xor U19848 (N_19848,N_15614,N_16811);
xnor U19849 (N_19849,N_17377,N_17181);
nand U19850 (N_19850,N_16241,N_15911);
or U19851 (N_19851,N_15008,N_16526);
nor U19852 (N_19852,N_15476,N_17444);
and U19853 (N_19853,N_16836,N_16657);
nand U19854 (N_19854,N_16405,N_15183);
nand U19855 (N_19855,N_15309,N_15674);
nand U19856 (N_19856,N_15934,N_15461);
xor U19857 (N_19857,N_16487,N_15987);
or U19858 (N_19858,N_15182,N_17050);
or U19859 (N_19859,N_15917,N_15552);
nand U19860 (N_19860,N_17296,N_17003);
and U19861 (N_19861,N_17082,N_17443);
xnor U19862 (N_19862,N_17458,N_15656);
nand U19863 (N_19863,N_16844,N_16973);
xor U19864 (N_19864,N_16426,N_15831);
and U19865 (N_19865,N_16716,N_15068);
or U19866 (N_19866,N_17388,N_16954);
nor U19867 (N_19867,N_16310,N_16796);
nor U19868 (N_19868,N_17490,N_17374);
or U19869 (N_19869,N_15493,N_15353);
nor U19870 (N_19870,N_15965,N_15260);
nand U19871 (N_19871,N_16541,N_17040);
nor U19872 (N_19872,N_17164,N_15574);
and U19873 (N_19873,N_17053,N_16856);
or U19874 (N_19874,N_15264,N_17266);
xor U19875 (N_19875,N_15498,N_15044);
nor U19876 (N_19876,N_16771,N_17079);
and U19877 (N_19877,N_17290,N_17423);
nand U19878 (N_19878,N_16912,N_16891);
and U19879 (N_19879,N_16876,N_15140);
nand U19880 (N_19880,N_15335,N_16696);
xor U19881 (N_19881,N_15020,N_16133);
xor U19882 (N_19882,N_16585,N_16035);
or U19883 (N_19883,N_15769,N_16042);
xor U19884 (N_19884,N_16723,N_17466);
nand U19885 (N_19885,N_16858,N_16390);
xor U19886 (N_19886,N_16774,N_17466);
nor U19887 (N_19887,N_17081,N_16014);
xnor U19888 (N_19888,N_17368,N_15178);
and U19889 (N_19889,N_16987,N_17298);
nor U19890 (N_19890,N_16059,N_17381);
or U19891 (N_19891,N_16197,N_15706);
nand U19892 (N_19892,N_15234,N_16318);
nor U19893 (N_19893,N_15930,N_16748);
nor U19894 (N_19894,N_17352,N_17483);
or U19895 (N_19895,N_15258,N_16800);
or U19896 (N_19896,N_16155,N_16631);
and U19897 (N_19897,N_17130,N_15708);
or U19898 (N_19898,N_16764,N_16677);
xor U19899 (N_19899,N_16016,N_15532);
nand U19900 (N_19900,N_15653,N_15144);
and U19901 (N_19901,N_15349,N_15247);
xnor U19902 (N_19902,N_15679,N_16732);
nor U19903 (N_19903,N_16977,N_16012);
or U19904 (N_19904,N_16185,N_15164);
or U19905 (N_19905,N_17333,N_16150);
nand U19906 (N_19906,N_16342,N_16565);
or U19907 (N_19907,N_16061,N_16847);
nand U19908 (N_19908,N_16461,N_17344);
xor U19909 (N_19909,N_15051,N_16017);
and U19910 (N_19910,N_16001,N_15116);
nand U19911 (N_19911,N_16953,N_17340);
nor U19912 (N_19912,N_16604,N_17461);
xor U19913 (N_19913,N_17498,N_15734);
xnor U19914 (N_19914,N_16850,N_15279);
nand U19915 (N_19915,N_16625,N_15669);
nor U19916 (N_19916,N_15150,N_16741);
nand U19917 (N_19917,N_15332,N_15091);
nand U19918 (N_19918,N_15937,N_17001);
nor U19919 (N_19919,N_17168,N_16298);
or U19920 (N_19920,N_17362,N_15122);
and U19921 (N_19921,N_17464,N_16209);
or U19922 (N_19922,N_16603,N_17156);
nand U19923 (N_19923,N_17395,N_15263);
nand U19924 (N_19924,N_15850,N_15539);
or U19925 (N_19925,N_16564,N_17184);
nor U19926 (N_19926,N_16280,N_15626);
nor U19927 (N_19927,N_17395,N_17236);
nor U19928 (N_19928,N_17393,N_15981);
xnor U19929 (N_19929,N_17084,N_16051);
and U19930 (N_19930,N_16213,N_16184);
nor U19931 (N_19931,N_17260,N_15335);
or U19932 (N_19932,N_15022,N_16943);
and U19933 (N_19933,N_15352,N_17121);
and U19934 (N_19934,N_16559,N_15685);
or U19935 (N_19935,N_15440,N_16117);
xnor U19936 (N_19936,N_17060,N_15073);
xor U19937 (N_19937,N_16818,N_15935);
nor U19938 (N_19938,N_16274,N_16366);
xor U19939 (N_19939,N_15082,N_15564);
xnor U19940 (N_19940,N_17293,N_15378);
and U19941 (N_19941,N_15170,N_17482);
and U19942 (N_19942,N_16491,N_15948);
and U19943 (N_19943,N_15939,N_16401);
or U19944 (N_19944,N_16470,N_16068);
or U19945 (N_19945,N_15036,N_16937);
nand U19946 (N_19946,N_15950,N_15304);
or U19947 (N_19947,N_17055,N_15406);
nand U19948 (N_19948,N_15571,N_16908);
nand U19949 (N_19949,N_16578,N_15112);
and U19950 (N_19950,N_15282,N_15352);
xor U19951 (N_19951,N_16654,N_16182);
xnor U19952 (N_19952,N_16239,N_15435);
and U19953 (N_19953,N_16312,N_17400);
or U19954 (N_19954,N_15684,N_16526);
xnor U19955 (N_19955,N_17097,N_15761);
nand U19956 (N_19956,N_15164,N_15697);
nor U19957 (N_19957,N_16458,N_15618);
xor U19958 (N_19958,N_17428,N_16814);
or U19959 (N_19959,N_15204,N_15784);
nand U19960 (N_19960,N_17295,N_16718);
and U19961 (N_19961,N_15288,N_16883);
and U19962 (N_19962,N_15771,N_15238);
nand U19963 (N_19963,N_16760,N_15977);
nand U19964 (N_19964,N_16088,N_15840);
nand U19965 (N_19965,N_15423,N_15204);
and U19966 (N_19966,N_15081,N_17205);
nor U19967 (N_19967,N_16208,N_16980);
nor U19968 (N_19968,N_15708,N_17321);
nor U19969 (N_19969,N_16590,N_15728);
nor U19970 (N_19970,N_17183,N_15877);
and U19971 (N_19971,N_16820,N_16640);
xnor U19972 (N_19972,N_17474,N_16686);
xor U19973 (N_19973,N_15499,N_15062);
and U19974 (N_19974,N_15346,N_16799);
nand U19975 (N_19975,N_16683,N_17228);
or U19976 (N_19976,N_16314,N_17361);
or U19977 (N_19977,N_16565,N_17493);
and U19978 (N_19978,N_15267,N_15498);
nor U19979 (N_19979,N_15540,N_15115);
or U19980 (N_19980,N_15449,N_16442);
nand U19981 (N_19981,N_16520,N_16264);
xnor U19982 (N_19982,N_16747,N_16920);
nand U19983 (N_19983,N_15416,N_16807);
and U19984 (N_19984,N_15428,N_15918);
xnor U19985 (N_19985,N_15798,N_16580);
or U19986 (N_19986,N_15376,N_16470);
nand U19987 (N_19987,N_15454,N_17256);
nand U19988 (N_19988,N_16652,N_16053);
nor U19989 (N_19989,N_16187,N_16472);
and U19990 (N_19990,N_16601,N_16638);
and U19991 (N_19991,N_17028,N_17312);
nor U19992 (N_19992,N_15724,N_15811);
nor U19993 (N_19993,N_15349,N_16698);
nand U19994 (N_19994,N_16700,N_16378);
xor U19995 (N_19995,N_16665,N_15668);
nor U19996 (N_19996,N_15461,N_16289);
nor U19997 (N_19997,N_15723,N_16283);
nor U19998 (N_19998,N_16059,N_15633);
nor U19999 (N_19999,N_17377,N_15344);
nor U20000 (N_20000,N_18719,N_18547);
nor U20001 (N_20001,N_18030,N_18854);
and U20002 (N_20002,N_17508,N_17768);
or U20003 (N_20003,N_19201,N_19118);
nor U20004 (N_20004,N_18818,N_19701);
and U20005 (N_20005,N_17570,N_19522);
nand U20006 (N_20006,N_18243,N_18885);
xor U20007 (N_20007,N_19133,N_18904);
or U20008 (N_20008,N_19098,N_17568);
xor U20009 (N_20009,N_19682,N_19848);
nand U20010 (N_20010,N_19899,N_17533);
xnor U20011 (N_20011,N_17879,N_17591);
or U20012 (N_20012,N_19725,N_18503);
or U20013 (N_20013,N_19526,N_19251);
and U20014 (N_20014,N_18008,N_18023);
and U20015 (N_20015,N_18408,N_18632);
or U20016 (N_20016,N_18371,N_19813);
xnor U20017 (N_20017,N_19002,N_18938);
nor U20018 (N_20018,N_19864,N_18360);
nand U20019 (N_20019,N_17601,N_19886);
nand U20020 (N_20020,N_19503,N_18742);
nor U20021 (N_20021,N_17620,N_19929);
xnor U20022 (N_20022,N_19532,N_19377);
nand U20023 (N_20023,N_19043,N_19507);
and U20024 (N_20024,N_19825,N_19148);
or U20025 (N_20025,N_19122,N_19268);
nor U20026 (N_20026,N_19070,N_18186);
nand U20027 (N_20027,N_18588,N_19850);
and U20028 (N_20028,N_18354,N_19315);
and U20029 (N_20029,N_18064,N_19077);
nor U20030 (N_20030,N_18836,N_19069);
nor U20031 (N_20031,N_17559,N_17563);
nor U20032 (N_20032,N_19390,N_19476);
and U20033 (N_20033,N_19036,N_19175);
and U20034 (N_20034,N_19634,N_18110);
and U20035 (N_20035,N_18123,N_18219);
nand U20036 (N_20036,N_18473,N_18669);
nor U20037 (N_20037,N_18966,N_18456);
xor U20038 (N_20038,N_17608,N_19966);
xor U20039 (N_20039,N_17839,N_19796);
xor U20040 (N_20040,N_19294,N_17866);
or U20041 (N_20041,N_19677,N_18848);
nand U20042 (N_20042,N_19557,N_17875);
xnor U20043 (N_20043,N_19244,N_18878);
nand U20044 (N_20044,N_18239,N_18006);
or U20045 (N_20045,N_18301,N_17564);
xor U20046 (N_20046,N_18240,N_19967);
xnor U20047 (N_20047,N_18271,N_17847);
or U20048 (N_20048,N_19593,N_18931);
or U20049 (N_20049,N_18325,N_19012);
xor U20050 (N_20050,N_19344,N_18055);
nor U20051 (N_20051,N_17710,N_17724);
nand U20052 (N_20052,N_18537,N_19766);
nor U20053 (N_20053,N_19424,N_19099);
nand U20054 (N_20054,N_17702,N_19924);
nor U20055 (N_20055,N_18142,N_17773);
or U20056 (N_20056,N_19194,N_17515);
xnor U20057 (N_20057,N_17987,N_19328);
or U20058 (N_20058,N_19159,N_18415);
nor U20059 (N_20059,N_19697,N_19604);
xnor U20060 (N_20060,N_19569,N_18351);
or U20061 (N_20061,N_17814,N_19025);
or U20062 (N_20062,N_17876,N_17948);
nand U20063 (N_20063,N_18617,N_17506);
or U20064 (N_20064,N_18831,N_17838);
xor U20065 (N_20065,N_19490,N_17593);
nand U20066 (N_20066,N_19680,N_18631);
and U20067 (N_20067,N_18377,N_19773);
nor U20068 (N_20068,N_18201,N_17906);
or U20069 (N_20069,N_18627,N_18167);
or U20070 (N_20070,N_19576,N_17534);
and U20071 (N_20071,N_19094,N_17926);
nand U20072 (N_20072,N_17758,N_18734);
nor U20073 (N_20073,N_18144,N_19510);
xor U20074 (N_20074,N_19664,N_17654);
nand U20075 (N_20075,N_19814,N_17784);
xnor U20076 (N_20076,N_17981,N_18444);
xnor U20077 (N_20077,N_17889,N_19193);
nor U20078 (N_20078,N_19411,N_19910);
or U20079 (N_20079,N_18450,N_19897);
or U20080 (N_20080,N_17578,N_19992);
nor U20081 (N_20081,N_17994,N_19700);
and U20082 (N_20082,N_19947,N_17543);
or U20083 (N_20083,N_18881,N_18375);
nor U20084 (N_20084,N_18768,N_19064);
or U20085 (N_20085,N_18474,N_18180);
xnor U20086 (N_20086,N_18838,N_17785);
and U20087 (N_20087,N_19902,N_19749);
or U20088 (N_20088,N_18879,N_18993);
or U20089 (N_20089,N_18391,N_18257);
or U20090 (N_20090,N_18772,N_19414);
xor U20091 (N_20091,N_19457,N_18769);
xnor U20092 (N_20092,N_17940,N_19284);
xnor U20093 (N_20093,N_17852,N_19347);
nor U20094 (N_20094,N_18693,N_18963);
or U20095 (N_20095,N_19354,N_18807);
nor U20096 (N_20096,N_17565,N_18234);
or U20097 (N_20097,N_17792,N_18428);
xnor U20098 (N_20098,N_19731,N_17943);
and U20099 (N_20099,N_18715,N_19780);
or U20100 (N_20100,N_19953,N_17918);
or U20101 (N_20101,N_19330,N_19331);
nor U20102 (N_20102,N_19007,N_19809);
or U20103 (N_20103,N_18821,N_19208);
nor U20104 (N_20104,N_18113,N_19633);
xor U20105 (N_20105,N_18935,N_18595);
nor U20106 (N_20106,N_18461,N_19101);
and U20107 (N_20107,N_18906,N_18107);
nand U20108 (N_20108,N_17603,N_19919);
nor U20109 (N_20109,N_17984,N_18267);
or U20110 (N_20110,N_19401,N_18546);
nand U20111 (N_20111,N_19446,N_19391);
nor U20112 (N_20112,N_19247,N_17642);
and U20113 (N_20113,N_19811,N_19669);
and U20114 (N_20114,N_18153,N_17811);
or U20115 (N_20115,N_19250,N_18798);
and U20116 (N_20116,N_17989,N_18463);
xnor U20117 (N_20117,N_19686,N_18216);
nand U20118 (N_20118,N_19514,N_19092);
nand U20119 (N_20119,N_18773,N_19292);
nand U20120 (N_20120,N_19191,N_18573);
xor U20121 (N_20121,N_19371,N_18388);
nand U20122 (N_20122,N_19548,N_18514);
nor U20123 (N_20123,N_18973,N_18845);
or U20124 (N_20124,N_18764,N_19234);
or U20125 (N_20125,N_17698,N_19581);
xor U20126 (N_20126,N_17867,N_18579);
or U20127 (N_20127,N_18012,N_19260);
nand U20128 (N_20128,N_18814,N_19640);
xor U20129 (N_20129,N_18407,N_19676);
and U20130 (N_20130,N_18007,N_19478);
nor U20131 (N_20131,N_18921,N_18675);
nor U20132 (N_20132,N_19829,N_18732);
and U20133 (N_20133,N_19795,N_18914);
xnor U20134 (N_20134,N_17854,N_18355);
or U20135 (N_20135,N_19129,N_18756);
nand U20136 (N_20136,N_18792,N_19135);
nand U20137 (N_20137,N_17697,N_18698);
xnor U20138 (N_20138,N_17979,N_18810);
nor U20139 (N_20139,N_18972,N_18908);
and U20140 (N_20140,N_17677,N_18762);
and U20141 (N_20141,N_19198,N_18259);
xnor U20142 (N_20142,N_18531,N_19710);
nor U20143 (N_20143,N_18997,N_19000);
nand U20144 (N_20144,N_17976,N_19555);
nor U20145 (N_20145,N_18600,N_17502);
and U20146 (N_20146,N_17978,N_19951);
and U20147 (N_20147,N_18302,N_17527);
or U20148 (N_20148,N_19982,N_19365);
or U20149 (N_20149,N_19463,N_19277);
nor U20150 (N_20150,N_19210,N_19496);
or U20151 (N_20151,N_18849,N_18034);
nor U20152 (N_20152,N_18620,N_18712);
or U20153 (N_20153,N_19560,N_18598);
nand U20154 (N_20154,N_17993,N_18690);
nand U20155 (N_20155,N_19591,N_19415);
xnor U20156 (N_20156,N_17621,N_19104);
and U20157 (N_20157,N_17835,N_17997);
xnor U20158 (N_20158,N_19888,N_18862);
nand U20159 (N_20159,N_19273,N_18209);
or U20160 (N_20160,N_18104,N_19097);
nor U20161 (N_20161,N_18535,N_19574);
or U20162 (N_20162,N_19934,N_19061);
nand U20163 (N_20163,N_17645,N_19649);
nor U20164 (N_20164,N_17592,N_19038);
nor U20165 (N_20165,N_19372,N_17911);
and U20166 (N_20166,N_18562,N_17575);
and U20167 (N_20167,N_19004,N_19040);
and U20168 (N_20168,N_18475,N_18074);
nor U20169 (N_20169,N_17942,N_19616);
or U20170 (N_20170,N_18635,N_18552);
or U20171 (N_20171,N_17514,N_18046);
or U20172 (N_20172,N_19985,N_18129);
nor U20173 (N_20173,N_17661,N_18379);
and U20174 (N_20174,N_19163,N_18888);
nand U20175 (N_20175,N_19445,N_19475);
nand U20176 (N_20176,N_18221,N_17830);
nor U20177 (N_20177,N_17795,N_18961);
nand U20178 (N_20178,N_19747,N_17779);
nor U20179 (N_20179,N_19971,N_19596);
xor U20180 (N_20180,N_19461,N_17500);
xor U20181 (N_20181,N_19804,N_17572);
xor U20182 (N_20182,N_19483,N_18057);
xnor U20183 (N_20183,N_19826,N_19263);
or U20184 (N_20184,N_18718,N_17726);
nor U20185 (N_20185,N_18198,N_18442);
and U20186 (N_20186,N_18670,N_19779);
and U20187 (N_20187,N_19525,N_17812);
and U20188 (N_20188,N_17837,N_19754);
nor U20189 (N_20189,N_18398,N_18062);
nor U20190 (N_20190,N_17713,N_18532);
or U20191 (N_20191,N_18162,N_17536);
or U20192 (N_20192,N_19736,N_19805);
nor U20193 (N_20193,N_18707,N_19958);
nand U20194 (N_20194,N_19918,N_19889);
and U20195 (N_20195,N_17870,N_19536);
and U20196 (N_20196,N_19110,N_18913);
nand U20197 (N_20197,N_19931,N_19699);
and U20198 (N_20198,N_19236,N_19681);
nor U20199 (N_20199,N_18636,N_19545);
or U20200 (N_20200,N_19213,N_18197);
and U20201 (N_20201,N_18946,N_17655);
nor U20202 (N_20202,N_18919,N_17715);
xor U20203 (N_20203,N_18068,N_18472);
or U20204 (N_20204,N_19540,N_18823);
nand U20205 (N_20205,N_17672,N_17694);
or U20206 (N_20206,N_18847,N_18050);
or U20207 (N_20207,N_19241,N_17902);
nor U20208 (N_20208,N_18362,N_19741);
xnor U20209 (N_20209,N_18136,N_18053);
nor U20210 (N_20210,N_17922,N_17759);
and U20211 (N_20211,N_17958,N_17826);
nand U20212 (N_20212,N_18655,N_18190);
and U20213 (N_20213,N_18643,N_17874);
xnor U20214 (N_20214,N_19647,N_19382);
or U20215 (N_20215,N_19824,N_19403);
nor U20216 (N_20216,N_18920,N_19949);
nand U20217 (N_20217,N_18549,N_18273);
xor U20218 (N_20218,N_19182,N_18395);
nor U20219 (N_20219,N_17813,N_19619);
or U20220 (N_20220,N_18811,N_18322);
nor U20221 (N_20221,N_19717,N_19753);
and U20222 (N_20222,N_17951,N_19821);
nor U20223 (N_20223,N_19146,N_19229);
and U20224 (N_20224,N_19047,N_18610);
or U20225 (N_20225,N_18424,N_18329);
and U20226 (N_20226,N_18895,N_18576);
nor U20227 (N_20227,N_18833,N_17703);
xor U20228 (N_20228,N_18029,N_19014);
nand U20229 (N_20229,N_19041,N_18173);
or U20230 (N_20230,N_17797,N_19960);
or U20231 (N_20231,N_19885,N_19205);
nand U20232 (N_20232,N_19959,N_18916);
and U20233 (N_20233,N_19552,N_19565);
or U20234 (N_20234,N_18366,N_18599);
xor U20235 (N_20235,N_19995,N_17615);
nor U20236 (N_20236,N_18800,N_18000);
nor U20237 (N_20237,N_18460,N_19480);
nand U20238 (N_20238,N_17845,N_19602);
and U20239 (N_20239,N_17964,N_19626);
xnor U20240 (N_20240,N_18128,N_18336);
xnor U20241 (N_20241,N_19610,N_19079);
nor U20242 (N_20242,N_18897,N_18349);
nand U20243 (N_20243,N_18727,N_19879);
or U20244 (N_20244,N_19857,N_17913);
nor U20245 (N_20245,N_19538,N_17765);
xor U20246 (N_20246,N_19563,N_18410);
xnor U20247 (N_20247,N_18297,N_19878);
nor U20248 (N_20248,N_17821,N_19876);
and U20249 (N_20249,N_19262,N_19454);
or U20250 (N_20250,N_18251,N_18891);
nor U20251 (N_20251,N_18134,N_17819);
xor U20252 (N_20252,N_19769,N_19368);
and U20253 (N_20253,N_18928,N_17684);
and U20254 (N_20254,N_18527,N_19109);
or U20255 (N_20255,N_18135,N_19989);
and U20256 (N_20256,N_17895,N_18303);
nand U20257 (N_20257,N_18193,N_18509);
nor U20258 (N_20258,N_18312,N_19239);
or U20259 (N_20259,N_18352,N_19645);
nand U20260 (N_20260,N_19008,N_18130);
nand U20261 (N_20261,N_19635,N_17587);
xor U20262 (N_20262,N_18277,N_19030);
xor U20263 (N_20263,N_19996,N_18274);
and U20264 (N_20264,N_17971,N_18445);
xnor U20265 (N_20265,N_18261,N_18014);
xnor U20266 (N_20266,N_18641,N_17598);
and U20267 (N_20267,N_19997,N_17573);
nand U20268 (N_20268,N_18479,N_19499);
and U20269 (N_20269,N_18944,N_18393);
and U20270 (N_20270,N_18044,N_18356);
or U20271 (N_20271,N_19531,N_18939);
xor U20272 (N_20272,N_17541,N_18105);
nor U20273 (N_20273,N_18866,N_19594);
nand U20274 (N_20274,N_19685,N_17516);
nand U20275 (N_20275,N_18634,N_19527);
xor U20276 (N_20276,N_17518,N_19866);
and U20277 (N_20277,N_17720,N_19867);
nor U20278 (N_20278,N_18047,N_19102);
nor U20279 (N_20279,N_19224,N_19636);
and U20280 (N_20280,N_17966,N_18604);
nor U20281 (N_20281,N_18868,N_19196);
xor U20282 (N_20282,N_18174,N_17968);
or U20283 (N_20283,N_18924,N_18813);
or U20284 (N_20284,N_18587,N_19801);
and U20285 (N_20285,N_19246,N_19984);
nor U20286 (N_20286,N_17531,N_18500);
nor U20287 (N_20287,N_18411,N_17687);
nor U20288 (N_20288,N_18668,N_19612);
or U20289 (N_20289,N_19827,N_19764);
nor U20290 (N_20290,N_18860,N_19045);
and U20291 (N_20291,N_17557,N_19788);
or U20292 (N_20292,N_19906,N_19187);
nor U20293 (N_20293,N_18640,N_19440);
xnor U20294 (N_20294,N_18704,N_17962);
or U20295 (N_20295,N_17562,N_19991);
or U20296 (N_20296,N_19189,N_19974);
nand U20297 (N_20297,N_19618,N_18199);
nand U20298 (N_20298,N_17663,N_18822);
xor U20299 (N_20299,N_17682,N_19154);
nand U20300 (N_20300,N_19617,N_18563);
xor U20301 (N_20301,N_19761,N_18625);
and U20302 (N_20302,N_17817,N_18466);
nand U20303 (N_20303,N_18231,N_18292);
nand U20304 (N_20304,N_18373,N_17673);
nor U20305 (N_20305,N_19571,N_18037);
and U20306 (N_20306,N_18540,N_19721);
xnor U20307 (N_20307,N_19477,N_18841);
and U20308 (N_20308,N_19376,N_17800);
and U20309 (N_20309,N_17719,N_18208);
xor U20310 (N_20310,N_18593,N_18035);
nand U20311 (N_20311,N_17772,N_19726);
xnor U20312 (N_20312,N_18580,N_18100);
or U20313 (N_20313,N_18941,N_17907);
or U20314 (N_20314,N_19957,N_18121);
or U20315 (N_20315,N_19310,N_19508);
nor U20316 (N_20316,N_18059,N_18320);
xnor U20317 (N_20317,N_18247,N_18323);
or U20318 (N_20318,N_17947,N_18770);
nor U20319 (N_20319,N_18217,N_18179);
nand U20320 (N_20320,N_18476,N_19511);
nand U20321 (N_20321,N_19184,N_18969);
nor U20322 (N_20322,N_19279,N_19111);
xnor U20323 (N_20323,N_19925,N_18067);
nor U20324 (N_20324,N_18898,N_18150);
and U20325 (N_20325,N_19880,N_19080);
xor U20326 (N_20326,N_18926,N_19816);
and U20327 (N_20327,N_18999,N_17883);
and U20328 (N_20328,N_18882,N_18390);
nand U20329 (N_20329,N_18052,N_19369);
xor U20330 (N_20330,N_18027,N_18279);
nor U20331 (N_20331,N_19871,N_17632);
and U20332 (N_20332,N_19218,N_18656);
xnor U20333 (N_20333,N_18975,N_18950);
nor U20334 (N_20334,N_18629,N_18771);
or U20335 (N_20335,N_17535,N_18559);
and U20336 (N_20336,N_19751,N_19068);
or U20337 (N_20337,N_18075,N_19358);
and U20338 (N_20338,N_19443,N_19287);
nand U20339 (N_20339,N_18872,N_18419);
nand U20340 (N_20340,N_19689,N_17748);
and U20341 (N_20341,N_18212,N_19684);
nand U20342 (N_20342,N_19978,N_17511);
and U20343 (N_20343,N_18420,N_17877);
or U20344 (N_20344,N_17594,N_18066);
nor U20345 (N_20345,N_18706,N_19137);
nor U20346 (N_20346,N_17658,N_18747);
and U20347 (N_20347,N_18242,N_18143);
nor U20348 (N_20348,N_18940,N_18948);
or U20349 (N_20349,N_19907,N_18233);
or U20350 (N_20350,N_19656,N_19426);
and U20351 (N_20351,N_18671,N_17991);
xnor U20352 (N_20352,N_19870,N_18076);
nand U20353 (N_20353,N_18571,N_19032);
nor U20354 (N_20354,N_18910,N_17676);
and U20355 (N_20355,N_18026,N_19474);
or U20356 (N_20356,N_18272,N_19072);
nand U20357 (N_20357,N_19348,N_19715);
or U20358 (N_20358,N_19679,N_19733);
nor U20359 (N_20359,N_19537,N_17609);
xnor U20360 (N_20360,N_19486,N_18477);
nand U20361 (N_20361,N_19627,N_17639);
nor U20362 (N_20362,N_19550,N_19453);
xor U20363 (N_20363,N_18763,N_17542);
nor U20364 (N_20364,N_18761,N_18427);
or U20365 (N_20365,N_19011,N_19089);
and U20366 (N_20366,N_17977,N_17600);
nand U20367 (N_20367,N_18799,N_18048);
or U20368 (N_20368,N_17745,N_18021);
nand U20369 (N_20369,N_19759,N_17999);
nor U20370 (N_20370,N_19297,N_17912);
or U20371 (N_20371,N_17622,N_19868);
nand U20372 (N_20372,N_19441,N_19784);
and U20373 (N_20373,N_18077,N_18894);
xor U20374 (N_20374,N_18266,N_19350);
or U20375 (N_20375,N_18953,N_18146);
and U20376 (N_20376,N_17569,N_17766);
or U20377 (N_20377,N_17771,N_18353);
or U20378 (N_20378,N_18019,N_19623);
nand U20379 (N_20379,N_18225,N_19559);
and U20380 (N_20380,N_19143,N_18803);
nor U20381 (N_20381,N_18850,N_18268);
and U20382 (N_20382,N_19026,N_19956);
or U20383 (N_20383,N_19854,N_18650);
nor U20384 (N_20384,N_17714,N_19006);
or U20385 (N_20385,N_18314,N_18499);
and U20386 (N_20386,N_19057,N_19506);
nor U20387 (N_20387,N_17865,N_19981);
and U20388 (N_20388,N_18839,N_19497);
nand U20389 (N_20389,N_18909,N_17789);
and U20390 (N_20390,N_17853,N_17956);
or U20391 (N_20391,N_19892,N_18396);
nand U20392 (N_20392,N_18929,N_18736);
or U20393 (N_20393,N_18932,N_19858);
or U20394 (N_20394,N_17747,N_19972);
or U20395 (N_20395,N_19245,N_18663);
and U20396 (N_20396,N_19615,N_17864);
and U20397 (N_20397,N_18607,N_18339);
nor U20398 (N_20398,N_17732,N_19819);
nand U20399 (N_20399,N_17783,N_18725);
xnor U20400 (N_20400,N_18346,N_19657);
nand U20401 (N_20401,N_17679,N_19065);
nand U20402 (N_20402,N_19039,N_19639);
xor U20403 (N_20403,N_18181,N_19933);
nor U20404 (N_20404,N_19975,N_17613);
xnor U20405 (N_20405,N_18729,N_19893);
xor U20406 (N_20406,N_18613,N_18166);
nor U20407 (N_20407,N_19744,N_19822);
or U20408 (N_20408,N_17945,N_19459);
nand U20409 (N_20409,N_18206,N_19087);
or U20410 (N_20410,N_19509,N_17588);
nor U20411 (N_20411,N_18102,N_19523);
nor U20412 (N_20412,N_18967,N_18542);
nor U20413 (N_20413,N_19394,N_18204);
and U20414 (N_20414,N_19249,N_17923);
nand U20415 (N_20415,N_18258,N_19692);
and U20416 (N_20416,N_18172,N_19573);
nand U20417 (N_20417,N_19123,N_18705);
xnor U20418 (N_20418,N_17558,N_18072);
or U20419 (N_20419,N_19387,N_18287);
xnor U20420 (N_20420,N_19712,N_19781);
and U20421 (N_20421,N_17775,N_18551);
nand U20422 (N_20422,N_18001,N_18115);
nand U20423 (N_20423,N_18911,N_18890);
xnor U20424 (N_20424,N_17844,N_18334);
nor U20425 (N_20425,N_19223,N_17651);
xnor U20426 (N_20426,N_18344,N_19530);
and U20427 (N_20427,N_19028,N_19071);
and U20428 (N_20428,N_19739,N_19803);
or U20429 (N_20429,N_19314,N_19683);
nor U20430 (N_20430,N_19388,N_19607);
and U20431 (N_20431,N_17802,N_18844);
or U20432 (N_20432,N_19861,N_19316);
nor U20433 (N_20433,N_18673,N_18589);
xnor U20434 (N_20434,N_18099,N_18917);
nand U20435 (N_20435,N_18383,N_18369);
or U20436 (N_20436,N_18748,N_17547);
nand U20437 (N_20437,N_19939,N_18545);
nor U20438 (N_20438,N_19547,N_18554);
xor U20439 (N_20439,N_19333,N_19504);
or U20440 (N_20440,N_18679,N_17794);
nor U20441 (N_20441,N_18449,N_17635);
xnor U20442 (N_20442,N_17842,N_17707);
nand U20443 (N_20443,N_18887,N_19326);
nand U20444 (N_20444,N_19702,N_18943);
nand U20445 (N_20445,N_19730,N_19887);
or U20446 (N_20446,N_19666,N_18095);
or U20447 (N_20447,N_18745,N_18223);
xnor U20448 (N_20448,N_18350,N_18686);
nor U20449 (N_20449,N_19663,N_19752);
or U20450 (N_20450,N_17970,N_18677);
nand U20451 (N_20451,N_17705,N_19017);
xnor U20452 (N_20452,N_18794,N_17728);
nor U20453 (N_20453,N_19301,N_19772);
nand U20454 (N_20454,N_19471,N_18009);
and U20455 (N_20455,N_17696,N_18505);
or U20456 (N_20456,N_18086,N_18318);
nor U20457 (N_20457,N_17920,N_19209);
nor U20458 (N_20458,N_19737,N_18653);
nor U20459 (N_20459,N_17888,N_18731);
or U20460 (N_20460,N_19820,N_19131);
or U20461 (N_20461,N_19589,N_19756);
nand U20462 (N_20462,N_18131,N_18605);
nor U20463 (N_20463,N_19240,N_18126);
nand U20464 (N_20464,N_18577,N_19812);
or U20465 (N_20465,N_18585,N_18294);
nand U20466 (N_20466,N_18092,N_19265);
xnor U20467 (N_20467,N_19668,N_19711);
nor U20468 (N_20468,N_18033,N_19170);
nor U20469 (N_20469,N_18192,N_19542);
nand U20470 (N_20470,N_18722,N_17823);
nor U20471 (N_20471,N_17688,N_18714);
or U20472 (N_20472,N_19300,N_18912);
or U20473 (N_20473,N_18555,N_19115);
xor U20474 (N_20474,N_18687,N_19944);
and U20475 (N_20475,N_19716,N_19270);
nor U20476 (N_20476,N_17751,N_19705);
nand U20477 (N_20477,N_17756,N_19206);
xor U20478 (N_20478,N_17992,N_19383);
nand U20479 (N_20479,N_19621,N_17884);
nor U20480 (N_20480,N_19601,N_18169);
xnor U20481 (N_20481,N_17526,N_18430);
nor U20482 (N_20482,N_19895,N_18017);
and U20483 (N_20483,N_18536,N_19179);
and U20484 (N_20484,N_18776,N_17626);
and U20485 (N_20485,N_19317,N_19738);
nor U20486 (N_20486,N_18766,N_18439);
nand U20487 (N_20487,N_19998,N_19145);
nor U20488 (N_20488,N_18141,N_18157);
or U20489 (N_20489,N_19144,N_18827);
nand U20490 (N_20490,N_17725,N_18214);
nand U20491 (N_20491,N_19112,N_18084);
nand U20492 (N_20492,N_18544,N_17544);
xnor U20493 (N_20493,N_19577,N_19815);
and U20494 (N_20494,N_17933,N_18140);
or U20495 (N_20495,N_17924,N_17693);
or U20496 (N_20496,N_18020,N_17723);
nor U20497 (N_20497,N_18253,N_17549);
and U20498 (N_20498,N_17825,N_18815);
or U20499 (N_20499,N_18222,N_17625);
and U20500 (N_20500,N_18385,N_18802);
or U20501 (N_20501,N_19272,N_19053);
nand U20502 (N_20502,N_19418,N_18399);
xor U20503 (N_20503,N_19787,N_19655);
or U20504 (N_20504,N_19035,N_19379);
nor U20505 (N_20505,N_19535,N_19905);
nand U20506 (N_20506,N_18469,N_18662);
and U20507 (N_20507,N_18413,N_19049);
or U20508 (N_20508,N_19161,N_18070);
nand U20509 (N_20509,N_19654,N_17735);
nor U20510 (N_20510,N_17555,N_18743);
nand U20511 (N_20511,N_18959,N_19740);
or U20512 (N_20512,N_18730,N_18754);
and U20513 (N_20513,N_18628,N_17636);
xor U20514 (N_20514,N_18416,N_19786);
nor U20515 (N_20515,N_17574,N_18746);
nand U20516 (N_20516,N_19427,N_18936);
xnor U20517 (N_20517,N_19912,N_18382);
and U20518 (N_20518,N_19139,N_19168);
or U20519 (N_20519,N_18389,N_17736);
nor U20520 (N_20520,N_18484,N_17669);
and U20521 (N_20521,N_19999,N_18089);
nand U20522 (N_20522,N_18394,N_17937);
nand U20523 (N_20523,N_17931,N_19846);
or U20524 (N_20524,N_17827,N_19853);
nand U20525 (N_20525,N_19295,N_17681);
xnor U20526 (N_20526,N_18981,N_18965);
or U20527 (N_20527,N_19431,N_17885);
xor U20528 (N_20528,N_18575,N_19637);
xor U20529 (N_20529,N_19732,N_18678);
and U20530 (N_20530,N_18567,N_18359);
nor U20531 (N_20531,N_18093,N_17953);
xnor U20532 (N_20532,N_18147,N_19728);
nor U20533 (N_20533,N_19930,N_19843);
xnor U20534 (N_20534,N_18249,N_18659);
and U20535 (N_20535,N_17754,N_19782);
nand U20536 (N_20536,N_17529,N_19450);
nor U20537 (N_20537,N_19817,N_18111);
or U20538 (N_20538,N_18530,N_19067);
nand U20539 (N_20539,N_19495,N_17757);
nand U20540 (N_20540,N_19117,N_18406);
and U20541 (N_20541,N_17843,N_19405);
and U20542 (N_20542,N_19373,N_19632);
or U20543 (N_20543,N_18361,N_19052);
xnor U20544 (N_20544,N_18561,N_17892);
or U20545 (N_20545,N_18989,N_17871);
xor U20546 (N_20546,N_18338,N_18189);
xnor U20547 (N_20547,N_17585,N_19136);
or U20548 (N_20548,N_17510,N_19298);
nand U20549 (N_20549,N_19969,N_19422);
nor U20550 (N_20550,N_19015,N_18786);
and U20551 (N_20551,N_18202,N_19018);
nor U20552 (N_20552,N_17634,N_19338);
and U20553 (N_20553,N_19884,N_18623);
or U20554 (N_20554,N_18210,N_18820);
and U20555 (N_20555,N_19493,N_18649);
nor U20556 (N_20556,N_18293,N_18592);
nand U20557 (N_20557,N_18624,N_17583);
nand U20558 (N_20558,N_18572,N_18478);
nor U20559 (N_20559,N_18630,N_17898);
nor U20560 (N_20560,N_18875,N_19166);
nor U20561 (N_20561,N_19652,N_18720);
xnor U20562 (N_20562,N_19554,N_19033);
or U20563 (N_20563,N_19438,N_18363);
nor U20564 (N_20564,N_19927,N_18884);
and U20565 (N_20565,N_18837,N_17650);
nand U20566 (N_20566,N_19955,N_18288);
and U20567 (N_20567,N_18237,N_18342);
nand U20568 (N_20568,N_18452,N_17612);
and U20569 (N_20569,N_18982,N_18435);
xor U20570 (N_20570,N_19950,N_19675);
xnor U20571 (N_20571,N_18211,N_18482);
and U20572 (N_20572,N_18263,N_17597);
and U20573 (N_20573,N_17815,N_18995);
and U20574 (N_20574,N_19755,N_19190);
or U20575 (N_20575,N_18175,N_18645);
nor U20576 (N_20576,N_19124,N_17624);
nand U20577 (N_20577,N_18073,N_19257);
or U20578 (N_20578,N_19696,N_19976);
and U20579 (N_20579,N_18096,N_18283);
and U20580 (N_20580,N_18332,N_19777);
nand U20581 (N_20581,N_19259,N_18918);
nor U20582 (N_20582,N_19396,N_18782);
nor U20583 (N_20583,N_18949,N_18735);
nand U20584 (N_20584,N_18248,N_17887);
nand U20585 (N_20585,N_19983,N_18937);
and U20586 (N_20586,N_17869,N_18235);
nand U20587 (N_20587,N_18467,N_18945);
nand U20588 (N_20588,N_18250,N_19409);
or U20589 (N_20589,N_19221,N_18560);
xor U20590 (N_20590,N_18685,N_19192);
xor U20591 (N_20591,N_19802,N_17530);
nand U20592 (N_20592,N_18695,N_18905);
or U20593 (N_20593,N_17855,N_19237);
xor U20594 (N_20594,N_18457,N_19703);
xor U20595 (N_20595,N_17798,N_18638);
xor U20596 (N_20596,N_18780,N_19911);
nor U20597 (N_20597,N_18319,N_19521);
xnor U20598 (N_20598,N_18925,N_17910);
nor U20599 (N_20599,N_17777,N_18788);
nand U20600 (N_20600,N_17683,N_18816);
and U20601 (N_20601,N_19162,N_19862);
and U20602 (N_20602,N_17739,N_17896);
xnor U20603 (N_20603,N_19100,N_19707);
or U20604 (N_20604,N_17695,N_17501);
xor U20605 (N_20605,N_19408,N_19171);
or U20606 (N_20606,N_17939,N_18443);
nand U20607 (N_20607,N_17599,N_19729);
xnor U20608 (N_20608,N_18321,N_19869);
xor U20609 (N_20609,N_18767,N_17656);
xor U20610 (N_20610,N_18139,N_19211);
nor U20611 (N_20611,N_17610,N_19890);
and U20612 (N_20612,N_19380,N_18384);
xor U20613 (N_20613,N_18117,N_17517);
nand U20614 (N_20614,N_19570,N_18985);
nor U20615 (N_20615,N_17662,N_19688);
and U20616 (N_20616,N_19667,N_18958);
nor U20617 (N_20617,N_17946,N_19600);
nand U20618 (N_20618,N_17787,N_18819);
nand U20619 (N_20619,N_19389,N_18570);
and U20620 (N_20620,N_18244,N_18791);
and U20621 (N_20621,N_18521,N_18612);
and U20622 (N_20622,N_19466,N_18529);
and U20623 (N_20623,N_18608,N_19197);
xor U20624 (N_20624,N_19765,N_18124);
and U20625 (N_20625,N_17752,N_19151);
xnor U20626 (N_20626,N_19622,N_18696);
and U20627 (N_20627,N_18633,N_18843);
nand U20628 (N_20628,N_19055,N_18094);
xor U20629 (N_20629,N_17718,N_17589);
or U20630 (N_20630,N_18606,N_17909);
and U20631 (N_20631,N_18808,N_19852);
and U20632 (N_20632,N_18619,N_19834);
or U20633 (N_20633,N_18749,N_19519);
and U20634 (N_20634,N_18038,N_17988);
nor U20635 (N_20635,N_18665,N_18041);
xor U20636 (N_20636,N_17652,N_19095);
or U20637 (N_20637,N_18036,N_18282);
or U20638 (N_20638,N_19125,N_18358);
xor U20639 (N_20639,N_18063,N_19349);
or U20640 (N_20640,N_18345,N_17810);
nor U20641 (N_20641,N_19695,N_17633);
xnor U20642 (N_20642,N_18045,N_19127);
nor U20643 (N_20643,N_19325,N_19384);
xor U20644 (N_20644,N_19278,N_17602);
nand U20645 (N_20645,N_17881,N_19840);
nand U20646 (N_20646,N_19945,N_18737);
nand U20647 (N_20647,N_17522,N_17954);
or U20648 (N_20648,N_18137,N_17742);
and U20649 (N_20649,N_18299,N_18507);
and U20650 (N_20650,N_19074,N_18992);
xor U20651 (N_20651,N_19926,N_19152);
or U20652 (N_20652,N_19472,N_19516);
and U20653 (N_20653,N_19776,N_18723);
nand U20654 (N_20654,N_18942,N_19367);
xor U20655 (N_20655,N_19407,N_18459);
nor U20656 (N_20656,N_19743,N_17807);
nand U20657 (N_20657,N_18708,N_19505);
and U20658 (N_20658,N_17778,N_19215);
and U20659 (N_20659,N_19108,N_19212);
and U20660 (N_20660,N_19083,N_18412);
and U20661 (N_20661,N_19285,N_17846);
nor U20662 (N_20662,N_19051,N_19021);
nand U20663 (N_20663,N_18340,N_19990);
xnor U20664 (N_20664,N_19771,N_17919);
nor U20665 (N_20665,N_18646,N_19722);
nand U20666 (N_20666,N_18738,N_18777);
or U20667 (N_20667,N_18976,N_18703);
and U20668 (N_20668,N_19149,N_18994);
or U20669 (N_20669,N_19385,N_18489);
xor U20670 (N_20670,N_19044,N_18717);
or U20671 (N_20671,N_17699,N_19544);
xnor U20672 (N_20672,N_17561,N_19322);
or U20673 (N_20673,N_19855,N_18446);
and U20674 (N_20674,N_19009,N_18471);
xor U20675 (N_20675,N_18755,N_19882);
xor U20676 (N_20676,N_19793,N_18934);
nand U20677 (N_20677,N_19219,N_18069);
xor U20678 (N_20678,N_19416,N_17670);
and U20679 (N_20679,N_19288,N_19010);
nand U20680 (N_20680,N_19464,N_18852);
or U20681 (N_20681,N_18785,N_18182);
or U20682 (N_20682,N_18331,N_19873);
and U20683 (N_20683,N_17708,N_18740);
nor U20684 (N_20684,N_19091,N_18960);
nand U20685 (N_20685,N_19833,N_19818);
nand U20686 (N_20686,N_17540,N_17927);
xnor U20687 (N_20687,N_19770,N_19164);
nand U20688 (N_20688,N_19296,N_19528);
nand U20689 (N_20689,N_19558,N_19183);
xor U20690 (N_20690,N_19020,N_17969);
nand U20691 (N_20691,N_17796,N_18028);
or U20692 (N_20692,N_19120,N_17749);
and U20693 (N_20693,N_18951,N_19147);
nor U20694 (N_20694,N_17750,N_19948);
nand U20695 (N_20695,N_18991,N_18005);
nor U20696 (N_20696,N_18315,N_19468);
nor U20697 (N_20697,N_19562,N_17706);
xnor U20698 (N_20698,N_19381,N_17985);
nor U20699 (N_20699,N_19276,N_17665);
xor U20700 (N_20700,N_18490,N_18024);
and U20701 (N_20701,N_18541,N_19132);
xor U20702 (N_20702,N_17646,N_19849);
xor U20703 (N_20703,N_19492,N_18481);
nand U20704 (N_20704,N_19674,N_17727);
and U20705 (N_20705,N_17955,N_18016);
nand U20706 (N_20706,N_19181,N_19231);
nor U20707 (N_20707,N_17781,N_19877);
nor U20708 (N_20708,N_17886,N_18787);
and U20709 (N_20709,N_18744,N_17618);
nand U20710 (N_20710,N_17744,N_17936);
nand U20711 (N_20711,N_19502,N_19534);
and U20712 (N_20712,N_18486,N_18526);
and U20713 (N_20713,N_18138,N_19073);
or U20714 (N_20714,N_18455,N_17963);
and U20715 (N_20715,N_19746,N_18152);
xnor U20716 (N_20716,N_19106,N_19253);
and U20717 (N_20717,N_18098,N_19436);
and U20718 (N_20718,N_18970,N_18378);
nand U20719 (N_20719,N_17716,N_19375);
or U20720 (N_20720,N_19363,N_19023);
nor U20721 (N_20721,N_19435,N_18185);
nand U20722 (N_20722,N_18083,N_19321);
nand U20723 (N_20723,N_18590,N_19928);
nor U20724 (N_20724,N_19341,N_19393);
nor U20725 (N_20725,N_18402,N_19922);
nand U20726 (N_20726,N_18870,N_19332);
nand U20727 (N_20727,N_19397,N_19103);
xnor U20728 (N_20728,N_19644,N_19351);
xnor U20729 (N_20729,N_18664,N_19580);
or U20730 (N_20730,N_17973,N_17580);
xor U20731 (N_20731,N_19113,N_18236);
nor U20732 (N_20732,N_18156,N_18421);
nand U20733 (N_20733,N_17957,N_18877);
or U20734 (N_20734,N_19230,N_19698);
and U20735 (N_20735,N_17586,N_17809);
or U20736 (N_20736,N_19714,N_19258);
or U20737 (N_20737,N_18433,N_19767);
and U20738 (N_20738,N_19760,N_19823);
or U20739 (N_20739,N_17860,N_18516);
or U20740 (N_20740,N_19086,N_19360);
nor U20741 (N_20741,N_18495,N_18178);
and U20742 (N_20742,N_17507,N_18004);
nand U20743 (N_20743,N_17689,N_18191);
and U20744 (N_20744,N_19107,N_17614);
or U20745 (N_20745,N_18165,N_17512);
nor U20746 (N_20746,N_18978,N_18539);
and U20747 (N_20747,N_18654,N_17764);
and U20748 (N_20748,N_19603,N_18502);
nand U20749 (N_20749,N_19309,N_18876);
nand U20750 (N_20750,N_19458,N_17900);
or U20751 (N_20751,N_17824,N_17850);
nand U20752 (N_20752,N_19671,N_19592);
or U20753 (N_20753,N_18962,N_18122);
xnor U20754 (N_20754,N_18423,N_18700);
nor U20755 (N_20755,N_17753,N_18324);
nor U20756 (N_20756,N_18642,N_19606);
nor U20757 (N_20757,N_18434,N_17803);
nor U20758 (N_20758,N_18553,N_18688);
nor U20759 (N_20759,N_18611,N_18689);
nand U20760 (N_20760,N_19423,N_19800);
nor U20761 (N_20761,N_19177,N_19690);
and U20762 (N_20762,N_17607,N_19727);
and U20763 (N_20763,N_18618,N_18080);
and U20764 (N_20764,N_18429,N_17929);
nor U20765 (N_20765,N_17667,N_19952);
and U20766 (N_20766,N_19965,N_17638);
and U20767 (N_20767,N_19165,N_19831);
xnor U20768 (N_20768,N_19203,N_17643);
nor U20769 (N_20769,N_18296,N_18071);
nor U20770 (N_20770,N_18907,N_18869);
nand U20771 (N_20771,N_19410,N_17930);
and U20772 (N_20772,N_19595,N_19362);
nor U20773 (N_20773,N_19515,N_19398);
xnor U20774 (N_20774,N_18269,N_19546);
nand U20775 (N_20775,N_19587,N_19762);
nand U20776 (N_20776,N_18367,N_17721);
nor U20777 (N_20777,N_17982,N_18586);
and U20778 (N_20778,N_18512,N_19932);
nand U20779 (N_20779,N_19799,N_19847);
and U20780 (N_20780,N_18133,N_19141);
or U20781 (N_20781,N_19076,N_19353);
and U20782 (N_20782,N_19789,N_19859);
nor U20783 (N_20783,N_18859,N_17581);
or U20784 (N_20784,N_19228,N_17660);
nand U20785 (N_20785,N_19172,N_19643);
xnor U20786 (N_20786,N_18900,N_18177);
or U20787 (N_20787,N_18892,N_17686);
and U20788 (N_20788,N_18414,N_19386);
nor U20789 (N_20789,N_18765,N_18603);
and U20790 (N_20790,N_18284,N_18082);
nand U20791 (N_20791,N_19900,N_18468);
xnor U20792 (N_20792,N_17972,N_18155);
or U20793 (N_20793,N_19160,N_18583);
nand U20794 (N_20794,N_17576,N_19792);
or U20795 (N_20795,N_18508,N_19188);
xnor U20796 (N_20796,N_17709,N_18087);
and U20797 (N_20797,N_19318,N_19961);
nor U20798 (N_20798,N_17551,N_19027);
nor U20799 (N_20799,N_18255,N_19517);
or U20800 (N_20800,N_19693,N_19708);
or U20801 (N_20801,N_19226,N_19320);
or U20802 (N_20802,N_17790,N_18386);
and U20803 (N_20803,N_17915,N_18733);
and U20804 (N_20804,N_18840,N_18025);
nand U20805 (N_20805,N_19114,N_17743);
nor U20806 (N_20806,N_19572,N_17509);
xor U20807 (N_20807,N_17938,N_17659);
xor U20808 (N_20808,N_19630,N_17629);
or U20809 (N_20809,N_19469,N_18795);
xnor U20810 (N_20810,N_18757,N_18661);
and U20811 (N_20811,N_18440,N_18518);
xnor U20812 (N_20812,N_18252,N_18116);
nor U20813 (N_20813,N_19556,N_19356);
xnor U20814 (N_20814,N_19938,N_19290);
nor U20815 (N_20815,N_19366,N_19419);
xnor U20816 (N_20816,N_19484,N_19691);
nor U20817 (N_20817,N_19339,N_18867);
nand U20818 (N_20818,N_19968,N_17767);
nand U20819 (N_20819,N_18660,N_18015);
xnor U20820 (N_20820,N_19417,N_18699);
and U20821 (N_20821,N_18711,N_19153);
nor U20822 (N_20822,N_19140,N_19896);
nor U20823 (N_20823,N_17755,N_19628);
nand U20824 (N_20824,N_17741,N_19970);
nor U20825 (N_20825,N_19227,N_17829);
and U20826 (N_20826,N_19261,N_18513);
or U20827 (N_20827,N_19845,N_19093);
xnor U20828 (N_20828,N_18873,N_18574);
and U20829 (N_20829,N_18285,N_18830);
xnor U20830 (N_20830,N_19993,N_19357);
nand U20831 (N_20831,N_19916,N_18256);
nand U20832 (N_20832,N_19611,N_17546);
nand U20833 (N_20833,N_17616,N_17882);
nor U20834 (N_20834,N_17627,N_18265);
and U20835 (N_20835,N_18793,N_19016);
xnor U20836 (N_20836,N_18853,N_19579);
nand U20837 (N_20837,N_18493,N_18657);
and U20838 (N_20838,N_18061,N_19158);
xnor U20839 (N_20839,N_18511,N_19444);
or U20840 (N_20840,N_19624,N_19904);
and U20841 (N_20841,N_17623,N_18829);
or U20842 (N_20842,N_18775,N_17995);
and U20843 (N_20843,N_19940,N_19582);
or U20844 (N_20844,N_19399,N_18404);
or U20845 (N_20845,N_19134,N_18042);
nor U20846 (N_20846,N_19758,N_17539);
nor U20847 (N_20847,N_17740,N_18750);
xnor U20848 (N_20848,N_18602,N_18114);
xor U20849 (N_20849,N_18056,N_18739);
xor U20850 (N_20850,N_19255,N_19048);
or U20851 (N_20851,N_18002,N_18227);
or U20852 (N_20852,N_18701,N_17566);
or U20853 (N_20853,N_18492,N_18262);
nor U20854 (N_20854,N_18328,N_17804);
and U20855 (N_20855,N_17950,N_19256);
or U20856 (N_20856,N_18317,N_17737);
and U20857 (N_20857,N_17862,N_18896);
and U20858 (N_20858,N_18713,N_18159);
nand U20859 (N_20859,N_19126,N_19839);
and U20860 (N_20860,N_19487,N_17722);
xor U20861 (N_20861,N_19432,N_17548);
xor U20862 (N_20862,N_18824,N_18333);
nor U20863 (N_20863,N_18145,N_17960);
and U20864 (N_20864,N_17730,N_18176);
nor U20865 (N_20865,N_19662,N_19345);
nor U20866 (N_20866,N_17674,N_19650);
xnor U20867 (N_20867,N_18432,N_18397);
nor U20868 (N_20868,N_18022,N_19807);
nand U20869 (N_20869,N_19670,N_19908);
nand U20870 (N_20870,N_18224,N_18902);
and U20871 (N_20871,N_17961,N_19937);
nand U20872 (N_20872,N_18010,N_19319);
xnor U20873 (N_20873,N_17584,N_17822);
nand U20874 (N_20874,N_18341,N_19060);
or U20875 (N_20875,N_19578,N_18409);
nor U20876 (N_20876,N_19413,N_18011);
nor U20877 (N_20877,N_19404,N_19116);
or U20878 (N_20878,N_17680,N_18779);
or U20879 (N_20879,N_18229,N_18564);
and U20880 (N_20880,N_19734,N_17628);
or U20881 (N_20881,N_18238,N_19901);
nand U20882 (N_20882,N_19402,N_17644);
nand U20883 (N_20883,N_17799,N_19551);
xor U20884 (N_20884,N_18639,N_19324);
nor U20885 (N_20885,N_18922,N_18522);
xor U20886 (N_20886,N_17917,N_18566);
nand U20887 (N_20887,N_19489,N_18971);
and U20888 (N_20888,N_17967,N_17712);
or U20889 (N_20889,N_18977,N_19174);
xnor U20890 (N_20890,N_19608,N_19653);
or U20891 (N_20891,N_19719,N_18667);
xor U20892 (N_20892,N_19275,N_18289);
nor U20893 (N_20893,N_19903,N_18874);
or U20894 (N_20894,N_18392,N_18680);
xnor U20895 (N_20895,N_18347,N_19941);
and U20896 (N_20896,N_18846,N_19835);
and U20897 (N_20897,N_18903,N_17596);
xnor U20898 (N_20898,N_18998,N_19625);
xnor U20899 (N_20899,N_19987,N_19620);
and U20900 (N_20900,N_19199,N_18626);
xnor U20901 (N_20901,N_19005,N_17657);
nand U20902 (N_20902,N_17890,N_18952);
and U20903 (N_20903,N_19019,N_19425);
or U20904 (N_20904,N_17554,N_19302);
nand U20905 (N_20905,N_19935,N_18832);
nand U20906 (N_20906,N_17769,N_18205);
or U20907 (N_20907,N_17832,N_18097);
and U20908 (N_20908,N_18154,N_19584);
or U20909 (N_20909,N_18863,N_17801);
or U20910 (N_20910,N_18652,N_17641);
or U20911 (N_20911,N_19613,N_19121);
or U20912 (N_20912,N_18127,N_19282);
or U20913 (N_20913,N_18809,N_18188);
or U20914 (N_20914,N_18374,N_19269);
xnor U20915 (N_20915,N_18309,N_18864);
nor U20916 (N_20916,N_18825,N_17537);
or U20917 (N_20917,N_18298,N_18264);
nand U20918 (N_20918,N_17934,N_19293);
xnor U20919 (N_20919,N_18515,N_18683);
or U20920 (N_20920,N_19874,N_18984);
nand U20921 (N_20921,N_19706,N_19790);
nand U20922 (N_20922,N_18609,N_18441);
nor U20923 (N_20923,N_17786,N_19745);
or U20924 (N_20924,N_19775,N_17605);
nand U20925 (N_20925,N_18497,N_17833);
xor U20926 (N_20926,N_19437,N_18381);
xnor U20927 (N_20927,N_18245,N_19274);
and U20928 (N_20928,N_17553,N_19173);
and U20929 (N_20929,N_19456,N_17532);
nor U20930 (N_20930,N_17770,N_19420);
xor U20931 (N_20931,N_17793,N_19586);
or U20932 (N_20932,N_18405,N_18343);
nor U20933 (N_20933,N_19750,N_17851);
or U20934 (N_20934,N_19303,N_19434);
xor U20935 (N_20935,N_19851,N_19359);
and U20936 (N_20936,N_19001,N_19883);
xor U20937 (N_20937,N_19894,N_17849);
or U20938 (N_20938,N_18581,N_19406);
or U20939 (N_20939,N_19022,N_17873);
or U20940 (N_20940,N_19252,N_18184);
nand U20941 (N_20941,N_18039,N_19678);
and U20942 (N_20942,N_17729,N_17701);
and U20943 (N_20943,N_19791,N_19448);
nand U20944 (N_20944,N_18207,N_17791);
nand U20945 (N_20945,N_19794,N_18741);
xnor U20946 (N_20946,N_18119,N_17731);
and U20947 (N_20947,N_19963,N_19378);
and U20948 (N_20948,N_19629,N_19810);
nor U20949 (N_20949,N_19337,N_19566);
nor U20950 (N_20950,N_17863,N_18364);
and U20951 (N_20951,N_17959,N_17782);
xor U20952 (N_20952,N_18893,N_17519);
xor U20953 (N_20953,N_19254,N_19264);
xor U20954 (N_20954,N_18728,N_17908);
xor U20955 (N_20955,N_19660,N_17816);
nor U20956 (N_20956,N_18278,N_18158);
nor U20957 (N_20957,N_19512,N_19832);
nand U20958 (N_20958,N_17836,N_17841);
nand U20959 (N_20959,N_17925,N_18565);
or U20960 (N_20960,N_19232,N_18692);
nand U20961 (N_20961,N_19713,N_18534);
xnor U20962 (N_20962,N_18709,N_18491);
xor U20963 (N_20963,N_19312,N_18401);
nand U20964 (N_20964,N_17788,N_19128);
nand U20965 (N_20965,N_17582,N_19964);
or U20966 (N_20966,N_18724,N_18681);
xnor U20967 (N_20967,N_18170,N_17935);
nor U20968 (N_20968,N_19421,N_17831);
nor U20969 (N_20969,N_18990,N_18558);
or U20970 (N_20970,N_19299,N_19479);
and U20971 (N_20971,N_17983,N_19305);
nor U20972 (N_20972,N_18702,N_17899);
or U20973 (N_20973,N_18524,N_18691);
nand U20974 (N_20974,N_18980,N_19501);
xor U20975 (N_20975,N_19225,N_19059);
or U20976 (N_20976,N_19768,N_19180);
xnor U20977 (N_20977,N_18753,N_18149);
or U20978 (N_20978,N_18241,N_19267);
nand U20979 (N_20979,N_18504,N_18417);
xor U20980 (N_20980,N_18120,N_18270);
and U20981 (N_20981,N_18160,N_18230);
nor U20982 (N_20982,N_19342,N_19178);
nor U20983 (N_20983,N_18710,N_19881);
nand U20984 (N_20984,N_19343,N_17653);
nand U20985 (N_20985,N_19195,N_18065);
xnor U20986 (N_20986,N_18403,N_17691);
nor U20987 (N_20987,N_18125,N_19266);
nor U20988 (N_20988,N_18760,N_18817);
or U20989 (N_20989,N_18510,N_18616);
xnor U20990 (N_20990,N_19979,N_19451);
or U20991 (N_20991,N_17949,N_18372);
and U20992 (N_20992,N_19156,N_18506);
nor U20993 (N_20993,N_19661,N_19046);
nor U20994 (N_20994,N_19541,N_17545);
nor U20995 (N_20995,N_17763,N_19216);
and U20996 (N_20996,N_18533,N_19513);
and U20997 (N_20997,N_17524,N_19155);
or U20998 (N_20998,N_18425,N_19271);
or U20999 (N_20999,N_19248,N_19543);
nand U21000 (N_21000,N_19860,N_19673);
nor U21001 (N_21001,N_18622,N_19837);
nand U21002 (N_21002,N_19449,N_18480);
or U21003 (N_21003,N_18964,N_19096);
and U21004 (N_21004,N_19936,N_17717);
or U21005 (N_21005,N_18276,N_19588);
nor U21006 (N_21006,N_18054,N_18987);
or U21007 (N_21007,N_18789,N_19485);
or U21008 (N_21008,N_17904,N_18889);
or U21009 (N_21009,N_18454,N_19105);
and U21010 (N_21010,N_18431,N_18758);
and U21011 (N_21011,N_18281,N_19797);
xnor U21012 (N_21012,N_19340,N_18196);
or U21013 (N_21013,N_19567,N_18148);
xor U21014 (N_21014,N_18956,N_19488);
nand U21015 (N_21015,N_17504,N_19281);
nor U21016 (N_21016,N_17675,N_19395);
xnor U21017 (N_21017,N_18164,N_19222);
and U21018 (N_21018,N_19742,N_19646);
and U21019 (N_21019,N_18517,N_17678);
nand U21020 (N_21020,N_17550,N_19042);
and U21021 (N_21021,N_17941,N_19757);
nand U21022 (N_21022,N_18927,N_17965);
and U21023 (N_21023,N_17668,N_19648);
and U21024 (N_21024,N_19599,N_19943);
nand U21025 (N_21025,N_19498,N_19917);
and U21026 (N_21026,N_19306,N_18957);
nor U21027 (N_21027,N_19085,N_19233);
nor U21028 (N_21028,N_19346,N_18260);
nor U21029 (N_21029,N_18751,N_17560);
and U21030 (N_21030,N_17880,N_19062);
nand U21031 (N_21031,N_19524,N_19066);
xnor U21032 (N_21032,N_18525,N_19167);
nor U21033 (N_21033,N_19709,N_19003);
or U21034 (N_21034,N_18203,N_18171);
and U21035 (N_21035,N_18436,N_17868);
xor U21036 (N_21036,N_18805,N_18311);
or U21037 (N_21037,N_19763,N_19783);
xor U21038 (N_21038,N_19614,N_18090);
and U21039 (N_21039,N_18726,N_17525);
or U21040 (N_21040,N_19439,N_19597);
nand U21041 (N_21041,N_18313,N_19238);
xnor U21042 (N_21042,N_18018,N_17848);
nand U21043 (N_21043,N_18658,N_17671);
nor U21044 (N_21044,N_17820,N_19291);
nand U21045 (N_21045,N_19176,N_19915);
and U21046 (N_21046,N_18003,N_19374);
nand U21047 (N_21047,N_17761,N_19923);
or U21048 (N_21048,N_18861,N_19962);
xor U21049 (N_21049,N_18721,N_18676);
nor U21050 (N_21050,N_19186,N_18582);
xor U21051 (N_21051,N_19609,N_17975);
nor U21052 (N_21052,N_18520,N_19467);
or U21053 (N_21053,N_18672,N_19054);
and U21054 (N_21054,N_18376,N_19641);
nand U21055 (N_21055,N_17664,N_18648);
nor U21056 (N_21056,N_19304,N_18246);
or U21057 (N_21057,N_19575,N_19429);
nor U21058 (N_21058,N_19056,N_19520);
and U21059 (N_21059,N_18306,N_18596);
nand U21060 (N_21060,N_19914,N_19204);
xor U21061 (N_21061,N_18865,N_18290);
nor U21062 (N_21062,N_19954,N_19058);
or U21063 (N_21063,N_19774,N_18784);
nand U21064 (N_21064,N_19034,N_19220);
or U21065 (N_21065,N_18218,N_18584);
and U21066 (N_21066,N_18183,N_19533);
nand U21067 (N_21067,N_18644,N_17760);
nor U21068 (N_21068,N_19024,N_18088);
nor U21069 (N_21069,N_19748,N_17996);
nand U21070 (N_21070,N_18983,N_18418);
nand U21071 (N_21071,N_19242,N_18357);
nor U21072 (N_21072,N_19977,N_18954);
and U21073 (N_21073,N_19031,N_19119);
and U21074 (N_21074,N_19549,N_18674);
xor U21075 (N_21075,N_18651,N_18834);
or U21076 (N_21076,N_18778,N_18031);
xor U21077 (N_21077,N_18858,N_19200);
or U21078 (N_21078,N_18307,N_19583);
nor U21079 (N_21079,N_17858,N_19084);
nor U21080 (N_21080,N_17746,N_19452);
xnor U21081 (N_21081,N_18759,N_19308);
and U21082 (N_21082,N_19082,N_18040);
nor U21083 (N_21083,N_18215,N_17521);
nor U21084 (N_21084,N_17630,N_18304);
and U21085 (N_21085,N_18774,N_19335);
nor U21086 (N_21086,N_19830,N_19286);
and U21087 (N_21087,N_17690,N_18451);
or U21088 (N_21088,N_19605,N_19355);
or U21089 (N_21089,N_18694,N_17974);
xor U21090 (N_21090,N_18226,N_19539);
nand U21091 (N_21091,N_19462,N_19202);
or U21092 (N_21092,N_18901,N_17631);
nand U21093 (N_21093,N_18326,N_19658);
and U21094 (N_21094,N_17648,N_18337);
and U21095 (N_21095,N_18538,N_18286);
xnor U21096 (N_21096,N_19909,N_19585);
nand U21097 (N_21097,N_17818,N_19720);
nor U21098 (N_21098,N_18871,N_18496);
xnor U21099 (N_21099,N_18783,N_18557);
xor U21100 (N_21100,N_19455,N_17692);
or U21101 (N_21101,N_18923,N_18327);
nor U21102 (N_21102,N_17914,N_18458);
xnor U21103 (N_21103,N_17776,N_19865);
or U21104 (N_21104,N_19169,N_17700);
nor U21105 (N_21105,N_17856,N_18308);
and U21106 (N_21106,N_19470,N_18812);
and U21107 (N_21107,N_19465,N_17738);
and U21108 (N_21108,N_18195,N_19921);
nand U21109 (N_21109,N_19568,N_19590);
xor U21110 (N_21110,N_17611,N_18335);
xnor U21111 (N_21111,N_18232,N_18621);
xor U21112 (N_21112,N_19460,N_17894);
nor U21113 (N_21113,N_17604,N_18453);
xnor U21114 (N_21114,N_18543,N_18880);
or U21115 (N_21115,N_17704,N_18058);
nand U21116 (N_21116,N_18883,N_19313);
and U21117 (N_21117,N_18220,N_19778);
or U21118 (N_21118,N_19430,N_19518);
and U21119 (N_21119,N_18804,N_17859);
xor U21120 (N_21120,N_19988,N_18835);
nand U21121 (N_21121,N_18591,N_18275);
xor U21122 (N_21122,N_17897,N_18200);
or U21123 (N_21123,N_18118,N_18826);
xnor U21124 (N_21124,N_17952,N_17579);
xnor U21125 (N_21125,N_19081,N_18194);
or U21126 (N_21126,N_19598,N_19694);
xor U21127 (N_21127,N_19704,N_17774);
and U21128 (N_21128,N_17944,N_18494);
nand U21129 (N_21129,N_17513,N_18213);
xnor U21130 (N_21130,N_18569,N_17916);
xor U21131 (N_21131,N_18933,N_18851);
nand U21132 (N_21132,N_18426,N_18310);
nor U21133 (N_21133,N_18955,N_19307);
nand U21134 (N_21134,N_18614,N_17649);
and U21135 (N_21135,N_19946,N_18085);
nand U21136 (N_21136,N_18796,N_18348);
nand U21137 (N_21137,N_17590,N_17640);
and U21138 (N_21138,N_19553,N_19078);
or U21139 (N_21139,N_18682,N_19090);
and U21140 (N_21140,N_17980,N_19013);
nand U21141 (N_21141,N_18316,N_19735);
or U21142 (N_21142,N_18081,N_19942);
nand U21143 (N_21143,N_17538,N_18106);
nand U21144 (N_21144,N_18151,N_18886);
nor U21145 (N_21145,N_19336,N_18109);
xnor U21146 (N_21146,N_17637,N_18187);
nor U21147 (N_21147,N_19207,N_18387);
and U21148 (N_21148,N_19412,N_18716);
xnor U21149 (N_21149,N_17861,N_17556);
and U21150 (N_21150,N_19672,N_19138);
or U21151 (N_21151,N_19844,N_18806);
nor U21152 (N_21152,N_18801,N_18550);
nand U21153 (N_21153,N_18448,N_17552);
xnor U21154 (N_21154,N_17921,N_17606);
xor U21155 (N_21155,N_19323,N_17503);
or U21156 (N_21156,N_19642,N_19875);
nand U21157 (N_21157,N_18400,N_18781);
nor U21158 (N_21158,N_18228,N_18501);
and U21159 (N_21159,N_18013,N_18974);
or U21160 (N_21160,N_18752,N_19150);
and U21161 (N_21161,N_18556,N_19838);
xor U21162 (N_21162,N_18996,N_19638);
nand U21163 (N_21163,N_19050,N_18078);
or U21164 (N_21164,N_18132,N_19659);
nand U21165 (N_21165,N_17571,N_18930);
and U21166 (N_21166,N_18594,N_18855);
xnor U21167 (N_21167,N_19973,N_18483);
or U21168 (N_21168,N_18828,N_18043);
nor U21169 (N_21169,N_19828,N_17805);
nand U21170 (N_21170,N_17528,N_18438);
and U21171 (N_21171,N_17523,N_17520);
or U21172 (N_21172,N_17998,N_18101);
and U21173 (N_21173,N_19142,N_18487);
and U21174 (N_21174,N_18254,N_19891);
and U21175 (N_21175,N_18790,N_17990);
xnor U21176 (N_21176,N_19529,N_17986);
nand U21177 (N_21177,N_19500,N_19785);
xor U21178 (N_21178,N_19561,N_17903);
and U21179 (N_21179,N_19564,N_17901);
and U21180 (N_21180,N_18523,N_18462);
nand U21181 (N_21181,N_18368,N_19364);
xnor U21182 (N_21182,N_18280,N_18797);
nand U21183 (N_21183,N_17577,N_18986);
and U21184 (N_21184,N_19913,N_18168);
nand U21185 (N_21185,N_18485,N_19863);
nand U21186 (N_21186,N_19898,N_19289);
xor U21187 (N_21187,N_19447,N_18305);
nor U21188 (N_21188,N_19428,N_19482);
or U21189 (N_21189,N_19280,N_19806);
nor U21190 (N_21190,N_19836,N_18163);
xnor U21191 (N_21191,N_19798,N_18437);
nand U21192 (N_21192,N_19283,N_17891);
and U21193 (N_21193,N_18528,N_19481);
xor U21194 (N_21194,N_19029,N_17595);
xor U21195 (N_21195,N_19994,N_17828);
or U21196 (N_21196,N_19392,N_17734);
and U21197 (N_21197,N_19400,N_18988);
nand U21198 (N_21198,N_18464,N_18647);
nor U21199 (N_21199,N_18291,N_18161);
nor U21200 (N_21200,N_18968,N_19665);
nor U21201 (N_21201,N_18295,N_19235);
and U21202 (N_21202,N_18051,N_18380);
nand U21203 (N_21203,N_19334,N_17666);
nor U21204 (N_21204,N_19442,N_18856);
and U21205 (N_21205,N_19494,N_19361);
or U21206 (N_21206,N_19842,N_19718);
nand U21207 (N_21207,N_18615,N_18470);
or U21208 (N_21208,N_17857,N_18519);
nand U21209 (N_21209,N_19311,N_19723);
nor U21210 (N_21210,N_17780,N_17928);
and U21211 (N_21211,N_19808,N_18032);
or U21212 (N_21212,N_19473,N_18422);
or U21213 (N_21213,N_19433,N_18112);
xor U21214 (N_21214,N_19214,N_18049);
nand U21215 (N_21215,N_17711,N_18498);
xnor U21216 (N_21216,N_17872,N_18979);
or U21217 (N_21217,N_19920,N_19185);
or U21218 (N_21218,N_18370,N_18684);
nand U21219 (N_21219,N_18915,N_17762);
and U21220 (N_21220,N_18060,N_19856);
or U21221 (N_21221,N_17878,N_19370);
nor U21222 (N_21222,N_18447,N_17834);
xor U21223 (N_21223,N_18601,N_17733);
and U21224 (N_21224,N_18842,N_17617);
nor U21225 (N_21225,N_19491,N_18666);
xnor U21226 (N_21226,N_17647,N_19872);
nand U21227 (N_21227,N_18597,N_18857);
or U21228 (N_21228,N_18103,N_18465);
xor U21229 (N_21229,N_19037,N_17806);
and U21230 (N_21230,N_17567,N_19687);
nor U21231 (N_21231,N_17505,N_19980);
or U21232 (N_21232,N_19631,N_19352);
xor U21233 (N_21233,N_18568,N_19063);
or U21234 (N_21234,N_19651,N_19088);
xor U21235 (N_21235,N_18697,N_19243);
nand U21236 (N_21236,N_17932,N_19329);
nor U21237 (N_21237,N_18330,N_17685);
nor U21238 (N_21238,N_17619,N_18108);
nand U21239 (N_21239,N_18300,N_19724);
nand U21240 (N_21240,N_18899,N_19075);
or U21241 (N_21241,N_18637,N_18488);
and U21242 (N_21242,N_18548,N_18365);
xnor U21243 (N_21243,N_17893,N_19157);
nand U21244 (N_21244,N_18079,N_19217);
nand U21245 (N_21245,N_17840,N_19327);
nor U21246 (N_21246,N_17905,N_19986);
xor U21247 (N_21247,N_17808,N_19841);
xnor U21248 (N_21248,N_18091,N_18947);
nand U21249 (N_21249,N_19130,N_18578);
xor U21250 (N_21250,N_17615,N_19992);
xor U21251 (N_21251,N_19006,N_19328);
nand U21252 (N_21252,N_18286,N_19400);
nor U21253 (N_21253,N_18346,N_19914);
and U21254 (N_21254,N_17502,N_17632);
nor U21255 (N_21255,N_17858,N_17575);
nand U21256 (N_21256,N_18205,N_18944);
nand U21257 (N_21257,N_19631,N_18464);
nor U21258 (N_21258,N_18126,N_18881);
xnor U21259 (N_21259,N_19532,N_17702);
nor U21260 (N_21260,N_18690,N_17852);
nor U21261 (N_21261,N_19979,N_18947);
nor U21262 (N_21262,N_18017,N_17848);
xor U21263 (N_21263,N_18545,N_19894);
nor U21264 (N_21264,N_19565,N_19206);
nor U21265 (N_21265,N_19725,N_19481);
nand U21266 (N_21266,N_19191,N_19222);
nor U21267 (N_21267,N_18064,N_18012);
nand U21268 (N_21268,N_19915,N_19494);
nand U21269 (N_21269,N_18108,N_17764);
or U21270 (N_21270,N_18775,N_18729);
or U21271 (N_21271,N_17702,N_18126);
nand U21272 (N_21272,N_19505,N_18567);
and U21273 (N_21273,N_19687,N_18002);
nand U21274 (N_21274,N_19847,N_17730);
xor U21275 (N_21275,N_17919,N_18186);
nand U21276 (N_21276,N_17677,N_18141);
and U21277 (N_21277,N_19887,N_17683);
and U21278 (N_21278,N_19012,N_17969);
xor U21279 (N_21279,N_18027,N_18999);
xnor U21280 (N_21280,N_18974,N_19877);
or U21281 (N_21281,N_19646,N_18099);
xnor U21282 (N_21282,N_17523,N_17644);
or U21283 (N_21283,N_18995,N_19324);
xor U21284 (N_21284,N_18175,N_17804);
xor U21285 (N_21285,N_19023,N_18492);
nand U21286 (N_21286,N_19286,N_18624);
nand U21287 (N_21287,N_19805,N_19921);
xor U21288 (N_21288,N_19990,N_18932);
or U21289 (N_21289,N_18853,N_17780);
or U21290 (N_21290,N_18916,N_18288);
xor U21291 (N_21291,N_18189,N_19180);
and U21292 (N_21292,N_18655,N_19966);
nor U21293 (N_21293,N_19800,N_18234);
and U21294 (N_21294,N_18579,N_18187);
xnor U21295 (N_21295,N_18210,N_18605);
or U21296 (N_21296,N_18765,N_19494);
and U21297 (N_21297,N_18940,N_19993);
or U21298 (N_21298,N_17597,N_17926);
nand U21299 (N_21299,N_18750,N_18850);
xor U21300 (N_21300,N_18156,N_18426);
nand U21301 (N_21301,N_19537,N_19150);
nor U21302 (N_21302,N_19547,N_17670);
nor U21303 (N_21303,N_19984,N_18661);
and U21304 (N_21304,N_19089,N_18150);
nor U21305 (N_21305,N_18656,N_18768);
and U21306 (N_21306,N_18683,N_19789);
nor U21307 (N_21307,N_18147,N_19239);
xnor U21308 (N_21308,N_17529,N_17830);
xor U21309 (N_21309,N_18577,N_17803);
or U21310 (N_21310,N_18311,N_19774);
or U21311 (N_21311,N_18832,N_18904);
and U21312 (N_21312,N_17500,N_18873);
or U21313 (N_21313,N_18506,N_19223);
nand U21314 (N_21314,N_19116,N_18571);
and U21315 (N_21315,N_17761,N_19442);
nand U21316 (N_21316,N_19770,N_18629);
nor U21317 (N_21317,N_19157,N_19076);
or U21318 (N_21318,N_19016,N_19908);
or U21319 (N_21319,N_18090,N_18922);
nor U21320 (N_21320,N_18822,N_19481);
and U21321 (N_21321,N_17783,N_17690);
xor U21322 (N_21322,N_18832,N_17832);
nand U21323 (N_21323,N_18442,N_19153);
nand U21324 (N_21324,N_17813,N_17672);
xor U21325 (N_21325,N_19281,N_19278);
or U21326 (N_21326,N_19311,N_19806);
xnor U21327 (N_21327,N_19762,N_17600);
xor U21328 (N_21328,N_19599,N_19929);
nand U21329 (N_21329,N_18125,N_19983);
and U21330 (N_21330,N_19963,N_19923);
xnor U21331 (N_21331,N_19251,N_19077);
or U21332 (N_21332,N_19361,N_19365);
nand U21333 (N_21333,N_19374,N_18901);
nor U21334 (N_21334,N_18446,N_18032);
and U21335 (N_21335,N_18852,N_17803);
or U21336 (N_21336,N_17685,N_17515);
xnor U21337 (N_21337,N_19083,N_18414);
nand U21338 (N_21338,N_17547,N_18947);
nor U21339 (N_21339,N_18160,N_18636);
nand U21340 (N_21340,N_18866,N_18027);
xnor U21341 (N_21341,N_18019,N_17744);
nor U21342 (N_21342,N_18261,N_18604);
xor U21343 (N_21343,N_18145,N_18302);
nand U21344 (N_21344,N_19768,N_19787);
or U21345 (N_21345,N_18869,N_18200);
nand U21346 (N_21346,N_17778,N_18259);
nand U21347 (N_21347,N_19303,N_17914);
nand U21348 (N_21348,N_18001,N_17862);
or U21349 (N_21349,N_19087,N_18555);
or U21350 (N_21350,N_17547,N_18318);
and U21351 (N_21351,N_19455,N_19704);
and U21352 (N_21352,N_18037,N_17570);
xor U21353 (N_21353,N_18311,N_18124);
nand U21354 (N_21354,N_18852,N_19856);
or U21355 (N_21355,N_19900,N_17796);
nand U21356 (N_21356,N_19566,N_19314);
xor U21357 (N_21357,N_18726,N_19257);
nand U21358 (N_21358,N_19816,N_19629);
and U21359 (N_21359,N_19251,N_18310);
and U21360 (N_21360,N_19510,N_19270);
xnor U21361 (N_21361,N_18001,N_18947);
or U21362 (N_21362,N_19991,N_19458);
nor U21363 (N_21363,N_18289,N_19592);
nor U21364 (N_21364,N_19956,N_18033);
xor U21365 (N_21365,N_18547,N_18931);
nor U21366 (N_21366,N_18699,N_19127);
nor U21367 (N_21367,N_17958,N_19921);
and U21368 (N_21368,N_18519,N_18430);
nand U21369 (N_21369,N_19679,N_18718);
or U21370 (N_21370,N_18147,N_17797);
xnor U21371 (N_21371,N_19428,N_18300);
nand U21372 (N_21372,N_17938,N_19367);
or U21373 (N_21373,N_18105,N_19285);
nor U21374 (N_21374,N_18500,N_18115);
or U21375 (N_21375,N_19961,N_18692);
and U21376 (N_21376,N_18121,N_18161);
and U21377 (N_21377,N_19278,N_17900);
and U21378 (N_21378,N_19754,N_18741);
nor U21379 (N_21379,N_18456,N_18278);
nor U21380 (N_21380,N_19573,N_18812);
xnor U21381 (N_21381,N_18197,N_18242);
nand U21382 (N_21382,N_19011,N_19002);
or U21383 (N_21383,N_19710,N_17869);
or U21384 (N_21384,N_18149,N_18168);
and U21385 (N_21385,N_19314,N_19185);
and U21386 (N_21386,N_19355,N_19538);
or U21387 (N_21387,N_18858,N_18550);
nor U21388 (N_21388,N_19241,N_18610);
xor U21389 (N_21389,N_19802,N_18527);
or U21390 (N_21390,N_19618,N_17773);
nand U21391 (N_21391,N_19259,N_18771);
xnor U21392 (N_21392,N_18049,N_18521);
and U21393 (N_21393,N_19982,N_17940);
xor U21394 (N_21394,N_17551,N_19780);
xor U21395 (N_21395,N_18491,N_19979);
or U21396 (N_21396,N_18424,N_17603);
xor U21397 (N_21397,N_18527,N_19959);
or U21398 (N_21398,N_18641,N_18343);
and U21399 (N_21399,N_17708,N_18206);
nor U21400 (N_21400,N_18362,N_19138);
and U21401 (N_21401,N_18368,N_18552);
and U21402 (N_21402,N_18663,N_18344);
xnor U21403 (N_21403,N_19400,N_17702);
nand U21404 (N_21404,N_19805,N_17979);
and U21405 (N_21405,N_19343,N_18557);
and U21406 (N_21406,N_17677,N_18185);
nor U21407 (N_21407,N_18109,N_18231);
nand U21408 (N_21408,N_19713,N_18081);
nand U21409 (N_21409,N_17756,N_17751);
nor U21410 (N_21410,N_19358,N_19271);
nor U21411 (N_21411,N_19314,N_18669);
or U21412 (N_21412,N_19090,N_19415);
or U21413 (N_21413,N_18912,N_19183);
nand U21414 (N_21414,N_18169,N_19339);
or U21415 (N_21415,N_18802,N_19150);
and U21416 (N_21416,N_17804,N_18990);
nor U21417 (N_21417,N_18747,N_19644);
nor U21418 (N_21418,N_18199,N_17661);
or U21419 (N_21419,N_18051,N_18562);
nor U21420 (N_21420,N_19106,N_19296);
nand U21421 (N_21421,N_19915,N_19471);
xnor U21422 (N_21422,N_17689,N_19490);
or U21423 (N_21423,N_19545,N_17636);
nor U21424 (N_21424,N_18418,N_18821);
nand U21425 (N_21425,N_18483,N_19436);
nand U21426 (N_21426,N_19597,N_17670);
nand U21427 (N_21427,N_17539,N_18823);
nor U21428 (N_21428,N_19845,N_19823);
nand U21429 (N_21429,N_19828,N_17561);
nor U21430 (N_21430,N_17813,N_19808);
nand U21431 (N_21431,N_17697,N_18582);
xor U21432 (N_21432,N_17522,N_19435);
and U21433 (N_21433,N_19319,N_19996);
nand U21434 (N_21434,N_18141,N_19230);
or U21435 (N_21435,N_19817,N_19340);
and U21436 (N_21436,N_18379,N_18947);
xnor U21437 (N_21437,N_19022,N_19174);
nor U21438 (N_21438,N_19216,N_17669);
nor U21439 (N_21439,N_18777,N_19741);
nor U21440 (N_21440,N_19883,N_19579);
xnor U21441 (N_21441,N_17522,N_18818);
or U21442 (N_21442,N_18621,N_19313);
or U21443 (N_21443,N_18903,N_18938);
xnor U21444 (N_21444,N_19830,N_19003);
and U21445 (N_21445,N_19055,N_17973);
nor U21446 (N_21446,N_19814,N_17513);
or U21447 (N_21447,N_17716,N_17987);
nor U21448 (N_21448,N_19953,N_19427);
and U21449 (N_21449,N_18695,N_18928);
nand U21450 (N_21450,N_18780,N_19432);
nand U21451 (N_21451,N_17703,N_19652);
or U21452 (N_21452,N_19473,N_17871);
xor U21453 (N_21453,N_18056,N_19341);
and U21454 (N_21454,N_19149,N_17589);
nor U21455 (N_21455,N_19503,N_18159);
nor U21456 (N_21456,N_18485,N_18450);
or U21457 (N_21457,N_17519,N_18913);
xor U21458 (N_21458,N_17551,N_19009);
xnor U21459 (N_21459,N_19778,N_18887);
xor U21460 (N_21460,N_18894,N_18883);
xor U21461 (N_21461,N_19627,N_17729);
nand U21462 (N_21462,N_18526,N_19421);
nand U21463 (N_21463,N_19407,N_18281);
nand U21464 (N_21464,N_18594,N_19736);
nor U21465 (N_21465,N_17630,N_18402);
xor U21466 (N_21466,N_17835,N_18021);
and U21467 (N_21467,N_19569,N_18039);
nand U21468 (N_21468,N_17740,N_19096);
xnor U21469 (N_21469,N_17527,N_19900);
xor U21470 (N_21470,N_18187,N_18534);
nor U21471 (N_21471,N_18745,N_19995);
xnor U21472 (N_21472,N_19727,N_17815);
nor U21473 (N_21473,N_19564,N_18204);
nor U21474 (N_21474,N_19623,N_18889);
nor U21475 (N_21475,N_19016,N_17615);
nand U21476 (N_21476,N_19847,N_18190);
and U21477 (N_21477,N_17689,N_19229);
or U21478 (N_21478,N_18766,N_17573);
or U21479 (N_21479,N_18693,N_17709);
xor U21480 (N_21480,N_17766,N_19621);
xnor U21481 (N_21481,N_17638,N_19054);
and U21482 (N_21482,N_18829,N_19678);
nor U21483 (N_21483,N_19760,N_17952);
or U21484 (N_21484,N_18998,N_19478);
or U21485 (N_21485,N_19626,N_19578);
or U21486 (N_21486,N_17597,N_18503);
and U21487 (N_21487,N_19591,N_19163);
xnor U21488 (N_21488,N_18988,N_18814);
and U21489 (N_21489,N_18146,N_19151);
xnor U21490 (N_21490,N_18948,N_18567);
xor U21491 (N_21491,N_19369,N_19314);
nand U21492 (N_21492,N_18348,N_18538);
and U21493 (N_21493,N_17693,N_18604);
nand U21494 (N_21494,N_17634,N_18061);
and U21495 (N_21495,N_19813,N_19202);
xor U21496 (N_21496,N_17529,N_19654);
nand U21497 (N_21497,N_18440,N_18465);
and U21498 (N_21498,N_19599,N_18346);
and U21499 (N_21499,N_19432,N_19400);
or U21500 (N_21500,N_19993,N_18117);
nand U21501 (N_21501,N_19241,N_17814);
nand U21502 (N_21502,N_19609,N_19114);
xnor U21503 (N_21503,N_17594,N_18808);
or U21504 (N_21504,N_19542,N_18525);
nor U21505 (N_21505,N_18778,N_19066);
or U21506 (N_21506,N_17689,N_19012);
and U21507 (N_21507,N_17518,N_19406);
or U21508 (N_21508,N_18125,N_18434);
nor U21509 (N_21509,N_17812,N_17672);
nor U21510 (N_21510,N_19389,N_19966);
nand U21511 (N_21511,N_19954,N_17975);
xor U21512 (N_21512,N_19475,N_18129);
nor U21513 (N_21513,N_18461,N_19418);
nand U21514 (N_21514,N_19848,N_18926);
nand U21515 (N_21515,N_17654,N_18236);
xor U21516 (N_21516,N_17833,N_19236);
and U21517 (N_21517,N_18420,N_18949);
and U21518 (N_21518,N_19316,N_18250);
and U21519 (N_21519,N_17680,N_17634);
and U21520 (N_21520,N_19005,N_18117);
or U21521 (N_21521,N_19516,N_19419);
nor U21522 (N_21522,N_19673,N_17888);
or U21523 (N_21523,N_18088,N_17759);
nand U21524 (N_21524,N_19468,N_19971);
nand U21525 (N_21525,N_19617,N_19124);
xnor U21526 (N_21526,N_18686,N_19990);
nand U21527 (N_21527,N_17559,N_17669);
xnor U21528 (N_21528,N_18636,N_18155);
xnor U21529 (N_21529,N_19192,N_19313);
nor U21530 (N_21530,N_18301,N_19442);
xnor U21531 (N_21531,N_19969,N_19281);
and U21532 (N_21532,N_19170,N_18827);
nor U21533 (N_21533,N_18225,N_19861);
nor U21534 (N_21534,N_19492,N_18565);
nor U21535 (N_21535,N_18663,N_19656);
or U21536 (N_21536,N_18110,N_17640);
or U21537 (N_21537,N_19589,N_17769);
or U21538 (N_21538,N_18190,N_17919);
or U21539 (N_21539,N_17755,N_19470);
and U21540 (N_21540,N_18438,N_18413);
and U21541 (N_21541,N_18036,N_18826);
nand U21542 (N_21542,N_18308,N_19048);
and U21543 (N_21543,N_19780,N_19314);
nor U21544 (N_21544,N_19305,N_19043);
or U21545 (N_21545,N_18477,N_19672);
or U21546 (N_21546,N_19312,N_19421);
nor U21547 (N_21547,N_18192,N_19846);
nand U21548 (N_21548,N_19658,N_18598);
nand U21549 (N_21549,N_19022,N_17992);
nand U21550 (N_21550,N_17678,N_18058);
nor U21551 (N_21551,N_19518,N_19197);
xnor U21552 (N_21552,N_18557,N_17980);
or U21553 (N_21553,N_19397,N_19081);
nor U21554 (N_21554,N_17758,N_17583);
nor U21555 (N_21555,N_19589,N_19022);
nand U21556 (N_21556,N_19084,N_18237);
xor U21557 (N_21557,N_18671,N_17531);
or U21558 (N_21558,N_17990,N_19317);
nand U21559 (N_21559,N_19433,N_18696);
nand U21560 (N_21560,N_18518,N_19276);
nor U21561 (N_21561,N_19404,N_19478);
xor U21562 (N_21562,N_17736,N_18217);
and U21563 (N_21563,N_17641,N_17777);
nand U21564 (N_21564,N_19576,N_18379);
or U21565 (N_21565,N_18755,N_19065);
and U21566 (N_21566,N_17806,N_17643);
nor U21567 (N_21567,N_18447,N_19262);
nand U21568 (N_21568,N_19297,N_19488);
or U21569 (N_21569,N_17683,N_18458);
nand U21570 (N_21570,N_19272,N_18445);
nor U21571 (N_21571,N_18431,N_17935);
nand U21572 (N_21572,N_18258,N_18754);
xor U21573 (N_21573,N_19731,N_19597);
or U21574 (N_21574,N_18711,N_18458);
or U21575 (N_21575,N_17585,N_18981);
xor U21576 (N_21576,N_18057,N_18864);
nand U21577 (N_21577,N_19359,N_18398);
xor U21578 (N_21578,N_18306,N_18301);
or U21579 (N_21579,N_17965,N_19082);
nand U21580 (N_21580,N_18008,N_17814);
nand U21581 (N_21581,N_19668,N_18149);
nor U21582 (N_21582,N_17872,N_18387);
or U21583 (N_21583,N_17907,N_19426);
xor U21584 (N_21584,N_19377,N_19615);
or U21585 (N_21585,N_18051,N_18572);
xnor U21586 (N_21586,N_17680,N_19697);
nand U21587 (N_21587,N_19791,N_19789);
and U21588 (N_21588,N_19690,N_18758);
and U21589 (N_21589,N_18241,N_17936);
nand U21590 (N_21590,N_19091,N_18871);
nand U21591 (N_21591,N_19777,N_19263);
and U21592 (N_21592,N_18890,N_17644);
and U21593 (N_21593,N_17687,N_19767);
xor U21594 (N_21594,N_18429,N_17692);
and U21595 (N_21595,N_19988,N_17516);
or U21596 (N_21596,N_18781,N_18939);
nor U21597 (N_21597,N_17921,N_18345);
or U21598 (N_21598,N_19932,N_17679);
nand U21599 (N_21599,N_19332,N_19492);
nand U21600 (N_21600,N_18082,N_19213);
xnor U21601 (N_21601,N_19741,N_18266);
nor U21602 (N_21602,N_17827,N_19961);
xnor U21603 (N_21603,N_18819,N_19445);
nor U21604 (N_21604,N_19220,N_17592);
and U21605 (N_21605,N_18607,N_19813);
and U21606 (N_21606,N_18170,N_18556);
xnor U21607 (N_21607,N_19736,N_18315);
nor U21608 (N_21608,N_19899,N_18924);
and U21609 (N_21609,N_17605,N_18805);
and U21610 (N_21610,N_18207,N_19913);
nand U21611 (N_21611,N_18588,N_19712);
or U21612 (N_21612,N_18024,N_18513);
xor U21613 (N_21613,N_17823,N_19487);
or U21614 (N_21614,N_19242,N_19707);
and U21615 (N_21615,N_19073,N_19532);
and U21616 (N_21616,N_17547,N_19528);
and U21617 (N_21617,N_19588,N_18228);
nor U21618 (N_21618,N_19670,N_19318);
nand U21619 (N_21619,N_18689,N_18017);
or U21620 (N_21620,N_18396,N_18823);
xor U21621 (N_21621,N_19297,N_19418);
nand U21622 (N_21622,N_18948,N_18738);
or U21623 (N_21623,N_18218,N_17635);
and U21624 (N_21624,N_17802,N_18447);
or U21625 (N_21625,N_19833,N_19837);
or U21626 (N_21626,N_18354,N_18365);
or U21627 (N_21627,N_19111,N_18604);
nand U21628 (N_21628,N_19934,N_18628);
xnor U21629 (N_21629,N_18481,N_19240);
or U21630 (N_21630,N_19477,N_18623);
nand U21631 (N_21631,N_18101,N_18794);
nor U21632 (N_21632,N_18593,N_17879);
nand U21633 (N_21633,N_19499,N_18256);
xnor U21634 (N_21634,N_18539,N_18701);
nand U21635 (N_21635,N_18516,N_19267);
nand U21636 (N_21636,N_17898,N_18560);
xnor U21637 (N_21637,N_18851,N_18459);
nor U21638 (N_21638,N_18657,N_19722);
nand U21639 (N_21639,N_19271,N_19941);
nand U21640 (N_21640,N_17919,N_19874);
and U21641 (N_21641,N_19735,N_19883);
nand U21642 (N_21642,N_17982,N_18877);
xor U21643 (N_21643,N_19760,N_17775);
nor U21644 (N_21644,N_19733,N_18757);
nor U21645 (N_21645,N_19500,N_19632);
nor U21646 (N_21646,N_19619,N_19865);
nand U21647 (N_21647,N_18033,N_18797);
or U21648 (N_21648,N_18941,N_18781);
xnor U21649 (N_21649,N_18850,N_18016);
nand U21650 (N_21650,N_17887,N_17903);
or U21651 (N_21651,N_18368,N_18109);
xor U21652 (N_21652,N_18582,N_19070);
nand U21653 (N_21653,N_19182,N_17518);
nand U21654 (N_21654,N_19109,N_18456);
nand U21655 (N_21655,N_19107,N_19608);
or U21656 (N_21656,N_19458,N_18841);
and U21657 (N_21657,N_19526,N_17974);
or U21658 (N_21658,N_18838,N_17635);
nor U21659 (N_21659,N_18244,N_18225);
xor U21660 (N_21660,N_18230,N_18520);
and U21661 (N_21661,N_18633,N_19456);
or U21662 (N_21662,N_18460,N_18123);
or U21663 (N_21663,N_17725,N_19422);
or U21664 (N_21664,N_18919,N_18931);
xnor U21665 (N_21665,N_18080,N_19464);
nand U21666 (N_21666,N_18828,N_18879);
xor U21667 (N_21667,N_18171,N_19484);
nor U21668 (N_21668,N_18349,N_19145);
nor U21669 (N_21669,N_19496,N_18620);
nor U21670 (N_21670,N_19768,N_18605);
nor U21671 (N_21671,N_18246,N_18619);
xor U21672 (N_21672,N_18979,N_19042);
and U21673 (N_21673,N_19295,N_18609);
and U21674 (N_21674,N_19826,N_18794);
nor U21675 (N_21675,N_17971,N_19746);
and U21676 (N_21676,N_19649,N_18968);
nor U21677 (N_21677,N_19319,N_17698);
or U21678 (N_21678,N_19150,N_19861);
and U21679 (N_21679,N_17866,N_18393);
nand U21680 (N_21680,N_18313,N_17546);
nor U21681 (N_21681,N_19223,N_19381);
nor U21682 (N_21682,N_18981,N_18831);
nand U21683 (N_21683,N_19237,N_18820);
nand U21684 (N_21684,N_19633,N_18615);
nor U21685 (N_21685,N_19357,N_19758);
xnor U21686 (N_21686,N_17674,N_18120);
xnor U21687 (N_21687,N_18193,N_19247);
or U21688 (N_21688,N_19859,N_18393);
nor U21689 (N_21689,N_19766,N_18412);
nor U21690 (N_21690,N_17815,N_17713);
and U21691 (N_21691,N_18716,N_19914);
and U21692 (N_21692,N_19064,N_18033);
nor U21693 (N_21693,N_19011,N_19949);
and U21694 (N_21694,N_18625,N_17673);
xor U21695 (N_21695,N_19972,N_18402);
and U21696 (N_21696,N_19944,N_18591);
nor U21697 (N_21697,N_17920,N_19646);
or U21698 (N_21698,N_18639,N_17930);
nor U21699 (N_21699,N_19885,N_19134);
and U21700 (N_21700,N_18602,N_19623);
and U21701 (N_21701,N_19743,N_17699);
xnor U21702 (N_21702,N_18760,N_18602);
nand U21703 (N_21703,N_17743,N_17879);
or U21704 (N_21704,N_18665,N_17591);
xnor U21705 (N_21705,N_19616,N_18368);
or U21706 (N_21706,N_19833,N_17529);
nand U21707 (N_21707,N_18197,N_19818);
and U21708 (N_21708,N_19193,N_18098);
and U21709 (N_21709,N_18143,N_19259);
nand U21710 (N_21710,N_18783,N_17735);
nor U21711 (N_21711,N_18999,N_17831);
nor U21712 (N_21712,N_17783,N_17901);
xnor U21713 (N_21713,N_19403,N_17757);
or U21714 (N_21714,N_17826,N_19873);
nand U21715 (N_21715,N_17620,N_19825);
or U21716 (N_21716,N_18783,N_18178);
nand U21717 (N_21717,N_17907,N_17547);
and U21718 (N_21718,N_18116,N_19102);
xnor U21719 (N_21719,N_18683,N_19446);
nand U21720 (N_21720,N_18810,N_19386);
or U21721 (N_21721,N_19338,N_19921);
nor U21722 (N_21722,N_18281,N_18528);
nand U21723 (N_21723,N_18217,N_19459);
xnor U21724 (N_21724,N_18114,N_19060);
nand U21725 (N_21725,N_18646,N_19999);
and U21726 (N_21726,N_18878,N_17681);
xnor U21727 (N_21727,N_18845,N_19349);
nand U21728 (N_21728,N_19487,N_17595);
xor U21729 (N_21729,N_18186,N_18544);
nand U21730 (N_21730,N_19203,N_17728);
or U21731 (N_21731,N_17736,N_18825);
nor U21732 (N_21732,N_19070,N_18142);
or U21733 (N_21733,N_19152,N_18801);
nor U21734 (N_21734,N_17839,N_18982);
and U21735 (N_21735,N_18710,N_17846);
nor U21736 (N_21736,N_18201,N_18735);
nand U21737 (N_21737,N_19629,N_19369);
nor U21738 (N_21738,N_17695,N_18682);
and U21739 (N_21739,N_19210,N_19558);
and U21740 (N_21740,N_18961,N_18077);
nand U21741 (N_21741,N_19012,N_18011);
xnor U21742 (N_21742,N_18922,N_17729);
nand U21743 (N_21743,N_19076,N_19239);
or U21744 (N_21744,N_18760,N_18732);
nor U21745 (N_21745,N_18034,N_19563);
xnor U21746 (N_21746,N_18818,N_19204);
xnor U21747 (N_21747,N_18371,N_18468);
nand U21748 (N_21748,N_17879,N_19795);
nor U21749 (N_21749,N_17532,N_19339);
or U21750 (N_21750,N_19070,N_19997);
nand U21751 (N_21751,N_19507,N_17651);
xor U21752 (N_21752,N_18849,N_19688);
nor U21753 (N_21753,N_18936,N_18187);
and U21754 (N_21754,N_19273,N_18330);
nor U21755 (N_21755,N_19616,N_18405);
nand U21756 (N_21756,N_18819,N_19172);
nor U21757 (N_21757,N_18515,N_19424);
nand U21758 (N_21758,N_18425,N_19421);
or U21759 (N_21759,N_18639,N_19745);
xor U21760 (N_21760,N_19720,N_18650);
nand U21761 (N_21761,N_18950,N_18649);
nor U21762 (N_21762,N_18357,N_19512);
nand U21763 (N_21763,N_17928,N_17840);
nor U21764 (N_21764,N_19586,N_19926);
or U21765 (N_21765,N_19590,N_19703);
or U21766 (N_21766,N_18231,N_18569);
and U21767 (N_21767,N_19373,N_18369);
and U21768 (N_21768,N_17989,N_17723);
or U21769 (N_21769,N_18537,N_19302);
xnor U21770 (N_21770,N_19792,N_19134);
xor U21771 (N_21771,N_19018,N_17897);
nor U21772 (N_21772,N_17709,N_18277);
and U21773 (N_21773,N_19940,N_19422);
xnor U21774 (N_21774,N_19004,N_18320);
nor U21775 (N_21775,N_19041,N_17886);
or U21776 (N_21776,N_17550,N_18808);
nor U21777 (N_21777,N_19767,N_19332);
nor U21778 (N_21778,N_18778,N_18976);
and U21779 (N_21779,N_19541,N_19863);
and U21780 (N_21780,N_17711,N_18909);
xor U21781 (N_21781,N_19517,N_19668);
nand U21782 (N_21782,N_19172,N_18050);
and U21783 (N_21783,N_19060,N_18815);
nand U21784 (N_21784,N_19068,N_18150);
and U21785 (N_21785,N_18658,N_18408);
or U21786 (N_21786,N_19486,N_18787);
nor U21787 (N_21787,N_19981,N_17904);
nor U21788 (N_21788,N_18745,N_17631);
and U21789 (N_21789,N_17650,N_17698);
xor U21790 (N_21790,N_18563,N_18370);
xor U21791 (N_21791,N_19932,N_19927);
nand U21792 (N_21792,N_18400,N_19496);
nor U21793 (N_21793,N_17767,N_19460);
or U21794 (N_21794,N_18603,N_17956);
nor U21795 (N_21795,N_19216,N_17850);
nor U21796 (N_21796,N_19972,N_17677);
xor U21797 (N_21797,N_19416,N_18582);
and U21798 (N_21798,N_19651,N_19084);
xnor U21799 (N_21799,N_17596,N_18102);
nor U21800 (N_21800,N_18983,N_19671);
and U21801 (N_21801,N_18674,N_17717);
xnor U21802 (N_21802,N_18488,N_19758);
or U21803 (N_21803,N_18672,N_18288);
nor U21804 (N_21804,N_18490,N_19732);
nor U21805 (N_21805,N_17662,N_19850);
nor U21806 (N_21806,N_19914,N_18786);
xnor U21807 (N_21807,N_19319,N_19202);
nor U21808 (N_21808,N_18010,N_18083);
and U21809 (N_21809,N_19682,N_19963);
xor U21810 (N_21810,N_19332,N_19665);
or U21811 (N_21811,N_17788,N_18136);
nand U21812 (N_21812,N_18027,N_19071);
xnor U21813 (N_21813,N_17726,N_18632);
and U21814 (N_21814,N_18706,N_18999);
nor U21815 (N_21815,N_19241,N_19138);
xnor U21816 (N_21816,N_18877,N_18600);
nand U21817 (N_21817,N_19708,N_19510);
nor U21818 (N_21818,N_19786,N_18883);
or U21819 (N_21819,N_19882,N_19815);
nand U21820 (N_21820,N_17934,N_19642);
nand U21821 (N_21821,N_17932,N_19449);
xor U21822 (N_21822,N_18895,N_18934);
xor U21823 (N_21823,N_19249,N_19220);
xnor U21824 (N_21824,N_17776,N_19833);
xor U21825 (N_21825,N_17675,N_19954);
nor U21826 (N_21826,N_19391,N_19680);
and U21827 (N_21827,N_19321,N_18558);
and U21828 (N_21828,N_17754,N_18531);
and U21829 (N_21829,N_18567,N_19105);
xor U21830 (N_21830,N_18868,N_18234);
nand U21831 (N_21831,N_17973,N_18581);
and U21832 (N_21832,N_19055,N_19566);
nand U21833 (N_21833,N_18042,N_18824);
nor U21834 (N_21834,N_19045,N_17603);
nand U21835 (N_21835,N_18268,N_17682);
nor U21836 (N_21836,N_19990,N_19806);
nor U21837 (N_21837,N_18921,N_18154);
and U21838 (N_21838,N_18530,N_19477);
nor U21839 (N_21839,N_18185,N_19530);
or U21840 (N_21840,N_17866,N_18956);
xnor U21841 (N_21841,N_19482,N_19533);
and U21842 (N_21842,N_18405,N_17745);
nor U21843 (N_21843,N_18856,N_19783);
nand U21844 (N_21844,N_18172,N_17591);
or U21845 (N_21845,N_19998,N_19435);
nor U21846 (N_21846,N_17588,N_18926);
and U21847 (N_21847,N_18617,N_19684);
xor U21848 (N_21848,N_19546,N_18707);
nor U21849 (N_21849,N_19479,N_18644);
and U21850 (N_21850,N_18882,N_17522);
and U21851 (N_21851,N_18856,N_19695);
nand U21852 (N_21852,N_17708,N_18704);
xnor U21853 (N_21853,N_19879,N_17970);
or U21854 (N_21854,N_19191,N_19992);
nor U21855 (N_21855,N_18441,N_19638);
nand U21856 (N_21856,N_18543,N_17774);
and U21857 (N_21857,N_18794,N_19761);
and U21858 (N_21858,N_18280,N_19798);
nor U21859 (N_21859,N_18151,N_19437);
nand U21860 (N_21860,N_19942,N_19040);
nor U21861 (N_21861,N_19265,N_17835);
and U21862 (N_21862,N_17503,N_18575);
and U21863 (N_21863,N_18938,N_19739);
or U21864 (N_21864,N_19317,N_19631);
nand U21865 (N_21865,N_19455,N_17776);
nor U21866 (N_21866,N_19032,N_19738);
xnor U21867 (N_21867,N_18914,N_19435);
or U21868 (N_21868,N_19459,N_17772);
nor U21869 (N_21869,N_19415,N_19165);
nor U21870 (N_21870,N_19983,N_17951);
xor U21871 (N_21871,N_19496,N_19355);
xor U21872 (N_21872,N_19330,N_18317);
nand U21873 (N_21873,N_18978,N_19385);
nor U21874 (N_21874,N_18753,N_19383);
xnor U21875 (N_21875,N_18466,N_18032);
nand U21876 (N_21876,N_19835,N_18334);
or U21877 (N_21877,N_18853,N_18192);
xor U21878 (N_21878,N_19353,N_19305);
nor U21879 (N_21879,N_17912,N_17803);
nand U21880 (N_21880,N_19548,N_19033);
nor U21881 (N_21881,N_19673,N_19392);
or U21882 (N_21882,N_19978,N_19133);
nand U21883 (N_21883,N_19211,N_18185);
nand U21884 (N_21884,N_18277,N_19740);
and U21885 (N_21885,N_19320,N_18777);
nand U21886 (N_21886,N_18090,N_17534);
xor U21887 (N_21887,N_17959,N_19654);
nor U21888 (N_21888,N_18507,N_18016);
and U21889 (N_21889,N_19273,N_18181);
nand U21890 (N_21890,N_18838,N_18504);
and U21891 (N_21891,N_17841,N_19862);
or U21892 (N_21892,N_19216,N_19330);
xnor U21893 (N_21893,N_18803,N_18189);
xor U21894 (N_21894,N_17646,N_19441);
xnor U21895 (N_21895,N_18193,N_18628);
xnor U21896 (N_21896,N_17759,N_17594);
nand U21897 (N_21897,N_17795,N_19498);
nor U21898 (N_21898,N_19693,N_18336);
xnor U21899 (N_21899,N_17766,N_18354);
nand U21900 (N_21900,N_18989,N_19032);
and U21901 (N_21901,N_19800,N_18076);
nor U21902 (N_21902,N_18569,N_18932);
nor U21903 (N_21903,N_18529,N_17778);
xor U21904 (N_21904,N_19115,N_18855);
nand U21905 (N_21905,N_17928,N_18449);
nor U21906 (N_21906,N_18331,N_18367);
and U21907 (N_21907,N_18768,N_19128);
nand U21908 (N_21908,N_19768,N_17705);
nor U21909 (N_21909,N_18915,N_19328);
nor U21910 (N_21910,N_19617,N_19280);
nor U21911 (N_21911,N_19928,N_19065);
nand U21912 (N_21912,N_19270,N_17586);
and U21913 (N_21913,N_17812,N_19717);
and U21914 (N_21914,N_17620,N_18745);
xnor U21915 (N_21915,N_18087,N_18950);
or U21916 (N_21916,N_19759,N_18869);
and U21917 (N_21917,N_18080,N_18097);
or U21918 (N_21918,N_18088,N_17597);
xnor U21919 (N_21919,N_19426,N_19122);
or U21920 (N_21920,N_18931,N_19047);
or U21921 (N_21921,N_19342,N_17711);
or U21922 (N_21922,N_18843,N_19601);
xor U21923 (N_21923,N_17698,N_18750);
nand U21924 (N_21924,N_19801,N_19048);
xnor U21925 (N_21925,N_19157,N_17976);
nor U21926 (N_21926,N_18287,N_19123);
or U21927 (N_21927,N_19966,N_18767);
nand U21928 (N_21928,N_18193,N_17854);
or U21929 (N_21929,N_18417,N_18535);
or U21930 (N_21930,N_18927,N_19349);
xor U21931 (N_21931,N_18355,N_19363);
and U21932 (N_21932,N_18196,N_19311);
nand U21933 (N_21933,N_18721,N_19128);
nor U21934 (N_21934,N_18667,N_17848);
and U21935 (N_21935,N_18880,N_17542);
or U21936 (N_21936,N_17989,N_18157);
nand U21937 (N_21937,N_19546,N_18706);
and U21938 (N_21938,N_17568,N_19095);
xor U21939 (N_21939,N_18711,N_18134);
nor U21940 (N_21940,N_19737,N_17873);
xnor U21941 (N_21941,N_18910,N_18732);
nand U21942 (N_21942,N_19224,N_19791);
nand U21943 (N_21943,N_19657,N_19374);
nand U21944 (N_21944,N_17964,N_18029);
nand U21945 (N_21945,N_18795,N_19288);
and U21946 (N_21946,N_19639,N_17621);
nand U21947 (N_21947,N_18479,N_19278);
or U21948 (N_21948,N_18649,N_18361);
nor U21949 (N_21949,N_18189,N_18780);
and U21950 (N_21950,N_18233,N_19377);
and U21951 (N_21951,N_18652,N_18755);
and U21952 (N_21952,N_18567,N_19886);
or U21953 (N_21953,N_17710,N_17642);
nor U21954 (N_21954,N_17983,N_18441);
xnor U21955 (N_21955,N_19786,N_18602);
or U21956 (N_21956,N_19765,N_18221);
and U21957 (N_21957,N_17991,N_17568);
and U21958 (N_21958,N_19673,N_18900);
nor U21959 (N_21959,N_19119,N_18832);
nor U21960 (N_21960,N_18522,N_18915);
or U21961 (N_21961,N_18187,N_18949);
or U21962 (N_21962,N_18088,N_17796);
nand U21963 (N_21963,N_18152,N_18058);
and U21964 (N_21964,N_17941,N_17693);
xnor U21965 (N_21965,N_19242,N_18521);
and U21966 (N_21966,N_17661,N_19284);
or U21967 (N_21967,N_19088,N_18967);
and U21968 (N_21968,N_18708,N_17639);
nor U21969 (N_21969,N_18806,N_19066);
nor U21970 (N_21970,N_19657,N_19589);
nand U21971 (N_21971,N_18092,N_18223);
or U21972 (N_21972,N_18848,N_19843);
and U21973 (N_21973,N_17837,N_18105);
xnor U21974 (N_21974,N_18958,N_18452);
or U21975 (N_21975,N_19833,N_18852);
or U21976 (N_21976,N_18816,N_17516);
nor U21977 (N_21977,N_18824,N_18481);
nor U21978 (N_21978,N_17727,N_18405);
and U21979 (N_21979,N_19984,N_17857);
and U21980 (N_21980,N_18868,N_18019);
and U21981 (N_21981,N_17597,N_18597);
nand U21982 (N_21982,N_19811,N_17618);
or U21983 (N_21983,N_17738,N_17879);
xor U21984 (N_21984,N_17659,N_17597);
nor U21985 (N_21985,N_18989,N_17923);
nor U21986 (N_21986,N_17843,N_17741);
nor U21987 (N_21987,N_17800,N_18075);
and U21988 (N_21988,N_19743,N_18465);
or U21989 (N_21989,N_18228,N_17530);
nor U21990 (N_21990,N_19141,N_18779);
xor U21991 (N_21991,N_18945,N_18966);
nor U21992 (N_21992,N_18141,N_18807);
or U21993 (N_21993,N_18198,N_19110);
and U21994 (N_21994,N_19670,N_18222);
xor U21995 (N_21995,N_18663,N_17802);
and U21996 (N_21996,N_18985,N_18382);
xnor U21997 (N_21997,N_19614,N_18670);
xnor U21998 (N_21998,N_19615,N_18293);
nor U21999 (N_21999,N_19983,N_19548);
nand U22000 (N_22000,N_19689,N_19454);
nor U22001 (N_22001,N_17630,N_19684);
xor U22002 (N_22002,N_19471,N_19136);
xnor U22003 (N_22003,N_19960,N_18167);
and U22004 (N_22004,N_19688,N_18596);
and U22005 (N_22005,N_19461,N_19065);
or U22006 (N_22006,N_18007,N_18692);
nor U22007 (N_22007,N_19879,N_17769);
nor U22008 (N_22008,N_18234,N_17589);
nor U22009 (N_22009,N_19832,N_18158);
or U22010 (N_22010,N_19105,N_18375);
or U22011 (N_22011,N_18436,N_18918);
nor U22012 (N_22012,N_18395,N_19984);
nor U22013 (N_22013,N_17608,N_18890);
xnor U22014 (N_22014,N_18516,N_17519);
xnor U22015 (N_22015,N_19126,N_17628);
nor U22016 (N_22016,N_19120,N_18620);
nor U22017 (N_22017,N_18235,N_17550);
nor U22018 (N_22018,N_17633,N_19043);
or U22019 (N_22019,N_17923,N_18040);
and U22020 (N_22020,N_19181,N_19737);
nand U22021 (N_22021,N_18004,N_19170);
xnor U22022 (N_22022,N_17565,N_18819);
xnor U22023 (N_22023,N_17932,N_17652);
and U22024 (N_22024,N_18292,N_19715);
nand U22025 (N_22025,N_19358,N_18468);
nor U22026 (N_22026,N_19794,N_18733);
or U22027 (N_22027,N_18588,N_17819);
nand U22028 (N_22028,N_19548,N_18583);
or U22029 (N_22029,N_19007,N_18832);
and U22030 (N_22030,N_17667,N_19518);
or U22031 (N_22031,N_18296,N_18650);
and U22032 (N_22032,N_19633,N_18077);
xor U22033 (N_22033,N_18882,N_18573);
and U22034 (N_22034,N_17816,N_18401);
or U22035 (N_22035,N_19170,N_18380);
xor U22036 (N_22036,N_19682,N_18671);
nor U22037 (N_22037,N_17699,N_18267);
or U22038 (N_22038,N_17535,N_18205);
nand U22039 (N_22039,N_17875,N_19906);
xnor U22040 (N_22040,N_17947,N_18662);
xor U22041 (N_22041,N_19546,N_19176);
or U22042 (N_22042,N_18501,N_18224);
nand U22043 (N_22043,N_19164,N_19735);
nor U22044 (N_22044,N_18615,N_18054);
nand U22045 (N_22045,N_19554,N_19986);
nor U22046 (N_22046,N_18150,N_19402);
nand U22047 (N_22047,N_19880,N_18797);
nor U22048 (N_22048,N_19497,N_19143);
xor U22049 (N_22049,N_19394,N_18936);
or U22050 (N_22050,N_18467,N_19103);
nand U22051 (N_22051,N_18868,N_18461);
and U22052 (N_22052,N_18197,N_18760);
nand U22053 (N_22053,N_19426,N_19325);
and U22054 (N_22054,N_18122,N_18427);
or U22055 (N_22055,N_19694,N_18918);
xnor U22056 (N_22056,N_19096,N_17501);
or U22057 (N_22057,N_18501,N_18334);
and U22058 (N_22058,N_19547,N_17623);
nor U22059 (N_22059,N_19766,N_17668);
or U22060 (N_22060,N_18083,N_17774);
nor U22061 (N_22061,N_18631,N_19449);
nand U22062 (N_22062,N_18447,N_19278);
nand U22063 (N_22063,N_19395,N_18921);
and U22064 (N_22064,N_19486,N_18478);
nor U22065 (N_22065,N_18139,N_18888);
nand U22066 (N_22066,N_18217,N_19013);
nor U22067 (N_22067,N_19783,N_19483);
xnor U22068 (N_22068,N_18261,N_19349);
nand U22069 (N_22069,N_19322,N_19963);
or U22070 (N_22070,N_19637,N_19317);
xnor U22071 (N_22071,N_19530,N_18122);
and U22072 (N_22072,N_19661,N_18890);
and U22073 (N_22073,N_17670,N_18260);
nor U22074 (N_22074,N_18427,N_19306);
and U22075 (N_22075,N_18134,N_18594);
xnor U22076 (N_22076,N_17807,N_17867);
nor U22077 (N_22077,N_19587,N_19880);
or U22078 (N_22078,N_18558,N_17651);
xor U22079 (N_22079,N_18273,N_19645);
nand U22080 (N_22080,N_17967,N_19574);
or U22081 (N_22081,N_19791,N_18559);
nand U22082 (N_22082,N_19467,N_19435);
and U22083 (N_22083,N_18702,N_18684);
nand U22084 (N_22084,N_19686,N_17598);
nor U22085 (N_22085,N_18248,N_19030);
nand U22086 (N_22086,N_19398,N_19958);
xor U22087 (N_22087,N_18133,N_17728);
and U22088 (N_22088,N_19855,N_19993);
or U22089 (N_22089,N_19229,N_19089);
and U22090 (N_22090,N_19386,N_17714);
nand U22091 (N_22091,N_17616,N_18899);
nand U22092 (N_22092,N_17721,N_17600);
or U22093 (N_22093,N_18340,N_17843);
or U22094 (N_22094,N_18774,N_17916);
nand U22095 (N_22095,N_17725,N_18475);
nand U22096 (N_22096,N_18787,N_19585);
and U22097 (N_22097,N_19869,N_18907);
or U22098 (N_22098,N_17552,N_17513);
and U22099 (N_22099,N_19812,N_19449);
or U22100 (N_22100,N_19066,N_19585);
nand U22101 (N_22101,N_17876,N_17919);
nand U22102 (N_22102,N_17628,N_19549);
or U22103 (N_22103,N_18572,N_18504);
and U22104 (N_22104,N_17866,N_18463);
xnor U22105 (N_22105,N_19333,N_18636);
and U22106 (N_22106,N_19737,N_18185);
nor U22107 (N_22107,N_18411,N_18328);
nand U22108 (N_22108,N_18004,N_18425);
nand U22109 (N_22109,N_19165,N_18438);
nor U22110 (N_22110,N_18439,N_18219);
nand U22111 (N_22111,N_18588,N_17908);
nor U22112 (N_22112,N_18134,N_19519);
nand U22113 (N_22113,N_19336,N_17681);
xnor U22114 (N_22114,N_18243,N_17719);
and U22115 (N_22115,N_19896,N_18995);
nand U22116 (N_22116,N_19811,N_17819);
xnor U22117 (N_22117,N_18489,N_18987);
or U22118 (N_22118,N_19783,N_19369);
nor U22119 (N_22119,N_18384,N_19536);
nor U22120 (N_22120,N_18451,N_18059);
xnor U22121 (N_22121,N_17817,N_18040);
nand U22122 (N_22122,N_17587,N_17982);
and U22123 (N_22123,N_18968,N_17884);
or U22124 (N_22124,N_19772,N_19993);
nor U22125 (N_22125,N_17685,N_17848);
and U22126 (N_22126,N_18785,N_19032);
or U22127 (N_22127,N_18054,N_19829);
or U22128 (N_22128,N_18861,N_19144);
and U22129 (N_22129,N_18224,N_19117);
nand U22130 (N_22130,N_18930,N_19336);
nand U22131 (N_22131,N_17739,N_18840);
nand U22132 (N_22132,N_18002,N_17845);
and U22133 (N_22133,N_18670,N_17961);
or U22134 (N_22134,N_17597,N_18879);
xor U22135 (N_22135,N_18806,N_17788);
xnor U22136 (N_22136,N_19867,N_19368);
nor U22137 (N_22137,N_17769,N_19136);
or U22138 (N_22138,N_18739,N_19461);
xnor U22139 (N_22139,N_18884,N_18461);
and U22140 (N_22140,N_18025,N_18531);
or U22141 (N_22141,N_19595,N_18087);
and U22142 (N_22142,N_19729,N_19267);
xnor U22143 (N_22143,N_18927,N_19596);
xor U22144 (N_22144,N_17729,N_18192);
and U22145 (N_22145,N_18553,N_18697);
nand U22146 (N_22146,N_17666,N_19424);
xnor U22147 (N_22147,N_19838,N_18725);
nor U22148 (N_22148,N_17644,N_17744);
nor U22149 (N_22149,N_17852,N_17797);
nand U22150 (N_22150,N_19450,N_18208);
and U22151 (N_22151,N_17983,N_19288);
nand U22152 (N_22152,N_17614,N_19054);
nor U22153 (N_22153,N_17701,N_19367);
or U22154 (N_22154,N_18369,N_18215);
and U22155 (N_22155,N_18449,N_19142);
nand U22156 (N_22156,N_19808,N_18668);
and U22157 (N_22157,N_19406,N_19024);
xnor U22158 (N_22158,N_17985,N_18744);
xnor U22159 (N_22159,N_18593,N_18723);
and U22160 (N_22160,N_18945,N_19547);
and U22161 (N_22161,N_18415,N_18935);
nand U22162 (N_22162,N_19273,N_19190);
xor U22163 (N_22163,N_19075,N_18202);
xor U22164 (N_22164,N_19972,N_19311);
nand U22165 (N_22165,N_19613,N_17773);
nand U22166 (N_22166,N_18821,N_19106);
and U22167 (N_22167,N_18708,N_19550);
xor U22168 (N_22168,N_19882,N_17900);
nand U22169 (N_22169,N_18819,N_18106);
or U22170 (N_22170,N_18784,N_18795);
nand U22171 (N_22171,N_18216,N_18188);
nand U22172 (N_22172,N_18599,N_17534);
nand U22173 (N_22173,N_19619,N_18701);
or U22174 (N_22174,N_18014,N_18514);
nor U22175 (N_22175,N_17918,N_18694);
or U22176 (N_22176,N_19314,N_19612);
and U22177 (N_22177,N_18398,N_18976);
or U22178 (N_22178,N_18074,N_17782);
and U22179 (N_22179,N_19761,N_19271);
nor U22180 (N_22180,N_18462,N_19670);
nand U22181 (N_22181,N_19385,N_18356);
or U22182 (N_22182,N_19237,N_19360);
or U22183 (N_22183,N_18876,N_18797);
xnor U22184 (N_22184,N_18446,N_18080);
nand U22185 (N_22185,N_18973,N_19814);
nand U22186 (N_22186,N_19538,N_18601);
xor U22187 (N_22187,N_18897,N_18158);
and U22188 (N_22188,N_18745,N_19530);
nand U22189 (N_22189,N_19433,N_19780);
and U22190 (N_22190,N_18031,N_17921);
nor U22191 (N_22191,N_18791,N_18596);
or U22192 (N_22192,N_18331,N_17624);
xor U22193 (N_22193,N_18418,N_17847);
nand U22194 (N_22194,N_19269,N_18664);
nor U22195 (N_22195,N_19240,N_19758);
or U22196 (N_22196,N_19652,N_18952);
xor U22197 (N_22197,N_18503,N_18395);
and U22198 (N_22198,N_19192,N_18734);
nand U22199 (N_22199,N_18746,N_18873);
or U22200 (N_22200,N_18281,N_18031);
nand U22201 (N_22201,N_19998,N_18066);
nand U22202 (N_22202,N_19173,N_18966);
xnor U22203 (N_22203,N_18584,N_17751);
or U22204 (N_22204,N_18258,N_18269);
xor U22205 (N_22205,N_18103,N_18412);
or U22206 (N_22206,N_19729,N_18952);
nand U22207 (N_22207,N_19421,N_17882);
xor U22208 (N_22208,N_19889,N_17736);
and U22209 (N_22209,N_18937,N_17773);
and U22210 (N_22210,N_19237,N_18247);
xnor U22211 (N_22211,N_19426,N_18435);
nand U22212 (N_22212,N_18822,N_18692);
nor U22213 (N_22213,N_18917,N_19715);
and U22214 (N_22214,N_18519,N_19354);
and U22215 (N_22215,N_18677,N_17749);
nand U22216 (N_22216,N_19598,N_17711);
nor U22217 (N_22217,N_17500,N_17835);
nor U22218 (N_22218,N_18523,N_18642);
nand U22219 (N_22219,N_19583,N_18313);
or U22220 (N_22220,N_19284,N_17985);
nor U22221 (N_22221,N_19414,N_17861);
nor U22222 (N_22222,N_18998,N_18362);
or U22223 (N_22223,N_19289,N_19410);
nor U22224 (N_22224,N_17627,N_17535);
and U22225 (N_22225,N_17772,N_17818);
nand U22226 (N_22226,N_17997,N_17531);
or U22227 (N_22227,N_19874,N_18207);
xor U22228 (N_22228,N_19579,N_18967);
xnor U22229 (N_22229,N_17818,N_17658);
xnor U22230 (N_22230,N_18577,N_18413);
xnor U22231 (N_22231,N_18621,N_18429);
and U22232 (N_22232,N_17919,N_19953);
nand U22233 (N_22233,N_19196,N_18154);
and U22234 (N_22234,N_19984,N_19963);
or U22235 (N_22235,N_18911,N_18845);
and U22236 (N_22236,N_19350,N_19141);
xor U22237 (N_22237,N_18083,N_19865);
or U22238 (N_22238,N_17677,N_18690);
nand U22239 (N_22239,N_17777,N_18130);
nand U22240 (N_22240,N_17832,N_18808);
or U22241 (N_22241,N_17856,N_19546);
and U22242 (N_22242,N_18269,N_17887);
xor U22243 (N_22243,N_18754,N_17740);
or U22244 (N_22244,N_17885,N_18014);
nor U22245 (N_22245,N_18639,N_18174);
and U22246 (N_22246,N_18532,N_19074);
and U22247 (N_22247,N_19180,N_17696);
nand U22248 (N_22248,N_19293,N_18765);
nand U22249 (N_22249,N_19795,N_18955);
or U22250 (N_22250,N_19433,N_18867);
nand U22251 (N_22251,N_19411,N_18143);
and U22252 (N_22252,N_18522,N_19443);
xor U22253 (N_22253,N_19595,N_18206);
nor U22254 (N_22254,N_19856,N_18882);
or U22255 (N_22255,N_18145,N_19250);
and U22256 (N_22256,N_18976,N_17627);
xnor U22257 (N_22257,N_17875,N_19937);
or U22258 (N_22258,N_18706,N_19440);
xnor U22259 (N_22259,N_18032,N_18640);
and U22260 (N_22260,N_18560,N_18964);
nor U22261 (N_22261,N_19083,N_18161);
or U22262 (N_22262,N_19033,N_17675);
xnor U22263 (N_22263,N_18388,N_18316);
nand U22264 (N_22264,N_19881,N_19440);
or U22265 (N_22265,N_18417,N_19482);
and U22266 (N_22266,N_18218,N_18132);
xor U22267 (N_22267,N_19690,N_18335);
or U22268 (N_22268,N_19426,N_17522);
xnor U22269 (N_22269,N_18780,N_18991);
and U22270 (N_22270,N_19444,N_19878);
nor U22271 (N_22271,N_19319,N_18532);
nand U22272 (N_22272,N_18657,N_19804);
or U22273 (N_22273,N_19124,N_18414);
nand U22274 (N_22274,N_17926,N_18401);
nor U22275 (N_22275,N_18606,N_18443);
nand U22276 (N_22276,N_19014,N_19775);
xor U22277 (N_22277,N_19348,N_19173);
or U22278 (N_22278,N_19610,N_18527);
xor U22279 (N_22279,N_18143,N_19520);
and U22280 (N_22280,N_19035,N_17871);
nor U22281 (N_22281,N_19324,N_18515);
and U22282 (N_22282,N_19470,N_19688);
and U22283 (N_22283,N_18482,N_17782);
xor U22284 (N_22284,N_19337,N_19887);
xnor U22285 (N_22285,N_18055,N_19801);
and U22286 (N_22286,N_19554,N_19754);
and U22287 (N_22287,N_17762,N_18398);
nor U22288 (N_22288,N_19098,N_18690);
nand U22289 (N_22289,N_17529,N_18512);
nand U22290 (N_22290,N_19932,N_18063);
xor U22291 (N_22291,N_19488,N_18079);
nand U22292 (N_22292,N_17657,N_18764);
nor U22293 (N_22293,N_18967,N_19215);
and U22294 (N_22294,N_17799,N_17984);
nand U22295 (N_22295,N_18092,N_18053);
and U22296 (N_22296,N_19574,N_18910);
and U22297 (N_22297,N_18052,N_18787);
xor U22298 (N_22298,N_18186,N_19655);
or U22299 (N_22299,N_18084,N_18780);
xnor U22300 (N_22300,N_17777,N_18429);
xor U22301 (N_22301,N_18723,N_19430);
and U22302 (N_22302,N_19844,N_17995);
or U22303 (N_22303,N_19193,N_19265);
nand U22304 (N_22304,N_18723,N_18904);
xor U22305 (N_22305,N_18064,N_18810);
xor U22306 (N_22306,N_18311,N_17732);
nor U22307 (N_22307,N_18778,N_19141);
or U22308 (N_22308,N_18143,N_17970);
or U22309 (N_22309,N_19288,N_19698);
xnor U22310 (N_22310,N_17884,N_19499);
nand U22311 (N_22311,N_18323,N_19204);
nand U22312 (N_22312,N_19739,N_17860);
nand U22313 (N_22313,N_19614,N_18143);
and U22314 (N_22314,N_18401,N_19196);
nand U22315 (N_22315,N_19961,N_17677);
nor U22316 (N_22316,N_17923,N_19577);
and U22317 (N_22317,N_19870,N_19059);
and U22318 (N_22318,N_19783,N_19160);
xor U22319 (N_22319,N_18027,N_17561);
xnor U22320 (N_22320,N_18080,N_19873);
nand U22321 (N_22321,N_19579,N_17780);
xor U22322 (N_22322,N_19588,N_19055);
nand U22323 (N_22323,N_19593,N_18442);
nand U22324 (N_22324,N_19080,N_18319);
or U22325 (N_22325,N_18673,N_18496);
nand U22326 (N_22326,N_18822,N_19784);
or U22327 (N_22327,N_18396,N_19024);
nand U22328 (N_22328,N_19824,N_19564);
nor U22329 (N_22329,N_19192,N_18067);
or U22330 (N_22330,N_17681,N_18016);
nand U22331 (N_22331,N_17629,N_19709);
nor U22332 (N_22332,N_18063,N_19852);
nor U22333 (N_22333,N_18344,N_18195);
or U22334 (N_22334,N_19792,N_19328);
nand U22335 (N_22335,N_18024,N_19895);
xor U22336 (N_22336,N_18407,N_19142);
and U22337 (N_22337,N_19115,N_18040);
and U22338 (N_22338,N_19219,N_19807);
and U22339 (N_22339,N_19617,N_18495);
nand U22340 (N_22340,N_18664,N_18250);
and U22341 (N_22341,N_19842,N_19305);
nand U22342 (N_22342,N_18058,N_18059);
xnor U22343 (N_22343,N_17837,N_17649);
or U22344 (N_22344,N_18167,N_19199);
and U22345 (N_22345,N_19974,N_18355);
nand U22346 (N_22346,N_18752,N_18011);
nor U22347 (N_22347,N_18817,N_17548);
xnor U22348 (N_22348,N_17517,N_19947);
or U22349 (N_22349,N_17595,N_19829);
nand U22350 (N_22350,N_18372,N_18384);
nor U22351 (N_22351,N_18795,N_18436);
xnor U22352 (N_22352,N_18772,N_19245);
nor U22353 (N_22353,N_19486,N_18494);
nand U22354 (N_22354,N_18062,N_18991);
and U22355 (N_22355,N_18646,N_18387);
or U22356 (N_22356,N_19611,N_18198);
nor U22357 (N_22357,N_19662,N_18351);
and U22358 (N_22358,N_19261,N_18984);
or U22359 (N_22359,N_19388,N_19654);
or U22360 (N_22360,N_19293,N_18003);
and U22361 (N_22361,N_19832,N_18213);
xor U22362 (N_22362,N_18114,N_18115);
and U22363 (N_22363,N_17529,N_19992);
or U22364 (N_22364,N_18210,N_19557);
and U22365 (N_22365,N_17503,N_17571);
xnor U22366 (N_22366,N_18201,N_19458);
nor U22367 (N_22367,N_19228,N_19241);
nand U22368 (N_22368,N_18286,N_18181);
and U22369 (N_22369,N_19599,N_19081);
and U22370 (N_22370,N_18883,N_19613);
and U22371 (N_22371,N_18654,N_19407);
xnor U22372 (N_22372,N_19750,N_17536);
nand U22373 (N_22373,N_19296,N_19576);
nand U22374 (N_22374,N_19090,N_17931);
and U22375 (N_22375,N_19831,N_18528);
nor U22376 (N_22376,N_19630,N_19837);
and U22377 (N_22377,N_19440,N_19738);
nand U22378 (N_22378,N_18526,N_19716);
nor U22379 (N_22379,N_17685,N_19966);
xnor U22380 (N_22380,N_18110,N_17683);
nand U22381 (N_22381,N_19276,N_17779);
xnor U22382 (N_22382,N_19714,N_18106);
or U22383 (N_22383,N_17817,N_19947);
nor U22384 (N_22384,N_18332,N_19518);
and U22385 (N_22385,N_19654,N_18364);
or U22386 (N_22386,N_18149,N_17669);
or U22387 (N_22387,N_18124,N_18169);
nor U22388 (N_22388,N_18349,N_19710);
xnor U22389 (N_22389,N_19062,N_19710);
xor U22390 (N_22390,N_17705,N_18800);
nand U22391 (N_22391,N_17784,N_19953);
xnor U22392 (N_22392,N_19509,N_18146);
xnor U22393 (N_22393,N_18921,N_17773);
or U22394 (N_22394,N_19226,N_17665);
or U22395 (N_22395,N_18768,N_19041);
nand U22396 (N_22396,N_19887,N_17529);
nor U22397 (N_22397,N_19250,N_18467);
xor U22398 (N_22398,N_18872,N_19087);
or U22399 (N_22399,N_19095,N_19479);
or U22400 (N_22400,N_18471,N_19310);
or U22401 (N_22401,N_18817,N_18439);
and U22402 (N_22402,N_18066,N_18847);
nand U22403 (N_22403,N_19946,N_19132);
xnor U22404 (N_22404,N_18432,N_17548);
and U22405 (N_22405,N_17631,N_19901);
xor U22406 (N_22406,N_18619,N_18216);
nand U22407 (N_22407,N_18338,N_19700);
and U22408 (N_22408,N_18031,N_18290);
and U22409 (N_22409,N_18218,N_19366);
nor U22410 (N_22410,N_19863,N_19924);
nand U22411 (N_22411,N_18219,N_19284);
xnor U22412 (N_22412,N_18201,N_19261);
or U22413 (N_22413,N_19807,N_18445);
or U22414 (N_22414,N_19810,N_18462);
xnor U22415 (N_22415,N_17544,N_18431);
and U22416 (N_22416,N_18167,N_17568);
xor U22417 (N_22417,N_18149,N_18960);
or U22418 (N_22418,N_19836,N_19125);
nand U22419 (N_22419,N_19196,N_17887);
or U22420 (N_22420,N_19213,N_19387);
or U22421 (N_22421,N_17701,N_17585);
or U22422 (N_22422,N_18546,N_19415);
and U22423 (N_22423,N_17519,N_17971);
xnor U22424 (N_22424,N_17812,N_19342);
xor U22425 (N_22425,N_19792,N_18558);
or U22426 (N_22426,N_18169,N_19556);
or U22427 (N_22427,N_19212,N_17549);
nand U22428 (N_22428,N_19753,N_17885);
and U22429 (N_22429,N_17627,N_18382);
or U22430 (N_22430,N_19538,N_19950);
and U22431 (N_22431,N_17575,N_18212);
xor U22432 (N_22432,N_19024,N_18589);
and U22433 (N_22433,N_19831,N_19586);
or U22434 (N_22434,N_19705,N_18325);
or U22435 (N_22435,N_19415,N_17751);
nor U22436 (N_22436,N_18423,N_19393);
nor U22437 (N_22437,N_18721,N_18192);
nand U22438 (N_22438,N_18918,N_19377);
and U22439 (N_22439,N_18992,N_18177);
xor U22440 (N_22440,N_17767,N_17758);
xor U22441 (N_22441,N_17881,N_19559);
and U22442 (N_22442,N_19215,N_18347);
nand U22443 (N_22443,N_18441,N_18461);
xnor U22444 (N_22444,N_19352,N_17644);
and U22445 (N_22445,N_19679,N_19062);
nand U22446 (N_22446,N_18961,N_17945);
nor U22447 (N_22447,N_19151,N_18045);
and U22448 (N_22448,N_17821,N_19874);
or U22449 (N_22449,N_18703,N_19384);
nor U22450 (N_22450,N_18253,N_19803);
or U22451 (N_22451,N_18559,N_18455);
or U22452 (N_22452,N_17817,N_18614);
xnor U22453 (N_22453,N_18825,N_19984);
or U22454 (N_22454,N_19329,N_18504);
or U22455 (N_22455,N_19732,N_19922);
nor U22456 (N_22456,N_19183,N_19710);
nor U22457 (N_22457,N_18509,N_19772);
nor U22458 (N_22458,N_18615,N_17662);
nand U22459 (N_22459,N_19525,N_19870);
nand U22460 (N_22460,N_18460,N_19714);
nor U22461 (N_22461,N_19198,N_18978);
or U22462 (N_22462,N_18665,N_18791);
xor U22463 (N_22463,N_17808,N_17899);
nand U22464 (N_22464,N_17681,N_18993);
nor U22465 (N_22465,N_18076,N_19041);
nand U22466 (N_22466,N_19713,N_19165);
or U22467 (N_22467,N_19439,N_19408);
and U22468 (N_22468,N_17750,N_17961);
or U22469 (N_22469,N_17899,N_18405);
or U22470 (N_22470,N_18972,N_18784);
or U22471 (N_22471,N_18800,N_18549);
xnor U22472 (N_22472,N_18716,N_19097);
xor U22473 (N_22473,N_18397,N_19398);
nand U22474 (N_22474,N_19673,N_18368);
and U22475 (N_22475,N_18327,N_17984);
nand U22476 (N_22476,N_19669,N_17597);
nor U22477 (N_22477,N_19223,N_18096);
or U22478 (N_22478,N_19312,N_19151);
or U22479 (N_22479,N_17745,N_19570);
xor U22480 (N_22480,N_18205,N_19710);
and U22481 (N_22481,N_18774,N_17873);
and U22482 (N_22482,N_19775,N_18799);
nand U22483 (N_22483,N_18759,N_18975);
or U22484 (N_22484,N_18369,N_17617);
and U22485 (N_22485,N_19279,N_18325);
nor U22486 (N_22486,N_18613,N_18814);
nand U22487 (N_22487,N_18415,N_19705);
or U22488 (N_22488,N_18876,N_17801);
or U22489 (N_22489,N_19924,N_19565);
and U22490 (N_22490,N_17798,N_17584);
nor U22491 (N_22491,N_18631,N_17545);
nand U22492 (N_22492,N_19712,N_17592);
nor U22493 (N_22493,N_19276,N_18250);
and U22494 (N_22494,N_19857,N_18758);
or U22495 (N_22495,N_18737,N_17986);
nor U22496 (N_22496,N_19776,N_19815);
and U22497 (N_22497,N_17946,N_18004);
or U22498 (N_22498,N_17514,N_17737);
or U22499 (N_22499,N_19888,N_19426);
xor U22500 (N_22500,N_20996,N_22352);
and U22501 (N_22501,N_20814,N_20526);
nand U22502 (N_22502,N_22070,N_21377);
nand U22503 (N_22503,N_20175,N_20945);
and U22504 (N_22504,N_22386,N_22321);
and U22505 (N_22505,N_20759,N_20829);
nand U22506 (N_22506,N_20582,N_22219);
or U22507 (N_22507,N_22283,N_21198);
or U22508 (N_22508,N_21858,N_20736);
nor U22509 (N_22509,N_22005,N_20283);
nor U22510 (N_22510,N_20568,N_21227);
xnor U22511 (N_22511,N_22054,N_21445);
nand U22512 (N_22512,N_20264,N_20366);
nand U22513 (N_22513,N_21717,N_20978);
xor U22514 (N_22514,N_20321,N_20145);
xnor U22515 (N_22515,N_20427,N_21658);
nand U22516 (N_22516,N_22017,N_20190);
nor U22517 (N_22517,N_21973,N_21228);
nand U22518 (N_22518,N_21213,N_20623);
and U22519 (N_22519,N_21698,N_21631);
or U22520 (N_22520,N_20154,N_21331);
xor U22521 (N_22521,N_21687,N_22039);
and U22522 (N_22522,N_21914,N_21723);
or U22523 (N_22523,N_20198,N_21451);
nor U22524 (N_22524,N_22072,N_21417);
nor U22525 (N_22525,N_21525,N_21839);
nand U22526 (N_22526,N_22288,N_20870);
or U22527 (N_22527,N_21849,N_22163);
nor U22528 (N_22528,N_21260,N_21838);
nand U22529 (N_22529,N_21581,N_21813);
or U22530 (N_22530,N_22284,N_22200);
nand U22531 (N_22531,N_20450,N_21767);
and U22532 (N_22532,N_20386,N_20948);
nor U22533 (N_22533,N_20312,N_21645);
xnor U22534 (N_22534,N_22271,N_20776);
nor U22535 (N_22535,N_21959,N_21514);
nand U22536 (N_22536,N_22334,N_21237);
or U22537 (N_22537,N_21828,N_21616);
or U22538 (N_22538,N_20749,N_20362);
and U22539 (N_22539,N_20067,N_20635);
or U22540 (N_22540,N_21136,N_21335);
xor U22541 (N_22541,N_20871,N_20713);
nand U22542 (N_22542,N_20303,N_22104);
and U22543 (N_22543,N_22137,N_21899);
nand U22544 (N_22544,N_22165,N_22216);
and U22545 (N_22545,N_22096,N_20624);
xor U22546 (N_22546,N_20464,N_21502);
or U22547 (N_22547,N_20345,N_20525);
and U22548 (N_22548,N_21062,N_20114);
nand U22549 (N_22549,N_21909,N_20703);
nor U22550 (N_22550,N_20798,N_22375);
xor U22551 (N_22551,N_21425,N_21726);
and U22552 (N_22552,N_20886,N_22304);
and U22553 (N_22553,N_20878,N_22022);
and U22554 (N_22554,N_20531,N_20295);
nand U22555 (N_22555,N_21665,N_21216);
nor U22556 (N_22556,N_21883,N_21326);
nor U22557 (N_22557,N_21463,N_21366);
nor U22558 (N_22558,N_20520,N_22045);
or U22559 (N_22559,N_21346,N_22437);
or U22560 (N_22560,N_20664,N_21117);
xnor U22561 (N_22561,N_21479,N_21499);
nand U22562 (N_22562,N_20758,N_22019);
xor U22563 (N_22563,N_22217,N_21403);
nand U22564 (N_22564,N_20428,N_21952);
nor U22565 (N_22565,N_20921,N_21755);
nor U22566 (N_22566,N_20355,N_20769);
nand U22567 (N_22567,N_20816,N_22139);
xnor U22568 (N_22568,N_21146,N_21236);
nand U22569 (N_22569,N_20002,N_21732);
xor U22570 (N_22570,N_21370,N_21742);
or U22571 (N_22571,N_20023,N_22004);
nand U22572 (N_22572,N_20139,N_20918);
and U22573 (N_22573,N_22348,N_20227);
nand U22574 (N_22574,N_21796,N_22394);
xor U22575 (N_22575,N_22023,N_21073);
nand U22576 (N_22576,N_22041,N_21411);
and U22577 (N_22577,N_21513,N_20044);
and U22578 (N_22578,N_20266,N_21476);
nor U22579 (N_22579,N_20509,N_21416);
nor U22580 (N_22580,N_21811,N_21148);
and U22581 (N_22581,N_20113,N_21162);
nand U22582 (N_22582,N_21786,N_22097);
and U22583 (N_22583,N_20179,N_21399);
or U22584 (N_22584,N_21298,N_20107);
nor U22585 (N_22585,N_20939,N_20319);
and U22586 (N_22586,N_20043,N_21307);
and U22587 (N_22587,N_22393,N_21946);
xor U22588 (N_22588,N_20208,N_21275);
nand U22589 (N_22589,N_20533,N_20108);
and U22590 (N_22590,N_20731,N_20835);
xor U22591 (N_22591,N_21409,N_21611);
nor U22592 (N_22592,N_22310,N_20923);
nor U22593 (N_22593,N_21894,N_20066);
or U22594 (N_22594,N_22114,N_21106);
or U22595 (N_22595,N_21531,N_20708);
nor U22596 (N_22596,N_20318,N_20560);
nor U22597 (N_22597,N_21803,N_22002);
or U22598 (N_22598,N_20964,N_21240);
and U22599 (N_22599,N_21563,N_20074);
xor U22600 (N_22600,N_20785,N_21745);
and U22601 (N_22601,N_20467,N_21920);
xnor U22602 (N_22602,N_21270,N_20137);
nand U22603 (N_22603,N_22102,N_20022);
xnor U22604 (N_22604,N_20183,N_21699);
and U22605 (N_22605,N_21972,N_22349);
and U22606 (N_22606,N_21245,N_22392);
nor U22607 (N_22607,N_20342,N_20550);
nand U22608 (N_22608,N_20609,N_20593);
nand U22609 (N_22609,N_20688,N_20005);
nand U22610 (N_22610,N_20647,N_22444);
xnor U22611 (N_22611,N_20129,N_20439);
nand U22612 (N_22612,N_21390,N_20955);
or U22613 (N_22613,N_20670,N_20608);
and U22614 (N_22614,N_20577,N_21814);
nand U22615 (N_22615,N_20810,N_22182);
or U22616 (N_22616,N_22178,N_21327);
or U22617 (N_22617,N_20984,N_20262);
xnor U22618 (N_22618,N_21166,N_21781);
and U22619 (N_22619,N_21915,N_20191);
nor U22620 (N_22620,N_21540,N_22308);
or U22621 (N_22621,N_22043,N_22458);
and U22622 (N_22622,N_21364,N_20335);
nand U22623 (N_22623,N_20363,N_21992);
xnor U22624 (N_22624,N_21931,N_20414);
nor U22625 (N_22625,N_21321,N_21614);
or U22626 (N_22626,N_20625,N_20028);
nand U22627 (N_22627,N_21780,N_21837);
and U22628 (N_22628,N_21217,N_22330);
and U22629 (N_22629,N_21609,N_22249);
nor U22630 (N_22630,N_20979,N_21765);
nand U22631 (N_22631,N_22235,N_21944);
and U22632 (N_22632,N_21273,N_21483);
or U22633 (N_22633,N_21398,N_20844);
and U22634 (N_22634,N_21109,N_20828);
nand U22635 (N_22635,N_20837,N_20725);
and U22636 (N_22636,N_20395,N_22478);
or U22637 (N_22637,N_22229,N_21963);
nor U22638 (N_22638,N_20834,N_20443);
nor U22639 (N_22639,N_21473,N_21646);
xor U22640 (N_22640,N_22058,N_22068);
nand U22641 (N_22641,N_22332,N_20019);
or U22642 (N_22642,N_20867,N_21223);
and U22643 (N_22643,N_21913,N_20890);
nand U22644 (N_22644,N_21529,N_20899);
nand U22645 (N_22645,N_21209,N_21748);
or U22646 (N_22646,N_21594,N_21075);
nand U22647 (N_22647,N_20633,N_21577);
and U22648 (N_22648,N_22358,N_21902);
nor U22649 (N_22649,N_21116,N_21674);
and U22650 (N_22650,N_22107,N_22177);
nor U22651 (N_22651,N_21661,N_21640);
or U22652 (N_22652,N_21842,N_21739);
nor U22653 (N_22653,N_22242,N_20528);
xor U22654 (N_22654,N_20046,N_21940);
nand U22655 (N_22655,N_22014,N_20212);
and U22656 (N_22656,N_21657,N_21941);
nor U22657 (N_22657,N_21664,N_22048);
xor U22658 (N_22658,N_20275,N_22300);
nor U22659 (N_22659,N_22465,N_21741);
xor U22660 (N_22660,N_20151,N_20185);
or U22661 (N_22661,N_22250,N_22038);
xor U22662 (N_22662,N_21979,N_21468);
nand U22663 (N_22663,N_21857,N_20135);
xor U22664 (N_22664,N_21266,N_21504);
nand U22665 (N_22665,N_21666,N_22422);
nor U22666 (N_22666,N_21045,N_21904);
xnor U22667 (N_22667,N_21945,N_21265);
nor U22668 (N_22668,N_20910,N_21309);
xnor U22669 (N_22669,N_22479,N_21010);
nor U22670 (N_22670,N_22150,N_20279);
xor U22671 (N_22671,N_22088,N_20237);
and U22672 (N_22672,N_20281,N_21603);
nand U22673 (N_22673,N_22003,N_20289);
xor U22674 (N_22674,N_22320,N_20874);
xnor U22675 (N_22675,N_21703,N_22362);
or U22676 (N_22676,N_21200,N_21668);
nand U22677 (N_22677,N_20308,N_22035);
xnor U22678 (N_22678,N_21402,N_22359);
xnor U22679 (N_22679,N_21597,N_22335);
xnor U22680 (N_22680,N_20296,N_22448);
xnor U22681 (N_22681,N_22383,N_22476);
or U22682 (N_22682,N_22025,N_22469);
or U22683 (N_22683,N_20375,N_22248);
and U22684 (N_22684,N_21080,N_20174);
and U22685 (N_22685,N_21926,N_21608);
nand U22686 (N_22686,N_21874,N_21546);
and U22687 (N_22687,N_20478,N_20203);
nand U22688 (N_22688,N_20906,N_22273);
xor U22689 (N_22689,N_20196,N_20681);
nor U22690 (N_22690,N_20573,N_22236);
and U22691 (N_22691,N_20711,N_20062);
xnor U22692 (N_22692,N_20805,N_21845);
and U22693 (N_22693,N_20990,N_20305);
nand U22694 (N_22694,N_22000,N_20150);
nor U22695 (N_22695,N_21675,N_22326);
nor U22696 (N_22696,N_22261,N_21610);
xor U22697 (N_22697,N_22255,N_20441);
or U22698 (N_22698,N_21547,N_20869);
xnor U22699 (N_22699,N_21667,N_21362);
nand U22700 (N_22700,N_21287,N_22001);
nand U22701 (N_22701,N_21113,N_20447);
xor U22702 (N_22702,N_21482,N_21450);
nor U22703 (N_22703,N_21636,N_21983);
nor U22704 (N_22704,N_20434,N_21691);
or U22705 (N_22705,N_22067,N_22061);
nand U22706 (N_22706,N_21255,N_20340);
nand U22707 (N_22707,N_20425,N_20142);
xor U22708 (N_22708,N_20314,N_21406);
and U22709 (N_22709,N_20784,N_22403);
nand U22710 (N_22710,N_21069,N_21215);
xor U22711 (N_22711,N_20975,N_20592);
and U22712 (N_22712,N_21981,N_20740);
or U22713 (N_22713,N_20039,N_20501);
or U22714 (N_22714,N_22312,N_20494);
or U22715 (N_22715,N_20463,N_22237);
nand U22716 (N_22716,N_20544,N_20933);
nand U22717 (N_22717,N_20802,N_21258);
nand U22718 (N_22718,N_21143,N_20796);
xor U22719 (N_22719,N_21163,N_21026);
nand U22720 (N_22720,N_21334,N_22474);
nand U22721 (N_22721,N_22207,N_21555);
nor U22722 (N_22722,N_21179,N_21071);
or U22723 (N_22723,N_22008,N_21624);
xor U22724 (N_22724,N_22034,N_21836);
and U22725 (N_22725,N_21960,N_20457);
or U22726 (N_22726,N_21787,N_21772);
nor U22727 (N_22727,N_20104,N_20376);
xnor U22728 (N_22728,N_22186,N_22057);
or U22729 (N_22729,N_21068,N_21271);
and U22730 (N_22730,N_21413,N_20885);
xor U22731 (N_22731,N_21040,N_20106);
nand U22732 (N_22732,N_21696,N_20205);
nor U22733 (N_22733,N_22099,N_21617);
and U22734 (N_22734,N_21683,N_20671);
nor U22735 (N_22735,N_21011,N_21572);
or U22736 (N_22736,N_20089,N_20707);
and U22737 (N_22737,N_21776,N_20685);
or U22738 (N_22738,N_20881,N_22292);
or U22739 (N_22739,N_20596,N_20686);
or U22740 (N_22740,N_22077,N_20604);
and U22741 (N_22741,N_21369,N_21191);
or U22742 (N_22742,N_22103,N_22372);
and U22743 (N_22743,N_21853,N_21596);
nor U22744 (N_22744,N_20995,N_21028);
nor U22745 (N_22745,N_21908,N_22371);
xor U22746 (N_22746,N_21170,N_20390);
and U22747 (N_22747,N_20513,N_21986);
or U22748 (N_22748,N_22342,N_21873);
and U22749 (N_22749,N_20717,N_21176);
nand U22750 (N_22750,N_20638,N_22244);
nand U22751 (N_22751,N_21840,N_21243);
or U22752 (N_22752,N_21322,N_21936);
xor U22753 (N_22753,N_20291,N_20288);
nor U22754 (N_22754,N_21344,N_22056);
nor U22755 (N_22755,N_20547,N_21269);
nor U22756 (N_22756,N_20620,N_20585);
nand U22757 (N_22757,N_22351,N_20859);
or U22758 (N_22758,N_20977,N_22411);
and U22759 (N_22759,N_20093,N_20158);
nand U22760 (N_22760,N_21948,N_20284);
nand U22761 (N_22761,N_21281,N_20430);
nor U22762 (N_22762,N_20863,N_21249);
xor U22763 (N_22763,N_21202,N_21194);
or U22764 (N_22764,N_20627,N_20925);
nand U22765 (N_22765,N_21893,N_20721);
xnor U22766 (N_22766,N_20591,N_21141);
nand U22767 (N_22767,N_20639,N_21112);
or U22768 (N_22768,N_20256,N_20141);
nand U22769 (N_22769,N_20897,N_21521);
nor U22770 (N_22770,N_20167,N_22282);
or U22771 (N_22771,N_21353,N_20613);
or U22772 (N_22772,N_22108,N_20389);
xnor U22773 (N_22773,N_20020,N_21711);
or U22774 (N_22774,N_20187,N_20770);
nor U22775 (N_22775,N_20619,N_21193);
nor U22776 (N_22776,N_20879,N_22029);
nand U22777 (N_22777,N_20603,N_22203);
nand U22778 (N_22778,N_20241,N_21349);
or U22779 (N_22779,N_21005,N_21092);
and U22780 (N_22780,N_20887,N_21918);
nand U22781 (N_22781,N_22126,N_21239);
and U22782 (N_22782,N_21804,N_21889);
or U22783 (N_22783,N_21312,N_21890);
or U22784 (N_22784,N_20912,N_22280);
xor U22785 (N_22785,N_22353,N_20626);
nor U22786 (N_22786,N_22460,N_22260);
and U22787 (N_22787,N_20157,N_21456);
or U22788 (N_22788,N_22245,N_21537);
or U22789 (N_22789,N_20667,N_20570);
and U22790 (N_22790,N_22129,N_21430);
nand U22791 (N_22791,N_20941,N_20750);
nand U22792 (N_22792,N_21713,N_21144);
xnor U22793 (N_22793,N_20644,N_21410);
nor U22794 (N_22794,N_20407,N_21458);
or U22795 (N_22795,N_21190,N_20850);
nor U22796 (N_22796,N_20722,N_20426);
nor U22797 (N_22797,N_20220,N_22286);
nor U22798 (N_22798,N_22291,N_20417);
or U22799 (N_22799,N_20460,N_22339);
nor U22800 (N_22800,N_20148,N_22447);
nand U22801 (N_22801,N_20254,N_20373);
xor U22802 (N_22802,N_20579,N_20502);
nor U22803 (N_22803,N_21051,N_20696);
xnor U22804 (N_22804,N_21851,N_20399);
or U22805 (N_22805,N_20632,N_20492);
nor U22806 (N_22806,N_20041,N_20586);
nor U22807 (N_22807,N_20383,N_21330);
xor U22808 (N_22808,N_21522,N_20689);
and U22809 (N_22809,N_22454,N_20301);
nand U22810 (N_22810,N_21001,N_20915);
and U22811 (N_22811,N_21488,N_22269);
or U22812 (N_22812,N_21137,N_22376);
xnor U22813 (N_22813,N_22445,N_20495);
nand U22814 (N_22814,N_20919,N_21453);
xnor U22815 (N_22815,N_21046,N_21881);
xor U22816 (N_22816,N_21622,N_22162);
nor U22817 (N_22817,N_21048,N_22153);
nand U22818 (N_22818,N_21098,N_22272);
and U22819 (N_22819,N_22031,N_20052);
or U22820 (N_22820,N_20672,N_21880);
xnor U22821 (N_22821,N_22404,N_21961);
nand U22822 (N_22822,N_20893,N_21434);
nor U22823 (N_22823,N_21626,N_20068);
or U22824 (N_22824,N_21724,N_20669);
and U22825 (N_22825,N_20000,N_20432);
xnor U22826 (N_22826,N_20600,N_20300);
nor U22827 (N_22827,N_20214,N_21279);
xor U22828 (N_22828,N_21559,N_22184);
nand U22829 (N_22829,N_22489,N_22477);
nand U22830 (N_22830,N_20133,N_21274);
nand U22831 (N_22831,N_22256,N_21388);
xnor U22832 (N_22832,N_21511,N_20377);
xor U22833 (N_22833,N_21774,N_21077);
nand U22834 (N_22834,N_20905,N_20246);
or U22835 (N_22835,N_21440,N_20599);
nand U22836 (N_22836,N_20775,N_21865);
nor U22837 (N_22837,N_20815,N_20987);
nand U22838 (N_22838,N_21498,N_21160);
nand U22839 (N_22839,N_22081,N_20116);
nand U22840 (N_22840,N_20841,N_22055);
nand U22841 (N_22841,N_20690,N_20752);
and U22842 (N_22842,N_20204,N_21916);
xor U22843 (N_22843,N_21167,N_20665);
or U22844 (N_22844,N_20315,N_21588);
or U22845 (N_22845,N_20287,N_21999);
or U22846 (N_22846,N_21474,N_21494);
and U22847 (N_22847,N_21705,N_20827);
nand U22848 (N_22848,N_22384,N_21182);
and U22849 (N_22849,N_21714,N_21431);
and U22850 (N_22850,N_21731,N_21013);
xnor U22851 (N_22851,N_22136,N_20602);
xor U22852 (N_22852,N_21812,N_20372);
and U22853 (N_22853,N_21805,N_20883);
xnor U22854 (N_22854,N_22295,N_21980);
xnor U22855 (N_22855,N_22487,N_20349);
nand U22856 (N_22856,N_22427,N_22241);
nor U22857 (N_22857,N_21517,N_21910);
and U22858 (N_22858,N_21574,N_21878);
or U22859 (N_22859,N_21058,N_21937);
nor U22860 (N_22860,N_22398,N_22264);
or U22861 (N_22861,N_21676,N_21497);
and U22862 (N_22862,N_22080,N_21820);
or U22863 (N_22863,N_22125,N_20419);
and U22864 (N_22864,N_21489,N_20452);
or U22865 (N_22865,N_21593,N_20038);
nor U22866 (N_22866,N_21565,N_21448);
xor U22867 (N_22867,N_21435,N_21746);
nand U22868 (N_22868,N_21222,N_21740);
xor U22869 (N_22869,N_22278,N_21201);
nor U22870 (N_22870,N_22197,N_21997);
nand U22871 (N_22871,N_20343,N_20476);
nand U22872 (N_22872,N_22231,N_21022);
xor U22873 (N_22873,N_21462,N_22052);
or U22874 (N_22874,N_21817,N_21464);
nor U22875 (N_22875,N_21442,N_20763);
and U22876 (N_22876,N_22410,N_22075);
or U22877 (N_22877,N_20817,N_20851);
xnor U22878 (N_22878,N_22144,N_20011);
nor U22879 (N_22879,N_20496,N_21523);
nand U22880 (N_22880,N_22305,N_20225);
or U22881 (N_22881,N_22463,N_20206);
xor U22882 (N_22882,N_22434,N_21292);
or U22883 (N_22883,N_22306,N_21949);
nor U22884 (N_22884,N_22311,N_21380);
nand U22885 (N_22885,N_20192,N_20292);
nor U22886 (N_22886,N_21354,N_22322);
or U22887 (N_22887,N_22324,N_20967);
nand U22888 (N_22888,N_20265,N_20741);
and U22889 (N_22889,N_21418,N_22405);
and U22890 (N_22890,N_21066,N_21841);
xor U22891 (N_22891,N_20566,N_22105);
xnor U22892 (N_22892,N_21998,N_20849);
nor U22893 (N_22893,N_21756,N_20551);
nor U22894 (N_22894,N_21911,N_21278);
nand U22895 (N_22895,N_20199,N_22363);
nor U22896 (N_22896,N_21184,N_20073);
xnor U22897 (N_22897,N_21050,N_21340);
nand U22898 (N_22898,N_21969,N_21304);
or U22899 (N_22899,N_21671,N_20025);
nor U22900 (N_22900,N_20037,N_20569);
xnor U22901 (N_22901,N_21719,N_20976);
or U22902 (N_22902,N_20486,N_21782);
and U22903 (N_22903,N_21749,N_20221);
or U22904 (N_22904,N_20917,N_21181);
nand U22905 (N_22905,N_21564,N_21103);
nor U22906 (N_22906,N_21656,N_20127);
nand U22907 (N_22907,N_21082,N_21528);
or U22908 (N_22908,N_20224,N_21807);
and U22909 (N_22909,N_20306,N_20488);
nor U22910 (N_22910,N_22147,N_22373);
nand U22911 (N_22911,N_20747,N_21306);
nor U22912 (N_22912,N_20705,N_21041);
and U22913 (N_22913,N_20401,N_21871);
or U22914 (N_22914,N_22166,N_21449);
xnor U22915 (N_22915,N_20103,N_20554);
nor U22916 (N_22916,N_21018,N_20251);
nand U22917 (N_22917,N_21283,N_21175);
xor U22918 (N_22918,N_21342,N_21568);
nand U22919 (N_22919,N_22227,N_20954);
nor U22920 (N_22920,N_20209,N_21233);
or U22921 (N_22921,N_21284,N_21690);
or U22922 (N_22922,N_21925,N_20821);
xor U22923 (N_22923,N_21538,N_21548);
nor U22924 (N_22924,N_21996,N_22344);
nand U22925 (N_22925,N_22254,N_20963);
nor U22926 (N_22926,N_21466,N_21150);
or U22927 (N_22927,N_21688,N_20553);
xnor U22928 (N_22928,N_21230,N_21131);
nand U22929 (N_22929,N_22268,N_21373);
nand U22930 (N_22930,N_22111,N_20244);
or U22931 (N_22931,N_20404,N_22095);
or U22932 (N_22932,N_22079,N_22356);
nor U22933 (N_22933,N_21171,N_20847);
or U22934 (N_22934,N_21766,N_21316);
nor U22935 (N_22935,N_21487,N_20369);
xnor U22936 (N_22936,N_20197,N_20971);
or U22937 (N_22937,N_22154,N_21095);
and U22938 (N_22938,N_22180,N_21024);
nor U22939 (N_22939,N_21951,N_21800);
nand U22940 (N_22940,N_21052,N_20822);
and U22941 (N_22941,N_21437,N_20410);
xnor U22942 (N_22942,N_20413,N_20588);
nor U22943 (N_22943,N_21552,N_22316);
xor U22944 (N_22944,N_20666,N_21056);
or U22945 (N_22945,N_22194,N_22090);
or U22946 (N_22946,N_20008,N_22436);
or U22947 (N_22947,N_22360,N_20911);
xnor U22948 (N_22948,N_21180,N_21947);
and U22949 (N_22949,N_20538,N_21161);
nor U22950 (N_22950,N_22262,N_22408);
or U22951 (N_22951,N_20615,N_21734);
and U22952 (N_22952,N_20048,N_21467);
and U22953 (N_22953,N_21738,N_20218);
xnor U22954 (N_22954,N_20571,N_22119);
nor U22955 (N_22955,N_20248,N_21672);
and U22956 (N_22956,N_21130,N_22085);
and U22957 (N_22957,N_20642,N_20200);
and U22958 (N_22958,N_21900,N_20004);
nor U22959 (N_22959,N_20966,N_21519);
and U22960 (N_22960,N_20641,N_20812);
or U22961 (N_22961,N_21185,N_21029);
and U22962 (N_22962,N_20493,N_22382);
and U22963 (N_22963,N_20807,N_20969);
or U22964 (N_22964,N_21345,N_20012);
nand U22965 (N_22965,N_21267,N_20344);
nand U22966 (N_22966,N_20272,N_21361);
nand U22967 (N_22967,N_20445,N_22497);
nor U22968 (N_22968,N_20764,N_21085);
and U22969 (N_22969,N_20354,N_20347);
xnor U22970 (N_22970,N_21427,N_20422);
and U22971 (N_22971,N_21653,N_22205);
and U22972 (N_22972,N_21114,N_20147);
or U22973 (N_22973,N_22457,N_21833);
xnor U22974 (N_22974,N_21825,N_20622);
nand U22975 (N_22975,N_20235,N_20247);
nor U22976 (N_22976,N_21806,N_22233);
and U22977 (N_22977,N_21987,N_20333);
and U22978 (N_22978,N_21660,N_20660);
and U22979 (N_22979,N_20574,N_21509);
and U22980 (N_22980,N_21632,N_21589);
nor U22981 (N_22981,N_20115,N_21966);
and U22982 (N_22982,N_21432,N_21967);
nor U22983 (N_22983,N_20781,N_21072);
nor U22984 (N_22984,N_20085,N_21244);
and U22985 (N_22985,N_21207,N_21587);
or U22986 (N_22986,N_20131,N_20676);
xnor U22987 (N_22987,N_21633,N_20732);
and U22988 (N_22988,N_20030,N_20448);
and U22989 (N_22989,N_21128,N_22201);
and U22990 (N_22990,N_21855,N_21280);
and U22991 (N_22991,N_22430,N_21950);
nor U22992 (N_22992,N_22073,N_20238);
nand U22993 (N_22993,N_22395,N_21580);
nor U22994 (N_22994,N_20324,N_21753);
xor U22995 (N_22995,N_20331,N_20719);
nand U22996 (N_22996,N_21197,N_22396);
nor U22997 (N_22997,N_22263,N_20216);
nor U22998 (N_22998,N_20437,N_21367);
xor U22999 (N_22999,N_20500,N_20485);
xor U23000 (N_23000,N_21879,N_21002);
nor U23001 (N_23001,N_21752,N_20779);
xor U23002 (N_23002,N_21219,N_22228);
nor U23003 (N_23003,N_21628,N_20534);
nor U23004 (N_23004,N_20589,N_20138);
and U23005 (N_23005,N_21481,N_22199);
xnor U23006 (N_23006,N_20724,N_22115);
xnor U23007 (N_23007,N_20972,N_21769);
or U23008 (N_23008,N_21870,N_20612);
or U23009 (N_23009,N_21682,N_20506);
xor U23010 (N_23010,N_21484,N_21534);
or U23011 (N_23011,N_20078,N_22234);
xnor U23012 (N_23012,N_20510,N_21921);
xor U23013 (N_23013,N_20675,N_21199);
xor U23014 (N_23014,N_22007,N_20015);
xor U23015 (N_23015,N_20845,N_20746);
nand U23016 (N_23016,N_20310,N_20226);
and U23017 (N_23017,N_21108,N_21599);
nand U23018 (N_23018,N_22499,N_21195);
or U23019 (N_23019,N_22062,N_20188);
nand U23020 (N_23020,N_22490,N_21063);
nor U23021 (N_23021,N_20800,N_22049);
or U23022 (N_23022,N_20516,N_22076);
xnor U23023 (N_23023,N_22270,N_20356);
xnor U23024 (N_23024,N_20367,N_20146);
and U23025 (N_23025,N_20514,N_22141);
nor U23026 (N_23026,N_20455,N_21794);
and U23027 (N_23027,N_22148,N_20999);
and U23028 (N_23028,N_20490,N_21567);
nand U23029 (N_23029,N_21037,N_20839);
or U23030 (N_23030,N_21384,N_22467);
nor U23031 (N_23031,N_22093,N_21810);
xor U23032 (N_23032,N_20580,N_21212);
and U23033 (N_23033,N_21365,N_21093);
nand U23034 (N_23034,N_20710,N_20018);
or U23035 (N_23035,N_20162,N_20338);
nor U23036 (N_23036,N_21654,N_20105);
nor U23037 (N_23037,N_21428,N_21635);
nand U23038 (N_23038,N_20403,N_20692);
or U23039 (N_23039,N_20332,N_22415);
nor U23040 (N_23040,N_20253,N_20014);
xnor U23041 (N_23041,N_20121,N_21604);
or U23042 (N_23042,N_21120,N_21272);
nor U23043 (N_23043,N_21897,N_22323);
and U23044 (N_23044,N_21027,N_21892);
and U23045 (N_23045,N_21697,N_20801);
and U23046 (N_23046,N_21070,N_21964);
xnor U23047 (N_23047,N_21721,N_20236);
nand U23048 (N_23048,N_20536,N_22494);
nor U23049 (N_23049,N_21332,N_20359);
xnor U23050 (N_23050,N_20090,N_22258);
and U23051 (N_23051,N_21206,N_20650);
xor U23052 (N_23052,N_20959,N_20962);
xor U23053 (N_23053,N_21057,N_22368);
nand U23054 (N_23054,N_20583,N_22220);
nand U23055 (N_23055,N_21186,N_22317);
nand U23056 (N_23056,N_21470,N_20695);
nor U23057 (N_23057,N_21263,N_22143);
xor U23058 (N_23058,N_21573,N_21701);
nand U23059 (N_23059,N_20313,N_22401);
or U23060 (N_23060,N_20584,N_20405);
and U23061 (N_23061,N_21562,N_20637);
xor U23062 (N_23062,N_20257,N_21295);
or U23063 (N_23063,N_21832,N_20512);
or U23064 (N_23064,N_20679,N_21720);
nand U23065 (N_23065,N_21627,N_21076);
nor U23066 (N_23066,N_20738,N_21324);
nand U23067 (N_23067,N_20143,N_20791);
xor U23068 (N_23068,N_21135,N_21030);
and U23069 (N_23069,N_21895,N_22350);
xnor U23070 (N_23070,N_20940,N_22021);
and U23071 (N_23071,N_21798,N_20128);
xnor U23072 (N_23072,N_21457,N_22071);
xnor U23073 (N_23073,N_21429,N_20652);
or U23074 (N_23074,N_22202,N_21715);
and U23075 (N_23075,N_20271,N_21877);
and U23076 (N_23076,N_20704,N_22206);
or U23077 (N_23077,N_22377,N_22390);
and U23078 (N_23078,N_21039,N_20709);
or U23079 (N_23079,N_20843,N_21294);
nor U23080 (N_23080,N_21606,N_21355);
and U23081 (N_23081,N_20755,N_20140);
and U23082 (N_23082,N_20875,N_21530);
or U23083 (N_23083,N_21578,N_20282);
or U23084 (N_23084,N_20595,N_22173);
and U23085 (N_23085,N_21882,N_20748);
and U23086 (N_23086,N_21704,N_21009);
nor U23087 (N_23087,N_21977,N_20891);
nor U23088 (N_23088,N_21225,N_21475);
and U23089 (N_23089,N_22328,N_21020);
and U23090 (N_23090,N_21939,N_20751);
nor U23091 (N_23091,N_20806,N_21360);
nor U23092 (N_23092,N_22400,N_21031);
and U23093 (N_23093,N_21495,N_20617);
xnor U23094 (N_23094,N_20070,N_22016);
and U23095 (N_23095,N_21460,N_21712);
nand U23096 (N_23096,N_21907,N_21091);
nand U23097 (N_23097,N_20754,N_20350);
nor U23098 (N_23098,N_21145,N_21919);
nor U23099 (N_23099,N_22294,N_20013);
xnor U23100 (N_23100,N_21864,N_20575);
nor U23101 (N_23101,N_22122,N_21038);
or U23102 (N_23102,N_22195,N_22092);
or U23103 (N_23103,N_21764,N_20936);
or U23104 (N_23104,N_21571,N_21854);
nand U23105 (N_23105,N_21313,N_22414);
nand U23106 (N_23106,N_21419,N_21134);
and U23107 (N_23107,N_20973,N_21935);
nor U23108 (N_23108,N_20491,N_21679);
or U23109 (N_23109,N_21081,N_21993);
xor U23110 (N_23110,N_20122,N_21550);
and U23111 (N_23111,N_20986,N_22232);
xor U23112 (N_23112,N_21337,N_21680);
nor U23113 (N_23113,N_20461,N_22425);
xnor U23114 (N_23114,N_22087,N_22452);
nor U23115 (N_23115,N_21097,N_21984);
or U23116 (N_23116,N_21455,N_20280);
or U23117 (N_23117,N_21681,N_22006);
xnor U23118 (N_23118,N_20032,N_20507);
xor U23119 (N_23119,N_22296,N_21142);
xor U23120 (N_23120,N_21750,N_21693);
nand U23121 (N_23121,N_21084,N_20123);
and U23122 (N_23122,N_21863,N_21507);
and U23123 (N_23123,N_21592,N_20339);
xor U23124 (N_23124,N_22208,N_22307);
xor U23125 (N_23125,N_21543,N_21709);
nand U23126 (N_23126,N_20927,N_20952);
nand U23127 (N_23127,N_21043,N_22413);
xor U23128 (N_23128,N_21382,N_22484);
nand U23129 (N_23129,N_20673,N_22127);
nand U23130 (N_23130,N_22406,N_22492);
and U23131 (N_23131,N_22024,N_22337);
xnor U23132 (N_23132,N_21105,N_20680);
xnor U23133 (N_23133,N_20657,N_20866);
and U23134 (N_23134,N_22433,N_21922);
nand U23135 (N_23135,N_21358,N_20483);
nor U23136 (N_23136,N_21644,N_20346);
nor U23137 (N_23137,N_20854,N_20868);
and U23138 (N_23138,N_20654,N_20826);
xor U23139 (N_23139,N_21107,N_21025);
nor U23140 (N_23140,N_21778,N_20273);
xnor U23141 (N_23141,N_22106,N_20130);
nor U23142 (N_23142,N_21485,N_20700);
nor U23143 (N_23143,N_22419,N_21634);
or U23144 (N_23144,N_20079,N_22329);
xnor U23145 (N_23145,N_21859,N_22252);
or U23146 (N_23146,N_20698,N_21843);
and U23147 (N_23147,N_20371,N_20440);
nand U23148 (N_23148,N_21503,N_21318);
xnor U23149 (N_23149,N_21770,N_21439);
xnor U23150 (N_23150,N_21183,N_21338);
nand U23151 (N_23151,N_21042,N_20756);
nand U23152 (N_23152,N_22428,N_21516);
nand U23153 (N_23153,N_21139,N_20031);
nand U23154 (N_23154,N_20396,N_22179);
xnor U23155 (N_23155,N_22462,N_20097);
nand U23156 (N_23156,N_20436,N_22407);
nor U23157 (N_23157,N_22379,N_22482);
or U23158 (N_23158,N_21823,N_21735);
and U23159 (N_23159,N_21788,N_20605);
nor U23160 (N_23160,N_20161,N_21618);
and U23161 (N_23161,N_21591,N_20982);
xor U23162 (N_23162,N_20683,N_21196);
or U23163 (N_23163,N_22120,N_21722);
and U23164 (N_23164,N_21310,N_20341);
nand U23165 (N_23165,N_20454,N_20518);
nand U23166 (N_23166,N_21831,N_22446);
nand U23167 (N_23167,N_20329,N_21971);
or U23168 (N_23168,N_21924,N_22149);
xnor U23169 (N_23169,N_21586,N_22060);
and U23170 (N_23170,N_20558,N_21637);
nor U23171 (N_23171,N_22481,N_20112);
nor U23172 (N_23172,N_20240,N_20092);
xnor U23173 (N_23173,N_22094,N_20076);
and U23174 (N_23174,N_20913,N_20471);
or U23175 (N_23175,N_21801,N_20922);
and U23176 (N_23176,N_22374,N_22211);
xnor U23177 (N_23177,N_20239,N_21536);
xor U23178 (N_23178,N_22160,N_20678);
and U23179 (N_23179,N_22193,N_20920);
or U23180 (N_23180,N_20252,N_21965);
xor U23181 (N_23181,N_21102,N_22333);
xor U23182 (N_23182,N_21235,N_21422);
nand U23183 (N_23183,N_20578,N_20661);
nor U23184 (N_23184,N_21156,N_20294);
nor U23185 (N_23185,N_21446,N_21686);
or U23186 (N_23186,N_21395,N_22253);
xnor U23187 (N_23187,N_21300,N_21089);
nand U23188 (N_23188,N_20634,N_22089);
and U23189 (N_23189,N_20034,N_21829);
nand U23190 (N_23190,N_20616,N_22293);
nand U23191 (N_23191,N_20118,N_20388);
or U23192 (N_23192,N_20446,N_22370);
nor U23193 (N_23193,N_21518,N_21790);
nand U23194 (N_23194,N_20177,N_20640);
nor U23195 (N_23195,N_21575,N_21783);
nand U23196 (N_23196,N_22069,N_21234);
xnor U23197 (N_23197,N_21898,N_21157);
or U23198 (N_23198,N_20409,N_20249);
nand U23199 (N_23199,N_21210,N_20336);
xor U23200 (N_23200,N_22276,N_20572);
xor U23201 (N_23201,N_21158,N_21876);
nand U23202 (N_23202,N_20047,N_21343);
xor U23203 (N_23203,N_21291,N_21133);
and U23204 (N_23204,N_21164,N_20864);
and U23205 (N_23205,N_21954,N_20957);
and U23206 (N_23206,N_20497,N_20900);
and U23207 (N_23207,N_21242,N_21702);
or U23208 (N_23208,N_20286,N_22461);
nor U23209 (N_23209,N_21647,N_21016);
and U23210 (N_23210,N_21584,N_20857);
xnor U23211 (N_23211,N_22417,N_21003);
nand U23212 (N_23212,N_21508,N_22140);
nor U23213 (N_23213,N_21869,N_21613);
and U23214 (N_23214,N_21775,N_20621);
or U23215 (N_23215,N_20487,N_21991);
and U23216 (N_23216,N_21426,N_21420);
and U23217 (N_23217,N_22064,N_21447);
nand U23218 (N_23218,N_20326,N_21505);
or U23219 (N_23219,N_21551,N_21743);
and U23220 (N_23220,N_22113,N_21598);
and U23221 (N_23221,N_21625,N_22498);
and U23222 (N_23222,N_20050,N_20521);
nor U23223 (N_23223,N_20958,N_20385);
nor U23224 (N_23224,N_20853,N_20223);
and U23225 (N_23225,N_20762,N_20610);
or U23226 (N_23226,N_21385,N_20803);
and U23227 (N_23227,N_21238,N_20479);
nor U23228 (N_23228,N_21669,N_20648);
or U23229 (N_23229,N_21371,N_21962);
nor U23230 (N_23230,N_21376,N_21861);
and U23231 (N_23231,N_20981,N_22485);
or U23232 (N_23232,N_22158,N_21884);
and U23233 (N_23233,N_21262,N_21761);
nand U23234 (N_23234,N_20484,N_21308);
nor U23235 (N_23235,N_20184,N_22218);
nor U23236 (N_23236,N_21760,N_20120);
or U23237 (N_23237,N_22145,N_20334);
nor U23238 (N_23238,N_21083,N_22385);
nor U23239 (N_23239,N_20646,N_20733);
xor U23240 (N_23240,N_20938,N_21621);
nor U23241 (N_23241,N_21314,N_20327);
nand U23242 (N_23242,N_20556,N_21465);
nand U23243 (N_23243,N_20029,N_20504);
nand U23244 (N_23244,N_20111,N_21491);
and U23245 (N_23245,N_21639,N_21506);
or U23246 (N_23246,N_22364,N_20086);
nand U23247 (N_23247,N_20387,N_21887);
or U23248 (N_23248,N_21968,N_20178);
xor U23249 (N_23249,N_21685,N_21023);
xor U23250 (N_23250,N_22033,N_21677);
or U23251 (N_23251,N_20459,N_20818);
and U23252 (N_23252,N_22409,N_21110);
nor U23253 (N_23253,N_21389,N_20777);
nor U23254 (N_23254,N_21566,N_21862);
nor U23255 (N_23255,N_21017,N_20049);
nand U23256 (N_23256,N_20472,N_20021);
or U23257 (N_23257,N_20993,N_21079);
nor U23258 (N_23258,N_20576,N_21320);
and U23259 (N_23259,N_22435,N_21477);
and U23260 (N_23260,N_21414,N_20559);
xnor U23261 (N_23261,N_22213,N_20003);
xnor U23262 (N_23262,N_20929,N_20475);
nor U23263 (N_23263,N_22161,N_22188);
nor U23264 (N_23264,N_21325,N_21652);
nor U23265 (N_23265,N_21736,N_20539);
nor U23266 (N_23266,N_20110,N_22109);
or U23267 (N_23267,N_21707,N_21459);
and U23268 (N_23268,N_20170,N_22313);
xnor U23269 (N_23269,N_21816,N_21121);
nor U23270 (N_23270,N_21988,N_20824);
and U23271 (N_23271,N_22083,N_22169);
nor U23272 (N_23272,N_21866,N_21372);
or U23273 (N_23273,N_20714,N_22443);
and U23274 (N_23274,N_21768,N_21848);
nor U23275 (N_23275,N_20380,N_20606);
or U23276 (N_23276,N_21044,N_22156);
or U23277 (N_23277,N_21220,N_21104);
nand U23278 (N_23278,N_20663,N_20087);
xnor U23279 (N_23279,N_20994,N_20465);
xor U23280 (N_23280,N_21779,N_21785);
nor U23281 (N_23281,N_21126,N_20228);
nor U23282 (N_23282,N_20523,N_20542);
nor U23283 (N_23283,N_21560,N_21297);
nand U23284 (N_23284,N_22074,N_21906);
or U23285 (N_23285,N_20453,N_21958);
nand U23286 (N_23286,N_20793,N_21096);
and U23287 (N_23287,N_20774,N_22128);
or U23288 (N_23288,N_21655,N_22309);
and U23289 (N_23289,N_21643,N_20594);
or U23290 (N_23290,N_21032,N_20983);
nor U23291 (N_23291,N_21891,N_20065);
or U23292 (N_23292,N_20862,N_20629);
and U23293 (N_23293,N_20761,N_22152);
xnor U23294 (N_23294,N_20293,N_20071);
nor U23295 (N_23295,N_21579,N_21725);
xnor U23296 (N_23296,N_21296,N_20988);
xnor U23297 (N_23297,N_21975,N_21718);
nor U23298 (N_23298,N_22267,N_22369);
xor U23299 (N_23299,N_21791,N_21100);
nand U23300 (N_23300,N_20530,N_22037);
or U23301 (N_23301,N_21099,N_20532);
nand U23302 (N_23302,N_21689,N_22151);
or U23303 (N_23303,N_20728,N_20132);
xnor U23304 (N_23304,N_20924,N_22391);
xor U23305 (N_23305,N_21847,N_22473);
nor U23306 (N_23306,N_21792,N_21155);
nand U23307 (N_23307,N_21533,N_20699);
nor U23308 (N_23308,N_21078,N_22491);
or U23309 (N_23309,N_21896,N_20655);
nor U23310 (N_23310,N_20360,N_21623);
xor U23311 (N_23311,N_21147,N_21014);
and U23312 (N_23312,N_21412,N_21251);
or U23313 (N_23313,N_22130,N_21558);
nor U23314 (N_23314,N_21648,N_21441);
or U23315 (N_23315,N_20790,N_21352);
nor U23316 (N_23316,N_20091,N_21357);
or U23317 (N_23317,N_22032,N_21049);
or U23318 (N_23318,N_20909,N_22439);
xnor U23319 (N_23319,N_22238,N_21424);
and U23320 (N_23320,N_20060,N_20543);
nand U23321 (N_23321,N_20587,N_21708);
nand U23322 (N_23322,N_22459,N_20581);
nor U23323 (N_23323,N_22325,N_20865);
or U23324 (N_23324,N_21802,N_20527);
and U23325 (N_23325,N_22171,N_20825);
xnor U23326 (N_23326,N_20242,N_20297);
and U23327 (N_23327,N_20951,N_20166);
nor U23328 (N_23328,N_21729,N_20194);
nor U23329 (N_23329,N_21315,N_21762);
nor U23330 (N_23330,N_21989,N_20213);
nor U23331 (N_23331,N_20261,N_20456);
nor U23332 (N_23332,N_21970,N_21374);
xor U23333 (N_23333,N_21241,N_20063);
xnor U23334 (N_23334,N_20771,N_20760);
or U23335 (N_23335,N_20649,N_20064);
nand U23336 (N_23336,N_20907,N_21629);
and U23337 (N_23337,N_20320,N_22230);
xnor U23338 (N_23338,N_20189,N_22246);
or U23339 (N_23339,N_22240,N_21151);
and U23340 (N_23340,N_20056,N_22225);
and U23341 (N_23341,N_20535,N_20499);
or U23342 (N_23342,N_22100,N_20101);
and U23343 (N_23343,N_20694,N_21602);
and U23344 (N_23344,N_21286,N_22495);
xnor U23345 (N_23345,N_21520,N_22167);
nand U23346 (N_23346,N_20232,N_20393);
nor U23347 (N_23347,N_20876,N_20838);
xor U23348 (N_23348,N_22274,N_20099);
nor U23349 (N_23349,N_22416,N_21247);
nor U23350 (N_23350,N_22265,N_22131);
nor U23351 (N_23351,N_22078,N_22488);
xnor U23352 (N_23352,N_21923,N_20937);
or U23353 (N_23353,N_21074,N_20082);
nor U23354 (N_23354,N_20451,N_20024);
xnor U23355 (N_23355,N_20304,N_21350);
and U23356 (N_23356,N_21351,N_20601);
xnor U23357 (N_23357,N_21822,N_21773);
nor U23358 (N_23358,N_22123,N_21757);
nor U23359 (N_23359,N_22496,N_20898);
nor U23360 (N_23360,N_21670,N_20159);
or U23361 (N_23361,N_21174,N_20186);
nor U23362 (N_23362,N_20054,N_22059);
or U23363 (N_23363,N_20953,N_22303);
nor U23364 (N_23364,N_22259,N_21728);
or U23365 (N_23365,N_21777,N_21730);
xnor U23366 (N_23366,N_20415,N_22299);
xnor U23367 (N_23367,N_22318,N_20872);
nor U23368 (N_23368,N_20381,N_21867);
and U23369 (N_23369,N_21188,N_20524);
nor U23370 (N_23370,N_21254,N_22204);
nand U23371 (N_23371,N_21404,N_22341);
nand U23372 (N_23372,N_20402,N_20787);
xor U23373 (N_23373,N_21808,N_21256);
or U23374 (N_23374,N_20902,N_22345);
xor U23375 (N_23375,N_20702,N_20201);
or U23376 (N_23376,N_21438,N_20808);
or U23377 (N_23377,N_20677,N_20658);
nor U23378 (N_23378,N_21047,N_21444);
xnor U23379 (N_23379,N_20960,N_21276);
xor U23380 (N_23380,N_20412,N_21510);
nor U23381 (N_23381,N_21830,N_20234);
nand U23382 (N_23382,N_20316,N_20384);
nand U23383 (N_23383,N_20337,N_20057);
or U23384 (N_23384,N_21751,N_20016);
and U23385 (N_23385,N_22018,N_20033);
nand U23386 (N_23386,N_22112,N_21169);
xor U23387 (N_23387,N_22146,N_21060);
or U23388 (N_23388,N_20180,N_20182);
xnor U23389 (N_23389,N_20726,N_21391);
xnor U23390 (N_23390,N_21605,N_22091);
xor U23391 (N_23391,N_21524,N_21339);
nor U23392 (N_23392,N_21111,N_21747);
or U23393 (N_23393,N_21386,N_21356);
and U23394 (N_23394,N_21615,N_22387);
and U23395 (N_23395,N_20370,N_20042);
xor U23396 (N_23396,N_22134,N_21526);
xnor U23397 (N_23397,N_20081,N_20420);
or U23398 (N_23398,N_21678,N_21153);
and U23399 (N_23399,N_22012,N_20716);
xor U23400 (N_23400,N_21570,N_21363);
and U23401 (N_23401,N_21641,N_22302);
nand U23402 (N_23402,N_21443,N_20053);
xor U23403 (N_23403,N_22456,N_22347);
nor U23404 (N_23404,N_21493,N_21299);
xor U23405 (N_23405,N_21659,N_20659);
and U23406 (N_23406,N_20211,N_20469);
nand U23407 (N_23407,N_21461,N_20519);
nand U23408 (N_23408,N_22367,N_20522);
nor U23409 (N_23409,N_20442,N_22483);
xnor U23410 (N_23410,N_21612,N_22486);
nor U23411 (N_23411,N_21815,N_20051);
or U23412 (N_23412,N_21771,N_20379);
xnor U23413 (N_23413,N_21257,N_20697);
nor U23414 (N_23414,N_21985,N_22009);
xor U23415 (N_23415,N_20651,N_22117);
nand U23416 (N_23416,N_22381,N_22338);
nor U23417 (N_23417,N_22315,N_20059);
xnor U23418 (N_23418,N_21059,N_21994);
and U23419 (N_23419,N_20991,N_21515);
nand U23420 (N_23420,N_21912,N_22159);
nand U23421 (N_23421,N_21917,N_20307);
and U23422 (N_23422,N_20489,N_21539);
or U23423 (N_23423,N_20809,N_22429);
or U23424 (N_23424,N_22441,N_22475);
nor U23425 (N_23425,N_20643,N_20449);
nand U23426 (N_23426,N_22196,N_20730);
nor U23427 (N_23427,N_22343,N_21393);
and U23428 (N_23428,N_20852,N_20357);
and U23429 (N_23429,N_22168,N_22455);
or U23430 (N_23430,N_21545,N_20124);
and U23431 (N_23431,N_21737,N_21246);
xor U23432 (N_23432,N_20358,N_22226);
nand U23433 (N_23433,N_20094,N_20684);
and U23434 (N_23434,N_20322,N_20563);
nand U23435 (N_23435,N_20255,N_20176);
nor U23436 (N_23436,N_21642,N_20259);
nand U23437 (N_23437,N_21478,N_20168);
xor U23438 (N_23438,N_20928,N_21323);
nand U23439 (N_23439,N_21694,N_22010);
or U23440 (N_23440,N_20916,N_22421);
or U23441 (N_23441,N_20207,N_21329);
xor U23442 (N_23442,N_22223,N_20552);
or U23443 (N_23443,N_20873,N_21159);
or U23444 (N_23444,N_21835,N_22036);
and U23445 (N_23445,N_21053,N_21496);
xnor U23446 (N_23446,N_20423,N_20382);
nand U23447 (N_23447,N_21285,N_22198);
or U23448 (N_23448,N_20152,N_22449);
nand U23449 (N_23449,N_21004,N_22040);
nand U23450 (N_23450,N_20365,N_21885);
xnor U23451 (N_23451,N_22042,N_20548);
nor U23452 (N_23452,N_22026,N_20274);
xor U23453 (N_23453,N_21684,N_20934);
nand U23454 (N_23454,N_20541,N_21132);
and U23455 (N_23455,N_22212,N_21261);
xor U23456 (N_23456,N_21224,N_22438);
or U23457 (N_23457,N_20149,N_20693);
nor U23458 (N_23458,N_21638,N_20511);
and U23459 (N_23459,N_20786,N_20328);
or U23460 (N_23460,N_21311,N_20795);
nand U23461 (N_23461,N_20231,N_21818);
and U23462 (N_23462,N_20546,N_21168);
or U23463 (N_23463,N_20561,N_21819);
nand U23464 (N_23464,N_21789,N_20778);
nand U23465 (N_23465,N_21221,N_20739);
nor U23466 (N_23466,N_20233,N_20299);
xor U23467 (N_23467,N_21903,N_20250);
nor U23468 (N_23468,N_22287,N_20564);
nor U23469 (N_23469,N_22013,N_21379);
xor U23470 (N_23470,N_22418,N_21557);
nand U23471 (N_23471,N_20323,N_20352);
nand U23472 (N_23472,N_21600,N_20408);
nand U23473 (N_23473,N_20540,N_22361);
xnor U23474 (N_23474,N_20947,N_20894);
nor U23475 (N_23475,N_21302,N_21317);
nand U23476 (N_23476,N_22297,N_20406);
or U23477 (N_23477,N_21875,N_21214);
or U23478 (N_23478,N_20477,N_22191);
nor U23479 (N_23479,N_22063,N_20895);
or U23480 (N_23480,N_20819,N_21187);
and U23481 (N_23481,N_20080,N_21152);
nor U23482 (N_23482,N_21204,N_22066);
or U23483 (N_23483,N_20706,N_22133);
or U23484 (N_23484,N_21928,N_21716);
nand U23485 (N_23485,N_20529,N_22065);
and U23486 (N_23486,N_22176,N_20173);
xor U23487 (N_23487,N_20797,N_20268);
nor U23488 (N_23488,N_22399,N_22275);
nand U23489 (N_23489,N_20302,N_21480);
or U23490 (N_23490,N_21569,N_20035);
and U23491 (N_23491,N_21938,N_20628);
nand U23492 (N_23492,N_20858,N_22121);
nor U23493 (N_23493,N_22210,N_20645);
nand U23494 (N_23494,N_21248,N_22336);
nand U23495 (N_23495,N_22050,N_21293);
xnor U23496 (N_23496,N_21333,N_21086);
nor U23497 (N_23497,N_21583,N_21348);
xnor U23498 (N_23498,N_21888,N_20416);
nand U23499 (N_23499,N_21303,N_20088);
or U23500 (N_23500,N_21192,N_20840);
nor U23501 (N_23501,N_20735,N_21305);
nor U23502 (N_23502,N_22243,N_20017);
nand U23503 (N_23503,N_22209,N_20290);
nand U23504 (N_23504,N_20590,N_22298);
xnor U23505 (N_23505,N_20230,N_21387);
nor U23506 (N_23506,N_20788,N_21990);
or U23507 (N_23507,N_21995,N_22319);
and U23508 (N_23508,N_22314,N_20470);
nor U23509 (N_23509,N_21692,N_20773);
or U23510 (N_23510,N_21021,N_22118);
or U23511 (N_23511,N_20715,N_20466);
xor U23512 (N_23512,N_21982,N_22366);
xnor U23513 (N_23513,N_20549,N_20848);
xor U23514 (N_23514,N_22257,N_20134);
nand U23515 (N_23515,N_20998,N_20903);
nor U23516 (N_23516,N_20330,N_21934);
and U23517 (N_23517,N_20742,N_22084);
or U23518 (N_23518,N_21375,N_21943);
or U23519 (N_23519,N_20505,N_22331);
xnor U23520 (N_23520,N_22020,N_21942);
nor U23521 (N_23521,N_20970,N_21259);
xnor U23522 (N_23522,N_21695,N_20896);
nand U23523 (N_23523,N_21601,N_22138);
xor U23524 (N_23524,N_20737,N_22222);
and U23525 (N_23525,N_22189,N_20718);
nor U23526 (N_23526,N_20508,N_21905);
nand U23527 (N_23527,N_20965,N_20745);
nand U23528 (N_23528,N_21490,N_20072);
nor U23529 (N_23529,N_20877,N_20098);
and U23530 (N_23530,N_21824,N_21763);
xor U23531 (N_23531,N_22170,N_20832);
nand U23532 (N_23532,N_21232,N_22142);
or U23533 (N_23533,N_21301,N_20435);
and U23534 (N_23534,N_21054,N_20429);
or U23535 (N_23535,N_21901,N_20222);
nor U23536 (N_23536,N_21036,N_20473);
or U23537 (N_23537,N_22086,N_20368);
nand U23538 (N_23538,N_20431,N_21205);
xnor U23539 (N_23539,N_20438,N_20084);
nand U23540 (N_23540,N_22285,N_20026);
and U23541 (N_23541,N_20095,N_20007);
or U23542 (N_23542,N_22426,N_20169);
and U23543 (N_23543,N_20270,N_21651);
or U23544 (N_23544,N_21034,N_20942);
nor U23545 (N_23545,N_22340,N_20245);
or U23546 (N_23546,N_21976,N_20481);
or U23547 (N_23547,N_20662,N_21544);
and U23548 (N_23548,N_20193,N_21512);
nor U23549 (N_23549,N_21290,N_22277);
nand U23550 (N_23550,N_20611,N_20636);
or U23551 (N_23551,N_21400,N_21033);
and U23552 (N_23552,N_21178,N_22027);
nor U23553 (N_23553,N_22011,N_22192);
nor U23554 (N_23554,N_20682,N_20263);
or U23555 (N_23555,N_21472,N_21930);
and U23556 (N_23556,N_20164,N_21590);
and U23557 (N_23557,N_20006,N_20418);
and U23558 (N_23558,N_22214,N_21177);
nor U23559 (N_23559,N_20317,N_20100);
and U23560 (N_23560,N_21341,N_22110);
nand U23561 (N_23561,N_21549,N_21328);
xor U23562 (N_23562,N_20083,N_21101);
nor U23563 (N_23563,N_21229,N_22082);
or U23564 (N_23564,N_20468,N_22279);
and U23565 (N_23565,N_20630,N_21061);
and U23566 (N_23566,N_22157,N_21154);
xnor U23567 (N_23567,N_20411,N_20215);
xor U23568 (N_23568,N_22247,N_20789);
nand U23569 (N_23569,N_20311,N_20217);
or U23570 (N_23570,N_21140,N_22116);
nor U23571 (N_23571,N_20424,N_21795);
or U23572 (N_23572,N_21012,N_20855);
and U23573 (N_23573,N_22301,N_21662);
or U23574 (N_23574,N_21253,N_20792);
xnor U23575 (N_23575,N_21784,N_21000);
and U23576 (N_23576,N_20557,N_20444);
and U23577 (N_23577,N_21436,N_21408);
xnor U23578 (N_23578,N_22365,N_21208);
nand U23579 (N_23579,N_22397,N_21122);
nand U23580 (N_23580,N_22378,N_20276);
or U23581 (N_23581,N_20989,N_21527);
nor U23582 (N_23582,N_21620,N_22053);
and U23583 (N_23583,N_22289,N_20398);
and U23584 (N_23584,N_20598,N_20219);
nand U23585 (N_23585,N_20618,N_20943);
or U23586 (N_23586,N_20944,N_20687);
or U23587 (N_23587,N_21556,N_20823);
or U23588 (N_23588,N_21932,N_20027);
nand U23589 (N_23589,N_20243,N_20856);
nand U23590 (N_23590,N_22464,N_21394);
nand U23591 (N_23591,N_22172,N_20565);
nand U23592 (N_23592,N_20378,N_20631);
nor U23593 (N_23593,N_20480,N_20309);
xnor U23594 (N_23594,N_20458,N_21576);
xnor U23595 (N_23595,N_20077,N_20668);
nor U23596 (N_23596,N_21268,N_21231);
xor U23597 (N_23597,N_21758,N_20055);
and U23598 (N_23598,N_20691,N_20861);
nor U23599 (N_23599,N_21452,N_21929);
nand U23600 (N_23600,N_22431,N_20361);
nor U23601 (N_23601,N_20260,N_22412);
nand U23602 (N_23602,N_22327,N_21850);
or U23603 (N_23603,N_20930,N_20780);
nand U23604 (N_23604,N_22239,N_20914);
and U23605 (N_23605,N_20811,N_22181);
nor U23606 (N_23606,N_21250,N_21663);
xor U23607 (N_23607,N_20946,N_20474);
and U23608 (N_23608,N_22290,N_20880);
or U23609 (N_23609,N_20968,N_21827);
nand U23610 (N_23610,N_21226,N_21172);
and U23611 (N_23611,N_21532,N_20153);
or U23612 (N_23612,N_21700,N_20842);
xor U23613 (N_23613,N_20799,N_21486);
nor U23614 (N_23614,N_21582,N_20997);
nand U23615 (N_23615,N_20172,N_20325);
or U23616 (N_23616,N_21727,N_22472);
and U23617 (N_23617,N_21368,N_20195);
or U23618 (N_23618,N_22471,N_20833);
nand U23619 (N_23619,N_20109,N_20956);
nand U23620 (N_23620,N_21797,N_22480);
nand U23621 (N_23621,N_21733,N_20394);
or U23622 (N_23622,N_21264,N_22221);
nor U23623 (N_23623,N_21846,N_22030);
nor U23624 (N_23624,N_20391,N_21125);
xor U23625 (N_23625,N_22046,N_21383);
nor U23626 (N_23626,N_20102,N_22047);
nor U23627 (N_23627,N_21927,N_20421);
and U23628 (N_23628,N_22423,N_22281);
and U23629 (N_23629,N_20075,N_21189);
nor U23630 (N_23630,N_21218,N_20045);
xnor U23631 (N_23631,N_20125,N_21319);
and U23632 (N_23632,N_21978,N_21649);
and U23633 (N_23633,N_21492,N_21821);
and U23634 (N_23634,N_22051,N_22224);
xor U23635 (N_23635,N_21336,N_21585);
or U23636 (N_23636,N_20555,N_22135);
or U23637 (N_23637,N_20482,N_21607);
nor U23638 (N_23638,N_22468,N_20278);
nor U23639 (N_23639,N_20351,N_20889);
or U23640 (N_23640,N_21433,N_21471);
xor U23641 (N_23641,N_21094,N_21421);
and U23642 (N_23642,N_20567,N_22044);
nor U23643 (N_23643,N_21956,N_20061);
xnor U23644 (N_23644,N_21454,N_21974);
or U23645 (N_23645,N_21868,N_20935);
or U23646 (N_23646,N_21542,N_21252);
or U23647 (N_23647,N_22453,N_20831);
and U23648 (N_23648,N_20860,N_20804);
or U23649 (N_23649,N_20400,N_21173);
nor U23650 (N_23650,N_22101,N_21055);
xnor U23651 (N_23651,N_20269,N_20181);
and U23652 (N_23652,N_20882,N_22174);
xor U23653 (N_23653,N_20950,N_21347);
xor U23654 (N_23654,N_21119,N_20392);
nor U23655 (N_23655,N_21015,N_20712);
and U23656 (N_23656,N_20901,N_20931);
nor U23657 (N_23657,N_21415,N_22442);
and U23658 (N_23658,N_22155,N_22215);
and U23659 (N_23659,N_22355,N_21138);
nand U23660 (N_23660,N_22266,N_20036);
and U23661 (N_23661,N_20846,N_21127);
xnor U23662 (N_23662,N_20772,N_22028);
and U23663 (N_23663,N_20813,N_20884);
or U23664 (N_23664,N_20298,N_21619);
or U23665 (N_23665,N_21541,N_20932);
and U23666 (N_23666,N_20374,N_21595);
and U23667 (N_23667,N_20607,N_22380);
xor U23668 (N_23668,N_22354,N_21203);
nand U23669 (N_23669,N_21955,N_20503);
nand U23670 (N_23670,N_21953,N_22450);
nand U23671 (N_23671,N_20992,N_20892);
and U23672 (N_23672,N_20009,N_20040);
and U23673 (N_23673,N_20498,N_22466);
nor U23674 (N_23674,N_20701,N_21008);
nor U23675 (N_23675,N_20753,N_20126);
and U23676 (N_23676,N_22346,N_20433);
or U23677 (N_23677,N_22470,N_21553);
nor U23678 (N_23678,N_21561,N_20720);
xnor U23679 (N_23679,N_20545,N_20904);
and U23680 (N_23680,N_20144,N_20210);
or U23681 (N_23681,N_21396,N_20462);
xnor U23682 (N_23682,N_21860,N_20653);
and U23683 (N_23683,N_22175,N_21277);
nand U23684 (N_23684,N_21289,N_20757);
or U23685 (N_23685,N_21852,N_20258);
nand U23686 (N_23686,N_21650,N_21500);
nor U23687 (N_23687,N_20069,N_20961);
or U23688 (N_23688,N_21407,N_22185);
and U23689 (N_23689,N_21359,N_22420);
nor U23690 (N_23690,N_21872,N_20515);
xnor U23691 (N_23691,N_20537,N_22451);
or U23692 (N_23692,N_20974,N_20836);
and U23693 (N_23693,N_21856,N_21826);
nand U23694 (N_23694,N_20155,N_21087);
nor U23695 (N_23695,N_21799,N_22432);
nor U23696 (N_23696,N_20743,N_20980);
nor U23697 (N_23697,N_21149,N_21834);
and U23698 (N_23698,N_22164,N_20119);
nand U23699 (N_23699,N_21123,N_21535);
xnor U23700 (N_23700,N_21381,N_21064);
or U23701 (N_23701,N_20723,N_22190);
or U23702 (N_23702,N_20364,N_20277);
nor U23703 (N_23703,N_21501,N_20656);
xnor U23704 (N_23704,N_20397,N_20926);
or U23705 (N_23705,N_20830,N_21035);
or U23706 (N_23706,N_20517,N_20727);
and U23707 (N_23707,N_22493,N_20767);
and U23708 (N_23708,N_20768,N_21809);
and U23709 (N_23709,N_20202,N_20171);
or U23710 (N_23710,N_21744,N_22015);
nand U23711 (N_23711,N_21397,N_21754);
nand U23712 (N_23712,N_21378,N_21710);
nand U23713 (N_23713,N_21793,N_20729);
nor U23714 (N_23714,N_20794,N_21554);
nand U23715 (N_23715,N_20562,N_20744);
nand U23716 (N_23716,N_21211,N_21067);
nor U23717 (N_23717,N_21124,N_21759);
nand U23718 (N_23718,N_21469,N_22124);
nand U23719 (N_23719,N_20908,N_21165);
or U23720 (N_23720,N_20160,N_20010);
nor U23721 (N_23721,N_20058,N_22357);
nor U23722 (N_23722,N_20985,N_21706);
nand U23723 (N_23723,N_22389,N_22440);
or U23724 (N_23724,N_21886,N_20888);
xnor U23725 (N_23725,N_20156,N_21090);
nand U23726 (N_23726,N_22183,N_20117);
or U23727 (N_23727,N_20136,N_20163);
xnor U23728 (N_23728,N_20614,N_20766);
and U23729 (N_23729,N_21282,N_20674);
nor U23730 (N_23730,N_20782,N_21065);
and U23731 (N_23731,N_22251,N_22402);
nand U23732 (N_23732,N_22187,N_22424);
nand U23733 (N_23733,N_20285,N_20949);
or U23734 (N_23734,N_21673,N_21392);
xnor U23735 (N_23735,N_20597,N_20353);
nor U23736 (N_23736,N_20165,N_21088);
or U23737 (N_23737,N_21006,N_21118);
xor U23738 (N_23738,N_22098,N_20001);
or U23739 (N_23739,N_20820,N_21405);
and U23740 (N_23740,N_20096,N_22388);
nor U23741 (N_23741,N_21933,N_20267);
nand U23742 (N_23742,N_20734,N_21630);
and U23743 (N_23743,N_21844,N_21129);
or U23744 (N_23744,N_21423,N_21401);
xor U23745 (N_23745,N_21288,N_21115);
xnor U23746 (N_23746,N_20348,N_20229);
and U23747 (N_23747,N_21957,N_21019);
or U23748 (N_23748,N_20765,N_21007);
nor U23749 (N_23749,N_22132,N_20783);
and U23750 (N_23750,N_21280,N_21592);
nand U23751 (N_23751,N_22201,N_22131);
nand U23752 (N_23752,N_20659,N_20573);
nand U23753 (N_23753,N_20248,N_20325);
and U23754 (N_23754,N_20366,N_20497);
xor U23755 (N_23755,N_20480,N_20512);
nand U23756 (N_23756,N_20180,N_22075);
nor U23757 (N_23757,N_21102,N_20908);
nand U23758 (N_23758,N_21555,N_20406);
nand U23759 (N_23759,N_20404,N_21881);
nor U23760 (N_23760,N_20531,N_20514);
xor U23761 (N_23761,N_21533,N_20927);
nor U23762 (N_23762,N_21566,N_22474);
and U23763 (N_23763,N_21753,N_22305);
xor U23764 (N_23764,N_21898,N_21254);
nand U23765 (N_23765,N_21676,N_20845);
and U23766 (N_23766,N_21347,N_22344);
or U23767 (N_23767,N_20905,N_21216);
or U23768 (N_23768,N_21262,N_20102);
nor U23769 (N_23769,N_21700,N_22212);
or U23770 (N_23770,N_20153,N_22259);
nor U23771 (N_23771,N_20104,N_21689);
nand U23772 (N_23772,N_21835,N_21498);
or U23773 (N_23773,N_21865,N_21396);
nor U23774 (N_23774,N_20399,N_21057);
and U23775 (N_23775,N_21196,N_22363);
xor U23776 (N_23776,N_22126,N_20620);
or U23777 (N_23777,N_20669,N_20352);
or U23778 (N_23778,N_20973,N_21329);
nand U23779 (N_23779,N_20982,N_20940);
nand U23780 (N_23780,N_21308,N_21631);
nand U23781 (N_23781,N_20175,N_20252);
and U23782 (N_23782,N_21305,N_21907);
or U23783 (N_23783,N_21922,N_21958);
xor U23784 (N_23784,N_22222,N_21952);
nor U23785 (N_23785,N_22335,N_20534);
xor U23786 (N_23786,N_21116,N_22091);
nor U23787 (N_23787,N_20163,N_20409);
and U23788 (N_23788,N_22233,N_21792);
or U23789 (N_23789,N_20702,N_21529);
nor U23790 (N_23790,N_20293,N_22483);
nand U23791 (N_23791,N_20510,N_21867);
xnor U23792 (N_23792,N_21262,N_20884);
nor U23793 (N_23793,N_20268,N_21815);
or U23794 (N_23794,N_21036,N_21430);
or U23795 (N_23795,N_20074,N_21577);
xnor U23796 (N_23796,N_22008,N_21319);
nor U23797 (N_23797,N_20010,N_22377);
and U23798 (N_23798,N_21310,N_20295);
and U23799 (N_23799,N_22013,N_20953);
and U23800 (N_23800,N_21114,N_20452);
and U23801 (N_23801,N_22287,N_20544);
and U23802 (N_23802,N_20881,N_21977);
nor U23803 (N_23803,N_20798,N_20394);
or U23804 (N_23804,N_20981,N_22065);
and U23805 (N_23805,N_21201,N_20182);
xor U23806 (N_23806,N_21677,N_20682);
and U23807 (N_23807,N_21006,N_22366);
nor U23808 (N_23808,N_22122,N_20555);
nor U23809 (N_23809,N_20670,N_20594);
nor U23810 (N_23810,N_21918,N_21986);
nor U23811 (N_23811,N_22382,N_22185);
nor U23812 (N_23812,N_20165,N_21904);
or U23813 (N_23813,N_22144,N_20813);
and U23814 (N_23814,N_21133,N_21164);
and U23815 (N_23815,N_20550,N_21536);
xnor U23816 (N_23816,N_21616,N_21444);
and U23817 (N_23817,N_21121,N_22209);
or U23818 (N_23818,N_20096,N_21589);
nor U23819 (N_23819,N_20596,N_21009);
and U23820 (N_23820,N_21886,N_21367);
nand U23821 (N_23821,N_20690,N_20938);
and U23822 (N_23822,N_20738,N_22000);
or U23823 (N_23823,N_21220,N_21900);
and U23824 (N_23824,N_20938,N_20183);
nand U23825 (N_23825,N_20529,N_20792);
xor U23826 (N_23826,N_21753,N_22047);
and U23827 (N_23827,N_21257,N_20124);
nand U23828 (N_23828,N_20688,N_21041);
nand U23829 (N_23829,N_22127,N_20273);
or U23830 (N_23830,N_20397,N_20619);
or U23831 (N_23831,N_20690,N_21902);
xnor U23832 (N_23832,N_21148,N_21436);
or U23833 (N_23833,N_20065,N_21154);
xor U23834 (N_23834,N_21766,N_20315);
or U23835 (N_23835,N_22236,N_20398);
or U23836 (N_23836,N_21467,N_20201);
or U23837 (N_23837,N_21091,N_20361);
or U23838 (N_23838,N_22438,N_20494);
nand U23839 (N_23839,N_20444,N_20946);
or U23840 (N_23840,N_21427,N_22135);
xnor U23841 (N_23841,N_21715,N_20296);
or U23842 (N_23842,N_21652,N_20331);
nand U23843 (N_23843,N_20107,N_20018);
nand U23844 (N_23844,N_21947,N_20265);
and U23845 (N_23845,N_20732,N_20205);
xor U23846 (N_23846,N_22372,N_21001);
xnor U23847 (N_23847,N_20613,N_21085);
nor U23848 (N_23848,N_21847,N_21549);
and U23849 (N_23849,N_22167,N_20524);
and U23850 (N_23850,N_22127,N_21376);
nand U23851 (N_23851,N_22399,N_21748);
nor U23852 (N_23852,N_20704,N_22417);
or U23853 (N_23853,N_20553,N_20830);
and U23854 (N_23854,N_21216,N_20363);
nand U23855 (N_23855,N_21301,N_21060);
xnor U23856 (N_23856,N_21411,N_20753);
or U23857 (N_23857,N_21610,N_21802);
nand U23858 (N_23858,N_22129,N_21250);
xor U23859 (N_23859,N_21970,N_21050);
nor U23860 (N_23860,N_20275,N_22433);
and U23861 (N_23861,N_21303,N_20147);
nor U23862 (N_23862,N_20284,N_21315);
or U23863 (N_23863,N_20577,N_21006);
nor U23864 (N_23864,N_21305,N_20302);
nor U23865 (N_23865,N_20221,N_20269);
and U23866 (N_23866,N_22202,N_22252);
nand U23867 (N_23867,N_21936,N_20198);
nor U23868 (N_23868,N_20179,N_22457);
and U23869 (N_23869,N_20582,N_21925);
xnor U23870 (N_23870,N_21288,N_22015);
nor U23871 (N_23871,N_21878,N_20803);
or U23872 (N_23872,N_20806,N_20549);
nor U23873 (N_23873,N_20045,N_21113);
xnor U23874 (N_23874,N_20056,N_20306);
and U23875 (N_23875,N_20142,N_22472);
or U23876 (N_23876,N_22342,N_20715);
nor U23877 (N_23877,N_20533,N_20921);
nand U23878 (N_23878,N_21496,N_20621);
nand U23879 (N_23879,N_21683,N_22259);
and U23880 (N_23880,N_20181,N_21309);
or U23881 (N_23881,N_21987,N_22177);
and U23882 (N_23882,N_20176,N_22045);
and U23883 (N_23883,N_21434,N_21604);
and U23884 (N_23884,N_21566,N_22343);
nand U23885 (N_23885,N_21138,N_21587);
or U23886 (N_23886,N_20417,N_20477);
nand U23887 (N_23887,N_20483,N_22402);
nor U23888 (N_23888,N_21624,N_21353);
xnor U23889 (N_23889,N_20533,N_21137);
xor U23890 (N_23890,N_20328,N_20576);
and U23891 (N_23891,N_20293,N_21058);
nor U23892 (N_23892,N_22323,N_21583);
nor U23893 (N_23893,N_20712,N_22297);
nor U23894 (N_23894,N_20111,N_21603);
xor U23895 (N_23895,N_20676,N_20640);
or U23896 (N_23896,N_20324,N_21817);
nand U23897 (N_23897,N_21450,N_20422);
or U23898 (N_23898,N_21550,N_21946);
xor U23899 (N_23899,N_22107,N_22280);
xor U23900 (N_23900,N_22419,N_20909);
or U23901 (N_23901,N_20129,N_22227);
xnor U23902 (N_23902,N_20234,N_22358);
or U23903 (N_23903,N_20675,N_21030);
or U23904 (N_23904,N_21541,N_21692);
and U23905 (N_23905,N_21750,N_21226);
or U23906 (N_23906,N_21985,N_20171);
nand U23907 (N_23907,N_20954,N_21624);
or U23908 (N_23908,N_20689,N_20893);
and U23909 (N_23909,N_21307,N_22225);
and U23910 (N_23910,N_20750,N_21187);
and U23911 (N_23911,N_21742,N_21575);
nor U23912 (N_23912,N_20685,N_20034);
xnor U23913 (N_23913,N_21578,N_20076);
or U23914 (N_23914,N_20702,N_20697);
or U23915 (N_23915,N_20427,N_21801);
or U23916 (N_23916,N_21682,N_20199);
nand U23917 (N_23917,N_22441,N_20282);
and U23918 (N_23918,N_21224,N_20516);
nor U23919 (N_23919,N_21336,N_21616);
nand U23920 (N_23920,N_21640,N_21596);
xor U23921 (N_23921,N_20515,N_20826);
or U23922 (N_23922,N_20182,N_21052);
nand U23923 (N_23923,N_20221,N_22490);
nand U23924 (N_23924,N_21920,N_20916);
nand U23925 (N_23925,N_21455,N_22094);
and U23926 (N_23926,N_21739,N_21423);
or U23927 (N_23927,N_20602,N_21302);
or U23928 (N_23928,N_20188,N_20557);
or U23929 (N_23929,N_20151,N_20646);
xnor U23930 (N_23930,N_20895,N_22358);
xor U23931 (N_23931,N_22149,N_20167);
nand U23932 (N_23932,N_21105,N_21533);
nand U23933 (N_23933,N_21092,N_22277);
xor U23934 (N_23934,N_22411,N_20611);
xnor U23935 (N_23935,N_21183,N_22053);
and U23936 (N_23936,N_20155,N_20701);
nor U23937 (N_23937,N_22286,N_20502);
nor U23938 (N_23938,N_20800,N_22093);
or U23939 (N_23939,N_21587,N_21519);
xor U23940 (N_23940,N_20531,N_20994);
nor U23941 (N_23941,N_21083,N_20016);
or U23942 (N_23942,N_22356,N_20113);
nand U23943 (N_23943,N_21866,N_21757);
nand U23944 (N_23944,N_20847,N_20295);
nor U23945 (N_23945,N_20587,N_22482);
and U23946 (N_23946,N_20799,N_21361);
nand U23947 (N_23947,N_22135,N_21648);
nand U23948 (N_23948,N_21493,N_20621);
or U23949 (N_23949,N_21784,N_20114);
xnor U23950 (N_23950,N_21742,N_21484);
and U23951 (N_23951,N_22054,N_21613);
and U23952 (N_23952,N_20342,N_22089);
or U23953 (N_23953,N_20535,N_20486);
nor U23954 (N_23954,N_21134,N_20716);
xnor U23955 (N_23955,N_21025,N_21153);
nand U23956 (N_23956,N_21178,N_21124);
or U23957 (N_23957,N_21811,N_21892);
xor U23958 (N_23958,N_20247,N_20526);
xnor U23959 (N_23959,N_21236,N_20628);
or U23960 (N_23960,N_21763,N_22256);
nor U23961 (N_23961,N_21961,N_22011);
xor U23962 (N_23962,N_21374,N_22436);
or U23963 (N_23963,N_22433,N_20239);
and U23964 (N_23964,N_21765,N_21795);
and U23965 (N_23965,N_21451,N_22454);
and U23966 (N_23966,N_21574,N_20657);
and U23967 (N_23967,N_22192,N_21116);
xor U23968 (N_23968,N_21514,N_20787);
or U23969 (N_23969,N_22445,N_22036);
nor U23970 (N_23970,N_21707,N_22040);
or U23971 (N_23971,N_20402,N_22098);
or U23972 (N_23972,N_20220,N_20190);
and U23973 (N_23973,N_22037,N_21443);
xnor U23974 (N_23974,N_20685,N_21938);
nor U23975 (N_23975,N_20529,N_21126);
and U23976 (N_23976,N_21408,N_20391);
nand U23977 (N_23977,N_22197,N_21891);
or U23978 (N_23978,N_21856,N_20304);
or U23979 (N_23979,N_22025,N_21897);
or U23980 (N_23980,N_20064,N_20510);
and U23981 (N_23981,N_21792,N_21104);
xnor U23982 (N_23982,N_20191,N_20290);
or U23983 (N_23983,N_20656,N_20591);
nor U23984 (N_23984,N_22447,N_22024);
and U23985 (N_23985,N_20961,N_22379);
xor U23986 (N_23986,N_20662,N_20512);
and U23987 (N_23987,N_21775,N_21805);
nor U23988 (N_23988,N_21090,N_21250);
xor U23989 (N_23989,N_22043,N_20946);
or U23990 (N_23990,N_22371,N_22246);
nor U23991 (N_23991,N_20844,N_20986);
or U23992 (N_23992,N_20183,N_21452);
or U23993 (N_23993,N_20344,N_20683);
xor U23994 (N_23994,N_20389,N_20949);
nor U23995 (N_23995,N_22364,N_20740);
nand U23996 (N_23996,N_22333,N_21862);
nand U23997 (N_23997,N_20006,N_22287);
and U23998 (N_23998,N_20645,N_20649);
nor U23999 (N_23999,N_21283,N_21758);
or U24000 (N_24000,N_20364,N_21939);
or U24001 (N_24001,N_21748,N_22366);
nor U24002 (N_24002,N_20376,N_20005);
and U24003 (N_24003,N_20347,N_22274);
nand U24004 (N_24004,N_20272,N_21122);
or U24005 (N_24005,N_22184,N_20182);
xnor U24006 (N_24006,N_21216,N_21036);
or U24007 (N_24007,N_22003,N_20070);
and U24008 (N_24008,N_20964,N_21891);
nand U24009 (N_24009,N_21014,N_20949);
and U24010 (N_24010,N_21854,N_20548);
or U24011 (N_24011,N_20953,N_20902);
or U24012 (N_24012,N_20760,N_22411);
nor U24013 (N_24013,N_22397,N_21982);
nand U24014 (N_24014,N_20518,N_21812);
nor U24015 (N_24015,N_21968,N_21288);
or U24016 (N_24016,N_20866,N_20170);
xor U24017 (N_24017,N_21652,N_20752);
xnor U24018 (N_24018,N_20760,N_21166);
xnor U24019 (N_24019,N_21151,N_22297);
nor U24020 (N_24020,N_20276,N_20556);
or U24021 (N_24021,N_20195,N_21791);
or U24022 (N_24022,N_21996,N_22032);
xnor U24023 (N_24023,N_21338,N_22060);
xor U24024 (N_24024,N_20237,N_22228);
nor U24025 (N_24025,N_20510,N_20992);
xnor U24026 (N_24026,N_20601,N_21973);
nand U24027 (N_24027,N_21294,N_22495);
nor U24028 (N_24028,N_20929,N_21345);
nand U24029 (N_24029,N_22475,N_22376);
nand U24030 (N_24030,N_22118,N_21290);
nor U24031 (N_24031,N_22435,N_21822);
nand U24032 (N_24032,N_22259,N_20835);
nor U24033 (N_24033,N_20064,N_20916);
or U24034 (N_24034,N_20516,N_22400);
or U24035 (N_24035,N_22250,N_21253);
xnor U24036 (N_24036,N_20221,N_20538);
xnor U24037 (N_24037,N_22150,N_20958);
nand U24038 (N_24038,N_21608,N_20979);
or U24039 (N_24039,N_22185,N_21839);
nand U24040 (N_24040,N_20160,N_22494);
nor U24041 (N_24041,N_20870,N_20992);
or U24042 (N_24042,N_20614,N_20521);
or U24043 (N_24043,N_21531,N_20086);
nor U24044 (N_24044,N_21558,N_20338);
or U24045 (N_24045,N_20138,N_21366);
nand U24046 (N_24046,N_21849,N_21369);
nor U24047 (N_24047,N_20821,N_22458);
xnor U24048 (N_24048,N_20106,N_21108);
nand U24049 (N_24049,N_21680,N_20964);
nor U24050 (N_24050,N_21430,N_21368);
nor U24051 (N_24051,N_21190,N_21844);
nand U24052 (N_24052,N_21957,N_20009);
and U24053 (N_24053,N_21184,N_21696);
or U24054 (N_24054,N_22465,N_21409);
nor U24055 (N_24055,N_20129,N_20794);
and U24056 (N_24056,N_21361,N_20915);
and U24057 (N_24057,N_22408,N_21600);
nor U24058 (N_24058,N_20304,N_22173);
nand U24059 (N_24059,N_21160,N_21000);
xor U24060 (N_24060,N_21385,N_21300);
xnor U24061 (N_24061,N_21469,N_20676);
or U24062 (N_24062,N_20930,N_21847);
and U24063 (N_24063,N_21658,N_20531);
nor U24064 (N_24064,N_21797,N_20981);
nand U24065 (N_24065,N_22487,N_20001);
and U24066 (N_24066,N_21799,N_21462);
nand U24067 (N_24067,N_21067,N_21235);
nand U24068 (N_24068,N_20310,N_21119);
nand U24069 (N_24069,N_20081,N_20123);
xnor U24070 (N_24070,N_21497,N_20236);
nand U24071 (N_24071,N_21273,N_21470);
xnor U24072 (N_24072,N_20979,N_20721);
nor U24073 (N_24073,N_21348,N_20219);
and U24074 (N_24074,N_21365,N_22203);
xor U24075 (N_24075,N_21144,N_21460);
nand U24076 (N_24076,N_21309,N_22198);
and U24077 (N_24077,N_20451,N_22140);
or U24078 (N_24078,N_20906,N_21993);
nand U24079 (N_24079,N_22052,N_21523);
nor U24080 (N_24080,N_20522,N_21076);
and U24081 (N_24081,N_20081,N_22159);
nor U24082 (N_24082,N_22052,N_22146);
xnor U24083 (N_24083,N_21500,N_20323);
xnor U24084 (N_24084,N_20523,N_20098);
xnor U24085 (N_24085,N_20775,N_21969);
xnor U24086 (N_24086,N_21832,N_20832);
or U24087 (N_24087,N_22337,N_21542);
nand U24088 (N_24088,N_21196,N_21441);
nand U24089 (N_24089,N_21263,N_20771);
xor U24090 (N_24090,N_21699,N_21354);
or U24091 (N_24091,N_22400,N_22466);
nor U24092 (N_24092,N_21989,N_21067);
nor U24093 (N_24093,N_21641,N_21755);
nor U24094 (N_24094,N_21038,N_20416);
nand U24095 (N_24095,N_20902,N_22280);
nand U24096 (N_24096,N_22312,N_21514);
nor U24097 (N_24097,N_22145,N_21107);
nor U24098 (N_24098,N_20046,N_22102);
and U24099 (N_24099,N_20093,N_20255);
and U24100 (N_24100,N_20449,N_21833);
nand U24101 (N_24101,N_20693,N_22235);
or U24102 (N_24102,N_20812,N_20236);
xnor U24103 (N_24103,N_20987,N_20914);
and U24104 (N_24104,N_20005,N_21583);
nand U24105 (N_24105,N_21365,N_21445);
xor U24106 (N_24106,N_20465,N_22432);
nor U24107 (N_24107,N_21706,N_22241);
xor U24108 (N_24108,N_22201,N_22121);
nand U24109 (N_24109,N_20216,N_20795);
and U24110 (N_24110,N_21781,N_22378);
or U24111 (N_24111,N_21983,N_20414);
and U24112 (N_24112,N_21862,N_22263);
xor U24113 (N_24113,N_20305,N_20484);
nand U24114 (N_24114,N_22186,N_22299);
and U24115 (N_24115,N_21052,N_21336);
xnor U24116 (N_24116,N_20313,N_20006);
or U24117 (N_24117,N_22277,N_20520);
nor U24118 (N_24118,N_20165,N_20115);
or U24119 (N_24119,N_21958,N_22351);
nor U24120 (N_24120,N_20847,N_21070);
nor U24121 (N_24121,N_20652,N_20202);
nand U24122 (N_24122,N_20933,N_20166);
nor U24123 (N_24123,N_20176,N_20382);
nor U24124 (N_24124,N_20356,N_20202);
or U24125 (N_24125,N_22146,N_21550);
nor U24126 (N_24126,N_21999,N_20227);
nor U24127 (N_24127,N_20271,N_21608);
and U24128 (N_24128,N_22255,N_20068);
nor U24129 (N_24129,N_20165,N_20229);
nor U24130 (N_24130,N_21714,N_20292);
and U24131 (N_24131,N_21024,N_20837);
and U24132 (N_24132,N_22006,N_20874);
nor U24133 (N_24133,N_20297,N_21524);
nand U24134 (N_24134,N_20089,N_22233);
xnor U24135 (N_24135,N_21618,N_20664);
xor U24136 (N_24136,N_20131,N_21249);
or U24137 (N_24137,N_20351,N_21967);
or U24138 (N_24138,N_20501,N_20110);
nor U24139 (N_24139,N_21361,N_21837);
nand U24140 (N_24140,N_21674,N_22070);
xnor U24141 (N_24141,N_21177,N_20339);
nor U24142 (N_24142,N_21064,N_21013);
and U24143 (N_24143,N_21095,N_22144);
xor U24144 (N_24144,N_22239,N_20303);
xnor U24145 (N_24145,N_22121,N_22027);
nand U24146 (N_24146,N_21400,N_20562);
nand U24147 (N_24147,N_20973,N_20655);
nand U24148 (N_24148,N_21477,N_21476);
or U24149 (N_24149,N_20406,N_21014);
nand U24150 (N_24150,N_20689,N_21594);
and U24151 (N_24151,N_21975,N_21439);
and U24152 (N_24152,N_21298,N_20427);
nand U24153 (N_24153,N_21065,N_20518);
and U24154 (N_24154,N_22144,N_22114);
or U24155 (N_24155,N_21367,N_21752);
and U24156 (N_24156,N_20737,N_21965);
and U24157 (N_24157,N_20123,N_22159);
nand U24158 (N_24158,N_21283,N_20075);
and U24159 (N_24159,N_21464,N_22113);
or U24160 (N_24160,N_21518,N_20654);
and U24161 (N_24161,N_21163,N_21623);
nand U24162 (N_24162,N_21365,N_20323);
or U24163 (N_24163,N_20228,N_21776);
xor U24164 (N_24164,N_21902,N_20023);
xnor U24165 (N_24165,N_20584,N_21026);
nor U24166 (N_24166,N_20545,N_20255);
or U24167 (N_24167,N_20408,N_21591);
nand U24168 (N_24168,N_21717,N_21707);
nor U24169 (N_24169,N_21349,N_21606);
nand U24170 (N_24170,N_21378,N_21365);
or U24171 (N_24171,N_22271,N_22435);
xnor U24172 (N_24172,N_21762,N_21035);
nand U24173 (N_24173,N_21412,N_20962);
nand U24174 (N_24174,N_21626,N_20558);
xnor U24175 (N_24175,N_21586,N_20073);
and U24176 (N_24176,N_22387,N_20318);
and U24177 (N_24177,N_20377,N_20432);
nor U24178 (N_24178,N_20946,N_21782);
or U24179 (N_24179,N_20346,N_20509);
xnor U24180 (N_24180,N_21734,N_21677);
and U24181 (N_24181,N_20448,N_21638);
or U24182 (N_24182,N_22041,N_20409);
nand U24183 (N_24183,N_22092,N_21609);
xor U24184 (N_24184,N_22088,N_20090);
and U24185 (N_24185,N_20531,N_20799);
or U24186 (N_24186,N_21650,N_21546);
nand U24187 (N_24187,N_21118,N_20434);
nand U24188 (N_24188,N_22251,N_21026);
and U24189 (N_24189,N_21236,N_22270);
or U24190 (N_24190,N_20494,N_22003);
nand U24191 (N_24191,N_21200,N_21699);
xor U24192 (N_24192,N_20984,N_20212);
nor U24193 (N_24193,N_20154,N_20524);
xor U24194 (N_24194,N_21843,N_20359);
xnor U24195 (N_24195,N_20705,N_20493);
or U24196 (N_24196,N_21056,N_20896);
and U24197 (N_24197,N_22169,N_20779);
nor U24198 (N_24198,N_21199,N_20203);
xnor U24199 (N_24199,N_21215,N_20827);
nand U24200 (N_24200,N_22304,N_21719);
nand U24201 (N_24201,N_20106,N_21194);
and U24202 (N_24202,N_21300,N_20927);
or U24203 (N_24203,N_20500,N_21152);
and U24204 (N_24204,N_20555,N_21480);
and U24205 (N_24205,N_21169,N_20428);
xor U24206 (N_24206,N_20736,N_21838);
xor U24207 (N_24207,N_21510,N_22399);
nor U24208 (N_24208,N_21604,N_21832);
xnor U24209 (N_24209,N_20132,N_21228);
xor U24210 (N_24210,N_22044,N_20378);
nor U24211 (N_24211,N_22434,N_22066);
nand U24212 (N_24212,N_20028,N_21605);
and U24213 (N_24213,N_22372,N_21140);
and U24214 (N_24214,N_22076,N_21135);
xor U24215 (N_24215,N_22061,N_21207);
and U24216 (N_24216,N_22085,N_21698);
nor U24217 (N_24217,N_21260,N_20125);
nor U24218 (N_24218,N_21112,N_21506);
nor U24219 (N_24219,N_20840,N_20633);
or U24220 (N_24220,N_20720,N_20701);
nand U24221 (N_24221,N_22371,N_20386);
nand U24222 (N_24222,N_21453,N_20686);
xor U24223 (N_24223,N_21266,N_20385);
nor U24224 (N_24224,N_21483,N_22269);
nor U24225 (N_24225,N_20080,N_22289);
or U24226 (N_24226,N_20662,N_21199);
or U24227 (N_24227,N_21766,N_20568);
xnor U24228 (N_24228,N_21279,N_21012);
or U24229 (N_24229,N_20201,N_22103);
or U24230 (N_24230,N_21812,N_22032);
or U24231 (N_24231,N_21171,N_20009);
nor U24232 (N_24232,N_21463,N_20068);
nor U24233 (N_24233,N_21757,N_21305);
or U24234 (N_24234,N_21331,N_22004);
xor U24235 (N_24235,N_20758,N_21717);
or U24236 (N_24236,N_22451,N_20381);
nor U24237 (N_24237,N_20731,N_21522);
nor U24238 (N_24238,N_20295,N_20911);
xor U24239 (N_24239,N_21246,N_22292);
and U24240 (N_24240,N_20344,N_20849);
nor U24241 (N_24241,N_20098,N_21707);
or U24242 (N_24242,N_20473,N_20098);
nand U24243 (N_24243,N_20509,N_21327);
nand U24244 (N_24244,N_21576,N_21179);
nand U24245 (N_24245,N_22139,N_20764);
and U24246 (N_24246,N_21910,N_21684);
xor U24247 (N_24247,N_20040,N_21265);
or U24248 (N_24248,N_21944,N_21100);
nand U24249 (N_24249,N_21347,N_22093);
and U24250 (N_24250,N_20317,N_22210);
and U24251 (N_24251,N_20111,N_20298);
nand U24252 (N_24252,N_22460,N_20783);
and U24253 (N_24253,N_20254,N_21713);
nand U24254 (N_24254,N_22146,N_20156);
nand U24255 (N_24255,N_21544,N_20463);
nand U24256 (N_24256,N_21389,N_20264);
nand U24257 (N_24257,N_22433,N_20245);
xor U24258 (N_24258,N_20185,N_21923);
xnor U24259 (N_24259,N_20329,N_20191);
and U24260 (N_24260,N_20217,N_21784);
xnor U24261 (N_24261,N_20369,N_20665);
xnor U24262 (N_24262,N_22046,N_20204);
nand U24263 (N_24263,N_20262,N_21525);
nor U24264 (N_24264,N_20610,N_20274);
nor U24265 (N_24265,N_21908,N_22473);
or U24266 (N_24266,N_20286,N_20672);
and U24267 (N_24267,N_21674,N_20233);
xnor U24268 (N_24268,N_21753,N_20994);
nand U24269 (N_24269,N_20816,N_20170);
xnor U24270 (N_24270,N_20332,N_21784);
or U24271 (N_24271,N_22010,N_21321);
or U24272 (N_24272,N_22401,N_20201);
xor U24273 (N_24273,N_21378,N_22402);
nor U24274 (N_24274,N_22160,N_22188);
nor U24275 (N_24275,N_20726,N_20566);
xor U24276 (N_24276,N_21383,N_20293);
or U24277 (N_24277,N_20660,N_20395);
or U24278 (N_24278,N_21583,N_21733);
nand U24279 (N_24279,N_21933,N_21951);
nand U24280 (N_24280,N_21544,N_21386);
nand U24281 (N_24281,N_21035,N_22023);
or U24282 (N_24282,N_20736,N_20101);
xnor U24283 (N_24283,N_21071,N_20474);
or U24284 (N_24284,N_21119,N_20625);
and U24285 (N_24285,N_22195,N_21074);
xor U24286 (N_24286,N_22179,N_20351);
xnor U24287 (N_24287,N_20128,N_21398);
nor U24288 (N_24288,N_20075,N_20400);
and U24289 (N_24289,N_21717,N_20236);
xor U24290 (N_24290,N_20690,N_22158);
xor U24291 (N_24291,N_20710,N_21874);
or U24292 (N_24292,N_21736,N_21265);
xnor U24293 (N_24293,N_20619,N_21288);
and U24294 (N_24294,N_21061,N_21222);
nand U24295 (N_24295,N_21498,N_21816);
xor U24296 (N_24296,N_20597,N_20842);
xnor U24297 (N_24297,N_20596,N_21820);
and U24298 (N_24298,N_20142,N_20694);
or U24299 (N_24299,N_21402,N_21884);
or U24300 (N_24300,N_21021,N_21812);
xnor U24301 (N_24301,N_20932,N_21316);
or U24302 (N_24302,N_21936,N_20802);
xnor U24303 (N_24303,N_22119,N_21700);
nor U24304 (N_24304,N_21201,N_20498);
and U24305 (N_24305,N_21614,N_21406);
xnor U24306 (N_24306,N_21796,N_21800);
xor U24307 (N_24307,N_20013,N_21033);
nand U24308 (N_24308,N_21909,N_21584);
xnor U24309 (N_24309,N_22150,N_21352);
and U24310 (N_24310,N_21437,N_22048);
nor U24311 (N_24311,N_22279,N_20671);
xnor U24312 (N_24312,N_21858,N_21346);
and U24313 (N_24313,N_22478,N_21376);
nand U24314 (N_24314,N_21734,N_21176);
and U24315 (N_24315,N_22009,N_21834);
or U24316 (N_24316,N_20114,N_20718);
and U24317 (N_24317,N_20800,N_21641);
or U24318 (N_24318,N_20337,N_21892);
xor U24319 (N_24319,N_21041,N_21348);
nand U24320 (N_24320,N_20088,N_20795);
or U24321 (N_24321,N_22010,N_21055);
and U24322 (N_24322,N_21282,N_21556);
or U24323 (N_24323,N_22479,N_21187);
xor U24324 (N_24324,N_21507,N_21301);
nand U24325 (N_24325,N_21107,N_22374);
and U24326 (N_24326,N_20635,N_22272);
nor U24327 (N_24327,N_22217,N_20504);
nand U24328 (N_24328,N_22254,N_20491);
nor U24329 (N_24329,N_22271,N_21880);
nand U24330 (N_24330,N_21768,N_21248);
nand U24331 (N_24331,N_20042,N_22316);
or U24332 (N_24332,N_20060,N_21452);
or U24333 (N_24333,N_20188,N_21644);
and U24334 (N_24334,N_21922,N_20725);
xor U24335 (N_24335,N_20536,N_21652);
and U24336 (N_24336,N_21875,N_21264);
nand U24337 (N_24337,N_21144,N_21934);
xor U24338 (N_24338,N_20480,N_20783);
nand U24339 (N_24339,N_20083,N_22468);
xor U24340 (N_24340,N_21332,N_20381);
xnor U24341 (N_24341,N_21132,N_22480);
nor U24342 (N_24342,N_20178,N_20738);
nor U24343 (N_24343,N_20516,N_21328);
xnor U24344 (N_24344,N_20314,N_20391);
nor U24345 (N_24345,N_22309,N_21615);
nand U24346 (N_24346,N_21433,N_20815);
nor U24347 (N_24347,N_20742,N_20752);
nor U24348 (N_24348,N_22170,N_22346);
and U24349 (N_24349,N_20866,N_21598);
or U24350 (N_24350,N_21752,N_22150);
nand U24351 (N_24351,N_20560,N_21819);
and U24352 (N_24352,N_20799,N_21785);
nand U24353 (N_24353,N_21888,N_20179);
or U24354 (N_24354,N_20955,N_20002);
nand U24355 (N_24355,N_21311,N_22298);
nor U24356 (N_24356,N_21252,N_20328);
and U24357 (N_24357,N_21708,N_20210);
or U24358 (N_24358,N_20612,N_21852);
xor U24359 (N_24359,N_20278,N_22462);
nand U24360 (N_24360,N_21817,N_21893);
xor U24361 (N_24361,N_21894,N_21454);
and U24362 (N_24362,N_20723,N_20449);
nand U24363 (N_24363,N_21328,N_21954);
nor U24364 (N_24364,N_20458,N_22103);
nand U24365 (N_24365,N_20630,N_21259);
nand U24366 (N_24366,N_20224,N_21853);
nand U24367 (N_24367,N_20535,N_20447);
nand U24368 (N_24368,N_22030,N_20920);
or U24369 (N_24369,N_22150,N_22231);
or U24370 (N_24370,N_21417,N_20894);
nand U24371 (N_24371,N_20584,N_21068);
and U24372 (N_24372,N_22094,N_21081);
nand U24373 (N_24373,N_21620,N_21855);
and U24374 (N_24374,N_20471,N_21689);
and U24375 (N_24375,N_22119,N_22425);
and U24376 (N_24376,N_21422,N_22275);
nor U24377 (N_24377,N_21473,N_21690);
and U24378 (N_24378,N_21740,N_20609);
nand U24379 (N_24379,N_20341,N_21766);
nand U24380 (N_24380,N_20495,N_21601);
nor U24381 (N_24381,N_20578,N_21647);
xor U24382 (N_24382,N_20813,N_22285);
xor U24383 (N_24383,N_20991,N_21876);
and U24384 (N_24384,N_21952,N_20160);
or U24385 (N_24385,N_22167,N_21384);
xnor U24386 (N_24386,N_20499,N_21358);
nand U24387 (N_24387,N_21226,N_21367);
xnor U24388 (N_24388,N_22049,N_20817);
nand U24389 (N_24389,N_21052,N_20439);
and U24390 (N_24390,N_20595,N_22255);
and U24391 (N_24391,N_20809,N_21286);
xnor U24392 (N_24392,N_21332,N_22186);
and U24393 (N_24393,N_20795,N_20417);
nor U24394 (N_24394,N_22121,N_22407);
nand U24395 (N_24395,N_22272,N_20639);
nor U24396 (N_24396,N_20651,N_21837);
and U24397 (N_24397,N_20479,N_20144);
or U24398 (N_24398,N_20474,N_20685);
and U24399 (N_24399,N_20323,N_22372);
xor U24400 (N_24400,N_20926,N_21570);
xor U24401 (N_24401,N_22132,N_20888);
xor U24402 (N_24402,N_20691,N_22142);
xor U24403 (N_24403,N_22400,N_20118);
or U24404 (N_24404,N_21295,N_22069);
nor U24405 (N_24405,N_21749,N_20782);
xor U24406 (N_24406,N_20099,N_21622);
nor U24407 (N_24407,N_22037,N_20891);
nand U24408 (N_24408,N_22076,N_20120);
nand U24409 (N_24409,N_20886,N_20726);
xor U24410 (N_24410,N_22001,N_20288);
xnor U24411 (N_24411,N_22038,N_20643);
xnor U24412 (N_24412,N_21117,N_21364);
or U24413 (N_24413,N_21774,N_20149);
nor U24414 (N_24414,N_20355,N_22391);
nand U24415 (N_24415,N_20149,N_20109);
nor U24416 (N_24416,N_20431,N_21117);
nand U24417 (N_24417,N_21013,N_21677);
xor U24418 (N_24418,N_20116,N_20024);
and U24419 (N_24419,N_21240,N_21895);
nor U24420 (N_24420,N_20687,N_21498);
nand U24421 (N_24421,N_22102,N_20168);
or U24422 (N_24422,N_21265,N_20752);
and U24423 (N_24423,N_20775,N_21774);
nand U24424 (N_24424,N_20992,N_21069);
xnor U24425 (N_24425,N_21926,N_21424);
xor U24426 (N_24426,N_22445,N_20885);
nor U24427 (N_24427,N_21034,N_20660);
and U24428 (N_24428,N_20093,N_20462);
nor U24429 (N_24429,N_20582,N_21939);
nor U24430 (N_24430,N_21114,N_20376);
xnor U24431 (N_24431,N_21043,N_20768);
or U24432 (N_24432,N_21563,N_22096);
nand U24433 (N_24433,N_22117,N_21526);
nand U24434 (N_24434,N_21948,N_21157);
nand U24435 (N_24435,N_20951,N_22432);
or U24436 (N_24436,N_20030,N_21784);
xnor U24437 (N_24437,N_21608,N_20810);
nand U24438 (N_24438,N_20313,N_22424);
or U24439 (N_24439,N_20205,N_22465);
or U24440 (N_24440,N_20658,N_20940);
nand U24441 (N_24441,N_21951,N_21263);
xnor U24442 (N_24442,N_20351,N_22064);
nor U24443 (N_24443,N_20197,N_21242);
nor U24444 (N_24444,N_21422,N_21305);
and U24445 (N_24445,N_21314,N_22253);
xor U24446 (N_24446,N_20465,N_21997);
xor U24447 (N_24447,N_21504,N_20197);
xor U24448 (N_24448,N_22451,N_20191);
nor U24449 (N_24449,N_20216,N_20499);
xor U24450 (N_24450,N_21358,N_21248);
xor U24451 (N_24451,N_21651,N_22417);
xor U24452 (N_24452,N_22141,N_20351);
or U24453 (N_24453,N_20965,N_20570);
xor U24454 (N_24454,N_21497,N_21341);
nand U24455 (N_24455,N_20818,N_20665);
and U24456 (N_24456,N_20083,N_21447);
and U24457 (N_24457,N_21655,N_21586);
or U24458 (N_24458,N_22266,N_20774);
nor U24459 (N_24459,N_22299,N_21339);
nand U24460 (N_24460,N_20214,N_21918);
nand U24461 (N_24461,N_21056,N_21416);
nor U24462 (N_24462,N_21950,N_22269);
xnor U24463 (N_24463,N_20577,N_21906);
nor U24464 (N_24464,N_21529,N_21632);
nor U24465 (N_24465,N_20744,N_20137);
xor U24466 (N_24466,N_21615,N_22493);
nor U24467 (N_24467,N_21887,N_21959);
or U24468 (N_24468,N_22281,N_20201);
xnor U24469 (N_24469,N_21493,N_21738);
or U24470 (N_24470,N_21387,N_20479);
nor U24471 (N_24471,N_20780,N_22058);
or U24472 (N_24472,N_20954,N_21280);
or U24473 (N_24473,N_20252,N_21895);
nor U24474 (N_24474,N_21640,N_20682);
nand U24475 (N_24475,N_20639,N_20955);
xor U24476 (N_24476,N_22472,N_21059);
or U24477 (N_24477,N_20682,N_21988);
nand U24478 (N_24478,N_20726,N_20311);
nand U24479 (N_24479,N_21576,N_21359);
xnor U24480 (N_24480,N_22490,N_21928);
nand U24481 (N_24481,N_20892,N_20337);
and U24482 (N_24482,N_21488,N_21273);
nor U24483 (N_24483,N_21496,N_20816);
and U24484 (N_24484,N_21022,N_20868);
nor U24485 (N_24485,N_20262,N_22456);
nand U24486 (N_24486,N_21201,N_20462);
or U24487 (N_24487,N_21436,N_21210);
xnor U24488 (N_24488,N_22261,N_21323);
and U24489 (N_24489,N_21361,N_21885);
or U24490 (N_24490,N_20190,N_22472);
nor U24491 (N_24491,N_21297,N_21505);
or U24492 (N_24492,N_21706,N_20352);
and U24493 (N_24493,N_20131,N_21328);
nor U24494 (N_24494,N_21700,N_21486);
or U24495 (N_24495,N_22150,N_21153);
xnor U24496 (N_24496,N_22130,N_21704);
nor U24497 (N_24497,N_22387,N_21614);
nor U24498 (N_24498,N_20844,N_20777);
nor U24499 (N_24499,N_20936,N_20339);
or U24500 (N_24500,N_21586,N_20968);
or U24501 (N_24501,N_20057,N_20529);
or U24502 (N_24502,N_22396,N_20555);
and U24503 (N_24503,N_20585,N_21476);
xor U24504 (N_24504,N_20747,N_20215);
and U24505 (N_24505,N_21711,N_21138);
or U24506 (N_24506,N_22332,N_21778);
nand U24507 (N_24507,N_22164,N_22354);
xor U24508 (N_24508,N_21359,N_20480);
nand U24509 (N_24509,N_21091,N_20033);
and U24510 (N_24510,N_20064,N_22353);
nand U24511 (N_24511,N_20921,N_21429);
xor U24512 (N_24512,N_20377,N_20537);
nand U24513 (N_24513,N_20817,N_21083);
and U24514 (N_24514,N_21086,N_21372);
xor U24515 (N_24515,N_21618,N_21930);
or U24516 (N_24516,N_20999,N_20858);
xnor U24517 (N_24517,N_20853,N_21829);
xnor U24518 (N_24518,N_21805,N_20760);
nor U24519 (N_24519,N_20287,N_21894);
nand U24520 (N_24520,N_22435,N_21144);
and U24521 (N_24521,N_21181,N_20139);
nand U24522 (N_24522,N_20670,N_21976);
and U24523 (N_24523,N_22182,N_22122);
nor U24524 (N_24524,N_20321,N_21874);
xor U24525 (N_24525,N_20659,N_20025);
nand U24526 (N_24526,N_22090,N_21533);
and U24527 (N_24527,N_22086,N_21456);
nor U24528 (N_24528,N_20934,N_21816);
xor U24529 (N_24529,N_21389,N_20033);
xor U24530 (N_24530,N_20108,N_20811);
xor U24531 (N_24531,N_20935,N_22190);
or U24532 (N_24532,N_20368,N_20491);
nor U24533 (N_24533,N_21836,N_22116);
xor U24534 (N_24534,N_22375,N_20536);
or U24535 (N_24535,N_21635,N_20674);
xor U24536 (N_24536,N_21184,N_20489);
nand U24537 (N_24537,N_20057,N_20834);
or U24538 (N_24538,N_20164,N_22058);
and U24539 (N_24539,N_20451,N_20123);
xor U24540 (N_24540,N_21295,N_21584);
nand U24541 (N_24541,N_21195,N_21226);
nand U24542 (N_24542,N_20705,N_22466);
xnor U24543 (N_24543,N_22331,N_20912);
nand U24544 (N_24544,N_21355,N_22035);
xnor U24545 (N_24545,N_21051,N_20433);
and U24546 (N_24546,N_21970,N_20712);
nand U24547 (N_24547,N_22095,N_22359);
nor U24548 (N_24548,N_21280,N_20616);
and U24549 (N_24549,N_22165,N_21063);
or U24550 (N_24550,N_22325,N_22353);
xor U24551 (N_24551,N_22373,N_21860);
or U24552 (N_24552,N_22431,N_21679);
nor U24553 (N_24553,N_22352,N_20277);
xor U24554 (N_24554,N_21531,N_22137);
or U24555 (N_24555,N_21242,N_20745);
and U24556 (N_24556,N_22410,N_21449);
and U24557 (N_24557,N_21136,N_20520);
nor U24558 (N_24558,N_20341,N_21490);
nor U24559 (N_24559,N_21523,N_20482);
and U24560 (N_24560,N_22369,N_20876);
xnor U24561 (N_24561,N_21891,N_21567);
and U24562 (N_24562,N_20526,N_21623);
xnor U24563 (N_24563,N_20158,N_20697);
or U24564 (N_24564,N_22193,N_20807);
nor U24565 (N_24565,N_22217,N_22258);
xor U24566 (N_24566,N_20991,N_21680);
nand U24567 (N_24567,N_21383,N_22028);
or U24568 (N_24568,N_20294,N_22285);
and U24569 (N_24569,N_22260,N_20734);
or U24570 (N_24570,N_21288,N_22010);
xnor U24571 (N_24571,N_20616,N_20983);
nor U24572 (N_24572,N_21228,N_21574);
xor U24573 (N_24573,N_22124,N_21849);
and U24574 (N_24574,N_21909,N_20493);
nor U24575 (N_24575,N_22214,N_20010);
or U24576 (N_24576,N_22384,N_22217);
nor U24577 (N_24577,N_21430,N_22348);
and U24578 (N_24578,N_21825,N_21352);
nand U24579 (N_24579,N_20071,N_21585);
nor U24580 (N_24580,N_21694,N_22264);
xnor U24581 (N_24581,N_21374,N_21057);
xor U24582 (N_24582,N_20991,N_22359);
and U24583 (N_24583,N_20941,N_20043);
xor U24584 (N_24584,N_21184,N_21212);
nor U24585 (N_24585,N_20998,N_20312);
or U24586 (N_24586,N_20638,N_21312);
and U24587 (N_24587,N_20010,N_22270);
and U24588 (N_24588,N_20842,N_21032);
and U24589 (N_24589,N_22305,N_20672);
nor U24590 (N_24590,N_22475,N_20208);
and U24591 (N_24591,N_22410,N_21367);
or U24592 (N_24592,N_21568,N_20945);
xnor U24593 (N_24593,N_22445,N_20733);
nand U24594 (N_24594,N_21477,N_21338);
nand U24595 (N_24595,N_21259,N_22081);
and U24596 (N_24596,N_21516,N_22027);
and U24597 (N_24597,N_20748,N_21423);
and U24598 (N_24598,N_21159,N_22471);
or U24599 (N_24599,N_21943,N_21143);
xor U24600 (N_24600,N_20907,N_20281);
and U24601 (N_24601,N_20644,N_21664);
nand U24602 (N_24602,N_20901,N_20095);
xnor U24603 (N_24603,N_22084,N_20027);
or U24604 (N_24604,N_21190,N_20366);
nand U24605 (N_24605,N_22474,N_20612);
nor U24606 (N_24606,N_21206,N_21698);
or U24607 (N_24607,N_21685,N_21862);
nor U24608 (N_24608,N_20819,N_22142);
xor U24609 (N_24609,N_21951,N_21011);
xor U24610 (N_24610,N_22254,N_20611);
and U24611 (N_24611,N_21186,N_22359);
nor U24612 (N_24612,N_21957,N_20921);
xnor U24613 (N_24613,N_20569,N_20786);
xor U24614 (N_24614,N_22498,N_21195);
nor U24615 (N_24615,N_20344,N_22259);
or U24616 (N_24616,N_22071,N_20166);
nor U24617 (N_24617,N_20495,N_20578);
nor U24618 (N_24618,N_21162,N_21426);
or U24619 (N_24619,N_22127,N_21990);
xnor U24620 (N_24620,N_22373,N_22187);
nand U24621 (N_24621,N_21225,N_21583);
and U24622 (N_24622,N_22304,N_20818);
nand U24623 (N_24623,N_21219,N_22117);
nor U24624 (N_24624,N_21267,N_20190);
nor U24625 (N_24625,N_21018,N_20467);
or U24626 (N_24626,N_21356,N_20075);
nand U24627 (N_24627,N_20223,N_21103);
and U24628 (N_24628,N_22283,N_22126);
xnor U24629 (N_24629,N_20297,N_21188);
nor U24630 (N_24630,N_21670,N_22226);
nand U24631 (N_24631,N_22439,N_21620);
or U24632 (N_24632,N_20123,N_22241);
nand U24633 (N_24633,N_21634,N_21909);
nand U24634 (N_24634,N_22191,N_21840);
xnor U24635 (N_24635,N_22044,N_21344);
or U24636 (N_24636,N_22368,N_21490);
or U24637 (N_24637,N_20800,N_21333);
nand U24638 (N_24638,N_21563,N_22274);
xnor U24639 (N_24639,N_21908,N_20652);
nand U24640 (N_24640,N_20212,N_22279);
and U24641 (N_24641,N_21938,N_20914);
and U24642 (N_24642,N_20853,N_21184);
xor U24643 (N_24643,N_22186,N_21133);
and U24644 (N_24644,N_20672,N_20852);
nor U24645 (N_24645,N_21297,N_21993);
nor U24646 (N_24646,N_21318,N_21501);
xnor U24647 (N_24647,N_20734,N_20390);
xor U24648 (N_24648,N_20486,N_21768);
nand U24649 (N_24649,N_20312,N_22214);
or U24650 (N_24650,N_20754,N_21471);
nand U24651 (N_24651,N_22051,N_21477);
and U24652 (N_24652,N_21213,N_21227);
and U24653 (N_24653,N_22336,N_22363);
nor U24654 (N_24654,N_21164,N_20516);
and U24655 (N_24655,N_21932,N_20774);
or U24656 (N_24656,N_20508,N_22351);
nor U24657 (N_24657,N_20859,N_22359);
nor U24658 (N_24658,N_20948,N_20185);
xor U24659 (N_24659,N_21132,N_22114);
or U24660 (N_24660,N_20111,N_21572);
xor U24661 (N_24661,N_21828,N_21231);
nand U24662 (N_24662,N_20211,N_20005);
and U24663 (N_24663,N_20315,N_20578);
xnor U24664 (N_24664,N_22206,N_21780);
nor U24665 (N_24665,N_22365,N_22453);
nor U24666 (N_24666,N_20124,N_20370);
nand U24667 (N_24667,N_20464,N_20283);
or U24668 (N_24668,N_21421,N_21135);
xnor U24669 (N_24669,N_22036,N_20568);
nand U24670 (N_24670,N_22087,N_22215);
xor U24671 (N_24671,N_22251,N_20083);
or U24672 (N_24672,N_21265,N_20568);
and U24673 (N_24673,N_20878,N_20589);
nand U24674 (N_24674,N_20959,N_20257);
xnor U24675 (N_24675,N_20103,N_21787);
xnor U24676 (N_24676,N_20826,N_22033);
nor U24677 (N_24677,N_21501,N_21637);
nand U24678 (N_24678,N_22179,N_22019);
nor U24679 (N_24679,N_22147,N_21759);
nand U24680 (N_24680,N_21536,N_21344);
nand U24681 (N_24681,N_20772,N_21247);
nor U24682 (N_24682,N_20984,N_21999);
nor U24683 (N_24683,N_22375,N_20548);
nor U24684 (N_24684,N_21738,N_22086);
and U24685 (N_24685,N_21282,N_20347);
and U24686 (N_24686,N_21040,N_21592);
and U24687 (N_24687,N_21975,N_21268);
xnor U24688 (N_24688,N_20012,N_20348);
nor U24689 (N_24689,N_20502,N_20041);
nand U24690 (N_24690,N_21337,N_22046);
and U24691 (N_24691,N_22043,N_21933);
xnor U24692 (N_24692,N_21428,N_20786);
xor U24693 (N_24693,N_22249,N_21894);
nor U24694 (N_24694,N_20554,N_20029);
or U24695 (N_24695,N_20021,N_20664);
nand U24696 (N_24696,N_22350,N_22030);
nand U24697 (N_24697,N_21349,N_21423);
or U24698 (N_24698,N_20408,N_22205);
nor U24699 (N_24699,N_22445,N_22341);
nor U24700 (N_24700,N_21019,N_21380);
nand U24701 (N_24701,N_22154,N_20627);
nor U24702 (N_24702,N_22298,N_20678);
nor U24703 (N_24703,N_22162,N_21901);
xor U24704 (N_24704,N_22323,N_20451);
nand U24705 (N_24705,N_21021,N_21271);
nor U24706 (N_24706,N_22075,N_21637);
nor U24707 (N_24707,N_20095,N_20162);
xnor U24708 (N_24708,N_21129,N_21477);
and U24709 (N_24709,N_22167,N_22224);
and U24710 (N_24710,N_21669,N_22193);
nor U24711 (N_24711,N_22485,N_22074);
nand U24712 (N_24712,N_21056,N_21068);
nand U24713 (N_24713,N_21111,N_20964);
and U24714 (N_24714,N_22252,N_21759);
and U24715 (N_24715,N_21474,N_20883);
xor U24716 (N_24716,N_20708,N_20944);
nor U24717 (N_24717,N_21359,N_22423);
xor U24718 (N_24718,N_21969,N_22193);
nand U24719 (N_24719,N_20248,N_21642);
xnor U24720 (N_24720,N_22491,N_22370);
xor U24721 (N_24721,N_21756,N_21688);
or U24722 (N_24722,N_21075,N_21941);
xnor U24723 (N_24723,N_21052,N_21558);
nor U24724 (N_24724,N_20940,N_21238);
nand U24725 (N_24725,N_20022,N_20153);
nor U24726 (N_24726,N_21693,N_21877);
and U24727 (N_24727,N_22433,N_20887);
nor U24728 (N_24728,N_22294,N_20499);
nand U24729 (N_24729,N_22152,N_22494);
or U24730 (N_24730,N_20243,N_21740);
xor U24731 (N_24731,N_20867,N_20475);
nand U24732 (N_24732,N_22380,N_20413);
xnor U24733 (N_24733,N_20511,N_21792);
nand U24734 (N_24734,N_21912,N_20642);
and U24735 (N_24735,N_20963,N_20528);
or U24736 (N_24736,N_21225,N_20946);
or U24737 (N_24737,N_20642,N_22463);
and U24738 (N_24738,N_20113,N_20138);
nand U24739 (N_24739,N_21618,N_20623);
nand U24740 (N_24740,N_21580,N_21494);
or U24741 (N_24741,N_22444,N_20138);
nor U24742 (N_24742,N_21007,N_20024);
xnor U24743 (N_24743,N_22444,N_20199);
and U24744 (N_24744,N_22117,N_22283);
xnor U24745 (N_24745,N_20754,N_21598);
nor U24746 (N_24746,N_22428,N_20682);
and U24747 (N_24747,N_21849,N_20896);
and U24748 (N_24748,N_21336,N_21755);
nor U24749 (N_24749,N_20133,N_21185);
or U24750 (N_24750,N_20733,N_20538);
nor U24751 (N_24751,N_21540,N_21729);
and U24752 (N_24752,N_20204,N_20256);
xnor U24753 (N_24753,N_20787,N_22403);
xnor U24754 (N_24754,N_20225,N_21721);
nand U24755 (N_24755,N_20910,N_20975);
nor U24756 (N_24756,N_20903,N_21245);
nand U24757 (N_24757,N_21569,N_21355);
nand U24758 (N_24758,N_20318,N_20866);
nor U24759 (N_24759,N_22494,N_22068);
or U24760 (N_24760,N_20362,N_20743);
nor U24761 (N_24761,N_20718,N_20497);
or U24762 (N_24762,N_20180,N_20891);
xor U24763 (N_24763,N_21169,N_21751);
nand U24764 (N_24764,N_20512,N_21870);
and U24765 (N_24765,N_20198,N_21654);
nand U24766 (N_24766,N_20440,N_21454);
or U24767 (N_24767,N_22125,N_22327);
nor U24768 (N_24768,N_20963,N_20096);
or U24769 (N_24769,N_21628,N_21706);
or U24770 (N_24770,N_22101,N_20941);
nand U24771 (N_24771,N_22160,N_20832);
or U24772 (N_24772,N_20595,N_20224);
and U24773 (N_24773,N_21548,N_20225);
nand U24774 (N_24774,N_20104,N_21612);
nand U24775 (N_24775,N_20696,N_21827);
nor U24776 (N_24776,N_20390,N_20586);
and U24777 (N_24777,N_22043,N_20106);
or U24778 (N_24778,N_21594,N_21382);
xnor U24779 (N_24779,N_21297,N_20258);
nor U24780 (N_24780,N_21570,N_21019);
xor U24781 (N_24781,N_20225,N_21926);
xnor U24782 (N_24782,N_20789,N_22332);
nor U24783 (N_24783,N_21851,N_21749);
xor U24784 (N_24784,N_21967,N_21684);
or U24785 (N_24785,N_20976,N_22397);
xnor U24786 (N_24786,N_21107,N_20734);
nand U24787 (N_24787,N_20537,N_20482);
and U24788 (N_24788,N_20704,N_22231);
or U24789 (N_24789,N_20491,N_21030);
or U24790 (N_24790,N_20944,N_22365);
nand U24791 (N_24791,N_21121,N_21042);
or U24792 (N_24792,N_21804,N_20810);
or U24793 (N_24793,N_20030,N_20534);
and U24794 (N_24794,N_22014,N_21182);
and U24795 (N_24795,N_21514,N_21932);
xor U24796 (N_24796,N_21815,N_22283);
or U24797 (N_24797,N_20118,N_20556);
nor U24798 (N_24798,N_22151,N_22073);
nand U24799 (N_24799,N_20121,N_21185);
or U24800 (N_24800,N_20562,N_22248);
nor U24801 (N_24801,N_21584,N_22155);
or U24802 (N_24802,N_21130,N_21624);
nand U24803 (N_24803,N_21306,N_20735);
or U24804 (N_24804,N_21714,N_21822);
nor U24805 (N_24805,N_21570,N_20719);
nand U24806 (N_24806,N_20580,N_20026);
and U24807 (N_24807,N_21138,N_20521);
xnor U24808 (N_24808,N_21549,N_22210);
nand U24809 (N_24809,N_21231,N_22103);
nand U24810 (N_24810,N_21883,N_21848);
or U24811 (N_24811,N_21648,N_20014);
and U24812 (N_24812,N_22308,N_22336);
or U24813 (N_24813,N_20791,N_21962);
xor U24814 (N_24814,N_21098,N_22419);
nand U24815 (N_24815,N_22100,N_20274);
xnor U24816 (N_24816,N_20145,N_21207);
or U24817 (N_24817,N_20514,N_20172);
or U24818 (N_24818,N_20960,N_20198);
xnor U24819 (N_24819,N_21370,N_21693);
xnor U24820 (N_24820,N_20347,N_21855);
or U24821 (N_24821,N_21712,N_21506);
xor U24822 (N_24822,N_21058,N_21607);
and U24823 (N_24823,N_21295,N_20709);
and U24824 (N_24824,N_21650,N_21256);
and U24825 (N_24825,N_20309,N_21008);
or U24826 (N_24826,N_21567,N_21322);
xor U24827 (N_24827,N_20365,N_20991);
nor U24828 (N_24828,N_21006,N_21084);
nor U24829 (N_24829,N_21397,N_21471);
xor U24830 (N_24830,N_22278,N_21232);
nor U24831 (N_24831,N_21521,N_21212);
xnor U24832 (N_24832,N_21437,N_20065);
xor U24833 (N_24833,N_20643,N_20454);
nor U24834 (N_24834,N_20600,N_21984);
nor U24835 (N_24835,N_21149,N_20926);
or U24836 (N_24836,N_21975,N_20786);
xnor U24837 (N_24837,N_20995,N_20185);
xnor U24838 (N_24838,N_21982,N_21551);
nor U24839 (N_24839,N_22468,N_22359);
or U24840 (N_24840,N_21856,N_21163);
and U24841 (N_24841,N_20040,N_21225);
nand U24842 (N_24842,N_22182,N_20073);
or U24843 (N_24843,N_20395,N_21417);
nand U24844 (N_24844,N_20507,N_21513);
nor U24845 (N_24845,N_22206,N_22227);
xor U24846 (N_24846,N_20847,N_22463);
xnor U24847 (N_24847,N_20781,N_20583);
xor U24848 (N_24848,N_22448,N_21809);
nand U24849 (N_24849,N_21956,N_21390);
nand U24850 (N_24850,N_22175,N_20763);
nor U24851 (N_24851,N_20834,N_21767);
or U24852 (N_24852,N_20832,N_22024);
or U24853 (N_24853,N_22191,N_20623);
nand U24854 (N_24854,N_20177,N_20396);
nor U24855 (N_24855,N_22484,N_20834);
and U24856 (N_24856,N_21963,N_20744);
and U24857 (N_24857,N_20325,N_21964);
and U24858 (N_24858,N_21202,N_21150);
nor U24859 (N_24859,N_20008,N_20592);
nand U24860 (N_24860,N_21252,N_20596);
nand U24861 (N_24861,N_20801,N_21915);
xor U24862 (N_24862,N_22183,N_20702);
xnor U24863 (N_24863,N_20533,N_21213);
nand U24864 (N_24864,N_20190,N_20841);
and U24865 (N_24865,N_22289,N_20471);
or U24866 (N_24866,N_22334,N_21907);
or U24867 (N_24867,N_20695,N_21053);
nand U24868 (N_24868,N_21961,N_22027);
nand U24869 (N_24869,N_21671,N_21366);
xnor U24870 (N_24870,N_21152,N_21901);
nand U24871 (N_24871,N_20259,N_20047);
or U24872 (N_24872,N_20215,N_20818);
xor U24873 (N_24873,N_20658,N_20645);
nand U24874 (N_24874,N_20040,N_22309);
nand U24875 (N_24875,N_21358,N_21589);
nand U24876 (N_24876,N_20203,N_21280);
xnor U24877 (N_24877,N_20326,N_20300);
nor U24878 (N_24878,N_21785,N_20690);
and U24879 (N_24879,N_21206,N_20785);
nand U24880 (N_24880,N_21105,N_22305);
nand U24881 (N_24881,N_22026,N_21708);
nand U24882 (N_24882,N_22494,N_20399);
and U24883 (N_24883,N_20837,N_22143);
or U24884 (N_24884,N_20020,N_20987);
or U24885 (N_24885,N_21590,N_21720);
xor U24886 (N_24886,N_21187,N_22164);
nor U24887 (N_24887,N_22141,N_21716);
nor U24888 (N_24888,N_20970,N_20991);
xor U24889 (N_24889,N_20133,N_22312);
xor U24890 (N_24890,N_20885,N_21259);
xor U24891 (N_24891,N_21092,N_22415);
nor U24892 (N_24892,N_20066,N_21018);
or U24893 (N_24893,N_20456,N_20250);
nor U24894 (N_24894,N_21022,N_20489);
xor U24895 (N_24895,N_20053,N_21564);
and U24896 (N_24896,N_21468,N_20519);
nor U24897 (N_24897,N_20167,N_20491);
nand U24898 (N_24898,N_22129,N_22283);
or U24899 (N_24899,N_20114,N_20516);
and U24900 (N_24900,N_20171,N_21235);
nand U24901 (N_24901,N_20623,N_22183);
and U24902 (N_24902,N_22059,N_21398);
and U24903 (N_24903,N_21110,N_20089);
nand U24904 (N_24904,N_21317,N_21894);
nor U24905 (N_24905,N_22361,N_20167);
or U24906 (N_24906,N_21487,N_22034);
nand U24907 (N_24907,N_22081,N_21815);
or U24908 (N_24908,N_22298,N_20891);
and U24909 (N_24909,N_22150,N_22123);
and U24910 (N_24910,N_22072,N_22397);
or U24911 (N_24911,N_22161,N_21167);
or U24912 (N_24912,N_21853,N_20478);
nand U24913 (N_24913,N_22219,N_22200);
nand U24914 (N_24914,N_20849,N_20245);
xnor U24915 (N_24915,N_21569,N_20065);
nand U24916 (N_24916,N_20018,N_20315);
nand U24917 (N_24917,N_20772,N_22144);
nand U24918 (N_24918,N_21211,N_22418);
xnor U24919 (N_24919,N_20399,N_20921);
or U24920 (N_24920,N_21160,N_21106);
nand U24921 (N_24921,N_21709,N_20336);
nor U24922 (N_24922,N_21334,N_20146);
xor U24923 (N_24923,N_22471,N_20588);
nand U24924 (N_24924,N_20800,N_21940);
xor U24925 (N_24925,N_21081,N_20356);
or U24926 (N_24926,N_20453,N_22358);
xor U24927 (N_24927,N_20524,N_20729);
nor U24928 (N_24928,N_20395,N_21163);
or U24929 (N_24929,N_22035,N_22145);
or U24930 (N_24930,N_20991,N_20239);
nand U24931 (N_24931,N_21725,N_20159);
nand U24932 (N_24932,N_22484,N_20963);
nor U24933 (N_24933,N_20398,N_22189);
nand U24934 (N_24934,N_22008,N_21550);
xor U24935 (N_24935,N_21690,N_22225);
or U24936 (N_24936,N_21794,N_22345);
xor U24937 (N_24937,N_20108,N_22407);
or U24938 (N_24938,N_20154,N_21587);
nor U24939 (N_24939,N_21953,N_20616);
or U24940 (N_24940,N_20238,N_21109);
xor U24941 (N_24941,N_22368,N_22481);
and U24942 (N_24942,N_21241,N_20126);
nor U24943 (N_24943,N_20455,N_20128);
xnor U24944 (N_24944,N_21811,N_20139);
nor U24945 (N_24945,N_20532,N_21114);
nand U24946 (N_24946,N_20166,N_22058);
and U24947 (N_24947,N_20155,N_21216);
or U24948 (N_24948,N_22002,N_20620);
or U24949 (N_24949,N_21583,N_20008);
or U24950 (N_24950,N_20079,N_20789);
nor U24951 (N_24951,N_21755,N_21790);
xnor U24952 (N_24952,N_20982,N_20662);
nor U24953 (N_24953,N_22490,N_21318);
nor U24954 (N_24954,N_21613,N_22356);
nand U24955 (N_24955,N_21735,N_21296);
or U24956 (N_24956,N_22212,N_21696);
and U24957 (N_24957,N_20228,N_21889);
or U24958 (N_24958,N_20511,N_20861);
and U24959 (N_24959,N_21646,N_20257);
or U24960 (N_24960,N_22417,N_20968);
or U24961 (N_24961,N_21209,N_20415);
or U24962 (N_24962,N_21491,N_22333);
xor U24963 (N_24963,N_20376,N_20601);
xor U24964 (N_24964,N_22453,N_22188);
or U24965 (N_24965,N_21076,N_20861);
nor U24966 (N_24966,N_22130,N_21468);
nand U24967 (N_24967,N_20614,N_20054);
nand U24968 (N_24968,N_20989,N_22289);
xnor U24969 (N_24969,N_20209,N_21878);
or U24970 (N_24970,N_20128,N_21875);
nor U24971 (N_24971,N_20344,N_21642);
or U24972 (N_24972,N_20337,N_21784);
nor U24973 (N_24973,N_22474,N_21591);
nand U24974 (N_24974,N_21975,N_20180);
nand U24975 (N_24975,N_21030,N_22468);
xor U24976 (N_24976,N_20885,N_21012);
xnor U24977 (N_24977,N_20372,N_20210);
xor U24978 (N_24978,N_22213,N_20657);
xnor U24979 (N_24979,N_21574,N_20599);
nor U24980 (N_24980,N_22390,N_21831);
nor U24981 (N_24981,N_20427,N_21968);
nand U24982 (N_24982,N_20376,N_20122);
nor U24983 (N_24983,N_20195,N_20941);
or U24984 (N_24984,N_21275,N_20869);
and U24985 (N_24985,N_21956,N_20957);
nand U24986 (N_24986,N_20444,N_20553);
nor U24987 (N_24987,N_20153,N_22377);
nor U24988 (N_24988,N_22369,N_20489);
and U24989 (N_24989,N_21456,N_22186);
or U24990 (N_24990,N_20791,N_20269);
or U24991 (N_24991,N_20122,N_21051);
xor U24992 (N_24992,N_21806,N_21757);
xor U24993 (N_24993,N_21980,N_21339);
nand U24994 (N_24994,N_21485,N_20256);
xnor U24995 (N_24995,N_22249,N_21974);
nor U24996 (N_24996,N_20597,N_21409);
and U24997 (N_24997,N_21062,N_21725);
or U24998 (N_24998,N_21189,N_21960);
nor U24999 (N_24999,N_20807,N_22002);
xnor UO_0 (O_0,N_24392,N_23227);
and UO_1 (O_1,N_24568,N_24286);
nand UO_2 (O_2,N_23148,N_24034);
nor UO_3 (O_3,N_24586,N_23353);
xor UO_4 (O_4,N_24380,N_23722);
or UO_5 (O_5,N_24203,N_23214);
nor UO_6 (O_6,N_23428,N_23316);
or UO_7 (O_7,N_22989,N_24759);
or UO_8 (O_8,N_23398,N_24545);
nand UO_9 (O_9,N_23321,N_23642);
xor UO_10 (O_10,N_22919,N_22986);
or UO_11 (O_11,N_24028,N_24997);
or UO_12 (O_12,N_24009,N_23651);
nand UO_13 (O_13,N_24577,N_23129);
or UO_14 (O_14,N_22605,N_24958);
and UO_15 (O_15,N_23328,N_23436);
xor UO_16 (O_16,N_23077,N_24030);
or UO_17 (O_17,N_24957,N_23983);
nor UO_18 (O_18,N_23828,N_23183);
xnor UO_19 (O_19,N_23569,N_23528);
and UO_20 (O_20,N_24932,N_23880);
nand UO_21 (O_21,N_24664,N_24907);
or UO_22 (O_22,N_24388,N_24963);
nand UO_23 (O_23,N_23974,N_24744);
and UO_24 (O_24,N_23846,N_24233);
xor UO_25 (O_25,N_24757,N_23351);
nand UO_26 (O_26,N_24273,N_22964);
nor UO_27 (O_27,N_23993,N_24040);
xor UO_28 (O_28,N_23422,N_23478);
xnor UO_29 (O_29,N_23168,N_24599);
nor UO_30 (O_30,N_24775,N_23190);
or UO_31 (O_31,N_23742,N_22898);
nor UO_32 (O_32,N_23821,N_24947);
or UO_33 (O_33,N_22563,N_23845);
nand UO_34 (O_34,N_24204,N_23242);
xor UO_35 (O_35,N_23295,N_24548);
nor UO_36 (O_36,N_24184,N_22994);
nand UO_37 (O_37,N_24588,N_23061);
or UO_38 (O_38,N_23411,N_24235);
nor UO_39 (O_39,N_23103,N_23511);
nor UO_40 (O_40,N_24325,N_24736);
or UO_41 (O_41,N_22777,N_23648);
xnor UO_42 (O_42,N_22683,N_24319);
xor UO_43 (O_43,N_24955,N_24129);
nor UO_44 (O_44,N_23432,N_24227);
xnor UO_45 (O_45,N_24027,N_23093);
and UO_46 (O_46,N_24169,N_24376);
xor UO_47 (O_47,N_24180,N_23581);
and UO_48 (O_48,N_23171,N_24289);
nand UO_49 (O_49,N_24343,N_23583);
nor UO_50 (O_50,N_24124,N_22584);
nor UO_51 (O_51,N_24277,N_22589);
xnor UO_52 (O_52,N_24991,N_24080);
nor UO_53 (O_53,N_24979,N_24803);
nor UO_54 (O_54,N_23865,N_22999);
or UO_55 (O_55,N_23289,N_23716);
and UO_56 (O_56,N_23764,N_23650);
or UO_57 (O_57,N_23453,N_22951);
xnor UO_58 (O_58,N_24906,N_23735);
nand UO_59 (O_59,N_23065,N_24560);
nor UO_60 (O_60,N_23384,N_22567);
and UO_61 (O_61,N_23693,N_23258);
xnor UO_62 (O_62,N_22914,N_23039);
or UO_63 (O_63,N_23607,N_24996);
nor UO_64 (O_64,N_23813,N_23443);
or UO_65 (O_65,N_23074,N_22513);
and UO_66 (O_66,N_24142,N_22514);
and UO_67 (O_67,N_23775,N_22786);
xor UO_68 (O_68,N_24770,N_24147);
or UO_69 (O_69,N_24972,N_24240);
and UO_70 (O_70,N_24182,N_23773);
nor UO_71 (O_71,N_23133,N_24054);
xnor UO_72 (O_72,N_23445,N_24778);
xor UO_73 (O_73,N_22834,N_22782);
nand UO_74 (O_74,N_23255,N_24871);
nand UO_75 (O_75,N_22756,N_24818);
xnor UO_76 (O_76,N_23842,N_22798);
nor UO_77 (O_77,N_23456,N_24158);
nand UO_78 (O_78,N_23799,N_23405);
nand UO_79 (O_79,N_23926,N_23052);
nor UO_80 (O_80,N_23404,N_23355);
nor UO_81 (O_81,N_23504,N_24475);
xnor UO_82 (O_82,N_22873,N_23394);
nor UO_83 (O_83,N_24107,N_23236);
nand UO_84 (O_84,N_23386,N_22506);
nand UO_85 (O_85,N_23507,N_24318);
nand UO_86 (O_86,N_22721,N_23347);
nor UO_87 (O_87,N_23348,N_24843);
and UO_88 (O_88,N_23589,N_22717);
nor UO_89 (O_89,N_24667,N_23446);
nor UO_90 (O_90,N_23667,N_23248);
or UO_91 (O_91,N_24193,N_22807);
xnor UO_92 (O_92,N_24780,N_24581);
or UO_93 (O_93,N_22733,N_22830);
nand UO_94 (O_94,N_23984,N_24561);
or UO_95 (O_95,N_23162,N_22885);
nand UO_96 (O_96,N_23068,N_22823);
nand UO_97 (O_97,N_23379,N_23803);
xnor UO_98 (O_98,N_24353,N_22858);
xor UO_99 (O_99,N_23125,N_24503);
and UO_100 (O_100,N_22825,N_24970);
nor UO_101 (O_101,N_23469,N_24317);
or UO_102 (O_102,N_24373,N_24303);
or UO_103 (O_103,N_24709,N_23201);
nor UO_104 (O_104,N_24478,N_22536);
nor UO_105 (O_105,N_23225,N_22525);
and UO_106 (O_106,N_24883,N_24562);
and UO_107 (O_107,N_23450,N_23408);
or UO_108 (O_108,N_24648,N_24713);
or UO_109 (O_109,N_23085,N_23585);
or UO_110 (O_110,N_23466,N_24519);
or UO_111 (O_111,N_22620,N_23892);
nand UO_112 (O_112,N_22663,N_23043);
nor UO_113 (O_113,N_24364,N_24755);
xor UO_114 (O_114,N_24569,N_22517);
nor UO_115 (O_115,N_23186,N_24237);
and UO_116 (O_116,N_24938,N_23151);
and UO_117 (O_117,N_22680,N_24062);
and UO_118 (O_118,N_24653,N_24333);
nor UO_119 (O_119,N_24496,N_24804);
nand UO_120 (O_120,N_22857,N_23646);
nand UO_121 (O_121,N_23196,N_23529);
xor UO_122 (O_122,N_24461,N_22741);
and UO_123 (O_123,N_24149,N_24377);
nor UO_124 (O_124,N_23672,N_24059);
xor UO_125 (O_125,N_22634,N_23914);
nor UO_126 (O_126,N_24595,N_24647);
nor UO_127 (O_127,N_22938,N_22572);
xor UO_128 (O_128,N_24490,N_23496);
xor UO_129 (O_129,N_23657,N_24742);
and UO_130 (O_130,N_22688,N_23666);
nand UO_131 (O_131,N_23038,N_23200);
or UO_132 (O_132,N_23671,N_23013);
nor UO_133 (O_133,N_23895,N_24756);
nand UO_134 (O_134,N_23156,N_23717);
and UO_135 (O_135,N_24911,N_24155);
or UO_136 (O_136,N_24265,N_24630);
nor UO_137 (O_137,N_24557,N_24251);
and UO_138 (O_138,N_24596,N_24181);
and UO_139 (O_139,N_23855,N_23545);
and UO_140 (O_140,N_23574,N_23121);
and UO_141 (O_141,N_24567,N_22615);
or UO_142 (O_142,N_23661,N_24532);
xnor UO_143 (O_143,N_23229,N_22690);
and UO_144 (O_144,N_22578,N_24481);
nor UO_145 (O_145,N_24716,N_23972);
nand UO_146 (O_146,N_24146,N_24666);
or UO_147 (O_147,N_23866,N_24914);
xor UO_148 (O_148,N_22622,N_24872);
and UO_149 (O_149,N_24224,N_23669);
and UO_150 (O_150,N_24538,N_24448);
xor UO_151 (O_151,N_23305,N_23461);
nand UO_152 (O_152,N_24086,N_22806);
or UO_153 (O_153,N_24899,N_23290);
and UO_154 (O_154,N_23425,N_22993);
nand UO_155 (O_155,N_24805,N_24572);
and UO_156 (O_156,N_24305,N_24156);
nand UO_157 (O_157,N_22743,N_24084);
nand UO_158 (O_158,N_24247,N_24882);
nand UO_159 (O_159,N_24358,N_24624);
nand UO_160 (O_160,N_22776,N_24485);
nand UO_161 (O_161,N_23144,N_24405);
or UO_162 (O_162,N_23877,N_24992);
or UO_163 (O_163,N_23811,N_24801);
nor UO_164 (O_164,N_23096,N_23746);
and UO_165 (O_165,N_23870,N_24998);
xor UO_166 (O_166,N_24593,N_23170);
and UO_167 (O_167,N_24681,N_24762);
nor UO_168 (O_168,N_23680,N_23908);
xnor UO_169 (O_169,N_22770,N_22939);
and UO_170 (O_170,N_24454,N_23415);
nor UO_171 (O_171,N_23387,N_23276);
nand UO_172 (O_172,N_22509,N_22828);
nor UO_173 (O_173,N_24937,N_23356);
nand UO_174 (O_174,N_23596,N_23910);
nor UO_175 (O_175,N_22793,N_23766);
and UO_176 (O_176,N_24087,N_24296);
nor UO_177 (O_177,N_23303,N_24961);
or UO_178 (O_178,N_24437,N_22976);
nor UO_179 (O_179,N_23844,N_24311);
and UO_180 (O_180,N_22610,N_24608);
nor UO_181 (O_181,N_22607,N_23304);
and UO_182 (O_182,N_22655,N_22730);
xor UO_183 (O_183,N_23023,N_23288);
nand UO_184 (O_184,N_22520,N_24137);
or UO_185 (O_185,N_22719,N_23904);
and UO_186 (O_186,N_23221,N_23881);
or UO_187 (O_187,N_24017,N_22819);
and UO_188 (O_188,N_22501,N_22727);
xnor UO_189 (O_189,N_23262,N_22987);
and UO_190 (O_190,N_24931,N_23176);
xor UO_191 (O_191,N_22712,N_24290);
or UO_192 (O_192,N_24426,N_24109);
or UO_193 (O_193,N_22542,N_24642);
xor UO_194 (O_194,N_23861,N_24293);
xnor UO_195 (O_195,N_23978,N_24272);
nor UO_196 (O_196,N_23625,N_23640);
xor UO_197 (O_197,N_23774,N_24045);
and UO_198 (O_198,N_24603,N_24754);
nor UO_199 (O_199,N_24400,N_23518);
and UO_200 (O_200,N_24993,N_24051);
and UO_201 (O_201,N_24795,N_24006);
nand UO_202 (O_202,N_23948,N_22748);
nor UO_203 (O_203,N_24005,N_23677);
nor UO_204 (O_204,N_24316,N_23543);
nand UO_205 (O_205,N_23195,N_23638);
nor UO_206 (O_206,N_24302,N_24238);
and UO_207 (O_207,N_22991,N_24905);
xor UO_208 (O_208,N_24786,N_24597);
and UO_209 (O_209,N_22720,N_24877);
nand UO_210 (O_210,N_24347,N_23519);
nand UO_211 (O_211,N_22639,N_24619);
or UO_212 (O_212,N_23956,N_23718);
nor UO_213 (O_213,N_22995,N_24835);
xor UO_214 (O_214,N_24055,N_24357);
xor UO_215 (O_215,N_23653,N_24136);
or UO_216 (O_216,N_23600,N_24760);
and UO_217 (O_217,N_23857,N_23191);
or UO_218 (O_218,N_23423,N_23066);
xor UO_219 (O_219,N_24611,N_23831);
nand UO_220 (O_220,N_23772,N_23322);
xor UO_221 (O_221,N_24585,N_24328);
and UO_222 (O_222,N_23198,N_22626);
or UO_223 (O_223,N_24102,N_24342);
and UO_224 (O_224,N_24960,N_23980);
and UO_225 (O_225,N_23476,N_23138);
or UO_226 (O_226,N_24999,N_22836);
nor UO_227 (O_227,N_23726,N_22545);
and UO_228 (O_228,N_23101,N_23762);
or UO_229 (O_229,N_24528,N_22670);
nand UO_230 (O_230,N_23498,N_23070);
nor UO_231 (O_231,N_24480,N_23576);
or UO_232 (O_232,N_24032,N_23577);
or UO_233 (O_233,N_23879,N_24816);
and UO_234 (O_234,N_24408,N_23922);
nand UO_235 (O_235,N_24679,N_24458);
xor UO_236 (O_236,N_23682,N_24913);
xor UO_237 (O_237,N_24120,N_24476);
nand UO_238 (O_238,N_23142,N_23494);
nand UO_239 (O_239,N_24135,N_24811);
nand UO_240 (O_240,N_24799,N_22903);
and UO_241 (O_241,N_23790,N_22551);
xnor UO_242 (O_242,N_23829,N_24011);
or UO_243 (O_243,N_22621,N_24506);
or UO_244 (O_244,N_23327,N_23343);
or UO_245 (O_245,N_22702,N_23439);
nor UO_246 (O_246,N_22638,N_24723);
xor UO_247 (O_247,N_24399,N_22511);
xor UO_248 (O_248,N_23767,N_24640);
and UO_249 (O_249,N_24049,N_22664);
or UO_250 (O_250,N_23301,N_24896);
and UO_251 (O_251,N_24351,N_23929);
nand UO_252 (O_252,N_24749,N_22869);
or UO_253 (O_253,N_24923,N_24382);
and UO_254 (O_254,N_24815,N_24675);
xor UO_255 (O_255,N_23024,N_23570);
xor UO_256 (O_256,N_23707,N_23639);
xnor UO_257 (O_257,N_24887,N_22791);
xor UO_258 (O_258,N_22848,N_22967);
or UO_259 (O_259,N_24101,N_24719);
or UO_260 (O_260,N_24607,N_24985);
nand UO_261 (O_261,N_23234,N_24910);
and UO_262 (O_262,N_22515,N_24518);
nand UO_263 (O_263,N_22636,N_24665);
xnor UO_264 (O_264,N_23155,N_23034);
and UO_265 (O_265,N_23223,N_23256);
xor UO_266 (O_266,N_23678,N_24278);
xnor UO_267 (O_267,N_22788,N_24326);
or UO_268 (O_268,N_23104,N_24340);
and UO_269 (O_269,N_22523,N_24209);
nor UO_270 (O_270,N_22594,N_23560);
or UO_271 (O_271,N_24922,N_22805);
nand UO_272 (O_272,N_23952,N_24023);
and UO_273 (O_273,N_23783,N_24934);
xor UO_274 (O_274,N_24618,N_24785);
and UO_275 (O_275,N_23864,N_24982);
nand UO_276 (O_276,N_23624,N_23284);
xor UO_277 (O_277,N_24151,N_23184);
and UO_278 (O_278,N_23481,N_22765);
nor UO_279 (O_279,N_23614,N_23662);
nand UO_280 (O_280,N_23324,N_23711);
nand UO_281 (O_281,N_23503,N_22998);
or UO_282 (O_282,N_24442,N_23369);
and UO_283 (O_283,N_23297,N_24254);
nor UO_284 (O_284,N_24003,N_24916);
nand UO_285 (O_285,N_24256,N_23032);
or UO_286 (O_286,N_23098,N_23599);
nand UO_287 (O_287,N_24395,N_23704);
and UO_288 (O_288,N_24735,N_24660);
nor UO_289 (O_289,N_24796,N_24867);
or UO_290 (O_290,N_24188,N_24178);
xor UO_291 (O_291,N_23733,N_23793);
and UO_292 (O_292,N_23235,N_24592);
xnor UO_293 (O_293,N_23350,N_24920);
and UO_294 (O_294,N_22527,N_22558);
nor UO_295 (O_295,N_23389,N_24969);
and UO_296 (O_296,N_24711,N_24443);
nand UO_297 (O_297,N_24241,N_24092);
and UO_298 (O_298,N_24891,N_22749);
nor UO_299 (O_299,N_24858,N_24396);
nor UO_300 (O_300,N_24537,N_23709);
nand UO_301 (O_301,N_22946,N_23721);
nand UO_302 (O_302,N_23636,N_24652);
nand UO_303 (O_303,N_22893,N_22772);
xor UO_304 (O_304,N_22985,N_24171);
or UO_305 (O_305,N_23216,N_24456);
nand UO_306 (O_306,N_24379,N_22959);
nand UO_307 (O_307,N_23137,N_24975);
nor UO_308 (O_308,N_23488,N_24421);
xnor UO_309 (O_309,N_23758,N_24067);
and UO_310 (O_310,N_23986,N_24141);
and UO_311 (O_311,N_24591,N_24952);
nor UO_312 (O_312,N_23253,N_22835);
nor UO_313 (O_313,N_23120,N_23808);
nor UO_314 (O_314,N_23563,N_24472);
and UO_315 (O_315,N_23932,N_23594);
or UO_316 (O_316,N_23388,N_22706);
xor UO_317 (O_317,N_22868,N_24898);
xor UO_318 (O_318,N_22981,N_23542);
and UO_319 (O_319,N_24840,N_23812);
and UO_320 (O_320,N_24236,N_24850);
nor UO_321 (O_321,N_23226,N_23713);
nand UO_322 (O_322,N_24980,N_23521);
nand UO_323 (O_323,N_24659,N_23994);
nor UO_324 (O_324,N_24800,N_24025);
nor UO_325 (O_325,N_24069,N_24439);
or UO_326 (O_326,N_22936,N_24383);
and UO_327 (O_327,N_23078,N_22662);
xnor UO_328 (O_328,N_23049,N_23022);
nor UO_329 (O_329,N_24688,N_23832);
nand UO_330 (O_330,N_24218,N_23957);
and UO_331 (O_331,N_23051,N_24190);
nand UO_332 (O_332,N_23161,N_23802);
xnor UO_333 (O_333,N_24411,N_24763);
nand UO_334 (O_334,N_24354,N_23177);
and UO_335 (O_335,N_23337,N_23946);
and UO_336 (O_336,N_24699,N_23800);
and UO_337 (O_337,N_24057,N_24707);
and UO_338 (O_338,N_24628,N_23958);
nand UO_339 (O_339,N_22625,N_24623);
and UO_340 (O_340,N_23701,N_24908);
xor UO_341 (O_341,N_23174,N_23862);
and UO_342 (O_342,N_23208,N_23925);
nand UO_343 (O_343,N_22643,N_23365);
nand UO_344 (O_344,N_22867,N_24787);
or UO_345 (O_345,N_23990,N_23329);
xnor UO_346 (O_346,N_22755,N_22879);
or UO_347 (O_347,N_24873,N_24473);
nand UO_348 (O_348,N_22897,N_24122);
or UO_349 (O_349,N_22812,N_23149);
and UO_350 (O_350,N_24708,N_24186);
xor UO_351 (O_351,N_24220,N_24440);
xnor UO_352 (O_352,N_24412,N_23033);
and UO_353 (O_353,N_22632,N_23076);
xnor UO_354 (O_354,N_24499,N_22775);
nor UO_355 (O_355,N_23499,N_22778);
or UO_356 (O_356,N_24206,N_24085);
nand UO_357 (O_357,N_24339,N_23407);
or UO_358 (O_358,N_23390,N_23686);
xor UO_359 (O_359,N_23668,N_22710);
nor UO_360 (O_360,N_23841,N_24616);
nor UO_361 (O_361,N_22773,N_22642);
nor UO_362 (O_362,N_24730,N_24935);
nand UO_363 (O_363,N_24876,N_23302);
and UO_364 (O_364,N_24862,N_24888);
nor UO_365 (O_365,N_23444,N_24686);
nand UO_366 (O_366,N_23243,N_24676);
nand UO_367 (O_367,N_23473,N_23826);
xnor UO_368 (O_368,N_23849,N_23601);
and UO_369 (O_369,N_24036,N_23246);
and UO_370 (O_370,N_24469,N_22887);
nor UO_371 (O_371,N_24825,N_23402);
xor UO_372 (O_372,N_23128,N_23482);
and UO_373 (O_373,N_24594,N_23745);
nor UO_374 (O_374,N_23515,N_24764);
and UO_375 (O_375,N_24988,N_24718);
xor UO_376 (O_376,N_23893,N_23426);
nand UO_377 (O_377,N_22974,N_24940);
xnor UO_378 (O_378,N_23205,N_23629);
and UO_379 (O_379,N_23558,N_24814);
or UO_380 (O_380,N_23417,N_24295);
nand UO_381 (O_381,N_23291,N_24821);
nor UO_382 (O_382,N_22950,N_23209);
or UO_383 (O_383,N_22676,N_23189);
and UO_384 (O_384,N_22923,N_24859);
nand UO_385 (O_385,N_24550,N_22612);
nor UO_386 (O_386,N_22774,N_24424);
nand UO_387 (O_387,N_23508,N_22571);
xnor UO_388 (O_388,N_23616,N_24621);
nand UO_389 (O_389,N_23771,N_23115);
nor UO_390 (O_390,N_22564,N_23058);
xor UO_391 (O_391,N_24995,N_24554);
xor UO_392 (O_392,N_22860,N_24977);
xnor UO_393 (O_393,N_24004,N_23840);
nor UO_394 (O_394,N_24198,N_24088);
nand UO_395 (O_395,N_23438,N_23557);
nor UO_396 (O_396,N_22792,N_22695);
nor UO_397 (O_397,N_22725,N_24580);
nand UO_398 (O_398,N_23935,N_23664);
nor UO_399 (O_399,N_23360,N_23238);
nand UO_400 (O_400,N_24651,N_24897);
nor UO_401 (O_401,N_22771,N_22649);
xnor UO_402 (O_402,N_24168,N_22601);
nand UO_403 (O_403,N_24909,N_23153);
nand UO_404 (O_404,N_23786,N_24987);
xor UO_405 (O_405,N_24646,N_24052);
nor UO_406 (O_406,N_23839,N_22644);
and UO_407 (O_407,N_23296,N_22685);
and UO_408 (O_408,N_24314,N_23108);
or UO_409 (O_409,N_24893,N_23382);
nor UO_410 (O_410,N_23951,N_24336);
or UO_411 (O_411,N_22602,N_24349);
nor UO_412 (O_412,N_23123,N_23736);
nor UO_413 (O_413,N_22837,N_23072);
and UO_414 (O_414,N_23173,N_24832);
and UO_415 (O_415,N_22968,N_23937);
and UO_416 (O_416,N_22539,N_24625);
and UO_417 (O_417,N_24470,N_22864);
nand UO_418 (O_418,N_23278,N_23838);
and UO_419 (O_419,N_23418,N_24522);
nor UO_420 (O_420,N_24422,N_23602);
nor UO_421 (O_421,N_23107,N_24981);
nand UO_422 (O_422,N_23975,N_24511);
nand UO_423 (O_423,N_23447,N_23210);
and UO_424 (O_424,N_22648,N_24292);
nand UO_425 (O_425,N_24263,N_23591);
and UO_426 (O_426,N_23606,N_24406);
xnor UO_427 (O_427,N_23323,N_23240);
xor UO_428 (O_428,N_24720,N_22958);
xnor UO_429 (O_429,N_22637,N_24018);
xor UO_430 (O_430,N_23002,N_23393);
xnor UO_431 (O_431,N_24279,N_24794);
xor UO_432 (O_432,N_24024,N_24747);
nand UO_433 (O_433,N_22894,N_24431);
nor UO_434 (O_434,N_23853,N_24615);
and UO_435 (O_435,N_23573,N_23941);
and UO_436 (O_436,N_22591,N_23333);
xor UO_437 (O_437,N_23409,N_24613);
nor UO_438 (O_438,N_23283,N_23193);
and UO_439 (O_439,N_23950,N_22631);
nor UO_440 (O_440,N_24978,N_23441);
or UO_441 (O_441,N_22746,N_24143);
nor UO_442 (O_442,N_24784,N_24090);
and UO_443 (O_443,N_23719,N_24185);
and UO_444 (O_444,N_23113,N_24394);
nand UO_445 (O_445,N_22983,N_24463);
nor UO_446 (O_446,N_24068,N_24728);
nand UO_447 (O_447,N_24435,N_23637);
and UO_448 (O_448,N_24753,N_24817);
nor UO_449 (O_449,N_23136,N_24638);
nand UO_450 (O_450,N_24971,N_22872);
and UO_451 (O_451,N_22884,N_22530);
nand UO_452 (O_452,N_23564,N_24890);
nand UO_453 (O_453,N_24103,N_24721);
xnor UO_454 (O_454,N_23856,N_23250);
nor UO_455 (O_455,N_24990,N_24732);
xor UO_456 (O_456,N_22789,N_23556);
nor UO_457 (O_457,N_22899,N_23780);
and UO_458 (O_458,N_24223,N_24523);
nand UO_459 (O_459,N_23674,N_22599);
xor UO_460 (O_460,N_23493,N_23213);
nor UO_461 (O_461,N_23754,N_22829);
nand UO_462 (O_462,N_22554,N_24967);
nor UO_463 (O_463,N_24945,N_23851);
nand UO_464 (O_464,N_23400,N_24270);
or UO_465 (O_465,N_23728,N_22549);
and UO_466 (O_466,N_23015,N_22814);
nor UO_467 (O_467,N_24584,N_24510);
nand UO_468 (O_468,N_24536,N_23111);
xor UO_469 (O_469,N_24576,N_24413);
nand UO_470 (O_470,N_22882,N_23867);
or UO_471 (O_471,N_24268,N_22767);
nand UO_472 (O_472,N_24612,N_24879);
nand UO_473 (O_473,N_24847,N_24674);
nor UO_474 (O_474,N_22616,N_23750);
and UO_475 (O_475,N_22992,N_22847);
and UO_476 (O_476,N_23366,N_24231);
and UO_477 (O_477,N_22930,N_22891);
and UO_478 (O_478,N_24702,N_23567);
nand UO_479 (O_479,N_22853,N_24868);
xnor UO_480 (O_480,N_22573,N_24133);
nor UO_481 (O_481,N_24253,N_24207);
and UO_482 (O_482,N_24035,N_24574);
xnor UO_483 (O_483,N_23269,N_22692);
or UO_484 (O_484,N_24874,N_23903);
nor UO_485 (O_485,N_24924,N_24459);
nand UO_486 (O_486,N_22962,N_24810);
and UO_487 (O_487,N_23268,N_24583);
nand UO_488 (O_488,N_22953,N_23424);
xor UO_489 (O_489,N_23035,N_23911);
nand UO_490 (O_490,N_23275,N_23339);
and UO_491 (O_491,N_23572,N_22769);
or UO_492 (O_492,N_24948,N_24410);
nand UO_493 (O_493,N_23056,N_23949);
xnor UO_494 (O_494,N_23943,N_22973);
and UO_495 (O_495,N_22606,N_24076);
and UO_496 (O_496,N_22679,N_24163);
xnor UO_497 (O_497,N_24176,N_24001);
nand UO_498 (O_498,N_23320,N_24629);
nor UO_499 (O_499,N_23059,N_23530);
nand UO_500 (O_500,N_23175,N_24403);
xnor UO_501 (O_501,N_24356,N_22831);
nor UO_502 (O_502,N_24285,N_23141);
or UO_503 (O_503,N_23681,N_24571);
or UO_504 (O_504,N_24782,N_23346);
xnor UO_505 (O_505,N_22790,N_22809);
nor UO_506 (O_506,N_24758,N_23685);
nor UO_507 (O_507,N_24007,N_23448);
nand UO_508 (O_508,N_22905,N_23938);
xor UO_509 (O_509,N_22659,N_23936);
xor UO_510 (O_510,N_23403,N_23480);
nor UO_511 (O_511,N_24724,N_24886);
nor UO_512 (O_512,N_24880,N_23126);
xor UO_513 (O_513,N_23756,N_23901);
or UO_514 (O_514,N_23309,N_24019);
xnor UO_515 (O_515,N_22531,N_22707);
and UO_516 (O_516,N_24857,N_23273);
nor UO_517 (O_517,N_22705,N_24094);
or UO_518 (O_518,N_22816,N_24205);
nor UO_519 (O_519,N_23734,N_23890);
and UO_520 (O_520,N_23124,N_24637);
and UO_521 (O_521,N_24418,N_23391);
or UO_522 (O_522,N_24631,N_24921);
nand UO_523 (O_523,N_23559,N_22768);
nor UO_524 (O_524,N_22943,N_24836);
xnor UO_525 (O_525,N_22543,N_24689);
nand UO_526 (O_526,N_24697,N_24260);
nand UO_527 (O_527,N_23314,N_23502);
or UO_528 (O_528,N_24460,N_23584);
nand UO_529 (O_529,N_22842,N_24474);
nand UO_530 (O_530,N_24234,N_23420);
nand UO_531 (O_531,N_23544,N_22896);
xor UO_532 (O_532,N_24492,N_24925);
nand UO_533 (O_533,N_24768,N_23160);
nand UO_534 (O_534,N_22925,N_22912);
and UO_535 (O_535,N_22512,N_23703);
and UO_536 (O_536,N_23012,N_24578);
xnor UO_537 (O_537,N_22575,N_24404);
or UO_538 (O_538,N_23286,N_23920);
nor UO_539 (O_539,N_23509,N_23966);
xnor UO_540 (O_540,N_23697,N_22802);
nor UO_541 (O_541,N_22592,N_24063);
or UO_542 (O_542,N_23359,N_24130);
nor UO_543 (O_543,N_23510,N_22552);
or UO_544 (O_544,N_23690,N_23921);
xnor UO_545 (O_545,N_24776,N_24968);
nand UO_546 (O_546,N_23267,N_22797);
and UO_547 (O_547,N_22966,N_24432);
and UO_548 (O_548,N_24949,N_23334);
and UO_549 (O_549,N_24037,N_24346);
or UO_550 (O_550,N_23338,N_24885);
xor UO_551 (O_551,N_23999,N_24287);
nand UO_552 (O_552,N_22561,N_24486);
nand UO_553 (O_553,N_23536,N_22876);
and UO_554 (O_554,N_23293,N_23706);
nor UO_555 (O_555,N_23539,N_22555);
nor UO_556 (O_556,N_23723,N_23399);
and UO_557 (O_557,N_23579,N_23540);
nand UO_558 (O_558,N_23976,N_24375);
nor UO_559 (O_559,N_24773,N_22750);
nand UO_560 (O_560,N_23206,N_23406);
nor UO_561 (O_561,N_23592,N_23687);
and UO_562 (O_562,N_24144,N_24722);
or UO_563 (O_563,N_23298,N_23612);
and UO_564 (O_564,N_23822,N_24627);
and UO_565 (O_565,N_24061,N_23410);
xnor UO_566 (O_566,N_24172,N_22731);
nor UO_567 (O_567,N_22582,N_23837);
nor UO_568 (O_568,N_22880,N_23797);
xor UO_569 (O_569,N_22529,N_23188);
or UO_570 (O_570,N_23825,N_24767);
nand UO_571 (O_571,N_24022,N_24113);
nand UO_572 (O_572,N_24153,N_23645);
or UO_573 (O_573,N_22955,N_23702);
and UO_574 (O_574,N_23451,N_24901);
nor UO_575 (O_575,N_23514,N_24179);
nand UO_576 (O_576,N_23725,N_23769);
xor UO_577 (O_577,N_24177,N_23484);
or UO_578 (O_578,N_23740,N_22658);
xnor UO_579 (O_579,N_24164,N_23942);
and UO_580 (O_580,N_23823,N_24108);
xnor UO_581 (O_581,N_22687,N_23930);
xnor UO_582 (O_582,N_24078,N_23850);
nand UO_583 (O_583,N_22518,N_24696);
or UO_584 (O_584,N_24495,N_23127);
and UO_585 (O_585,N_23491,N_24604);
xnor UO_586 (O_586,N_23277,N_22675);
xor UO_587 (O_587,N_23971,N_23376);
nor UO_588 (O_588,N_22794,N_23795);
and UO_589 (O_589,N_24831,N_23730);
or UO_590 (O_590,N_22559,N_23122);
xnor UO_591 (O_591,N_22617,N_23165);
and UO_592 (O_592,N_23859,N_23714);
or UO_593 (O_593,N_23112,N_23460);
and UO_594 (O_594,N_23279,N_22906);
nand UO_595 (O_595,N_24337,N_23894);
and UO_596 (O_596,N_24582,N_23010);
and UO_597 (O_597,N_23094,N_22841);
or UO_598 (O_598,N_23241,N_22883);
nor UO_599 (O_599,N_24429,N_24355);
xnor UO_600 (O_600,N_23915,N_22988);
or UO_601 (O_601,N_23219,N_22997);
nor UO_602 (O_602,N_22971,N_24517);
nand UO_603 (O_603,N_22927,N_22533);
and UO_604 (O_604,N_24116,N_24081);
nand UO_605 (O_605,N_23414,N_22961);
and UO_606 (O_606,N_23526,N_24366);
and UO_607 (O_607,N_23179,N_24544);
xnor UO_608 (O_608,N_22604,N_24479);
or UO_609 (O_609,N_23315,N_23228);
nor UO_610 (O_610,N_24291,N_23737);
or UO_611 (O_611,N_23025,N_23048);
nand UO_612 (O_612,N_24798,N_22895);
and UO_613 (O_613,N_23030,N_23457);
nor UO_614 (O_614,N_23089,N_23064);
and UO_615 (O_615,N_24918,N_24944);
nor UO_616 (O_616,N_22764,N_24793);
xor UO_617 (O_617,N_23341,N_24327);
nor UO_618 (O_618,N_22624,N_24643);
nand UO_619 (O_619,N_24710,N_24507);
nand UO_620 (O_620,N_22863,N_23421);
or UO_621 (O_621,N_23374,N_24259);
nand UO_622 (O_622,N_23281,N_23532);
nor UO_623 (O_623,N_24219,N_22724);
and UO_624 (O_624,N_24974,N_24526);
xor UO_625 (O_625,N_24419,N_22541);
and UO_626 (O_626,N_23694,N_24515);
or UO_627 (O_627,N_24261,N_22783);
xor UO_628 (O_628,N_24098,N_24501);
xnor UO_629 (O_629,N_22656,N_23470);
nor UO_630 (O_630,N_23836,N_22628);
nand UO_631 (O_631,N_23259,N_24157);
or UO_632 (O_632,N_23500,N_23118);
or UO_633 (O_633,N_22603,N_24042);
or UO_634 (O_634,N_23185,N_23537);
or UO_635 (O_635,N_23044,N_24895);
and UO_636 (O_636,N_24669,N_22874);
nor UO_637 (O_637,N_23760,N_23081);
nand UO_638 (O_638,N_23827,N_23207);
and UO_639 (O_639,N_24622,N_24717);
nor UO_640 (O_640,N_24397,N_23474);
xor UO_641 (O_641,N_22726,N_22557);
and UO_642 (O_642,N_23968,N_23801);
and UO_643 (O_643,N_23084,N_22979);
nand UO_644 (O_644,N_24573,N_22579);
and UO_645 (O_645,N_23882,N_24387);
or UO_646 (O_646,N_23732,N_22941);
and UO_647 (O_647,N_23342,N_24195);
and UO_648 (O_648,N_23785,N_24712);
nor UO_649 (O_649,N_23245,N_24199);
or UO_650 (O_650,N_24213,N_24772);
and UO_651 (O_651,N_22671,N_22700);
nand UO_652 (O_652,N_23396,N_22540);
and UO_653 (O_653,N_22660,N_23231);
nor UO_654 (O_654,N_24225,N_22654);
or UO_655 (O_655,N_22875,N_22978);
nor UO_656 (O_656,N_24950,N_24264);
or UO_657 (O_657,N_24726,N_23373);
and UO_658 (O_658,N_23419,N_23715);
nand UO_659 (O_659,N_23658,N_24280);
and UO_660 (O_660,N_22852,N_22694);
and UO_661 (O_661,N_24482,N_23203);
or UO_662 (O_662,N_23164,N_23900);
xor UO_663 (O_663,N_23489,N_24769);
nand UO_664 (O_664,N_24790,N_23166);
nand UO_665 (O_665,N_24943,N_24527);
nand UO_666 (O_666,N_24508,N_23782);
or UO_667 (O_667,N_24700,N_23872);
or UO_668 (O_668,N_23110,N_24487);
nor UO_669 (O_669,N_22916,N_24680);
and UO_670 (O_670,N_24750,N_22866);
xor UO_671 (O_671,N_23271,N_23998);
nor UO_672 (O_672,N_23747,N_23363);
nand UO_673 (O_673,N_22948,N_24020);
nand UO_674 (O_674,N_22917,N_22699);
nor UO_675 (O_675,N_22566,N_24900);
and UO_676 (O_676,N_24493,N_23906);
nand UO_677 (O_677,N_23001,N_24512);
nand UO_678 (O_678,N_22753,N_24809);
or UO_679 (O_679,N_24566,N_24834);
nand UO_680 (O_680,N_22510,N_24912);
xor UO_681 (O_681,N_23163,N_23566);
nor UO_682 (O_682,N_24986,N_24075);
nand UO_683 (O_683,N_22739,N_23805);
or UO_684 (O_684,N_22901,N_22975);
nand UO_685 (O_685,N_24352,N_22900);
or UO_686 (O_686,N_24852,N_23610);
and UO_687 (O_687,N_22516,N_24425);
nand UO_688 (O_688,N_24064,N_24520);
or UO_689 (O_689,N_24731,N_24324);
and UO_690 (O_690,N_23244,N_23644);
or UO_691 (O_691,N_24058,N_22677);
nor UO_692 (O_692,N_24682,N_24601);
or UO_693 (O_693,N_23464,N_22766);
and UO_694 (O_694,N_23683,N_22910);
xnor UO_695 (O_695,N_22562,N_24315);
xnor UO_696 (O_696,N_24632,N_23100);
and UO_697 (O_697,N_24704,N_23139);
nor UO_698 (O_698,N_23595,N_24690);
xnor UO_699 (O_699,N_23416,N_22701);
or UO_700 (O_700,N_23613,N_23158);
xnor UO_701 (O_701,N_24533,N_24008);
xnor UO_702 (O_702,N_24082,N_23562);
or UO_703 (O_703,N_24192,N_24232);
nor UO_704 (O_704,N_23251,N_24255);
or UO_705 (O_705,N_22546,N_22704);
or UO_706 (O_706,N_24468,N_24808);
and UO_707 (O_707,N_22934,N_23326);
and UO_708 (O_708,N_23313,N_24239);
xnor UO_709 (O_709,N_23997,N_22849);
or UO_710 (O_710,N_24984,N_23551);
and UO_711 (O_711,N_23307,N_23744);
nor UO_712 (O_712,N_24864,N_23134);
nor UO_713 (O_713,N_23549,N_23868);
xnor UO_714 (O_714,N_24602,N_23913);
or UO_715 (O_715,N_22673,N_23898);
or UO_716 (O_716,N_24838,N_24587);
nand UO_717 (O_717,N_23370,N_23934);
and UO_718 (O_718,N_24189,N_24903);
nor UO_719 (O_719,N_22503,N_23940);
xor UO_720 (O_720,N_24010,N_23883);
xor UO_721 (O_721,N_23615,N_24513);
and UO_722 (O_722,N_23538,N_23252);
or UO_723 (O_723,N_23731,N_23886);
and UO_724 (O_724,N_22888,N_23729);
and UO_725 (O_725,N_23345,N_24370);
and UO_726 (O_726,N_24444,N_24668);
or UO_727 (O_727,N_23858,N_22640);
or UO_728 (O_728,N_24274,N_24134);
nand UO_729 (O_729,N_22785,N_23654);
nand UO_730 (O_730,N_24451,N_23254);
or UO_731 (O_731,N_24409,N_23380);
and UO_732 (O_732,N_24284,N_22821);
nor UO_733 (O_733,N_24521,N_23586);
nor UO_734 (O_734,N_23779,N_24781);
nor UO_735 (O_735,N_24367,N_23172);
nor UO_736 (O_736,N_24617,N_24338);
nor UO_737 (O_737,N_23517,N_23099);
nand UO_738 (O_738,N_24670,N_24777);
nand UO_739 (O_739,N_23608,N_24106);
xor UO_740 (O_740,N_23117,N_24677);
or UO_741 (O_741,N_23979,N_23472);
nand UO_742 (O_742,N_23019,N_24365);
and UO_743 (O_743,N_23796,N_22840);
and UO_744 (O_744,N_22583,N_23553);
and UO_745 (O_745,N_23568,N_24031);
and UO_746 (O_746,N_22686,N_23230);
and UO_747 (O_747,N_24673,N_23712);
or UO_748 (O_748,N_22742,N_24516);
nor UO_749 (O_749,N_22815,N_23768);
nor UO_750 (O_750,N_22878,N_24826);
or UO_751 (O_751,N_24854,N_23989);
and UO_752 (O_752,N_24563,N_24266);
or UO_753 (O_753,N_24048,N_22697);
nor UO_754 (O_754,N_24514,N_24807);
nor UO_755 (O_755,N_24226,N_23757);
nand UO_756 (O_756,N_24542,N_24091);
and UO_757 (O_757,N_24332,N_22751);
nand UO_758 (O_758,N_24994,N_24620);
xor UO_759 (O_759,N_23287,N_24654);
or UO_760 (O_760,N_23215,N_24348);
nor UO_761 (O_761,N_24417,N_24655);
or UO_762 (O_762,N_24446,N_24727);
and UO_763 (O_763,N_22990,N_24283);
or UO_764 (O_764,N_23021,N_24217);
xor UO_765 (O_765,N_22928,N_23977);
or UO_766 (O_766,N_24691,N_23847);
xor UO_767 (O_767,N_24079,N_24471);
nor UO_768 (O_768,N_22889,N_23280);
nand UO_769 (O_769,N_24941,N_24350);
nor UO_770 (O_770,N_23459,N_24884);
or UO_771 (O_771,N_23835,N_23748);
nand UO_772 (O_772,N_24741,N_23598);
or UO_773 (O_773,N_24095,N_24927);
nand UO_774 (O_774,N_23905,N_22728);
xnor UO_775 (O_775,N_23300,N_24099);
nand UO_776 (O_776,N_24806,N_24959);
or UO_777 (O_777,N_23580,N_23804);
nand UO_778 (O_778,N_24308,N_23197);
xor UO_779 (O_779,N_23427,N_24430);
nand UO_780 (O_780,N_24634,N_23582);
xnor UO_781 (O_781,N_22913,N_24257);
or UO_782 (O_782,N_22996,N_24307);
nor UO_783 (O_783,N_23097,N_24118);
and UO_784 (O_784,N_24374,N_23860);
xor UO_785 (O_785,N_22611,N_24525);
nand UO_786 (O_786,N_23140,N_24973);
xor UO_787 (O_787,N_22521,N_24535);
or UO_788 (O_788,N_24252,N_22909);
or UO_789 (O_789,N_23285,N_23053);
or UO_790 (O_790,N_24498,N_24294);
xor UO_791 (O_791,N_22784,N_22886);
and UO_792 (O_792,N_23055,N_23969);
xnor UO_793 (O_793,N_24589,N_22956);
nand UO_794 (O_794,N_23311,N_24415);
nand UO_795 (O_795,N_24737,N_24715);
nand UO_796 (O_796,N_24733,N_24752);
or UO_797 (O_797,N_23434,N_24965);
nor UO_798 (O_798,N_24433,N_23741);
nand UO_799 (O_799,N_24249,N_23781);
and UO_800 (O_800,N_23159,N_23217);
or UO_801 (O_801,N_22691,N_24687);
xor UO_802 (O_802,N_23116,N_23344);
xnor UO_803 (O_803,N_24071,N_23431);
nor UO_804 (O_804,N_23617,N_24276);
or UO_805 (O_805,N_23308,N_23132);
or UO_806 (O_806,N_24694,N_23330);
xnor UO_807 (O_807,N_23357,N_23381);
or UO_808 (O_808,N_23959,N_22580);
xnor UO_809 (O_809,N_22629,N_23525);
nand UO_810 (O_810,N_24894,N_23753);
nand UO_811 (O_811,N_23609,N_23670);
nand UO_812 (O_812,N_23257,N_22653);
xnor UO_813 (O_813,N_24765,N_22667);
or UO_814 (O_814,N_24013,N_22661);
xnor UO_815 (O_815,N_23260,N_22922);
nand UO_816 (O_816,N_23531,N_23501);
nor UO_817 (O_817,N_22709,N_23294);
nand UO_818 (O_818,N_23486,N_22877);
xnor UO_819 (O_819,N_24853,N_24441);
nand UO_820 (O_820,N_22587,N_24539);
or UO_821 (O_821,N_24695,N_22758);
or UO_822 (O_822,N_24488,N_24070);
nand UO_823 (O_823,N_22586,N_23306);
xnor UO_824 (O_824,N_23180,N_22657);
and UO_825 (O_825,N_23724,N_24917);
nand UO_826 (O_826,N_23045,N_24457);
and UO_827 (O_827,N_24115,N_23806);
nand UO_828 (O_828,N_24320,N_22581);
nor UO_829 (O_829,N_24626,N_24309);
xnor UO_830 (O_830,N_22759,N_23479);
and UO_831 (O_831,N_24869,N_24391);
or UO_832 (O_832,N_23863,N_23987);
nand UO_833 (O_833,N_23069,N_24505);
or UO_834 (O_834,N_23080,N_24494);
or UO_835 (O_835,N_24739,N_24014);
nand UO_836 (O_836,N_22668,N_23899);
xor UO_837 (O_837,N_24951,N_24407);
and UO_838 (O_838,N_23752,N_24792);
and UO_839 (O_839,N_24771,N_24196);
and UO_840 (O_840,N_22781,N_22635);
and UO_841 (O_841,N_23909,N_24066);
nand UO_842 (O_842,N_22678,N_22881);
nand UO_843 (O_843,N_24683,N_24117);
nor UO_844 (O_844,N_23788,N_24401);
xor UO_845 (O_845,N_23810,N_22824);
nand UO_846 (O_846,N_24165,N_23916);
or UO_847 (O_847,N_23082,N_23927);
nor UO_848 (O_848,N_24111,N_23961);
or UO_849 (O_849,N_24275,N_24530);
or UO_850 (O_850,N_24540,N_23202);
nor UO_851 (O_851,N_23887,N_24000);
nand UO_852 (O_852,N_23776,N_24614);
xor UO_853 (O_853,N_23454,N_23816);
xnor UO_854 (O_854,N_22547,N_23211);
and UO_855 (O_855,N_23008,N_24046);
nand UO_856 (O_856,N_22723,N_23371);
xnor UO_857 (O_857,N_23027,N_24962);
and UO_858 (O_858,N_23621,N_22597);
xnor UO_859 (O_859,N_22870,N_23708);
nor UO_860 (O_860,N_24645,N_24322);
or UO_861 (O_861,N_23848,N_24788);
nor UO_862 (O_862,N_24851,N_24600);
nor UO_863 (O_863,N_24725,N_24371);
xnor UO_864 (O_864,N_22519,N_24248);
and UO_865 (O_865,N_22576,N_22862);
nor UO_866 (O_866,N_24021,N_22920);
xor UO_867 (O_867,N_22669,N_23282);
and UO_868 (O_868,N_24222,N_24685);
and UO_869 (O_869,N_24112,N_22904);
nand UO_870 (O_870,N_23169,N_23970);
xnor UO_871 (O_871,N_24751,N_24693);
or UO_872 (O_872,N_23761,N_23603);
nand UO_873 (O_873,N_24477,N_23960);
nor UO_874 (O_874,N_24579,N_22652);
nor UO_875 (O_875,N_23440,N_23871);
nand UO_876 (O_876,N_24823,N_23485);
or UO_877 (O_877,N_23820,N_23014);
and UO_878 (O_878,N_24230,N_24892);
nor UO_879 (O_879,N_24827,N_24841);
or UO_880 (O_880,N_24465,N_24829);
or UO_881 (O_881,N_23009,N_24384);
xor UO_882 (O_882,N_23042,N_24402);
nor UO_883 (O_883,N_23385,N_23057);
xnor UO_884 (O_884,N_22647,N_22940);
xnor UO_885 (O_885,N_22526,N_23145);
or UO_886 (O_886,N_22623,N_24489);
nor UO_887 (O_887,N_24246,N_24845);
or UO_888 (O_888,N_23495,N_23524);
nor UO_889 (O_889,N_22908,N_23335);
or UO_890 (O_890,N_23981,N_23325);
xnor UO_891 (O_891,N_23204,N_23655);
or UO_892 (O_892,N_24200,N_24930);
nand UO_893 (O_893,N_24047,N_24590);
nand UO_894 (O_894,N_23604,N_24002);
or UO_895 (O_895,N_23477,N_24096);
nand UO_896 (O_896,N_23513,N_23954);
nor UO_897 (O_897,N_23264,N_23955);
nand UO_898 (O_898,N_23896,N_24902);
nand UO_899 (O_899,N_23988,N_24766);
xnor UO_900 (O_900,N_22954,N_24541);
xnor UO_901 (O_901,N_23888,N_22796);
xnor UO_902 (O_902,N_23548,N_23352);
or UO_903 (O_903,N_22822,N_24714);
xnor UO_904 (O_904,N_23547,N_24946);
xor UO_905 (O_905,N_22550,N_23095);
nand UO_906 (O_906,N_23917,N_23266);
xnor UO_907 (O_907,N_24954,N_24449);
or UO_908 (O_908,N_24789,N_23364);
and UO_909 (O_909,N_23727,N_23814);
nor UO_910 (O_910,N_23194,N_22929);
xnor UO_911 (O_911,N_24928,N_23088);
nand UO_912 (O_912,N_22960,N_24761);
or UO_913 (O_913,N_24166,N_22813);
xnor UO_914 (O_914,N_24484,N_23947);
xor UO_915 (O_915,N_22565,N_24870);
xnor UO_916 (O_916,N_24875,N_22734);
and UO_917 (O_917,N_22508,N_23005);
and UO_918 (O_918,N_24455,N_23554);
nor UO_919 (O_919,N_23050,N_24509);
and UO_920 (O_920,N_24662,N_22722);
or UO_921 (O_921,N_23630,N_23224);
nand UO_922 (O_922,N_23696,N_24229);
or UO_923 (O_923,N_23041,N_22556);
and UO_924 (O_924,N_23429,N_23392);
and UO_925 (O_925,N_24904,N_23340);
and UO_926 (O_926,N_23458,N_24428);
or UO_927 (O_927,N_23361,N_24746);
or UO_928 (O_928,N_23789,N_22651);
nand UO_929 (O_929,N_23751,N_22803);
or UO_930 (O_930,N_24672,N_24703);
nand UO_931 (O_931,N_22538,N_24547);
nor UO_932 (O_932,N_23433,N_24097);
nand UO_933 (O_933,N_22633,N_24830);
or UO_934 (O_934,N_24639,N_24605);
and UO_935 (O_935,N_24104,N_23036);
nand UO_936 (O_936,N_24779,N_24644);
or UO_937 (O_937,N_23923,N_23641);
xor UO_938 (O_938,N_24445,N_24983);
or UO_939 (O_939,N_24706,N_24243);
nand UO_940 (O_940,N_24372,N_23063);
xor UO_941 (O_941,N_23046,N_22646);
xnor UO_942 (O_942,N_23028,N_23649);
xnor UO_943 (O_943,N_22799,N_23412);
xor UO_944 (O_944,N_23794,N_24497);
nand UO_945 (O_945,N_22818,N_23738);
nor UO_946 (O_946,N_22708,N_22665);
nand UO_947 (O_947,N_23815,N_22711);
or UO_948 (O_948,N_24734,N_23889);
xnor UO_949 (O_949,N_23995,N_22570);
and UO_950 (O_950,N_22614,N_24221);
nor UO_951 (O_951,N_24956,N_24197);
xor UO_952 (O_952,N_22744,N_23310);
or UO_953 (O_953,N_22590,N_23247);
nor UO_954 (O_954,N_24363,N_22952);
or UO_955 (O_955,N_22931,N_24029);
nand UO_956 (O_956,N_23263,N_23854);
xnor UO_957 (O_957,N_24502,N_23552);
xnor UO_958 (O_958,N_24833,N_22850);
nand UO_959 (O_959,N_23090,N_23798);
or UO_960 (O_960,N_24558,N_23368);
or UO_961 (O_961,N_23222,N_22963);
nor UO_962 (O_962,N_24531,N_22524);
nor UO_963 (O_963,N_23071,N_23073);
and UO_964 (O_964,N_23852,N_22832);
xor UO_965 (O_965,N_24245,N_22833);
xor UO_966 (O_966,N_23218,N_23541);
xor UO_967 (O_967,N_24414,N_24390);
xnor UO_968 (O_968,N_23628,N_24663);
and UO_969 (O_969,N_24026,N_22859);
nor UO_970 (O_970,N_22504,N_23597);
nand UO_971 (O_971,N_23109,N_24077);
or UO_972 (O_972,N_23944,N_22747);
or UO_973 (O_973,N_23765,N_23054);
or UO_974 (O_974,N_22548,N_23212);
nor UO_975 (O_975,N_24201,N_23755);
nand UO_976 (O_976,N_23575,N_23083);
xor UO_977 (O_977,N_24132,N_23931);
or UO_978 (O_978,N_23710,N_22738);
nor UO_979 (O_979,N_23699,N_24636);
xor UO_980 (O_980,N_22693,N_24416);
nand UO_981 (O_981,N_24543,N_22745);
xnor UO_982 (O_982,N_23331,N_24127);
nand UO_983 (O_983,N_22532,N_22820);
xor UO_984 (O_984,N_22810,N_23237);
xor UO_985 (O_985,N_23985,N_22609);
nand UO_986 (O_986,N_22984,N_24161);
nand UO_987 (O_987,N_23605,N_24423);
nand UO_988 (O_988,N_23187,N_24128);
and UO_989 (O_989,N_24466,N_23632);
or UO_990 (O_990,N_22801,N_24126);
xor UO_991 (O_991,N_24926,N_23375);
nand UO_992 (O_992,N_23199,N_23587);
or UO_993 (O_993,N_24861,N_24570);
nand UO_994 (O_994,N_22535,N_23698);
nand UO_995 (O_995,N_23830,N_24878);
nor UO_996 (O_996,N_24976,N_24546);
and UO_997 (O_997,N_23467,N_22608);
nor UO_998 (O_998,N_24123,N_23152);
and UO_999 (O_999,N_23953,N_24989);
nand UO_1000 (O_1000,N_24160,N_22871);
and UO_1001 (O_1001,N_23809,N_23475);
and UO_1002 (O_1002,N_24483,N_24140);
nand UO_1003 (O_1003,N_23274,N_24641);
xor UO_1004 (O_1004,N_23663,N_24150);
and UO_1005 (O_1005,N_24551,N_23182);
or UO_1006 (O_1006,N_22544,N_22732);
nand UO_1007 (O_1007,N_24500,N_24849);
and UO_1008 (O_1008,N_23679,N_24114);
nand UO_1009 (O_1009,N_23912,N_22932);
nor UO_1010 (O_1010,N_22736,N_23505);
nor UO_1011 (O_1011,N_23395,N_24450);
nand UO_1012 (O_1012,N_24698,N_24942);
nand UO_1013 (O_1013,N_24050,N_24215);
nor UO_1014 (O_1014,N_24297,N_22838);
nor UO_1015 (O_1015,N_24748,N_24797);
nand UO_1016 (O_1016,N_24889,N_23588);
or UO_1017 (O_1017,N_23824,N_22977);
nand UO_1018 (O_1018,N_24167,N_24012);
or UO_1019 (O_1019,N_24738,N_23565);
xor UO_1020 (O_1020,N_22729,N_23817);
or UO_1021 (O_1021,N_23317,N_22970);
nand UO_1022 (O_1022,N_22811,N_23759);
xnor UO_1023 (O_1023,N_24812,N_24555);
xnor UO_1024 (O_1024,N_23627,N_24389);
nand UO_1025 (O_1025,N_23659,N_23869);
nand UO_1026 (O_1026,N_24073,N_23618);
xnor UO_1027 (O_1027,N_24609,N_23623);
nand UO_1028 (O_1028,N_22740,N_22844);
nand UO_1029 (O_1029,N_24262,N_24214);
nor UO_1030 (O_1030,N_22569,N_24183);
nand UO_1031 (O_1031,N_22856,N_24863);
or UO_1032 (O_1032,N_23673,N_23692);
and UO_1033 (O_1033,N_24119,N_24298);
nor UO_1034 (O_1034,N_23020,N_24145);
nand UO_1035 (O_1035,N_24341,N_24359);
nand UO_1036 (O_1036,N_24335,N_24881);
or UO_1037 (O_1037,N_22595,N_23875);
nand UO_1038 (O_1038,N_22937,N_24105);
nor UO_1039 (O_1039,N_24865,N_23818);
nor UO_1040 (O_1040,N_23018,N_24791);
nor UO_1041 (O_1041,N_23665,N_23086);
and UO_1042 (O_1042,N_23622,N_23272);
xor UO_1043 (O_1043,N_23114,N_24039);
nand UO_1044 (O_1044,N_22965,N_24553);
or UO_1045 (O_1045,N_23919,N_24745);
nor UO_1046 (O_1046,N_24299,N_23819);
nor UO_1047 (O_1047,N_24534,N_23131);
nand UO_1048 (O_1048,N_22944,N_22826);
nand UO_1049 (O_1049,N_24774,N_23017);
xor UO_1050 (O_1050,N_23029,N_24649);
nor UO_1051 (O_1051,N_22808,N_23354);
nor UO_1052 (O_1052,N_23964,N_24267);
or UO_1053 (O_1053,N_24964,N_23590);
and UO_1054 (O_1054,N_23777,N_24304);
or UO_1055 (O_1055,N_23261,N_22627);
nand UO_1056 (O_1056,N_24321,N_22613);
or UO_1057 (O_1057,N_23520,N_24919);
and UO_1058 (O_1058,N_24202,N_22682);
or UO_1059 (O_1059,N_23533,N_23233);
nand UO_1060 (O_1060,N_23873,N_23550);
nand UO_1061 (O_1061,N_22528,N_23265);
xnor UO_1062 (O_1062,N_23792,N_23401);
or UO_1063 (O_1063,N_24661,N_24855);
xnor UO_1064 (O_1064,N_24860,N_23527);
nor UO_1065 (O_1065,N_23635,N_24301);
nand UO_1066 (O_1066,N_22754,N_22596);
or UO_1067 (O_1067,N_24828,N_24125);
or UO_1068 (O_1068,N_24658,N_22982);
xnor UO_1069 (O_1069,N_24856,N_23430);
nor UO_1070 (O_1070,N_24565,N_23192);
or UO_1071 (O_1071,N_24056,N_24953);
xor UO_1072 (O_1072,N_24173,N_23619);
and UO_1073 (O_1073,N_24598,N_22924);
and UO_1074 (O_1074,N_23631,N_24344);
nand UO_1075 (O_1075,N_23620,N_24438);
xnor UO_1076 (O_1076,N_23312,N_23060);
and UO_1077 (O_1077,N_23611,N_23383);
nand UO_1078 (O_1078,N_24334,N_23876);
xnor UO_1079 (O_1079,N_24740,N_23497);
nand UO_1080 (O_1080,N_23874,N_24110);
xnor UO_1081 (O_1081,N_23483,N_24966);
or UO_1082 (O_1082,N_24842,N_22714);
and UO_1083 (O_1083,N_23091,N_22674);
xor UO_1084 (O_1084,N_24705,N_24452);
nand UO_1085 (O_1085,N_24813,N_23626);
nand UO_1086 (O_1086,N_23037,N_24083);
nand UO_1087 (O_1087,N_23232,N_23907);
or UO_1088 (O_1088,N_24072,N_23939);
nand UO_1089 (O_1089,N_23991,N_24839);
and UO_1090 (O_1090,N_24837,N_23154);
and UO_1091 (O_1091,N_24212,N_23902);
or UO_1092 (O_1092,N_23787,N_24915);
or UO_1093 (O_1093,N_23449,N_23555);
xor UO_1094 (O_1094,N_23578,N_22787);
or UO_1095 (O_1095,N_23092,N_24250);
or UO_1096 (O_1096,N_24398,N_23918);
or UO_1097 (O_1097,N_22865,N_23593);
and UO_1098 (O_1098,N_23743,N_23534);
nand UO_1099 (O_1099,N_23358,N_24361);
and UO_1100 (O_1100,N_23143,N_22577);
nor UO_1101 (O_1101,N_22534,N_23075);
or UO_1102 (O_1102,N_23778,N_23181);
nor UO_1103 (O_1103,N_23791,N_24329);
xor UO_1104 (O_1104,N_22505,N_23963);
nor UO_1105 (O_1105,N_24360,N_24939);
and UO_1106 (O_1106,N_22553,N_23647);
xor UO_1107 (O_1107,N_22846,N_24453);
and UO_1108 (O_1108,N_24529,N_23016);
xor UO_1109 (O_1109,N_24552,N_22735);
nor UO_1110 (O_1110,N_24242,N_23362);
and UO_1111 (O_1111,N_23378,N_22619);
or UO_1112 (O_1112,N_24684,N_24100);
xnor UO_1113 (O_1113,N_24678,N_24866);
nor UO_1114 (O_1114,N_23372,N_22762);
xnor UO_1115 (O_1115,N_24313,N_22500);
xor UO_1116 (O_1116,N_24933,N_23643);
nand UO_1117 (O_1117,N_23026,N_24936);
or UO_1118 (O_1118,N_22618,N_24844);
xor UO_1119 (O_1119,N_23996,N_24743);
nand UO_1120 (O_1120,N_24170,N_22779);
nand UO_1121 (O_1121,N_24139,N_24162);
nand UO_1122 (O_1122,N_22902,N_23220);
nor UO_1123 (O_1123,N_22945,N_23062);
nor UO_1124 (O_1124,N_22933,N_24244);
or UO_1125 (O_1125,N_24386,N_23377);
nor UO_1126 (O_1126,N_24323,N_22827);
or UO_1127 (O_1127,N_23633,N_23047);
xor UO_1128 (O_1128,N_24074,N_23167);
nor UO_1129 (O_1129,N_23157,N_22718);
and UO_1130 (O_1130,N_24564,N_22921);
nand UO_1131 (O_1131,N_23739,N_24491);
or UO_1132 (O_1132,N_24330,N_24362);
xor UO_1133 (O_1133,N_23452,N_24187);
and UO_1134 (O_1134,N_23967,N_22502);
and UO_1135 (O_1135,N_24635,N_22926);
or UO_1136 (O_1136,N_23455,N_24381);
nor UO_1137 (O_1137,N_24258,N_22942);
nor UO_1138 (O_1138,N_23332,N_22641);
or UO_1139 (O_1139,N_22666,N_24368);
xor UO_1140 (O_1140,N_24671,N_24210);
or UO_1141 (O_1141,N_23897,N_23437);
or UO_1142 (O_1142,N_24269,N_24434);
nand UO_1143 (O_1143,N_24420,N_23535);
nand UO_1144 (O_1144,N_22907,N_24033);
xnor UO_1145 (O_1145,N_24093,N_24089);
nand UO_1146 (O_1146,N_23150,N_22752);
nand UO_1147 (O_1147,N_24121,N_24393);
nor UO_1148 (O_1148,N_24556,N_24174);
xor UO_1149 (O_1149,N_23770,N_23367);
xor UO_1150 (O_1150,N_22703,N_24929);
and UO_1151 (O_1151,N_22684,N_23004);
and UO_1152 (O_1152,N_24138,N_22861);
xnor UO_1153 (O_1153,N_24216,N_22574);
or UO_1154 (O_1154,N_22737,N_22804);
xor UO_1155 (O_1155,N_23878,N_22845);
nand UO_1156 (O_1156,N_24288,N_22568);
nand UO_1157 (O_1157,N_24041,N_22918);
xor UO_1158 (O_1158,N_24729,N_24159);
and UO_1159 (O_1159,N_23933,N_22892);
or UO_1160 (O_1160,N_23336,N_23105);
nor UO_1161 (O_1161,N_22843,N_24148);
nand UO_1162 (O_1162,N_22585,N_23884);
or UO_1163 (O_1163,N_22522,N_23891);
nand UO_1164 (O_1164,N_22817,N_23292);
nand UO_1165 (O_1165,N_24822,N_23924);
nand UO_1166 (O_1166,N_22645,N_23106);
nand UO_1167 (O_1167,N_23270,N_23546);
or UO_1168 (O_1168,N_23349,N_24053);
nor UO_1169 (O_1169,N_23249,N_22650);
xnor UO_1170 (O_1170,N_23178,N_24281);
nor UO_1171 (O_1171,N_24211,N_23965);
nand UO_1172 (O_1172,N_23634,N_23749);
and UO_1173 (O_1173,N_23571,N_23885);
nand UO_1174 (O_1174,N_22560,N_23003);
nor UO_1175 (O_1175,N_22588,N_24282);
nand UO_1176 (O_1176,N_23319,N_23135);
and UO_1177 (O_1177,N_24824,N_24633);
and UO_1178 (O_1178,N_23413,N_24559);
and UO_1179 (O_1179,N_22537,N_22760);
xor UO_1180 (O_1180,N_22761,N_23487);
nand UO_1181 (O_1181,N_23720,N_24271);
nand UO_1182 (O_1182,N_22507,N_23807);
nand UO_1183 (O_1183,N_23031,N_23945);
nor UO_1184 (O_1184,N_23239,N_23462);
or UO_1185 (O_1185,N_23523,N_23512);
xnor UO_1186 (O_1186,N_24462,N_22713);
and UO_1187 (O_1187,N_23982,N_23006);
nand UO_1188 (O_1188,N_22757,N_22698);
nor UO_1189 (O_1189,N_23397,N_23691);
nand UO_1190 (O_1190,N_23675,N_23992);
nor UO_1191 (O_1191,N_24369,N_22689);
or UO_1192 (O_1192,N_24447,N_23011);
nand UO_1193 (O_1193,N_23465,N_23522);
nor UO_1194 (O_1194,N_22947,N_23516);
or UO_1195 (O_1195,N_23087,N_24191);
or UO_1196 (O_1196,N_24467,N_23763);
and UO_1197 (O_1197,N_23102,N_24656);
or UO_1198 (O_1198,N_23834,N_22800);
xnor UO_1199 (O_1199,N_22600,N_23705);
nor UO_1200 (O_1200,N_22980,N_24310);
xor UO_1201 (O_1201,N_24783,N_22780);
nor UO_1202 (O_1202,N_22681,N_24692);
and UO_1203 (O_1203,N_23973,N_22598);
xnor UO_1204 (O_1204,N_23067,N_23656);
xnor UO_1205 (O_1205,N_24300,N_23000);
xor UO_1206 (O_1206,N_23079,N_22839);
or UO_1207 (O_1207,N_22855,N_23471);
and UO_1208 (O_1208,N_24549,N_23700);
and UO_1209 (O_1209,N_23784,N_22935);
nor UO_1210 (O_1210,N_22696,N_22715);
or UO_1211 (O_1211,N_24464,N_24436);
or UO_1212 (O_1212,N_24152,N_24175);
and UO_1213 (O_1213,N_24504,N_22672);
and UO_1214 (O_1214,N_23962,N_23007);
xor UO_1215 (O_1215,N_22957,N_24208);
or UO_1216 (O_1216,N_23689,N_24427);
or UO_1217 (O_1217,N_24065,N_22949);
nor UO_1218 (O_1218,N_23442,N_24043);
xor UO_1219 (O_1219,N_24657,N_24331);
nand UO_1220 (O_1220,N_24015,N_23299);
nand UO_1221 (O_1221,N_24802,N_23506);
nor UO_1222 (O_1222,N_23843,N_23147);
nand UO_1223 (O_1223,N_24131,N_22763);
nand UO_1224 (O_1224,N_24650,N_24044);
and UO_1225 (O_1225,N_23684,N_22851);
and UO_1226 (O_1226,N_24378,N_24345);
xor UO_1227 (O_1227,N_23040,N_24575);
nor UO_1228 (O_1228,N_22795,N_23492);
xnor UO_1229 (O_1229,N_22969,N_22890);
nor UO_1230 (O_1230,N_23318,N_24306);
xnor UO_1231 (O_1231,N_23833,N_24701);
and UO_1232 (O_1232,N_24312,N_24038);
or UO_1233 (O_1233,N_23660,N_22972);
xnor UO_1234 (O_1234,N_24060,N_24846);
nor UO_1235 (O_1235,N_23928,N_23130);
and UO_1236 (O_1236,N_23463,N_24194);
and UO_1237 (O_1237,N_24610,N_23561);
or UO_1238 (O_1238,N_23435,N_22716);
and UO_1239 (O_1239,N_22854,N_23146);
xor UO_1240 (O_1240,N_24848,N_22630);
nor UO_1241 (O_1241,N_23468,N_24819);
or UO_1242 (O_1242,N_23695,N_23119);
nand UO_1243 (O_1243,N_24385,N_23652);
and UO_1244 (O_1244,N_22911,N_24820);
and UO_1245 (O_1245,N_23490,N_23688);
and UO_1246 (O_1246,N_22593,N_24524);
nand UO_1247 (O_1247,N_22915,N_24016);
nor UO_1248 (O_1248,N_23676,N_24154);
or UO_1249 (O_1249,N_24606,N_24228);
or UO_1250 (O_1250,N_24502,N_22683);
nor UO_1251 (O_1251,N_23891,N_23915);
or UO_1252 (O_1252,N_23483,N_22969);
nand UO_1253 (O_1253,N_22866,N_24630);
or UO_1254 (O_1254,N_23544,N_23104);
nor UO_1255 (O_1255,N_23068,N_24932);
nand UO_1256 (O_1256,N_23577,N_23963);
nand UO_1257 (O_1257,N_23911,N_24803);
or UO_1258 (O_1258,N_24204,N_24292);
or UO_1259 (O_1259,N_24104,N_24214);
xnor UO_1260 (O_1260,N_23596,N_23980);
nor UO_1261 (O_1261,N_24051,N_24887);
nor UO_1262 (O_1262,N_23581,N_22867);
xnor UO_1263 (O_1263,N_24931,N_23141);
and UO_1264 (O_1264,N_24667,N_24004);
nor UO_1265 (O_1265,N_24869,N_23637);
or UO_1266 (O_1266,N_22745,N_23546);
nand UO_1267 (O_1267,N_22560,N_24565);
or UO_1268 (O_1268,N_24277,N_22551);
xnor UO_1269 (O_1269,N_24766,N_24556);
and UO_1270 (O_1270,N_24915,N_22804);
nand UO_1271 (O_1271,N_23539,N_24724);
nor UO_1272 (O_1272,N_23593,N_23669);
nor UO_1273 (O_1273,N_24180,N_22815);
nand UO_1274 (O_1274,N_24089,N_24643);
and UO_1275 (O_1275,N_22724,N_23604);
nand UO_1276 (O_1276,N_22710,N_24030);
and UO_1277 (O_1277,N_24305,N_23394);
nand UO_1278 (O_1278,N_24960,N_23578);
or UO_1279 (O_1279,N_23065,N_23830);
and UO_1280 (O_1280,N_24699,N_22581);
nand UO_1281 (O_1281,N_22563,N_22961);
xnor UO_1282 (O_1282,N_24104,N_23794);
or UO_1283 (O_1283,N_24567,N_22991);
or UO_1284 (O_1284,N_22574,N_22839);
xnor UO_1285 (O_1285,N_24025,N_23776);
or UO_1286 (O_1286,N_22525,N_24688);
or UO_1287 (O_1287,N_23910,N_23724);
or UO_1288 (O_1288,N_24642,N_23026);
nand UO_1289 (O_1289,N_23610,N_24460);
or UO_1290 (O_1290,N_23241,N_24568);
xnor UO_1291 (O_1291,N_24517,N_23432);
xor UO_1292 (O_1292,N_23125,N_24938);
nor UO_1293 (O_1293,N_24880,N_22909);
or UO_1294 (O_1294,N_24552,N_23581);
and UO_1295 (O_1295,N_23849,N_24841);
nor UO_1296 (O_1296,N_22941,N_23184);
xnor UO_1297 (O_1297,N_23129,N_24196);
nand UO_1298 (O_1298,N_23829,N_23674);
xnor UO_1299 (O_1299,N_22924,N_23103);
xor UO_1300 (O_1300,N_24876,N_23655);
or UO_1301 (O_1301,N_22636,N_24169);
or UO_1302 (O_1302,N_23607,N_24552);
nand UO_1303 (O_1303,N_22929,N_23118);
nand UO_1304 (O_1304,N_23382,N_22583);
or UO_1305 (O_1305,N_23163,N_23417);
and UO_1306 (O_1306,N_24100,N_24873);
nand UO_1307 (O_1307,N_23300,N_24451);
and UO_1308 (O_1308,N_23295,N_22626);
or UO_1309 (O_1309,N_23509,N_24632);
xor UO_1310 (O_1310,N_22926,N_24456);
or UO_1311 (O_1311,N_22740,N_22703);
nand UO_1312 (O_1312,N_24771,N_22698);
nand UO_1313 (O_1313,N_24948,N_23912);
nand UO_1314 (O_1314,N_23125,N_22573);
nor UO_1315 (O_1315,N_23359,N_24948);
nand UO_1316 (O_1316,N_24748,N_24610);
or UO_1317 (O_1317,N_24334,N_22626);
and UO_1318 (O_1318,N_22940,N_24699);
or UO_1319 (O_1319,N_22713,N_24290);
xor UO_1320 (O_1320,N_24545,N_23759);
or UO_1321 (O_1321,N_23160,N_24780);
nor UO_1322 (O_1322,N_23549,N_23278);
or UO_1323 (O_1323,N_23935,N_24217);
nor UO_1324 (O_1324,N_24170,N_22987);
or UO_1325 (O_1325,N_23100,N_23014);
xnor UO_1326 (O_1326,N_22955,N_24599);
or UO_1327 (O_1327,N_24489,N_23193);
nor UO_1328 (O_1328,N_23385,N_23453);
nor UO_1329 (O_1329,N_22747,N_24213);
or UO_1330 (O_1330,N_23768,N_22559);
xnor UO_1331 (O_1331,N_23679,N_24997);
nand UO_1332 (O_1332,N_24979,N_23849);
nand UO_1333 (O_1333,N_24612,N_24215);
xor UO_1334 (O_1334,N_24865,N_23935);
or UO_1335 (O_1335,N_22916,N_22892);
and UO_1336 (O_1336,N_22589,N_23535);
or UO_1337 (O_1337,N_22968,N_22662);
nand UO_1338 (O_1338,N_23088,N_22979);
nand UO_1339 (O_1339,N_22873,N_23765);
xnor UO_1340 (O_1340,N_24143,N_24216);
nor UO_1341 (O_1341,N_24500,N_22604);
or UO_1342 (O_1342,N_24473,N_24400);
and UO_1343 (O_1343,N_24148,N_24346);
nor UO_1344 (O_1344,N_23853,N_23687);
and UO_1345 (O_1345,N_24912,N_24275);
nand UO_1346 (O_1346,N_24767,N_24238);
or UO_1347 (O_1347,N_23742,N_24450);
nand UO_1348 (O_1348,N_22681,N_24634);
nand UO_1349 (O_1349,N_23950,N_24306);
xor UO_1350 (O_1350,N_23435,N_23756);
xnor UO_1351 (O_1351,N_24317,N_24723);
xor UO_1352 (O_1352,N_22814,N_23733);
and UO_1353 (O_1353,N_24504,N_22804);
nand UO_1354 (O_1354,N_24235,N_23431);
nand UO_1355 (O_1355,N_23842,N_23605);
and UO_1356 (O_1356,N_23868,N_22611);
xor UO_1357 (O_1357,N_23651,N_24666);
xor UO_1358 (O_1358,N_24497,N_24444);
or UO_1359 (O_1359,N_24125,N_23593);
nor UO_1360 (O_1360,N_22742,N_23762);
nand UO_1361 (O_1361,N_23380,N_22981);
xnor UO_1362 (O_1362,N_22516,N_24733);
nor UO_1363 (O_1363,N_23769,N_24714);
nor UO_1364 (O_1364,N_24911,N_23302);
xnor UO_1365 (O_1365,N_23421,N_24904);
nor UO_1366 (O_1366,N_24197,N_23472);
or UO_1367 (O_1367,N_22595,N_23803);
or UO_1368 (O_1368,N_24135,N_22861);
or UO_1369 (O_1369,N_24124,N_23982);
xnor UO_1370 (O_1370,N_22972,N_22790);
and UO_1371 (O_1371,N_24053,N_23548);
xnor UO_1372 (O_1372,N_24627,N_24232);
nor UO_1373 (O_1373,N_23743,N_23366);
xnor UO_1374 (O_1374,N_23164,N_24254);
nand UO_1375 (O_1375,N_24131,N_24417);
xor UO_1376 (O_1376,N_24592,N_23980);
xor UO_1377 (O_1377,N_22732,N_23158);
or UO_1378 (O_1378,N_24162,N_24252);
and UO_1379 (O_1379,N_23480,N_23149);
nand UO_1380 (O_1380,N_24921,N_23984);
nand UO_1381 (O_1381,N_24584,N_24509);
or UO_1382 (O_1382,N_22576,N_22829);
nor UO_1383 (O_1383,N_24084,N_23230);
or UO_1384 (O_1384,N_24631,N_24015);
or UO_1385 (O_1385,N_24453,N_23625);
xnor UO_1386 (O_1386,N_24497,N_22656);
nor UO_1387 (O_1387,N_24699,N_22570);
or UO_1388 (O_1388,N_24325,N_23982);
or UO_1389 (O_1389,N_22712,N_23480);
nor UO_1390 (O_1390,N_23844,N_22526);
nand UO_1391 (O_1391,N_23824,N_24929);
and UO_1392 (O_1392,N_23025,N_24586);
nand UO_1393 (O_1393,N_24113,N_24046);
xnor UO_1394 (O_1394,N_24959,N_24766);
nor UO_1395 (O_1395,N_24559,N_22814);
and UO_1396 (O_1396,N_24287,N_24562);
and UO_1397 (O_1397,N_22826,N_24083);
nor UO_1398 (O_1398,N_24192,N_23812);
nor UO_1399 (O_1399,N_23247,N_24745);
nor UO_1400 (O_1400,N_22622,N_22649);
and UO_1401 (O_1401,N_22728,N_24120);
and UO_1402 (O_1402,N_23864,N_24721);
nand UO_1403 (O_1403,N_24214,N_23038);
nand UO_1404 (O_1404,N_23241,N_24327);
nor UO_1405 (O_1405,N_22528,N_23400);
and UO_1406 (O_1406,N_22954,N_22635);
and UO_1407 (O_1407,N_24369,N_24875);
nor UO_1408 (O_1408,N_23031,N_22989);
or UO_1409 (O_1409,N_23396,N_22793);
nand UO_1410 (O_1410,N_23217,N_23069);
nand UO_1411 (O_1411,N_23032,N_22876);
and UO_1412 (O_1412,N_24789,N_24381);
and UO_1413 (O_1413,N_23384,N_24704);
nand UO_1414 (O_1414,N_23435,N_24172);
nor UO_1415 (O_1415,N_24045,N_24253);
nand UO_1416 (O_1416,N_22707,N_23224);
nand UO_1417 (O_1417,N_23997,N_24777);
nor UO_1418 (O_1418,N_24334,N_24199);
nor UO_1419 (O_1419,N_24262,N_24369);
and UO_1420 (O_1420,N_23527,N_24490);
nor UO_1421 (O_1421,N_24842,N_23070);
and UO_1422 (O_1422,N_24394,N_24289);
nand UO_1423 (O_1423,N_23366,N_22948);
xor UO_1424 (O_1424,N_23341,N_24475);
and UO_1425 (O_1425,N_24572,N_23078);
nor UO_1426 (O_1426,N_23384,N_23403);
or UO_1427 (O_1427,N_23886,N_24100);
nor UO_1428 (O_1428,N_22513,N_24755);
and UO_1429 (O_1429,N_24549,N_23551);
nor UO_1430 (O_1430,N_24746,N_22541);
xnor UO_1431 (O_1431,N_24927,N_22753);
nor UO_1432 (O_1432,N_23291,N_24909);
and UO_1433 (O_1433,N_24090,N_24003);
nand UO_1434 (O_1434,N_24876,N_22515);
nand UO_1435 (O_1435,N_22695,N_24822);
and UO_1436 (O_1436,N_23820,N_23093);
nor UO_1437 (O_1437,N_23177,N_23855);
or UO_1438 (O_1438,N_23536,N_23712);
xor UO_1439 (O_1439,N_24947,N_22554);
or UO_1440 (O_1440,N_24992,N_24007);
xnor UO_1441 (O_1441,N_24012,N_23754);
xor UO_1442 (O_1442,N_24765,N_24067);
xnor UO_1443 (O_1443,N_24439,N_23738);
nand UO_1444 (O_1444,N_22774,N_22785);
nor UO_1445 (O_1445,N_24878,N_24010);
nor UO_1446 (O_1446,N_24301,N_24640);
nand UO_1447 (O_1447,N_24578,N_24390);
nor UO_1448 (O_1448,N_23964,N_23197);
or UO_1449 (O_1449,N_24408,N_23669);
nand UO_1450 (O_1450,N_23941,N_24729);
xnor UO_1451 (O_1451,N_24047,N_23705);
or UO_1452 (O_1452,N_23351,N_23366);
nor UO_1453 (O_1453,N_23829,N_23208);
nor UO_1454 (O_1454,N_23632,N_23424);
nand UO_1455 (O_1455,N_24945,N_24258);
nand UO_1456 (O_1456,N_24076,N_24553);
nor UO_1457 (O_1457,N_23597,N_24797);
or UO_1458 (O_1458,N_23952,N_22752);
and UO_1459 (O_1459,N_23751,N_23803);
nand UO_1460 (O_1460,N_24825,N_23748);
xor UO_1461 (O_1461,N_24402,N_22802);
nand UO_1462 (O_1462,N_24045,N_23638);
xor UO_1463 (O_1463,N_23353,N_24595);
and UO_1464 (O_1464,N_22659,N_22904);
nor UO_1465 (O_1465,N_23582,N_24171);
or UO_1466 (O_1466,N_24898,N_23500);
nand UO_1467 (O_1467,N_24645,N_24582);
nand UO_1468 (O_1468,N_24180,N_23385);
and UO_1469 (O_1469,N_22615,N_23051);
xor UO_1470 (O_1470,N_24385,N_23825);
nand UO_1471 (O_1471,N_23898,N_24473);
nand UO_1472 (O_1472,N_23007,N_23719);
nor UO_1473 (O_1473,N_23280,N_24149);
and UO_1474 (O_1474,N_22650,N_23974);
nand UO_1475 (O_1475,N_24226,N_23693);
nor UO_1476 (O_1476,N_23101,N_22710);
or UO_1477 (O_1477,N_23811,N_22542);
or UO_1478 (O_1478,N_23456,N_24883);
nor UO_1479 (O_1479,N_23180,N_23629);
and UO_1480 (O_1480,N_23672,N_22947);
xor UO_1481 (O_1481,N_23929,N_24430);
nand UO_1482 (O_1482,N_23183,N_24448);
xnor UO_1483 (O_1483,N_24477,N_24804);
or UO_1484 (O_1484,N_24966,N_23978);
or UO_1485 (O_1485,N_22660,N_24837);
nor UO_1486 (O_1486,N_24104,N_24072);
nor UO_1487 (O_1487,N_24732,N_24500);
or UO_1488 (O_1488,N_23802,N_24438);
or UO_1489 (O_1489,N_22580,N_24184);
and UO_1490 (O_1490,N_22796,N_23606);
xnor UO_1491 (O_1491,N_24459,N_23107);
nor UO_1492 (O_1492,N_23540,N_22849);
xnor UO_1493 (O_1493,N_24868,N_23734);
and UO_1494 (O_1494,N_24071,N_24447);
xnor UO_1495 (O_1495,N_22964,N_23103);
nand UO_1496 (O_1496,N_23264,N_23797);
or UO_1497 (O_1497,N_24545,N_22811);
or UO_1498 (O_1498,N_23642,N_24990);
and UO_1499 (O_1499,N_23290,N_23617);
or UO_1500 (O_1500,N_23506,N_23754);
and UO_1501 (O_1501,N_22663,N_23433);
nor UO_1502 (O_1502,N_23470,N_23116);
and UO_1503 (O_1503,N_24268,N_22855);
or UO_1504 (O_1504,N_23496,N_23997);
or UO_1505 (O_1505,N_24242,N_24546);
and UO_1506 (O_1506,N_24554,N_24916);
xnor UO_1507 (O_1507,N_23343,N_22982);
nor UO_1508 (O_1508,N_24605,N_22834);
and UO_1509 (O_1509,N_23160,N_24442);
and UO_1510 (O_1510,N_22813,N_23229);
nand UO_1511 (O_1511,N_23115,N_24365);
and UO_1512 (O_1512,N_24320,N_22538);
nor UO_1513 (O_1513,N_23489,N_23290);
nand UO_1514 (O_1514,N_22625,N_24179);
xor UO_1515 (O_1515,N_24764,N_23731);
nand UO_1516 (O_1516,N_23751,N_24874);
nand UO_1517 (O_1517,N_24667,N_24555);
nand UO_1518 (O_1518,N_23998,N_24247);
or UO_1519 (O_1519,N_24594,N_22708);
nand UO_1520 (O_1520,N_23273,N_23724);
xor UO_1521 (O_1521,N_23729,N_24316);
or UO_1522 (O_1522,N_22656,N_22716);
nor UO_1523 (O_1523,N_24838,N_22959);
and UO_1524 (O_1524,N_24940,N_23899);
and UO_1525 (O_1525,N_23225,N_23446);
nand UO_1526 (O_1526,N_23337,N_24517);
or UO_1527 (O_1527,N_22582,N_22565);
and UO_1528 (O_1528,N_24794,N_24154);
nor UO_1529 (O_1529,N_23143,N_22783);
or UO_1530 (O_1530,N_22793,N_22617);
nand UO_1531 (O_1531,N_24041,N_24444);
nor UO_1532 (O_1532,N_22773,N_24023);
xor UO_1533 (O_1533,N_23648,N_23860);
or UO_1534 (O_1534,N_22976,N_24446);
xnor UO_1535 (O_1535,N_24044,N_22923);
and UO_1536 (O_1536,N_22915,N_22836);
or UO_1537 (O_1537,N_24061,N_23527);
nor UO_1538 (O_1538,N_24644,N_24151);
xor UO_1539 (O_1539,N_22534,N_24187);
nand UO_1540 (O_1540,N_23982,N_24668);
or UO_1541 (O_1541,N_22741,N_24178);
xnor UO_1542 (O_1542,N_23847,N_24573);
xnor UO_1543 (O_1543,N_23145,N_23610);
nor UO_1544 (O_1544,N_23543,N_22546);
nor UO_1545 (O_1545,N_22621,N_23038);
xor UO_1546 (O_1546,N_22940,N_23495);
or UO_1547 (O_1547,N_23056,N_24970);
nor UO_1548 (O_1548,N_23275,N_22581);
and UO_1549 (O_1549,N_24405,N_23230);
or UO_1550 (O_1550,N_23313,N_24153);
nor UO_1551 (O_1551,N_23574,N_23643);
xor UO_1552 (O_1552,N_22815,N_24654);
or UO_1553 (O_1553,N_22757,N_23330);
nand UO_1554 (O_1554,N_24944,N_23298);
nor UO_1555 (O_1555,N_23632,N_22577);
nor UO_1556 (O_1556,N_24059,N_23651);
xnor UO_1557 (O_1557,N_24090,N_24409);
or UO_1558 (O_1558,N_23976,N_24637);
xnor UO_1559 (O_1559,N_24670,N_23982);
xnor UO_1560 (O_1560,N_24991,N_23700);
and UO_1561 (O_1561,N_22648,N_24219);
and UO_1562 (O_1562,N_24308,N_23628);
or UO_1563 (O_1563,N_22639,N_22658);
nand UO_1564 (O_1564,N_24141,N_24645);
nor UO_1565 (O_1565,N_23746,N_23392);
and UO_1566 (O_1566,N_22878,N_24300);
nand UO_1567 (O_1567,N_22733,N_22835);
and UO_1568 (O_1568,N_24216,N_24981);
or UO_1569 (O_1569,N_24889,N_24209);
nor UO_1570 (O_1570,N_23421,N_24525);
nand UO_1571 (O_1571,N_24424,N_22979);
xnor UO_1572 (O_1572,N_24807,N_22559);
nand UO_1573 (O_1573,N_23821,N_23744);
and UO_1574 (O_1574,N_24034,N_23705);
nor UO_1575 (O_1575,N_22888,N_23332);
nand UO_1576 (O_1576,N_23232,N_22651);
or UO_1577 (O_1577,N_23642,N_22855);
nand UO_1578 (O_1578,N_24086,N_23851);
and UO_1579 (O_1579,N_24351,N_24961);
or UO_1580 (O_1580,N_22988,N_24397);
nand UO_1581 (O_1581,N_23901,N_24407);
or UO_1582 (O_1582,N_24902,N_24565);
or UO_1583 (O_1583,N_24861,N_23977);
xnor UO_1584 (O_1584,N_24327,N_23750);
nor UO_1585 (O_1585,N_24736,N_24726);
nand UO_1586 (O_1586,N_24653,N_22836);
and UO_1587 (O_1587,N_24468,N_24447);
nand UO_1588 (O_1588,N_24330,N_23641);
or UO_1589 (O_1589,N_24782,N_24027);
xor UO_1590 (O_1590,N_23656,N_22955);
nor UO_1591 (O_1591,N_24649,N_23695);
xor UO_1592 (O_1592,N_23487,N_24089);
and UO_1593 (O_1593,N_23322,N_23787);
nor UO_1594 (O_1594,N_22820,N_23614);
or UO_1595 (O_1595,N_22856,N_23432);
nand UO_1596 (O_1596,N_23257,N_23015);
xor UO_1597 (O_1597,N_22681,N_24322);
xnor UO_1598 (O_1598,N_24559,N_23417);
nor UO_1599 (O_1599,N_24422,N_24924);
nor UO_1600 (O_1600,N_24816,N_24587);
and UO_1601 (O_1601,N_24088,N_23468);
xor UO_1602 (O_1602,N_24464,N_24300);
xnor UO_1603 (O_1603,N_23824,N_24661);
xnor UO_1604 (O_1604,N_23623,N_23019);
and UO_1605 (O_1605,N_23298,N_24253);
xor UO_1606 (O_1606,N_23885,N_24993);
or UO_1607 (O_1607,N_24400,N_23932);
nand UO_1608 (O_1608,N_24797,N_24067);
and UO_1609 (O_1609,N_23127,N_24443);
xnor UO_1610 (O_1610,N_24910,N_23482);
xnor UO_1611 (O_1611,N_23001,N_24782);
and UO_1612 (O_1612,N_24156,N_22763);
and UO_1613 (O_1613,N_23980,N_23069);
or UO_1614 (O_1614,N_23955,N_23496);
nand UO_1615 (O_1615,N_23298,N_23059);
xor UO_1616 (O_1616,N_24854,N_23231);
nand UO_1617 (O_1617,N_24553,N_22543);
nand UO_1618 (O_1618,N_23052,N_24287);
xnor UO_1619 (O_1619,N_24476,N_23581);
and UO_1620 (O_1620,N_23767,N_24072);
and UO_1621 (O_1621,N_23710,N_24464);
nor UO_1622 (O_1622,N_23065,N_24712);
nor UO_1623 (O_1623,N_23606,N_23161);
or UO_1624 (O_1624,N_24823,N_24859);
xor UO_1625 (O_1625,N_24470,N_23380);
nor UO_1626 (O_1626,N_22769,N_22989);
and UO_1627 (O_1627,N_24062,N_23296);
nor UO_1628 (O_1628,N_23836,N_23703);
nor UO_1629 (O_1629,N_24421,N_22955);
xor UO_1630 (O_1630,N_24603,N_24055);
xnor UO_1631 (O_1631,N_24998,N_24297);
nor UO_1632 (O_1632,N_23586,N_23564);
nor UO_1633 (O_1633,N_24733,N_23408);
xnor UO_1634 (O_1634,N_24990,N_23193);
xor UO_1635 (O_1635,N_23110,N_23276);
nor UO_1636 (O_1636,N_23396,N_24794);
or UO_1637 (O_1637,N_24718,N_23112);
nand UO_1638 (O_1638,N_23789,N_23959);
and UO_1639 (O_1639,N_24111,N_23724);
xnor UO_1640 (O_1640,N_23985,N_23157);
nand UO_1641 (O_1641,N_22973,N_23035);
and UO_1642 (O_1642,N_24640,N_23559);
nand UO_1643 (O_1643,N_23227,N_23766);
and UO_1644 (O_1644,N_23720,N_22915);
xor UO_1645 (O_1645,N_23260,N_22691);
nor UO_1646 (O_1646,N_23504,N_23300);
or UO_1647 (O_1647,N_24680,N_23806);
xor UO_1648 (O_1648,N_24165,N_23859);
nand UO_1649 (O_1649,N_24305,N_24262);
nor UO_1650 (O_1650,N_24038,N_23127);
nor UO_1651 (O_1651,N_23218,N_24893);
or UO_1652 (O_1652,N_22924,N_23392);
and UO_1653 (O_1653,N_24582,N_23107);
nor UO_1654 (O_1654,N_24782,N_23920);
xor UO_1655 (O_1655,N_23485,N_23735);
nand UO_1656 (O_1656,N_24975,N_24484);
or UO_1657 (O_1657,N_23435,N_24522);
and UO_1658 (O_1658,N_22806,N_24080);
nand UO_1659 (O_1659,N_24284,N_24483);
and UO_1660 (O_1660,N_23577,N_22882);
and UO_1661 (O_1661,N_23118,N_23223);
xnor UO_1662 (O_1662,N_23737,N_22729);
or UO_1663 (O_1663,N_23500,N_24056);
or UO_1664 (O_1664,N_22931,N_24251);
or UO_1665 (O_1665,N_23400,N_23362);
nor UO_1666 (O_1666,N_23768,N_23722);
nand UO_1667 (O_1667,N_23832,N_23724);
and UO_1668 (O_1668,N_22999,N_23796);
and UO_1669 (O_1669,N_24378,N_22553);
nand UO_1670 (O_1670,N_23363,N_24923);
nor UO_1671 (O_1671,N_23164,N_24407);
nor UO_1672 (O_1672,N_23485,N_22672);
or UO_1673 (O_1673,N_23540,N_23131);
xnor UO_1674 (O_1674,N_22554,N_23100);
nor UO_1675 (O_1675,N_24738,N_24296);
and UO_1676 (O_1676,N_23607,N_23792);
xor UO_1677 (O_1677,N_24811,N_24180);
and UO_1678 (O_1678,N_22577,N_22847);
and UO_1679 (O_1679,N_23145,N_23505);
xor UO_1680 (O_1680,N_24225,N_24457);
nor UO_1681 (O_1681,N_23273,N_22950);
or UO_1682 (O_1682,N_23292,N_23421);
xor UO_1683 (O_1683,N_22768,N_24153);
nor UO_1684 (O_1684,N_24810,N_24087);
or UO_1685 (O_1685,N_24990,N_23051);
or UO_1686 (O_1686,N_24444,N_22747);
xor UO_1687 (O_1687,N_24437,N_23844);
xnor UO_1688 (O_1688,N_23034,N_23454);
nand UO_1689 (O_1689,N_24180,N_24338);
xor UO_1690 (O_1690,N_23933,N_23347);
and UO_1691 (O_1691,N_22530,N_23550);
or UO_1692 (O_1692,N_23687,N_23759);
or UO_1693 (O_1693,N_24005,N_23450);
nand UO_1694 (O_1694,N_24395,N_24257);
nor UO_1695 (O_1695,N_23527,N_24819);
or UO_1696 (O_1696,N_22703,N_22943);
nand UO_1697 (O_1697,N_22960,N_24218);
or UO_1698 (O_1698,N_23011,N_23692);
or UO_1699 (O_1699,N_23924,N_24561);
xnor UO_1700 (O_1700,N_22782,N_22832);
or UO_1701 (O_1701,N_23589,N_23558);
nand UO_1702 (O_1702,N_24178,N_22659);
nand UO_1703 (O_1703,N_22541,N_24412);
nor UO_1704 (O_1704,N_24586,N_22931);
nand UO_1705 (O_1705,N_24453,N_24577);
nor UO_1706 (O_1706,N_24351,N_24262);
nor UO_1707 (O_1707,N_23629,N_23716);
nor UO_1708 (O_1708,N_23435,N_23947);
and UO_1709 (O_1709,N_23675,N_24917);
nand UO_1710 (O_1710,N_24484,N_24897);
and UO_1711 (O_1711,N_24103,N_23899);
and UO_1712 (O_1712,N_24056,N_24688);
and UO_1713 (O_1713,N_22537,N_22627);
and UO_1714 (O_1714,N_24017,N_23353);
or UO_1715 (O_1715,N_22740,N_24533);
nand UO_1716 (O_1716,N_23639,N_22878);
nor UO_1717 (O_1717,N_22608,N_22845);
nand UO_1718 (O_1718,N_23923,N_23269);
nand UO_1719 (O_1719,N_23183,N_23772);
and UO_1720 (O_1720,N_24098,N_23116);
nand UO_1721 (O_1721,N_24883,N_23453);
nor UO_1722 (O_1722,N_22727,N_22543);
nand UO_1723 (O_1723,N_22534,N_22977);
nor UO_1724 (O_1724,N_24919,N_22816);
xnor UO_1725 (O_1725,N_24689,N_23692);
or UO_1726 (O_1726,N_24014,N_22767);
nor UO_1727 (O_1727,N_22803,N_23567);
nor UO_1728 (O_1728,N_24084,N_24960);
nand UO_1729 (O_1729,N_24827,N_22542);
xnor UO_1730 (O_1730,N_23211,N_22882);
nand UO_1731 (O_1731,N_24661,N_24524);
or UO_1732 (O_1732,N_24764,N_24176);
xnor UO_1733 (O_1733,N_24046,N_22732);
nand UO_1734 (O_1734,N_24418,N_22825);
nor UO_1735 (O_1735,N_24654,N_24266);
nand UO_1736 (O_1736,N_24175,N_22739);
nand UO_1737 (O_1737,N_23314,N_24451);
nand UO_1738 (O_1738,N_22656,N_24119);
nand UO_1739 (O_1739,N_23083,N_24958);
xor UO_1740 (O_1740,N_23283,N_24039);
or UO_1741 (O_1741,N_23246,N_24950);
nor UO_1742 (O_1742,N_23947,N_24948);
or UO_1743 (O_1743,N_24143,N_23262);
nand UO_1744 (O_1744,N_23102,N_24903);
nand UO_1745 (O_1745,N_23990,N_22520);
nor UO_1746 (O_1746,N_23054,N_22900);
or UO_1747 (O_1747,N_24286,N_24462);
nand UO_1748 (O_1748,N_23930,N_24515);
nor UO_1749 (O_1749,N_24549,N_24064);
nand UO_1750 (O_1750,N_23042,N_23076);
or UO_1751 (O_1751,N_23174,N_23346);
nand UO_1752 (O_1752,N_23224,N_23120);
nand UO_1753 (O_1753,N_23110,N_22912);
nor UO_1754 (O_1754,N_24248,N_24609);
or UO_1755 (O_1755,N_23934,N_23983);
nand UO_1756 (O_1756,N_22672,N_23548);
nor UO_1757 (O_1757,N_23390,N_24422);
nor UO_1758 (O_1758,N_24117,N_24501);
nor UO_1759 (O_1759,N_22656,N_22782);
or UO_1760 (O_1760,N_24754,N_22848);
nor UO_1761 (O_1761,N_24149,N_24348);
nand UO_1762 (O_1762,N_24288,N_24822);
and UO_1763 (O_1763,N_24468,N_23559);
nor UO_1764 (O_1764,N_23449,N_23158);
and UO_1765 (O_1765,N_24582,N_22837);
nand UO_1766 (O_1766,N_23777,N_23164);
nand UO_1767 (O_1767,N_23724,N_24234);
nand UO_1768 (O_1768,N_23371,N_22996);
xor UO_1769 (O_1769,N_22957,N_22538);
nand UO_1770 (O_1770,N_23746,N_22891);
xnor UO_1771 (O_1771,N_23291,N_23481);
or UO_1772 (O_1772,N_23800,N_23322);
nor UO_1773 (O_1773,N_22749,N_24253);
nor UO_1774 (O_1774,N_23579,N_23363);
xor UO_1775 (O_1775,N_24832,N_24599);
or UO_1776 (O_1776,N_24946,N_23069);
and UO_1777 (O_1777,N_23566,N_24410);
nand UO_1778 (O_1778,N_22890,N_24113);
xnor UO_1779 (O_1779,N_23665,N_22729);
nor UO_1780 (O_1780,N_23177,N_24821);
nor UO_1781 (O_1781,N_23262,N_22680);
and UO_1782 (O_1782,N_24458,N_23951);
and UO_1783 (O_1783,N_23688,N_24772);
and UO_1784 (O_1784,N_23714,N_24112);
xnor UO_1785 (O_1785,N_22845,N_23882);
xor UO_1786 (O_1786,N_24851,N_23629);
nor UO_1787 (O_1787,N_22992,N_23655);
or UO_1788 (O_1788,N_24053,N_23300);
xor UO_1789 (O_1789,N_23304,N_23835);
nor UO_1790 (O_1790,N_24832,N_24673);
and UO_1791 (O_1791,N_24097,N_24684);
nand UO_1792 (O_1792,N_24470,N_23504);
or UO_1793 (O_1793,N_23965,N_22835);
and UO_1794 (O_1794,N_22996,N_24037);
xnor UO_1795 (O_1795,N_23966,N_22806);
and UO_1796 (O_1796,N_23251,N_23094);
xnor UO_1797 (O_1797,N_23722,N_24694);
nor UO_1798 (O_1798,N_24324,N_23713);
nor UO_1799 (O_1799,N_24726,N_23032);
and UO_1800 (O_1800,N_24977,N_24704);
xor UO_1801 (O_1801,N_23467,N_22798);
or UO_1802 (O_1802,N_23845,N_24907);
or UO_1803 (O_1803,N_22735,N_22676);
or UO_1804 (O_1804,N_24626,N_24072);
nand UO_1805 (O_1805,N_24909,N_23697);
nand UO_1806 (O_1806,N_22533,N_23176);
nand UO_1807 (O_1807,N_24624,N_23618);
and UO_1808 (O_1808,N_24085,N_23046);
xnor UO_1809 (O_1809,N_24846,N_22856);
and UO_1810 (O_1810,N_24911,N_23613);
nand UO_1811 (O_1811,N_22646,N_24295);
xnor UO_1812 (O_1812,N_22821,N_24977);
nand UO_1813 (O_1813,N_24107,N_24998);
nand UO_1814 (O_1814,N_23347,N_22611);
nor UO_1815 (O_1815,N_24938,N_24478);
xnor UO_1816 (O_1816,N_24843,N_22930);
nand UO_1817 (O_1817,N_23944,N_22633);
and UO_1818 (O_1818,N_23182,N_22975);
nor UO_1819 (O_1819,N_22673,N_22993);
or UO_1820 (O_1820,N_24379,N_23433);
and UO_1821 (O_1821,N_23278,N_23518);
and UO_1822 (O_1822,N_23804,N_22741);
nand UO_1823 (O_1823,N_24853,N_22952);
or UO_1824 (O_1824,N_24494,N_24164);
nor UO_1825 (O_1825,N_23137,N_24333);
nor UO_1826 (O_1826,N_22895,N_23150);
and UO_1827 (O_1827,N_23248,N_24864);
or UO_1828 (O_1828,N_23971,N_24479);
xnor UO_1829 (O_1829,N_24030,N_24696);
xor UO_1830 (O_1830,N_24341,N_23477);
xor UO_1831 (O_1831,N_24745,N_24676);
nor UO_1832 (O_1832,N_24135,N_24537);
nor UO_1833 (O_1833,N_24061,N_23903);
nand UO_1834 (O_1834,N_24384,N_23678);
nand UO_1835 (O_1835,N_22598,N_24023);
or UO_1836 (O_1836,N_23991,N_23171);
or UO_1837 (O_1837,N_24950,N_24738);
and UO_1838 (O_1838,N_22536,N_24779);
nor UO_1839 (O_1839,N_22503,N_22638);
and UO_1840 (O_1840,N_23020,N_23781);
and UO_1841 (O_1841,N_24774,N_22523);
xor UO_1842 (O_1842,N_22695,N_23687);
nand UO_1843 (O_1843,N_23628,N_23687);
xor UO_1844 (O_1844,N_23472,N_24684);
and UO_1845 (O_1845,N_24489,N_22803);
xnor UO_1846 (O_1846,N_23743,N_24737);
or UO_1847 (O_1847,N_24223,N_23771);
nor UO_1848 (O_1848,N_24507,N_24704);
and UO_1849 (O_1849,N_23460,N_24433);
or UO_1850 (O_1850,N_22658,N_24109);
or UO_1851 (O_1851,N_24666,N_24701);
nor UO_1852 (O_1852,N_22803,N_24774);
or UO_1853 (O_1853,N_23215,N_24290);
nand UO_1854 (O_1854,N_24808,N_23679);
nand UO_1855 (O_1855,N_22681,N_22637);
and UO_1856 (O_1856,N_22534,N_23564);
and UO_1857 (O_1857,N_22774,N_24176);
nor UO_1858 (O_1858,N_22621,N_23379);
nor UO_1859 (O_1859,N_23138,N_24568);
nor UO_1860 (O_1860,N_24091,N_24891);
xor UO_1861 (O_1861,N_24611,N_23188);
nand UO_1862 (O_1862,N_23211,N_24499);
nor UO_1863 (O_1863,N_24138,N_23930);
nand UO_1864 (O_1864,N_23613,N_23616);
or UO_1865 (O_1865,N_24317,N_24379);
xor UO_1866 (O_1866,N_23672,N_23304);
and UO_1867 (O_1867,N_23067,N_22767);
xnor UO_1868 (O_1868,N_22540,N_24374);
nand UO_1869 (O_1869,N_24496,N_23211);
or UO_1870 (O_1870,N_24873,N_22971);
and UO_1871 (O_1871,N_23874,N_24162);
nand UO_1872 (O_1872,N_24078,N_23798);
xor UO_1873 (O_1873,N_24814,N_22712);
nor UO_1874 (O_1874,N_23362,N_23299);
nor UO_1875 (O_1875,N_24793,N_22997);
nand UO_1876 (O_1876,N_22854,N_23341);
and UO_1877 (O_1877,N_22635,N_23198);
nand UO_1878 (O_1878,N_23525,N_24042);
nor UO_1879 (O_1879,N_23448,N_23459);
nand UO_1880 (O_1880,N_24118,N_24006);
and UO_1881 (O_1881,N_24222,N_23337);
or UO_1882 (O_1882,N_24214,N_22512);
xor UO_1883 (O_1883,N_23141,N_22575);
xor UO_1884 (O_1884,N_24765,N_24457);
and UO_1885 (O_1885,N_23139,N_22679);
xnor UO_1886 (O_1886,N_24302,N_23031);
nand UO_1887 (O_1887,N_24048,N_23949);
nor UO_1888 (O_1888,N_24555,N_22725);
nor UO_1889 (O_1889,N_23646,N_24063);
or UO_1890 (O_1890,N_24155,N_24613);
xnor UO_1891 (O_1891,N_22903,N_24245);
nand UO_1892 (O_1892,N_22952,N_23802);
or UO_1893 (O_1893,N_23902,N_22946);
or UO_1894 (O_1894,N_22872,N_23711);
xor UO_1895 (O_1895,N_23873,N_23503);
or UO_1896 (O_1896,N_24242,N_24851);
or UO_1897 (O_1897,N_23122,N_23341);
nand UO_1898 (O_1898,N_23305,N_24910);
nand UO_1899 (O_1899,N_24006,N_23149);
xor UO_1900 (O_1900,N_23040,N_24246);
and UO_1901 (O_1901,N_23549,N_23791);
xnor UO_1902 (O_1902,N_22822,N_23131);
or UO_1903 (O_1903,N_23640,N_24022);
nand UO_1904 (O_1904,N_24668,N_23809);
nor UO_1905 (O_1905,N_24980,N_24692);
nand UO_1906 (O_1906,N_24899,N_24600);
and UO_1907 (O_1907,N_24722,N_24372);
xnor UO_1908 (O_1908,N_23244,N_22887);
nor UO_1909 (O_1909,N_24811,N_23863);
nor UO_1910 (O_1910,N_24759,N_23059);
nor UO_1911 (O_1911,N_23339,N_22571);
or UO_1912 (O_1912,N_22951,N_23251);
xnor UO_1913 (O_1913,N_23400,N_24606);
or UO_1914 (O_1914,N_22879,N_24372);
xnor UO_1915 (O_1915,N_23198,N_22846);
and UO_1916 (O_1916,N_22795,N_23219);
xor UO_1917 (O_1917,N_24685,N_23111);
nand UO_1918 (O_1918,N_23285,N_24023);
and UO_1919 (O_1919,N_22588,N_24896);
nor UO_1920 (O_1920,N_23641,N_24541);
and UO_1921 (O_1921,N_23218,N_24598);
nor UO_1922 (O_1922,N_24486,N_24124);
and UO_1923 (O_1923,N_23585,N_23240);
nor UO_1924 (O_1924,N_23071,N_23031);
xnor UO_1925 (O_1925,N_24616,N_24502);
or UO_1926 (O_1926,N_24976,N_23862);
or UO_1927 (O_1927,N_24140,N_24649);
nand UO_1928 (O_1928,N_22804,N_24528);
or UO_1929 (O_1929,N_24123,N_24627);
nand UO_1930 (O_1930,N_22525,N_23347);
nor UO_1931 (O_1931,N_23210,N_22501);
or UO_1932 (O_1932,N_24923,N_24575);
xnor UO_1933 (O_1933,N_23710,N_22927);
xnor UO_1934 (O_1934,N_22536,N_23674);
xor UO_1935 (O_1935,N_24483,N_22743);
nand UO_1936 (O_1936,N_23192,N_23818);
xnor UO_1937 (O_1937,N_23812,N_24004);
or UO_1938 (O_1938,N_22916,N_24053);
or UO_1939 (O_1939,N_24238,N_24747);
nor UO_1940 (O_1940,N_23559,N_23222);
or UO_1941 (O_1941,N_24437,N_23007);
and UO_1942 (O_1942,N_22604,N_24603);
nand UO_1943 (O_1943,N_22803,N_24168);
or UO_1944 (O_1944,N_24010,N_23749);
nand UO_1945 (O_1945,N_24388,N_24970);
nand UO_1946 (O_1946,N_23943,N_23866);
and UO_1947 (O_1947,N_23603,N_23744);
nor UO_1948 (O_1948,N_23396,N_24371);
and UO_1949 (O_1949,N_24063,N_22700);
nand UO_1950 (O_1950,N_22883,N_24813);
nand UO_1951 (O_1951,N_23736,N_24665);
nand UO_1952 (O_1952,N_23482,N_23794);
nor UO_1953 (O_1953,N_24124,N_23693);
xor UO_1954 (O_1954,N_24357,N_22912);
nor UO_1955 (O_1955,N_24251,N_24566);
xor UO_1956 (O_1956,N_23049,N_23486);
nand UO_1957 (O_1957,N_23110,N_24722);
or UO_1958 (O_1958,N_24786,N_24401);
nand UO_1959 (O_1959,N_22934,N_23955);
nor UO_1960 (O_1960,N_24673,N_23368);
or UO_1961 (O_1961,N_24581,N_23661);
nor UO_1962 (O_1962,N_24083,N_22983);
nand UO_1963 (O_1963,N_22789,N_23931);
nor UO_1964 (O_1964,N_23806,N_23415);
xnor UO_1965 (O_1965,N_23302,N_24929);
xnor UO_1966 (O_1966,N_23119,N_22541);
or UO_1967 (O_1967,N_23184,N_24199);
nand UO_1968 (O_1968,N_24178,N_23576);
nor UO_1969 (O_1969,N_24714,N_24106);
or UO_1970 (O_1970,N_24481,N_23868);
or UO_1971 (O_1971,N_23183,N_23005);
nor UO_1972 (O_1972,N_22552,N_24617);
and UO_1973 (O_1973,N_23749,N_24687);
or UO_1974 (O_1974,N_23324,N_24776);
nand UO_1975 (O_1975,N_23245,N_24920);
nor UO_1976 (O_1976,N_24672,N_24092);
nand UO_1977 (O_1977,N_22883,N_22976);
nor UO_1978 (O_1978,N_22812,N_24255);
and UO_1979 (O_1979,N_23608,N_24949);
or UO_1980 (O_1980,N_23990,N_22768);
nand UO_1981 (O_1981,N_24558,N_24871);
or UO_1982 (O_1982,N_23682,N_24123);
xnor UO_1983 (O_1983,N_23297,N_23051);
xnor UO_1984 (O_1984,N_23240,N_24659);
nand UO_1985 (O_1985,N_23690,N_22637);
and UO_1986 (O_1986,N_24783,N_22967);
or UO_1987 (O_1987,N_22638,N_24683);
nand UO_1988 (O_1988,N_22609,N_22918);
xor UO_1989 (O_1989,N_24402,N_23131);
and UO_1990 (O_1990,N_22810,N_24854);
and UO_1991 (O_1991,N_24731,N_24699);
xnor UO_1992 (O_1992,N_22709,N_23832);
or UO_1993 (O_1993,N_22813,N_23963);
nor UO_1994 (O_1994,N_23947,N_23047);
or UO_1995 (O_1995,N_23213,N_24817);
or UO_1996 (O_1996,N_23648,N_24774);
xnor UO_1997 (O_1997,N_23436,N_23265);
nand UO_1998 (O_1998,N_23746,N_23352);
nor UO_1999 (O_1999,N_24594,N_23976);
nor UO_2000 (O_2000,N_24802,N_23416);
xnor UO_2001 (O_2001,N_24133,N_22550);
and UO_2002 (O_2002,N_23096,N_24749);
xor UO_2003 (O_2003,N_24709,N_23134);
and UO_2004 (O_2004,N_22687,N_24936);
xor UO_2005 (O_2005,N_22710,N_22531);
xor UO_2006 (O_2006,N_24231,N_24194);
or UO_2007 (O_2007,N_22703,N_22728);
nand UO_2008 (O_2008,N_22616,N_24280);
nor UO_2009 (O_2009,N_23937,N_22672);
nor UO_2010 (O_2010,N_24961,N_22915);
or UO_2011 (O_2011,N_23864,N_22808);
and UO_2012 (O_2012,N_22899,N_23992);
or UO_2013 (O_2013,N_24573,N_23609);
and UO_2014 (O_2014,N_24439,N_24881);
and UO_2015 (O_2015,N_22877,N_23767);
nor UO_2016 (O_2016,N_23598,N_22638);
and UO_2017 (O_2017,N_22519,N_23578);
and UO_2018 (O_2018,N_24115,N_23068);
nand UO_2019 (O_2019,N_24315,N_24113);
xnor UO_2020 (O_2020,N_23658,N_22808);
xor UO_2021 (O_2021,N_22906,N_24832);
nor UO_2022 (O_2022,N_22850,N_23700);
xor UO_2023 (O_2023,N_24743,N_23264);
and UO_2024 (O_2024,N_23645,N_23981);
nor UO_2025 (O_2025,N_23905,N_24756);
nor UO_2026 (O_2026,N_23720,N_24185);
or UO_2027 (O_2027,N_22741,N_23258);
xnor UO_2028 (O_2028,N_22563,N_24285);
or UO_2029 (O_2029,N_24505,N_23369);
nand UO_2030 (O_2030,N_24278,N_23672);
nor UO_2031 (O_2031,N_24849,N_22985);
and UO_2032 (O_2032,N_23570,N_24280);
and UO_2033 (O_2033,N_23960,N_24781);
xnor UO_2034 (O_2034,N_24571,N_23376);
nand UO_2035 (O_2035,N_24111,N_24967);
and UO_2036 (O_2036,N_23463,N_24712);
xnor UO_2037 (O_2037,N_23052,N_23167);
xor UO_2038 (O_2038,N_23057,N_23370);
nand UO_2039 (O_2039,N_22714,N_23643);
xor UO_2040 (O_2040,N_22737,N_22538);
or UO_2041 (O_2041,N_22583,N_24774);
or UO_2042 (O_2042,N_23333,N_22775);
xor UO_2043 (O_2043,N_23867,N_23208);
nor UO_2044 (O_2044,N_24616,N_24466);
xnor UO_2045 (O_2045,N_23651,N_24969);
xnor UO_2046 (O_2046,N_24940,N_23251);
or UO_2047 (O_2047,N_23483,N_23905);
and UO_2048 (O_2048,N_24166,N_22665);
xnor UO_2049 (O_2049,N_23569,N_24830);
nand UO_2050 (O_2050,N_22519,N_24496);
and UO_2051 (O_2051,N_24758,N_22672);
nor UO_2052 (O_2052,N_23691,N_24137);
and UO_2053 (O_2053,N_23880,N_24963);
and UO_2054 (O_2054,N_24132,N_23778);
xnor UO_2055 (O_2055,N_24219,N_22842);
and UO_2056 (O_2056,N_22538,N_23251);
and UO_2057 (O_2057,N_23236,N_24416);
nor UO_2058 (O_2058,N_23056,N_23675);
and UO_2059 (O_2059,N_23560,N_23730);
and UO_2060 (O_2060,N_23187,N_23663);
xnor UO_2061 (O_2061,N_24931,N_22569);
or UO_2062 (O_2062,N_23371,N_22986);
xor UO_2063 (O_2063,N_24350,N_24598);
nor UO_2064 (O_2064,N_24786,N_23893);
and UO_2065 (O_2065,N_24159,N_24917);
xor UO_2066 (O_2066,N_24487,N_23547);
nor UO_2067 (O_2067,N_22885,N_22897);
nor UO_2068 (O_2068,N_24917,N_24125);
and UO_2069 (O_2069,N_23483,N_24544);
nand UO_2070 (O_2070,N_24102,N_24484);
or UO_2071 (O_2071,N_24445,N_22578);
nand UO_2072 (O_2072,N_23052,N_24989);
and UO_2073 (O_2073,N_23104,N_22858);
and UO_2074 (O_2074,N_24057,N_23525);
and UO_2075 (O_2075,N_22528,N_23426);
xor UO_2076 (O_2076,N_22556,N_24734);
or UO_2077 (O_2077,N_23431,N_22686);
nand UO_2078 (O_2078,N_24871,N_23569);
nor UO_2079 (O_2079,N_24556,N_23322);
nor UO_2080 (O_2080,N_24643,N_24315);
and UO_2081 (O_2081,N_23786,N_24963);
or UO_2082 (O_2082,N_23937,N_23137);
and UO_2083 (O_2083,N_24734,N_23150);
and UO_2084 (O_2084,N_24824,N_24755);
or UO_2085 (O_2085,N_23924,N_22819);
nor UO_2086 (O_2086,N_22857,N_24471);
nor UO_2087 (O_2087,N_23426,N_22934);
or UO_2088 (O_2088,N_22746,N_22512);
or UO_2089 (O_2089,N_24016,N_24560);
nand UO_2090 (O_2090,N_24303,N_23035);
nor UO_2091 (O_2091,N_24314,N_24436);
nor UO_2092 (O_2092,N_24987,N_23537);
nand UO_2093 (O_2093,N_23344,N_24572);
and UO_2094 (O_2094,N_24138,N_24567);
xnor UO_2095 (O_2095,N_23594,N_23050);
nor UO_2096 (O_2096,N_23731,N_23272);
nand UO_2097 (O_2097,N_23596,N_23886);
or UO_2098 (O_2098,N_22592,N_24810);
and UO_2099 (O_2099,N_23473,N_24420);
and UO_2100 (O_2100,N_23776,N_22818);
nor UO_2101 (O_2101,N_22646,N_22933);
nor UO_2102 (O_2102,N_24116,N_24115);
or UO_2103 (O_2103,N_23930,N_23905);
xnor UO_2104 (O_2104,N_22969,N_23563);
and UO_2105 (O_2105,N_24819,N_23025);
nand UO_2106 (O_2106,N_22851,N_23290);
xor UO_2107 (O_2107,N_23669,N_22553);
or UO_2108 (O_2108,N_24150,N_24055);
nor UO_2109 (O_2109,N_23804,N_24769);
or UO_2110 (O_2110,N_24084,N_23451);
or UO_2111 (O_2111,N_22804,N_23412);
nor UO_2112 (O_2112,N_24813,N_24265);
nand UO_2113 (O_2113,N_24390,N_23456);
xnor UO_2114 (O_2114,N_23174,N_24737);
xnor UO_2115 (O_2115,N_23422,N_23603);
xnor UO_2116 (O_2116,N_24984,N_24005);
xnor UO_2117 (O_2117,N_23680,N_22724);
xor UO_2118 (O_2118,N_23383,N_24088);
and UO_2119 (O_2119,N_24249,N_24192);
and UO_2120 (O_2120,N_23946,N_23727);
or UO_2121 (O_2121,N_24067,N_24165);
nor UO_2122 (O_2122,N_24918,N_24344);
nand UO_2123 (O_2123,N_22825,N_22855);
or UO_2124 (O_2124,N_23189,N_22891);
xor UO_2125 (O_2125,N_23375,N_22733);
or UO_2126 (O_2126,N_24077,N_24520);
nand UO_2127 (O_2127,N_22643,N_23012);
xnor UO_2128 (O_2128,N_22864,N_23263);
and UO_2129 (O_2129,N_23716,N_23284);
and UO_2130 (O_2130,N_24217,N_24748);
nand UO_2131 (O_2131,N_23398,N_22968);
xor UO_2132 (O_2132,N_24249,N_22687);
and UO_2133 (O_2133,N_24332,N_24217);
and UO_2134 (O_2134,N_23126,N_24628);
nor UO_2135 (O_2135,N_22942,N_24216);
nor UO_2136 (O_2136,N_24303,N_22705);
or UO_2137 (O_2137,N_24429,N_22670);
nor UO_2138 (O_2138,N_24386,N_24318);
nor UO_2139 (O_2139,N_23327,N_22737);
nand UO_2140 (O_2140,N_22606,N_24667);
and UO_2141 (O_2141,N_24531,N_23639);
xnor UO_2142 (O_2142,N_24462,N_24531);
and UO_2143 (O_2143,N_22500,N_23863);
nor UO_2144 (O_2144,N_24066,N_23794);
and UO_2145 (O_2145,N_24670,N_23913);
and UO_2146 (O_2146,N_24505,N_22678);
nor UO_2147 (O_2147,N_23920,N_22880);
nand UO_2148 (O_2148,N_22597,N_22857);
and UO_2149 (O_2149,N_23722,N_22911);
xnor UO_2150 (O_2150,N_24781,N_24947);
xor UO_2151 (O_2151,N_22703,N_23191);
nand UO_2152 (O_2152,N_24147,N_24337);
nand UO_2153 (O_2153,N_23987,N_23606);
and UO_2154 (O_2154,N_22795,N_23694);
xnor UO_2155 (O_2155,N_23472,N_24735);
xor UO_2156 (O_2156,N_22679,N_23764);
nand UO_2157 (O_2157,N_22983,N_23929);
nand UO_2158 (O_2158,N_22708,N_24981);
nor UO_2159 (O_2159,N_24090,N_23205);
xnor UO_2160 (O_2160,N_23070,N_23621);
nand UO_2161 (O_2161,N_24281,N_22643);
nand UO_2162 (O_2162,N_24192,N_22573);
nand UO_2163 (O_2163,N_24593,N_23929);
and UO_2164 (O_2164,N_24335,N_23685);
nand UO_2165 (O_2165,N_24328,N_24296);
xnor UO_2166 (O_2166,N_24475,N_22846);
nor UO_2167 (O_2167,N_23930,N_23764);
and UO_2168 (O_2168,N_23549,N_22908);
or UO_2169 (O_2169,N_24575,N_24895);
and UO_2170 (O_2170,N_23831,N_23692);
xnor UO_2171 (O_2171,N_24223,N_22864);
and UO_2172 (O_2172,N_24926,N_24381);
and UO_2173 (O_2173,N_24203,N_23099);
nand UO_2174 (O_2174,N_24496,N_24453);
nand UO_2175 (O_2175,N_23194,N_22703);
or UO_2176 (O_2176,N_23172,N_22847);
xor UO_2177 (O_2177,N_23413,N_23766);
or UO_2178 (O_2178,N_22994,N_22597);
nor UO_2179 (O_2179,N_23886,N_23539);
and UO_2180 (O_2180,N_24306,N_22607);
and UO_2181 (O_2181,N_22660,N_23937);
nor UO_2182 (O_2182,N_24924,N_24507);
xnor UO_2183 (O_2183,N_23278,N_23399);
or UO_2184 (O_2184,N_24449,N_24835);
and UO_2185 (O_2185,N_24744,N_24792);
or UO_2186 (O_2186,N_24419,N_23375);
nor UO_2187 (O_2187,N_24532,N_24925);
and UO_2188 (O_2188,N_23013,N_23416);
or UO_2189 (O_2189,N_24626,N_24102);
and UO_2190 (O_2190,N_24901,N_24585);
and UO_2191 (O_2191,N_22601,N_22932);
and UO_2192 (O_2192,N_23057,N_22636);
nor UO_2193 (O_2193,N_24378,N_23687);
and UO_2194 (O_2194,N_22501,N_24904);
or UO_2195 (O_2195,N_22923,N_23257);
or UO_2196 (O_2196,N_23852,N_22886);
xor UO_2197 (O_2197,N_23642,N_24741);
or UO_2198 (O_2198,N_22986,N_23302);
or UO_2199 (O_2199,N_23088,N_23543);
nor UO_2200 (O_2200,N_23831,N_23467);
xor UO_2201 (O_2201,N_23676,N_22834);
or UO_2202 (O_2202,N_24064,N_24327);
xor UO_2203 (O_2203,N_24053,N_24184);
nor UO_2204 (O_2204,N_24431,N_24199);
and UO_2205 (O_2205,N_23809,N_23618);
nand UO_2206 (O_2206,N_24283,N_23372);
and UO_2207 (O_2207,N_23777,N_23818);
nor UO_2208 (O_2208,N_22660,N_23298);
or UO_2209 (O_2209,N_24898,N_24623);
and UO_2210 (O_2210,N_24902,N_23364);
xnor UO_2211 (O_2211,N_22719,N_23230);
nand UO_2212 (O_2212,N_23454,N_23367);
or UO_2213 (O_2213,N_24558,N_23870);
xor UO_2214 (O_2214,N_23770,N_24042);
and UO_2215 (O_2215,N_23733,N_24359);
nor UO_2216 (O_2216,N_24181,N_24191);
nor UO_2217 (O_2217,N_24799,N_22674);
xnor UO_2218 (O_2218,N_24260,N_23176);
nor UO_2219 (O_2219,N_24678,N_24951);
or UO_2220 (O_2220,N_23218,N_24760);
or UO_2221 (O_2221,N_23820,N_24369);
or UO_2222 (O_2222,N_24775,N_22924);
or UO_2223 (O_2223,N_23756,N_22529);
or UO_2224 (O_2224,N_23956,N_23202);
or UO_2225 (O_2225,N_24444,N_24829);
and UO_2226 (O_2226,N_24497,N_23925);
xor UO_2227 (O_2227,N_23906,N_24118);
nand UO_2228 (O_2228,N_24051,N_23504);
or UO_2229 (O_2229,N_24193,N_24011);
or UO_2230 (O_2230,N_23003,N_24054);
or UO_2231 (O_2231,N_24894,N_22517);
nand UO_2232 (O_2232,N_23775,N_23372);
xnor UO_2233 (O_2233,N_22656,N_24390);
and UO_2234 (O_2234,N_24312,N_24791);
xnor UO_2235 (O_2235,N_23462,N_24756);
xnor UO_2236 (O_2236,N_24731,N_23418);
or UO_2237 (O_2237,N_23581,N_23739);
nand UO_2238 (O_2238,N_23021,N_24689);
nand UO_2239 (O_2239,N_23360,N_24523);
nor UO_2240 (O_2240,N_24498,N_24760);
or UO_2241 (O_2241,N_24550,N_22845);
or UO_2242 (O_2242,N_24801,N_22975);
and UO_2243 (O_2243,N_24216,N_23935);
or UO_2244 (O_2244,N_22717,N_23278);
xnor UO_2245 (O_2245,N_23089,N_23182);
and UO_2246 (O_2246,N_22892,N_24721);
and UO_2247 (O_2247,N_23777,N_22740);
or UO_2248 (O_2248,N_23659,N_22645);
xnor UO_2249 (O_2249,N_22596,N_24052);
and UO_2250 (O_2250,N_23102,N_22580);
or UO_2251 (O_2251,N_23064,N_24223);
or UO_2252 (O_2252,N_23463,N_23442);
nor UO_2253 (O_2253,N_23018,N_24468);
nand UO_2254 (O_2254,N_24540,N_24386);
and UO_2255 (O_2255,N_23809,N_24239);
or UO_2256 (O_2256,N_24819,N_24032);
and UO_2257 (O_2257,N_23350,N_23650);
nor UO_2258 (O_2258,N_23648,N_23921);
or UO_2259 (O_2259,N_24070,N_24734);
and UO_2260 (O_2260,N_23456,N_22638);
nor UO_2261 (O_2261,N_24327,N_22580);
and UO_2262 (O_2262,N_23024,N_24537);
xnor UO_2263 (O_2263,N_23111,N_23075);
and UO_2264 (O_2264,N_23633,N_23177);
or UO_2265 (O_2265,N_24913,N_24485);
nand UO_2266 (O_2266,N_23945,N_22517);
or UO_2267 (O_2267,N_22596,N_22953);
nor UO_2268 (O_2268,N_23595,N_24386);
and UO_2269 (O_2269,N_24320,N_23498);
nor UO_2270 (O_2270,N_22673,N_24671);
and UO_2271 (O_2271,N_23645,N_24291);
xor UO_2272 (O_2272,N_22795,N_24098);
nand UO_2273 (O_2273,N_23047,N_24536);
and UO_2274 (O_2274,N_23967,N_23447);
nand UO_2275 (O_2275,N_24788,N_23353);
and UO_2276 (O_2276,N_24284,N_24161);
xor UO_2277 (O_2277,N_24581,N_23948);
or UO_2278 (O_2278,N_23804,N_23143);
or UO_2279 (O_2279,N_24840,N_24951);
nand UO_2280 (O_2280,N_24146,N_23913);
nand UO_2281 (O_2281,N_24534,N_22559);
xnor UO_2282 (O_2282,N_24503,N_22844);
nand UO_2283 (O_2283,N_24375,N_24298);
and UO_2284 (O_2284,N_23415,N_23310);
or UO_2285 (O_2285,N_24050,N_23487);
nor UO_2286 (O_2286,N_24749,N_24993);
nor UO_2287 (O_2287,N_23549,N_24730);
and UO_2288 (O_2288,N_23584,N_22688);
nor UO_2289 (O_2289,N_23755,N_23304);
and UO_2290 (O_2290,N_22749,N_23413);
and UO_2291 (O_2291,N_24511,N_24691);
xnor UO_2292 (O_2292,N_22850,N_23354);
xor UO_2293 (O_2293,N_23988,N_23907);
or UO_2294 (O_2294,N_23024,N_22775);
or UO_2295 (O_2295,N_24673,N_23017);
nor UO_2296 (O_2296,N_23157,N_24989);
and UO_2297 (O_2297,N_23441,N_23143);
xnor UO_2298 (O_2298,N_23194,N_22958);
or UO_2299 (O_2299,N_24712,N_23016);
or UO_2300 (O_2300,N_22950,N_23902);
nand UO_2301 (O_2301,N_23314,N_22799);
nand UO_2302 (O_2302,N_22801,N_23002);
nand UO_2303 (O_2303,N_23066,N_24817);
nor UO_2304 (O_2304,N_24107,N_22849);
or UO_2305 (O_2305,N_23519,N_23114);
and UO_2306 (O_2306,N_24789,N_23893);
nand UO_2307 (O_2307,N_24285,N_24049);
or UO_2308 (O_2308,N_22902,N_23284);
or UO_2309 (O_2309,N_23812,N_22701);
nor UO_2310 (O_2310,N_23100,N_22918);
and UO_2311 (O_2311,N_23268,N_24298);
xor UO_2312 (O_2312,N_23873,N_24004);
xor UO_2313 (O_2313,N_22633,N_24105);
or UO_2314 (O_2314,N_23977,N_24721);
and UO_2315 (O_2315,N_23022,N_24199);
nand UO_2316 (O_2316,N_24911,N_22649);
xor UO_2317 (O_2317,N_24046,N_22532);
xnor UO_2318 (O_2318,N_24835,N_24442);
nor UO_2319 (O_2319,N_24574,N_23716);
nand UO_2320 (O_2320,N_24788,N_23063);
nand UO_2321 (O_2321,N_22803,N_23369);
nor UO_2322 (O_2322,N_24564,N_23655);
xnor UO_2323 (O_2323,N_24033,N_23502);
nor UO_2324 (O_2324,N_22582,N_22906);
nand UO_2325 (O_2325,N_23077,N_22588);
or UO_2326 (O_2326,N_24497,N_23056);
or UO_2327 (O_2327,N_23425,N_23353);
nor UO_2328 (O_2328,N_24629,N_23512);
nor UO_2329 (O_2329,N_23522,N_22578);
and UO_2330 (O_2330,N_24489,N_23895);
xor UO_2331 (O_2331,N_23480,N_23920);
nand UO_2332 (O_2332,N_23281,N_24314);
nor UO_2333 (O_2333,N_23722,N_22862);
or UO_2334 (O_2334,N_24412,N_23692);
or UO_2335 (O_2335,N_22896,N_23729);
or UO_2336 (O_2336,N_24432,N_22916);
and UO_2337 (O_2337,N_23540,N_24029);
nor UO_2338 (O_2338,N_23207,N_24689);
xor UO_2339 (O_2339,N_24643,N_22588);
or UO_2340 (O_2340,N_24294,N_24652);
nor UO_2341 (O_2341,N_23572,N_22550);
nor UO_2342 (O_2342,N_24778,N_22907);
or UO_2343 (O_2343,N_23589,N_24006);
nand UO_2344 (O_2344,N_24434,N_24646);
xor UO_2345 (O_2345,N_24840,N_22521);
and UO_2346 (O_2346,N_22569,N_22658);
nand UO_2347 (O_2347,N_24152,N_24432);
nand UO_2348 (O_2348,N_23396,N_22900);
xnor UO_2349 (O_2349,N_23009,N_23775);
and UO_2350 (O_2350,N_23996,N_22667);
xnor UO_2351 (O_2351,N_24023,N_23499);
or UO_2352 (O_2352,N_24841,N_24881);
xnor UO_2353 (O_2353,N_22746,N_24462);
and UO_2354 (O_2354,N_23445,N_23708);
or UO_2355 (O_2355,N_23803,N_23352);
and UO_2356 (O_2356,N_22616,N_22721);
nand UO_2357 (O_2357,N_23484,N_24357);
nand UO_2358 (O_2358,N_23964,N_23802);
or UO_2359 (O_2359,N_24539,N_22921);
nand UO_2360 (O_2360,N_24526,N_22779);
and UO_2361 (O_2361,N_24653,N_22978);
or UO_2362 (O_2362,N_23376,N_24290);
and UO_2363 (O_2363,N_23643,N_23831);
or UO_2364 (O_2364,N_23582,N_23255);
xor UO_2365 (O_2365,N_23128,N_23102);
and UO_2366 (O_2366,N_23920,N_24523);
or UO_2367 (O_2367,N_22671,N_23689);
nand UO_2368 (O_2368,N_23882,N_23274);
nor UO_2369 (O_2369,N_22568,N_23800);
xnor UO_2370 (O_2370,N_23804,N_24640);
or UO_2371 (O_2371,N_23217,N_23063);
and UO_2372 (O_2372,N_22700,N_24054);
nand UO_2373 (O_2373,N_24167,N_24184);
nand UO_2374 (O_2374,N_23972,N_24647);
and UO_2375 (O_2375,N_23299,N_23209);
nor UO_2376 (O_2376,N_23876,N_24109);
and UO_2377 (O_2377,N_24934,N_22666);
nand UO_2378 (O_2378,N_23895,N_24499);
or UO_2379 (O_2379,N_22507,N_23326);
xor UO_2380 (O_2380,N_23161,N_23426);
nand UO_2381 (O_2381,N_22719,N_24483);
or UO_2382 (O_2382,N_24417,N_24831);
or UO_2383 (O_2383,N_23987,N_22929);
and UO_2384 (O_2384,N_23782,N_24402);
nor UO_2385 (O_2385,N_22833,N_24565);
xnor UO_2386 (O_2386,N_23630,N_22548);
xnor UO_2387 (O_2387,N_23310,N_22545);
or UO_2388 (O_2388,N_22706,N_22536);
nand UO_2389 (O_2389,N_23239,N_24813);
nor UO_2390 (O_2390,N_23093,N_23415);
nor UO_2391 (O_2391,N_23772,N_23930);
and UO_2392 (O_2392,N_23844,N_24412);
xor UO_2393 (O_2393,N_23379,N_24376);
xnor UO_2394 (O_2394,N_23595,N_24435);
or UO_2395 (O_2395,N_24026,N_24956);
xnor UO_2396 (O_2396,N_23379,N_24540);
and UO_2397 (O_2397,N_24008,N_24980);
or UO_2398 (O_2398,N_24893,N_24466);
xnor UO_2399 (O_2399,N_23695,N_23223);
nand UO_2400 (O_2400,N_23227,N_23529);
xnor UO_2401 (O_2401,N_24581,N_24259);
or UO_2402 (O_2402,N_23276,N_23054);
or UO_2403 (O_2403,N_24094,N_24460);
and UO_2404 (O_2404,N_23613,N_23478);
and UO_2405 (O_2405,N_24470,N_24557);
nor UO_2406 (O_2406,N_24335,N_23462);
nand UO_2407 (O_2407,N_22571,N_22629);
xor UO_2408 (O_2408,N_24856,N_22667);
nor UO_2409 (O_2409,N_23366,N_24797);
or UO_2410 (O_2410,N_23064,N_23195);
or UO_2411 (O_2411,N_22609,N_24999);
and UO_2412 (O_2412,N_22694,N_24611);
nor UO_2413 (O_2413,N_23083,N_24099);
and UO_2414 (O_2414,N_24935,N_22542);
nand UO_2415 (O_2415,N_24784,N_24793);
and UO_2416 (O_2416,N_23224,N_24613);
nor UO_2417 (O_2417,N_22601,N_23257);
and UO_2418 (O_2418,N_23373,N_23176);
xor UO_2419 (O_2419,N_23285,N_23837);
nor UO_2420 (O_2420,N_23627,N_22562);
nand UO_2421 (O_2421,N_24079,N_23909);
and UO_2422 (O_2422,N_23816,N_24451);
or UO_2423 (O_2423,N_22506,N_22662);
or UO_2424 (O_2424,N_22789,N_24432);
and UO_2425 (O_2425,N_24095,N_22573);
nor UO_2426 (O_2426,N_22718,N_22911);
nor UO_2427 (O_2427,N_22737,N_23384);
or UO_2428 (O_2428,N_23813,N_24399);
and UO_2429 (O_2429,N_24211,N_24575);
or UO_2430 (O_2430,N_23136,N_23830);
or UO_2431 (O_2431,N_22784,N_23722);
and UO_2432 (O_2432,N_23530,N_22729);
xnor UO_2433 (O_2433,N_24396,N_22532);
xor UO_2434 (O_2434,N_22801,N_24162);
nor UO_2435 (O_2435,N_22968,N_23260);
nor UO_2436 (O_2436,N_22528,N_23917);
or UO_2437 (O_2437,N_22964,N_23533);
xnor UO_2438 (O_2438,N_22855,N_24188);
nor UO_2439 (O_2439,N_23251,N_23620);
xnor UO_2440 (O_2440,N_23309,N_23698);
nor UO_2441 (O_2441,N_24295,N_22542);
nand UO_2442 (O_2442,N_23365,N_23635);
nand UO_2443 (O_2443,N_24486,N_24156);
or UO_2444 (O_2444,N_24828,N_24719);
and UO_2445 (O_2445,N_24621,N_23858);
nor UO_2446 (O_2446,N_23057,N_23903);
nor UO_2447 (O_2447,N_24608,N_23598);
xor UO_2448 (O_2448,N_23925,N_22544);
nor UO_2449 (O_2449,N_23206,N_24653);
and UO_2450 (O_2450,N_24619,N_24113);
or UO_2451 (O_2451,N_24671,N_23991);
and UO_2452 (O_2452,N_24586,N_24619);
nor UO_2453 (O_2453,N_22798,N_24743);
xnor UO_2454 (O_2454,N_22761,N_23408);
nand UO_2455 (O_2455,N_24718,N_24315);
and UO_2456 (O_2456,N_22659,N_24408);
xnor UO_2457 (O_2457,N_23917,N_24075);
and UO_2458 (O_2458,N_24223,N_23582);
nand UO_2459 (O_2459,N_23235,N_23543);
nand UO_2460 (O_2460,N_22633,N_22914);
or UO_2461 (O_2461,N_22699,N_22638);
and UO_2462 (O_2462,N_24574,N_24079);
or UO_2463 (O_2463,N_22945,N_23540);
xnor UO_2464 (O_2464,N_22702,N_23708);
or UO_2465 (O_2465,N_24568,N_23289);
xnor UO_2466 (O_2466,N_23891,N_24725);
nand UO_2467 (O_2467,N_24796,N_23173);
nand UO_2468 (O_2468,N_23623,N_24710);
and UO_2469 (O_2469,N_24986,N_22895);
nand UO_2470 (O_2470,N_22842,N_23662);
nand UO_2471 (O_2471,N_23241,N_24351);
nand UO_2472 (O_2472,N_23867,N_24785);
nand UO_2473 (O_2473,N_23182,N_23412);
xor UO_2474 (O_2474,N_23744,N_23204);
or UO_2475 (O_2475,N_24841,N_23802);
or UO_2476 (O_2476,N_23698,N_24191);
and UO_2477 (O_2477,N_24243,N_22508);
or UO_2478 (O_2478,N_24065,N_24283);
or UO_2479 (O_2479,N_24626,N_23113);
nand UO_2480 (O_2480,N_24827,N_23691);
or UO_2481 (O_2481,N_24755,N_23183);
nand UO_2482 (O_2482,N_23497,N_23982);
or UO_2483 (O_2483,N_24060,N_22713);
nor UO_2484 (O_2484,N_24622,N_23237);
nor UO_2485 (O_2485,N_23892,N_23201);
xor UO_2486 (O_2486,N_22787,N_24822);
nand UO_2487 (O_2487,N_22887,N_22833);
nor UO_2488 (O_2488,N_23871,N_23117);
and UO_2489 (O_2489,N_23232,N_24692);
nor UO_2490 (O_2490,N_23107,N_22616);
nor UO_2491 (O_2491,N_23026,N_22652);
or UO_2492 (O_2492,N_23138,N_23471);
nor UO_2493 (O_2493,N_22699,N_24129);
and UO_2494 (O_2494,N_23051,N_24916);
nor UO_2495 (O_2495,N_24994,N_24052);
nor UO_2496 (O_2496,N_22688,N_23415);
nand UO_2497 (O_2497,N_24359,N_23753);
nand UO_2498 (O_2498,N_24261,N_22526);
nand UO_2499 (O_2499,N_23596,N_23840);
or UO_2500 (O_2500,N_23375,N_22886);
nand UO_2501 (O_2501,N_24508,N_23263);
xor UO_2502 (O_2502,N_22552,N_23517);
xor UO_2503 (O_2503,N_24670,N_23883);
and UO_2504 (O_2504,N_23923,N_24610);
xor UO_2505 (O_2505,N_24638,N_24879);
xor UO_2506 (O_2506,N_24820,N_24304);
and UO_2507 (O_2507,N_22988,N_23186);
nand UO_2508 (O_2508,N_23084,N_24595);
nand UO_2509 (O_2509,N_23353,N_24416);
nand UO_2510 (O_2510,N_23805,N_23368);
xor UO_2511 (O_2511,N_22579,N_23515);
nand UO_2512 (O_2512,N_24312,N_24682);
and UO_2513 (O_2513,N_23329,N_24631);
or UO_2514 (O_2514,N_23163,N_23073);
nand UO_2515 (O_2515,N_22767,N_24184);
xor UO_2516 (O_2516,N_23444,N_24300);
nand UO_2517 (O_2517,N_24587,N_23138);
or UO_2518 (O_2518,N_24149,N_22637);
or UO_2519 (O_2519,N_24652,N_22954);
nor UO_2520 (O_2520,N_22563,N_23654);
nand UO_2521 (O_2521,N_24074,N_23598);
and UO_2522 (O_2522,N_23790,N_24296);
xnor UO_2523 (O_2523,N_24528,N_23870);
or UO_2524 (O_2524,N_24705,N_24156);
nand UO_2525 (O_2525,N_23076,N_23522);
xnor UO_2526 (O_2526,N_23328,N_23539);
nand UO_2527 (O_2527,N_23298,N_22814);
or UO_2528 (O_2528,N_23017,N_24362);
nor UO_2529 (O_2529,N_23433,N_22850);
nand UO_2530 (O_2530,N_24784,N_22823);
and UO_2531 (O_2531,N_24134,N_22611);
xnor UO_2532 (O_2532,N_24228,N_24670);
nor UO_2533 (O_2533,N_24661,N_23414);
nand UO_2534 (O_2534,N_24390,N_23055);
xnor UO_2535 (O_2535,N_24231,N_22917);
xor UO_2536 (O_2536,N_23760,N_23400);
and UO_2537 (O_2537,N_22853,N_22708);
xor UO_2538 (O_2538,N_22610,N_23741);
and UO_2539 (O_2539,N_24404,N_24816);
nor UO_2540 (O_2540,N_24399,N_22987);
nor UO_2541 (O_2541,N_24341,N_24292);
xnor UO_2542 (O_2542,N_23407,N_24556);
xor UO_2543 (O_2543,N_23814,N_24445);
xor UO_2544 (O_2544,N_22506,N_23102);
xnor UO_2545 (O_2545,N_24866,N_24978);
nand UO_2546 (O_2546,N_23856,N_22562);
nor UO_2547 (O_2547,N_23348,N_23373);
nand UO_2548 (O_2548,N_24391,N_23718);
nor UO_2549 (O_2549,N_24504,N_23033);
nand UO_2550 (O_2550,N_23136,N_24467);
nand UO_2551 (O_2551,N_22984,N_24277);
and UO_2552 (O_2552,N_23124,N_24543);
nand UO_2553 (O_2553,N_23445,N_23179);
or UO_2554 (O_2554,N_23991,N_22827);
nor UO_2555 (O_2555,N_24389,N_23671);
and UO_2556 (O_2556,N_23019,N_23110);
nor UO_2557 (O_2557,N_24726,N_24689);
xor UO_2558 (O_2558,N_23957,N_22705);
or UO_2559 (O_2559,N_23941,N_23444);
nand UO_2560 (O_2560,N_23350,N_22792);
xor UO_2561 (O_2561,N_24257,N_24857);
or UO_2562 (O_2562,N_24205,N_22991);
xor UO_2563 (O_2563,N_23483,N_23756);
or UO_2564 (O_2564,N_23006,N_23870);
or UO_2565 (O_2565,N_22787,N_24297);
nand UO_2566 (O_2566,N_23578,N_22909);
or UO_2567 (O_2567,N_24829,N_24016);
and UO_2568 (O_2568,N_24161,N_24609);
nand UO_2569 (O_2569,N_24418,N_24764);
xor UO_2570 (O_2570,N_23837,N_24124);
nor UO_2571 (O_2571,N_22721,N_24035);
xnor UO_2572 (O_2572,N_22693,N_23033);
nand UO_2573 (O_2573,N_23833,N_22973);
xnor UO_2574 (O_2574,N_23683,N_24938);
nand UO_2575 (O_2575,N_22642,N_22838);
nor UO_2576 (O_2576,N_22652,N_23910);
and UO_2577 (O_2577,N_24482,N_23779);
nand UO_2578 (O_2578,N_24970,N_24745);
nor UO_2579 (O_2579,N_23169,N_22756);
or UO_2580 (O_2580,N_24480,N_24115);
or UO_2581 (O_2581,N_24025,N_24975);
and UO_2582 (O_2582,N_23287,N_22714);
xnor UO_2583 (O_2583,N_24898,N_24011);
xor UO_2584 (O_2584,N_23445,N_23494);
and UO_2585 (O_2585,N_23319,N_23250);
or UO_2586 (O_2586,N_23977,N_23539);
nand UO_2587 (O_2587,N_23737,N_23798);
nand UO_2588 (O_2588,N_22899,N_23916);
and UO_2589 (O_2589,N_24806,N_22546);
nand UO_2590 (O_2590,N_23280,N_24536);
nand UO_2591 (O_2591,N_22846,N_22718);
nand UO_2592 (O_2592,N_23070,N_22885);
or UO_2593 (O_2593,N_22662,N_23069);
nor UO_2594 (O_2594,N_23895,N_23821);
xnor UO_2595 (O_2595,N_23947,N_23441);
nor UO_2596 (O_2596,N_24660,N_23151);
nor UO_2597 (O_2597,N_24460,N_23077);
nand UO_2598 (O_2598,N_24728,N_22579);
xor UO_2599 (O_2599,N_24439,N_23661);
and UO_2600 (O_2600,N_24093,N_24407);
and UO_2601 (O_2601,N_23183,N_23339);
and UO_2602 (O_2602,N_23425,N_23867);
or UO_2603 (O_2603,N_24490,N_24236);
or UO_2604 (O_2604,N_22627,N_24720);
nand UO_2605 (O_2605,N_22995,N_24844);
nand UO_2606 (O_2606,N_23843,N_24125);
nand UO_2607 (O_2607,N_24639,N_24775);
and UO_2608 (O_2608,N_23453,N_22973);
nor UO_2609 (O_2609,N_24811,N_24720);
xnor UO_2610 (O_2610,N_23436,N_23264);
nand UO_2611 (O_2611,N_23841,N_23094);
and UO_2612 (O_2612,N_24492,N_23013);
and UO_2613 (O_2613,N_23700,N_22593);
or UO_2614 (O_2614,N_22955,N_24806);
nand UO_2615 (O_2615,N_22756,N_24174);
nor UO_2616 (O_2616,N_23356,N_23347);
or UO_2617 (O_2617,N_23363,N_23148);
or UO_2618 (O_2618,N_22842,N_24144);
xor UO_2619 (O_2619,N_22985,N_24483);
and UO_2620 (O_2620,N_23250,N_24186);
or UO_2621 (O_2621,N_23993,N_22828);
nor UO_2622 (O_2622,N_23659,N_24877);
or UO_2623 (O_2623,N_23899,N_23312);
xor UO_2624 (O_2624,N_24118,N_23630);
or UO_2625 (O_2625,N_24572,N_24881);
or UO_2626 (O_2626,N_24544,N_22801);
xor UO_2627 (O_2627,N_22734,N_24233);
nor UO_2628 (O_2628,N_23952,N_24672);
xor UO_2629 (O_2629,N_24876,N_23954);
xor UO_2630 (O_2630,N_23598,N_24491);
or UO_2631 (O_2631,N_23543,N_23900);
and UO_2632 (O_2632,N_23879,N_22900);
nor UO_2633 (O_2633,N_24094,N_24395);
xnor UO_2634 (O_2634,N_24737,N_23530);
or UO_2635 (O_2635,N_24450,N_24839);
or UO_2636 (O_2636,N_22788,N_24037);
nor UO_2637 (O_2637,N_24199,N_23106);
and UO_2638 (O_2638,N_22855,N_22630);
xnor UO_2639 (O_2639,N_24519,N_23627);
nor UO_2640 (O_2640,N_24826,N_24315);
or UO_2641 (O_2641,N_24634,N_23991);
or UO_2642 (O_2642,N_23562,N_24172);
and UO_2643 (O_2643,N_24858,N_24301);
and UO_2644 (O_2644,N_22732,N_24848);
nand UO_2645 (O_2645,N_24677,N_22558);
or UO_2646 (O_2646,N_22596,N_24226);
nand UO_2647 (O_2647,N_24802,N_23224);
nor UO_2648 (O_2648,N_23827,N_23721);
nor UO_2649 (O_2649,N_24644,N_24423);
nand UO_2650 (O_2650,N_24728,N_24181);
xor UO_2651 (O_2651,N_23357,N_24258);
nand UO_2652 (O_2652,N_23149,N_23088);
nor UO_2653 (O_2653,N_23333,N_22989);
nand UO_2654 (O_2654,N_24912,N_24104);
or UO_2655 (O_2655,N_23219,N_22688);
xor UO_2656 (O_2656,N_22722,N_23744);
xnor UO_2657 (O_2657,N_22754,N_24660);
nor UO_2658 (O_2658,N_24174,N_23422);
or UO_2659 (O_2659,N_24269,N_22764);
or UO_2660 (O_2660,N_23445,N_24298);
xnor UO_2661 (O_2661,N_23828,N_23922);
or UO_2662 (O_2662,N_24264,N_22978);
and UO_2663 (O_2663,N_22865,N_23525);
nor UO_2664 (O_2664,N_23463,N_24999);
xnor UO_2665 (O_2665,N_22841,N_24057);
and UO_2666 (O_2666,N_22840,N_22632);
nor UO_2667 (O_2667,N_24904,N_23769);
nor UO_2668 (O_2668,N_24013,N_24305);
xnor UO_2669 (O_2669,N_22545,N_24061);
or UO_2670 (O_2670,N_24073,N_22801);
or UO_2671 (O_2671,N_24407,N_23018);
nor UO_2672 (O_2672,N_24274,N_24453);
and UO_2673 (O_2673,N_24740,N_24817);
xnor UO_2674 (O_2674,N_24994,N_24422);
nand UO_2675 (O_2675,N_23731,N_23399);
nand UO_2676 (O_2676,N_24294,N_24248);
xnor UO_2677 (O_2677,N_23657,N_23120);
and UO_2678 (O_2678,N_23352,N_23754);
nor UO_2679 (O_2679,N_23948,N_23237);
or UO_2680 (O_2680,N_22714,N_24226);
xor UO_2681 (O_2681,N_23975,N_24249);
nand UO_2682 (O_2682,N_23212,N_23757);
xnor UO_2683 (O_2683,N_23327,N_23199);
or UO_2684 (O_2684,N_23763,N_24331);
nand UO_2685 (O_2685,N_23175,N_24451);
nor UO_2686 (O_2686,N_23678,N_22681);
nand UO_2687 (O_2687,N_22716,N_24285);
and UO_2688 (O_2688,N_22767,N_23020);
nand UO_2689 (O_2689,N_24636,N_23336);
and UO_2690 (O_2690,N_23596,N_23587);
nand UO_2691 (O_2691,N_24574,N_24643);
nand UO_2692 (O_2692,N_24767,N_23275);
or UO_2693 (O_2693,N_23886,N_22550);
xnor UO_2694 (O_2694,N_23936,N_23803);
nor UO_2695 (O_2695,N_23498,N_23535);
xnor UO_2696 (O_2696,N_22573,N_22818);
and UO_2697 (O_2697,N_23678,N_23182);
nor UO_2698 (O_2698,N_22938,N_24385);
nand UO_2699 (O_2699,N_22742,N_24238);
nor UO_2700 (O_2700,N_24520,N_23490);
and UO_2701 (O_2701,N_24296,N_23912);
xnor UO_2702 (O_2702,N_24636,N_23043);
and UO_2703 (O_2703,N_22622,N_22757);
or UO_2704 (O_2704,N_22865,N_24693);
or UO_2705 (O_2705,N_23104,N_23312);
xnor UO_2706 (O_2706,N_22938,N_24395);
and UO_2707 (O_2707,N_24721,N_24146);
nor UO_2708 (O_2708,N_24189,N_23758);
and UO_2709 (O_2709,N_23585,N_22787);
xor UO_2710 (O_2710,N_24197,N_23366);
xnor UO_2711 (O_2711,N_22784,N_24564);
and UO_2712 (O_2712,N_22574,N_24975);
xnor UO_2713 (O_2713,N_23782,N_22952);
nor UO_2714 (O_2714,N_24537,N_22958);
or UO_2715 (O_2715,N_23496,N_22637);
nand UO_2716 (O_2716,N_22839,N_22954);
nand UO_2717 (O_2717,N_24959,N_22693);
nand UO_2718 (O_2718,N_23950,N_23535);
nor UO_2719 (O_2719,N_22641,N_24111);
xor UO_2720 (O_2720,N_23360,N_24662);
xnor UO_2721 (O_2721,N_23682,N_24590);
nor UO_2722 (O_2722,N_23828,N_22756);
nand UO_2723 (O_2723,N_22830,N_23417);
nor UO_2724 (O_2724,N_24595,N_23837);
nor UO_2725 (O_2725,N_24779,N_23690);
or UO_2726 (O_2726,N_24074,N_24929);
nor UO_2727 (O_2727,N_24682,N_23688);
xnor UO_2728 (O_2728,N_24321,N_24119);
xnor UO_2729 (O_2729,N_24637,N_24311);
xor UO_2730 (O_2730,N_23526,N_22611);
or UO_2731 (O_2731,N_24346,N_23179);
nand UO_2732 (O_2732,N_23245,N_22927);
or UO_2733 (O_2733,N_23031,N_22834);
nand UO_2734 (O_2734,N_24741,N_24450);
or UO_2735 (O_2735,N_23282,N_24335);
or UO_2736 (O_2736,N_23390,N_22956);
nand UO_2737 (O_2737,N_24647,N_23608);
nand UO_2738 (O_2738,N_24496,N_24252);
nand UO_2739 (O_2739,N_24862,N_24185);
nand UO_2740 (O_2740,N_23371,N_23001);
and UO_2741 (O_2741,N_24140,N_24978);
and UO_2742 (O_2742,N_22822,N_23927);
or UO_2743 (O_2743,N_24798,N_23280);
nor UO_2744 (O_2744,N_24959,N_23767);
nor UO_2745 (O_2745,N_24667,N_24095);
xor UO_2746 (O_2746,N_24718,N_24944);
nand UO_2747 (O_2747,N_22713,N_22725);
nor UO_2748 (O_2748,N_24051,N_22989);
or UO_2749 (O_2749,N_22996,N_24811);
nand UO_2750 (O_2750,N_24713,N_24985);
xnor UO_2751 (O_2751,N_23533,N_24848);
nor UO_2752 (O_2752,N_23877,N_24130);
xnor UO_2753 (O_2753,N_23093,N_24817);
nor UO_2754 (O_2754,N_23252,N_22777);
or UO_2755 (O_2755,N_24752,N_24686);
xnor UO_2756 (O_2756,N_23820,N_24589);
nor UO_2757 (O_2757,N_23348,N_24233);
nand UO_2758 (O_2758,N_24933,N_23424);
or UO_2759 (O_2759,N_24587,N_24206);
xor UO_2760 (O_2760,N_24190,N_24185);
or UO_2761 (O_2761,N_23844,N_24162);
xor UO_2762 (O_2762,N_24717,N_23222);
xor UO_2763 (O_2763,N_24243,N_22502);
nor UO_2764 (O_2764,N_24101,N_23103);
or UO_2765 (O_2765,N_23043,N_23522);
and UO_2766 (O_2766,N_22605,N_23247);
nor UO_2767 (O_2767,N_23539,N_23118);
or UO_2768 (O_2768,N_24219,N_22594);
nor UO_2769 (O_2769,N_24114,N_24600);
or UO_2770 (O_2770,N_23443,N_23676);
and UO_2771 (O_2771,N_24501,N_23114);
xor UO_2772 (O_2772,N_22703,N_24209);
nand UO_2773 (O_2773,N_23727,N_24677);
nand UO_2774 (O_2774,N_24906,N_24968);
nand UO_2775 (O_2775,N_23514,N_22621);
nand UO_2776 (O_2776,N_22804,N_24747);
nand UO_2777 (O_2777,N_23901,N_24701);
xor UO_2778 (O_2778,N_23018,N_24166);
nor UO_2779 (O_2779,N_23099,N_22631);
xor UO_2780 (O_2780,N_23711,N_24806);
and UO_2781 (O_2781,N_23811,N_22647);
and UO_2782 (O_2782,N_23647,N_24201);
nor UO_2783 (O_2783,N_24838,N_24819);
and UO_2784 (O_2784,N_22605,N_23101);
or UO_2785 (O_2785,N_24507,N_23533);
and UO_2786 (O_2786,N_23153,N_24514);
or UO_2787 (O_2787,N_24864,N_24225);
xor UO_2788 (O_2788,N_23030,N_23878);
and UO_2789 (O_2789,N_24911,N_24424);
xor UO_2790 (O_2790,N_24404,N_24151);
nor UO_2791 (O_2791,N_23809,N_24678);
and UO_2792 (O_2792,N_24422,N_24012);
nand UO_2793 (O_2793,N_23518,N_24030);
and UO_2794 (O_2794,N_24005,N_23674);
nor UO_2795 (O_2795,N_22909,N_22831);
nand UO_2796 (O_2796,N_23471,N_24874);
nand UO_2797 (O_2797,N_23677,N_24581);
nand UO_2798 (O_2798,N_23846,N_23665);
or UO_2799 (O_2799,N_24406,N_23727);
nand UO_2800 (O_2800,N_23172,N_22592);
xor UO_2801 (O_2801,N_22610,N_23559);
xnor UO_2802 (O_2802,N_23898,N_24228);
nand UO_2803 (O_2803,N_23165,N_23563);
nand UO_2804 (O_2804,N_23538,N_23595);
and UO_2805 (O_2805,N_23166,N_23896);
nand UO_2806 (O_2806,N_23168,N_24558);
xnor UO_2807 (O_2807,N_24299,N_22793);
xnor UO_2808 (O_2808,N_22598,N_22932);
xor UO_2809 (O_2809,N_23799,N_24035);
nand UO_2810 (O_2810,N_22560,N_24938);
or UO_2811 (O_2811,N_24641,N_24405);
nand UO_2812 (O_2812,N_24168,N_24826);
xnor UO_2813 (O_2813,N_24877,N_24651);
nor UO_2814 (O_2814,N_23229,N_24316);
and UO_2815 (O_2815,N_24621,N_24142);
nand UO_2816 (O_2816,N_22810,N_23535);
nor UO_2817 (O_2817,N_22990,N_23715);
and UO_2818 (O_2818,N_23255,N_24906);
or UO_2819 (O_2819,N_23232,N_23022);
and UO_2820 (O_2820,N_22594,N_24709);
nor UO_2821 (O_2821,N_23500,N_22783);
and UO_2822 (O_2822,N_23081,N_24021);
xor UO_2823 (O_2823,N_24680,N_24086);
or UO_2824 (O_2824,N_24738,N_24841);
and UO_2825 (O_2825,N_23018,N_24063);
and UO_2826 (O_2826,N_23394,N_24178);
nor UO_2827 (O_2827,N_24213,N_23013);
or UO_2828 (O_2828,N_23890,N_24535);
nor UO_2829 (O_2829,N_23841,N_23157);
nor UO_2830 (O_2830,N_23479,N_22768);
nand UO_2831 (O_2831,N_23276,N_23076);
nor UO_2832 (O_2832,N_23419,N_24819);
or UO_2833 (O_2833,N_24087,N_22896);
xnor UO_2834 (O_2834,N_23151,N_23865);
or UO_2835 (O_2835,N_24668,N_23766);
or UO_2836 (O_2836,N_24114,N_24301);
xnor UO_2837 (O_2837,N_24531,N_23670);
and UO_2838 (O_2838,N_23624,N_22603);
and UO_2839 (O_2839,N_22690,N_24070);
nor UO_2840 (O_2840,N_24817,N_23016);
nor UO_2841 (O_2841,N_24092,N_23969);
or UO_2842 (O_2842,N_24498,N_22770);
xor UO_2843 (O_2843,N_22989,N_24668);
nor UO_2844 (O_2844,N_24594,N_22854);
or UO_2845 (O_2845,N_23359,N_24333);
or UO_2846 (O_2846,N_23290,N_23497);
and UO_2847 (O_2847,N_24535,N_24556);
or UO_2848 (O_2848,N_23348,N_24083);
nand UO_2849 (O_2849,N_24993,N_24165);
xnor UO_2850 (O_2850,N_23580,N_23715);
and UO_2851 (O_2851,N_22854,N_24045);
nand UO_2852 (O_2852,N_22626,N_24303);
or UO_2853 (O_2853,N_24515,N_23100);
and UO_2854 (O_2854,N_24733,N_24102);
or UO_2855 (O_2855,N_23340,N_22863);
and UO_2856 (O_2856,N_24849,N_24113);
xor UO_2857 (O_2857,N_22853,N_22768);
nand UO_2858 (O_2858,N_23439,N_22582);
nand UO_2859 (O_2859,N_23629,N_23502);
and UO_2860 (O_2860,N_22500,N_23988);
and UO_2861 (O_2861,N_23489,N_23442);
nand UO_2862 (O_2862,N_22688,N_24401);
or UO_2863 (O_2863,N_24277,N_23383);
and UO_2864 (O_2864,N_22559,N_24746);
or UO_2865 (O_2865,N_22609,N_23359);
nand UO_2866 (O_2866,N_23545,N_22801);
xnor UO_2867 (O_2867,N_24148,N_24488);
nor UO_2868 (O_2868,N_24827,N_24642);
xor UO_2869 (O_2869,N_23749,N_23440);
nor UO_2870 (O_2870,N_24518,N_23515);
nand UO_2871 (O_2871,N_23025,N_23973);
and UO_2872 (O_2872,N_24739,N_24782);
xor UO_2873 (O_2873,N_24724,N_24955);
nand UO_2874 (O_2874,N_24264,N_23955);
xnor UO_2875 (O_2875,N_24279,N_24668);
or UO_2876 (O_2876,N_23409,N_23182);
nand UO_2877 (O_2877,N_24520,N_23780);
or UO_2878 (O_2878,N_22624,N_24665);
xnor UO_2879 (O_2879,N_22697,N_22896);
or UO_2880 (O_2880,N_24460,N_22511);
nand UO_2881 (O_2881,N_24481,N_24126);
or UO_2882 (O_2882,N_24333,N_24056);
and UO_2883 (O_2883,N_23018,N_24994);
and UO_2884 (O_2884,N_22987,N_24527);
and UO_2885 (O_2885,N_23450,N_23068);
nand UO_2886 (O_2886,N_22849,N_22962);
nor UO_2887 (O_2887,N_23225,N_24336);
and UO_2888 (O_2888,N_22832,N_23060);
nor UO_2889 (O_2889,N_23996,N_22599);
nor UO_2890 (O_2890,N_24963,N_23409);
nor UO_2891 (O_2891,N_22781,N_23610);
and UO_2892 (O_2892,N_22618,N_22974);
nand UO_2893 (O_2893,N_22625,N_23014);
or UO_2894 (O_2894,N_24609,N_23972);
or UO_2895 (O_2895,N_23100,N_22507);
nor UO_2896 (O_2896,N_24022,N_24037);
nor UO_2897 (O_2897,N_23473,N_22993);
nand UO_2898 (O_2898,N_23947,N_24811);
nor UO_2899 (O_2899,N_24485,N_22532);
and UO_2900 (O_2900,N_23562,N_23540);
or UO_2901 (O_2901,N_24735,N_24548);
and UO_2902 (O_2902,N_23119,N_24407);
nand UO_2903 (O_2903,N_24234,N_24291);
nand UO_2904 (O_2904,N_24064,N_24961);
nand UO_2905 (O_2905,N_24384,N_24374);
and UO_2906 (O_2906,N_23906,N_24579);
nand UO_2907 (O_2907,N_24919,N_23708);
and UO_2908 (O_2908,N_22853,N_24877);
and UO_2909 (O_2909,N_24906,N_24077);
nand UO_2910 (O_2910,N_23021,N_23785);
nand UO_2911 (O_2911,N_24296,N_22886);
nand UO_2912 (O_2912,N_24278,N_23187);
nand UO_2913 (O_2913,N_23530,N_24887);
xor UO_2914 (O_2914,N_23204,N_23338);
or UO_2915 (O_2915,N_24084,N_23136);
and UO_2916 (O_2916,N_22967,N_23861);
or UO_2917 (O_2917,N_23552,N_23402);
or UO_2918 (O_2918,N_23177,N_23563);
nand UO_2919 (O_2919,N_23276,N_24449);
or UO_2920 (O_2920,N_23977,N_22864);
or UO_2921 (O_2921,N_22821,N_24747);
nand UO_2922 (O_2922,N_24077,N_24812);
and UO_2923 (O_2923,N_24950,N_23237);
xor UO_2924 (O_2924,N_24222,N_22546);
and UO_2925 (O_2925,N_23113,N_23296);
nand UO_2926 (O_2926,N_22804,N_23487);
nor UO_2927 (O_2927,N_24877,N_23824);
nand UO_2928 (O_2928,N_23616,N_24838);
xor UO_2929 (O_2929,N_24736,N_22559);
and UO_2930 (O_2930,N_22767,N_23187);
and UO_2931 (O_2931,N_24740,N_22538);
and UO_2932 (O_2932,N_23374,N_23123);
or UO_2933 (O_2933,N_22628,N_23441);
nand UO_2934 (O_2934,N_23061,N_24775);
xor UO_2935 (O_2935,N_23706,N_24884);
xor UO_2936 (O_2936,N_23809,N_23068);
xnor UO_2937 (O_2937,N_22518,N_24490);
or UO_2938 (O_2938,N_22551,N_23802);
and UO_2939 (O_2939,N_23466,N_24567);
xnor UO_2940 (O_2940,N_24960,N_24345);
nand UO_2941 (O_2941,N_22717,N_24988);
xor UO_2942 (O_2942,N_22864,N_24631);
nor UO_2943 (O_2943,N_24624,N_22530);
and UO_2944 (O_2944,N_23371,N_24879);
nor UO_2945 (O_2945,N_23001,N_22587);
nand UO_2946 (O_2946,N_23246,N_24570);
nor UO_2947 (O_2947,N_22674,N_24785);
xor UO_2948 (O_2948,N_23429,N_24068);
xnor UO_2949 (O_2949,N_24972,N_22704);
nor UO_2950 (O_2950,N_22799,N_23454);
xnor UO_2951 (O_2951,N_24498,N_23618);
nand UO_2952 (O_2952,N_23961,N_23298);
xor UO_2953 (O_2953,N_24150,N_24443);
nand UO_2954 (O_2954,N_23675,N_24494);
nor UO_2955 (O_2955,N_24854,N_24702);
nand UO_2956 (O_2956,N_22949,N_23636);
nor UO_2957 (O_2957,N_24609,N_24408);
nand UO_2958 (O_2958,N_24307,N_22786);
nor UO_2959 (O_2959,N_23907,N_24659);
nor UO_2960 (O_2960,N_23747,N_24656);
nor UO_2961 (O_2961,N_24767,N_24604);
nor UO_2962 (O_2962,N_22876,N_24149);
and UO_2963 (O_2963,N_22629,N_24706);
xnor UO_2964 (O_2964,N_23952,N_22915);
nand UO_2965 (O_2965,N_24481,N_24537);
xor UO_2966 (O_2966,N_24495,N_23305);
xnor UO_2967 (O_2967,N_23325,N_24783);
nor UO_2968 (O_2968,N_23389,N_22953);
nor UO_2969 (O_2969,N_23112,N_24249);
nand UO_2970 (O_2970,N_23400,N_22610);
nor UO_2971 (O_2971,N_24756,N_24790);
or UO_2972 (O_2972,N_22742,N_24304);
or UO_2973 (O_2973,N_22610,N_23587);
nor UO_2974 (O_2974,N_24376,N_23562);
nor UO_2975 (O_2975,N_24160,N_24101);
nand UO_2976 (O_2976,N_23649,N_24144);
xor UO_2977 (O_2977,N_23919,N_23431);
xor UO_2978 (O_2978,N_23976,N_22787);
or UO_2979 (O_2979,N_22520,N_23960);
or UO_2980 (O_2980,N_24340,N_24362);
and UO_2981 (O_2981,N_24667,N_24216);
or UO_2982 (O_2982,N_23944,N_23761);
xnor UO_2983 (O_2983,N_24030,N_22643);
or UO_2984 (O_2984,N_24222,N_22863);
and UO_2985 (O_2985,N_24543,N_22688);
or UO_2986 (O_2986,N_22738,N_23597);
or UO_2987 (O_2987,N_24540,N_23768);
nor UO_2988 (O_2988,N_24414,N_22587);
or UO_2989 (O_2989,N_22519,N_23446);
nand UO_2990 (O_2990,N_23023,N_22851);
and UO_2991 (O_2991,N_22766,N_23543);
and UO_2992 (O_2992,N_24024,N_23437);
and UO_2993 (O_2993,N_22714,N_24638);
nor UO_2994 (O_2994,N_23167,N_23307);
and UO_2995 (O_2995,N_24209,N_23227);
nor UO_2996 (O_2996,N_23275,N_24322);
xor UO_2997 (O_2997,N_22720,N_23681);
nand UO_2998 (O_2998,N_22596,N_22563);
nand UO_2999 (O_2999,N_23770,N_24735);
endmodule