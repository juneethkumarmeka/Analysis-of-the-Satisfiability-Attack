module basic_1500_15000_2000_30_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1358,In_158);
xor U1 (N_1,In_1213,In_592);
or U2 (N_2,In_564,In_1490);
nor U3 (N_3,In_576,In_555);
nor U4 (N_4,In_1172,In_1120);
or U5 (N_5,In_1248,In_957);
nand U6 (N_6,In_385,In_1168);
nand U7 (N_7,In_1133,In_228);
xnor U8 (N_8,In_1206,In_207);
nor U9 (N_9,In_1016,In_5);
nand U10 (N_10,In_302,In_110);
and U11 (N_11,In_1029,In_753);
nor U12 (N_12,In_279,In_674);
and U13 (N_13,In_1318,In_618);
and U14 (N_14,In_244,In_1410);
nor U15 (N_15,In_819,In_1121);
or U16 (N_16,In_536,In_870);
or U17 (N_17,In_141,In_583);
or U18 (N_18,In_632,In_152);
nand U19 (N_19,In_30,In_976);
nand U20 (N_20,In_1209,In_1063);
or U21 (N_21,In_645,In_788);
and U22 (N_22,In_86,In_613);
nand U23 (N_23,In_1239,In_972);
xor U24 (N_24,In_122,In_1230);
and U25 (N_25,In_792,In_915);
nor U26 (N_26,In_802,In_81);
and U27 (N_27,In_1424,In_1295);
nor U28 (N_28,In_474,In_1357);
nand U29 (N_29,In_1182,In_66);
nand U30 (N_30,In_1186,In_1200);
nand U31 (N_31,In_734,In_1233);
nand U32 (N_32,In_960,In_318);
nor U33 (N_33,In_305,In_378);
nor U34 (N_34,In_1210,In_360);
or U35 (N_35,In_1151,In_439);
nand U36 (N_36,In_1044,In_1095);
and U37 (N_37,In_420,In_376);
nor U38 (N_38,In_1045,In_804);
and U39 (N_39,In_1485,In_742);
nor U40 (N_40,In_1379,In_824);
xnor U41 (N_41,In_400,In_186);
nor U42 (N_42,In_896,In_574);
or U43 (N_43,In_172,In_151);
nor U44 (N_44,In_402,In_954);
and U45 (N_45,In_1269,In_994);
nor U46 (N_46,In_337,In_398);
or U47 (N_47,In_1264,In_1378);
or U48 (N_48,In_774,In_356);
and U49 (N_49,In_1388,In_1347);
xnor U50 (N_50,In_869,In_68);
nor U51 (N_51,In_1166,In_98);
nand U52 (N_52,In_547,In_161);
nor U53 (N_53,In_473,In_1080);
nor U54 (N_54,In_46,In_1475);
nor U55 (N_55,In_35,In_812);
nand U56 (N_56,In_1272,In_1008);
nand U57 (N_57,In_362,In_1089);
xnor U58 (N_58,In_897,In_380);
and U59 (N_59,In_893,In_1196);
or U60 (N_60,In_894,In_531);
nand U61 (N_61,In_1279,In_73);
and U62 (N_62,In_1428,In_488);
or U63 (N_63,In_1390,In_1283);
or U64 (N_64,In_233,In_649);
xor U65 (N_65,In_1250,In_1115);
xor U66 (N_66,In_1051,In_1418);
nor U67 (N_67,In_1065,In_231);
or U68 (N_68,In_1436,In_200);
nand U69 (N_69,In_715,In_1132);
or U70 (N_70,In_1241,In_225);
nor U71 (N_71,In_1340,In_783);
nor U72 (N_72,In_740,In_1282);
xnor U73 (N_73,In_1001,In_1111);
xnor U74 (N_74,In_220,In_1060);
or U75 (N_75,In_1126,In_1040);
and U76 (N_76,In_955,In_164);
nand U77 (N_77,In_549,In_1078);
xnor U78 (N_78,In_963,In_218);
and U79 (N_79,In_993,In_1258);
or U80 (N_80,In_0,In_44);
xnor U81 (N_81,In_1434,In_1136);
and U82 (N_82,In_977,In_210);
nor U83 (N_83,In_193,In_899);
or U84 (N_84,In_1232,In_138);
nor U85 (N_85,In_258,In_588);
nand U86 (N_86,In_806,In_47);
xor U87 (N_87,In_521,In_304);
nor U88 (N_88,In_1130,In_340);
xor U89 (N_89,In_744,In_1161);
or U90 (N_90,In_842,In_898);
and U91 (N_91,In_939,In_985);
xnor U92 (N_92,In_884,In_1299);
nor U93 (N_93,In_1467,In_1408);
and U94 (N_94,In_289,In_619);
and U95 (N_95,In_837,In_442);
and U96 (N_96,In_568,In_518);
nor U97 (N_97,In_1013,In_91);
xor U98 (N_98,In_701,In_598);
xnor U99 (N_99,In_758,In_390);
nand U100 (N_100,In_121,In_187);
or U101 (N_101,In_1298,In_1105);
and U102 (N_102,In_1356,In_617);
nor U103 (N_103,In_1302,In_650);
nor U104 (N_104,In_638,In_154);
nand U105 (N_105,In_299,In_907);
nand U106 (N_106,In_106,In_309);
nand U107 (N_107,In_779,In_345);
and U108 (N_108,In_206,In_404);
nor U109 (N_109,In_24,In_428);
and U110 (N_110,In_1039,In_1135);
nor U111 (N_111,In_382,In_543);
and U112 (N_112,In_780,In_996);
nor U113 (N_113,In_216,In_155);
nor U114 (N_114,In_560,In_448);
xnor U115 (N_115,In_59,In_1253);
or U116 (N_116,In_325,In_671);
nor U117 (N_117,In_841,In_666);
xor U118 (N_118,In_48,In_522);
nand U119 (N_119,In_293,In_863);
xor U120 (N_120,In_1369,In_782);
nor U121 (N_121,In_498,In_1441);
and U122 (N_122,In_527,In_654);
or U123 (N_123,In_876,In_656);
nand U124 (N_124,In_445,In_1177);
and U125 (N_125,In_580,In_845);
nand U126 (N_126,In_381,In_1447);
or U127 (N_127,In_548,In_871);
nor U128 (N_128,In_331,In_1028);
nor U129 (N_129,In_131,In_601);
xnor U130 (N_130,In_1061,In_860);
and U131 (N_131,In_369,In_1495);
and U132 (N_132,In_291,In_659);
nand U133 (N_133,In_970,In_1224);
and U134 (N_134,In_310,In_1327);
nand U135 (N_135,In_992,In_1123);
and U136 (N_136,In_37,In_29);
xor U137 (N_137,In_596,In_1073);
nand U138 (N_138,In_1124,In_436);
xnor U139 (N_139,In_460,In_1406);
nor U140 (N_140,In_705,In_41);
nand U141 (N_141,In_998,In_567);
nor U142 (N_142,In_828,In_677);
nor U143 (N_143,In_883,In_139);
nand U144 (N_144,In_317,In_865);
nand U145 (N_145,In_278,In_700);
nand U146 (N_146,In_1421,In_388);
nor U147 (N_147,In_602,In_1464);
xnor U148 (N_148,In_107,In_112);
xor U149 (N_149,In_1353,In_22);
or U150 (N_150,In_1499,In_205);
nand U151 (N_151,In_146,In_1399);
xor U152 (N_152,In_680,In_1127);
and U153 (N_153,In_1189,In_1114);
xnor U154 (N_154,In_1303,In_1382);
nand U155 (N_155,In_123,In_287);
nand U156 (N_156,In_1398,In_1243);
nand U157 (N_157,In_1497,In_492);
and U158 (N_158,In_720,In_1043);
nor U159 (N_159,In_437,In_777);
or U160 (N_160,In_209,In_413);
nand U161 (N_161,In_1306,In_1351);
and U162 (N_162,In_1448,In_34);
nor U163 (N_163,In_471,In_1096);
or U164 (N_164,In_354,In_691);
and U165 (N_165,In_563,In_74);
nand U166 (N_166,In_213,In_214);
or U167 (N_167,In_581,In_810);
nand U168 (N_168,In_821,In_964);
nor U169 (N_169,In_558,In_485);
xor U170 (N_170,In_840,In_409);
xnor U171 (N_171,In_647,In_347);
or U172 (N_172,In_1307,In_55);
xnor U173 (N_173,In_1336,In_1350);
or U174 (N_174,In_653,In_1059);
nand U175 (N_175,In_495,In_1249);
and U176 (N_176,In_1184,In_475);
and U177 (N_177,In_743,In_257);
and U178 (N_178,In_807,In_1394);
nor U179 (N_179,In_178,In_1149);
nand U180 (N_180,In_94,In_562);
nand U181 (N_181,In_573,In_956);
nand U182 (N_182,In_1217,In_319);
nand U183 (N_183,In_533,In_750);
nor U184 (N_184,In_117,In_1483);
and U185 (N_185,In_1375,In_891);
nor U186 (N_186,In_1031,In_230);
nand U187 (N_187,In_509,In_1407);
nand U188 (N_188,In_90,In_585);
xor U189 (N_189,In_366,In_446);
or U190 (N_190,In_1075,In_377);
nor U191 (N_191,In_92,In_1471);
or U192 (N_192,In_1103,In_84);
xnor U193 (N_193,In_1486,In_415);
and U194 (N_194,In_113,In_517);
xnor U195 (N_195,In_261,In_245);
and U196 (N_196,In_361,In_940);
nand U197 (N_197,In_1138,In_769);
or U198 (N_198,In_1192,In_173);
nand U199 (N_199,In_843,In_313);
or U200 (N_200,In_771,In_524);
or U201 (N_201,In_1383,In_754);
xor U202 (N_202,In_1147,In_1456);
nor U203 (N_203,In_1226,In_729);
nor U204 (N_204,In_1163,In_1215);
and U205 (N_205,In_594,In_1081);
or U206 (N_206,In_1393,In_526);
nor U207 (N_207,In_599,In_1055);
and U208 (N_208,In_484,In_4);
nor U209 (N_209,In_367,In_429);
xnor U210 (N_210,In_1087,In_657);
xor U211 (N_211,In_868,In_222);
xnor U212 (N_212,In_639,In_1181);
xnor U213 (N_213,In_1162,In_1417);
or U214 (N_214,In_307,In_730);
nor U215 (N_215,In_835,In_462);
and U216 (N_216,In_269,In_125);
nor U217 (N_217,In_833,In_221);
or U218 (N_218,In_1141,In_1320);
or U219 (N_219,In_1247,In_888);
nand U220 (N_220,In_530,In_709);
xor U221 (N_221,In_759,In_793);
nor U222 (N_222,In_39,In_127);
xnor U223 (N_223,In_1468,In_809);
nand U224 (N_224,In_503,In_147);
or U225 (N_225,In_660,In_505);
xnor U226 (N_226,In_1085,In_1068);
or U227 (N_227,In_1329,In_1321);
nor U228 (N_228,In_1062,In_322);
xor U229 (N_229,In_1294,In_844);
nand U230 (N_230,In_983,In_1277);
nor U231 (N_231,In_126,In_167);
nor U232 (N_232,In_937,In_520);
nor U233 (N_233,In_616,In_1481);
or U234 (N_234,In_1405,In_431);
nand U235 (N_235,In_633,In_384);
xor U236 (N_236,In_798,In_1129);
or U237 (N_237,In_1183,In_383);
nor U238 (N_238,In_773,In_515);
xor U239 (N_239,In_764,In_137);
nand U240 (N_240,In_334,In_194);
and U241 (N_241,In_699,In_1131);
xnor U242 (N_242,In_546,In_738);
or U243 (N_243,In_1091,In_746);
xnor U244 (N_244,In_180,In_1324);
nand U245 (N_245,In_1443,In_1034);
or U246 (N_246,In_561,In_1292);
or U247 (N_247,In_28,In_295);
or U248 (N_248,In_504,In_288);
nor U249 (N_249,In_223,In_990);
xnor U250 (N_250,In_1194,In_1171);
and U251 (N_251,In_1025,In_829);
xnor U252 (N_252,In_593,In_423);
nand U253 (N_253,In_1064,In_1159);
or U254 (N_254,In_1066,In_1385);
and U255 (N_255,In_831,In_1396);
or U256 (N_256,In_1409,In_272);
nand U257 (N_257,In_283,In_1144);
xor U258 (N_258,In_85,In_589);
xnor U259 (N_259,In_967,In_962);
or U260 (N_260,In_8,In_145);
or U261 (N_261,In_766,In_432);
and U262 (N_262,In_1009,In_1387);
xnor U263 (N_263,In_668,In_532);
or U264 (N_264,In_344,In_1098);
nand U265 (N_265,In_1208,In_1088);
and U266 (N_266,In_1010,In_756);
xor U267 (N_267,In_805,In_519);
xor U268 (N_268,In_124,In_1234);
or U269 (N_269,In_324,In_978);
or U270 (N_270,In_36,In_501);
and U271 (N_271,In_794,In_359);
xor U272 (N_272,In_249,In_1257);
and U273 (N_273,In_1411,In_1440);
or U274 (N_274,In_1195,In_1370);
or U275 (N_275,In_394,In_40);
xnor U276 (N_276,In_1015,In_627);
xnor U277 (N_277,In_1032,In_748);
nor U278 (N_278,In_575,In_251);
or U279 (N_279,In_1309,In_1432);
and U280 (N_280,In_197,In_243);
nand U281 (N_281,In_236,In_1401);
or U282 (N_282,In_168,In_637);
xor U283 (N_283,In_268,In_215);
nand U284 (N_284,In_490,In_1496);
xor U285 (N_285,In_1187,In_1153);
xnor U286 (N_286,In_685,In_10);
and U287 (N_287,In_45,In_1037);
nand U288 (N_288,In_900,In_1276);
xnor U289 (N_289,In_447,In_421);
nor U290 (N_290,In_1170,In_1487);
or U291 (N_291,In_919,In_1445);
xor U292 (N_292,In_968,In_669);
nor U293 (N_293,In_468,In_1344);
and U294 (N_294,In_578,In_1325);
xor U295 (N_295,In_487,In_143);
nand U296 (N_296,In_1110,In_1083);
and U297 (N_297,In_718,In_456);
or U298 (N_298,In_1197,In_1079);
or U299 (N_299,In_1216,In_634);
or U300 (N_300,In_401,In_1498);
and U301 (N_301,In_452,In_1374);
and U302 (N_302,In_1176,In_239);
nand U303 (N_303,In_1152,In_1218);
nand U304 (N_304,In_177,In_343);
nand U305 (N_305,In_211,In_872);
xor U306 (N_306,In_529,In_449);
or U307 (N_307,In_1000,In_1316);
xor U308 (N_308,In_1386,In_1265);
nor U309 (N_309,In_969,In_1266);
nor U310 (N_310,In_670,In_714);
and U311 (N_311,In_1425,In_329);
xnor U312 (N_312,In_181,In_169);
or U313 (N_313,In_732,In_69);
xnor U314 (N_314,In_1235,In_166);
nor U315 (N_315,In_1284,In_948);
nor U316 (N_316,In_1287,In_237);
and U317 (N_317,In_537,In_148);
and U318 (N_318,In_609,In_1117);
nor U319 (N_319,In_1459,In_1326);
or U320 (N_320,In_623,In_328);
xor U321 (N_321,In_1288,In_1202);
nor U322 (N_322,In_440,In_1104);
nand U323 (N_323,In_1165,In_1455);
or U324 (N_324,In_1173,In_997);
or U325 (N_325,In_799,In_557);
nand U326 (N_326,In_1330,In_789);
xnor U327 (N_327,In_945,In_1041);
xor U328 (N_328,In_695,In_1204);
xnor U329 (N_329,In_476,In_1289);
nand U330 (N_330,In_959,In_502);
nand U331 (N_331,In_1221,In_414);
or U332 (N_332,In_1304,In_82);
nand U333 (N_333,In_1164,In_469);
nand U334 (N_334,In_1271,In_716);
or U335 (N_335,In_1431,In_1439);
xor U336 (N_336,In_1429,In_1494);
or U337 (N_337,In_817,In_1140);
and U338 (N_338,In_444,In_1052);
nor U339 (N_339,In_910,In_947);
nor U340 (N_340,In_751,In_921);
and U341 (N_341,In_1364,In_1036);
or U342 (N_342,In_1315,In_64);
nand U343 (N_343,In_877,In_483);
or U344 (N_344,In_591,In_1054);
or U345 (N_345,In_973,In_932);
nand U346 (N_346,In_62,In_597);
and U347 (N_347,In_1011,In_1179);
and U348 (N_348,In_652,In_312);
nor U349 (N_349,In_586,In_1106);
and U350 (N_350,In_1480,In_118);
xor U351 (N_351,In_75,In_570);
nor U352 (N_352,In_1403,In_908);
nand U353 (N_353,In_507,In_464);
xor U354 (N_354,In_739,In_296);
xnor U355 (N_355,In_1201,In_419);
or U356 (N_356,In_1268,In_864);
nand U357 (N_357,In_1229,In_918);
or U358 (N_358,In_1048,In_905);
and U359 (N_359,In_202,In_1005);
nand U360 (N_360,In_1301,In_813);
nor U361 (N_361,In_849,In_629);
nor U362 (N_362,In_255,In_1363);
nand U363 (N_363,In_50,In_1156);
nor U364 (N_364,In_506,In_227);
nand U365 (N_365,In_626,In_486);
nor U366 (N_366,In_1077,In_160);
and U367 (N_367,In_373,In_545);
xnor U368 (N_368,In_1033,In_1017);
or U369 (N_369,In_672,In_760);
or U370 (N_370,In_370,In_49);
and U371 (N_371,In_1312,In_403);
xnor U372 (N_372,In_203,In_1118);
xnor U373 (N_373,In_881,In_1222);
or U374 (N_374,In_426,In_1372);
or U375 (N_375,In_605,In_97);
nand U376 (N_376,In_89,In_830);
nand U377 (N_377,In_1076,In_353);
or U378 (N_378,In_1021,In_895);
or U379 (N_379,In_280,In_284);
nand U380 (N_380,In_630,In_234);
and U381 (N_381,In_96,In_424);
or U382 (N_382,In_1489,In_768);
nor U383 (N_383,In_1442,In_103);
nand U384 (N_384,In_1102,In_1446);
nand U385 (N_385,In_451,In_866);
nand U386 (N_386,In_534,In_1157);
nand U387 (N_387,In_1296,In_389);
nand U388 (N_388,In_676,In_153);
nand U389 (N_389,In_608,In_1006);
nand U390 (N_390,In_511,In_1155);
nor U391 (N_391,In_775,In_1384);
nand U392 (N_392,In_942,In_1175);
xnor U393 (N_393,In_516,In_33);
nand U394 (N_394,In_265,In_1478);
xor U395 (N_395,In_286,In_87);
xor U396 (N_396,In_374,In_784);
xnor U397 (N_397,In_162,In_1273);
nor U398 (N_398,In_352,In_479);
xnor U399 (N_399,In_628,In_566);
nand U400 (N_400,In_15,In_338);
and U401 (N_401,In_544,In_60);
and U402 (N_402,In_300,In_1328);
xnor U403 (N_403,In_1158,In_1391);
xnor U404 (N_404,In_19,In_1154);
xnor U405 (N_405,In_326,In_1337);
xor U406 (N_406,In_335,In_470);
or U407 (N_407,In_80,In_229);
and U408 (N_408,In_878,In_410);
or U409 (N_409,In_1047,In_355);
nand U410 (N_410,In_349,In_681);
nor U411 (N_411,In_248,In_952);
nor U412 (N_412,In_651,In_1214);
and U413 (N_413,In_737,In_267);
or U414 (N_414,In_102,In_727);
or U415 (N_415,In_600,In_457);
and U416 (N_416,In_816,In_1113);
nand U417 (N_417,In_1404,In_185);
xor U418 (N_418,In_801,In_1122);
and U419 (N_419,In_551,In_879);
nand U420 (N_420,In_408,In_54);
and U421 (N_421,In_1274,In_242);
nand U422 (N_422,In_1207,In_1473);
and U423 (N_423,In_684,In_93);
xor U424 (N_424,In_375,In_542);
and U425 (N_425,In_31,In_854);
or U426 (N_426,In_933,In_980);
nor U427 (N_427,In_867,In_1090);
or U428 (N_428,In_853,In_901);
or U429 (N_429,In_282,In_358);
nor U430 (N_430,In_620,In_391);
or U431 (N_431,In_1286,In_1291);
nand U432 (N_432,In_422,In_1360);
nor U433 (N_433,In_667,In_294);
xnor U434 (N_434,In_1430,In_489);
nor U435 (N_435,In_1335,In_478);
xor U436 (N_436,In_1451,In_949);
nor U437 (N_437,In_1342,In_664);
nor U438 (N_438,In_1125,In_508);
nor U439 (N_439,In_472,In_61);
and U440 (N_440,In_514,In_850);
and U441 (N_441,In_971,In_770);
nor U442 (N_442,In_232,In_1313);
nand U443 (N_443,In_1339,In_65);
nand U444 (N_444,In_1465,In_1018);
and U445 (N_445,In_682,In_1338);
nand U446 (N_446,In_1050,In_1323);
and U447 (N_447,In_1220,In_902);
and U448 (N_448,In_642,In_1180);
nor U449 (N_449,In_621,In_434);
xnor U450 (N_450,In_1492,In_1479);
and U451 (N_451,In_1420,In_722);
xnor U452 (N_452,In_938,In_1345);
nand U453 (N_453,In_1435,In_1469);
or U454 (N_454,In_698,In_17);
xnor U455 (N_455,In_277,In_208);
and U456 (N_456,In_624,In_862);
nor U457 (N_457,In_1026,In_70);
nor U458 (N_458,In_364,In_1367);
nor U459 (N_459,In_1108,In_995);
xor U460 (N_460,In_95,In_199);
nor U461 (N_461,In_974,In_182);
nand U462 (N_462,In_79,In_306);
and U463 (N_463,In_253,In_11);
nor U464 (N_464,In_1493,In_1365);
and U465 (N_465,In_625,In_1057);
and U466 (N_466,In_1193,In_512);
xor U467 (N_467,In_688,In_822);
xor U468 (N_468,In_644,In_467);
or U469 (N_469,In_1426,In_767);
or U470 (N_470,In_610,In_281);
nand U471 (N_471,In_16,In_814);
nand U472 (N_472,In_875,In_1228);
and U473 (N_473,In_1285,In_412);
or U474 (N_474,In_441,In_297);
nand U475 (N_475,In_1244,In_839);
xor U476 (N_476,In_387,In_20);
or U477 (N_477,In_710,In_923);
or U478 (N_478,In_724,In_786);
xor U479 (N_479,In_1174,In_1053);
nor U480 (N_480,In_880,In_1160);
or U481 (N_481,In_961,In_406);
xnor U482 (N_482,In_934,In_1236);
or U483 (N_483,In_238,In_858);
or U484 (N_484,In_1415,In_1362);
and U485 (N_485,In_1463,In_1354);
and U486 (N_486,In_697,In_966);
or U487 (N_487,In_1262,In_582);
nand U488 (N_488,In_192,In_252);
and U489 (N_489,In_776,In_991);
nor U490 (N_490,In_550,In_1416);
and U491 (N_491,In_1072,In_273);
nand U492 (N_492,In_1150,In_285);
nand U493 (N_493,In_808,In_1452);
and U494 (N_494,In_116,In_890);
or U495 (N_495,In_196,In_1116);
nand U496 (N_496,In_797,In_1069);
xnor U497 (N_497,In_1314,In_266);
and U498 (N_498,In_453,In_72);
or U499 (N_499,In_790,In_678);
nor U500 (N_500,In_663,In_27);
nand U501 (N_501,N_143,N_98);
nand U502 (N_502,N_330,In_1185);
nand U503 (N_503,In_590,In_395);
or U504 (N_504,In_694,N_59);
and U505 (N_505,In_1256,In_513);
xnor U506 (N_506,In_1263,In_1438);
nand U507 (N_507,N_226,In_397);
or U508 (N_508,N_498,N_47);
or U509 (N_509,N_80,In_38);
nand U510 (N_510,N_395,In_165);
xnor U511 (N_511,In_14,In_604);
and U512 (N_512,In_926,In_240);
nand U513 (N_513,In_1454,In_1119);
nor U514 (N_514,N_191,In_88);
nor U515 (N_515,N_322,In_941);
and U516 (N_516,N_207,N_400);
xnor U517 (N_517,In_851,N_377);
or U518 (N_518,In_713,In_1449);
and U519 (N_519,In_611,N_405);
xor U520 (N_520,N_192,In_1332);
or U521 (N_521,N_205,N_289);
or U522 (N_522,In_466,N_83);
or U523 (N_523,N_89,N_431);
and U524 (N_524,In_577,In_260);
nor U525 (N_525,N_203,N_197);
nand U526 (N_526,In_465,N_389);
and U527 (N_527,N_491,In_1474);
nor U528 (N_528,N_42,In_405);
nor U529 (N_529,In_1260,In_259);
xor U530 (N_530,In_539,N_167);
nor U531 (N_531,In_741,N_294);
or U532 (N_532,N_362,N_333);
and U533 (N_533,In_1143,N_107);
or U534 (N_534,N_272,In_846);
and U535 (N_535,In_128,In_332);
and U536 (N_536,N_78,In_379);
nand U537 (N_537,In_1007,N_18);
nand U538 (N_538,In_1317,N_221);
xor U539 (N_539,N_369,N_396);
nor U540 (N_540,N_470,N_261);
nor U541 (N_541,In_914,N_303);
or U542 (N_542,In_690,In_104);
nand U543 (N_543,In_717,In_1366);
and U544 (N_544,In_946,N_124);
and U545 (N_545,In_132,In_341);
or U546 (N_546,In_1444,In_658);
nand U547 (N_547,N_53,N_184);
or U548 (N_548,In_1112,N_229);
xnor U549 (N_549,In_1427,N_0);
or U550 (N_550,N_6,N_196);
and U551 (N_551,N_230,In_393);
or U552 (N_552,N_108,In_1056);
xnor U553 (N_553,N_131,In_747);
or U554 (N_554,N_390,N_284);
and U555 (N_555,N_129,In_930);
nor U556 (N_556,N_141,N_324);
nand U557 (N_557,N_401,In_953);
nand U558 (N_558,N_337,In_556);
or U559 (N_559,N_217,In_989);
and U560 (N_560,N_479,In_904);
nand U561 (N_561,In_538,In_825);
xnor U562 (N_562,N_29,N_465);
or U563 (N_563,N_402,N_356);
nand U564 (N_564,N_305,N_264);
or U565 (N_565,N_90,N_74);
xor U566 (N_566,In_612,In_321);
or U567 (N_567,In_1397,N_318);
xor U568 (N_568,N_25,In_241);
xnor U569 (N_569,In_1199,N_429);
nor U570 (N_570,In_301,In_981);
or U571 (N_571,In_702,N_104);
or U572 (N_572,N_457,N_100);
or U573 (N_573,In_348,N_443);
nand U574 (N_574,N_32,N_286);
or U575 (N_575,N_71,N_73);
nand U576 (N_576,In_823,In_392);
xnor U577 (N_577,N_291,N_288);
and U578 (N_578,N_478,In_12);
and U579 (N_579,In_712,N_148);
and U580 (N_580,In_719,N_281);
or U581 (N_581,N_418,N_342);
nand U582 (N_582,In_482,In_271);
nand U583 (N_583,N_296,In_411);
or U584 (N_584,N_157,In_728);
or U585 (N_585,In_1242,In_540);
nand U586 (N_586,N_338,N_138);
nor U587 (N_587,In_246,In_1252);
and U588 (N_588,In_76,In_443);
nand U589 (N_589,In_1310,In_703);
xor U590 (N_590,In_368,In_795);
nor U591 (N_591,In_219,N_233);
nor U592 (N_592,In_1297,In_140);
xor U593 (N_593,N_411,N_391);
xor U594 (N_594,In_1484,N_16);
nand U595 (N_595,N_359,In_330);
nand U596 (N_596,In_496,N_308);
and U597 (N_597,In_572,In_603);
xor U598 (N_598,In_1245,N_476);
nand U599 (N_599,In_1027,N_152);
nand U600 (N_600,In_1035,In_198);
nand U601 (N_601,In_1462,N_420);
or U602 (N_602,In_916,N_494);
nor U603 (N_603,N_285,N_436);
xor U604 (N_604,N_248,In_936);
xor U605 (N_605,N_379,In_417);
and U606 (N_606,N_119,In_292);
or U607 (N_607,N_2,N_113);
or U608 (N_608,In_655,In_1389);
nand U609 (N_609,N_309,N_497);
nor U610 (N_610,N_162,N_215);
nor U611 (N_611,In_1101,In_646);
nor U612 (N_612,N_433,In_1093);
nor U613 (N_613,In_435,In_497);
and U614 (N_614,In_958,In_1240);
nand U615 (N_615,N_154,In_987);
or U616 (N_616,N_245,N_188);
or U617 (N_617,In_1142,N_106);
and U618 (N_618,N_256,In_274);
nand U619 (N_619,N_327,In_1437);
and U620 (N_620,In_493,In_979);
and U621 (N_621,In_726,In_584);
nor U622 (N_622,In_63,N_246);
and U623 (N_623,N_354,N_387);
and U624 (N_624,N_358,N_234);
and U625 (N_625,N_101,N_344);
or U626 (N_626,N_22,N_121);
xor U627 (N_627,N_187,N_332);
nand U628 (N_628,N_475,In_836);
nand U629 (N_629,N_4,N_7);
nor U630 (N_630,In_778,N_15);
and U631 (N_631,In_1311,N_331);
or U632 (N_632,N_111,N_118);
xnor U633 (N_633,In_480,N_65);
and U634 (N_634,In_263,N_414);
nand U635 (N_635,N_399,N_232);
xor U636 (N_636,N_46,In_950);
and U637 (N_637,N_45,In_351);
nand U638 (N_638,In_1082,N_373);
xnor U639 (N_639,N_441,In_1278);
or U640 (N_640,In_924,In_1191);
or U641 (N_641,N_365,N_440);
and U642 (N_642,In_1084,In_622);
or U643 (N_643,In_765,In_665);
or U644 (N_644,N_142,In_6);
nand U645 (N_645,N_202,N_198);
nor U646 (N_646,In_1134,In_696);
nor U647 (N_647,N_166,N_406);
or U648 (N_648,In_1024,N_381);
or U649 (N_649,In_372,In_270);
nor U650 (N_650,In_336,In_927);
or U651 (N_651,N_276,In_1128);
xnor U652 (N_652,N_147,In_761);
or U653 (N_653,In_510,N_145);
nand U654 (N_654,N_383,N_149);
nand U655 (N_655,N_277,In_188);
nand U656 (N_656,In_1167,N_123);
or U657 (N_657,In_114,N_370);
nand U658 (N_658,N_258,N_378);
and U659 (N_659,In_43,In_1371);
xor U660 (N_660,N_304,In_418);
nand U661 (N_661,In_71,In_1460);
nor U662 (N_662,In_250,N_39);
nand U663 (N_663,In_1331,N_485);
nor U664 (N_664,In_1472,N_102);
xnor U665 (N_665,In_416,In_1);
xor U666 (N_666,N_220,N_14);
nor U667 (N_667,N_360,In_1343);
or U668 (N_668,In_105,In_791);
nor U669 (N_669,In_1198,In_53);
and U670 (N_670,N_326,N_403);
or U671 (N_671,In_1349,N_48);
and U672 (N_672,N_77,In_675);
nand U673 (N_673,In_150,N_404);
nor U674 (N_674,In_931,N_193);
and U675 (N_675,N_355,N_435);
xor U676 (N_676,N_92,N_170);
nor U677 (N_677,In_1280,In_553);
or U678 (N_678,In_1178,N_487);
nand U679 (N_679,In_461,N_320);
xor U680 (N_680,In_925,In_1169);
and U681 (N_681,N_125,In_1205);
nor U682 (N_682,N_474,N_456);
and U683 (N_683,N_267,N_164);
nor U684 (N_684,N_237,In_1254);
or U685 (N_685,In_224,N_386);
or U686 (N_686,N_481,In_943);
nor U687 (N_687,In_78,N_225);
or U688 (N_688,In_679,N_117);
xor U689 (N_689,In_763,In_640);
nand U690 (N_690,In_1225,N_375);
and U691 (N_691,In_320,In_1377);
nand U692 (N_692,In_1275,In_316);
and U693 (N_693,In_1461,In_3);
nand U694 (N_694,In_175,In_425);
and U695 (N_695,N_109,N_323);
xnor U696 (N_696,N_51,N_273);
xor U697 (N_697,N_130,In_882);
xnor U698 (N_698,In_569,N_325);
nor U699 (N_699,In_708,N_366);
or U700 (N_700,In_988,In_606);
nor U701 (N_701,In_752,N_12);
and U702 (N_702,In_909,N_54);
xnor U703 (N_703,In_859,In_523);
and U704 (N_704,N_484,N_75);
nand U705 (N_705,In_1419,N_467);
or U706 (N_706,N_447,N_460);
nor U707 (N_707,In_120,In_827);
nor U708 (N_708,N_96,N_278);
or U709 (N_709,N_329,N_115);
nand U710 (N_710,N_274,In_1097);
or U711 (N_711,In_189,N_409);
xor U712 (N_712,In_142,N_128);
and U713 (N_713,N_415,N_82);
nor U714 (N_714,In_903,N_171);
nor U715 (N_715,N_10,In_1413);
nand U716 (N_716,N_260,In_365);
or U717 (N_717,In_183,In_855);
nor U718 (N_718,In_308,N_69);
xnor U719 (N_719,N_156,N_471);
or U720 (N_720,N_295,In_499);
nor U721 (N_721,N_445,In_342);
and U722 (N_722,In_149,In_184);
nand U723 (N_723,N_301,In_458);
or U724 (N_724,N_252,In_427);
nor U725 (N_725,In_944,N_419);
and U726 (N_726,In_1300,N_434);
xnor U727 (N_727,In_857,In_815);
nor U728 (N_728,In_975,N_492);
nand U729 (N_729,In_796,In_136);
and U730 (N_730,In_254,In_913);
and U731 (N_731,N_186,In_1246);
nand U732 (N_732,N_228,N_3);
and U733 (N_733,N_263,In_1067);
xnor U734 (N_734,In_1392,In_204);
nor U735 (N_735,N_63,N_163);
xnor U736 (N_736,In_686,In_1211);
nor U737 (N_737,N_194,N_133);
and U738 (N_738,N_413,In_1476);
or U739 (N_739,In_303,In_57);
and U740 (N_740,In_749,N_62);
or U741 (N_741,In_951,In_1450);
and U742 (N_742,In_636,N_271);
nor U743 (N_743,In_1380,N_1);
xor U744 (N_744,N_79,N_158);
xor U745 (N_745,In_1470,N_316);
and U746 (N_746,In_1433,N_255);
nand U747 (N_747,In_535,In_371);
nor U748 (N_748,In_163,N_95);
xor U749 (N_749,N_417,N_336);
xor U750 (N_750,N_56,N_268);
xor U751 (N_751,In_595,N_208);
and U752 (N_752,In_433,N_345);
nand U753 (N_753,In_463,In_450);
xor U754 (N_754,N_270,In_986);
xor U755 (N_755,N_126,In_1453);
nand U756 (N_756,In_363,In_1361);
or U757 (N_757,N_81,N_20);
xor U758 (N_758,In_984,N_247);
xnor U759 (N_759,In_459,N_64);
nand U760 (N_760,N_210,N_227);
xnor U761 (N_761,N_76,N_132);
nand U762 (N_762,In_755,In_212);
xor U763 (N_763,N_176,In_787);
nand U764 (N_764,N_201,In_201);
nand U765 (N_765,N_266,In_1412);
nand U766 (N_766,N_195,N_212);
and U767 (N_767,In_982,In_886);
nor U768 (N_768,In_500,In_1109);
and U769 (N_769,N_361,N_116);
and U770 (N_770,In_1022,N_213);
nand U771 (N_771,In_554,N_68);
or U772 (N_772,N_11,In_179);
or U773 (N_773,N_463,In_579);
xnor U774 (N_774,In_811,N_340);
and U775 (N_775,In_820,In_1348);
nor U776 (N_776,In_1070,In_1281);
nor U777 (N_777,In_826,N_483);
xor U778 (N_778,In_1042,In_1019);
xor U779 (N_779,N_33,In_99);
or U780 (N_780,N_97,In_1293);
and U781 (N_781,N_394,In_115);
and U782 (N_782,N_40,In_101);
or U783 (N_783,N_493,N_426);
and U784 (N_784,N_346,In_438);
nand U785 (N_785,N_453,N_466);
and U786 (N_786,N_67,N_218);
nor U787 (N_787,N_464,In_1003);
nand U788 (N_788,In_662,N_8);
or U789 (N_789,N_462,In_687);
and U790 (N_790,In_191,N_490);
nor U791 (N_791,N_350,N_292);
nor U792 (N_792,In_1227,In_781);
xnor U793 (N_793,In_528,N_249);
nand U794 (N_794,N_444,N_178);
nand U795 (N_795,In_1251,N_150);
and U796 (N_796,In_129,In_1014);
or U797 (N_797,N_449,In_77);
xnor U798 (N_798,N_204,In_323);
or U799 (N_799,N_85,In_735);
nand U800 (N_800,In_1352,In_108);
nor U801 (N_801,N_250,In_314);
xor U802 (N_802,In_1457,In_1376);
nand U803 (N_803,N_482,N_161);
and U804 (N_804,In_174,N_9);
nand U805 (N_805,N_472,N_446);
or U806 (N_806,In_1482,N_328);
or U807 (N_807,In_327,In_1100);
xor U808 (N_808,N_41,N_120);
nand U809 (N_809,N_349,In_832);
nor U810 (N_810,In_1107,N_279);
or U811 (N_811,N_282,In_704);
nor U812 (N_812,In_929,N_24);
and U813 (N_813,In_1458,In_615);
nand U814 (N_814,In_733,N_58);
xnor U815 (N_815,In_922,N_459);
and U816 (N_816,N_306,N_242);
nor U817 (N_817,In_23,N_135);
or U818 (N_818,N_380,In_159);
nand U819 (N_819,N_262,In_1422);
and U820 (N_820,N_88,In_1491);
nand U821 (N_821,In_1137,N_280);
nor U822 (N_822,N_384,In_1381);
nor U823 (N_823,N_155,In_803);
and U824 (N_824,In_889,N_87);
or U825 (N_825,N_496,In_693);
and U826 (N_826,In_762,N_151);
or U827 (N_827,In_1414,N_236);
nor U828 (N_828,In_689,N_432);
or U829 (N_829,In_276,N_223);
nand U830 (N_830,N_442,N_19);
nor U831 (N_831,In_1020,N_240);
xnor U832 (N_832,In_1030,In_892);
and U833 (N_833,In_1099,N_31);
nor U834 (N_834,In_217,N_136);
or U835 (N_835,In_32,N_146);
and U836 (N_836,N_334,In_852);
or U837 (N_837,N_38,N_70);
or U838 (N_838,In_494,N_181);
nand U839 (N_839,N_57,N_49);
or U840 (N_840,N_37,In_176);
xnor U841 (N_841,N_177,In_1058);
nand U842 (N_842,N_105,N_454);
nor U843 (N_843,In_631,N_60);
and U844 (N_844,N_352,In_1466);
or U845 (N_845,In_707,N_259);
nor U846 (N_846,N_99,In_315);
nand U847 (N_847,N_110,In_481);
nor U848 (N_848,In_1146,N_319);
nor U849 (N_849,In_1071,In_917);
or U850 (N_850,In_9,In_111);
nand U851 (N_851,N_347,In_861);
and U852 (N_852,N_297,In_56);
nand U853 (N_853,N_293,N_93);
nand U854 (N_854,N_190,N_91);
nor U855 (N_855,In_455,N_219);
and U856 (N_856,N_372,N_13);
xnor U857 (N_857,N_86,N_139);
and U858 (N_858,In_156,In_607);
or U859 (N_859,In_133,In_311);
nand U860 (N_860,N_314,In_614);
and U861 (N_861,In_26,N_175);
or U862 (N_862,N_312,N_214);
nor U863 (N_863,In_430,In_887);
nand U864 (N_864,N_28,In_58);
nand U865 (N_865,In_454,N_290);
nor U866 (N_866,N_23,In_838);
nor U867 (N_867,N_423,In_1086);
or U868 (N_868,N_385,In_1203);
nand U869 (N_869,In_109,N_317);
nand U870 (N_870,N_34,N_458);
xor U871 (N_871,N_451,In_912);
and U872 (N_872,N_84,N_439);
and U873 (N_873,In_635,In_171);
and U874 (N_874,N_182,In_1212);
and U875 (N_875,N_275,N_437);
nand U876 (N_876,N_160,N_5);
nand U877 (N_877,N_367,In_226);
nand U878 (N_878,In_333,In_1402);
xnor U879 (N_879,N_165,N_448);
xnor U880 (N_880,In_262,N_427);
xor U881 (N_881,In_643,In_745);
or U882 (N_882,N_199,N_222);
nor U883 (N_883,In_648,N_172);
nor U884 (N_884,In_1223,N_300);
nor U885 (N_885,In_1023,In_785);
and U886 (N_886,In_83,In_1359);
or U887 (N_887,N_343,N_103);
and U888 (N_888,In_920,N_238);
or U889 (N_889,In_1308,In_1094);
or U890 (N_890,N_231,In_736);
or U891 (N_891,In_1148,In_2);
xor U892 (N_892,In_1261,N_241);
xnor U893 (N_893,N_94,In_1237);
nor U894 (N_894,In_190,N_36);
nand U895 (N_895,In_42,N_408);
nor U896 (N_896,N_243,In_641);
and U897 (N_897,In_1322,N_269);
or U898 (N_898,In_1333,N_209);
xor U899 (N_899,N_315,In_757);
and U900 (N_900,N_174,In_298);
and U901 (N_901,In_559,N_489);
or U902 (N_902,In_357,In_134);
or U903 (N_903,N_335,In_350);
or U904 (N_904,N_17,In_1002);
or U905 (N_905,N_397,In_264);
and U906 (N_906,In_135,N_43);
nand U907 (N_907,N_159,In_541);
and U908 (N_908,N_180,In_1074);
nor U909 (N_909,In_1346,N_307);
nand U910 (N_910,In_565,In_386);
nand U911 (N_911,In_1423,N_311);
or U912 (N_912,N_488,In_1395);
and U913 (N_913,N_127,In_885);
nor U914 (N_914,N_137,In_721);
nand U915 (N_915,In_935,In_25);
nor U916 (N_916,N_393,N_421);
nand U917 (N_917,In_1319,In_1238);
nor U918 (N_918,N_339,N_341);
nand U919 (N_919,In_290,N_265);
and U920 (N_920,N_388,N_351);
xor U921 (N_921,N_185,In_1259);
nand U922 (N_922,In_1341,In_256);
nand U923 (N_923,In_1038,N_254);
and U924 (N_924,In_407,N_216);
nand U925 (N_925,N_310,In_1270);
xnor U926 (N_926,N_425,In_772);
and U927 (N_927,In_1400,In_1190);
xnor U928 (N_928,In_130,In_928);
nand U929 (N_929,N_353,In_911);
or U930 (N_930,N_224,In_723);
and U931 (N_931,N_398,N_189);
xor U932 (N_932,N_179,N_368);
nand U933 (N_933,N_452,N_55);
nor U934 (N_934,N_407,In_906);
nand U935 (N_935,In_661,In_247);
nor U936 (N_936,In_834,N_299);
xnor U937 (N_937,In_1355,N_52);
nor U938 (N_938,N_251,N_72);
nor U939 (N_939,In_552,In_1267);
or U940 (N_940,N_499,In_1049);
and U941 (N_941,N_416,N_438);
or U942 (N_942,N_153,N_168);
nand U943 (N_943,N_450,In_51);
xnor U944 (N_944,In_477,N_183);
and U945 (N_945,In_235,N_61);
and U946 (N_946,N_206,In_1219);
nor U947 (N_947,In_1188,N_122);
and U948 (N_948,In_673,N_371);
nand U949 (N_949,In_1373,N_211);
nand U950 (N_950,N_287,N_480);
or U951 (N_951,N_477,In_874);
or U952 (N_952,In_491,N_495);
and U953 (N_953,In_1334,N_44);
nand U954 (N_954,N_374,In_195);
nor U955 (N_955,In_7,N_134);
nor U956 (N_956,N_26,N_455);
xor U957 (N_957,In_1231,In_706);
or U958 (N_958,In_525,N_112);
nand U959 (N_959,N_357,N_30);
nand U960 (N_960,N_376,In_21);
nor U961 (N_961,In_692,In_847);
nor U962 (N_962,N_114,In_731);
nor U963 (N_963,N_313,In_1290);
xor U964 (N_964,In_1139,In_1488);
or U965 (N_965,In_100,N_382);
nor U966 (N_966,N_473,In_67);
xnor U967 (N_967,In_157,In_1368);
or U968 (N_968,N_302,In_1145);
and U969 (N_969,In_18,In_13);
xnor U970 (N_970,In_52,N_412);
nand U971 (N_971,In_1046,In_571);
xor U972 (N_972,N_392,In_683);
xor U973 (N_973,In_1004,N_27);
nand U974 (N_974,In_999,N_66);
xnor U975 (N_975,In_1305,In_1477);
nor U976 (N_976,N_486,N_253);
nand U977 (N_977,In_396,In_1092);
and U978 (N_978,In_725,N_169);
or U979 (N_979,N_140,In_275);
or U980 (N_980,In_339,In_873);
nand U981 (N_981,N_239,N_50);
xor U982 (N_982,In_346,N_298);
xnor U983 (N_983,In_818,In_399);
nor U984 (N_984,N_461,In_587);
xnor U985 (N_985,In_711,N_257);
or U986 (N_986,In_848,N_428);
xor U987 (N_987,In_119,In_965);
and U988 (N_988,N_422,In_170);
nor U989 (N_989,N_173,N_200);
nor U990 (N_990,N_424,N_363);
nor U991 (N_991,N_235,In_1255);
nand U992 (N_992,In_1012,N_321);
or U993 (N_993,N_283,N_468);
nor U994 (N_994,N_21,In_856);
and U995 (N_995,N_469,N_348);
nand U996 (N_996,N_364,N_430);
and U997 (N_997,N_410,N_144);
nand U998 (N_998,In_144,In_800);
and U999 (N_999,N_244,N_35);
xnor U1000 (N_1000,N_692,N_835);
nor U1001 (N_1001,N_763,N_811);
nand U1002 (N_1002,N_874,N_676);
or U1003 (N_1003,N_813,N_974);
and U1004 (N_1004,N_681,N_607);
nor U1005 (N_1005,N_520,N_512);
nand U1006 (N_1006,N_637,N_724);
nand U1007 (N_1007,N_820,N_816);
and U1008 (N_1008,N_620,N_933);
xnor U1009 (N_1009,N_690,N_927);
or U1010 (N_1010,N_897,N_998);
and U1011 (N_1011,N_719,N_671);
and U1012 (N_1012,N_852,N_505);
nand U1013 (N_1013,N_901,N_652);
and U1014 (N_1014,N_696,N_950);
nand U1015 (N_1015,N_986,N_904);
and U1016 (N_1016,N_643,N_632);
and U1017 (N_1017,N_994,N_844);
nand U1018 (N_1018,N_554,N_794);
and U1019 (N_1019,N_604,N_859);
or U1020 (N_1020,N_513,N_899);
nor U1021 (N_1021,N_656,N_526);
nand U1022 (N_1022,N_629,N_702);
and U1023 (N_1023,N_806,N_644);
nand U1024 (N_1024,N_990,N_535);
or U1025 (N_1025,N_945,N_548);
and U1026 (N_1026,N_837,N_679);
or U1027 (N_1027,N_583,N_880);
nand U1028 (N_1028,N_853,N_865);
or U1029 (N_1029,N_660,N_570);
and U1030 (N_1030,N_868,N_791);
nor U1031 (N_1031,N_747,N_515);
nor U1032 (N_1032,N_939,N_675);
nand U1033 (N_1033,N_966,N_805);
and U1034 (N_1034,N_595,N_944);
or U1035 (N_1035,N_665,N_797);
and U1036 (N_1036,N_888,N_686);
nor U1037 (N_1037,N_642,N_650);
nor U1038 (N_1038,N_889,N_543);
nor U1039 (N_1039,N_908,N_792);
xnor U1040 (N_1040,N_736,N_824);
xnor U1041 (N_1041,N_674,N_598);
and U1042 (N_1042,N_864,N_815);
xor U1043 (N_1043,N_909,N_552);
nor U1044 (N_1044,N_694,N_788);
and U1045 (N_1045,N_663,N_553);
xnor U1046 (N_1046,N_761,N_819);
or U1047 (N_1047,N_712,N_978);
or U1048 (N_1048,N_551,N_539);
nor U1049 (N_1049,N_749,N_817);
or U1050 (N_1050,N_758,N_695);
xnor U1051 (N_1051,N_959,N_963);
and U1052 (N_1052,N_947,N_587);
nand U1053 (N_1053,N_508,N_930);
nor U1054 (N_1054,N_731,N_661);
xor U1055 (N_1055,N_634,N_854);
and U1056 (N_1056,N_659,N_910);
nor U1057 (N_1057,N_953,N_725);
xor U1058 (N_1058,N_795,N_765);
xnor U1059 (N_1059,N_918,N_952);
nand U1060 (N_1060,N_649,N_654);
and U1061 (N_1061,N_914,N_895);
or U1062 (N_1062,N_563,N_970);
or U1063 (N_1063,N_684,N_962);
or U1064 (N_1064,N_796,N_743);
nor U1065 (N_1065,N_705,N_774);
or U1066 (N_1066,N_999,N_834);
xnor U1067 (N_1067,N_872,N_677);
and U1068 (N_1068,N_510,N_704);
and U1069 (N_1069,N_667,N_697);
xor U1070 (N_1070,N_562,N_750);
xnor U1071 (N_1071,N_532,N_893);
and U1072 (N_1072,N_603,N_900);
nand U1073 (N_1073,N_975,N_716);
xor U1074 (N_1074,N_685,N_584);
nand U1075 (N_1075,N_809,N_589);
nand U1076 (N_1076,N_746,N_862);
nor U1077 (N_1077,N_582,N_720);
nor U1078 (N_1078,N_845,N_992);
xnor U1079 (N_1079,N_803,N_730);
and U1080 (N_1080,N_640,N_879);
nor U1081 (N_1081,N_519,N_954);
nor U1082 (N_1082,N_514,N_549);
nor U1083 (N_1083,N_613,N_842);
nand U1084 (N_1084,N_506,N_576);
or U1085 (N_1085,N_504,N_622);
and U1086 (N_1086,N_848,N_925);
or U1087 (N_1087,N_734,N_556);
nand U1088 (N_1088,N_524,N_631);
xnor U1089 (N_1089,N_830,N_832);
and U1090 (N_1090,N_827,N_594);
nor U1091 (N_1091,N_718,N_534);
nand U1092 (N_1092,N_866,N_841);
nor U1093 (N_1093,N_687,N_799);
or U1094 (N_1094,N_801,N_711);
and U1095 (N_1095,N_503,N_657);
or U1096 (N_1096,N_957,N_780);
nand U1097 (N_1097,N_574,N_863);
nor U1098 (N_1098,N_522,N_575);
and U1099 (N_1099,N_883,N_988);
xnor U1100 (N_1100,N_516,N_915);
or U1101 (N_1101,N_818,N_599);
nand U1102 (N_1102,N_886,N_931);
or U1103 (N_1103,N_987,N_728);
nand U1104 (N_1104,N_804,N_639);
xor U1105 (N_1105,N_776,N_766);
and U1106 (N_1106,N_942,N_849);
and U1107 (N_1107,N_767,N_628);
or U1108 (N_1108,N_569,N_567);
nand U1109 (N_1109,N_860,N_713);
and U1110 (N_1110,N_536,N_960);
or U1111 (N_1111,N_977,N_938);
and U1112 (N_1112,N_601,N_892);
nor U1113 (N_1113,N_839,N_826);
xnor U1114 (N_1114,N_688,N_588);
nor U1115 (N_1115,N_608,N_903);
xor U1116 (N_1116,N_623,N_840);
or U1117 (N_1117,N_614,N_812);
or U1118 (N_1118,N_611,N_814);
and U1119 (N_1119,N_609,N_670);
nand U1120 (N_1120,N_760,N_751);
or U1121 (N_1121,N_937,N_956);
and U1122 (N_1122,N_983,N_870);
and U1123 (N_1123,N_579,N_691);
nor U1124 (N_1124,N_600,N_754);
xor U1125 (N_1125,N_559,N_615);
nor U1126 (N_1126,N_861,N_917);
nor U1127 (N_1127,N_778,N_920);
and U1128 (N_1128,N_528,N_672);
nor U1129 (N_1129,N_737,N_913);
xnor U1130 (N_1130,N_891,N_568);
xor U1131 (N_1131,N_597,N_878);
xor U1132 (N_1132,N_932,N_748);
and U1133 (N_1133,N_790,N_919);
or U1134 (N_1134,N_785,N_664);
and U1135 (N_1135,N_969,N_668);
and U1136 (N_1136,N_653,N_940);
xor U1137 (N_1137,N_698,N_936);
and U1138 (N_1138,N_928,N_961);
or U1139 (N_1139,N_838,N_735);
nor U1140 (N_1140,N_565,N_523);
xnor U1141 (N_1141,N_828,N_509);
or U1142 (N_1142,N_592,N_912);
xor U1143 (N_1143,N_924,N_922);
or U1144 (N_1144,N_547,N_773);
xor U1145 (N_1145,N_545,N_745);
xnor U1146 (N_1146,N_882,N_984);
or U1147 (N_1147,N_951,N_602);
nor U1148 (N_1148,N_772,N_666);
nor U1149 (N_1149,N_875,N_525);
nor U1150 (N_1150,N_511,N_911);
nand U1151 (N_1151,N_890,N_810);
nand U1152 (N_1152,N_981,N_612);
xnor U1153 (N_1153,N_829,N_896);
nand U1154 (N_1154,N_968,N_802);
nand U1155 (N_1155,N_560,N_630);
or U1156 (N_1156,N_771,N_831);
nor U1157 (N_1157,N_616,N_996);
or U1158 (N_1158,N_775,N_501);
and U1159 (N_1159,N_926,N_581);
and U1160 (N_1160,N_707,N_573);
nand U1161 (N_1161,N_699,N_965);
xor U1162 (N_1162,N_625,N_894);
nor U1163 (N_1163,N_757,N_836);
nor U1164 (N_1164,N_706,N_997);
xnor U1165 (N_1165,N_590,N_738);
nor U1166 (N_1166,N_651,N_557);
and U1167 (N_1167,N_858,N_921);
and U1168 (N_1168,N_729,N_638);
or U1169 (N_1169,N_800,N_610);
xnor U1170 (N_1170,N_876,N_626);
xnor U1171 (N_1171,N_873,N_821);
nor U1172 (N_1172,N_700,N_782);
nand U1173 (N_1173,N_578,N_744);
xor U1174 (N_1174,N_635,N_722);
xor U1175 (N_1175,N_732,N_564);
nand U1176 (N_1176,N_518,N_558);
or U1177 (N_1177,N_784,N_586);
nand U1178 (N_1178,N_807,N_976);
xor U1179 (N_1179,N_647,N_869);
or U1180 (N_1180,N_833,N_636);
nand U1181 (N_1181,N_934,N_658);
nor U1182 (N_1182,N_871,N_777);
nand U1183 (N_1183,N_979,N_742);
xor U1184 (N_1184,N_881,N_789);
nor U1185 (N_1185,N_566,N_943);
nand U1186 (N_1186,N_645,N_958);
or U1187 (N_1187,N_843,N_980);
xor U1188 (N_1188,N_972,N_624);
xor U1189 (N_1189,N_714,N_884);
nand U1190 (N_1190,N_708,N_544);
nand U1191 (N_1191,N_507,N_641);
nor U1192 (N_1192,N_759,N_529);
or U1193 (N_1193,N_948,N_701);
xnor U1194 (N_1194,N_825,N_537);
and U1195 (N_1195,N_605,N_500);
and U1196 (N_1196,N_929,N_682);
or U1197 (N_1197,N_689,N_521);
xnor U1198 (N_1198,N_550,N_787);
xnor U1199 (N_1199,N_546,N_561);
xor U1200 (N_1200,N_555,N_793);
and U1201 (N_1201,N_762,N_517);
or U1202 (N_1202,N_973,N_887);
xnor U1203 (N_1203,N_709,N_715);
or U1204 (N_1204,N_619,N_673);
nor U1205 (N_1205,N_741,N_606);
or U1206 (N_1206,N_867,N_955);
nor U1207 (N_1207,N_571,N_753);
nor U1208 (N_1208,N_991,N_769);
and U1209 (N_1209,N_627,N_898);
and U1210 (N_1210,N_935,N_527);
xor U1211 (N_1211,N_541,N_967);
nand U1212 (N_1212,N_971,N_633);
nand U1213 (N_1213,N_764,N_655);
nor U1214 (N_1214,N_693,N_617);
xor U1215 (N_1215,N_993,N_855);
xnor U1216 (N_1216,N_577,N_538);
nor U1217 (N_1217,N_739,N_982);
xnor U1218 (N_1218,N_591,N_808);
nand U1219 (N_1219,N_856,N_733);
nor U1220 (N_1220,N_727,N_946);
or U1221 (N_1221,N_740,N_781);
nand U1222 (N_1222,N_540,N_851);
nor U1223 (N_1223,N_596,N_580);
and U1224 (N_1224,N_857,N_768);
xor U1225 (N_1225,N_985,N_779);
nand U1226 (N_1226,N_905,N_621);
xor U1227 (N_1227,N_846,N_786);
nor U1228 (N_1228,N_585,N_822);
nor U1229 (N_1229,N_531,N_907);
or U1230 (N_1230,N_648,N_723);
xnor U1231 (N_1231,N_783,N_703);
and U1232 (N_1232,N_756,N_916);
nand U1233 (N_1233,N_923,N_502);
and U1234 (N_1234,N_906,N_533);
nand U1235 (N_1235,N_850,N_710);
or U1236 (N_1236,N_646,N_572);
nor U1237 (N_1237,N_964,N_662);
and U1238 (N_1238,N_717,N_680);
and U1239 (N_1239,N_755,N_721);
and U1240 (N_1240,N_669,N_798);
and U1241 (N_1241,N_989,N_678);
nor U1242 (N_1242,N_941,N_530);
or U1243 (N_1243,N_618,N_877);
and U1244 (N_1244,N_683,N_770);
xor U1245 (N_1245,N_752,N_902);
nand U1246 (N_1246,N_949,N_847);
or U1247 (N_1247,N_885,N_593);
nor U1248 (N_1248,N_823,N_726);
and U1249 (N_1249,N_542,N_995);
nand U1250 (N_1250,N_796,N_558);
and U1251 (N_1251,N_676,N_554);
or U1252 (N_1252,N_904,N_626);
nand U1253 (N_1253,N_645,N_984);
nor U1254 (N_1254,N_842,N_979);
and U1255 (N_1255,N_940,N_893);
nor U1256 (N_1256,N_688,N_526);
xor U1257 (N_1257,N_547,N_529);
nor U1258 (N_1258,N_705,N_533);
nor U1259 (N_1259,N_791,N_700);
or U1260 (N_1260,N_630,N_864);
xor U1261 (N_1261,N_660,N_739);
and U1262 (N_1262,N_777,N_547);
or U1263 (N_1263,N_996,N_984);
or U1264 (N_1264,N_669,N_609);
xor U1265 (N_1265,N_541,N_896);
nor U1266 (N_1266,N_984,N_849);
nor U1267 (N_1267,N_912,N_862);
nor U1268 (N_1268,N_574,N_771);
xor U1269 (N_1269,N_846,N_594);
or U1270 (N_1270,N_914,N_907);
nor U1271 (N_1271,N_848,N_675);
and U1272 (N_1272,N_546,N_729);
nand U1273 (N_1273,N_522,N_917);
nand U1274 (N_1274,N_776,N_688);
nor U1275 (N_1275,N_636,N_601);
and U1276 (N_1276,N_833,N_558);
xnor U1277 (N_1277,N_786,N_644);
and U1278 (N_1278,N_587,N_559);
nor U1279 (N_1279,N_617,N_760);
xnor U1280 (N_1280,N_542,N_985);
and U1281 (N_1281,N_752,N_857);
xor U1282 (N_1282,N_590,N_835);
nor U1283 (N_1283,N_683,N_935);
nor U1284 (N_1284,N_956,N_810);
nor U1285 (N_1285,N_819,N_635);
and U1286 (N_1286,N_910,N_707);
nand U1287 (N_1287,N_911,N_700);
or U1288 (N_1288,N_902,N_726);
nand U1289 (N_1289,N_935,N_825);
nand U1290 (N_1290,N_957,N_784);
nor U1291 (N_1291,N_678,N_631);
xnor U1292 (N_1292,N_587,N_891);
or U1293 (N_1293,N_546,N_754);
or U1294 (N_1294,N_811,N_849);
and U1295 (N_1295,N_811,N_585);
xnor U1296 (N_1296,N_717,N_771);
or U1297 (N_1297,N_613,N_560);
xnor U1298 (N_1298,N_521,N_528);
nand U1299 (N_1299,N_992,N_543);
xor U1300 (N_1300,N_836,N_978);
xor U1301 (N_1301,N_680,N_838);
nand U1302 (N_1302,N_802,N_908);
nor U1303 (N_1303,N_644,N_932);
and U1304 (N_1304,N_607,N_819);
xnor U1305 (N_1305,N_987,N_851);
or U1306 (N_1306,N_544,N_609);
or U1307 (N_1307,N_626,N_964);
nor U1308 (N_1308,N_838,N_628);
and U1309 (N_1309,N_627,N_835);
xor U1310 (N_1310,N_511,N_714);
nand U1311 (N_1311,N_674,N_859);
or U1312 (N_1312,N_913,N_912);
nor U1313 (N_1313,N_504,N_976);
and U1314 (N_1314,N_694,N_837);
or U1315 (N_1315,N_842,N_898);
nand U1316 (N_1316,N_827,N_768);
nor U1317 (N_1317,N_958,N_975);
nand U1318 (N_1318,N_788,N_676);
nor U1319 (N_1319,N_630,N_872);
xnor U1320 (N_1320,N_577,N_833);
nand U1321 (N_1321,N_833,N_506);
nand U1322 (N_1322,N_705,N_854);
and U1323 (N_1323,N_973,N_890);
and U1324 (N_1324,N_619,N_971);
nor U1325 (N_1325,N_555,N_969);
and U1326 (N_1326,N_977,N_948);
or U1327 (N_1327,N_522,N_814);
or U1328 (N_1328,N_972,N_623);
or U1329 (N_1329,N_983,N_576);
nor U1330 (N_1330,N_564,N_892);
xnor U1331 (N_1331,N_579,N_526);
nor U1332 (N_1332,N_993,N_610);
nand U1333 (N_1333,N_644,N_564);
and U1334 (N_1334,N_917,N_799);
or U1335 (N_1335,N_666,N_678);
nand U1336 (N_1336,N_976,N_845);
nand U1337 (N_1337,N_989,N_776);
or U1338 (N_1338,N_672,N_538);
nor U1339 (N_1339,N_521,N_549);
nor U1340 (N_1340,N_748,N_596);
xor U1341 (N_1341,N_742,N_874);
or U1342 (N_1342,N_867,N_844);
nand U1343 (N_1343,N_685,N_964);
and U1344 (N_1344,N_851,N_819);
and U1345 (N_1345,N_610,N_541);
nand U1346 (N_1346,N_550,N_873);
and U1347 (N_1347,N_557,N_789);
and U1348 (N_1348,N_994,N_556);
and U1349 (N_1349,N_942,N_896);
xnor U1350 (N_1350,N_583,N_884);
nor U1351 (N_1351,N_607,N_639);
or U1352 (N_1352,N_718,N_951);
xnor U1353 (N_1353,N_578,N_803);
nor U1354 (N_1354,N_598,N_717);
xor U1355 (N_1355,N_515,N_979);
xnor U1356 (N_1356,N_986,N_782);
nor U1357 (N_1357,N_899,N_550);
nor U1358 (N_1358,N_605,N_869);
xnor U1359 (N_1359,N_696,N_561);
nor U1360 (N_1360,N_536,N_997);
nor U1361 (N_1361,N_539,N_953);
xnor U1362 (N_1362,N_744,N_561);
or U1363 (N_1363,N_810,N_634);
xnor U1364 (N_1364,N_528,N_830);
and U1365 (N_1365,N_736,N_727);
or U1366 (N_1366,N_749,N_546);
or U1367 (N_1367,N_786,N_855);
nand U1368 (N_1368,N_508,N_573);
or U1369 (N_1369,N_580,N_963);
nor U1370 (N_1370,N_681,N_933);
nor U1371 (N_1371,N_953,N_939);
nand U1372 (N_1372,N_723,N_612);
or U1373 (N_1373,N_889,N_687);
and U1374 (N_1374,N_510,N_605);
xor U1375 (N_1375,N_981,N_683);
nor U1376 (N_1376,N_957,N_894);
xor U1377 (N_1377,N_767,N_582);
nand U1378 (N_1378,N_891,N_992);
nor U1379 (N_1379,N_730,N_630);
nand U1380 (N_1380,N_655,N_651);
nand U1381 (N_1381,N_609,N_692);
nand U1382 (N_1382,N_810,N_513);
xnor U1383 (N_1383,N_719,N_935);
and U1384 (N_1384,N_941,N_960);
and U1385 (N_1385,N_947,N_661);
and U1386 (N_1386,N_549,N_935);
or U1387 (N_1387,N_618,N_857);
and U1388 (N_1388,N_851,N_814);
nand U1389 (N_1389,N_674,N_785);
nand U1390 (N_1390,N_852,N_845);
xor U1391 (N_1391,N_615,N_845);
xnor U1392 (N_1392,N_530,N_836);
xor U1393 (N_1393,N_680,N_668);
or U1394 (N_1394,N_623,N_797);
or U1395 (N_1395,N_815,N_953);
or U1396 (N_1396,N_893,N_753);
nand U1397 (N_1397,N_758,N_875);
nor U1398 (N_1398,N_856,N_608);
nor U1399 (N_1399,N_522,N_903);
nand U1400 (N_1400,N_698,N_848);
or U1401 (N_1401,N_675,N_883);
xor U1402 (N_1402,N_747,N_658);
xnor U1403 (N_1403,N_709,N_774);
and U1404 (N_1404,N_726,N_942);
or U1405 (N_1405,N_685,N_794);
nor U1406 (N_1406,N_932,N_738);
and U1407 (N_1407,N_718,N_695);
nand U1408 (N_1408,N_748,N_749);
xnor U1409 (N_1409,N_609,N_561);
or U1410 (N_1410,N_967,N_765);
nor U1411 (N_1411,N_986,N_643);
nor U1412 (N_1412,N_981,N_826);
xor U1413 (N_1413,N_720,N_706);
and U1414 (N_1414,N_863,N_787);
nand U1415 (N_1415,N_507,N_776);
nand U1416 (N_1416,N_744,N_870);
nand U1417 (N_1417,N_771,N_544);
nand U1418 (N_1418,N_846,N_892);
or U1419 (N_1419,N_966,N_723);
nand U1420 (N_1420,N_705,N_902);
nand U1421 (N_1421,N_508,N_675);
xor U1422 (N_1422,N_907,N_624);
or U1423 (N_1423,N_999,N_883);
or U1424 (N_1424,N_778,N_981);
nor U1425 (N_1425,N_764,N_788);
and U1426 (N_1426,N_585,N_632);
and U1427 (N_1427,N_588,N_959);
nand U1428 (N_1428,N_738,N_674);
and U1429 (N_1429,N_961,N_597);
and U1430 (N_1430,N_861,N_950);
nor U1431 (N_1431,N_637,N_596);
or U1432 (N_1432,N_785,N_995);
nor U1433 (N_1433,N_922,N_648);
nor U1434 (N_1434,N_662,N_874);
nand U1435 (N_1435,N_681,N_722);
and U1436 (N_1436,N_875,N_878);
xnor U1437 (N_1437,N_842,N_892);
nor U1438 (N_1438,N_718,N_873);
nand U1439 (N_1439,N_561,N_899);
and U1440 (N_1440,N_818,N_640);
xnor U1441 (N_1441,N_910,N_552);
nand U1442 (N_1442,N_697,N_888);
xor U1443 (N_1443,N_947,N_577);
and U1444 (N_1444,N_907,N_518);
or U1445 (N_1445,N_833,N_925);
xor U1446 (N_1446,N_569,N_592);
and U1447 (N_1447,N_622,N_933);
or U1448 (N_1448,N_780,N_767);
nor U1449 (N_1449,N_563,N_880);
nand U1450 (N_1450,N_607,N_863);
or U1451 (N_1451,N_530,N_827);
xnor U1452 (N_1452,N_730,N_704);
nand U1453 (N_1453,N_962,N_987);
xor U1454 (N_1454,N_906,N_802);
xor U1455 (N_1455,N_691,N_680);
nor U1456 (N_1456,N_551,N_822);
nor U1457 (N_1457,N_781,N_962);
nor U1458 (N_1458,N_592,N_892);
nand U1459 (N_1459,N_774,N_518);
and U1460 (N_1460,N_609,N_764);
and U1461 (N_1461,N_811,N_868);
nand U1462 (N_1462,N_967,N_893);
nor U1463 (N_1463,N_663,N_974);
nand U1464 (N_1464,N_603,N_806);
xnor U1465 (N_1465,N_997,N_649);
xnor U1466 (N_1466,N_754,N_519);
xnor U1467 (N_1467,N_903,N_638);
or U1468 (N_1468,N_814,N_920);
nor U1469 (N_1469,N_742,N_515);
nor U1470 (N_1470,N_577,N_890);
nor U1471 (N_1471,N_607,N_510);
xor U1472 (N_1472,N_514,N_668);
and U1473 (N_1473,N_833,N_663);
or U1474 (N_1474,N_839,N_888);
and U1475 (N_1475,N_641,N_602);
nor U1476 (N_1476,N_640,N_634);
and U1477 (N_1477,N_873,N_857);
nor U1478 (N_1478,N_737,N_788);
nand U1479 (N_1479,N_864,N_661);
nor U1480 (N_1480,N_746,N_559);
nand U1481 (N_1481,N_737,N_574);
nor U1482 (N_1482,N_896,N_603);
or U1483 (N_1483,N_683,N_730);
nand U1484 (N_1484,N_636,N_594);
nor U1485 (N_1485,N_755,N_840);
nand U1486 (N_1486,N_932,N_559);
nand U1487 (N_1487,N_629,N_613);
and U1488 (N_1488,N_535,N_979);
xor U1489 (N_1489,N_873,N_529);
and U1490 (N_1490,N_546,N_932);
xor U1491 (N_1491,N_942,N_548);
or U1492 (N_1492,N_766,N_876);
and U1493 (N_1493,N_628,N_641);
or U1494 (N_1494,N_969,N_831);
nor U1495 (N_1495,N_624,N_640);
and U1496 (N_1496,N_934,N_912);
or U1497 (N_1497,N_903,N_516);
or U1498 (N_1498,N_836,N_636);
and U1499 (N_1499,N_545,N_704);
nor U1500 (N_1500,N_1441,N_1292);
nor U1501 (N_1501,N_1159,N_1415);
nand U1502 (N_1502,N_1240,N_1016);
and U1503 (N_1503,N_1022,N_1008);
or U1504 (N_1504,N_1066,N_1107);
nor U1505 (N_1505,N_1295,N_1336);
or U1506 (N_1506,N_1084,N_1301);
and U1507 (N_1507,N_1327,N_1053);
xnor U1508 (N_1508,N_1223,N_1451);
and U1509 (N_1509,N_1179,N_1438);
or U1510 (N_1510,N_1421,N_1333);
nand U1511 (N_1511,N_1461,N_1472);
or U1512 (N_1512,N_1483,N_1235);
nand U1513 (N_1513,N_1044,N_1102);
or U1514 (N_1514,N_1152,N_1145);
or U1515 (N_1515,N_1028,N_1458);
or U1516 (N_1516,N_1432,N_1116);
nand U1517 (N_1517,N_1471,N_1436);
or U1518 (N_1518,N_1250,N_1137);
nand U1519 (N_1519,N_1479,N_1229);
xor U1520 (N_1520,N_1157,N_1495);
or U1521 (N_1521,N_1004,N_1334);
or U1522 (N_1522,N_1218,N_1249);
or U1523 (N_1523,N_1193,N_1474);
xor U1524 (N_1524,N_1040,N_1306);
xnor U1525 (N_1525,N_1353,N_1352);
or U1526 (N_1526,N_1307,N_1076);
and U1527 (N_1527,N_1287,N_1389);
xnor U1528 (N_1528,N_1175,N_1452);
nor U1529 (N_1529,N_1164,N_1330);
nor U1530 (N_1530,N_1363,N_1395);
nor U1531 (N_1531,N_1455,N_1464);
or U1532 (N_1532,N_1026,N_1337);
and U1533 (N_1533,N_1125,N_1408);
nand U1534 (N_1534,N_1232,N_1124);
xnor U1535 (N_1535,N_1132,N_1372);
and U1536 (N_1536,N_1380,N_1282);
nand U1537 (N_1537,N_1067,N_1156);
nor U1538 (N_1538,N_1216,N_1423);
and U1539 (N_1539,N_1106,N_1196);
nand U1540 (N_1540,N_1104,N_1001);
xnor U1541 (N_1541,N_1447,N_1412);
nand U1542 (N_1542,N_1148,N_1168);
xor U1543 (N_1543,N_1414,N_1043);
and U1544 (N_1544,N_1222,N_1362);
nand U1545 (N_1545,N_1042,N_1058);
nand U1546 (N_1546,N_1254,N_1169);
or U1547 (N_1547,N_1392,N_1069);
nand U1548 (N_1548,N_1129,N_1335);
nand U1549 (N_1549,N_1142,N_1101);
nand U1550 (N_1550,N_1338,N_1258);
nand U1551 (N_1551,N_1271,N_1018);
and U1552 (N_1552,N_1417,N_1002);
nand U1553 (N_1553,N_1439,N_1093);
nor U1554 (N_1554,N_1329,N_1313);
and U1555 (N_1555,N_1041,N_1300);
xor U1556 (N_1556,N_1375,N_1099);
nand U1557 (N_1557,N_1165,N_1138);
and U1558 (N_1558,N_1314,N_1082);
or U1559 (N_1559,N_1317,N_1344);
or U1560 (N_1560,N_1115,N_1469);
nor U1561 (N_1561,N_1114,N_1476);
xor U1562 (N_1562,N_1005,N_1089);
nor U1563 (N_1563,N_1341,N_1063);
nand U1564 (N_1564,N_1224,N_1091);
nor U1565 (N_1565,N_1209,N_1266);
or U1566 (N_1566,N_1297,N_1387);
or U1567 (N_1567,N_1012,N_1396);
xor U1568 (N_1568,N_1413,N_1398);
xnor U1569 (N_1569,N_1025,N_1096);
nand U1570 (N_1570,N_1397,N_1326);
xor U1571 (N_1571,N_1355,N_1298);
nor U1572 (N_1572,N_1290,N_1094);
xor U1573 (N_1573,N_1068,N_1368);
xnor U1574 (N_1574,N_1202,N_1460);
nor U1575 (N_1575,N_1299,N_1260);
and U1576 (N_1576,N_1331,N_1303);
xnor U1577 (N_1577,N_1081,N_1146);
nor U1578 (N_1578,N_1225,N_1324);
nor U1579 (N_1579,N_1172,N_1228);
xnor U1580 (N_1580,N_1493,N_1286);
xnor U1581 (N_1581,N_1070,N_1230);
and U1582 (N_1582,N_1238,N_1236);
nand U1583 (N_1583,N_1251,N_1090);
or U1584 (N_1584,N_1021,N_1373);
and U1585 (N_1585,N_1377,N_1374);
nor U1586 (N_1586,N_1348,N_1247);
or U1587 (N_1587,N_1477,N_1003);
nor U1588 (N_1588,N_1219,N_1481);
and U1589 (N_1589,N_1088,N_1231);
or U1590 (N_1590,N_1265,N_1204);
or U1591 (N_1591,N_1079,N_1369);
and U1592 (N_1592,N_1178,N_1391);
nor U1593 (N_1593,N_1029,N_1205);
xor U1594 (N_1594,N_1035,N_1478);
and U1595 (N_1595,N_1015,N_1055);
nand U1596 (N_1596,N_1416,N_1288);
xor U1597 (N_1597,N_1241,N_1083);
xnor U1598 (N_1598,N_1210,N_1130);
xnor U1599 (N_1599,N_1098,N_1147);
and U1600 (N_1600,N_1234,N_1281);
nor U1601 (N_1601,N_1456,N_1381);
nand U1602 (N_1602,N_1267,N_1332);
and U1603 (N_1603,N_1459,N_1047);
nand U1604 (N_1604,N_1182,N_1302);
or U1605 (N_1605,N_1486,N_1166);
nand U1606 (N_1606,N_1401,N_1211);
nand U1607 (N_1607,N_1346,N_1194);
xnor U1608 (N_1608,N_1468,N_1140);
or U1609 (N_1609,N_1402,N_1061);
nor U1610 (N_1610,N_1033,N_1122);
nor U1611 (N_1611,N_1113,N_1126);
and U1612 (N_1612,N_1394,N_1197);
nor U1613 (N_1613,N_1188,N_1428);
or U1614 (N_1614,N_1074,N_1463);
nand U1615 (N_1615,N_1246,N_1499);
nor U1616 (N_1616,N_1273,N_1162);
xnor U1617 (N_1617,N_1268,N_1127);
nand U1618 (N_1618,N_1252,N_1328);
nand U1619 (N_1619,N_1285,N_1470);
xor U1620 (N_1620,N_1272,N_1426);
or U1621 (N_1621,N_1195,N_1347);
nand U1622 (N_1622,N_1430,N_1110);
and U1623 (N_1623,N_1131,N_1085);
or U1624 (N_1624,N_1013,N_1027);
nor U1625 (N_1625,N_1345,N_1045);
nor U1626 (N_1626,N_1259,N_1108);
and U1627 (N_1627,N_1060,N_1278);
and U1628 (N_1628,N_1453,N_1019);
nor U1629 (N_1629,N_1057,N_1358);
and U1630 (N_1630,N_1242,N_1233);
and U1631 (N_1631,N_1201,N_1404);
xor U1632 (N_1632,N_1444,N_1189);
or U1633 (N_1633,N_1489,N_1289);
or U1634 (N_1634,N_1457,N_1312);
or U1635 (N_1635,N_1220,N_1192);
xor U1636 (N_1636,N_1462,N_1118);
xor U1637 (N_1637,N_1212,N_1245);
nor U1638 (N_1638,N_1150,N_1440);
xor U1639 (N_1639,N_1429,N_1186);
nand U1640 (N_1640,N_1181,N_1139);
or U1641 (N_1641,N_1318,N_1466);
nand U1642 (N_1642,N_1171,N_1121);
and U1643 (N_1643,N_1308,N_1160);
or U1644 (N_1644,N_1445,N_1161);
nand U1645 (N_1645,N_1239,N_1354);
and U1646 (N_1646,N_1071,N_1274);
xor U1647 (N_1647,N_1151,N_1092);
or U1648 (N_1648,N_1385,N_1010);
or U1649 (N_1649,N_1420,N_1153);
xnor U1650 (N_1650,N_1497,N_1384);
nor U1651 (N_1651,N_1050,N_1134);
nand U1652 (N_1652,N_1255,N_1325);
nor U1653 (N_1653,N_1418,N_1062);
and U1654 (N_1654,N_1262,N_1080);
nand U1655 (N_1655,N_1304,N_1073);
and U1656 (N_1656,N_1422,N_1097);
or U1657 (N_1657,N_1437,N_1263);
nand U1658 (N_1658,N_1487,N_1103);
xnor U1659 (N_1659,N_1149,N_1185);
nand U1660 (N_1660,N_1320,N_1128);
xor U1661 (N_1661,N_1244,N_1275);
xnor U1662 (N_1662,N_1490,N_1227);
nand U1663 (N_1663,N_1356,N_1410);
and U1664 (N_1664,N_1279,N_1064);
nand U1665 (N_1665,N_1494,N_1078);
nand U1666 (N_1666,N_1388,N_1133);
xnor U1667 (N_1667,N_1120,N_1180);
nor U1668 (N_1668,N_1020,N_1480);
nor U1669 (N_1669,N_1361,N_1383);
and U1670 (N_1670,N_1434,N_1293);
nand U1671 (N_1671,N_1379,N_1277);
or U1672 (N_1672,N_1054,N_1340);
xor U1673 (N_1673,N_1370,N_1492);
xor U1674 (N_1674,N_1427,N_1177);
and U1675 (N_1675,N_1316,N_1167);
nand U1676 (N_1676,N_1403,N_1339);
nor U1677 (N_1677,N_1376,N_1399);
nand U1678 (N_1678,N_1400,N_1498);
nor U1679 (N_1679,N_1009,N_1111);
or U1680 (N_1680,N_1206,N_1184);
nor U1681 (N_1681,N_1024,N_1243);
and U1682 (N_1682,N_1419,N_1390);
and U1683 (N_1683,N_1046,N_1357);
and U1684 (N_1684,N_1170,N_1207);
and U1685 (N_1685,N_1321,N_1269);
or U1686 (N_1686,N_1039,N_1311);
or U1687 (N_1687,N_1109,N_1284);
or U1688 (N_1688,N_1208,N_1248);
nor U1689 (N_1689,N_1261,N_1237);
or U1690 (N_1690,N_1023,N_1032);
nand U1691 (N_1691,N_1409,N_1296);
or U1692 (N_1692,N_1256,N_1393);
and U1693 (N_1693,N_1049,N_1488);
xnor U1694 (N_1694,N_1112,N_1482);
nand U1695 (N_1695,N_1264,N_1433);
or U1696 (N_1696,N_1359,N_1117);
and U1697 (N_1697,N_1349,N_1496);
nand U1698 (N_1698,N_1123,N_1011);
nor U1699 (N_1699,N_1473,N_1309);
nand U1700 (N_1700,N_1214,N_1425);
xnor U1701 (N_1701,N_1382,N_1305);
xnor U1702 (N_1702,N_1037,N_1014);
or U1703 (N_1703,N_1052,N_1283);
or U1704 (N_1704,N_1367,N_1100);
and U1705 (N_1705,N_1360,N_1351);
xor U1706 (N_1706,N_1176,N_1454);
xnor U1707 (N_1707,N_1484,N_1141);
nor U1708 (N_1708,N_1365,N_1407);
and U1709 (N_1709,N_1294,N_1031);
nor U1710 (N_1710,N_1217,N_1143);
nand U1711 (N_1711,N_1036,N_1000);
nor U1712 (N_1712,N_1007,N_1077);
and U1713 (N_1713,N_1072,N_1190);
xnor U1714 (N_1714,N_1411,N_1350);
nand U1715 (N_1715,N_1135,N_1203);
nor U1716 (N_1716,N_1405,N_1030);
nand U1717 (N_1717,N_1270,N_1276);
or U1718 (N_1718,N_1343,N_1280);
and U1719 (N_1719,N_1448,N_1017);
xnor U1720 (N_1720,N_1065,N_1174);
nand U1721 (N_1721,N_1406,N_1191);
or U1722 (N_1722,N_1087,N_1442);
and U1723 (N_1723,N_1155,N_1291);
nand U1724 (N_1724,N_1215,N_1173);
nor U1725 (N_1725,N_1465,N_1034);
nor U1726 (N_1726,N_1485,N_1200);
nand U1727 (N_1727,N_1475,N_1467);
and U1728 (N_1728,N_1006,N_1221);
nor U1729 (N_1729,N_1213,N_1136);
nand U1730 (N_1730,N_1386,N_1154);
or U1731 (N_1731,N_1051,N_1144);
or U1732 (N_1732,N_1491,N_1105);
or U1733 (N_1733,N_1443,N_1323);
nor U1734 (N_1734,N_1366,N_1319);
and U1735 (N_1735,N_1163,N_1095);
xnor U1736 (N_1736,N_1253,N_1257);
nor U1737 (N_1737,N_1199,N_1075);
or U1738 (N_1738,N_1086,N_1322);
xnor U1739 (N_1739,N_1342,N_1435);
nand U1740 (N_1740,N_1424,N_1198);
xor U1741 (N_1741,N_1431,N_1450);
and U1742 (N_1742,N_1449,N_1119);
nor U1743 (N_1743,N_1378,N_1310);
nor U1744 (N_1744,N_1315,N_1056);
xor U1745 (N_1745,N_1371,N_1226);
nor U1746 (N_1746,N_1187,N_1158);
or U1747 (N_1747,N_1364,N_1446);
and U1748 (N_1748,N_1059,N_1183);
nor U1749 (N_1749,N_1038,N_1048);
nand U1750 (N_1750,N_1498,N_1382);
nand U1751 (N_1751,N_1217,N_1089);
xor U1752 (N_1752,N_1106,N_1382);
or U1753 (N_1753,N_1253,N_1369);
nand U1754 (N_1754,N_1181,N_1369);
nor U1755 (N_1755,N_1132,N_1375);
nand U1756 (N_1756,N_1430,N_1454);
nor U1757 (N_1757,N_1003,N_1270);
xnor U1758 (N_1758,N_1178,N_1476);
xnor U1759 (N_1759,N_1334,N_1139);
or U1760 (N_1760,N_1386,N_1057);
or U1761 (N_1761,N_1005,N_1045);
and U1762 (N_1762,N_1243,N_1172);
nor U1763 (N_1763,N_1426,N_1408);
nor U1764 (N_1764,N_1407,N_1245);
xor U1765 (N_1765,N_1464,N_1012);
nand U1766 (N_1766,N_1053,N_1019);
nand U1767 (N_1767,N_1253,N_1147);
xor U1768 (N_1768,N_1415,N_1220);
or U1769 (N_1769,N_1211,N_1339);
nor U1770 (N_1770,N_1491,N_1283);
and U1771 (N_1771,N_1119,N_1359);
nand U1772 (N_1772,N_1427,N_1170);
or U1773 (N_1773,N_1393,N_1274);
or U1774 (N_1774,N_1126,N_1170);
nand U1775 (N_1775,N_1496,N_1400);
nor U1776 (N_1776,N_1189,N_1432);
or U1777 (N_1777,N_1191,N_1200);
and U1778 (N_1778,N_1030,N_1128);
or U1779 (N_1779,N_1444,N_1251);
nand U1780 (N_1780,N_1479,N_1373);
nor U1781 (N_1781,N_1034,N_1397);
nand U1782 (N_1782,N_1045,N_1090);
xor U1783 (N_1783,N_1215,N_1272);
nor U1784 (N_1784,N_1300,N_1012);
or U1785 (N_1785,N_1357,N_1077);
xor U1786 (N_1786,N_1129,N_1302);
or U1787 (N_1787,N_1079,N_1019);
and U1788 (N_1788,N_1108,N_1104);
and U1789 (N_1789,N_1468,N_1365);
or U1790 (N_1790,N_1407,N_1002);
nand U1791 (N_1791,N_1409,N_1404);
nor U1792 (N_1792,N_1243,N_1038);
xnor U1793 (N_1793,N_1480,N_1408);
or U1794 (N_1794,N_1317,N_1287);
xnor U1795 (N_1795,N_1041,N_1019);
nand U1796 (N_1796,N_1485,N_1213);
or U1797 (N_1797,N_1065,N_1146);
or U1798 (N_1798,N_1338,N_1028);
and U1799 (N_1799,N_1257,N_1270);
and U1800 (N_1800,N_1442,N_1093);
and U1801 (N_1801,N_1359,N_1327);
nand U1802 (N_1802,N_1162,N_1241);
nand U1803 (N_1803,N_1115,N_1321);
nand U1804 (N_1804,N_1065,N_1393);
nor U1805 (N_1805,N_1208,N_1323);
and U1806 (N_1806,N_1260,N_1324);
or U1807 (N_1807,N_1319,N_1380);
nand U1808 (N_1808,N_1082,N_1078);
xnor U1809 (N_1809,N_1189,N_1456);
nor U1810 (N_1810,N_1329,N_1308);
or U1811 (N_1811,N_1360,N_1386);
and U1812 (N_1812,N_1291,N_1054);
and U1813 (N_1813,N_1475,N_1363);
and U1814 (N_1814,N_1221,N_1331);
xor U1815 (N_1815,N_1215,N_1065);
and U1816 (N_1816,N_1114,N_1390);
xor U1817 (N_1817,N_1263,N_1019);
and U1818 (N_1818,N_1038,N_1146);
nand U1819 (N_1819,N_1116,N_1322);
xor U1820 (N_1820,N_1412,N_1244);
and U1821 (N_1821,N_1250,N_1291);
and U1822 (N_1822,N_1144,N_1382);
and U1823 (N_1823,N_1377,N_1056);
or U1824 (N_1824,N_1115,N_1422);
and U1825 (N_1825,N_1348,N_1043);
nor U1826 (N_1826,N_1380,N_1039);
nor U1827 (N_1827,N_1040,N_1354);
xnor U1828 (N_1828,N_1471,N_1324);
xnor U1829 (N_1829,N_1005,N_1324);
or U1830 (N_1830,N_1022,N_1000);
nor U1831 (N_1831,N_1100,N_1417);
nand U1832 (N_1832,N_1004,N_1450);
xor U1833 (N_1833,N_1378,N_1046);
and U1834 (N_1834,N_1063,N_1237);
and U1835 (N_1835,N_1191,N_1309);
xnor U1836 (N_1836,N_1001,N_1408);
or U1837 (N_1837,N_1306,N_1478);
nand U1838 (N_1838,N_1390,N_1025);
nor U1839 (N_1839,N_1460,N_1247);
or U1840 (N_1840,N_1268,N_1052);
or U1841 (N_1841,N_1451,N_1358);
and U1842 (N_1842,N_1169,N_1266);
xor U1843 (N_1843,N_1410,N_1119);
and U1844 (N_1844,N_1429,N_1480);
nand U1845 (N_1845,N_1086,N_1165);
or U1846 (N_1846,N_1213,N_1284);
xnor U1847 (N_1847,N_1259,N_1265);
or U1848 (N_1848,N_1372,N_1369);
nor U1849 (N_1849,N_1301,N_1136);
nor U1850 (N_1850,N_1147,N_1278);
or U1851 (N_1851,N_1493,N_1181);
and U1852 (N_1852,N_1167,N_1433);
nor U1853 (N_1853,N_1064,N_1036);
nand U1854 (N_1854,N_1471,N_1222);
nor U1855 (N_1855,N_1066,N_1361);
nand U1856 (N_1856,N_1075,N_1448);
or U1857 (N_1857,N_1288,N_1424);
and U1858 (N_1858,N_1381,N_1110);
xor U1859 (N_1859,N_1059,N_1362);
nand U1860 (N_1860,N_1382,N_1434);
xor U1861 (N_1861,N_1137,N_1083);
nand U1862 (N_1862,N_1028,N_1125);
or U1863 (N_1863,N_1332,N_1106);
xor U1864 (N_1864,N_1168,N_1377);
or U1865 (N_1865,N_1034,N_1003);
xnor U1866 (N_1866,N_1393,N_1207);
or U1867 (N_1867,N_1385,N_1035);
nand U1868 (N_1868,N_1285,N_1208);
and U1869 (N_1869,N_1012,N_1340);
xor U1870 (N_1870,N_1283,N_1339);
and U1871 (N_1871,N_1266,N_1101);
or U1872 (N_1872,N_1199,N_1215);
or U1873 (N_1873,N_1466,N_1178);
nand U1874 (N_1874,N_1365,N_1354);
or U1875 (N_1875,N_1367,N_1357);
nor U1876 (N_1876,N_1038,N_1160);
xor U1877 (N_1877,N_1309,N_1419);
and U1878 (N_1878,N_1063,N_1013);
nor U1879 (N_1879,N_1479,N_1392);
nand U1880 (N_1880,N_1280,N_1085);
nand U1881 (N_1881,N_1061,N_1443);
and U1882 (N_1882,N_1111,N_1323);
xor U1883 (N_1883,N_1092,N_1174);
nor U1884 (N_1884,N_1072,N_1320);
nor U1885 (N_1885,N_1232,N_1359);
or U1886 (N_1886,N_1376,N_1456);
and U1887 (N_1887,N_1266,N_1315);
or U1888 (N_1888,N_1083,N_1253);
nand U1889 (N_1889,N_1213,N_1292);
nand U1890 (N_1890,N_1169,N_1069);
nand U1891 (N_1891,N_1429,N_1073);
or U1892 (N_1892,N_1179,N_1166);
nand U1893 (N_1893,N_1114,N_1267);
xnor U1894 (N_1894,N_1452,N_1370);
or U1895 (N_1895,N_1212,N_1100);
nand U1896 (N_1896,N_1327,N_1362);
nand U1897 (N_1897,N_1272,N_1051);
and U1898 (N_1898,N_1236,N_1216);
or U1899 (N_1899,N_1065,N_1415);
nor U1900 (N_1900,N_1415,N_1184);
nand U1901 (N_1901,N_1319,N_1099);
nand U1902 (N_1902,N_1286,N_1428);
nor U1903 (N_1903,N_1007,N_1099);
nor U1904 (N_1904,N_1300,N_1297);
or U1905 (N_1905,N_1059,N_1180);
nand U1906 (N_1906,N_1013,N_1047);
and U1907 (N_1907,N_1372,N_1053);
nand U1908 (N_1908,N_1488,N_1212);
and U1909 (N_1909,N_1331,N_1422);
or U1910 (N_1910,N_1196,N_1088);
and U1911 (N_1911,N_1130,N_1235);
xor U1912 (N_1912,N_1208,N_1458);
nand U1913 (N_1913,N_1192,N_1352);
xor U1914 (N_1914,N_1268,N_1024);
or U1915 (N_1915,N_1053,N_1473);
or U1916 (N_1916,N_1236,N_1409);
or U1917 (N_1917,N_1366,N_1010);
and U1918 (N_1918,N_1363,N_1053);
xnor U1919 (N_1919,N_1249,N_1321);
xor U1920 (N_1920,N_1264,N_1358);
and U1921 (N_1921,N_1341,N_1379);
xnor U1922 (N_1922,N_1085,N_1250);
xnor U1923 (N_1923,N_1329,N_1493);
nand U1924 (N_1924,N_1413,N_1466);
and U1925 (N_1925,N_1416,N_1207);
and U1926 (N_1926,N_1154,N_1437);
nor U1927 (N_1927,N_1046,N_1196);
and U1928 (N_1928,N_1014,N_1015);
xnor U1929 (N_1929,N_1350,N_1163);
nand U1930 (N_1930,N_1186,N_1480);
and U1931 (N_1931,N_1049,N_1239);
nor U1932 (N_1932,N_1055,N_1290);
and U1933 (N_1933,N_1060,N_1294);
nand U1934 (N_1934,N_1075,N_1030);
nor U1935 (N_1935,N_1181,N_1344);
nor U1936 (N_1936,N_1069,N_1495);
and U1937 (N_1937,N_1346,N_1315);
nand U1938 (N_1938,N_1492,N_1219);
xnor U1939 (N_1939,N_1055,N_1393);
or U1940 (N_1940,N_1174,N_1295);
nor U1941 (N_1941,N_1236,N_1458);
nor U1942 (N_1942,N_1446,N_1015);
nor U1943 (N_1943,N_1318,N_1146);
xor U1944 (N_1944,N_1260,N_1309);
and U1945 (N_1945,N_1453,N_1433);
or U1946 (N_1946,N_1474,N_1391);
xor U1947 (N_1947,N_1367,N_1421);
and U1948 (N_1948,N_1078,N_1017);
and U1949 (N_1949,N_1093,N_1389);
nand U1950 (N_1950,N_1340,N_1001);
or U1951 (N_1951,N_1104,N_1451);
or U1952 (N_1952,N_1325,N_1389);
and U1953 (N_1953,N_1165,N_1275);
and U1954 (N_1954,N_1499,N_1428);
nor U1955 (N_1955,N_1391,N_1330);
and U1956 (N_1956,N_1137,N_1369);
and U1957 (N_1957,N_1475,N_1087);
nand U1958 (N_1958,N_1475,N_1438);
xor U1959 (N_1959,N_1106,N_1162);
or U1960 (N_1960,N_1274,N_1455);
nand U1961 (N_1961,N_1281,N_1089);
and U1962 (N_1962,N_1082,N_1128);
xor U1963 (N_1963,N_1487,N_1446);
and U1964 (N_1964,N_1497,N_1429);
nand U1965 (N_1965,N_1114,N_1276);
nand U1966 (N_1966,N_1186,N_1453);
nor U1967 (N_1967,N_1398,N_1218);
and U1968 (N_1968,N_1485,N_1340);
nor U1969 (N_1969,N_1199,N_1062);
nor U1970 (N_1970,N_1377,N_1368);
and U1971 (N_1971,N_1360,N_1237);
or U1972 (N_1972,N_1247,N_1163);
xor U1973 (N_1973,N_1352,N_1312);
or U1974 (N_1974,N_1144,N_1288);
xor U1975 (N_1975,N_1338,N_1198);
nand U1976 (N_1976,N_1229,N_1194);
nand U1977 (N_1977,N_1155,N_1462);
xor U1978 (N_1978,N_1378,N_1220);
xnor U1979 (N_1979,N_1216,N_1494);
or U1980 (N_1980,N_1489,N_1229);
or U1981 (N_1981,N_1308,N_1224);
nand U1982 (N_1982,N_1429,N_1070);
nand U1983 (N_1983,N_1402,N_1333);
nor U1984 (N_1984,N_1488,N_1351);
xnor U1985 (N_1985,N_1206,N_1420);
xnor U1986 (N_1986,N_1426,N_1141);
nand U1987 (N_1987,N_1222,N_1127);
nor U1988 (N_1988,N_1159,N_1018);
nor U1989 (N_1989,N_1293,N_1236);
xnor U1990 (N_1990,N_1026,N_1388);
nand U1991 (N_1991,N_1395,N_1438);
and U1992 (N_1992,N_1022,N_1075);
or U1993 (N_1993,N_1199,N_1281);
xor U1994 (N_1994,N_1123,N_1245);
xnor U1995 (N_1995,N_1309,N_1139);
nor U1996 (N_1996,N_1195,N_1278);
nand U1997 (N_1997,N_1239,N_1247);
nor U1998 (N_1998,N_1292,N_1076);
xnor U1999 (N_1999,N_1372,N_1314);
or U2000 (N_2000,N_1884,N_1620);
nor U2001 (N_2001,N_1778,N_1731);
xnor U2002 (N_2002,N_1513,N_1627);
or U2003 (N_2003,N_1548,N_1775);
nor U2004 (N_2004,N_1827,N_1857);
xor U2005 (N_2005,N_1754,N_1546);
and U2006 (N_2006,N_1647,N_1804);
nand U2007 (N_2007,N_1583,N_1988);
nor U2008 (N_2008,N_1985,N_1738);
or U2009 (N_2009,N_1830,N_1862);
nand U2010 (N_2010,N_1734,N_1605);
nand U2011 (N_2011,N_1685,N_1616);
nand U2012 (N_2012,N_1611,N_1791);
nor U2013 (N_2013,N_1562,N_1649);
and U2014 (N_2014,N_1765,N_1746);
nor U2015 (N_2015,N_1809,N_1690);
and U2016 (N_2016,N_1969,N_1593);
and U2017 (N_2017,N_1828,N_1903);
nor U2018 (N_2018,N_1590,N_1766);
or U2019 (N_2019,N_1912,N_1522);
nand U2020 (N_2020,N_1956,N_1661);
or U2021 (N_2021,N_1859,N_1878);
nand U2022 (N_2022,N_1640,N_1626);
and U2023 (N_2023,N_1994,N_1952);
and U2024 (N_2024,N_1686,N_1713);
nor U2025 (N_2025,N_1904,N_1675);
or U2026 (N_2026,N_1561,N_1960);
and U2027 (N_2027,N_1719,N_1648);
and U2028 (N_2028,N_1907,N_1650);
or U2029 (N_2029,N_1813,N_1573);
or U2030 (N_2030,N_1992,N_1806);
or U2031 (N_2031,N_1564,N_1659);
and U2032 (N_2032,N_1625,N_1964);
nand U2033 (N_2033,N_1824,N_1705);
and U2034 (N_2034,N_1788,N_1787);
xnor U2035 (N_2035,N_1744,N_1505);
xnor U2036 (N_2036,N_1785,N_1883);
nand U2037 (N_2037,N_1727,N_1945);
and U2038 (N_2038,N_1818,N_1556);
nand U2039 (N_2039,N_1540,N_1973);
or U2040 (N_2040,N_1702,N_1831);
or U2041 (N_2041,N_1846,N_1608);
or U2042 (N_2042,N_1998,N_1684);
xnor U2043 (N_2043,N_1925,N_1643);
xor U2044 (N_2044,N_1936,N_1800);
nand U2045 (N_2045,N_1689,N_1624);
xnor U2046 (N_2046,N_1595,N_1970);
nand U2047 (N_2047,N_1968,N_1697);
and U2048 (N_2048,N_1929,N_1858);
nand U2049 (N_2049,N_1639,N_1550);
xor U2050 (N_2050,N_1645,N_1844);
nor U2051 (N_2051,N_1959,N_1981);
and U2052 (N_2052,N_1826,N_1676);
nor U2053 (N_2053,N_1515,N_1655);
xnor U2054 (N_2054,N_1946,N_1758);
and U2055 (N_2055,N_1617,N_1773);
or U2056 (N_2056,N_1810,N_1926);
xor U2057 (N_2057,N_1591,N_1779);
nand U2058 (N_2058,N_1716,N_1602);
or U2059 (N_2059,N_1874,N_1918);
and U2060 (N_2060,N_1641,N_1833);
xnor U2061 (N_2061,N_1500,N_1604);
or U2062 (N_2062,N_1993,N_1563);
xor U2063 (N_2063,N_1701,N_1569);
xnor U2064 (N_2064,N_1843,N_1967);
and U2065 (N_2065,N_1978,N_1769);
and U2066 (N_2066,N_1948,N_1750);
or U2067 (N_2067,N_1721,N_1951);
and U2068 (N_2068,N_1603,N_1802);
and U2069 (N_2069,N_1877,N_1632);
nor U2070 (N_2070,N_1555,N_1980);
xnor U2071 (N_2071,N_1572,N_1982);
and U2072 (N_2072,N_1635,N_1658);
nor U2073 (N_2073,N_1847,N_1733);
nor U2074 (N_2074,N_1782,N_1710);
and U2075 (N_2075,N_1911,N_1558);
xnor U2076 (N_2076,N_1977,N_1580);
and U2077 (N_2077,N_1966,N_1680);
nor U2078 (N_2078,N_1694,N_1614);
xor U2079 (N_2079,N_1720,N_1509);
nor U2080 (N_2080,N_1983,N_1607);
and U2081 (N_2081,N_1913,N_1881);
and U2082 (N_2082,N_1792,N_1871);
nor U2083 (N_2083,N_1629,N_1693);
xnor U2084 (N_2084,N_1610,N_1514);
or U2085 (N_2085,N_1503,N_1814);
and U2086 (N_2086,N_1866,N_1707);
nor U2087 (N_2087,N_1681,N_1906);
xnor U2088 (N_2088,N_1533,N_1527);
and U2089 (N_2089,N_1708,N_1501);
and U2090 (N_2090,N_1660,N_1816);
and U2091 (N_2091,N_1612,N_1762);
and U2092 (N_2092,N_1714,N_1891);
xnor U2093 (N_2093,N_1835,N_1803);
or U2094 (N_2094,N_1520,N_1875);
nor U2095 (N_2095,N_1999,N_1772);
xor U2096 (N_2096,N_1848,N_1979);
nand U2097 (N_2097,N_1905,N_1896);
and U2098 (N_2098,N_1751,N_1609);
and U2099 (N_2099,N_1971,N_1799);
or U2100 (N_2100,N_1972,N_1776);
nor U2101 (N_2101,N_1886,N_1837);
or U2102 (N_2102,N_1990,N_1718);
or U2103 (N_2103,N_1790,N_1667);
and U2104 (N_2104,N_1834,N_1613);
and U2105 (N_2105,N_1670,N_1922);
or U2106 (N_2106,N_1786,N_1728);
and U2107 (N_2107,N_1674,N_1856);
xor U2108 (N_2108,N_1691,N_1914);
xnor U2109 (N_2109,N_1724,N_1579);
or U2110 (N_2110,N_1943,N_1975);
xnor U2111 (N_2111,N_1717,N_1600);
and U2112 (N_2112,N_1642,N_1568);
nor U2113 (N_2113,N_1656,N_1901);
xor U2114 (N_2114,N_1927,N_1822);
or U2115 (N_2115,N_1506,N_1794);
and U2116 (N_2116,N_1736,N_1745);
and U2117 (N_2117,N_1811,N_1598);
and U2118 (N_2118,N_1618,N_1991);
xor U2119 (N_2119,N_1666,N_1698);
nor U2120 (N_2120,N_1832,N_1938);
xor U2121 (N_2121,N_1541,N_1545);
or U2122 (N_2122,N_1796,N_1920);
or U2123 (N_2123,N_1654,N_1517);
nor U2124 (N_2124,N_1863,N_1899);
nor U2125 (N_2125,N_1829,N_1588);
nand U2126 (N_2126,N_1567,N_1543);
nor U2127 (N_2127,N_1930,N_1537);
and U2128 (N_2128,N_1931,N_1849);
xnor U2129 (N_2129,N_1646,N_1795);
nor U2130 (N_2130,N_1557,N_1512);
nand U2131 (N_2131,N_1673,N_1547);
or U2132 (N_2132,N_1840,N_1711);
or U2133 (N_2133,N_1651,N_1730);
or U2134 (N_2134,N_1934,N_1759);
nand U2135 (N_2135,N_1551,N_1633);
or U2136 (N_2136,N_1908,N_1757);
nand U2137 (N_2137,N_1984,N_1542);
nor U2138 (N_2138,N_1735,N_1574);
and U2139 (N_2139,N_1688,N_1560);
nor U2140 (N_2140,N_1669,N_1783);
xor U2141 (N_2141,N_1909,N_1836);
xnor U2142 (N_2142,N_1887,N_1737);
or U2143 (N_2143,N_1861,N_1663);
or U2144 (N_2144,N_1808,N_1894);
or U2145 (N_2145,N_1784,N_1882);
and U2146 (N_2146,N_1867,N_1644);
and U2147 (N_2147,N_1665,N_1578);
nand U2148 (N_2148,N_1987,N_1662);
nor U2149 (N_2149,N_1854,N_1622);
or U2150 (N_2150,N_1630,N_1636);
or U2151 (N_2151,N_1531,N_1774);
and U2152 (N_2152,N_1823,N_1584);
xor U2153 (N_2153,N_1864,N_1544);
or U2154 (N_2154,N_1812,N_1763);
or U2155 (N_2155,N_1534,N_1652);
xor U2156 (N_2156,N_1853,N_1789);
and U2157 (N_2157,N_1671,N_1915);
nor U2158 (N_2158,N_1825,N_1923);
or U2159 (N_2159,N_1621,N_1860);
or U2160 (N_2160,N_1585,N_1932);
xor U2161 (N_2161,N_1937,N_1725);
and U2162 (N_2162,N_1741,N_1756);
xor U2163 (N_2163,N_1597,N_1890);
and U2164 (N_2164,N_1615,N_1703);
nand U2165 (N_2165,N_1963,N_1530);
nand U2166 (N_2166,N_1753,N_1582);
xnor U2167 (N_2167,N_1781,N_1510);
or U2168 (N_2168,N_1897,N_1526);
and U2169 (N_2169,N_1965,N_1594);
or U2170 (N_2170,N_1596,N_1538);
or U2171 (N_2171,N_1748,N_1895);
or U2172 (N_2172,N_1755,N_1672);
and U2173 (N_2173,N_1589,N_1957);
nor U2174 (N_2174,N_1525,N_1687);
nor U2175 (N_2175,N_1521,N_1700);
or U2176 (N_2176,N_1518,N_1511);
and U2177 (N_2177,N_1601,N_1577);
or U2178 (N_2178,N_1761,N_1706);
nand U2179 (N_2179,N_1723,N_1869);
nor U2180 (N_2180,N_1732,N_1868);
nor U2181 (N_2181,N_1516,N_1553);
nor U2182 (N_2182,N_1910,N_1628);
nor U2183 (N_2183,N_1587,N_1872);
nand U2184 (N_2184,N_1696,N_1815);
nand U2185 (N_2185,N_1508,N_1528);
and U2186 (N_2186,N_1851,N_1532);
and U2187 (N_2187,N_1668,N_1954);
and U2188 (N_2188,N_1747,N_1539);
nand U2189 (N_2189,N_1797,N_1892);
xnor U2190 (N_2190,N_1780,N_1638);
or U2191 (N_2191,N_1742,N_1880);
xor U2192 (N_2192,N_1935,N_1599);
xnor U2193 (N_2193,N_1889,N_1683);
and U2194 (N_2194,N_1726,N_1722);
nand U2195 (N_2195,N_1739,N_1677);
nor U2196 (N_2196,N_1850,N_1917);
nor U2197 (N_2197,N_1947,N_1958);
nor U2198 (N_2198,N_1606,N_1933);
or U2199 (N_2199,N_1870,N_1712);
and U2200 (N_2200,N_1950,N_1807);
xnor U2201 (N_2201,N_1502,N_1565);
and U2202 (N_2202,N_1507,N_1549);
xor U2203 (N_2203,N_1821,N_1995);
and U2204 (N_2204,N_1657,N_1819);
and U2205 (N_2205,N_1529,N_1801);
nand U2206 (N_2206,N_1852,N_1519);
xor U2207 (N_2207,N_1879,N_1941);
nor U2208 (N_2208,N_1749,N_1942);
xor U2209 (N_2209,N_1845,N_1841);
nand U2210 (N_2210,N_1898,N_1571);
and U2211 (N_2211,N_1692,N_1928);
and U2212 (N_2212,N_1939,N_1752);
or U2213 (N_2213,N_1523,N_1842);
or U2214 (N_2214,N_1699,N_1623);
and U2215 (N_2215,N_1709,N_1570);
xnor U2216 (N_2216,N_1592,N_1940);
and U2217 (N_2217,N_1634,N_1974);
and U2218 (N_2218,N_1664,N_1949);
or U2219 (N_2219,N_1760,N_1865);
nand U2220 (N_2220,N_1961,N_1777);
or U2221 (N_2221,N_1962,N_1873);
or U2222 (N_2222,N_1885,N_1955);
xor U2223 (N_2223,N_1715,N_1916);
or U2224 (N_2224,N_1924,N_1536);
nor U2225 (N_2225,N_1793,N_1771);
or U2226 (N_2226,N_1919,N_1944);
nor U2227 (N_2227,N_1767,N_1888);
and U2228 (N_2228,N_1552,N_1996);
or U2229 (N_2229,N_1989,N_1900);
nand U2230 (N_2230,N_1876,N_1575);
xor U2231 (N_2231,N_1986,N_1576);
nand U2232 (N_2232,N_1953,N_1704);
and U2233 (N_2233,N_1921,N_1805);
and U2234 (N_2234,N_1619,N_1504);
and U2235 (N_2235,N_1524,N_1695);
and U2236 (N_2236,N_1770,N_1679);
nor U2237 (N_2237,N_1554,N_1740);
nor U2238 (N_2238,N_1768,N_1817);
and U2239 (N_2239,N_1798,N_1535);
or U2240 (N_2240,N_1976,N_1637);
and U2241 (N_2241,N_1566,N_1743);
and U2242 (N_2242,N_1839,N_1586);
and U2243 (N_2243,N_1764,N_1581);
xor U2244 (N_2244,N_1559,N_1997);
and U2245 (N_2245,N_1855,N_1729);
nor U2246 (N_2246,N_1902,N_1893);
nand U2247 (N_2247,N_1631,N_1838);
nand U2248 (N_2248,N_1653,N_1820);
nor U2249 (N_2249,N_1678,N_1682);
nor U2250 (N_2250,N_1981,N_1974);
nand U2251 (N_2251,N_1666,N_1733);
xor U2252 (N_2252,N_1722,N_1811);
xor U2253 (N_2253,N_1952,N_1532);
nor U2254 (N_2254,N_1938,N_1946);
or U2255 (N_2255,N_1652,N_1605);
nand U2256 (N_2256,N_1948,N_1853);
nand U2257 (N_2257,N_1501,N_1995);
nor U2258 (N_2258,N_1891,N_1540);
xor U2259 (N_2259,N_1736,N_1776);
and U2260 (N_2260,N_1858,N_1945);
and U2261 (N_2261,N_1562,N_1825);
and U2262 (N_2262,N_1898,N_1524);
xnor U2263 (N_2263,N_1735,N_1825);
nor U2264 (N_2264,N_1806,N_1769);
and U2265 (N_2265,N_1850,N_1528);
xnor U2266 (N_2266,N_1716,N_1987);
nor U2267 (N_2267,N_1925,N_1799);
or U2268 (N_2268,N_1903,N_1686);
nor U2269 (N_2269,N_1847,N_1884);
xor U2270 (N_2270,N_1922,N_1917);
or U2271 (N_2271,N_1574,N_1776);
xor U2272 (N_2272,N_1660,N_1821);
nand U2273 (N_2273,N_1531,N_1938);
and U2274 (N_2274,N_1673,N_1760);
xor U2275 (N_2275,N_1788,N_1789);
and U2276 (N_2276,N_1705,N_1723);
and U2277 (N_2277,N_1953,N_1538);
xor U2278 (N_2278,N_1615,N_1566);
or U2279 (N_2279,N_1811,N_1829);
or U2280 (N_2280,N_1720,N_1856);
nand U2281 (N_2281,N_1547,N_1821);
nor U2282 (N_2282,N_1570,N_1817);
or U2283 (N_2283,N_1710,N_1745);
nor U2284 (N_2284,N_1857,N_1858);
nor U2285 (N_2285,N_1739,N_1572);
xor U2286 (N_2286,N_1596,N_1558);
nand U2287 (N_2287,N_1732,N_1695);
nor U2288 (N_2288,N_1800,N_1899);
nor U2289 (N_2289,N_1842,N_1604);
nor U2290 (N_2290,N_1884,N_1646);
nor U2291 (N_2291,N_1601,N_1639);
nor U2292 (N_2292,N_1906,N_1926);
xnor U2293 (N_2293,N_1827,N_1948);
nor U2294 (N_2294,N_1575,N_1661);
nor U2295 (N_2295,N_1833,N_1871);
xor U2296 (N_2296,N_1939,N_1542);
nand U2297 (N_2297,N_1764,N_1906);
nor U2298 (N_2298,N_1589,N_1537);
and U2299 (N_2299,N_1718,N_1963);
xor U2300 (N_2300,N_1701,N_1542);
xnor U2301 (N_2301,N_1888,N_1797);
or U2302 (N_2302,N_1804,N_1703);
and U2303 (N_2303,N_1828,N_1954);
and U2304 (N_2304,N_1800,N_1549);
nor U2305 (N_2305,N_1627,N_1910);
nand U2306 (N_2306,N_1687,N_1657);
nor U2307 (N_2307,N_1985,N_1583);
or U2308 (N_2308,N_1518,N_1934);
or U2309 (N_2309,N_1707,N_1776);
or U2310 (N_2310,N_1810,N_1973);
or U2311 (N_2311,N_1830,N_1926);
or U2312 (N_2312,N_1988,N_1501);
nand U2313 (N_2313,N_1582,N_1535);
xnor U2314 (N_2314,N_1824,N_1820);
xnor U2315 (N_2315,N_1988,N_1975);
xor U2316 (N_2316,N_1747,N_1903);
or U2317 (N_2317,N_1518,N_1580);
xnor U2318 (N_2318,N_1731,N_1797);
and U2319 (N_2319,N_1957,N_1929);
nand U2320 (N_2320,N_1848,N_1830);
nor U2321 (N_2321,N_1844,N_1629);
nor U2322 (N_2322,N_1962,N_1628);
xor U2323 (N_2323,N_1551,N_1721);
or U2324 (N_2324,N_1781,N_1504);
nand U2325 (N_2325,N_1530,N_1817);
nor U2326 (N_2326,N_1552,N_1780);
nor U2327 (N_2327,N_1904,N_1829);
nor U2328 (N_2328,N_1970,N_1515);
nor U2329 (N_2329,N_1843,N_1829);
nor U2330 (N_2330,N_1591,N_1862);
nand U2331 (N_2331,N_1735,N_1647);
nand U2332 (N_2332,N_1763,N_1528);
nand U2333 (N_2333,N_1554,N_1771);
nor U2334 (N_2334,N_1583,N_1969);
or U2335 (N_2335,N_1560,N_1521);
nand U2336 (N_2336,N_1801,N_1745);
and U2337 (N_2337,N_1955,N_1933);
and U2338 (N_2338,N_1545,N_1776);
or U2339 (N_2339,N_1739,N_1933);
and U2340 (N_2340,N_1759,N_1575);
nor U2341 (N_2341,N_1736,N_1986);
or U2342 (N_2342,N_1795,N_1590);
nand U2343 (N_2343,N_1992,N_1501);
or U2344 (N_2344,N_1822,N_1750);
nor U2345 (N_2345,N_1755,N_1591);
xnor U2346 (N_2346,N_1988,N_1898);
or U2347 (N_2347,N_1931,N_1746);
or U2348 (N_2348,N_1631,N_1713);
and U2349 (N_2349,N_1745,N_1598);
or U2350 (N_2350,N_1638,N_1988);
or U2351 (N_2351,N_1539,N_1964);
xor U2352 (N_2352,N_1578,N_1939);
nor U2353 (N_2353,N_1991,N_1921);
xnor U2354 (N_2354,N_1818,N_1906);
xnor U2355 (N_2355,N_1604,N_1641);
and U2356 (N_2356,N_1518,N_1761);
and U2357 (N_2357,N_1791,N_1923);
nor U2358 (N_2358,N_1621,N_1807);
or U2359 (N_2359,N_1624,N_1733);
nand U2360 (N_2360,N_1785,N_1597);
nand U2361 (N_2361,N_1616,N_1933);
or U2362 (N_2362,N_1861,N_1546);
xnor U2363 (N_2363,N_1577,N_1608);
and U2364 (N_2364,N_1713,N_1958);
and U2365 (N_2365,N_1555,N_1999);
nor U2366 (N_2366,N_1607,N_1741);
nor U2367 (N_2367,N_1992,N_1900);
and U2368 (N_2368,N_1857,N_1923);
or U2369 (N_2369,N_1780,N_1569);
or U2370 (N_2370,N_1719,N_1525);
and U2371 (N_2371,N_1558,N_1671);
nor U2372 (N_2372,N_1633,N_1506);
nand U2373 (N_2373,N_1812,N_1628);
and U2374 (N_2374,N_1677,N_1844);
nand U2375 (N_2375,N_1996,N_1724);
nand U2376 (N_2376,N_1952,N_1650);
and U2377 (N_2377,N_1895,N_1873);
or U2378 (N_2378,N_1670,N_1552);
xnor U2379 (N_2379,N_1942,N_1720);
and U2380 (N_2380,N_1664,N_1563);
and U2381 (N_2381,N_1837,N_1923);
or U2382 (N_2382,N_1880,N_1903);
xnor U2383 (N_2383,N_1632,N_1542);
nor U2384 (N_2384,N_1907,N_1979);
xnor U2385 (N_2385,N_1802,N_1990);
nand U2386 (N_2386,N_1917,N_1921);
and U2387 (N_2387,N_1695,N_1751);
or U2388 (N_2388,N_1632,N_1620);
or U2389 (N_2389,N_1541,N_1975);
nand U2390 (N_2390,N_1728,N_1794);
or U2391 (N_2391,N_1982,N_1642);
nor U2392 (N_2392,N_1938,N_1508);
nor U2393 (N_2393,N_1805,N_1880);
or U2394 (N_2394,N_1813,N_1994);
or U2395 (N_2395,N_1933,N_1848);
nand U2396 (N_2396,N_1846,N_1573);
xnor U2397 (N_2397,N_1501,N_1827);
or U2398 (N_2398,N_1772,N_1839);
and U2399 (N_2399,N_1737,N_1842);
and U2400 (N_2400,N_1903,N_1996);
nor U2401 (N_2401,N_1589,N_1701);
xor U2402 (N_2402,N_1640,N_1771);
or U2403 (N_2403,N_1848,N_1542);
nor U2404 (N_2404,N_1967,N_1918);
nand U2405 (N_2405,N_1698,N_1500);
or U2406 (N_2406,N_1757,N_1889);
nor U2407 (N_2407,N_1946,N_1557);
nand U2408 (N_2408,N_1593,N_1547);
xor U2409 (N_2409,N_1843,N_1643);
xor U2410 (N_2410,N_1533,N_1926);
nand U2411 (N_2411,N_1583,N_1718);
or U2412 (N_2412,N_1953,N_1571);
nand U2413 (N_2413,N_1942,N_1507);
xor U2414 (N_2414,N_1632,N_1696);
nor U2415 (N_2415,N_1520,N_1773);
xor U2416 (N_2416,N_1777,N_1841);
or U2417 (N_2417,N_1603,N_1766);
xnor U2418 (N_2418,N_1804,N_1905);
nand U2419 (N_2419,N_1515,N_1888);
nor U2420 (N_2420,N_1997,N_1531);
nor U2421 (N_2421,N_1870,N_1521);
or U2422 (N_2422,N_1561,N_1634);
or U2423 (N_2423,N_1949,N_1692);
nor U2424 (N_2424,N_1883,N_1514);
and U2425 (N_2425,N_1578,N_1727);
nand U2426 (N_2426,N_1864,N_1712);
or U2427 (N_2427,N_1904,N_1670);
xor U2428 (N_2428,N_1848,N_1662);
nand U2429 (N_2429,N_1556,N_1917);
xor U2430 (N_2430,N_1909,N_1885);
and U2431 (N_2431,N_1720,N_1991);
and U2432 (N_2432,N_1800,N_1676);
nor U2433 (N_2433,N_1575,N_1803);
and U2434 (N_2434,N_1806,N_1860);
nand U2435 (N_2435,N_1866,N_1867);
nor U2436 (N_2436,N_1939,N_1993);
nor U2437 (N_2437,N_1968,N_1825);
nand U2438 (N_2438,N_1657,N_1921);
or U2439 (N_2439,N_1522,N_1963);
nor U2440 (N_2440,N_1720,N_1630);
or U2441 (N_2441,N_1754,N_1713);
or U2442 (N_2442,N_1635,N_1999);
and U2443 (N_2443,N_1853,N_1906);
nand U2444 (N_2444,N_1896,N_1713);
xnor U2445 (N_2445,N_1616,N_1560);
nand U2446 (N_2446,N_1861,N_1930);
nor U2447 (N_2447,N_1606,N_1557);
or U2448 (N_2448,N_1507,N_1666);
xnor U2449 (N_2449,N_1612,N_1557);
or U2450 (N_2450,N_1798,N_1879);
nand U2451 (N_2451,N_1809,N_1754);
and U2452 (N_2452,N_1858,N_1533);
and U2453 (N_2453,N_1735,N_1949);
or U2454 (N_2454,N_1697,N_1874);
nor U2455 (N_2455,N_1866,N_1608);
or U2456 (N_2456,N_1833,N_1620);
nand U2457 (N_2457,N_1545,N_1792);
and U2458 (N_2458,N_1669,N_1901);
xnor U2459 (N_2459,N_1626,N_1914);
nor U2460 (N_2460,N_1514,N_1973);
and U2461 (N_2461,N_1693,N_1927);
and U2462 (N_2462,N_1636,N_1503);
nand U2463 (N_2463,N_1941,N_1734);
nor U2464 (N_2464,N_1587,N_1920);
nand U2465 (N_2465,N_1741,N_1963);
nand U2466 (N_2466,N_1833,N_1522);
nand U2467 (N_2467,N_1719,N_1796);
or U2468 (N_2468,N_1579,N_1916);
and U2469 (N_2469,N_1762,N_1692);
nor U2470 (N_2470,N_1783,N_1623);
nor U2471 (N_2471,N_1714,N_1967);
or U2472 (N_2472,N_1731,N_1908);
nor U2473 (N_2473,N_1644,N_1625);
nand U2474 (N_2474,N_1650,N_1773);
or U2475 (N_2475,N_1940,N_1967);
xor U2476 (N_2476,N_1870,N_1593);
and U2477 (N_2477,N_1590,N_1813);
nand U2478 (N_2478,N_1649,N_1948);
or U2479 (N_2479,N_1979,N_1502);
nand U2480 (N_2480,N_1560,N_1693);
nor U2481 (N_2481,N_1524,N_1910);
or U2482 (N_2482,N_1699,N_1502);
nand U2483 (N_2483,N_1804,N_1780);
nand U2484 (N_2484,N_1869,N_1718);
xnor U2485 (N_2485,N_1780,N_1590);
nor U2486 (N_2486,N_1827,N_1848);
nand U2487 (N_2487,N_1805,N_1762);
and U2488 (N_2488,N_1664,N_1944);
nand U2489 (N_2489,N_1977,N_1547);
or U2490 (N_2490,N_1967,N_1764);
nand U2491 (N_2491,N_1788,N_1899);
xor U2492 (N_2492,N_1529,N_1686);
nand U2493 (N_2493,N_1542,N_1882);
nor U2494 (N_2494,N_1774,N_1619);
and U2495 (N_2495,N_1778,N_1543);
xor U2496 (N_2496,N_1798,N_1773);
nand U2497 (N_2497,N_1909,N_1625);
xor U2498 (N_2498,N_1990,N_1684);
nand U2499 (N_2499,N_1524,N_1614);
and U2500 (N_2500,N_2077,N_2187);
or U2501 (N_2501,N_2194,N_2450);
nor U2502 (N_2502,N_2211,N_2462);
xnor U2503 (N_2503,N_2089,N_2029);
nor U2504 (N_2504,N_2488,N_2276);
nor U2505 (N_2505,N_2304,N_2205);
and U2506 (N_2506,N_2197,N_2442);
nand U2507 (N_2507,N_2421,N_2107);
nor U2508 (N_2508,N_2141,N_2299);
and U2509 (N_2509,N_2114,N_2380);
or U2510 (N_2510,N_2310,N_2127);
nand U2511 (N_2511,N_2149,N_2035);
and U2512 (N_2512,N_2398,N_2013);
and U2513 (N_2513,N_2212,N_2484);
xnor U2514 (N_2514,N_2167,N_2108);
xor U2515 (N_2515,N_2243,N_2447);
and U2516 (N_2516,N_2102,N_2278);
and U2517 (N_2517,N_2349,N_2277);
or U2518 (N_2518,N_2483,N_2291);
nand U2519 (N_2519,N_2423,N_2021);
nand U2520 (N_2520,N_2088,N_2409);
xnor U2521 (N_2521,N_2361,N_2174);
nand U2522 (N_2522,N_2461,N_2069);
nand U2523 (N_2523,N_2455,N_2377);
and U2524 (N_2524,N_2147,N_2078);
and U2525 (N_2525,N_2416,N_2001);
nor U2526 (N_2526,N_2287,N_2363);
nand U2527 (N_2527,N_2010,N_2360);
and U2528 (N_2528,N_2378,N_2262);
xor U2529 (N_2529,N_2312,N_2414);
xor U2530 (N_2530,N_2123,N_2148);
nand U2531 (N_2531,N_2240,N_2048);
nor U2532 (N_2532,N_2324,N_2269);
nor U2533 (N_2533,N_2237,N_2456);
nand U2534 (N_2534,N_2444,N_2096);
nand U2535 (N_2535,N_2161,N_2176);
nor U2536 (N_2536,N_2028,N_2224);
nand U2537 (N_2537,N_2087,N_2449);
xor U2538 (N_2538,N_2375,N_2045);
nor U2539 (N_2539,N_2352,N_2079);
and U2540 (N_2540,N_2027,N_2284);
nor U2541 (N_2541,N_2266,N_2286);
nand U2542 (N_2542,N_2439,N_2471);
xor U2543 (N_2543,N_2465,N_2156);
xor U2544 (N_2544,N_2334,N_2393);
and U2545 (N_2545,N_2175,N_2158);
nand U2546 (N_2546,N_2358,N_2374);
nor U2547 (N_2547,N_2204,N_2384);
and U2548 (N_2548,N_2343,N_2353);
or U2549 (N_2549,N_2354,N_2301);
nor U2550 (N_2550,N_2101,N_2184);
and U2551 (N_2551,N_2056,N_2073);
and U2552 (N_2552,N_2064,N_2259);
nor U2553 (N_2553,N_2281,N_2136);
or U2554 (N_2554,N_2189,N_2081);
and U2555 (N_2555,N_2402,N_2198);
xor U2556 (N_2556,N_2459,N_2083);
xor U2557 (N_2557,N_2411,N_2248);
xnor U2558 (N_2558,N_2494,N_2199);
or U2559 (N_2559,N_2196,N_2124);
and U2560 (N_2560,N_2043,N_2115);
and U2561 (N_2561,N_2121,N_2093);
and U2562 (N_2562,N_2366,N_2231);
and U2563 (N_2563,N_2020,N_2009);
nor U2564 (N_2564,N_2249,N_2368);
nor U2565 (N_2565,N_2475,N_2213);
and U2566 (N_2566,N_2033,N_2234);
nand U2567 (N_2567,N_2319,N_2162);
or U2568 (N_2568,N_2091,N_2433);
or U2569 (N_2569,N_2489,N_2422);
xor U2570 (N_2570,N_2216,N_2195);
and U2571 (N_2571,N_2235,N_2372);
or U2572 (N_2572,N_2007,N_2206);
nand U2573 (N_2573,N_2133,N_2347);
xnor U2574 (N_2574,N_2453,N_2344);
nor U2575 (N_2575,N_2496,N_2024);
nand U2576 (N_2576,N_2185,N_2247);
nor U2577 (N_2577,N_2221,N_2082);
xor U2578 (N_2578,N_2467,N_2332);
nand U2579 (N_2579,N_2061,N_2367);
and U2580 (N_2580,N_2164,N_2267);
or U2581 (N_2581,N_2057,N_2296);
nor U2582 (N_2582,N_2392,N_2431);
nor U2583 (N_2583,N_2341,N_2111);
and U2584 (N_2584,N_2053,N_2445);
nor U2585 (N_2585,N_2457,N_2118);
and U2586 (N_2586,N_2345,N_2292);
xnor U2587 (N_2587,N_2413,N_2289);
nand U2588 (N_2588,N_2389,N_2298);
nor U2589 (N_2589,N_2485,N_2207);
xnor U2590 (N_2590,N_2321,N_2381);
xor U2591 (N_2591,N_2160,N_2498);
or U2592 (N_2592,N_2443,N_2113);
xor U2593 (N_2593,N_2428,N_2151);
or U2594 (N_2594,N_2364,N_2138);
nand U2595 (N_2595,N_2327,N_2255);
and U2596 (N_2596,N_2331,N_2210);
nand U2597 (N_2597,N_2408,N_2290);
or U2598 (N_2598,N_2186,N_2282);
or U2599 (N_2599,N_2429,N_2309);
and U2600 (N_2600,N_2018,N_2351);
xor U2601 (N_2601,N_2337,N_2085);
or U2602 (N_2602,N_2106,N_2242);
and U2603 (N_2603,N_2265,N_2190);
or U2604 (N_2604,N_2066,N_2239);
nand U2605 (N_2605,N_2365,N_2168);
nand U2606 (N_2606,N_2094,N_2244);
nand U2607 (N_2607,N_2068,N_2371);
and U2608 (N_2608,N_2335,N_2464);
nand U2609 (N_2609,N_2328,N_2050);
nand U2610 (N_2610,N_2256,N_2359);
or U2611 (N_2611,N_2006,N_2300);
and U2612 (N_2612,N_2280,N_2410);
and U2613 (N_2613,N_2135,N_2223);
xor U2614 (N_2614,N_2140,N_2474);
or U2615 (N_2615,N_2209,N_2193);
and U2616 (N_2616,N_2131,N_2323);
nor U2617 (N_2617,N_2454,N_2070);
xor U2618 (N_2618,N_2178,N_2480);
xor U2619 (N_2619,N_2188,N_2487);
or U2620 (N_2620,N_2143,N_2095);
and U2621 (N_2621,N_2134,N_2037);
or U2622 (N_2622,N_2306,N_2017);
nand U2623 (N_2623,N_2023,N_2369);
and U2624 (N_2624,N_2192,N_2099);
nor U2625 (N_2625,N_2499,N_2258);
xor U2626 (N_2626,N_2448,N_2452);
or U2627 (N_2627,N_2038,N_2391);
xnor U2628 (N_2628,N_2318,N_2217);
xor U2629 (N_2629,N_2002,N_2424);
xor U2630 (N_2630,N_2036,N_2051);
xor U2631 (N_2631,N_2098,N_2003);
nor U2632 (N_2632,N_2418,N_2376);
nand U2633 (N_2633,N_2202,N_2104);
nand U2634 (N_2634,N_2288,N_2152);
and U2635 (N_2635,N_2400,N_2092);
nor U2636 (N_2636,N_2451,N_2263);
nor U2637 (N_2637,N_2072,N_2463);
nand U2638 (N_2638,N_2016,N_2316);
or U2639 (N_2639,N_2407,N_2420);
or U2640 (N_2640,N_2103,N_2435);
and U2641 (N_2641,N_2307,N_2159);
and U2642 (N_2642,N_2271,N_2097);
or U2643 (N_2643,N_2170,N_2157);
nand U2644 (N_2644,N_2294,N_2226);
and U2645 (N_2645,N_2330,N_2283);
nor U2646 (N_2646,N_2386,N_2490);
and U2647 (N_2647,N_2139,N_2019);
nor U2648 (N_2648,N_2419,N_2075);
nand U2649 (N_2649,N_2253,N_2026);
nor U2650 (N_2650,N_2426,N_2339);
nand U2651 (N_2651,N_2396,N_2394);
nor U2652 (N_2652,N_2236,N_2432);
xor U2653 (N_2653,N_2275,N_2220);
nand U2654 (N_2654,N_2116,N_2179);
xor U2655 (N_2655,N_2145,N_2401);
nand U2656 (N_2656,N_2071,N_2491);
or U2657 (N_2657,N_2183,N_2122);
nand U2658 (N_2658,N_2142,N_2434);
nand U2659 (N_2659,N_2025,N_2273);
nand U2660 (N_2660,N_2405,N_2387);
nand U2661 (N_2661,N_2150,N_2350);
and U2662 (N_2662,N_2356,N_2427);
and U2663 (N_2663,N_2065,N_2305);
nor U2664 (N_2664,N_2482,N_2246);
or U2665 (N_2665,N_2117,N_2203);
and U2666 (N_2666,N_2446,N_2479);
nand U2667 (N_2667,N_2302,N_2497);
and U2668 (N_2668,N_2060,N_2348);
and U2669 (N_2669,N_2279,N_2132);
nand U2670 (N_2670,N_2342,N_2052);
and U2671 (N_2671,N_2336,N_2466);
and U2672 (N_2672,N_2397,N_2425);
nor U2673 (N_2673,N_2146,N_2406);
xor U2674 (N_2674,N_2412,N_2214);
or U2675 (N_2675,N_2308,N_2100);
nor U2676 (N_2676,N_2493,N_2090);
or U2677 (N_2677,N_2208,N_2333);
nor U2678 (N_2678,N_2005,N_2062);
nor U2679 (N_2679,N_2272,N_2254);
nand U2680 (N_2680,N_2233,N_2441);
or U2681 (N_2681,N_2125,N_2163);
nand U2682 (N_2682,N_2251,N_2346);
xor U2683 (N_2683,N_2313,N_2268);
xnor U2684 (N_2684,N_2382,N_2201);
nand U2685 (N_2685,N_2225,N_2458);
and U2686 (N_2686,N_2477,N_2469);
or U2687 (N_2687,N_2171,N_2270);
nor U2688 (N_2688,N_2227,N_2034);
or U2689 (N_2689,N_2044,N_2370);
nor U2690 (N_2690,N_2438,N_2440);
xor U2691 (N_2691,N_2297,N_2388);
nor U2692 (N_2692,N_2200,N_2495);
xnor U2693 (N_2693,N_2076,N_2385);
and U2694 (N_2694,N_2074,N_2063);
xor U2695 (N_2695,N_2436,N_2230);
nor U2696 (N_2696,N_2067,N_2228);
nand U2697 (N_2697,N_2481,N_2031);
or U2698 (N_2698,N_2177,N_2165);
nor U2699 (N_2699,N_2059,N_2395);
nand U2700 (N_2700,N_2112,N_2215);
nand U2701 (N_2701,N_2362,N_2460);
nand U2702 (N_2702,N_2169,N_2144);
nor U2703 (N_2703,N_2218,N_2229);
nand U2704 (N_2704,N_2172,N_2417);
nand U2705 (N_2705,N_2084,N_2014);
xnor U2706 (N_2706,N_2478,N_2315);
xnor U2707 (N_2707,N_2264,N_2015);
or U2708 (N_2708,N_2390,N_2430);
and U2709 (N_2709,N_2011,N_2238);
nand U2710 (N_2710,N_2154,N_2004);
nand U2711 (N_2711,N_2041,N_2317);
nor U2712 (N_2712,N_2252,N_2415);
and U2713 (N_2713,N_2293,N_2022);
nand U2714 (N_2714,N_2379,N_2054);
and U2715 (N_2715,N_2049,N_2329);
or U2716 (N_2716,N_2008,N_2047);
nand U2717 (N_2717,N_2325,N_2080);
nor U2718 (N_2718,N_2314,N_2399);
and U2719 (N_2719,N_2357,N_2285);
and U2720 (N_2720,N_2320,N_2295);
and U2721 (N_2721,N_2404,N_2241);
and U2722 (N_2722,N_2109,N_2338);
xnor U2723 (N_2723,N_2486,N_2470);
xnor U2724 (N_2724,N_2126,N_2303);
nor U2725 (N_2725,N_2472,N_2166);
nor U2726 (N_2726,N_2000,N_2222);
nand U2727 (N_2727,N_2110,N_2245);
xor U2728 (N_2728,N_2120,N_2274);
xor U2729 (N_2729,N_2191,N_2130);
nor U2730 (N_2730,N_2232,N_2119);
nand U2731 (N_2731,N_2340,N_2181);
or U2732 (N_2732,N_2492,N_2155);
nand U2733 (N_2733,N_2403,N_2153);
nor U2734 (N_2734,N_2129,N_2032);
nand U2735 (N_2735,N_2086,N_2257);
nor U2736 (N_2736,N_2355,N_2311);
and U2737 (N_2737,N_2173,N_2219);
or U2738 (N_2738,N_2039,N_2046);
nor U2739 (N_2739,N_2326,N_2030);
and U2740 (N_2740,N_2058,N_2473);
or U2741 (N_2741,N_2137,N_2437);
and U2742 (N_2742,N_2040,N_2128);
nor U2743 (N_2743,N_2250,N_2042);
nor U2744 (N_2744,N_2261,N_2373);
and U2745 (N_2745,N_2012,N_2182);
or U2746 (N_2746,N_2383,N_2322);
nand U2747 (N_2747,N_2476,N_2105);
and U2748 (N_2748,N_2260,N_2468);
or U2749 (N_2749,N_2180,N_2055);
xnor U2750 (N_2750,N_2343,N_2294);
xor U2751 (N_2751,N_2138,N_2127);
xor U2752 (N_2752,N_2290,N_2073);
nand U2753 (N_2753,N_2408,N_2388);
nand U2754 (N_2754,N_2191,N_2430);
xnor U2755 (N_2755,N_2141,N_2382);
and U2756 (N_2756,N_2447,N_2241);
xor U2757 (N_2757,N_2322,N_2271);
xor U2758 (N_2758,N_2103,N_2022);
xnor U2759 (N_2759,N_2258,N_2024);
and U2760 (N_2760,N_2204,N_2295);
nor U2761 (N_2761,N_2294,N_2231);
and U2762 (N_2762,N_2405,N_2267);
nor U2763 (N_2763,N_2438,N_2126);
nor U2764 (N_2764,N_2218,N_2217);
xnor U2765 (N_2765,N_2425,N_2298);
or U2766 (N_2766,N_2197,N_2299);
or U2767 (N_2767,N_2000,N_2325);
and U2768 (N_2768,N_2024,N_2105);
nand U2769 (N_2769,N_2273,N_2444);
or U2770 (N_2770,N_2401,N_2192);
and U2771 (N_2771,N_2205,N_2253);
or U2772 (N_2772,N_2342,N_2353);
and U2773 (N_2773,N_2141,N_2206);
xnor U2774 (N_2774,N_2108,N_2137);
xnor U2775 (N_2775,N_2445,N_2267);
nor U2776 (N_2776,N_2141,N_2459);
nand U2777 (N_2777,N_2312,N_2046);
nor U2778 (N_2778,N_2377,N_2146);
or U2779 (N_2779,N_2329,N_2361);
xnor U2780 (N_2780,N_2210,N_2004);
nand U2781 (N_2781,N_2041,N_2204);
xor U2782 (N_2782,N_2226,N_2135);
xnor U2783 (N_2783,N_2444,N_2392);
nand U2784 (N_2784,N_2418,N_2401);
nand U2785 (N_2785,N_2485,N_2208);
nor U2786 (N_2786,N_2370,N_2454);
or U2787 (N_2787,N_2021,N_2113);
and U2788 (N_2788,N_2066,N_2339);
xor U2789 (N_2789,N_2331,N_2232);
and U2790 (N_2790,N_2058,N_2290);
xor U2791 (N_2791,N_2240,N_2010);
xnor U2792 (N_2792,N_2322,N_2220);
nand U2793 (N_2793,N_2257,N_2320);
or U2794 (N_2794,N_2408,N_2059);
nand U2795 (N_2795,N_2196,N_2468);
and U2796 (N_2796,N_2492,N_2427);
nand U2797 (N_2797,N_2354,N_2487);
xor U2798 (N_2798,N_2365,N_2103);
or U2799 (N_2799,N_2039,N_2000);
nor U2800 (N_2800,N_2364,N_2348);
and U2801 (N_2801,N_2286,N_2260);
xor U2802 (N_2802,N_2417,N_2407);
and U2803 (N_2803,N_2139,N_2170);
and U2804 (N_2804,N_2259,N_2320);
or U2805 (N_2805,N_2469,N_2096);
or U2806 (N_2806,N_2108,N_2332);
and U2807 (N_2807,N_2310,N_2249);
or U2808 (N_2808,N_2186,N_2161);
and U2809 (N_2809,N_2038,N_2095);
or U2810 (N_2810,N_2276,N_2477);
and U2811 (N_2811,N_2446,N_2164);
and U2812 (N_2812,N_2125,N_2093);
nand U2813 (N_2813,N_2104,N_2417);
nand U2814 (N_2814,N_2051,N_2479);
or U2815 (N_2815,N_2269,N_2225);
or U2816 (N_2816,N_2390,N_2034);
xnor U2817 (N_2817,N_2330,N_2174);
or U2818 (N_2818,N_2405,N_2444);
and U2819 (N_2819,N_2251,N_2075);
nand U2820 (N_2820,N_2200,N_2335);
nor U2821 (N_2821,N_2102,N_2094);
nand U2822 (N_2822,N_2456,N_2160);
nor U2823 (N_2823,N_2185,N_2419);
or U2824 (N_2824,N_2258,N_2447);
nand U2825 (N_2825,N_2046,N_2241);
or U2826 (N_2826,N_2045,N_2010);
and U2827 (N_2827,N_2178,N_2283);
nand U2828 (N_2828,N_2205,N_2069);
xnor U2829 (N_2829,N_2407,N_2218);
nand U2830 (N_2830,N_2043,N_2012);
xnor U2831 (N_2831,N_2171,N_2184);
or U2832 (N_2832,N_2248,N_2377);
and U2833 (N_2833,N_2312,N_2197);
xor U2834 (N_2834,N_2159,N_2244);
nand U2835 (N_2835,N_2395,N_2477);
or U2836 (N_2836,N_2435,N_2260);
nor U2837 (N_2837,N_2004,N_2014);
or U2838 (N_2838,N_2069,N_2043);
nor U2839 (N_2839,N_2031,N_2051);
nand U2840 (N_2840,N_2334,N_2359);
nor U2841 (N_2841,N_2077,N_2101);
nor U2842 (N_2842,N_2150,N_2493);
nor U2843 (N_2843,N_2145,N_2000);
nor U2844 (N_2844,N_2346,N_2161);
nand U2845 (N_2845,N_2282,N_2226);
and U2846 (N_2846,N_2351,N_2345);
nand U2847 (N_2847,N_2309,N_2252);
nor U2848 (N_2848,N_2030,N_2308);
nand U2849 (N_2849,N_2260,N_2492);
nand U2850 (N_2850,N_2406,N_2486);
nand U2851 (N_2851,N_2007,N_2031);
and U2852 (N_2852,N_2496,N_2365);
and U2853 (N_2853,N_2484,N_2130);
xnor U2854 (N_2854,N_2350,N_2009);
nand U2855 (N_2855,N_2412,N_2064);
or U2856 (N_2856,N_2221,N_2106);
or U2857 (N_2857,N_2142,N_2299);
nor U2858 (N_2858,N_2444,N_2351);
nand U2859 (N_2859,N_2370,N_2147);
nor U2860 (N_2860,N_2194,N_2209);
nor U2861 (N_2861,N_2409,N_2413);
nor U2862 (N_2862,N_2428,N_2417);
nor U2863 (N_2863,N_2356,N_2057);
xor U2864 (N_2864,N_2359,N_2164);
xor U2865 (N_2865,N_2080,N_2162);
nor U2866 (N_2866,N_2084,N_2035);
nor U2867 (N_2867,N_2049,N_2067);
xnor U2868 (N_2868,N_2187,N_2170);
nand U2869 (N_2869,N_2167,N_2224);
nor U2870 (N_2870,N_2038,N_2411);
and U2871 (N_2871,N_2200,N_2028);
xor U2872 (N_2872,N_2411,N_2016);
xor U2873 (N_2873,N_2118,N_2027);
xor U2874 (N_2874,N_2073,N_2093);
and U2875 (N_2875,N_2101,N_2367);
or U2876 (N_2876,N_2336,N_2003);
and U2877 (N_2877,N_2484,N_2460);
nand U2878 (N_2878,N_2363,N_2390);
nor U2879 (N_2879,N_2042,N_2444);
or U2880 (N_2880,N_2000,N_2455);
or U2881 (N_2881,N_2468,N_2158);
nand U2882 (N_2882,N_2435,N_2004);
xnor U2883 (N_2883,N_2142,N_2403);
or U2884 (N_2884,N_2329,N_2119);
xor U2885 (N_2885,N_2324,N_2246);
or U2886 (N_2886,N_2462,N_2189);
or U2887 (N_2887,N_2333,N_2088);
and U2888 (N_2888,N_2273,N_2339);
nor U2889 (N_2889,N_2409,N_2288);
and U2890 (N_2890,N_2261,N_2213);
or U2891 (N_2891,N_2007,N_2393);
xnor U2892 (N_2892,N_2332,N_2088);
xor U2893 (N_2893,N_2434,N_2178);
and U2894 (N_2894,N_2157,N_2276);
and U2895 (N_2895,N_2446,N_2499);
or U2896 (N_2896,N_2269,N_2391);
xnor U2897 (N_2897,N_2481,N_2319);
nand U2898 (N_2898,N_2493,N_2401);
or U2899 (N_2899,N_2439,N_2026);
nor U2900 (N_2900,N_2191,N_2438);
or U2901 (N_2901,N_2243,N_2498);
nand U2902 (N_2902,N_2347,N_2255);
nand U2903 (N_2903,N_2283,N_2449);
nand U2904 (N_2904,N_2154,N_2464);
nand U2905 (N_2905,N_2435,N_2198);
and U2906 (N_2906,N_2200,N_2249);
xnor U2907 (N_2907,N_2495,N_2409);
nand U2908 (N_2908,N_2087,N_2135);
nand U2909 (N_2909,N_2140,N_2373);
and U2910 (N_2910,N_2256,N_2237);
xor U2911 (N_2911,N_2140,N_2039);
nand U2912 (N_2912,N_2104,N_2333);
or U2913 (N_2913,N_2133,N_2346);
xor U2914 (N_2914,N_2037,N_2289);
xnor U2915 (N_2915,N_2463,N_2015);
xnor U2916 (N_2916,N_2453,N_2063);
xnor U2917 (N_2917,N_2394,N_2389);
and U2918 (N_2918,N_2393,N_2442);
nand U2919 (N_2919,N_2243,N_2018);
nand U2920 (N_2920,N_2200,N_2086);
or U2921 (N_2921,N_2081,N_2006);
xnor U2922 (N_2922,N_2185,N_2007);
nand U2923 (N_2923,N_2301,N_2235);
nor U2924 (N_2924,N_2278,N_2045);
nand U2925 (N_2925,N_2206,N_2438);
or U2926 (N_2926,N_2425,N_2272);
or U2927 (N_2927,N_2393,N_2154);
and U2928 (N_2928,N_2102,N_2320);
or U2929 (N_2929,N_2153,N_2055);
nor U2930 (N_2930,N_2137,N_2059);
and U2931 (N_2931,N_2219,N_2167);
or U2932 (N_2932,N_2472,N_2494);
xor U2933 (N_2933,N_2369,N_2408);
nand U2934 (N_2934,N_2314,N_2076);
nor U2935 (N_2935,N_2168,N_2095);
or U2936 (N_2936,N_2053,N_2156);
nor U2937 (N_2937,N_2234,N_2174);
xor U2938 (N_2938,N_2490,N_2400);
nor U2939 (N_2939,N_2078,N_2442);
nor U2940 (N_2940,N_2111,N_2143);
and U2941 (N_2941,N_2491,N_2360);
and U2942 (N_2942,N_2437,N_2268);
and U2943 (N_2943,N_2492,N_2416);
nor U2944 (N_2944,N_2488,N_2044);
and U2945 (N_2945,N_2089,N_2050);
or U2946 (N_2946,N_2255,N_2161);
nand U2947 (N_2947,N_2464,N_2209);
and U2948 (N_2948,N_2032,N_2051);
nand U2949 (N_2949,N_2169,N_2007);
nand U2950 (N_2950,N_2376,N_2006);
nand U2951 (N_2951,N_2026,N_2340);
xor U2952 (N_2952,N_2286,N_2402);
nor U2953 (N_2953,N_2364,N_2091);
or U2954 (N_2954,N_2393,N_2229);
nor U2955 (N_2955,N_2403,N_2303);
and U2956 (N_2956,N_2247,N_2316);
nand U2957 (N_2957,N_2250,N_2452);
or U2958 (N_2958,N_2468,N_2487);
nor U2959 (N_2959,N_2032,N_2222);
or U2960 (N_2960,N_2471,N_2410);
nor U2961 (N_2961,N_2246,N_2445);
and U2962 (N_2962,N_2376,N_2387);
xnor U2963 (N_2963,N_2265,N_2385);
nor U2964 (N_2964,N_2070,N_2439);
nor U2965 (N_2965,N_2414,N_2435);
and U2966 (N_2966,N_2012,N_2014);
xor U2967 (N_2967,N_2387,N_2186);
xnor U2968 (N_2968,N_2152,N_2314);
and U2969 (N_2969,N_2111,N_2060);
nand U2970 (N_2970,N_2475,N_2472);
or U2971 (N_2971,N_2350,N_2345);
xnor U2972 (N_2972,N_2045,N_2296);
nor U2973 (N_2973,N_2002,N_2187);
xor U2974 (N_2974,N_2465,N_2313);
nand U2975 (N_2975,N_2171,N_2428);
nor U2976 (N_2976,N_2195,N_2439);
or U2977 (N_2977,N_2161,N_2340);
nor U2978 (N_2978,N_2229,N_2447);
nand U2979 (N_2979,N_2190,N_2204);
and U2980 (N_2980,N_2402,N_2290);
xnor U2981 (N_2981,N_2261,N_2140);
nor U2982 (N_2982,N_2074,N_2303);
xnor U2983 (N_2983,N_2089,N_2033);
xnor U2984 (N_2984,N_2157,N_2315);
or U2985 (N_2985,N_2383,N_2310);
and U2986 (N_2986,N_2382,N_2438);
xor U2987 (N_2987,N_2145,N_2462);
and U2988 (N_2988,N_2348,N_2425);
and U2989 (N_2989,N_2187,N_2205);
and U2990 (N_2990,N_2185,N_2355);
xnor U2991 (N_2991,N_2307,N_2358);
and U2992 (N_2992,N_2034,N_2167);
xor U2993 (N_2993,N_2296,N_2134);
nor U2994 (N_2994,N_2179,N_2339);
nor U2995 (N_2995,N_2229,N_2284);
and U2996 (N_2996,N_2351,N_2096);
and U2997 (N_2997,N_2144,N_2368);
nand U2998 (N_2998,N_2035,N_2007);
nand U2999 (N_2999,N_2254,N_2396);
and U3000 (N_3000,N_2690,N_2804);
nand U3001 (N_3001,N_2735,N_2964);
xnor U3002 (N_3002,N_2669,N_2889);
nand U3003 (N_3003,N_2558,N_2780);
nand U3004 (N_3004,N_2700,N_2732);
or U3005 (N_3005,N_2525,N_2740);
and U3006 (N_3006,N_2787,N_2881);
xnor U3007 (N_3007,N_2941,N_2693);
xnor U3008 (N_3008,N_2504,N_2500);
nand U3009 (N_3009,N_2791,N_2789);
or U3010 (N_3010,N_2798,N_2619);
nand U3011 (N_3011,N_2710,N_2810);
nor U3012 (N_3012,N_2826,N_2726);
xnor U3013 (N_3013,N_2648,N_2664);
nor U3014 (N_3014,N_2893,N_2679);
or U3015 (N_3015,N_2905,N_2630);
nand U3016 (N_3016,N_2886,N_2501);
xnor U3017 (N_3017,N_2821,N_2784);
nand U3018 (N_3018,N_2622,N_2918);
or U3019 (N_3019,N_2720,N_2706);
or U3020 (N_3020,N_2541,N_2729);
nor U3021 (N_3021,N_2528,N_2951);
or U3022 (N_3022,N_2503,N_2713);
nand U3023 (N_3023,N_2976,N_2639);
or U3024 (N_3024,N_2761,N_2954);
or U3025 (N_3025,N_2590,N_2997);
or U3026 (N_3026,N_2596,N_2862);
xnor U3027 (N_3027,N_2757,N_2717);
xnor U3028 (N_3028,N_2623,N_2513);
xnor U3029 (N_3029,N_2828,N_2745);
nor U3030 (N_3030,N_2545,N_2966);
xor U3031 (N_3031,N_2856,N_2742);
nor U3032 (N_3032,N_2800,N_2666);
nand U3033 (N_3033,N_2988,N_2878);
and U3034 (N_3034,N_2536,N_2860);
xor U3035 (N_3035,N_2896,N_2550);
xnor U3036 (N_3036,N_2831,N_2527);
nor U3037 (N_3037,N_2770,N_2543);
xnor U3038 (N_3038,N_2689,N_2707);
xnor U3039 (N_3039,N_2978,N_2508);
nor U3040 (N_3040,N_2506,N_2743);
and U3041 (N_3041,N_2759,N_2876);
nand U3042 (N_3042,N_2637,N_2792);
nand U3043 (N_3043,N_2645,N_2986);
nand U3044 (N_3044,N_2950,N_2704);
nor U3045 (N_3045,N_2822,N_2939);
and U3046 (N_3046,N_2725,N_2677);
and U3047 (N_3047,N_2942,N_2534);
nand U3048 (N_3048,N_2989,N_2829);
or U3049 (N_3049,N_2892,N_2775);
xor U3050 (N_3050,N_2785,N_2842);
xor U3051 (N_3051,N_2825,N_2540);
xnor U3052 (N_3052,N_2772,N_2620);
nand U3053 (N_3053,N_2934,N_2808);
and U3054 (N_3054,N_2588,N_2994);
nand U3055 (N_3055,N_2511,N_2799);
or U3056 (N_3056,N_2952,N_2882);
and U3057 (N_3057,N_2972,N_2643);
nor U3058 (N_3058,N_2647,N_2510);
or U3059 (N_3059,N_2771,N_2667);
nand U3060 (N_3060,N_2718,N_2533);
nand U3061 (N_3061,N_2701,N_2955);
nor U3062 (N_3062,N_2776,N_2749);
nand U3063 (N_3063,N_2566,N_2613);
or U3064 (N_3064,N_2801,N_2922);
and U3065 (N_3065,N_2849,N_2688);
nor U3066 (N_3066,N_2662,N_2845);
or U3067 (N_3067,N_2968,N_2995);
nand U3068 (N_3068,N_2857,N_2562);
xnor U3069 (N_3069,N_2736,N_2556);
nand U3070 (N_3070,N_2547,N_2817);
xnor U3071 (N_3071,N_2607,N_2908);
and U3072 (N_3072,N_2769,N_2699);
nand U3073 (N_3073,N_2575,N_2595);
xnor U3074 (N_3074,N_2778,N_2609);
or U3075 (N_3075,N_2919,N_2832);
xnor U3076 (N_3076,N_2820,N_2601);
nand U3077 (N_3077,N_2879,N_2658);
nor U3078 (N_3078,N_2549,N_2577);
and U3079 (N_3079,N_2616,N_2844);
and U3080 (N_3080,N_2923,N_2611);
nand U3081 (N_3081,N_2962,N_2873);
xor U3082 (N_3082,N_2910,N_2816);
nor U3083 (N_3083,N_2523,N_2764);
nand U3084 (N_3084,N_2684,N_2965);
xnor U3085 (N_3085,N_2608,N_2552);
and U3086 (N_3086,N_2531,N_2945);
and U3087 (N_3087,N_2629,N_2716);
or U3088 (N_3088,N_2937,N_2793);
nor U3089 (N_3089,N_2765,N_2651);
xnor U3090 (N_3090,N_2561,N_2573);
or U3091 (N_3091,N_2766,N_2872);
nor U3092 (N_3092,N_2723,N_2703);
or U3093 (N_3093,N_2712,N_2806);
or U3094 (N_3094,N_2655,N_2640);
nor U3095 (N_3095,N_2756,N_2839);
or U3096 (N_3096,N_2695,N_2884);
nor U3097 (N_3097,N_2734,N_2912);
nand U3098 (N_3098,N_2551,N_2850);
nor U3099 (N_3099,N_2657,N_2610);
xor U3100 (N_3100,N_2960,N_2582);
nor U3101 (N_3101,N_2578,N_2516);
and U3102 (N_3102,N_2676,N_2781);
nand U3103 (N_3103,N_2899,N_2754);
or U3104 (N_3104,N_2870,N_2587);
and U3105 (N_3105,N_2834,N_2904);
xor U3106 (N_3106,N_2730,N_2977);
nor U3107 (N_3107,N_2709,N_2874);
nor U3108 (N_3108,N_2931,N_2867);
and U3109 (N_3109,N_2967,N_2841);
xnor U3110 (N_3110,N_2627,N_2599);
and U3111 (N_3111,N_2885,N_2948);
nand U3112 (N_3112,N_2762,N_2568);
or U3113 (N_3113,N_2519,N_2797);
nor U3114 (N_3114,N_2612,N_2634);
nor U3115 (N_3115,N_2901,N_2586);
nand U3116 (N_3116,N_2836,N_2815);
nand U3117 (N_3117,N_2748,N_2788);
and U3118 (N_3118,N_2803,N_2838);
or U3119 (N_3119,N_2936,N_2539);
and U3120 (N_3120,N_2628,N_2584);
or U3121 (N_3121,N_2542,N_2935);
and U3122 (N_3122,N_2530,N_2509);
xnor U3123 (N_3123,N_2665,N_2891);
or U3124 (N_3124,N_2564,N_2774);
nand U3125 (N_3125,N_2767,N_2524);
or U3126 (N_3126,N_2557,N_2760);
xor U3127 (N_3127,N_2544,N_2959);
or U3128 (N_3128,N_2593,N_2833);
or U3129 (N_3129,N_2970,N_2777);
nand U3130 (N_3130,N_2894,N_2859);
or U3131 (N_3131,N_2569,N_2546);
and U3132 (N_3132,N_2768,N_2642);
nor U3133 (N_3133,N_2840,N_2917);
xor U3134 (N_3134,N_2698,N_2824);
nor U3135 (N_3135,N_2920,N_2852);
or U3136 (N_3136,N_2890,N_2830);
nand U3137 (N_3137,N_2554,N_2636);
nand U3138 (N_3138,N_2871,N_2813);
and U3139 (N_3139,N_2933,N_2783);
or U3140 (N_3140,N_2606,N_2980);
and U3141 (N_3141,N_2866,N_2624);
or U3142 (N_3142,N_2855,N_2515);
or U3143 (N_3143,N_2773,N_2921);
xnor U3144 (N_3144,N_2650,N_2719);
nor U3145 (N_3145,N_2671,N_2927);
nor U3146 (N_3146,N_2538,N_2938);
xnor U3147 (N_3147,N_2751,N_2535);
and U3148 (N_3148,N_2579,N_2696);
xor U3149 (N_3149,N_2576,N_2680);
or U3150 (N_3150,N_2758,N_2805);
and U3151 (N_3151,N_2843,N_2570);
or U3152 (N_3152,N_2812,N_2752);
and U3153 (N_3153,N_2883,N_2915);
or U3154 (N_3154,N_2600,N_2998);
nor U3155 (N_3155,N_2739,N_2949);
nand U3156 (N_3156,N_2673,N_2807);
and U3157 (N_3157,N_2633,N_2656);
and U3158 (N_3158,N_2727,N_2721);
nand U3159 (N_3159,N_2691,N_2814);
nor U3160 (N_3160,N_2926,N_2895);
nand U3161 (N_3161,N_2672,N_2750);
nand U3162 (N_3162,N_2646,N_2532);
nor U3163 (N_3163,N_2818,N_2733);
or U3164 (N_3164,N_2641,N_2786);
nand U3165 (N_3165,N_2746,N_2802);
or U3166 (N_3166,N_2763,N_2731);
and U3167 (N_3167,N_2553,N_2548);
xnor U3168 (N_3168,N_2888,N_2858);
xor U3169 (N_3169,N_2694,N_2574);
or U3170 (N_3170,N_2795,N_2993);
and U3171 (N_3171,N_2971,N_2559);
xnor U3172 (N_3172,N_2631,N_2681);
and U3173 (N_3173,N_2529,N_2944);
nand U3174 (N_3174,N_2617,N_2592);
or U3175 (N_3175,N_2603,N_2682);
or U3176 (N_3176,N_2953,N_2794);
nor U3177 (N_3177,N_2686,N_2969);
or U3178 (N_3178,N_2903,N_2809);
nand U3179 (N_3179,N_2711,N_2875);
nor U3180 (N_3180,N_2823,N_2626);
nand U3181 (N_3181,N_2835,N_2796);
and U3182 (N_3182,N_2683,N_2512);
xnor U3183 (N_3183,N_2963,N_2979);
nor U3184 (N_3184,N_2644,N_2956);
xnor U3185 (N_3185,N_2753,N_2913);
nor U3186 (N_3186,N_2705,N_2880);
nor U3187 (N_3187,N_2660,N_2741);
nand U3188 (N_3188,N_2678,N_2846);
xnor U3189 (N_3189,N_2911,N_2598);
and U3190 (N_3190,N_2591,N_2565);
and U3191 (N_3191,N_2602,N_2654);
xor U3192 (N_3192,N_2987,N_2659);
nand U3193 (N_3193,N_2618,N_2974);
and U3194 (N_3194,N_2670,N_2580);
and U3195 (N_3195,N_2779,N_2929);
xnor U3196 (N_3196,N_2865,N_2708);
nor U3197 (N_3197,N_2853,N_2632);
xor U3198 (N_3198,N_2958,N_2991);
nor U3199 (N_3199,N_2811,N_2521);
xnor U3200 (N_3200,N_2907,N_2635);
and U3201 (N_3201,N_2502,N_2737);
xor U3202 (N_3202,N_2567,N_2861);
nand U3203 (N_3203,N_2932,N_2663);
nor U3204 (N_3204,N_2668,N_2687);
nor U3205 (N_3205,N_2928,N_2661);
or U3206 (N_3206,N_2854,N_2982);
or U3207 (N_3207,N_2992,N_2924);
nor U3208 (N_3208,N_2990,N_2702);
or U3209 (N_3209,N_2714,N_2674);
xnor U3210 (N_3210,N_2851,N_2887);
or U3211 (N_3211,N_2946,N_2537);
and U3212 (N_3212,N_2722,N_2827);
and U3213 (N_3213,N_2518,N_2563);
or U3214 (N_3214,N_2555,N_2925);
xor U3215 (N_3215,N_2692,N_2615);
or U3216 (N_3216,N_2975,N_2755);
or U3217 (N_3217,N_2930,N_2863);
xnor U3218 (N_3218,N_2984,N_2526);
nand U3219 (N_3219,N_2864,N_2909);
xnor U3220 (N_3220,N_2868,N_2605);
nor U3221 (N_3221,N_2621,N_2877);
and U3222 (N_3222,N_2520,N_2715);
xnor U3223 (N_3223,N_2507,N_2738);
nor U3224 (N_3224,N_2996,N_2819);
nand U3225 (N_3225,N_2973,N_2589);
xnor U3226 (N_3226,N_2837,N_2614);
nor U3227 (N_3227,N_2957,N_2947);
and U3228 (N_3228,N_2869,N_2697);
nor U3229 (N_3229,N_2685,N_2571);
nor U3230 (N_3230,N_2943,N_2572);
nor U3231 (N_3231,N_2983,N_2514);
xnor U3232 (N_3232,N_2898,N_2649);
or U3233 (N_3233,N_2594,N_2675);
xor U3234 (N_3234,N_2848,N_2505);
or U3235 (N_3235,N_2597,N_2747);
nor U3236 (N_3236,N_2560,N_2847);
or U3237 (N_3237,N_2604,N_2583);
xnor U3238 (N_3238,N_2790,N_2981);
or U3239 (N_3239,N_2940,N_2581);
or U3240 (N_3240,N_2999,N_2782);
and U3241 (N_3241,N_2914,N_2900);
or U3242 (N_3242,N_2744,N_2522);
xor U3243 (N_3243,N_2625,N_2638);
nand U3244 (N_3244,N_2652,N_2517);
or U3245 (N_3245,N_2585,N_2724);
nand U3246 (N_3246,N_2906,N_2728);
xor U3247 (N_3247,N_2897,N_2985);
nand U3248 (N_3248,N_2902,N_2653);
xnor U3249 (N_3249,N_2916,N_2961);
or U3250 (N_3250,N_2929,N_2791);
nand U3251 (N_3251,N_2984,N_2997);
and U3252 (N_3252,N_2859,N_2574);
nor U3253 (N_3253,N_2747,N_2951);
xnor U3254 (N_3254,N_2553,N_2891);
nand U3255 (N_3255,N_2531,N_2585);
and U3256 (N_3256,N_2685,N_2752);
xor U3257 (N_3257,N_2790,N_2641);
nand U3258 (N_3258,N_2818,N_2654);
and U3259 (N_3259,N_2658,N_2914);
xor U3260 (N_3260,N_2969,N_2616);
or U3261 (N_3261,N_2565,N_2616);
or U3262 (N_3262,N_2931,N_2962);
or U3263 (N_3263,N_2627,N_2885);
xor U3264 (N_3264,N_2504,N_2525);
and U3265 (N_3265,N_2646,N_2934);
nor U3266 (N_3266,N_2568,N_2640);
and U3267 (N_3267,N_2891,N_2901);
xor U3268 (N_3268,N_2833,N_2676);
nand U3269 (N_3269,N_2993,N_2743);
nand U3270 (N_3270,N_2555,N_2657);
nand U3271 (N_3271,N_2887,N_2663);
nand U3272 (N_3272,N_2710,N_2743);
nand U3273 (N_3273,N_2520,N_2536);
and U3274 (N_3274,N_2951,N_2776);
nand U3275 (N_3275,N_2683,N_2945);
nor U3276 (N_3276,N_2905,N_2898);
and U3277 (N_3277,N_2759,N_2802);
or U3278 (N_3278,N_2512,N_2841);
xor U3279 (N_3279,N_2873,N_2978);
nor U3280 (N_3280,N_2935,N_2751);
or U3281 (N_3281,N_2615,N_2706);
and U3282 (N_3282,N_2722,N_2540);
or U3283 (N_3283,N_2635,N_2904);
and U3284 (N_3284,N_2763,N_2756);
nor U3285 (N_3285,N_2931,N_2988);
nor U3286 (N_3286,N_2792,N_2893);
xnor U3287 (N_3287,N_2514,N_2507);
nand U3288 (N_3288,N_2873,N_2912);
nor U3289 (N_3289,N_2719,N_2987);
or U3290 (N_3290,N_2617,N_2861);
nor U3291 (N_3291,N_2998,N_2871);
nor U3292 (N_3292,N_2671,N_2703);
and U3293 (N_3293,N_2859,N_2769);
xnor U3294 (N_3294,N_2864,N_2606);
xnor U3295 (N_3295,N_2842,N_2754);
and U3296 (N_3296,N_2613,N_2748);
xor U3297 (N_3297,N_2565,N_2747);
nand U3298 (N_3298,N_2726,N_2827);
xor U3299 (N_3299,N_2941,N_2507);
xnor U3300 (N_3300,N_2902,N_2854);
nand U3301 (N_3301,N_2533,N_2594);
nor U3302 (N_3302,N_2680,N_2720);
nand U3303 (N_3303,N_2910,N_2953);
or U3304 (N_3304,N_2719,N_2992);
xnor U3305 (N_3305,N_2777,N_2959);
nor U3306 (N_3306,N_2650,N_2596);
nand U3307 (N_3307,N_2978,N_2906);
or U3308 (N_3308,N_2708,N_2561);
nand U3309 (N_3309,N_2896,N_2542);
nand U3310 (N_3310,N_2658,N_2951);
nor U3311 (N_3311,N_2995,N_2632);
nand U3312 (N_3312,N_2788,N_2967);
or U3313 (N_3313,N_2767,N_2565);
and U3314 (N_3314,N_2579,N_2801);
and U3315 (N_3315,N_2672,N_2778);
xor U3316 (N_3316,N_2744,N_2933);
xor U3317 (N_3317,N_2938,N_2936);
nor U3318 (N_3318,N_2918,N_2639);
and U3319 (N_3319,N_2803,N_2596);
or U3320 (N_3320,N_2855,N_2942);
xnor U3321 (N_3321,N_2717,N_2743);
nor U3322 (N_3322,N_2984,N_2582);
xnor U3323 (N_3323,N_2823,N_2660);
and U3324 (N_3324,N_2732,N_2622);
or U3325 (N_3325,N_2645,N_2952);
xor U3326 (N_3326,N_2699,N_2522);
nand U3327 (N_3327,N_2922,N_2908);
nor U3328 (N_3328,N_2623,N_2759);
nor U3329 (N_3329,N_2653,N_2714);
xor U3330 (N_3330,N_2910,N_2858);
nand U3331 (N_3331,N_2771,N_2858);
nor U3332 (N_3332,N_2727,N_2670);
nand U3333 (N_3333,N_2536,N_2718);
or U3334 (N_3334,N_2874,N_2929);
nand U3335 (N_3335,N_2736,N_2661);
xor U3336 (N_3336,N_2986,N_2825);
xnor U3337 (N_3337,N_2954,N_2880);
xor U3338 (N_3338,N_2876,N_2854);
and U3339 (N_3339,N_2821,N_2856);
or U3340 (N_3340,N_2905,N_2931);
and U3341 (N_3341,N_2798,N_2670);
or U3342 (N_3342,N_2962,N_2771);
nand U3343 (N_3343,N_2595,N_2630);
nand U3344 (N_3344,N_2716,N_2778);
or U3345 (N_3345,N_2842,N_2543);
nor U3346 (N_3346,N_2994,N_2540);
nand U3347 (N_3347,N_2548,N_2937);
nor U3348 (N_3348,N_2866,N_2629);
or U3349 (N_3349,N_2791,N_2742);
nand U3350 (N_3350,N_2799,N_2974);
nand U3351 (N_3351,N_2737,N_2625);
nor U3352 (N_3352,N_2963,N_2780);
xor U3353 (N_3353,N_2522,N_2842);
or U3354 (N_3354,N_2990,N_2577);
xnor U3355 (N_3355,N_2551,N_2921);
and U3356 (N_3356,N_2631,N_2535);
and U3357 (N_3357,N_2957,N_2751);
nor U3358 (N_3358,N_2914,N_2609);
nand U3359 (N_3359,N_2748,N_2936);
nor U3360 (N_3360,N_2910,N_2619);
or U3361 (N_3361,N_2508,N_2734);
xor U3362 (N_3362,N_2916,N_2664);
xor U3363 (N_3363,N_2567,N_2868);
nor U3364 (N_3364,N_2673,N_2859);
xor U3365 (N_3365,N_2943,N_2573);
xnor U3366 (N_3366,N_2572,N_2965);
xor U3367 (N_3367,N_2935,N_2623);
and U3368 (N_3368,N_2814,N_2854);
and U3369 (N_3369,N_2717,N_2667);
xor U3370 (N_3370,N_2938,N_2821);
or U3371 (N_3371,N_2520,N_2845);
xnor U3372 (N_3372,N_2904,N_2806);
nand U3373 (N_3373,N_2913,N_2703);
and U3374 (N_3374,N_2749,N_2864);
and U3375 (N_3375,N_2598,N_2729);
nand U3376 (N_3376,N_2791,N_2900);
nor U3377 (N_3377,N_2884,N_2997);
or U3378 (N_3378,N_2760,N_2584);
or U3379 (N_3379,N_2579,N_2703);
xnor U3380 (N_3380,N_2663,N_2783);
nand U3381 (N_3381,N_2783,N_2606);
nand U3382 (N_3382,N_2779,N_2770);
xnor U3383 (N_3383,N_2683,N_2949);
nor U3384 (N_3384,N_2894,N_2542);
and U3385 (N_3385,N_2646,N_2533);
xor U3386 (N_3386,N_2565,N_2772);
nand U3387 (N_3387,N_2784,N_2647);
or U3388 (N_3388,N_2555,N_2777);
and U3389 (N_3389,N_2747,N_2815);
and U3390 (N_3390,N_2642,N_2675);
xor U3391 (N_3391,N_2597,N_2674);
xor U3392 (N_3392,N_2602,N_2938);
nor U3393 (N_3393,N_2732,N_2907);
or U3394 (N_3394,N_2627,N_2788);
xor U3395 (N_3395,N_2932,N_2624);
or U3396 (N_3396,N_2542,N_2798);
nand U3397 (N_3397,N_2724,N_2647);
and U3398 (N_3398,N_2979,N_2671);
and U3399 (N_3399,N_2617,N_2793);
or U3400 (N_3400,N_2940,N_2925);
nor U3401 (N_3401,N_2653,N_2655);
and U3402 (N_3402,N_2990,N_2505);
nor U3403 (N_3403,N_2597,N_2844);
or U3404 (N_3404,N_2500,N_2736);
xor U3405 (N_3405,N_2677,N_2964);
or U3406 (N_3406,N_2641,N_2603);
xor U3407 (N_3407,N_2702,N_2897);
nor U3408 (N_3408,N_2693,N_2664);
nand U3409 (N_3409,N_2818,N_2861);
and U3410 (N_3410,N_2931,N_2733);
xnor U3411 (N_3411,N_2663,N_2936);
or U3412 (N_3412,N_2741,N_2568);
nor U3413 (N_3413,N_2897,N_2714);
nor U3414 (N_3414,N_2641,N_2813);
nor U3415 (N_3415,N_2790,N_2685);
xnor U3416 (N_3416,N_2908,N_2872);
and U3417 (N_3417,N_2879,N_2799);
xor U3418 (N_3418,N_2629,N_2517);
or U3419 (N_3419,N_2608,N_2556);
xnor U3420 (N_3420,N_2646,N_2775);
and U3421 (N_3421,N_2931,N_2525);
or U3422 (N_3422,N_2524,N_2693);
or U3423 (N_3423,N_2523,N_2826);
and U3424 (N_3424,N_2780,N_2971);
and U3425 (N_3425,N_2642,N_2543);
nand U3426 (N_3426,N_2924,N_2701);
nand U3427 (N_3427,N_2559,N_2529);
and U3428 (N_3428,N_2987,N_2684);
nor U3429 (N_3429,N_2772,N_2841);
and U3430 (N_3430,N_2893,N_2729);
or U3431 (N_3431,N_2616,N_2815);
xnor U3432 (N_3432,N_2676,N_2621);
xnor U3433 (N_3433,N_2871,N_2500);
xor U3434 (N_3434,N_2786,N_2813);
nor U3435 (N_3435,N_2552,N_2940);
nand U3436 (N_3436,N_2946,N_2726);
xnor U3437 (N_3437,N_2570,N_2782);
nand U3438 (N_3438,N_2797,N_2904);
nor U3439 (N_3439,N_2612,N_2763);
or U3440 (N_3440,N_2664,N_2731);
or U3441 (N_3441,N_2925,N_2754);
or U3442 (N_3442,N_2894,N_2590);
nor U3443 (N_3443,N_2844,N_2858);
or U3444 (N_3444,N_2885,N_2777);
or U3445 (N_3445,N_2681,N_2748);
xnor U3446 (N_3446,N_2844,N_2988);
nor U3447 (N_3447,N_2790,N_2551);
nand U3448 (N_3448,N_2747,N_2717);
xor U3449 (N_3449,N_2998,N_2639);
nor U3450 (N_3450,N_2638,N_2933);
xnor U3451 (N_3451,N_2617,N_2764);
nand U3452 (N_3452,N_2858,N_2624);
nand U3453 (N_3453,N_2825,N_2614);
xor U3454 (N_3454,N_2913,N_2902);
nor U3455 (N_3455,N_2824,N_2670);
or U3456 (N_3456,N_2819,N_2920);
nand U3457 (N_3457,N_2875,N_2503);
nand U3458 (N_3458,N_2573,N_2511);
and U3459 (N_3459,N_2904,N_2543);
xor U3460 (N_3460,N_2712,N_2563);
and U3461 (N_3461,N_2955,N_2801);
and U3462 (N_3462,N_2598,N_2800);
nand U3463 (N_3463,N_2683,N_2970);
xnor U3464 (N_3464,N_2605,N_2987);
nor U3465 (N_3465,N_2503,N_2954);
and U3466 (N_3466,N_2766,N_2817);
xor U3467 (N_3467,N_2832,N_2707);
nor U3468 (N_3468,N_2617,N_2932);
xor U3469 (N_3469,N_2525,N_2694);
xor U3470 (N_3470,N_2661,N_2625);
and U3471 (N_3471,N_2897,N_2973);
or U3472 (N_3472,N_2525,N_2619);
xor U3473 (N_3473,N_2660,N_2503);
xnor U3474 (N_3474,N_2663,N_2503);
or U3475 (N_3475,N_2514,N_2656);
or U3476 (N_3476,N_2583,N_2887);
xor U3477 (N_3477,N_2726,N_2758);
nand U3478 (N_3478,N_2945,N_2624);
or U3479 (N_3479,N_2654,N_2658);
nor U3480 (N_3480,N_2779,N_2549);
or U3481 (N_3481,N_2977,N_2822);
nand U3482 (N_3482,N_2799,N_2560);
or U3483 (N_3483,N_2802,N_2841);
xor U3484 (N_3484,N_2989,N_2732);
and U3485 (N_3485,N_2882,N_2891);
xnor U3486 (N_3486,N_2884,N_2908);
xnor U3487 (N_3487,N_2951,N_2913);
xor U3488 (N_3488,N_2518,N_2507);
nand U3489 (N_3489,N_2996,N_2541);
and U3490 (N_3490,N_2760,N_2547);
xor U3491 (N_3491,N_2802,N_2790);
and U3492 (N_3492,N_2831,N_2960);
nor U3493 (N_3493,N_2528,N_2988);
and U3494 (N_3494,N_2869,N_2725);
or U3495 (N_3495,N_2652,N_2692);
nor U3496 (N_3496,N_2948,N_2631);
xnor U3497 (N_3497,N_2756,N_2771);
nand U3498 (N_3498,N_2990,N_2996);
nand U3499 (N_3499,N_2954,N_2864);
and U3500 (N_3500,N_3046,N_3067);
xor U3501 (N_3501,N_3160,N_3448);
xnor U3502 (N_3502,N_3224,N_3281);
nand U3503 (N_3503,N_3494,N_3049);
xor U3504 (N_3504,N_3241,N_3014);
and U3505 (N_3505,N_3223,N_3198);
or U3506 (N_3506,N_3444,N_3272);
nand U3507 (N_3507,N_3047,N_3188);
nand U3508 (N_3508,N_3112,N_3481);
and U3509 (N_3509,N_3383,N_3086);
nand U3510 (N_3510,N_3017,N_3107);
or U3511 (N_3511,N_3460,N_3474);
or U3512 (N_3512,N_3393,N_3249);
nand U3513 (N_3513,N_3080,N_3176);
nand U3514 (N_3514,N_3171,N_3173);
xnor U3515 (N_3515,N_3259,N_3394);
and U3516 (N_3516,N_3002,N_3335);
or U3517 (N_3517,N_3234,N_3099);
nor U3518 (N_3518,N_3385,N_3058);
nand U3519 (N_3519,N_3120,N_3125);
or U3520 (N_3520,N_3206,N_3359);
xnor U3521 (N_3521,N_3384,N_3435);
or U3522 (N_3522,N_3380,N_3311);
or U3523 (N_3523,N_3273,N_3271);
xnor U3524 (N_3524,N_3289,N_3456);
and U3525 (N_3525,N_3468,N_3091);
nor U3526 (N_3526,N_3346,N_3033);
or U3527 (N_3527,N_3462,N_3278);
or U3528 (N_3528,N_3236,N_3454);
and U3529 (N_3529,N_3111,N_3436);
nor U3530 (N_3530,N_3313,N_3212);
xor U3531 (N_3531,N_3180,N_3239);
and U3532 (N_3532,N_3297,N_3088);
or U3533 (N_3533,N_3178,N_3485);
nor U3534 (N_3534,N_3416,N_3177);
or U3535 (N_3535,N_3317,N_3333);
or U3536 (N_3536,N_3170,N_3071);
and U3537 (N_3537,N_3194,N_3202);
nand U3538 (N_3538,N_3362,N_3439);
or U3539 (N_3539,N_3341,N_3077);
nand U3540 (N_3540,N_3122,N_3219);
and U3541 (N_3541,N_3034,N_3050);
or U3542 (N_3542,N_3225,N_3497);
xnor U3543 (N_3543,N_3179,N_3300);
or U3544 (N_3544,N_3447,N_3493);
xnor U3545 (N_3545,N_3193,N_3132);
or U3546 (N_3546,N_3325,N_3477);
or U3547 (N_3547,N_3004,N_3262);
nor U3548 (N_3548,N_3440,N_3312);
nor U3549 (N_3549,N_3103,N_3204);
nor U3550 (N_3550,N_3075,N_3213);
nor U3551 (N_3551,N_3216,N_3282);
or U3552 (N_3552,N_3141,N_3404);
nand U3553 (N_3553,N_3438,N_3410);
xnor U3554 (N_3554,N_3471,N_3061);
and U3555 (N_3555,N_3016,N_3274);
or U3556 (N_3556,N_3126,N_3302);
and U3557 (N_3557,N_3339,N_3064);
and U3558 (N_3558,N_3015,N_3108);
or U3559 (N_3559,N_3328,N_3028);
or U3560 (N_3560,N_3123,N_3130);
nand U3561 (N_3561,N_3473,N_3310);
and U3562 (N_3562,N_3109,N_3463);
or U3563 (N_3563,N_3348,N_3402);
nand U3564 (N_3564,N_3025,N_3000);
xor U3565 (N_3565,N_3467,N_3442);
nor U3566 (N_3566,N_3258,N_3137);
xnor U3567 (N_3567,N_3165,N_3490);
or U3568 (N_3568,N_3452,N_3391);
or U3569 (N_3569,N_3327,N_3048);
or U3570 (N_3570,N_3323,N_3063);
nand U3571 (N_3571,N_3221,N_3181);
or U3572 (N_3572,N_3389,N_3106);
nor U3573 (N_3573,N_3466,N_3405);
and U3574 (N_3574,N_3338,N_3066);
nor U3575 (N_3575,N_3035,N_3269);
or U3576 (N_3576,N_3461,N_3101);
or U3577 (N_3577,N_3255,N_3018);
nand U3578 (N_3578,N_3465,N_3403);
and U3579 (N_3579,N_3052,N_3070);
nand U3580 (N_3580,N_3128,N_3147);
xor U3581 (N_3581,N_3256,N_3475);
or U3582 (N_3582,N_3043,N_3265);
nand U3583 (N_3583,N_3295,N_3069);
or U3584 (N_3584,N_3051,N_3476);
nand U3585 (N_3585,N_3196,N_3482);
nand U3586 (N_3586,N_3175,N_3149);
and U3587 (N_3587,N_3232,N_3378);
and U3588 (N_3588,N_3270,N_3499);
nand U3589 (N_3589,N_3084,N_3250);
nand U3590 (N_3590,N_3329,N_3153);
nand U3591 (N_3591,N_3395,N_3315);
nand U3592 (N_3592,N_3230,N_3089);
or U3593 (N_3593,N_3087,N_3429);
nor U3594 (N_3594,N_3209,N_3027);
nor U3595 (N_3595,N_3427,N_3010);
nand U3596 (N_3596,N_3409,N_3116);
and U3597 (N_3597,N_3286,N_3261);
and U3598 (N_3598,N_3100,N_3082);
nor U3599 (N_3599,N_3483,N_3486);
xor U3600 (N_3600,N_3334,N_3370);
nand U3601 (N_3601,N_3218,N_3055);
nor U3602 (N_3602,N_3365,N_3222);
or U3603 (N_3603,N_3372,N_3161);
xnor U3604 (N_3604,N_3131,N_3321);
nor U3605 (N_3605,N_3013,N_3214);
or U3606 (N_3606,N_3062,N_3023);
nor U3607 (N_3607,N_3157,N_3280);
xor U3608 (N_3608,N_3158,N_3314);
nor U3609 (N_3609,N_3022,N_3294);
nor U3610 (N_3610,N_3428,N_3257);
nor U3611 (N_3611,N_3470,N_3492);
or U3612 (N_3612,N_3182,N_3146);
nor U3613 (N_3613,N_3226,N_3277);
or U3614 (N_3614,N_3453,N_3105);
xor U3615 (N_3615,N_3041,N_3469);
nor U3616 (N_3616,N_3373,N_3331);
nor U3617 (N_3617,N_3162,N_3386);
xor U3618 (N_3618,N_3129,N_3392);
xnor U3619 (N_3619,N_3491,N_3079);
xnor U3620 (N_3620,N_3039,N_3056);
nand U3621 (N_3621,N_3285,N_3478);
or U3622 (N_3622,N_3387,N_3356);
or U3623 (N_3623,N_3431,N_3361);
nor U3624 (N_3624,N_3007,N_3498);
and U3625 (N_3625,N_3237,N_3235);
and U3626 (N_3626,N_3065,N_3008);
nand U3627 (N_3627,N_3211,N_3276);
and U3628 (N_3628,N_3368,N_3375);
or U3629 (N_3629,N_3284,N_3293);
nor U3630 (N_3630,N_3441,N_3119);
nor U3631 (N_3631,N_3135,N_3296);
xnor U3632 (N_3632,N_3220,N_3417);
and U3633 (N_3633,N_3369,N_3190);
xnor U3634 (N_3634,N_3053,N_3267);
and U3635 (N_3635,N_3248,N_3037);
or U3636 (N_3636,N_3426,N_3005);
xor U3637 (N_3637,N_3060,N_3117);
and U3638 (N_3638,N_3420,N_3174);
or U3639 (N_3639,N_3200,N_3412);
nand U3640 (N_3640,N_3422,N_3085);
and U3641 (N_3641,N_3287,N_3186);
nand U3642 (N_3642,N_3183,N_3118);
or U3643 (N_3643,N_3152,N_3090);
and U3644 (N_3644,N_3093,N_3367);
or U3645 (N_3645,N_3187,N_3144);
nand U3646 (N_3646,N_3078,N_3419);
and U3647 (N_3647,N_3390,N_3299);
nor U3648 (N_3648,N_3363,N_3487);
or U3649 (N_3649,N_3399,N_3217);
or U3650 (N_3650,N_3038,N_3414);
and U3651 (N_3651,N_3283,N_3247);
xnor U3652 (N_3652,N_3164,N_3104);
or U3653 (N_3653,N_3057,N_3244);
nor U3654 (N_3654,N_3203,N_3102);
or U3655 (N_3655,N_3288,N_3360);
xor U3656 (N_3656,N_3148,N_3446);
nand U3657 (N_3657,N_3115,N_3199);
xnor U3658 (N_3658,N_3326,N_3336);
nor U3659 (N_3659,N_3352,N_3423);
xor U3660 (N_3660,N_3024,N_3318);
or U3661 (N_3661,N_3309,N_3266);
nand U3662 (N_3662,N_3430,N_3154);
and U3663 (N_3663,N_3113,N_3040);
or U3664 (N_3664,N_3425,N_3434);
and U3665 (N_3665,N_3401,N_3011);
xnor U3666 (N_3666,N_3340,N_3207);
nand U3667 (N_3667,N_3397,N_3030);
or U3668 (N_3668,N_3001,N_3324);
nand U3669 (N_3669,N_3254,N_3026);
xnor U3670 (N_3670,N_3081,N_3455);
or U3671 (N_3671,N_3459,N_3305);
and U3672 (N_3672,N_3201,N_3308);
and U3673 (N_3673,N_3012,N_3433);
nor U3674 (N_3674,N_3134,N_3437);
nand U3675 (N_3675,N_3243,N_3238);
or U3676 (N_3676,N_3095,N_3320);
nor U3677 (N_3677,N_3197,N_3036);
nor U3678 (N_3678,N_3054,N_3127);
xnor U3679 (N_3679,N_3142,N_3381);
or U3680 (N_3680,N_3354,N_3306);
or U3681 (N_3681,N_3139,N_3457);
xor U3682 (N_3682,N_3076,N_3143);
nor U3683 (N_3683,N_3421,N_3019);
or U3684 (N_3684,N_3489,N_3145);
nand U3685 (N_3685,N_3020,N_3364);
and U3686 (N_3686,N_3316,N_3353);
xnor U3687 (N_3687,N_3445,N_3045);
nor U3688 (N_3688,N_3229,N_3150);
and U3689 (N_3689,N_3322,N_3344);
xnor U3690 (N_3690,N_3097,N_3059);
xor U3691 (N_3691,N_3379,N_3227);
and U3692 (N_3692,N_3319,N_3138);
and U3693 (N_3693,N_3291,N_3396);
xnor U3694 (N_3694,N_3382,N_3228);
xor U3695 (N_3695,N_3342,N_3156);
or U3696 (N_3696,N_3124,N_3031);
xor U3697 (N_3697,N_3407,N_3068);
nand U3698 (N_3698,N_3184,N_3350);
and U3699 (N_3699,N_3275,N_3424);
nor U3700 (N_3700,N_3133,N_3358);
and U3701 (N_3701,N_3376,N_3083);
nand U3702 (N_3702,N_3121,N_3406);
nand U3703 (N_3703,N_3480,N_3377);
or U3704 (N_3704,N_3345,N_3073);
or U3705 (N_3705,N_3195,N_3307);
xnor U3706 (N_3706,N_3298,N_3208);
or U3707 (N_3707,N_3398,N_3233);
and U3708 (N_3708,N_3355,N_3450);
nor U3709 (N_3709,N_3029,N_3451);
xnor U3710 (N_3710,N_3003,N_3242);
xnor U3711 (N_3711,N_3264,N_3246);
xor U3712 (N_3712,N_3290,N_3151);
and U3713 (N_3713,N_3432,N_3496);
nor U3714 (N_3714,N_3495,N_3303);
nor U3715 (N_3715,N_3166,N_3260);
nor U3716 (N_3716,N_3374,N_3279);
and U3717 (N_3717,N_3413,N_3400);
and U3718 (N_3718,N_3245,N_3332);
or U3719 (N_3719,N_3009,N_3163);
nor U3720 (N_3720,N_3098,N_3159);
xor U3721 (N_3721,N_3240,N_3172);
nor U3722 (N_3722,N_3268,N_3330);
xor U3723 (N_3723,N_3415,N_3168);
xnor U3724 (N_3724,N_3251,N_3167);
and U3725 (N_3725,N_3304,N_3337);
nor U3726 (N_3726,N_3351,N_3458);
nor U3727 (N_3727,N_3408,N_3140);
or U3728 (N_3728,N_3231,N_3044);
and U3729 (N_3729,N_3371,N_3136);
nor U3730 (N_3730,N_3347,N_3210);
xnor U3731 (N_3731,N_3411,N_3094);
and U3732 (N_3732,N_3114,N_3449);
or U3733 (N_3733,N_3074,N_3484);
and U3734 (N_3734,N_3189,N_3418);
nor U3735 (N_3735,N_3472,N_3192);
nand U3736 (N_3736,N_3349,N_3191);
and U3737 (N_3737,N_3479,N_3253);
nand U3738 (N_3738,N_3072,N_3464);
nor U3739 (N_3739,N_3292,N_3042);
xnor U3740 (N_3740,N_3092,N_3215);
nand U3741 (N_3741,N_3021,N_3006);
and U3742 (N_3742,N_3032,N_3096);
or U3743 (N_3743,N_3343,N_3357);
or U3744 (N_3744,N_3169,N_3205);
nand U3745 (N_3745,N_3488,N_3301);
xnor U3746 (N_3746,N_3263,N_3366);
xnor U3747 (N_3747,N_3388,N_3443);
nor U3748 (N_3748,N_3185,N_3155);
nand U3749 (N_3749,N_3110,N_3252);
nand U3750 (N_3750,N_3026,N_3043);
nand U3751 (N_3751,N_3221,N_3469);
and U3752 (N_3752,N_3461,N_3287);
or U3753 (N_3753,N_3163,N_3154);
or U3754 (N_3754,N_3386,N_3063);
or U3755 (N_3755,N_3062,N_3426);
xnor U3756 (N_3756,N_3004,N_3190);
nor U3757 (N_3757,N_3211,N_3444);
nor U3758 (N_3758,N_3215,N_3111);
nand U3759 (N_3759,N_3264,N_3427);
or U3760 (N_3760,N_3354,N_3400);
nand U3761 (N_3761,N_3075,N_3207);
nand U3762 (N_3762,N_3383,N_3234);
and U3763 (N_3763,N_3157,N_3253);
or U3764 (N_3764,N_3024,N_3166);
or U3765 (N_3765,N_3377,N_3421);
nand U3766 (N_3766,N_3481,N_3211);
nor U3767 (N_3767,N_3249,N_3151);
nor U3768 (N_3768,N_3427,N_3316);
xnor U3769 (N_3769,N_3161,N_3371);
nor U3770 (N_3770,N_3109,N_3406);
or U3771 (N_3771,N_3208,N_3318);
nor U3772 (N_3772,N_3282,N_3371);
xnor U3773 (N_3773,N_3225,N_3170);
and U3774 (N_3774,N_3415,N_3170);
nor U3775 (N_3775,N_3349,N_3359);
nor U3776 (N_3776,N_3308,N_3456);
or U3777 (N_3777,N_3121,N_3060);
xnor U3778 (N_3778,N_3301,N_3080);
nand U3779 (N_3779,N_3080,N_3407);
nor U3780 (N_3780,N_3370,N_3078);
nand U3781 (N_3781,N_3001,N_3493);
xnor U3782 (N_3782,N_3416,N_3038);
and U3783 (N_3783,N_3473,N_3416);
nand U3784 (N_3784,N_3195,N_3358);
and U3785 (N_3785,N_3260,N_3170);
or U3786 (N_3786,N_3306,N_3303);
or U3787 (N_3787,N_3064,N_3300);
or U3788 (N_3788,N_3224,N_3023);
xnor U3789 (N_3789,N_3277,N_3047);
or U3790 (N_3790,N_3320,N_3377);
and U3791 (N_3791,N_3062,N_3494);
nor U3792 (N_3792,N_3396,N_3107);
nand U3793 (N_3793,N_3322,N_3302);
and U3794 (N_3794,N_3453,N_3011);
nand U3795 (N_3795,N_3373,N_3460);
and U3796 (N_3796,N_3054,N_3342);
xnor U3797 (N_3797,N_3271,N_3483);
and U3798 (N_3798,N_3419,N_3289);
xnor U3799 (N_3799,N_3115,N_3219);
and U3800 (N_3800,N_3479,N_3246);
or U3801 (N_3801,N_3345,N_3093);
nor U3802 (N_3802,N_3170,N_3424);
and U3803 (N_3803,N_3154,N_3499);
or U3804 (N_3804,N_3411,N_3141);
nand U3805 (N_3805,N_3450,N_3196);
and U3806 (N_3806,N_3381,N_3217);
nand U3807 (N_3807,N_3078,N_3099);
or U3808 (N_3808,N_3408,N_3122);
nand U3809 (N_3809,N_3207,N_3102);
xor U3810 (N_3810,N_3344,N_3404);
and U3811 (N_3811,N_3105,N_3097);
and U3812 (N_3812,N_3273,N_3481);
nor U3813 (N_3813,N_3118,N_3177);
nor U3814 (N_3814,N_3130,N_3083);
nor U3815 (N_3815,N_3280,N_3419);
xor U3816 (N_3816,N_3326,N_3296);
nor U3817 (N_3817,N_3055,N_3379);
or U3818 (N_3818,N_3265,N_3377);
or U3819 (N_3819,N_3077,N_3319);
or U3820 (N_3820,N_3306,N_3153);
nor U3821 (N_3821,N_3112,N_3400);
or U3822 (N_3822,N_3098,N_3131);
and U3823 (N_3823,N_3022,N_3290);
nand U3824 (N_3824,N_3143,N_3095);
xnor U3825 (N_3825,N_3351,N_3023);
nand U3826 (N_3826,N_3040,N_3268);
xnor U3827 (N_3827,N_3325,N_3429);
xor U3828 (N_3828,N_3238,N_3164);
or U3829 (N_3829,N_3287,N_3214);
nor U3830 (N_3830,N_3450,N_3147);
nor U3831 (N_3831,N_3381,N_3306);
nand U3832 (N_3832,N_3271,N_3042);
and U3833 (N_3833,N_3484,N_3199);
xnor U3834 (N_3834,N_3037,N_3253);
nor U3835 (N_3835,N_3298,N_3125);
xnor U3836 (N_3836,N_3473,N_3480);
or U3837 (N_3837,N_3097,N_3108);
or U3838 (N_3838,N_3087,N_3483);
nor U3839 (N_3839,N_3034,N_3306);
xnor U3840 (N_3840,N_3077,N_3278);
and U3841 (N_3841,N_3344,N_3372);
or U3842 (N_3842,N_3060,N_3003);
nand U3843 (N_3843,N_3199,N_3381);
xor U3844 (N_3844,N_3198,N_3287);
nor U3845 (N_3845,N_3085,N_3426);
nand U3846 (N_3846,N_3204,N_3342);
nand U3847 (N_3847,N_3317,N_3395);
nand U3848 (N_3848,N_3317,N_3352);
xor U3849 (N_3849,N_3170,N_3349);
xor U3850 (N_3850,N_3143,N_3080);
and U3851 (N_3851,N_3146,N_3195);
nand U3852 (N_3852,N_3204,N_3442);
or U3853 (N_3853,N_3434,N_3209);
nor U3854 (N_3854,N_3294,N_3130);
xnor U3855 (N_3855,N_3332,N_3178);
nor U3856 (N_3856,N_3314,N_3027);
or U3857 (N_3857,N_3218,N_3221);
xor U3858 (N_3858,N_3122,N_3180);
nand U3859 (N_3859,N_3020,N_3277);
nand U3860 (N_3860,N_3171,N_3055);
and U3861 (N_3861,N_3283,N_3147);
nor U3862 (N_3862,N_3127,N_3344);
xor U3863 (N_3863,N_3201,N_3377);
or U3864 (N_3864,N_3257,N_3497);
xor U3865 (N_3865,N_3463,N_3310);
and U3866 (N_3866,N_3392,N_3203);
and U3867 (N_3867,N_3140,N_3490);
or U3868 (N_3868,N_3180,N_3245);
xnor U3869 (N_3869,N_3430,N_3092);
or U3870 (N_3870,N_3300,N_3070);
or U3871 (N_3871,N_3321,N_3365);
or U3872 (N_3872,N_3192,N_3405);
nor U3873 (N_3873,N_3424,N_3354);
xor U3874 (N_3874,N_3134,N_3178);
and U3875 (N_3875,N_3268,N_3404);
or U3876 (N_3876,N_3444,N_3467);
nor U3877 (N_3877,N_3428,N_3415);
nand U3878 (N_3878,N_3398,N_3307);
or U3879 (N_3879,N_3005,N_3126);
nand U3880 (N_3880,N_3315,N_3097);
and U3881 (N_3881,N_3178,N_3192);
nand U3882 (N_3882,N_3407,N_3057);
nor U3883 (N_3883,N_3232,N_3497);
xnor U3884 (N_3884,N_3028,N_3082);
or U3885 (N_3885,N_3475,N_3127);
nand U3886 (N_3886,N_3023,N_3196);
and U3887 (N_3887,N_3352,N_3347);
or U3888 (N_3888,N_3228,N_3236);
or U3889 (N_3889,N_3415,N_3479);
xor U3890 (N_3890,N_3122,N_3290);
nor U3891 (N_3891,N_3145,N_3415);
and U3892 (N_3892,N_3188,N_3488);
nand U3893 (N_3893,N_3385,N_3325);
and U3894 (N_3894,N_3321,N_3259);
xnor U3895 (N_3895,N_3394,N_3320);
nor U3896 (N_3896,N_3030,N_3390);
and U3897 (N_3897,N_3321,N_3104);
nor U3898 (N_3898,N_3476,N_3463);
nor U3899 (N_3899,N_3104,N_3390);
nor U3900 (N_3900,N_3070,N_3013);
or U3901 (N_3901,N_3358,N_3013);
xnor U3902 (N_3902,N_3328,N_3436);
and U3903 (N_3903,N_3232,N_3127);
nand U3904 (N_3904,N_3469,N_3185);
nor U3905 (N_3905,N_3064,N_3370);
xnor U3906 (N_3906,N_3269,N_3226);
xnor U3907 (N_3907,N_3222,N_3346);
xor U3908 (N_3908,N_3341,N_3027);
nand U3909 (N_3909,N_3253,N_3012);
or U3910 (N_3910,N_3090,N_3070);
and U3911 (N_3911,N_3258,N_3322);
or U3912 (N_3912,N_3350,N_3118);
or U3913 (N_3913,N_3497,N_3410);
and U3914 (N_3914,N_3376,N_3369);
or U3915 (N_3915,N_3352,N_3222);
and U3916 (N_3916,N_3494,N_3375);
nand U3917 (N_3917,N_3118,N_3277);
or U3918 (N_3918,N_3065,N_3048);
or U3919 (N_3919,N_3114,N_3342);
or U3920 (N_3920,N_3355,N_3239);
nand U3921 (N_3921,N_3175,N_3257);
nor U3922 (N_3922,N_3332,N_3220);
xnor U3923 (N_3923,N_3230,N_3187);
nor U3924 (N_3924,N_3176,N_3200);
nor U3925 (N_3925,N_3365,N_3461);
xor U3926 (N_3926,N_3199,N_3278);
and U3927 (N_3927,N_3253,N_3318);
xor U3928 (N_3928,N_3006,N_3241);
nand U3929 (N_3929,N_3259,N_3101);
or U3930 (N_3930,N_3224,N_3456);
and U3931 (N_3931,N_3457,N_3173);
nor U3932 (N_3932,N_3453,N_3415);
nor U3933 (N_3933,N_3081,N_3039);
or U3934 (N_3934,N_3098,N_3158);
nor U3935 (N_3935,N_3350,N_3217);
and U3936 (N_3936,N_3054,N_3319);
or U3937 (N_3937,N_3007,N_3172);
nand U3938 (N_3938,N_3214,N_3452);
nor U3939 (N_3939,N_3046,N_3240);
xnor U3940 (N_3940,N_3101,N_3269);
nor U3941 (N_3941,N_3230,N_3062);
nor U3942 (N_3942,N_3317,N_3104);
nor U3943 (N_3943,N_3475,N_3012);
nor U3944 (N_3944,N_3349,N_3204);
and U3945 (N_3945,N_3470,N_3175);
nand U3946 (N_3946,N_3210,N_3460);
and U3947 (N_3947,N_3057,N_3155);
xnor U3948 (N_3948,N_3080,N_3345);
nand U3949 (N_3949,N_3235,N_3010);
nor U3950 (N_3950,N_3122,N_3205);
xnor U3951 (N_3951,N_3221,N_3345);
xnor U3952 (N_3952,N_3076,N_3405);
xor U3953 (N_3953,N_3263,N_3056);
nand U3954 (N_3954,N_3489,N_3247);
or U3955 (N_3955,N_3262,N_3381);
and U3956 (N_3956,N_3437,N_3385);
nor U3957 (N_3957,N_3383,N_3162);
nor U3958 (N_3958,N_3119,N_3313);
nor U3959 (N_3959,N_3361,N_3385);
nor U3960 (N_3960,N_3071,N_3436);
and U3961 (N_3961,N_3339,N_3190);
nor U3962 (N_3962,N_3489,N_3345);
nand U3963 (N_3963,N_3037,N_3207);
or U3964 (N_3964,N_3459,N_3162);
nand U3965 (N_3965,N_3148,N_3373);
xnor U3966 (N_3966,N_3461,N_3125);
nand U3967 (N_3967,N_3392,N_3052);
or U3968 (N_3968,N_3387,N_3003);
nor U3969 (N_3969,N_3486,N_3239);
xor U3970 (N_3970,N_3398,N_3434);
or U3971 (N_3971,N_3292,N_3366);
nand U3972 (N_3972,N_3147,N_3032);
nor U3973 (N_3973,N_3025,N_3260);
nor U3974 (N_3974,N_3190,N_3403);
or U3975 (N_3975,N_3380,N_3384);
xnor U3976 (N_3976,N_3361,N_3281);
nand U3977 (N_3977,N_3428,N_3125);
nor U3978 (N_3978,N_3315,N_3470);
xor U3979 (N_3979,N_3097,N_3167);
and U3980 (N_3980,N_3205,N_3440);
and U3981 (N_3981,N_3238,N_3372);
xor U3982 (N_3982,N_3029,N_3411);
xor U3983 (N_3983,N_3497,N_3020);
xnor U3984 (N_3984,N_3233,N_3165);
nor U3985 (N_3985,N_3445,N_3388);
or U3986 (N_3986,N_3464,N_3299);
and U3987 (N_3987,N_3210,N_3486);
nor U3988 (N_3988,N_3248,N_3266);
or U3989 (N_3989,N_3025,N_3209);
or U3990 (N_3990,N_3220,N_3222);
nand U3991 (N_3991,N_3347,N_3259);
xnor U3992 (N_3992,N_3308,N_3400);
nor U3993 (N_3993,N_3023,N_3445);
and U3994 (N_3994,N_3123,N_3038);
and U3995 (N_3995,N_3419,N_3196);
xnor U3996 (N_3996,N_3102,N_3116);
and U3997 (N_3997,N_3373,N_3431);
nand U3998 (N_3998,N_3344,N_3170);
and U3999 (N_3999,N_3024,N_3284);
nand U4000 (N_4000,N_3772,N_3950);
xnor U4001 (N_4001,N_3522,N_3862);
nand U4002 (N_4002,N_3547,N_3952);
xor U4003 (N_4003,N_3753,N_3821);
nor U4004 (N_4004,N_3894,N_3733);
nor U4005 (N_4005,N_3904,N_3725);
nor U4006 (N_4006,N_3805,N_3984);
and U4007 (N_4007,N_3909,N_3689);
and U4008 (N_4008,N_3568,N_3793);
nand U4009 (N_4009,N_3856,N_3743);
nand U4010 (N_4010,N_3691,N_3855);
nand U4011 (N_4011,N_3640,N_3515);
nor U4012 (N_4012,N_3641,N_3738);
and U4013 (N_4013,N_3523,N_3732);
nand U4014 (N_4014,N_3591,N_3869);
nand U4015 (N_4015,N_3915,N_3673);
nand U4016 (N_4016,N_3835,N_3863);
nand U4017 (N_4017,N_3584,N_3867);
nand U4018 (N_4018,N_3590,N_3596);
nor U4019 (N_4019,N_3723,N_3634);
nand U4020 (N_4020,N_3840,N_3620);
xor U4021 (N_4021,N_3581,N_3875);
and U4022 (N_4022,N_3938,N_3779);
or U4023 (N_4023,N_3657,N_3531);
xnor U4024 (N_4024,N_3714,N_3746);
nand U4025 (N_4025,N_3643,N_3841);
or U4026 (N_4026,N_3517,N_3559);
and U4027 (N_4027,N_3928,N_3503);
nor U4028 (N_4028,N_3701,N_3994);
or U4029 (N_4029,N_3731,N_3852);
xnor U4030 (N_4030,N_3843,N_3958);
or U4031 (N_4031,N_3567,N_3504);
or U4032 (N_4032,N_3987,N_3902);
and U4033 (N_4033,N_3622,N_3942);
xnor U4034 (N_4034,N_3914,N_3651);
nor U4035 (N_4035,N_3955,N_3853);
or U4036 (N_4036,N_3839,N_3703);
and U4037 (N_4037,N_3786,N_3740);
or U4038 (N_4038,N_3500,N_3600);
nor U4039 (N_4039,N_3789,N_3586);
or U4040 (N_4040,N_3913,N_3879);
xor U4041 (N_4041,N_3918,N_3822);
nand U4042 (N_4042,N_3501,N_3607);
xnor U4043 (N_4043,N_3937,N_3744);
or U4044 (N_4044,N_3564,N_3580);
and U4045 (N_4045,N_3718,N_3811);
xor U4046 (N_4046,N_3550,N_3907);
or U4047 (N_4047,N_3849,N_3830);
or U4048 (N_4048,N_3627,N_3604);
xor U4049 (N_4049,N_3923,N_3502);
and U4050 (N_4050,N_3516,N_3979);
or U4051 (N_4051,N_3870,N_3606);
or U4052 (N_4052,N_3750,N_3807);
and U4053 (N_4053,N_3927,N_3621);
and U4054 (N_4054,N_3966,N_3892);
nand U4055 (N_4055,N_3921,N_3792);
and U4056 (N_4056,N_3990,N_3774);
nor U4057 (N_4057,N_3755,N_3859);
xnor U4058 (N_4058,N_3934,N_3794);
nand U4059 (N_4059,N_3616,N_3730);
nand U4060 (N_4060,N_3542,N_3813);
nand U4061 (N_4061,N_3615,N_3825);
xor U4062 (N_4062,N_3814,N_3770);
xor U4063 (N_4063,N_3727,N_3880);
xor U4064 (N_4064,N_3737,N_3963);
nor U4065 (N_4065,N_3671,N_3687);
or U4066 (N_4066,N_3765,N_3534);
or U4067 (N_4067,N_3818,N_3574);
or U4068 (N_4068,N_3512,N_3526);
nand U4069 (N_4069,N_3575,N_3832);
xnor U4070 (N_4070,N_3635,N_3837);
or U4071 (N_4071,N_3595,N_3989);
or U4072 (N_4072,N_3901,N_3650);
xnor U4073 (N_4073,N_3612,N_3578);
or U4074 (N_4074,N_3809,N_3783);
xor U4075 (N_4075,N_3722,N_3777);
or U4076 (N_4076,N_3636,N_3652);
nor U4077 (N_4077,N_3509,N_3583);
nor U4078 (N_4078,N_3639,N_3508);
and U4079 (N_4079,N_3827,N_3897);
nand U4080 (N_4080,N_3977,N_3957);
xor U4081 (N_4081,N_3956,N_3898);
and U4082 (N_4082,N_3976,N_3728);
nor U4083 (N_4083,N_3557,N_3624);
nor U4084 (N_4084,N_3954,N_3647);
xor U4085 (N_4085,N_3781,N_3947);
xor U4086 (N_4086,N_3973,N_3514);
xnor U4087 (N_4087,N_3886,N_3552);
and U4088 (N_4088,N_3775,N_3510);
xor U4089 (N_4089,N_3721,N_3688);
nor U4090 (N_4090,N_3748,N_3716);
or U4091 (N_4091,N_3800,N_3533);
xor U4092 (N_4092,N_3563,N_3911);
and U4093 (N_4093,N_3823,N_3625);
xnor U4094 (N_4094,N_3637,N_3613);
xnor U4095 (N_4095,N_3890,N_3573);
or U4096 (N_4096,N_3538,N_3618);
xnor U4097 (N_4097,N_3626,N_3601);
nand U4098 (N_4098,N_3645,N_3819);
nor U4099 (N_4099,N_3702,N_3697);
nor U4100 (N_4100,N_3536,N_3521);
xnor U4101 (N_4101,N_3762,N_3706);
nor U4102 (N_4102,N_3922,N_3598);
xor U4103 (N_4103,N_3945,N_3812);
or U4104 (N_4104,N_3924,N_3910);
nor U4105 (N_4105,N_3848,N_3642);
xor U4106 (N_4106,N_3695,N_3760);
nor U4107 (N_4107,N_3638,N_3736);
and U4108 (N_4108,N_3798,N_3519);
nand U4109 (N_4109,N_3739,N_3677);
or U4110 (N_4110,N_3797,N_3816);
nor U4111 (N_4111,N_3588,N_3998);
or U4112 (N_4112,N_3566,N_3530);
or U4113 (N_4113,N_3541,N_3784);
or U4114 (N_4114,N_3864,N_3971);
or U4115 (N_4115,N_3930,N_3693);
nor U4116 (N_4116,N_3719,N_3929);
nor U4117 (N_4117,N_3527,N_3611);
nor U4118 (N_4118,N_3696,N_3558);
xor U4119 (N_4119,N_3658,N_3836);
xor U4120 (N_4120,N_3726,N_3883);
or U4121 (N_4121,N_3919,N_3745);
or U4122 (N_4122,N_3665,N_3632);
or U4123 (N_4123,N_3985,N_3948);
nor U4124 (N_4124,N_3756,N_3799);
or U4125 (N_4125,N_3565,N_3824);
nand U4126 (N_4126,N_3978,N_3614);
nand U4127 (N_4127,N_3655,N_3965);
xor U4128 (N_4128,N_3916,N_3953);
xnor U4129 (N_4129,N_3939,N_3734);
and U4130 (N_4130,N_3704,N_3513);
nand U4131 (N_4131,N_3815,N_3751);
or U4132 (N_4132,N_3943,N_3758);
or U4133 (N_4133,N_3708,N_3710);
or U4134 (N_4134,N_3866,N_3975);
and U4135 (N_4135,N_3788,N_3858);
nand U4136 (N_4136,N_3659,N_3617);
and U4137 (N_4137,N_3742,N_3868);
nand U4138 (N_4138,N_3969,N_3847);
and U4139 (N_4139,N_3991,N_3996);
or U4140 (N_4140,N_3999,N_3810);
and U4141 (N_4141,N_3713,N_3663);
nor U4142 (N_4142,N_3549,N_3608);
and U4143 (N_4143,N_3576,N_3780);
and U4144 (N_4144,N_3675,N_3838);
nor U4145 (N_4145,N_3850,N_3861);
nand U4146 (N_4146,N_3680,N_3917);
xor U4147 (N_4147,N_3562,N_3993);
nor U4148 (N_4148,N_3878,N_3628);
xnor U4149 (N_4149,N_3769,N_3944);
or U4150 (N_4150,N_3763,N_3796);
nor U4151 (N_4151,N_3946,N_3594);
nor U4152 (N_4152,N_3699,N_3553);
and U4153 (N_4153,N_3694,N_3511);
nor U4154 (N_4154,N_3666,N_3585);
xor U4155 (N_4155,N_3540,N_3603);
or U4156 (N_4156,N_3980,N_3941);
or U4157 (N_4157,N_3709,N_3662);
nor U4158 (N_4158,N_3757,N_3854);
or U4159 (N_4159,N_3808,N_3895);
nor U4160 (N_4160,N_3820,N_3685);
or U4161 (N_4161,N_3949,N_3525);
or U4162 (N_4162,N_3881,N_3754);
xor U4163 (N_4163,N_3556,N_3964);
nor U4164 (N_4164,N_3690,N_3972);
xnor U4165 (N_4165,N_3676,N_3717);
and U4166 (N_4166,N_3968,N_3899);
or U4167 (N_4167,N_3981,N_3587);
nand U4168 (N_4168,N_3873,N_3661);
nor U4169 (N_4169,N_3729,N_3962);
nor U4170 (N_4170,N_3782,N_3806);
nor U4171 (N_4171,N_3630,N_3790);
and U4172 (N_4172,N_3507,N_3747);
or U4173 (N_4173,N_3992,N_3700);
nor U4174 (N_4174,N_3982,N_3582);
or U4175 (N_4175,N_3560,N_3933);
and U4176 (N_4176,N_3936,N_3764);
or U4177 (N_4177,N_3874,N_3967);
nand U4178 (N_4178,N_3678,N_3579);
xnor U4179 (N_4179,N_3599,N_3766);
nor U4180 (N_4180,N_3749,N_3698);
and U4181 (N_4181,N_3610,N_3983);
and U4182 (N_4182,N_3932,N_3773);
and U4183 (N_4183,N_3970,N_3644);
and U4184 (N_4184,N_3768,N_3571);
or U4185 (N_4185,N_3593,N_3561);
nand U4186 (N_4186,N_3851,N_3844);
and U4187 (N_4187,N_3683,N_3506);
and U4188 (N_4188,N_3537,N_3759);
nand U4189 (N_4189,N_3785,N_3995);
or U4190 (N_4190,N_3570,N_3834);
and U4191 (N_4191,N_3988,N_3857);
and U4192 (N_4192,N_3884,N_3872);
or U4193 (N_4193,N_3997,N_3654);
nand U4194 (N_4194,N_3707,N_3860);
and U4195 (N_4195,N_3896,N_3631);
and U4196 (N_4196,N_3926,N_3532);
nand U4197 (N_4197,N_3674,N_3801);
and U4198 (N_4198,N_3778,N_3961);
nand U4199 (N_4199,N_3649,N_3705);
and U4200 (N_4200,N_3524,N_3891);
and U4201 (N_4201,N_3935,N_3672);
nor U4202 (N_4202,N_3545,N_3529);
xnor U4203 (N_4203,N_3605,N_3931);
or U4204 (N_4204,N_3776,N_3905);
and U4205 (N_4205,N_3555,N_3893);
or U4206 (N_4206,N_3539,N_3889);
nand U4207 (N_4207,N_3828,N_3940);
xor U4208 (N_4208,N_3920,N_3960);
or U4209 (N_4209,N_3826,N_3900);
and U4210 (N_4210,N_3629,N_3882);
or U4211 (N_4211,N_3528,N_3633);
nand U4212 (N_4212,N_3842,N_3865);
and U4213 (N_4213,N_3974,N_3720);
or U4214 (N_4214,N_3569,N_3546);
nor U4215 (N_4215,N_3572,N_3711);
nand U4216 (N_4216,N_3876,N_3589);
xnor U4217 (N_4217,N_3551,N_3925);
nor U4218 (N_4218,N_3597,N_3518);
xnor U4219 (N_4219,N_3846,N_3505);
and U4220 (N_4220,N_3648,N_3715);
and U4221 (N_4221,N_3623,N_3653);
or U4222 (N_4222,N_3795,N_3535);
xor U4223 (N_4223,N_3544,N_3887);
or U4224 (N_4224,N_3752,N_3771);
xor U4225 (N_4225,N_3554,N_3791);
xor U4226 (N_4226,N_3906,N_3669);
nor U4227 (N_4227,N_3829,N_3619);
nor U4228 (N_4228,N_3986,N_3670);
nor U4229 (N_4229,N_3833,N_3803);
or U4230 (N_4230,N_3831,N_3602);
and U4231 (N_4231,N_3735,N_3802);
xor U4232 (N_4232,N_3646,N_3845);
nor U4233 (N_4233,N_3684,N_3682);
nand U4234 (N_4234,N_3871,N_3548);
xor U4235 (N_4235,N_3520,N_3686);
or U4236 (N_4236,N_3679,N_3787);
nor U4237 (N_4237,N_3724,N_3908);
xor U4238 (N_4238,N_3959,N_3885);
and U4239 (N_4239,N_3877,N_3888);
nand U4240 (N_4240,N_3681,N_3804);
and U4241 (N_4241,N_3543,N_3668);
and U4242 (N_4242,N_3903,N_3712);
nor U4243 (N_4243,N_3592,N_3741);
nor U4244 (N_4244,N_3912,N_3577);
and U4245 (N_4245,N_3817,N_3951);
and U4246 (N_4246,N_3767,N_3664);
and U4247 (N_4247,N_3656,N_3609);
or U4248 (N_4248,N_3660,N_3692);
xnor U4249 (N_4249,N_3761,N_3667);
xor U4250 (N_4250,N_3753,N_3960);
nand U4251 (N_4251,N_3685,N_3854);
and U4252 (N_4252,N_3812,N_3604);
nor U4253 (N_4253,N_3656,N_3637);
xor U4254 (N_4254,N_3716,N_3508);
nand U4255 (N_4255,N_3621,N_3803);
or U4256 (N_4256,N_3860,N_3742);
xnor U4257 (N_4257,N_3849,N_3734);
nand U4258 (N_4258,N_3801,N_3671);
and U4259 (N_4259,N_3947,N_3884);
nand U4260 (N_4260,N_3610,N_3747);
nand U4261 (N_4261,N_3770,N_3877);
nor U4262 (N_4262,N_3806,N_3597);
nand U4263 (N_4263,N_3823,N_3587);
xnor U4264 (N_4264,N_3685,N_3715);
and U4265 (N_4265,N_3873,N_3663);
and U4266 (N_4266,N_3908,N_3590);
xnor U4267 (N_4267,N_3669,N_3930);
nand U4268 (N_4268,N_3523,N_3763);
or U4269 (N_4269,N_3865,N_3798);
or U4270 (N_4270,N_3930,N_3731);
or U4271 (N_4271,N_3955,N_3643);
or U4272 (N_4272,N_3960,N_3732);
and U4273 (N_4273,N_3899,N_3988);
nand U4274 (N_4274,N_3954,N_3725);
nand U4275 (N_4275,N_3534,N_3722);
nor U4276 (N_4276,N_3921,N_3586);
or U4277 (N_4277,N_3528,N_3547);
nor U4278 (N_4278,N_3796,N_3795);
or U4279 (N_4279,N_3805,N_3787);
xnor U4280 (N_4280,N_3954,N_3906);
or U4281 (N_4281,N_3847,N_3999);
nor U4282 (N_4282,N_3542,N_3960);
nor U4283 (N_4283,N_3799,N_3688);
nand U4284 (N_4284,N_3614,N_3724);
nor U4285 (N_4285,N_3937,N_3829);
or U4286 (N_4286,N_3881,N_3891);
xor U4287 (N_4287,N_3545,N_3914);
nand U4288 (N_4288,N_3810,N_3863);
or U4289 (N_4289,N_3807,N_3596);
or U4290 (N_4290,N_3591,N_3627);
or U4291 (N_4291,N_3627,N_3518);
nand U4292 (N_4292,N_3594,N_3702);
nand U4293 (N_4293,N_3933,N_3554);
nand U4294 (N_4294,N_3845,N_3827);
nor U4295 (N_4295,N_3854,N_3844);
nor U4296 (N_4296,N_3687,N_3790);
nand U4297 (N_4297,N_3990,N_3612);
nor U4298 (N_4298,N_3563,N_3714);
nor U4299 (N_4299,N_3969,N_3682);
nor U4300 (N_4300,N_3919,N_3654);
xnor U4301 (N_4301,N_3598,N_3588);
xor U4302 (N_4302,N_3964,N_3870);
nand U4303 (N_4303,N_3539,N_3883);
or U4304 (N_4304,N_3522,N_3852);
xor U4305 (N_4305,N_3910,N_3649);
nor U4306 (N_4306,N_3575,N_3530);
or U4307 (N_4307,N_3828,N_3906);
nor U4308 (N_4308,N_3776,N_3921);
nand U4309 (N_4309,N_3563,N_3915);
xor U4310 (N_4310,N_3944,N_3801);
nor U4311 (N_4311,N_3835,N_3545);
nor U4312 (N_4312,N_3859,N_3795);
or U4313 (N_4313,N_3660,N_3887);
and U4314 (N_4314,N_3504,N_3844);
xnor U4315 (N_4315,N_3597,N_3592);
nor U4316 (N_4316,N_3952,N_3931);
or U4317 (N_4317,N_3630,N_3911);
nand U4318 (N_4318,N_3558,N_3819);
xnor U4319 (N_4319,N_3812,N_3836);
or U4320 (N_4320,N_3729,N_3889);
nand U4321 (N_4321,N_3816,N_3514);
or U4322 (N_4322,N_3720,N_3822);
nand U4323 (N_4323,N_3736,N_3825);
and U4324 (N_4324,N_3601,N_3525);
nor U4325 (N_4325,N_3506,N_3925);
and U4326 (N_4326,N_3664,N_3534);
nand U4327 (N_4327,N_3524,N_3710);
and U4328 (N_4328,N_3541,N_3608);
nor U4329 (N_4329,N_3705,N_3635);
nand U4330 (N_4330,N_3895,N_3536);
xnor U4331 (N_4331,N_3694,N_3665);
nor U4332 (N_4332,N_3965,N_3688);
xor U4333 (N_4333,N_3891,N_3721);
and U4334 (N_4334,N_3672,N_3791);
nand U4335 (N_4335,N_3558,N_3850);
xor U4336 (N_4336,N_3941,N_3575);
or U4337 (N_4337,N_3778,N_3981);
and U4338 (N_4338,N_3737,N_3729);
nor U4339 (N_4339,N_3940,N_3853);
and U4340 (N_4340,N_3562,N_3996);
and U4341 (N_4341,N_3970,N_3556);
or U4342 (N_4342,N_3612,N_3773);
xor U4343 (N_4343,N_3596,N_3532);
nor U4344 (N_4344,N_3612,N_3980);
nand U4345 (N_4345,N_3975,N_3546);
xnor U4346 (N_4346,N_3662,N_3887);
xnor U4347 (N_4347,N_3818,N_3570);
xnor U4348 (N_4348,N_3872,N_3984);
nand U4349 (N_4349,N_3941,N_3594);
or U4350 (N_4350,N_3594,N_3895);
xnor U4351 (N_4351,N_3717,N_3532);
or U4352 (N_4352,N_3948,N_3544);
or U4353 (N_4353,N_3539,N_3588);
nand U4354 (N_4354,N_3919,N_3723);
and U4355 (N_4355,N_3772,N_3783);
xnor U4356 (N_4356,N_3944,N_3524);
xor U4357 (N_4357,N_3827,N_3990);
or U4358 (N_4358,N_3833,N_3504);
xnor U4359 (N_4359,N_3891,N_3980);
xnor U4360 (N_4360,N_3768,N_3921);
nand U4361 (N_4361,N_3844,N_3606);
nor U4362 (N_4362,N_3567,N_3754);
nand U4363 (N_4363,N_3626,N_3972);
xor U4364 (N_4364,N_3735,N_3639);
nor U4365 (N_4365,N_3875,N_3882);
and U4366 (N_4366,N_3685,N_3659);
nor U4367 (N_4367,N_3879,N_3607);
and U4368 (N_4368,N_3561,N_3689);
and U4369 (N_4369,N_3558,N_3554);
nand U4370 (N_4370,N_3652,N_3501);
nor U4371 (N_4371,N_3674,N_3625);
nand U4372 (N_4372,N_3923,N_3640);
nand U4373 (N_4373,N_3706,N_3527);
and U4374 (N_4374,N_3835,N_3711);
xor U4375 (N_4375,N_3984,N_3870);
xor U4376 (N_4376,N_3523,N_3711);
and U4377 (N_4377,N_3645,N_3830);
xnor U4378 (N_4378,N_3876,N_3586);
and U4379 (N_4379,N_3586,N_3763);
nor U4380 (N_4380,N_3553,N_3714);
and U4381 (N_4381,N_3845,N_3988);
and U4382 (N_4382,N_3561,N_3614);
nor U4383 (N_4383,N_3944,N_3908);
and U4384 (N_4384,N_3735,N_3530);
nor U4385 (N_4385,N_3979,N_3921);
or U4386 (N_4386,N_3840,N_3950);
nand U4387 (N_4387,N_3803,N_3838);
xor U4388 (N_4388,N_3566,N_3861);
nor U4389 (N_4389,N_3718,N_3857);
nor U4390 (N_4390,N_3953,N_3991);
and U4391 (N_4391,N_3690,N_3611);
or U4392 (N_4392,N_3612,N_3800);
xor U4393 (N_4393,N_3815,N_3562);
nor U4394 (N_4394,N_3798,N_3959);
nand U4395 (N_4395,N_3722,N_3762);
and U4396 (N_4396,N_3567,N_3843);
or U4397 (N_4397,N_3597,N_3624);
or U4398 (N_4398,N_3948,N_3572);
or U4399 (N_4399,N_3651,N_3881);
or U4400 (N_4400,N_3800,N_3883);
or U4401 (N_4401,N_3971,N_3614);
or U4402 (N_4402,N_3522,N_3918);
and U4403 (N_4403,N_3753,N_3547);
and U4404 (N_4404,N_3962,N_3847);
nor U4405 (N_4405,N_3503,N_3780);
nor U4406 (N_4406,N_3627,N_3687);
xnor U4407 (N_4407,N_3631,N_3584);
xor U4408 (N_4408,N_3524,N_3824);
nor U4409 (N_4409,N_3761,N_3923);
and U4410 (N_4410,N_3946,N_3820);
nand U4411 (N_4411,N_3528,N_3525);
or U4412 (N_4412,N_3817,N_3541);
nor U4413 (N_4413,N_3812,N_3530);
xor U4414 (N_4414,N_3742,N_3919);
nand U4415 (N_4415,N_3788,N_3789);
and U4416 (N_4416,N_3611,N_3808);
or U4417 (N_4417,N_3766,N_3603);
xnor U4418 (N_4418,N_3928,N_3684);
nor U4419 (N_4419,N_3565,N_3673);
and U4420 (N_4420,N_3810,N_3596);
nor U4421 (N_4421,N_3785,N_3709);
nor U4422 (N_4422,N_3826,N_3576);
nor U4423 (N_4423,N_3780,N_3772);
or U4424 (N_4424,N_3908,N_3522);
xnor U4425 (N_4425,N_3911,N_3726);
and U4426 (N_4426,N_3678,N_3581);
nand U4427 (N_4427,N_3751,N_3711);
and U4428 (N_4428,N_3679,N_3547);
nor U4429 (N_4429,N_3601,N_3722);
and U4430 (N_4430,N_3885,N_3526);
nand U4431 (N_4431,N_3893,N_3704);
nand U4432 (N_4432,N_3730,N_3755);
nor U4433 (N_4433,N_3510,N_3895);
nor U4434 (N_4434,N_3980,N_3513);
nand U4435 (N_4435,N_3929,N_3870);
or U4436 (N_4436,N_3519,N_3651);
or U4437 (N_4437,N_3869,N_3545);
nor U4438 (N_4438,N_3746,N_3723);
and U4439 (N_4439,N_3626,N_3874);
xor U4440 (N_4440,N_3799,N_3664);
and U4441 (N_4441,N_3727,N_3947);
xnor U4442 (N_4442,N_3826,N_3976);
nand U4443 (N_4443,N_3996,N_3921);
nor U4444 (N_4444,N_3903,N_3997);
and U4445 (N_4445,N_3997,N_3847);
nor U4446 (N_4446,N_3645,N_3554);
or U4447 (N_4447,N_3801,N_3542);
or U4448 (N_4448,N_3652,N_3704);
nor U4449 (N_4449,N_3591,N_3548);
xor U4450 (N_4450,N_3909,N_3685);
nand U4451 (N_4451,N_3545,N_3980);
or U4452 (N_4452,N_3523,N_3546);
or U4453 (N_4453,N_3881,N_3924);
or U4454 (N_4454,N_3706,N_3684);
nor U4455 (N_4455,N_3580,N_3804);
nand U4456 (N_4456,N_3642,N_3745);
nor U4457 (N_4457,N_3570,N_3749);
xnor U4458 (N_4458,N_3588,N_3983);
or U4459 (N_4459,N_3577,N_3842);
or U4460 (N_4460,N_3755,N_3686);
and U4461 (N_4461,N_3652,N_3860);
xnor U4462 (N_4462,N_3816,N_3539);
and U4463 (N_4463,N_3513,N_3921);
nand U4464 (N_4464,N_3746,N_3676);
xor U4465 (N_4465,N_3889,N_3634);
and U4466 (N_4466,N_3616,N_3569);
nor U4467 (N_4467,N_3632,N_3760);
or U4468 (N_4468,N_3790,N_3723);
nor U4469 (N_4469,N_3774,N_3726);
nor U4470 (N_4470,N_3581,N_3755);
and U4471 (N_4471,N_3997,N_3716);
nor U4472 (N_4472,N_3530,N_3629);
xnor U4473 (N_4473,N_3524,N_3858);
xnor U4474 (N_4474,N_3694,N_3571);
xnor U4475 (N_4475,N_3730,N_3682);
xor U4476 (N_4476,N_3571,N_3832);
nand U4477 (N_4477,N_3570,N_3710);
nand U4478 (N_4478,N_3707,N_3771);
nand U4479 (N_4479,N_3589,N_3822);
nand U4480 (N_4480,N_3509,N_3981);
nand U4481 (N_4481,N_3796,N_3658);
nor U4482 (N_4482,N_3869,N_3577);
and U4483 (N_4483,N_3647,N_3637);
xnor U4484 (N_4484,N_3976,N_3618);
nor U4485 (N_4485,N_3749,N_3884);
and U4486 (N_4486,N_3806,N_3826);
and U4487 (N_4487,N_3637,N_3917);
or U4488 (N_4488,N_3781,N_3830);
or U4489 (N_4489,N_3719,N_3969);
and U4490 (N_4490,N_3736,N_3500);
or U4491 (N_4491,N_3655,N_3885);
nor U4492 (N_4492,N_3584,N_3803);
or U4493 (N_4493,N_3979,N_3730);
or U4494 (N_4494,N_3500,N_3771);
xnor U4495 (N_4495,N_3701,N_3989);
nand U4496 (N_4496,N_3987,N_3763);
nand U4497 (N_4497,N_3671,N_3928);
or U4498 (N_4498,N_3872,N_3896);
or U4499 (N_4499,N_3959,N_3670);
or U4500 (N_4500,N_4260,N_4037);
xor U4501 (N_4501,N_4192,N_4278);
xor U4502 (N_4502,N_4333,N_4395);
or U4503 (N_4503,N_4332,N_4183);
or U4504 (N_4504,N_4447,N_4417);
nand U4505 (N_4505,N_4190,N_4067);
and U4506 (N_4506,N_4055,N_4053);
xnor U4507 (N_4507,N_4062,N_4164);
xor U4508 (N_4508,N_4083,N_4025);
nand U4509 (N_4509,N_4430,N_4357);
nand U4510 (N_4510,N_4097,N_4474);
or U4511 (N_4511,N_4234,N_4342);
and U4512 (N_4512,N_4271,N_4168);
or U4513 (N_4513,N_4216,N_4242);
nor U4514 (N_4514,N_4444,N_4470);
nand U4515 (N_4515,N_4004,N_4279);
nand U4516 (N_4516,N_4445,N_4026);
or U4517 (N_4517,N_4128,N_4132);
nand U4518 (N_4518,N_4370,N_4096);
or U4519 (N_4519,N_4018,N_4410);
nor U4520 (N_4520,N_4195,N_4496);
xnor U4521 (N_4521,N_4135,N_4283);
xnor U4522 (N_4522,N_4100,N_4339);
or U4523 (N_4523,N_4011,N_4274);
xnor U4524 (N_4524,N_4019,N_4034);
nor U4525 (N_4525,N_4375,N_4400);
nand U4526 (N_4526,N_4264,N_4323);
and U4527 (N_4527,N_4028,N_4251);
nor U4528 (N_4528,N_4494,N_4321);
nor U4529 (N_4529,N_4121,N_4194);
and U4530 (N_4530,N_4058,N_4127);
and U4531 (N_4531,N_4098,N_4404);
nor U4532 (N_4532,N_4080,N_4134);
or U4533 (N_4533,N_4463,N_4009);
and U4534 (N_4534,N_4180,N_4289);
nand U4535 (N_4535,N_4467,N_4078);
nor U4536 (N_4536,N_4262,N_4420);
xor U4537 (N_4537,N_4077,N_4220);
xor U4538 (N_4538,N_4191,N_4046);
xnor U4539 (N_4539,N_4306,N_4416);
xnor U4540 (N_4540,N_4189,N_4273);
or U4541 (N_4541,N_4305,N_4409);
and U4542 (N_4542,N_4297,N_4140);
xor U4543 (N_4543,N_4090,N_4287);
and U4544 (N_4544,N_4255,N_4272);
and U4545 (N_4545,N_4147,N_4117);
xnor U4546 (N_4546,N_4040,N_4143);
xnor U4547 (N_4547,N_4091,N_4405);
nand U4548 (N_4548,N_4330,N_4356);
nor U4549 (N_4549,N_4010,N_4182);
nor U4550 (N_4550,N_4466,N_4041);
or U4551 (N_4551,N_4099,N_4437);
or U4552 (N_4552,N_4173,N_4243);
nor U4553 (N_4553,N_4208,N_4406);
nor U4554 (N_4554,N_4031,N_4081);
nor U4555 (N_4555,N_4382,N_4086);
or U4556 (N_4556,N_4142,N_4365);
xnor U4557 (N_4557,N_4071,N_4257);
or U4558 (N_4558,N_4145,N_4222);
nor U4559 (N_4559,N_4263,N_4150);
and U4560 (N_4560,N_4448,N_4221);
nand U4561 (N_4561,N_4450,N_4172);
xnor U4562 (N_4562,N_4228,N_4157);
or U4563 (N_4563,N_4057,N_4211);
nor U4564 (N_4564,N_4105,N_4353);
or U4565 (N_4565,N_4452,N_4288);
and U4566 (N_4566,N_4389,N_4000);
and U4567 (N_4567,N_4472,N_4166);
or U4568 (N_4568,N_4475,N_4126);
and U4569 (N_4569,N_4468,N_4006);
nor U4570 (N_4570,N_4301,N_4350);
and U4571 (N_4571,N_4439,N_4207);
nor U4572 (N_4572,N_4200,N_4027);
and U4573 (N_4573,N_4314,N_4013);
and U4574 (N_4574,N_4313,N_4462);
xor U4575 (N_4575,N_4138,N_4317);
xnor U4576 (N_4576,N_4203,N_4245);
or U4577 (N_4577,N_4438,N_4109);
xnor U4578 (N_4578,N_4413,N_4129);
nand U4579 (N_4579,N_4252,N_4111);
nand U4580 (N_4580,N_4014,N_4493);
and U4581 (N_4581,N_4036,N_4137);
and U4582 (N_4582,N_4484,N_4181);
nand U4583 (N_4583,N_4104,N_4276);
nor U4584 (N_4584,N_4225,N_4331);
or U4585 (N_4585,N_4022,N_4295);
nor U4586 (N_4586,N_4372,N_4308);
nor U4587 (N_4587,N_4212,N_4315);
nor U4588 (N_4588,N_4311,N_4108);
nand U4589 (N_4589,N_4451,N_4478);
or U4590 (N_4590,N_4326,N_4328);
and U4591 (N_4591,N_4303,N_4015);
and U4592 (N_4592,N_4029,N_4177);
nor U4593 (N_4593,N_4284,N_4193);
xnor U4594 (N_4594,N_4116,N_4407);
or U4595 (N_4595,N_4052,N_4076);
or U4596 (N_4596,N_4453,N_4455);
and U4597 (N_4597,N_4369,N_4336);
nor U4598 (N_4598,N_4280,N_4123);
and U4599 (N_4599,N_4304,N_4151);
nand U4600 (N_4600,N_4256,N_4367);
xor U4601 (N_4601,N_4481,N_4073);
and U4602 (N_4602,N_4485,N_4039);
nand U4603 (N_4603,N_4477,N_4114);
nor U4604 (N_4604,N_4202,N_4032);
nand U4605 (N_4605,N_4310,N_4049);
nand U4606 (N_4606,N_4146,N_4258);
and U4607 (N_4607,N_4392,N_4411);
xnor U4608 (N_4608,N_4456,N_4275);
nor U4609 (N_4609,N_4153,N_4425);
and U4610 (N_4610,N_4363,N_4259);
and U4611 (N_4611,N_4060,N_4106);
nand U4612 (N_4612,N_4385,N_4423);
and U4613 (N_4613,N_4327,N_4435);
nor U4614 (N_4614,N_4377,N_4042);
xnor U4615 (N_4615,N_4307,N_4038);
nor U4616 (N_4616,N_4346,N_4139);
nor U4617 (N_4617,N_4464,N_4499);
nor U4618 (N_4618,N_4185,N_4473);
and U4619 (N_4619,N_4426,N_4337);
xor U4620 (N_4620,N_4254,N_4422);
xnor U4621 (N_4621,N_4270,N_4461);
nor U4622 (N_4622,N_4489,N_4112);
or U4623 (N_4623,N_4092,N_4159);
nand U4624 (N_4624,N_4249,N_4240);
nand U4625 (N_4625,N_4329,N_4209);
and U4626 (N_4626,N_4075,N_4204);
xnor U4627 (N_4627,N_4383,N_4088);
xnor U4628 (N_4628,N_4047,N_4084);
and U4629 (N_4629,N_4324,N_4379);
and U4630 (N_4630,N_4428,N_4397);
nand U4631 (N_4631,N_4446,N_4196);
and U4632 (N_4632,N_4399,N_4424);
and U4633 (N_4633,N_4393,N_4162);
xnor U4634 (N_4634,N_4286,N_4418);
xnor U4635 (N_4635,N_4005,N_4267);
xnor U4636 (N_4636,N_4441,N_4197);
and U4637 (N_4637,N_4226,N_4050);
nand U4638 (N_4638,N_4188,N_4497);
nand U4639 (N_4639,N_4246,N_4002);
or U4640 (N_4640,N_4224,N_4170);
or U4641 (N_4641,N_4349,N_4338);
and U4642 (N_4642,N_4219,N_4089);
nor U4643 (N_4643,N_4431,N_4231);
nand U4644 (N_4644,N_4210,N_4459);
nand U4645 (N_4645,N_4229,N_4239);
nand U4646 (N_4646,N_4309,N_4347);
xnor U4647 (N_4647,N_4381,N_4486);
nand U4648 (N_4648,N_4218,N_4061);
nor U4649 (N_4649,N_4348,N_4119);
xnor U4650 (N_4650,N_4113,N_4294);
and U4651 (N_4651,N_4175,N_4103);
or U4652 (N_4652,N_4325,N_4176);
or U4653 (N_4653,N_4244,N_4107);
nor U4654 (N_4654,N_4386,N_4390);
and U4655 (N_4655,N_4487,N_4199);
or U4656 (N_4656,N_4415,N_4238);
or U4657 (N_4657,N_4449,N_4457);
nor U4658 (N_4658,N_4482,N_4490);
xnor U4659 (N_4659,N_4359,N_4102);
nor U4660 (N_4660,N_4265,N_4133);
nor U4661 (N_4661,N_4118,N_4394);
xnor U4662 (N_4662,N_4201,N_4023);
nand U4663 (N_4663,N_4085,N_4291);
nand U4664 (N_4664,N_4414,N_4371);
or U4665 (N_4665,N_4035,N_4269);
or U4666 (N_4666,N_4033,N_4261);
nor U4667 (N_4667,N_4072,N_4312);
or U4668 (N_4668,N_4427,N_4095);
and U4669 (N_4669,N_4454,N_4421);
and U4670 (N_4670,N_4458,N_4378);
nor U4671 (N_4671,N_4178,N_4056);
or U4672 (N_4672,N_4292,N_4282);
and U4673 (N_4673,N_4302,N_4479);
xnor U4674 (N_4674,N_4412,N_4131);
nand U4675 (N_4675,N_4087,N_4024);
nand U4676 (N_4676,N_4322,N_4169);
nand U4677 (N_4677,N_4094,N_4008);
nand U4678 (N_4678,N_4167,N_4429);
and U4679 (N_4679,N_4293,N_4360);
or U4680 (N_4680,N_4277,N_4124);
xor U4681 (N_4681,N_4480,N_4374);
nor U4682 (N_4682,N_4115,N_4398);
nand U4683 (N_4683,N_4161,N_4043);
nand U4684 (N_4684,N_4433,N_4391);
and U4685 (N_4685,N_4290,N_4373);
xor U4686 (N_4686,N_4432,N_4299);
and U4687 (N_4687,N_4149,N_4232);
xor U4688 (N_4688,N_4044,N_4155);
and U4689 (N_4689,N_4401,N_4334);
nor U4690 (N_4690,N_4492,N_4048);
nor U4691 (N_4691,N_4122,N_4384);
and U4692 (N_4692,N_4074,N_4030);
and U4693 (N_4693,N_4465,N_4165);
xor U4694 (N_4694,N_4408,N_4021);
nand U4695 (N_4695,N_4236,N_4316);
xor U4696 (N_4696,N_4483,N_4434);
and U4697 (N_4697,N_4174,N_4355);
nand U4698 (N_4698,N_4110,N_4380);
and U4699 (N_4699,N_4476,N_4186);
and U4700 (N_4700,N_4362,N_4051);
xnor U4701 (N_4701,N_4233,N_4230);
xor U4702 (N_4702,N_4156,N_4498);
and U4703 (N_4703,N_4388,N_4012);
and U4704 (N_4704,N_4340,N_4247);
xnor U4705 (N_4705,N_4064,N_4136);
and U4706 (N_4706,N_4396,N_4361);
nand U4707 (N_4707,N_4152,N_4069);
nor U4708 (N_4708,N_4351,N_4419);
nand U4709 (N_4709,N_4491,N_4001);
and U4710 (N_4710,N_4068,N_4079);
and U4711 (N_4711,N_4460,N_4266);
xor U4712 (N_4712,N_4045,N_4059);
or U4713 (N_4713,N_4187,N_4184);
or U4714 (N_4714,N_4120,N_4148);
or U4715 (N_4715,N_4471,N_4368);
and U4716 (N_4716,N_4341,N_4366);
nand U4717 (N_4717,N_4130,N_4281);
and U4718 (N_4718,N_4125,N_4319);
nor U4719 (N_4719,N_4402,N_4007);
nor U4720 (N_4720,N_4354,N_4345);
or U4721 (N_4721,N_4440,N_4248);
or U4722 (N_4722,N_4285,N_4344);
nor U4723 (N_4723,N_4154,N_4158);
or U4724 (N_4724,N_4442,N_4387);
and U4725 (N_4725,N_4237,N_4054);
and U4726 (N_4726,N_4101,N_4320);
and U4727 (N_4727,N_4436,N_4241);
xnor U4728 (N_4728,N_4358,N_4198);
nand U4729 (N_4729,N_4093,N_4250);
or U4730 (N_4730,N_4495,N_4017);
nand U4731 (N_4731,N_4070,N_4335);
nor U4732 (N_4732,N_4065,N_4443);
xnor U4733 (N_4733,N_4205,N_4300);
nand U4734 (N_4734,N_4020,N_4343);
or U4735 (N_4735,N_4235,N_4376);
xor U4736 (N_4736,N_4063,N_4144);
or U4737 (N_4737,N_4214,N_4082);
nor U4738 (N_4738,N_4163,N_4213);
nor U4739 (N_4739,N_4217,N_4160);
nor U4740 (N_4740,N_4179,N_4469);
or U4741 (N_4741,N_4227,N_4268);
xor U4742 (N_4742,N_4364,N_4003);
xor U4743 (N_4743,N_4488,N_4352);
or U4744 (N_4744,N_4318,N_4066);
nor U4745 (N_4745,N_4403,N_4298);
xnor U4746 (N_4746,N_4223,N_4171);
and U4747 (N_4747,N_4206,N_4141);
and U4748 (N_4748,N_4253,N_4215);
and U4749 (N_4749,N_4296,N_4016);
and U4750 (N_4750,N_4268,N_4220);
nor U4751 (N_4751,N_4480,N_4385);
nor U4752 (N_4752,N_4458,N_4497);
nor U4753 (N_4753,N_4176,N_4083);
nand U4754 (N_4754,N_4448,N_4310);
nor U4755 (N_4755,N_4472,N_4125);
and U4756 (N_4756,N_4359,N_4320);
xnor U4757 (N_4757,N_4228,N_4207);
and U4758 (N_4758,N_4020,N_4075);
nand U4759 (N_4759,N_4024,N_4056);
nand U4760 (N_4760,N_4033,N_4136);
or U4761 (N_4761,N_4238,N_4214);
and U4762 (N_4762,N_4224,N_4341);
xor U4763 (N_4763,N_4342,N_4458);
xor U4764 (N_4764,N_4073,N_4036);
nor U4765 (N_4765,N_4250,N_4434);
and U4766 (N_4766,N_4034,N_4120);
nor U4767 (N_4767,N_4499,N_4433);
nand U4768 (N_4768,N_4137,N_4425);
nand U4769 (N_4769,N_4342,N_4481);
and U4770 (N_4770,N_4325,N_4097);
or U4771 (N_4771,N_4386,N_4408);
xnor U4772 (N_4772,N_4105,N_4045);
and U4773 (N_4773,N_4153,N_4285);
and U4774 (N_4774,N_4007,N_4336);
or U4775 (N_4775,N_4483,N_4431);
and U4776 (N_4776,N_4114,N_4452);
or U4777 (N_4777,N_4158,N_4082);
or U4778 (N_4778,N_4057,N_4422);
nor U4779 (N_4779,N_4342,N_4477);
nor U4780 (N_4780,N_4392,N_4102);
and U4781 (N_4781,N_4149,N_4018);
nand U4782 (N_4782,N_4031,N_4315);
xor U4783 (N_4783,N_4084,N_4477);
or U4784 (N_4784,N_4242,N_4269);
nor U4785 (N_4785,N_4257,N_4120);
nor U4786 (N_4786,N_4487,N_4437);
nor U4787 (N_4787,N_4319,N_4081);
nand U4788 (N_4788,N_4106,N_4341);
or U4789 (N_4789,N_4279,N_4341);
xnor U4790 (N_4790,N_4204,N_4425);
and U4791 (N_4791,N_4054,N_4273);
and U4792 (N_4792,N_4353,N_4372);
and U4793 (N_4793,N_4127,N_4350);
xor U4794 (N_4794,N_4094,N_4128);
nand U4795 (N_4795,N_4009,N_4348);
and U4796 (N_4796,N_4465,N_4295);
xor U4797 (N_4797,N_4008,N_4205);
xor U4798 (N_4798,N_4005,N_4150);
and U4799 (N_4799,N_4384,N_4311);
xor U4800 (N_4800,N_4377,N_4242);
xor U4801 (N_4801,N_4370,N_4166);
or U4802 (N_4802,N_4043,N_4260);
nand U4803 (N_4803,N_4187,N_4365);
nor U4804 (N_4804,N_4453,N_4313);
nand U4805 (N_4805,N_4235,N_4085);
or U4806 (N_4806,N_4071,N_4141);
nor U4807 (N_4807,N_4189,N_4012);
nand U4808 (N_4808,N_4256,N_4158);
xnor U4809 (N_4809,N_4481,N_4065);
or U4810 (N_4810,N_4256,N_4239);
nand U4811 (N_4811,N_4368,N_4115);
nand U4812 (N_4812,N_4187,N_4060);
nor U4813 (N_4813,N_4461,N_4020);
nor U4814 (N_4814,N_4146,N_4154);
or U4815 (N_4815,N_4075,N_4039);
nor U4816 (N_4816,N_4428,N_4432);
or U4817 (N_4817,N_4336,N_4268);
or U4818 (N_4818,N_4085,N_4481);
or U4819 (N_4819,N_4153,N_4016);
nand U4820 (N_4820,N_4165,N_4068);
and U4821 (N_4821,N_4113,N_4146);
nand U4822 (N_4822,N_4114,N_4252);
nor U4823 (N_4823,N_4105,N_4164);
nand U4824 (N_4824,N_4147,N_4250);
xor U4825 (N_4825,N_4142,N_4273);
or U4826 (N_4826,N_4487,N_4267);
and U4827 (N_4827,N_4149,N_4314);
nor U4828 (N_4828,N_4115,N_4053);
and U4829 (N_4829,N_4085,N_4286);
or U4830 (N_4830,N_4358,N_4146);
nor U4831 (N_4831,N_4319,N_4182);
nor U4832 (N_4832,N_4414,N_4256);
and U4833 (N_4833,N_4258,N_4175);
nand U4834 (N_4834,N_4176,N_4264);
xor U4835 (N_4835,N_4104,N_4089);
nand U4836 (N_4836,N_4316,N_4434);
or U4837 (N_4837,N_4362,N_4298);
nor U4838 (N_4838,N_4045,N_4054);
xnor U4839 (N_4839,N_4470,N_4316);
xor U4840 (N_4840,N_4451,N_4075);
and U4841 (N_4841,N_4111,N_4408);
or U4842 (N_4842,N_4315,N_4472);
nor U4843 (N_4843,N_4395,N_4497);
nor U4844 (N_4844,N_4248,N_4095);
xnor U4845 (N_4845,N_4462,N_4222);
nor U4846 (N_4846,N_4069,N_4307);
and U4847 (N_4847,N_4114,N_4186);
xor U4848 (N_4848,N_4100,N_4406);
nor U4849 (N_4849,N_4111,N_4064);
or U4850 (N_4850,N_4032,N_4286);
xor U4851 (N_4851,N_4108,N_4044);
and U4852 (N_4852,N_4297,N_4332);
nor U4853 (N_4853,N_4193,N_4268);
nand U4854 (N_4854,N_4096,N_4164);
nand U4855 (N_4855,N_4369,N_4155);
and U4856 (N_4856,N_4048,N_4200);
nor U4857 (N_4857,N_4286,N_4168);
nor U4858 (N_4858,N_4237,N_4493);
xor U4859 (N_4859,N_4479,N_4029);
nor U4860 (N_4860,N_4213,N_4379);
xnor U4861 (N_4861,N_4182,N_4482);
or U4862 (N_4862,N_4098,N_4018);
nor U4863 (N_4863,N_4311,N_4178);
xor U4864 (N_4864,N_4449,N_4259);
or U4865 (N_4865,N_4179,N_4115);
nor U4866 (N_4866,N_4129,N_4234);
and U4867 (N_4867,N_4438,N_4407);
xor U4868 (N_4868,N_4194,N_4004);
and U4869 (N_4869,N_4285,N_4037);
or U4870 (N_4870,N_4320,N_4121);
nor U4871 (N_4871,N_4178,N_4449);
xnor U4872 (N_4872,N_4446,N_4120);
and U4873 (N_4873,N_4367,N_4203);
nor U4874 (N_4874,N_4490,N_4363);
xnor U4875 (N_4875,N_4295,N_4433);
or U4876 (N_4876,N_4218,N_4014);
nand U4877 (N_4877,N_4447,N_4480);
nor U4878 (N_4878,N_4004,N_4229);
xnor U4879 (N_4879,N_4483,N_4407);
nor U4880 (N_4880,N_4130,N_4030);
nand U4881 (N_4881,N_4366,N_4126);
xor U4882 (N_4882,N_4293,N_4390);
xor U4883 (N_4883,N_4311,N_4058);
nor U4884 (N_4884,N_4357,N_4079);
nor U4885 (N_4885,N_4187,N_4024);
nand U4886 (N_4886,N_4000,N_4304);
nand U4887 (N_4887,N_4212,N_4439);
or U4888 (N_4888,N_4082,N_4039);
and U4889 (N_4889,N_4320,N_4302);
xor U4890 (N_4890,N_4200,N_4493);
and U4891 (N_4891,N_4113,N_4249);
nand U4892 (N_4892,N_4449,N_4450);
nand U4893 (N_4893,N_4363,N_4450);
xnor U4894 (N_4894,N_4213,N_4290);
and U4895 (N_4895,N_4489,N_4175);
or U4896 (N_4896,N_4454,N_4343);
xnor U4897 (N_4897,N_4044,N_4258);
xor U4898 (N_4898,N_4412,N_4236);
xnor U4899 (N_4899,N_4498,N_4260);
nand U4900 (N_4900,N_4206,N_4178);
and U4901 (N_4901,N_4023,N_4291);
and U4902 (N_4902,N_4189,N_4258);
nand U4903 (N_4903,N_4445,N_4345);
nand U4904 (N_4904,N_4278,N_4157);
nor U4905 (N_4905,N_4440,N_4127);
nor U4906 (N_4906,N_4450,N_4048);
and U4907 (N_4907,N_4493,N_4147);
xor U4908 (N_4908,N_4467,N_4026);
xnor U4909 (N_4909,N_4324,N_4418);
xor U4910 (N_4910,N_4291,N_4152);
xor U4911 (N_4911,N_4189,N_4295);
nor U4912 (N_4912,N_4159,N_4490);
nor U4913 (N_4913,N_4371,N_4276);
nor U4914 (N_4914,N_4498,N_4338);
or U4915 (N_4915,N_4227,N_4301);
and U4916 (N_4916,N_4157,N_4096);
nand U4917 (N_4917,N_4175,N_4340);
and U4918 (N_4918,N_4455,N_4493);
and U4919 (N_4919,N_4360,N_4345);
nor U4920 (N_4920,N_4345,N_4137);
nor U4921 (N_4921,N_4072,N_4248);
and U4922 (N_4922,N_4170,N_4390);
nor U4923 (N_4923,N_4193,N_4368);
and U4924 (N_4924,N_4172,N_4217);
or U4925 (N_4925,N_4364,N_4081);
xor U4926 (N_4926,N_4411,N_4453);
nand U4927 (N_4927,N_4071,N_4034);
nor U4928 (N_4928,N_4463,N_4476);
xnor U4929 (N_4929,N_4305,N_4122);
nor U4930 (N_4930,N_4183,N_4202);
or U4931 (N_4931,N_4335,N_4446);
nand U4932 (N_4932,N_4276,N_4171);
or U4933 (N_4933,N_4081,N_4156);
and U4934 (N_4934,N_4211,N_4386);
and U4935 (N_4935,N_4064,N_4332);
nor U4936 (N_4936,N_4220,N_4193);
nor U4937 (N_4937,N_4388,N_4336);
nand U4938 (N_4938,N_4027,N_4332);
and U4939 (N_4939,N_4250,N_4321);
xnor U4940 (N_4940,N_4313,N_4063);
nor U4941 (N_4941,N_4249,N_4330);
xor U4942 (N_4942,N_4068,N_4001);
nor U4943 (N_4943,N_4216,N_4232);
nor U4944 (N_4944,N_4473,N_4140);
xnor U4945 (N_4945,N_4340,N_4213);
or U4946 (N_4946,N_4183,N_4124);
nand U4947 (N_4947,N_4433,N_4302);
or U4948 (N_4948,N_4241,N_4225);
xnor U4949 (N_4949,N_4215,N_4465);
nand U4950 (N_4950,N_4051,N_4378);
and U4951 (N_4951,N_4441,N_4396);
or U4952 (N_4952,N_4318,N_4391);
xor U4953 (N_4953,N_4416,N_4252);
or U4954 (N_4954,N_4044,N_4112);
nand U4955 (N_4955,N_4074,N_4378);
and U4956 (N_4956,N_4166,N_4034);
and U4957 (N_4957,N_4245,N_4295);
or U4958 (N_4958,N_4111,N_4441);
and U4959 (N_4959,N_4047,N_4442);
or U4960 (N_4960,N_4178,N_4026);
xor U4961 (N_4961,N_4297,N_4110);
or U4962 (N_4962,N_4049,N_4200);
nand U4963 (N_4963,N_4379,N_4134);
or U4964 (N_4964,N_4458,N_4128);
nand U4965 (N_4965,N_4208,N_4156);
nor U4966 (N_4966,N_4203,N_4071);
xor U4967 (N_4967,N_4001,N_4311);
nand U4968 (N_4968,N_4034,N_4188);
xnor U4969 (N_4969,N_4014,N_4447);
xor U4970 (N_4970,N_4182,N_4317);
or U4971 (N_4971,N_4429,N_4490);
nand U4972 (N_4972,N_4321,N_4239);
xor U4973 (N_4973,N_4053,N_4108);
nand U4974 (N_4974,N_4435,N_4271);
and U4975 (N_4975,N_4250,N_4291);
nand U4976 (N_4976,N_4324,N_4151);
nor U4977 (N_4977,N_4290,N_4031);
xnor U4978 (N_4978,N_4113,N_4445);
nand U4979 (N_4979,N_4011,N_4260);
nor U4980 (N_4980,N_4174,N_4442);
nor U4981 (N_4981,N_4490,N_4192);
and U4982 (N_4982,N_4339,N_4352);
nor U4983 (N_4983,N_4307,N_4033);
xnor U4984 (N_4984,N_4461,N_4392);
nor U4985 (N_4985,N_4167,N_4060);
xor U4986 (N_4986,N_4147,N_4350);
nand U4987 (N_4987,N_4177,N_4286);
and U4988 (N_4988,N_4340,N_4323);
nand U4989 (N_4989,N_4072,N_4170);
nand U4990 (N_4990,N_4033,N_4163);
nand U4991 (N_4991,N_4134,N_4007);
or U4992 (N_4992,N_4095,N_4160);
nor U4993 (N_4993,N_4495,N_4456);
or U4994 (N_4994,N_4114,N_4410);
and U4995 (N_4995,N_4377,N_4429);
nor U4996 (N_4996,N_4434,N_4032);
and U4997 (N_4997,N_4456,N_4144);
xor U4998 (N_4998,N_4262,N_4292);
and U4999 (N_4999,N_4176,N_4207);
and U5000 (N_5000,N_4653,N_4987);
nand U5001 (N_5001,N_4569,N_4608);
and U5002 (N_5002,N_4756,N_4913);
xor U5003 (N_5003,N_4500,N_4627);
or U5004 (N_5004,N_4744,N_4914);
and U5005 (N_5005,N_4945,N_4741);
and U5006 (N_5006,N_4875,N_4957);
and U5007 (N_5007,N_4534,N_4934);
nand U5008 (N_5008,N_4678,N_4975);
xnor U5009 (N_5009,N_4733,N_4859);
and U5010 (N_5010,N_4713,N_4829);
nand U5011 (N_5011,N_4911,N_4916);
nand U5012 (N_5012,N_4867,N_4902);
or U5013 (N_5013,N_4577,N_4929);
xnor U5014 (N_5014,N_4587,N_4662);
nand U5015 (N_5015,N_4924,N_4621);
nand U5016 (N_5016,N_4755,N_4827);
or U5017 (N_5017,N_4887,N_4894);
or U5018 (N_5018,N_4882,N_4920);
nand U5019 (N_5019,N_4554,N_4697);
nand U5020 (N_5020,N_4922,N_4556);
nor U5021 (N_5021,N_4823,N_4617);
xor U5022 (N_5022,N_4630,N_4502);
nand U5023 (N_5023,N_4970,N_4580);
and U5024 (N_5024,N_4901,N_4763);
xnor U5025 (N_5025,N_4739,N_4611);
nand U5026 (N_5026,N_4984,N_4988);
nand U5027 (N_5027,N_4535,N_4948);
nand U5028 (N_5028,N_4863,N_4727);
nor U5029 (N_5029,N_4681,N_4512);
nand U5030 (N_5030,N_4819,N_4790);
or U5031 (N_5031,N_4700,N_4707);
nand U5032 (N_5032,N_4889,N_4895);
and U5033 (N_5033,N_4812,N_4985);
and U5034 (N_5034,N_4892,N_4563);
nand U5035 (N_5035,N_4710,N_4840);
or U5036 (N_5036,N_4719,N_4677);
or U5037 (N_5037,N_4848,N_4992);
or U5038 (N_5038,N_4631,N_4915);
nor U5039 (N_5039,N_4644,N_4619);
nor U5040 (N_5040,N_4952,N_4841);
and U5041 (N_5041,N_4699,N_4981);
xnor U5042 (N_5042,N_4717,N_4565);
and U5043 (N_5043,N_4628,N_4856);
or U5044 (N_5044,N_4849,N_4966);
nand U5045 (N_5045,N_4685,N_4560);
xor U5046 (N_5046,N_4590,N_4964);
nand U5047 (N_5047,N_4711,N_4573);
xnor U5048 (N_5048,N_4839,N_4938);
xnor U5049 (N_5049,N_4650,N_4602);
or U5050 (N_5050,N_4910,N_4735);
nand U5051 (N_5051,N_4998,N_4657);
xor U5052 (N_5052,N_4523,N_4624);
nor U5053 (N_5053,N_4972,N_4898);
or U5054 (N_5054,N_4629,N_4956);
nand U5055 (N_5055,N_4568,N_4990);
xor U5056 (N_5056,N_4521,N_4724);
nand U5057 (N_5057,N_4664,N_4557);
nand U5058 (N_5058,N_4991,N_4514);
nand U5059 (N_5059,N_4953,N_4814);
and U5060 (N_5060,N_4708,N_4809);
or U5061 (N_5061,N_4919,N_4676);
nand U5062 (N_5062,N_4638,N_4932);
or U5063 (N_5063,N_4963,N_4528);
and U5064 (N_5064,N_4779,N_4515);
and U5065 (N_5065,N_4738,N_4601);
xor U5066 (N_5066,N_4616,N_4722);
xor U5067 (N_5067,N_4674,N_4960);
nor U5068 (N_5068,N_4788,N_4586);
nand U5069 (N_5069,N_4643,N_4761);
nor U5070 (N_5070,N_4931,N_4885);
nor U5071 (N_5071,N_4530,N_4725);
nand U5072 (N_5072,N_4647,N_4706);
nor U5073 (N_5073,N_4547,N_4858);
nand U5074 (N_5074,N_4787,N_4747);
nand U5075 (N_5075,N_4749,N_4552);
nor U5076 (N_5076,N_4874,N_4965);
xnor U5077 (N_5077,N_4730,N_4670);
xor U5078 (N_5078,N_4933,N_4632);
xnor U5079 (N_5079,N_4750,N_4732);
nor U5080 (N_5080,N_4857,N_4594);
nand U5081 (N_5081,N_4831,N_4701);
xnor U5082 (N_5082,N_4789,N_4836);
nor U5083 (N_5083,N_4751,N_4891);
nand U5084 (N_5084,N_4811,N_4773);
or U5085 (N_5085,N_4654,N_4687);
and U5086 (N_5086,N_4620,N_4529);
and U5087 (N_5087,N_4806,N_4612);
nor U5088 (N_5088,N_4917,N_4539);
nor U5089 (N_5089,N_4548,N_4704);
or U5090 (N_5090,N_4908,N_4683);
xor U5091 (N_5091,N_4610,N_4757);
nand U5092 (N_5092,N_4595,N_4899);
or U5093 (N_5093,N_4516,N_4625);
xnor U5094 (N_5094,N_4559,N_4513);
and U5095 (N_5095,N_4698,N_4663);
nor U5096 (N_5096,N_4690,N_4748);
and U5097 (N_5097,N_4682,N_4838);
nor U5098 (N_5098,N_4506,N_4684);
and U5099 (N_5099,N_4967,N_4928);
or U5100 (N_5100,N_4549,N_4696);
or U5101 (N_5101,N_4871,N_4959);
nand U5102 (N_5102,N_4776,N_4770);
nor U5103 (N_5103,N_4614,N_4589);
xor U5104 (N_5104,N_4525,N_4607);
or U5105 (N_5105,N_4833,N_4927);
nand U5106 (N_5106,N_4646,N_4883);
nand U5107 (N_5107,N_4937,N_4845);
nand U5108 (N_5108,N_4842,N_4855);
or U5109 (N_5109,N_4762,N_4921);
xor U5110 (N_5110,N_4862,N_4983);
and U5111 (N_5111,N_4672,N_4656);
nor U5112 (N_5112,N_4718,N_4618);
nor U5113 (N_5113,N_4571,N_4692);
and U5114 (N_5114,N_4879,N_4907);
or U5115 (N_5115,N_4782,N_4830);
nor U5116 (N_5116,N_4906,N_4726);
xnor U5117 (N_5117,N_4815,N_4796);
and U5118 (N_5118,N_4760,N_4888);
and U5119 (N_5119,N_4832,N_4818);
nor U5120 (N_5120,N_4716,N_4604);
xor U5121 (N_5121,N_4872,N_4686);
and U5122 (N_5122,N_4508,N_4799);
xnor U5123 (N_5123,N_4997,N_4540);
nor U5124 (N_5124,N_4825,N_4731);
and U5125 (N_5125,N_4843,N_4923);
nor U5126 (N_5126,N_4742,N_4802);
and U5127 (N_5127,N_4543,N_4926);
nand U5128 (N_5128,N_4769,N_4942);
and U5129 (N_5129,N_4592,N_4962);
or U5130 (N_5130,N_4768,N_4979);
nor U5131 (N_5131,N_4775,N_4994);
and U5132 (N_5132,N_4582,N_4579);
nand U5133 (N_5133,N_4864,N_4820);
or U5134 (N_5134,N_4572,N_4645);
nand U5135 (N_5135,N_4941,N_4736);
xnor U5136 (N_5136,N_4581,N_4740);
xnor U5137 (N_5137,N_4961,N_4835);
nand U5138 (N_5138,N_4993,N_4780);
and U5139 (N_5139,N_4860,N_4566);
xnor U5140 (N_5140,N_4537,N_4570);
and U5141 (N_5141,N_4821,N_4847);
nor U5142 (N_5142,N_4752,N_4615);
xor U5143 (N_5143,N_4712,N_4852);
nand U5144 (N_5144,N_4791,N_4526);
nand U5145 (N_5145,N_4890,N_4669);
nand U5146 (N_5146,N_4642,N_4605);
xor U5147 (N_5147,N_4817,N_4743);
xnor U5148 (N_5148,N_4986,N_4652);
xor U5149 (N_5149,N_4764,N_4969);
xor U5150 (N_5150,N_4505,N_4520);
nand U5151 (N_5151,N_4801,N_4828);
xnor U5152 (N_5152,N_4511,N_4754);
xor U5153 (N_5153,N_4714,N_4596);
xor U5154 (N_5154,N_4772,N_4968);
nor U5155 (N_5155,N_4804,N_4781);
or U5156 (N_5156,N_4777,N_4971);
or U5157 (N_5157,N_4824,N_4778);
xor U5158 (N_5158,N_4974,N_4689);
nand U5159 (N_5159,N_4658,N_4784);
and U5160 (N_5160,N_4637,N_4536);
nor U5161 (N_5161,N_4576,N_4567);
and U5162 (N_5162,N_4649,N_4542);
xor U5163 (N_5163,N_4854,N_4504);
nand U5164 (N_5164,N_4622,N_4798);
nor U5165 (N_5165,N_4999,N_4583);
and U5166 (N_5166,N_4640,N_4765);
xnor U5167 (N_5167,N_4939,N_4794);
nand U5168 (N_5168,N_4510,N_4976);
nand U5169 (N_5169,N_4869,N_4723);
or U5170 (N_5170,N_4980,N_4878);
or U5171 (N_5171,N_4578,N_4667);
xnor U5172 (N_5172,N_4673,N_4977);
and U5173 (N_5173,N_4598,N_4729);
xnor U5174 (N_5174,N_4593,N_4606);
or U5175 (N_5175,N_4655,N_4588);
nor U5176 (N_5176,N_4517,N_4721);
nand U5177 (N_5177,N_4575,N_4603);
nand U5178 (N_5178,N_4861,N_4865);
xor U5179 (N_5179,N_4786,N_4703);
nand U5180 (N_5180,N_4648,N_4944);
or U5181 (N_5181,N_4954,N_4550);
nand U5182 (N_5182,N_4635,N_4533);
nor U5183 (N_5183,N_4745,N_4715);
or U5184 (N_5184,N_4936,N_4800);
or U5185 (N_5185,N_4783,N_4955);
xor U5186 (N_5186,N_4702,N_4626);
nand U5187 (N_5187,N_4759,N_4884);
and U5188 (N_5188,N_4519,N_4893);
and U5189 (N_5189,N_4584,N_4978);
nor U5190 (N_5190,N_4558,N_4767);
nor U5191 (N_5191,N_4774,N_4940);
xnor U5192 (N_5192,N_4989,N_4679);
or U5193 (N_5193,N_4501,N_4668);
and U5194 (N_5194,N_4973,N_4561);
or U5195 (N_5195,N_4659,N_4666);
nor U5196 (N_5196,N_4897,N_4671);
nand U5197 (N_5197,N_4746,N_4639);
or U5198 (N_5198,N_4912,N_4870);
nor U5199 (N_5199,N_4597,N_4562);
or U5200 (N_5200,N_4636,N_4609);
xnor U5201 (N_5201,N_4958,N_4951);
xor U5202 (N_5202,N_4660,N_4705);
and U5203 (N_5203,N_4795,N_4691);
and U5204 (N_5204,N_4574,N_4946);
nor U5205 (N_5205,N_4600,N_4675);
or U5206 (N_5206,N_4753,N_4518);
or U5207 (N_5207,N_4544,N_4551);
xor U5208 (N_5208,N_4950,N_4737);
nor U5209 (N_5209,N_4538,N_4531);
nand U5210 (N_5210,N_4873,N_4507);
nor U5211 (N_5211,N_4524,N_4641);
xnor U5212 (N_5212,N_4947,N_4813);
nand U5213 (N_5213,N_4996,N_4868);
and U5214 (N_5214,N_4949,N_4680);
xnor U5215 (N_5215,N_4816,N_4943);
nand U5216 (N_5216,N_4758,N_4797);
nand U5217 (N_5217,N_4785,N_4633);
xnor U5218 (N_5218,N_4564,N_4613);
or U5219 (N_5219,N_4896,N_4880);
nand U5220 (N_5220,N_4623,N_4903);
or U5221 (N_5221,N_4982,N_4503);
xnor U5222 (N_5222,N_4930,N_4527);
nand U5223 (N_5223,N_4850,N_4853);
nand U5224 (N_5224,N_4851,N_4834);
nand U5225 (N_5225,N_4709,N_4822);
nand U5226 (N_5226,N_4665,N_4900);
and U5227 (N_5227,N_4837,N_4585);
xor U5228 (N_5228,N_4509,N_4810);
nand U5229 (N_5229,N_4793,N_4877);
nor U5230 (N_5230,N_4541,N_4661);
and U5231 (N_5231,N_4771,N_4909);
xnor U5232 (N_5232,N_4553,N_4591);
nand U5233 (N_5233,N_4734,N_4545);
or U5234 (N_5234,N_4803,N_4905);
or U5235 (N_5235,N_4693,N_4694);
nand U5236 (N_5236,N_4766,N_4695);
and U5237 (N_5237,N_4688,N_4826);
nor U5238 (N_5238,N_4808,N_4792);
xnor U5239 (N_5239,N_4866,N_4720);
and U5240 (N_5240,N_4846,N_4728);
nand U5241 (N_5241,N_4805,N_4634);
nor U5242 (N_5242,N_4904,N_4844);
or U5243 (N_5243,N_4522,N_4995);
xnor U5244 (N_5244,N_4925,N_4935);
nand U5245 (N_5245,N_4886,N_4555);
or U5246 (N_5246,N_4599,N_4651);
xnor U5247 (N_5247,N_4807,N_4532);
nor U5248 (N_5248,N_4546,N_4876);
xnor U5249 (N_5249,N_4918,N_4881);
xor U5250 (N_5250,N_4525,N_4679);
xnor U5251 (N_5251,N_4920,N_4623);
xnor U5252 (N_5252,N_4903,N_4639);
xor U5253 (N_5253,N_4582,N_4819);
nand U5254 (N_5254,N_4581,N_4790);
nor U5255 (N_5255,N_4723,N_4779);
and U5256 (N_5256,N_4532,N_4943);
or U5257 (N_5257,N_4656,N_4569);
nor U5258 (N_5258,N_4692,N_4625);
or U5259 (N_5259,N_4875,N_4834);
nor U5260 (N_5260,N_4936,N_4585);
nor U5261 (N_5261,N_4935,N_4796);
nor U5262 (N_5262,N_4849,N_4593);
and U5263 (N_5263,N_4783,N_4606);
xnor U5264 (N_5264,N_4709,N_4583);
nand U5265 (N_5265,N_4516,N_4591);
or U5266 (N_5266,N_4601,N_4688);
or U5267 (N_5267,N_4900,N_4818);
and U5268 (N_5268,N_4658,N_4765);
or U5269 (N_5269,N_4588,N_4955);
and U5270 (N_5270,N_4934,N_4926);
nor U5271 (N_5271,N_4523,N_4978);
or U5272 (N_5272,N_4786,N_4568);
and U5273 (N_5273,N_4964,N_4754);
nor U5274 (N_5274,N_4505,N_4997);
or U5275 (N_5275,N_4960,N_4700);
nand U5276 (N_5276,N_4756,N_4632);
nand U5277 (N_5277,N_4789,N_4660);
nand U5278 (N_5278,N_4786,N_4659);
xnor U5279 (N_5279,N_4966,N_4728);
and U5280 (N_5280,N_4545,N_4884);
or U5281 (N_5281,N_4548,N_4911);
xor U5282 (N_5282,N_4697,N_4591);
nor U5283 (N_5283,N_4510,N_4968);
or U5284 (N_5284,N_4532,N_4867);
xnor U5285 (N_5285,N_4655,N_4722);
nand U5286 (N_5286,N_4968,N_4973);
and U5287 (N_5287,N_4586,N_4673);
xnor U5288 (N_5288,N_4745,N_4524);
xnor U5289 (N_5289,N_4655,N_4870);
or U5290 (N_5290,N_4917,N_4890);
xnor U5291 (N_5291,N_4876,N_4765);
xnor U5292 (N_5292,N_4779,N_4819);
nand U5293 (N_5293,N_4681,N_4963);
nand U5294 (N_5294,N_4665,N_4782);
xnor U5295 (N_5295,N_4804,N_4788);
nor U5296 (N_5296,N_4914,N_4529);
or U5297 (N_5297,N_4659,N_4684);
nor U5298 (N_5298,N_4701,N_4664);
xor U5299 (N_5299,N_4940,N_4788);
and U5300 (N_5300,N_4507,N_4536);
nand U5301 (N_5301,N_4561,N_4830);
or U5302 (N_5302,N_4758,N_4819);
nor U5303 (N_5303,N_4733,N_4700);
nand U5304 (N_5304,N_4698,N_4863);
or U5305 (N_5305,N_4933,N_4685);
xnor U5306 (N_5306,N_4572,N_4950);
nand U5307 (N_5307,N_4765,N_4696);
nand U5308 (N_5308,N_4698,N_4560);
and U5309 (N_5309,N_4856,N_4514);
nor U5310 (N_5310,N_4604,N_4800);
nor U5311 (N_5311,N_4566,N_4970);
nor U5312 (N_5312,N_4804,N_4847);
nand U5313 (N_5313,N_4646,N_4799);
nor U5314 (N_5314,N_4984,N_4719);
or U5315 (N_5315,N_4584,N_4683);
nand U5316 (N_5316,N_4985,N_4974);
and U5317 (N_5317,N_4921,N_4733);
or U5318 (N_5318,N_4657,N_4789);
nor U5319 (N_5319,N_4908,N_4782);
nor U5320 (N_5320,N_4877,N_4628);
and U5321 (N_5321,N_4759,N_4930);
or U5322 (N_5322,N_4910,N_4992);
or U5323 (N_5323,N_4818,N_4576);
nand U5324 (N_5324,N_4922,N_4581);
and U5325 (N_5325,N_4556,N_4989);
and U5326 (N_5326,N_4905,N_4675);
or U5327 (N_5327,N_4904,N_4946);
and U5328 (N_5328,N_4853,N_4973);
nor U5329 (N_5329,N_4631,N_4853);
xnor U5330 (N_5330,N_4691,N_4792);
or U5331 (N_5331,N_4591,N_4706);
or U5332 (N_5332,N_4660,N_4678);
xor U5333 (N_5333,N_4611,N_4855);
nand U5334 (N_5334,N_4808,N_4733);
nand U5335 (N_5335,N_4810,N_4992);
xnor U5336 (N_5336,N_4587,N_4686);
xor U5337 (N_5337,N_4640,N_4857);
nand U5338 (N_5338,N_4719,N_4915);
and U5339 (N_5339,N_4704,N_4944);
nand U5340 (N_5340,N_4636,N_4913);
nor U5341 (N_5341,N_4883,N_4754);
and U5342 (N_5342,N_4768,N_4870);
xor U5343 (N_5343,N_4571,N_4914);
and U5344 (N_5344,N_4649,N_4886);
nor U5345 (N_5345,N_4516,N_4922);
or U5346 (N_5346,N_4879,N_4828);
nor U5347 (N_5347,N_4782,N_4873);
or U5348 (N_5348,N_4648,N_4813);
or U5349 (N_5349,N_4886,N_4931);
nor U5350 (N_5350,N_4917,N_4574);
xor U5351 (N_5351,N_4551,N_4899);
nand U5352 (N_5352,N_4880,N_4535);
nand U5353 (N_5353,N_4732,N_4743);
or U5354 (N_5354,N_4581,N_4921);
nor U5355 (N_5355,N_4893,N_4934);
nand U5356 (N_5356,N_4887,N_4989);
nor U5357 (N_5357,N_4893,N_4850);
xnor U5358 (N_5358,N_4626,N_4793);
and U5359 (N_5359,N_4940,N_4678);
nand U5360 (N_5360,N_4870,N_4907);
nand U5361 (N_5361,N_4532,N_4705);
xor U5362 (N_5362,N_4769,N_4967);
and U5363 (N_5363,N_4549,N_4588);
nor U5364 (N_5364,N_4599,N_4965);
or U5365 (N_5365,N_4768,N_4831);
xor U5366 (N_5366,N_4775,N_4735);
or U5367 (N_5367,N_4707,N_4928);
nand U5368 (N_5368,N_4848,N_4525);
or U5369 (N_5369,N_4514,N_4946);
and U5370 (N_5370,N_4984,N_4920);
and U5371 (N_5371,N_4594,N_4726);
and U5372 (N_5372,N_4958,N_4673);
nor U5373 (N_5373,N_4875,N_4548);
xnor U5374 (N_5374,N_4858,N_4827);
nor U5375 (N_5375,N_4722,N_4720);
and U5376 (N_5376,N_4701,N_4850);
nor U5377 (N_5377,N_4587,N_4740);
xnor U5378 (N_5378,N_4662,N_4734);
xnor U5379 (N_5379,N_4944,N_4749);
nor U5380 (N_5380,N_4722,N_4595);
and U5381 (N_5381,N_4982,N_4884);
nand U5382 (N_5382,N_4627,N_4825);
and U5383 (N_5383,N_4899,N_4842);
and U5384 (N_5384,N_4813,N_4989);
and U5385 (N_5385,N_4728,N_4957);
xor U5386 (N_5386,N_4902,N_4522);
xnor U5387 (N_5387,N_4504,N_4784);
or U5388 (N_5388,N_4852,N_4855);
or U5389 (N_5389,N_4999,N_4815);
nor U5390 (N_5390,N_4818,N_4697);
or U5391 (N_5391,N_4944,N_4854);
and U5392 (N_5392,N_4974,N_4926);
xor U5393 (N_5393,N_4734,N_4762);
xor U5394 (N_5394,N_4655,N_4973);
nor U5395 (N_5395,N_4720,N_4879);
and U5396 (N_5396,N_4878,N_4867);
nand U5397 (N_5397,N_4894,N_4722);
and U5398 (N_5398,N_4531,N_4789);
or U5399 (N_5399,N_4879,N_4692);
or U5400 (N_5400,N_4767,N_4798);
or U5401 (N_5401,N_4632,N_4925);
nor U5402 (N_5402,N_4871,N_4638);
nor U5403 (N_5403,N_4777,N_4560);
nand U5404 (N_5404,N_4528,N_4803);
nor U5405 (N_5405,N_4806,N_4704);
xnor U5406 (N_5406,N_4622,N_4724);
or U5407 (N_5407,N_4977,N_4963);
or U5408 (N_5408,N_4773,N_4610);
xor U5409 (N_5409,N_4664,N_4718);
and U5410 (N_5410,N_4553,N_4507);
xnor U5411 (N_5411,N_4750,N_4805);
nor U5412 (N_5412,N_4501,N_4793);
xnor U5413 (N_5413,N_4994,N_4862);
nand U5414 (N_5414,N_4645,N_4573);
nand U5415 (N_5415,N_4628,N_4629);
xor U5416 (N_5416,N_4590,N_4504);
or U5417 (N_5417,N_4568,N_4778);
and U5418 (N_5418,N_4503,N_4578);
xnor U5419 (N_5419,N_4519,N_4680);
and U5420 (N_5420,N_4770,N_4762);
nand U5421 (N_5421,N_4842,N_4992);
or U5422 (N_5422,N_4968,N_4869);
and U5423 (N_5423,N_4735,N_4610);
nor U5424 (N_5424,N_4958,N_4897);
xnor U5425 (N_5425,N_4913,N_4559);
nand U5426 (N_5426,N_4550,N_4626);
or U5427 (N_5427,N_4993,N_4777);
and U5428 (N_5428,N_4524,N_4738);
nand U5429 (N_5429,N_4549,N_4672);
nor U5430 (N_5430,N_4520,N_4646);
or U5431 (N_5431,N_4819,N_4905);
nand U5432 (N_5432,N_4701,N_4882);
nand U5433 (N_5433,N_4737,N_4906);
nand U5434 (N_5434,N_4891,N_4847);
nor U5435 (N_5435,N_4678,N_4550);
and U5436 (N_5436,N_4754,N_4645);
nand U5437 (N_5437,N_4849,N_4808);
nand U5438 (N_5438,N_4628,N_4724);
and U5439 (N_5439,N_4516,N_4864);
or U5440 (N_5440,N_4796,N_4648);
nor U5441 (N_5441,N_4844,N_4691);
xor U5442 (N_5442,N_4537,N_4569);
nor U5443 (N_5443,N_4923,N_4611);
xnor U5444 (N_5444,N_4939,N_4884);
nor U5445 (N_5445,N_4946,N_4711);
nor U5446 (N_5446,N_4961,N_4773);
xnor U5447 (N_5447,N_4908,N_4892);
nand U5448 (N_5448,N_4936,N_4503);
nand U5449 (N_5449,N_4604,N_4761);
and U5450 (N_5450,N_4578,N_4502);
nor U5451 (N_5451,N_4747,N_4732);
nor U5452 (N_5452,N_4960,N_4766);
nand U5453 (N_5453,N_4547,N_4743);
nand U5454 (N_5454,N_4843,N_4892);
nand U5455 (N_5455,N_4852,N_4995);
nor U5456 (N_5456,N_4931,N_4988);
nand U5457 (N_5457,N_4675,N_4980);
nor U5458 (N_5458,N_4524,N_4577);
or U5459 (N_5459,N_4735,N_4948);
and U5460 (N_5460,N_4880,N_4537);
and U5461 (N_5461,N_4587,N_4883);
or U5462 (N_5462,N_4653,N_4593);
xor U5463 (N_5463,N_4995,N_4924);
or U5464 (N_5464,N_4964,N_4533);
and U5465 (N_5465,N_4655,N_4651);
or U5466 (N_5466,N_4515,N_4736);
and U5467 (N_5467,N_4998,N_4514);
nand U5468 (N_5468,N_4793,N_4651);
nor U5469 (N_5469,N_4722,N_4564);
or U5470 (N_5470,N_4952,N_4899);
nor U5471 (N_5471,N_4504,N_4898);
xor U5472 (N_5472,N_4951,N_4774);
or U5473 (N_5473,N_4658,N_4567);
or U5474 (N_5474,N_4877,N_4590);
xnor U5475 (N_5475,N_4628,N_4940);
xnor U5476 (N_5476,N_4937,N_4653);
nor U5477 (N_5477,N_4918,N_4726);
nand U5478 (N_5478,N_4919,N_4817);
xnor U5479 (N_5479,N_4999,N_4661);
nand U5480 (N_5480,N_4584,N_4899);
or U5481 (N_5481,N_4932,N_4906);
and U5482 (N_5482,N_4728,N_4832);
nor U5483 (N_5483,N_4806,N_4559);
or U5484 (N_5484,N_4608,N_4771);
nand U5485 (N_5485,N_4567,N_4896);
nand U5486 (N_5486,N_4513,N_4825);
xor U5487 (N_5487,N_4891,N_4600);
nand U5488 (N_5488,N_4895,N_4708);
and U5489 (N_5489,N_4887,N_4833);
and U5490 (N_5490,N_4654,N_4990);
or U5491 (N_5491,N_4961,N_4615);
and U5492 (N_5492,N_4676,N_4957);
nand U5493 (N_5493,N_4750,N_4840);
nand U5494 (N_5494,N_4648,N_4641);
or U5495 (N_5495,N_4747,N_4963);
or U5496 (N_5496,N_4753,N_4733);
and U5497 (N_5497,N_4783,N_4745);
nor U5498 (N_5498,N_4758,N_4614);
or U5499 (N_5499,N_4986,N_4815);
and U5500 (N_5500,N_5262,N_5411);
nand U5501 (N_5501,N_5213,N_5166);
nor U5502 (N_5502,N_5015,N_5410);
xor U5503 (N_5503,N_5081,N_5119);
or U5504 (N_5504,N_5342,N_5293);
or U5505 (N_5505,N_5209,N_5247);
and U5506 (N_5506,N_5196,N_5235);
or U5507 (N_5507,N_5321,N_5215);
xor U5508 (N_5508,N_5490,N_5201);
nand U5509 (N_5509,N_5358,N_5181);
nand U5510 (N_5510,N_5044,N_5036);
xnor U5511 (N_5511,N_5335,N_5354);
and U5512 (N_5512,N_5090,N_5259);
nor U5513 (N_5513,N_5161,N_5296);
or U5514 (N_5514,N_5195,N_5052);
nor U5515 (N_5515,N_5420,N_5272);
nand U5516 (N_5516,N_5186,N_5025);
nor U5517 (N_5517,N_5417,N_5289);
or U5518 (N_5518,N_5388,N_5101);
or U5519 (N_5519,N_5111,N_5476);
and U5520 (N_5520,N_5375,N_5386);
nand U5521 (N_5521,N_5024,N_5487);
nand U5522 (N_5522,N_5395,N_5359);
and U5523 (N_5523,N_5002,N_5422);
or U5524 (N_5524,N_5057,N_5326);
and U5525 (N_5525,N_5205,N_5010);
and U5526 (N_5526,N_5017,N_5404);
nand U5527 (N_5527,N_5441,N_5049);
or U5528 (N_5528,N_5117,N_5221);
or U5529 (N_5529,N_5059,N_5261);
nor U5530 (N_5530,N_5435,N_5290);
nor U5531 (N_5531,N_5430,N_5495);
nor U5532 (N_5532,N_5477,N_5131);
nor U5533 (N_5533,N_5100,N_5268);
or U5534 (N_5534,N_5418,N_5093);
nand U5535 (N_5535,N_5264,N_5120);
nand U5536 (N_5536,N_5297,N_5462);
nand U5537 (N_5537,N_5083,N_5498);
or U5538 (N_5538,N_5373,N_5333);
xor U5539 (N_5539,N_5063,N_5160);
xor U5540 (N_5540,N_5271,N_5366);
xor U5541 (N_5541,N_5048,N_5400);
nand U5542 (N_5542,N_5095,N_5133);
xor U5543 (N_5543,N_5172,N_5338);
xor U5544 (N_5544,N_5184,N_5113);
xnor U5545 (N_5545,N_5029,N_5364);
or U5546 (N_5546,N_5428,N_5141);
nor U5547 (N_5547,N_5469,N_5125);
nor U5548 (N_5548,N_5445,N_5233);
nor U5549 (N_5549,N_5085,N_5301);
xnor U5550 (N_5550,N_5287,N_5202);
xor U5551 (N_5551,N_5176,N_5454);
nand U5552 (N_5552,N_5362,N_5001);
and U5553 (N_5553,N_5391,N_5199);
nor U5554 (N_5554,N_5070,N_5088);
xor U5555 (N_5555,N_5258,N_5414);
xnor U5556 (N_5556,N_5347,N_5171);
or U5557 (N_5557,N_5427,N_5452);
and U5558 (N_5558,N_5304,N_5041);
and U5559 (N_5559,N_5279,N_5046);
nand U5560 (N_5560,N_5352,N_5457);
and U5561 (N_5561,N_5311,N_5345);
and U5562 (N_5562,N_5156,N_5045);
and U5563 (N_5563,N_5327,N_5034);
nand U5564 (N_5564,N_5084,N_5329);
xnor U5565 (N_5565,N_5478,N_5399);
nand U5566 (N_5566,N_5053,N_5191);
nand U5567 (N_5567,N_5456,N_5488);
or U5568 (N_5568,N_5305,N_5320);
xor U5569 (N_5569,N_5365,N_5265);
nor U5570 (N_5570,N_5163,N_5474);
nand U5571 (N_5571,N_5148,N_5109);
nor U5572 (N_5572,N_5402,N_5256);
or U5573 (N_5573,N_5374,N_5357);
and U5574 (N_5574,N_5096,N_5130);
or U5575 (N_5575,N_5413,N_5466);
nor U5576 (N_5576,N_5447,N_5037);
nor U5577 (N_5577,N_5192,N_5419);
nand U5578 (N_5578,N_5206,N_5153);
xor U5579 (N_5579,N_5177,N_5401);
nand U5580 (N_5580,N_5231,N_5112);
and U5581 (N_5581,N_5019,N_5481);
or U5582 (N_5582,N_5239,N_5079);
and U5583 (N_5583,N_5137,N_5162);
and U5584 (N_5584,N_5406,N_5115);
or U5585 (N_5585,N_5307,N_5405);
nand U5586 (N_5586,N_5439,N_5281);
and U5587 (N_5587,N_5018,N_5444);
or U5588 (N_5588,N_5341,N_5194);
nand U5589 (N_5589,N_5464,N_5066);
nor U5590 (N_5590,N_5016,N_5087);
xor U5591 (N_5591,N_5227,N_5328);
xor U5592 (N_5592,N_5183,N_5243);
and U5593 (N_5593,N_5343,N_5050);
or U5594 (N_5594,N_5003,N_5266);
xor U5595 (N_5595,N_5425,N_5108);
nand U5596 (N_5596,N_5121,N_5260);
xnor U5597 (N_5597,N_5122,N_5179);
or U5598 (N_5598,N_5180,N_5159);
xor U5599 (N_5599,N_5127,N_5069);
nand U5600 (N_5600,N_5021,N_5074);
nor U5601 (N_5601,N_5339,N_5222);
nor U5602 (N_5602,N_5241,N_5030);
and U5603 (N_5603,N_5229,N_5434);
nor U5604 (N_5604,N_5203,N_5000);
xnor U5605 (N_5605,N_5197,N_5255);
nor U5606 (N_5606,N_5378,N_5032);
and U5607 (N_5607,N_5223,N_5237);
nand U5608 (N_5608,N_5035,N_5463);
nand U5609 (N_5609,N_5094,N_5234);
nor U5610 (N_5610,N_5154,N_5064);
and U5611 (N_5611,N_5062,N_5453);
and U5612 (N_5612,N_5383,N_5449);
and U5613 (N_5613,N_5368,N_5140);
and U5614 (N_5614,N_5280,N_5249);
nor U5615 (N_5615,N_5139,N_5150);
or U5616 (N_5616,N_5104,N_5496);
xnor U5617 (N_5617,N_5007,N_5220);
xnor U5618 (N_5618,N_5110,N_5322);
nor U5619 (N_5619,N_5011,N_5344);
nor U5620 (N_5620,N_5319,N_5274);
or U5621 (N_5621,N_5284,N_5068);
or U5622 (N_5622,N_5313,N_5144);
nand U5623 (N_5623,N_5306,N_5379);
nor U5624 (N_5624,N_5269,N_5408);
nand U5625 (N_5625,N_5424,N_5291);
nand U5626 (N_5626,N_5372,N_5027);
or U5627 (N_5627,N_5497,N_5086);
or U5628 (N_5628,N_5253,N_5031);
nor U5629 (N_5629,N_5216,N_5361);
nand U5630 (N_5630,N_5055,N_5043);
nor U5631 (N_5631,N_5080,N_5494);
or U5632 (N_5632,N_5299,N_5270);
and U5633 (N_5633,N_5136,N_5302);
xnor U5634 (N_5634,N_5168,N_5423);
nand U5635 (N_5635,N_5242,N_5483);
and U5636 (N_5636,N_5022,N_5263);
xor U5637 (N_5637,N_5039,N_5026);
nor U5638 (N_5638,N_5089,N_5170);
nor U5639 (N_5639,N_5492,N_5240);
and U5640 (N_5640,N_5105,N_5285);
xor U5641 (N_5641,N_5409,N_5218);
nand U5642 (N_5642,N_5288,N_5437);
nand U5643 (N_5643,N_5292,N_5228);
xor U5644 (N_5644,N_5387,N_5325);
xor U5645 (N_5645,N_5047,N_5350);
xnor U5646 (N_5646,N_5470,N_5097);
or U5647 (N_5647,N_5107,N_5219);
or U5648 (N_5648,N_5480,N_5340);
nor U5649 (N_5649,N_5278,N_5232);
nor U5650 (N_5650,N_5076,N_5479);
nor U5651 (N_5651,N_5275,N_5252);
nand U5652 (N_5652,N_5316,N_5167);
nand U5653 (N_5653,N_5389,N_5468);
nor U5654 (N_5654,N_5182,N_5407);
or U5655 (N_5655,N_5248,N_5214);
nand U5656 (N_5656,N_5436,N_5385);
or U5657 (N_5657,N_5426,N_5005);
and U5658 (N_5658,N_5099,N_5072);
and U5659 (N_5659,N_5075,N_5152);
and U5660 (N_5660,N_5224,N_5384);
and U5661 (N_5661,N_5324,N_5295);
nand U5662 (N_5662,N_5028,N_5103);
xnor U5663 (N_5663,N_5416,N_5377);
or U5664 (N_5664,N_5082,N_5450);
or U5665 (N_5665,N_5403,N_5443);
xnor U5666 (N_5666,N_5489,N_5485);
or U5667 (N_5667,N_5225,N_5370);
nand U5668 (N_5668,N_5106,N_5472);
or U5669 (N_5669,N_5286,N_5363);
nor U5670 (N_5670,N_5174,N_5189);
nor U5671 (N_5671,N_5315,N_5238);
nor U5672 (N_5672,N_5008,N_5397);
xor U5673 (N_5673,N_5376,N_5020);
and U5674 (N_5674,N_5294,N_5356);
nand U5675 (N_5675,N_5346,N_5198);
and U5676 (N_5676,N_5337,N_5440);
and U5677 (N_5677,N_5250,N_5467);
nor U5678 (N_5678,N_5254,N_5132);
and U5679 (N_5679,N_5078,N_5398);
nor U5680 (N_5680,N_5267,N_5102);
or U5681 (N_5681,N_5207,N_5392);
or U5682 (N_5682,N_5067,N_5382);
xnor U5683 (N_5683,N_5381,N_5369);
or U5684 (N_5684,N_5204,N_5282);
and U5685 (N_5685,N_5330,N_5458);
or U5686 (N_5686,N_5236,N_5116);
or U5687 (N_5687,N_5190,N_5200);
or U5688 (N_5688,N_5394,N_5465);
and U5689 (N_5689,N_5367,N_5165);
and U5690 (N_5690,N_5226,N_5033);
nand U5691 (N_5691,N_5147,N_5134);
nor U5692 (N_5692,N_5124,N_5118);
nor U5693 (N_5693,N_5128,N_5298);
nand U5694 (N_5694,N_5210,N_5460);
nor U5695 (N_5695,N_5332,N_5091);
nand U5696 (N_5696,N_5331,N_5155);
and U5697 (N_5697,N_5244,N_5175);
and U5698 (N_5698,N_5169,N_5303);
or U5699 (N_5699,N_5421,N_5014);
nand U5700 (N_5700,N_5123,N_5491);
nand U5701 (N_5701,N_5459,N_5114);
nand U5702 (N_5702,N_5396,N_5451);
nor U5703 (N_5703,N_5349,N_5173);
nand U5704 (N_5704,N_5318,N_5390);
and U5705 (N_5705,N_5438,N_5212);
nor U5706 (N_5706,N_5217,N_5208);
xnor U5707 (N_5707,N_5486,N_5146);
and U5708 (N_5708,N_5245,N_5393);
nor U5709 (N_5709,N_5251,N_5273);
xor U5710 (N_5710,N_5211,N_5433);
xor U5711 (N_5711,N_5060,N_5073);
nor U5712 (N_5712,N_5092,N_5126);
nand U5713 (N_5713,N_5071,N_5009);
nor U5714 (N_5714,N_5355,N_5371);
and U5715 (N_5715,N_5360,N_5429);
nor U5716 (N_5716,N_5277,N_5164);
and U5717 (N_5717,N_5006,N_5038);
nand U5718 (N_5718,N_5455,N_5246);
nor U5719 (N_5719,N_5143,N_5415);
or U5720 (N_5720,N_5061,N_5446);
and U5721 (N_5721,N_5051,N_5230);
nor U5722 (N_5722,N_5484,N_5351);
xor U5723 (N_5723,N_5471,N_5151);
nand U5724 (N_5724,N_5135,N_5158);
xnor U5725 (N_5725,N_5193,N_5310);
and U5726 (N_5726,N_5475,N_5187);
xor U5727 (N_5727,N_5129,N_5185);
nor U5728 (N_5728,N_5145,N_5336);
nor U5729 (N_5729,N_5257,N_5323);
nand U5730 (N_5730,N_5334,N_5442);
nor U5731 (N_5731,N_5013,N_5142);
nand U5732 (N_5732,N_5283,N_5380);
and U5733 (N_5733,N_5098,N_5065);
and U5734 (N_5734,N_5461,N_5314);
nand U5735 (N_5735,N_5188,N_5012);
nand U5736 (N_5736,N_5308,N_5040);
nor U5737 (N_5737,N_5448,N_5312);
and U5738 (N_5738,N_5348,N_5077);
and U5739 (N_5739,N_5300,N_5023);
nand U5740 (N_5740,N_5493,N_5054);
nand U5741 (N_5741,N_5276,N_5309);
and U5742 (N_5742,N_5431,N_5149);
nand U5743 (N_5743,N_5499,N_5157);
xnor U5744 (N_5744,N_5473,N_5058);
or U5745 (N_5745,N_5138,N_5412);
nand U5746 (N_5746,N_5056,N_5004);
xor U5747 (N_5747,N_5482,N_5432);
nand U5748 (N_5748,N_5042,N_5353);
nor U5749 (N_5749,N_5317,N_5178);
or U5750 (N_5750,N_5196,N_5444);
nor U5751 (N_5751,N_5472,N_5341);
xor U5752 (N_5752,N_5225,N_5080);
and U5753 (N_5753,N_5380,N_5068);
xor U5754 (N_5754,N_5007,N_5469);
xnor U5755 (N_5755,N_5477,N_5068);
and U5756 (N_5756,N_5083,N_5281);
xnor U5757 (N_5757,N_5434,N_5123);
and U5758 (N_5758,N_5235,N_5140);
xor U5759 (N_5759,N_5027,N_5211);
and U5760 (N_5760,N_5036,N_5390);
xor U5761 (N_5761,N_5158,N_5210);
nand U5762 (N_5762,N_5445,N_5018);
xor U5763 (N_5763,N_5314,N_5449);
xor U5764 (N_5764,N_5320,N_5308);
or U5765 (N_5765,N_5181,N_5279);
nand U5766 (N_5766,N_5345,N_5150);
nand U5767 (N_5767,N_5095,N_5357);
nand U5768 (N_5768,N_5100,N_5235);
nand U5769 (N_5769,N_5050,N_5196);
nor U5770 (N_5770,N_5085,N_5459);
nand U5771 (N_5771,N_5124,N_5402);
and U5772 (N_5772,N_5163,N_5224);
nor U5773 (N_5773,N_5051,N_5459);
xor U5774 (N_5774,N_5237,N_5010);
xnor U5775 (N_5775,N_5428,N_5348);
and U5776 (N_5776,N_5130,N_5157);
and U5777 (N_5777,N_5205,N_5287);
and U5778 (N_5778,N_5465,N_5199);
or U5779 (N_5779,N_5059,N_5262);
or U5780 (N_5780,N_5254,N_5396);
and U5781 (N_5781,N_5066,N_5183);
nor U5782 (N_5782,N_5442,N_5359);
or U5783 (N_5783,N_5327,N_5467);
nor U5784 (N_5784,N_5247,N_5268);
nor U5785 (N_5785,N_5171,N_5196);
and U5786 (N_5786,N_5118,N_5347);
or U5787 (N_5787,N_5197,N_5406);
or U5788 (N_5788,N_5170,N_5491);
xor U5789 (N_5789,N_5105,N_5464);
nand U5790 (N_5790,N_5418,N_5487);
nand U5791 (N_5791,N_5044,N_5037);
or U5792 (N_5792,N_5005,N_5235);
and U5793 (N_5793,N_5046,N_5421);
xnor U5794 (N_5794,N_5313,N_5158);
and U5795 (N_5795,N_5262,N_5235);
nand U5796 (N_5796,N_5231,N_5105);
and U5797 (N_5797,N_5420,N_5449);
xor U5798 (N_5798,N_5020,N_5406);
nor U5799 (N_5799,N_5055,N_5241);
xnor U5800 (N_5800,N_5499,N_5230);
xor U5801 (N_5801,N_5255,N_5305);
or U5802 (N_5802,N_5358,N_5150);
nand U5803 (N_5803,N_5042,N_5014);
and U5804 (N_5804,N_5317,N_5320);
nor U5805 (N_5805,N_5187,N_5143);
or U5806 (N_5806,N_5407,N_5144);
xnor U5807 (N_5807,N_5212,N_5202);
and U5808 (N_5808,N_5174,N_5050);
xor U5809 (N_5809,N_5131,N_5379);
xor U5810 (N_5810,N_5163,N_5406);
and U5811 (N_5811,N_5143,N_5038);
xnor U5812 (N_5812,N_5176,N_5320);
nand U5813 (N_5813,N_5478,N_5475);
nand U5814 (N_5814,N_5353,N_5133);
xnor U5815 (N_5815,N_5186,N_5257);
nand U5816 (N_5816,N_5459,N_5005);
and U5817 (N_5817,N_5463,N_5247);
and U5818 (N_5818,N_5380,N_5274);
or U5819 (N_5819,N_5127,N_5199);
nor U5820 (N_5820,N_5294,N_5026);
xor U5821 (N_5821,N_5078,N_5313);
xnor U5822 (N_5822,N_5392,N_5476);
nand U5823 (N_5823,N_5306,N_5033);
nand U5824 (N_5824,N_5192,N_5140);
nand U5825 (N_5825,N_5383,N_5281);
xor U5826 (N_5826,N_5253,N_5280);
xnor U5827 (N_5827,N_5128,N_5062);
xor U5828 (N_5828,N_5180,N_5103);
or U5829 (N_5829,N_5047,N_5214);
xnor U5830 (N_5830,N_5255,N_5466);
and U5831 (N_5831,N_5499,N_5055);
and U5832 (N_5832,N_5033,N_5338);
and U5833 (N_5833,N_5207,N_5024);
or U5834 (N_5834,N_5396,N_5210);
nor U5835 (N_5835,N_5465,N_5370);
nand U5836 (N_5836,N_5080,N_5023);
xor U5837 (N_5837,N_5023,N_5038);
and U5838 (N_5838,N_5469,N_5466);
xor U5839 (N_5839,N_5426,N_5164);
or U5840 (N_5840,N_5024,N_5026);
or U5841 (N_5841,N_5305,N_5435);
or U5842 (N_5842,N_5181,N_5250);
nor U5843 (N_5843,N_5345,N_5467);
nand U5844 (N_5844,N_5162,N_5348);
xnor U5845 (N_5845,N_5294,N_5087);
or U5846 (N_5846,N_5328,N_5074);
xor U5847 (N_5847,N_5398,N_5304);
or U5848 (N_5848,N_5091,N_5441);
nor U5849 (N_5849,N_5293,N_5303);
nor U5850 (N_5850,N_5275,N_5410);
or U5851 (N_5851,N_5349,N_5291);
xor U5852 (N_5852,N_5208,N_5463);
or U5853 (N_5853,N_5045,N_5220);
nand U5854 (N_5854,N_5392,N_5054);
and U5855 (N_5855,N_5029,N_5146);
and U5856 (N_5856,N_5311,N_5273);
nor U5857 (N_5857,N_5434,N_5300);
and U5858 (N_5858,N_5189,N_5138);
and U5859 (N_5859,N_5175,N_5180);
xor U5860 (N_5860,N_5442,N_5424);
nand U5861 (N_5861,N_5033,N_5086);
or U5862 (N_5862,N_5064,N_5438);
nor U5863 (N_5863,N_5453,N_5414);
and U5864 (N_5864,N_5004,N_5453);
or U5865 (N_5865,N_5349,N_5073);
or U5866 (N_5866,N_5351,N_5333);
nand U5867 (N_5867,N_5172,N_5002);
xnor U5868 (N_5868,N_5127,N_5146);
or U5869 (N_5869,N_5206,N_5202);
or U5870 (N_5870,N_5388,N_5402);
xor U5871 (N_5871,N_5461,N_5266);
xor U5872 (N_5872,N_5241,N_5187);
or U5873 (N_5873,N_5405,N_5302);
or U5874 (N_5874,N_5036,N_5487);
nor U5875 (N_5875,N_5137,N_5448);
nand U5876 (N_5876,N_5476,N_5090);
xnor U5877 (N_5877,N_5158,N_5439);
nor U5878 (N_5878,N_5211,N_5011);
xor U5879 (N_5879,N_5446,N_5257);
or U5880 (N_5880,N_5379,N_5404);
nand U5881 (N_5881,N_5152,N_5228);
or U5882 (N_5882,N_5227,N_5396);
and U5883 (N_5883,N_5040,N_5174);
or U5884 (N_5884,N_5270,N_5463);
or U5885 (N_5885,N_5283,N_5389);
xor U5886 (N_5886,N_5468,N_5117);
and U5887 (N_5887,N_5140,N_5185);
nor U5888 (N_5888,N_5211,N_5381);
nand U5889 (N_5889,N_5070,N_5242);
nand U5890 (N_5890,N_5302,N_5076);
nand U5891 (N_5891,N_5347,N_5357);
nand U5892 (N_5892,N_5066,N_5018);
xor U5893 (N_5893,N_5067,N_5470);
xnor U5894 (N_5894,N_5182,N_5051);
nor U5895 (N_5895,N_5377,N_5280);
and U5896 (N_5896,N_5459,N_5453);
or U5897 (N_5897,N_5277,N_5317);
or U5898 (N_5898,N_5245,N_5063);
and U5899 (N_5899,N_5121,N_5111);
xnor U5900 (N_5900,N_5041,N_5472);
or U5901 (N_5901,N_5368,N_5297);
nor U5902 (N_5902,N_5134,N_5010);
or U5903 (N_5903,N_5480,N_5003);
nor U5904 (N_5904,N_5311,N_5485);
nor U5905 (N_5905,N_5019,N_5479);
xnor U5906 (N_5906,N_5081,N_5438);
and U5907 (N_5907,N_5178,N_5203);
or U5908 (N_5908,N_5406,N_5243);
xor U5909 (N_5909,N_5428,N_5234);
nor U5910 (N_5910,N_5372,N_5192);
or U5911 (N_5911,N_5330,N_5315);
nand U5912 (N_5912,N_5049,N_5488);
and U5913 (N_5913,N_5351,N_5364);
nand U5914 (N_5914,N_5029,N_5410);
xor U5915 (N_5915,N_5186,N_5283);
xnor U5916 (N_5916,N_5211,N_5476);
and U5917 (N_5917,N_5357,N_5493);
nor U5918 (N_5918,N_5489,N_5494);
and U5919 (N_5919,N_5119,N_5406);
nand U5920 (N_5920,N_5098,N_5017);
nand U5921 (N_5921,N_5494,N_5049);
or U5922 (N_5922,N_5218,N_5472);
and U5923 (N_5923,N_5312,N_5286);
or U5924 (N_5924,N_5087,N_5160);
xor U5925 (N_5925,N_5174,N_5148);
xnor U5926 (N_5926,N_5260,N_5072);
or U5927 (N_5927,N_5112,N_5115);
nand U5928 (N_5928,N_5408,N_5186);
or U5929 (N_5929,N_5387,N_5366);
xor U5930 (N_5930,N_5283,N_5282);
nor U5931 (N_5931,N_5056,N_5259);
or U5932 (N_5932,N_5458,N_5126);
nor U5933 (N_5933,N_5341,N_5238);
nand U5934 (N_5934,N_5313,N_5361);
or U5935 (N_5935,N_5491,N_5075);
nand U5936 (N_5936,N_5123,N_5068);
or U5937 (N_5937,N_5399,N_5363);
xnor U5938 (N_5938,N_5073,N_5259);
nand U5939 (N_5939,N_5370,N_5316);
and U5940 (N_5940,N_5151,N_5187);
xnor U5941 (N_5941,N_5484,N_5134);
xnor U5942 (N_5942,N_5028,N_5078);
and U5943 (N_5943,N_5030,N_5285);
nor U5944 (N_5944,N_5170,N_5052);
and U5945 (N_5945,N_5157,N_5173);
or U5946 (N_5946,N_5034,N_5072);
xnor U5947 (N_5947,N_5381,N_5493);
nor U5948 (N_5948,N_5329,N_5185);
xor U5949 (N_5949,N_5470,N_5045);
or U5950 (N_5950,N_5139,N_5321);
nor U5951 (N_5951,N_5281,N_5328);
xnor U5952 (N_5952,N_5474,N_5189);
and U5953 (N_5953,N_5182,N_5472);
and U5954 (N_5954,N_5196,N_5095);
or U5955 (N_5955,N_5256,N_5012);
xnor U5956 (N_5956,N_5315,N_5230);
or U5957 (N_5957,N_5326,N_5146);
nor U5958 (N_5958,N_5277,N_5089);
xnor U5959 (N_5959,N_5243,N_5437);
nor U5960 (N_5960,N_5356,N_5256);
or U5961 (N_5961,N_5174,N_5348);
nor U5962 (N_5962,N_5058,N_5420);
nand U5963 (N_5963,N_5313,N_5151);
xor U5964 (N_5964,N_5267,N_5355);
nand U5965 (N_5965,N_5486,N_5135);
or U5966 (N_5966,N_5357,N_5301);
and U5967 (N_5967,N_5435,N_5445);
nor U5968 (N_5968,N_5449,N_5254);
or U5969 (N_5969,N_5174,N_5001);
nand U5970 (N_5970,N_5168,N_5183);
or U5971 (N_5971,N_5420,N_5268);
or U5972 (N_5972,N_5208,N_5404);
or U5973 (N_5973,N_5129,N_5463);
and U5974 (N_5974,N_5342,N_5093);
nor U5975 (N_5975,N_5124,N_5441);
xor U5976 (N_5976,N_5094,N_5316);
nand U5977 (N_5977,N_5048,N_5288);
xor U5978 (N_5978,N_5140,N_5226);
xor U5979 (N_5979,N_5336,N_5455);
or U5980 (N_5980,N_5022,N_5314);
xnor U5981 (N_5981,N_5328,N_5365);
nor U5982 (N_5982,N_5317,N_5130);
xnor U5983 (N_5983,N_5224,N_5084);
nand U5984 (N_5984,N_5234,N_5114);
and U5985 (N_5985,N_5075,N_5267);
nand U5986 (N_5986,N_5089,N_5356);
nand U5987 (N_5987,N_5401,N_5065);
xor U5988 (N_5988,N_5408,N_5120);
nor U5989 (N_5989,N_5253,N_5402);
nand U5990 (N_5990,N_5453,N_5404);
xor U5991 (N_5991,N_5336,N_5202);
and U5992 (N_5992,N_5189,N_5376);
xnor U5993 (N_5993,N_5239,N_5163);
nand U5994 (N_5994,N_5499,N_5069);
or U5995 (N_5995,N_5226,N_5343);
nand U5996 (N_5996,N_5004,N_5154);
or U5997 (N_5997,N_5065,N_5042);
and U5998 (N_5998,N_5165,N_5041);
nor U5999 (N_5999,N_5073,N_5174);
and U6000 (N_6000,N_5854,N_5735);
and U6001 (N_6001,N_5538,N_5624);
nor U6002 (N_6002,N_5699,N_5981);
nor U6003 (N_6003,N_5669,N_5713);
xor U6004 (N_6004,N_5800,N_5761);
xor U6005 (N_6005,N_5519,N_5500);
nor U6006 (N_6006,N_5998,N_5868);
and U6007 (N_6007,N_5781,N_5550);
xor U6008 (N_6008,N_5652,N_5999);
nand U6009 (N_6009,N_5689,N_5967);
or U6010 (N_6010,N_5590,N_5930);
and U6011 (N_6011,N_5929,N_5912);
or U6012 (N_6012,N_5531,N_5984);
xor U6013 (N_6013,N_5804,N_5522);
xor U6014 (N_6014,N_5567,N_5941);
xor U6015 (N_6015,N_5973,N_5805);
nor U6016 (N_6016,N_5958,N_5839);
or U6017 (N_6017,N_5851,N_5797);
nor U6018 (N_6018,N_5926,N_5748);
and U6019 (N_6019,N_5970,N_5589);
or U6020 (N_6020,N_5777,N_5892);
nor U6021 (N_6021,N_5622,N_5584);
xor U6022 (N_6022,N_5977,N_5582);
and U6023 (N_6023,N_5558,N_5943);
and U6024 (N_6024,N_5983,N_5738);
or U6025 (N_6025,N_5524,N_5721);
nand U6026 (N_6026,N_5974,N_5563);
or U6027 (N_6027,N_5936,N_5593);
xnor U6028 (N_6028,N_5730,N_5850);
or U6029 (N_6029,N_5802,N_5686);
and U6030 (N_6030,N_5661,N_5893);
nor U6031 (N_6031,N_5934,N_5980);
and U6032 (N_6032,N_5752,N_5557);
xnor U6033 (N_6033,N_5782,N_5501);
nor U6034 (N_6034,N_5874,N_5681);
xnor U6035 (N_6035,N_5731,N_5931);
nand U6036 (N_6036,N_5578,N_5732);
or U6037 (N_6037,N_5809,N_5822);
nor U6038 (N_6038,N_5801,N_5823);
nor U6039 (N_6039,N_5751,N_5609);
xor U6040 (N_6040,N_5543,N_5827);
nor U6041 (N_6041,N_5895,N_5862);
xnor U6042 (N_6042,N_5636,N_5789);
nand U6043 (N_6043,N_5896,N_5647);
or U6044 (N_6044,N_5964,N_5716);
nand U6045 (N_6045,N_5966,N_5860);
nor U6046 (N_6046,N_5544,N_5599);
nand U6047 (N_6047,N_5553,N_5588);
or U6048 (N_6048,N_5598,N_5665);
or U6049 (N_6049,N_5712,N_5743);
nand U6050 (N_6050,N_5855,N_5794);
xnor U6051 (N_6051,N_5734,N_5549);
or U6052 (N_6052,N_5595,N_5872);
and U6053 (N_6053,N_5662,N_5910);
nor U6054 (N_6054,N_5791,N_5900);
xor U6055 (N_6055,N_5675,N_5744);
xnor U6056 (N_6056,N_5869,N_5724);
and U6057 (N_6057,N_5736,N_5775);
or U6058 (N_6058,N_5506,N_5733);
and U6059 (N_6059,N_5603,N_5754);
or U6060 (N_6060,N_5905,N_5678);
nand U6061 (N_6061,N_5503,N_5663);
or U6062 (N_6062,N_5608,N_5798);
or U6063 (N_6063,N_5556,N_5659);
or U6064 (N_6064,N_5753,N_5693);
nand U6065 (N_6065,N_5774,N_5705);
xnor U6066 (N_6066,N_5568,N_5921);
and U6067 (N_6067,N_5684,N_5762);
or U6068 (N_6068,N_5671,N_5803);
xnor U6069 (N_6069,N_5740,N_5903);
and U6070 (N_6070,N_5668,N_5745);
or U6071 (N_6071,N_5529,N_5637);
nand U6072 (N_6072,N_5674,N_5810);
and U6073 (N_6073,N_5517,N_5985);
or U6074 (N_6074,N_5513,N_5554);
xnor U6075 (N_6075,N_5703,N_5946);
nand U6076 (N_6076,N_5757,N_5894);
nand U6077 (N_6077,N_5766,N_5989);
and U6078 (N_6078,N_5932,N_5516);
xor U6079 (N_6079,N_5913,N_5954);
and U6080 (N_6080,N_5790,N_5945);
and U6081 (N_6081,N_5642,N_5651);
nand U6082 (N_6082,N_5807,N_5683);
xor U6083 (N_6083,N_5539,N_5961);
or U6084 (N_6084,N_5886,N_5555);
and U6085 (N_6085,N_5650,N_5701);
nand U6086 (N_6086,N_5623,N_5887);
xnor U6087 (N_6087,N_5843,N_5914);
and U6088 (N_6088,N_5715,N_5867);
or U6089 (N_6089,N_5725,N_5580);
xnor U6090 (N_6090,N_5570,N_5658);
nand U6091 (N_6091,N_5645,N_5955);
xor U6092 (N_6092,N_5680,N_5648);
nor U6093 (N_6093,N_5849,N_5585);
xor U6094 (N_6094,N_5847,N_5879);
or U6095 (N_6095,N_5817,N_5948);
or U6096 (N_6096,N_5676,N_5882);
xor U6097 (N_6097,N_5793,N_5950);
xnor U6098 (N_6098,N_5631,N_5508);
and U6099 (N_6099,N_5911,N_5546);
nand U6100 (N_6100,N_5877,N_5820);
and U6101 (N_6101,N_5937,N_5942);
xor U6102 (N_6102,N_5884,N_5861);
or U6103 (N_6103,N_5602,N_5617);
or U6104 (N_6104,N_5548,N_5646);
xor U6105 (N_6105,N_5933,N_5959);
and U6106 (N_6106,N_5677,N_5763);
xnor U6107 (N_6107,N_5523,N_5512);
and U6108 (N_6108,N_5864,N_5635);
nand U6109 (N_6109,N_5845,N_5878);
and U6110 (N_6110,N_5880,N_5504);
and U6111 (N_6111,N_5962,N_5526);
nor U6112 (N_6112,N_5530,N_5644);
or U6113 (N_6113,N_5653,N_5951);
and U6114 (N_6114,N_5547,N_5904);
xor U6115 (N_6115,N_5828,N_5729);
nor U6116 (N_6116,N_5708,N_5856);
xor U6117 (N_6117,N_5525,N_5520);
nand U6118 (N_6118,N_5627,N_5566);
nand U6119 (N_6119,N_5924,N_5840);
or U6120 (N_6120,N_5632,N_5865);
xor U6121 (N_6121,N_5891,N_5577);
and U6122 (N_6122,N_5965,N_5618);
nand U6123 (N_6123,N_5605,N_5808);
or U6124 (N_6124,N_5755,N_5818);
nor U6125 (N_6125,N_5906,N_5717);
nor U6126 (N_6126,N_5837,N_5611);
nand U6127 (N_6127,N_5770,N_5572);
or U6128 (N_6128,N_5772,N_5586);
nor U6129 (N_6129,N_5614,N_5919);
and U6130 (N_6130,N_5502,N_5515);
nor U6131 (N_6131,N_5534,N_5667);
xnor U6132 (N_6132,N_5816,N_5690);
xnor U6133 (N_6133,N_5838,N_5995);
xnor U6134 (N_6134,N_5704,N_5971);
nand U6135 (N_6135,N_5537,N_5511);
and U6136 (N_6136,N_5994,N_5835);
and U6137 (N_6137,N_5698,N_5747);
xnor U6138 (N_6138,N_5830,N_5792);
nor U6139 (N_6139,N_5842,N_5706);
and U6140 (N_6140,N_5888,N_5982);
nor U6141 (N_6141,N_5996,N_5988);
xnor U6142 (N_6142,N_5746,N_5758);
nor U6143 (N_6143,N_5533,N_5779);
nand U6144 (N_6144,N_5821,N_5923);
xnor U6145 (N_6145,N_5815,N_5814);
or U6146 (N_6146,N_5682,N_5969);
and U6147 (N_6147,N_5521,N_5574);
xor U6148 (N_6148,N_5741,N_5949);
and U6149 (N_6149,N_5944,N_5938);
and U6150 (N_6150,N_5700,N_5709);
nand U6151 (N_6151,N_5960,N_5569);
or U6152 (N_6152,N_5812,N_5990);
nand U6153 (N_6153,N_5863,N_5633);
and U6154 (N_6154,N_5691,N_5890);
xnor U6155 (N_6155,N_5979,N_5728);
nand U6156 (N_6156,N_5655,N_5552);
xor U6157 (N_6157,N_5848,N_5707);
xnor U6158 (N_6158,N_5952,N_5873);
or U6159 (N_6159,N_5889,N_5718);
nand U6160 (N_6160,N_5976,N_5768);
or U6161 (N_6161,N_5902,N_5875);
nor U6162 (N_6162,N_5612,N_5759);
nor U6163 (N_6163,N_5784,N_5920);
or U6164 (N_6164,N_5630,N_5714);
and U6165 (N_6165,N_5615,N_5947);
and U6166 (N_6166,N_5688,N_5831);
and U6167 (N_6167,N_5829,N_5592);
xor U6168 (N_6168,N_5819,N_5532);
nor U6169 (N_6169,N_5601,N_5799);
and U6170 (N_6170,N_5634,N_5695);
nand U6171 (N_6171,N_5510,N_5901);
and U6172 (N_6172,N_5899,N_5720);
nand U6173 (N_6173,N_5997,N_5987);
and U6174 (N_6174,N_5579,N_5885);
nand U6175 (N_6175,N_5771,N_5639);
nor U6176 (N_6176,N_5992,N_5576);
or U6177 (N_6177,N_5916,N_5927);
nor U6178 (N_6178,N_5654,N_5514);
xnor U6179 (N_6179,N_5583,N_5649);
xnor U6180 (N_6180,N_5666,N_5737);
nor U6181 (N_6181,N_5581,N_5600);
and U6182 (N_6182,N_5641,N_5968);
or U6183 (N_6183,N_5859,N_5536);
and U6184 (N_6184,N_5858,N_5697);
xnor U6185 (N_6185,N_5626,N_5594);
nand U6186 (N_6186,N_5972,N_5638);
nand U6187 (N_6187,N_5841,N_5767);
and U6188 (N_6188,N_5540,N_5940);
and U6189 (N_6189,N_5897,N_5773);
xor U6190 (N_6190,N_5750,N_5852);
nor U6191 (N_6191,N_5551,N_5760);
nor U6192 (N_6192,N_5723,N_5857);
xnor U6193 (N_6193,N_5727,N_5694);
or U6194 (N_6194,N_5765,N_5620);
xnor U6195 (N_6195,N_5573,N_5660);
nand U6196 (N_6196,N_5535,N_5957);
xnor U6197 (N_6197,N_5991,N_5670);
or U6198 (N_6198,N_5883,N_5559);
nor U6199 (N_6199,N_5813,N_5832);
or U6200 (N_6200,N_5918,N_5625);
xor U6201 (N_6201,N_5778,N_5953);
nor U6202 (N_6202,N_5518,N_5505);
or U6203 (N_6203,N_5898,N_5780);
xnor U6204 (N_6204,N_5788,N_5978);
and U6205 (N_6205,N_5591,N_5795);
nand U6206 (N_6206,N_5769,N_5825);
xnor U6207 (N_6207,N_5610,N_5606);
nand U6208 (N_6208,N_5710,N_5664);
or U6209 (N_6209,N_5975,N_5672);
and U6210 (N_6210,N_5836,N_5542);
xor U6211 (N_6211,N_5607,N_5613);
nor U6212 (N_6212,N_5719,N_5696);
xor U6213 (N_6213,N_5564,N_5939);
or U6214 (N_6214,N_5679,N_5756);
or U6215 (N_6215,N_5871,N_5673);
and U6216 (N_6216,N_5742,N_5925);
nand U6217 (N_6217,N_5783,N_5587);
and U6218 (N_6218,N_5796,N_5749);
xor U6219 (N_6219,N_5776,N_5619);
nand U6220 (N_6220,N_5687,N_5956);
and U6221 (N_6221,N_5509,N_5565);
or U6222 (N_6222,N_5571,N_5908);
and U6223 (N_6223,N_5657,N_5824);
xnor U6224 (N_6224,N_5575,N_5811);
or U6225 (N_6225,N_5621,N_5907);
or U6226 (N_6226,N_5785,N_5935);
nand U6227 (N_6227,N_5876,N_5870);
nand U6228 (N_6228,N_5881,N_5764);
or U6229 (N_6229,N_5643,N_5993);
or U6230 (N_6230,N_5833,N_5561);
nand U6231 (N_6231,N_5853,N_5826);
xnor U6232 (N_6232,N_5986,N_5541);
and U6233 (N_6233,N_5702,N_5560);
or U6234 (N_6234,N_5806,N_5656);
nand U6235 (N_6235,N_5739,N_5545);
nor U6236 (N_6236,N_5616,N_5928);
xnor U6237 (N_6237,N_5866,N_5640);
xnor U6238 (N_6238,N_5628,N_5629);
xor U6239 (N_6239,N_5909,N_5787);
and U6240 (N_6240,N_5604,N_5846);
or U6241 (N_6241,N_5722,N_5685);
xor U6242 (N_6242,N_5726,N_5692);
nand U6243 (N_6243,N_5786,N_5596);
or U6244 (N_6244,N_5711,N_5917);
nand U6245 (N_6245,N_5834,N_5922);
nand U6246 (N_6246,N_5562,N_5963);
xor U6247 (N_6247,N_5507,N_5527);
nand U6248 (N_6248,N_5597,N_5915);
and U6249 (N_6249,N_5844,N_5528);
and U6250 (N_6250,N_5959,N_5976);
nand U6251 (N_6251,N_5525,N_5557);
xnor U6252 (N_6252,N_5568,N_5896);
or U6253 (N_6253,N_5996,N_5846);
and U6254 (N_6254,N_5723,N_5962);
nor U6255 (N_6255,N_5672,N_5874);
or U6256 (N_6256,N_5784,N_5862);
nor U6257 (N_6257,N_5717,N_5540);
nor U6258 (N_6258,N_5577,N_5640);
and U6259 (N_6259,N_5977,N_5957);
nor U6260 (N_6260,N_5619,N_5789);
xnor U6261 (N_6261,N_5933,N_5765);
nor U6262 (N_6262,N_5950,N_5742);
nand U6263 (N_6263,N_5641,N_5787);
xnor U6264 (N_6264,N_5508,N_5665);
and U6265 (N_6265,N_5647,N_5545);
nor U6266 (N_6266,N_5599,N_5956);
xnor U6267 (N_6267,N_5709,N_5891);
nand U6268 (N_6268,N_5506,N_5936);
or U6269 (N_6269,N_5896,N_5984);
xor U6270 (N_6270,N_5718,N_5516);
nand U6271 (N_6271,N_5872,N_5949);
and U6272 (N_6272,N_5674,N_5587);
or U6273 (N_6273,N_5974,N_5773);
nand U6274 (N_6274,N_5926,N_5834);
and U6275 (N_6275,N_5669,N_5831);
or U6276 (N_6276,N_5881,N_5510);
nand U6277 (N_6277,N_5971,N_5840);
nor U6278 (N_6278,N_5687,N_5937);
xor U6279 (N_6279,N_5678,N_5698);
and U6280 (N_6280,N_5550,N_5933);
nor U6281 (N_6281,N_5512,N_5973);
and U6282 (N_6282,N_5966,N_5974);
and U6283 (N_6283,N_5623,N_5558);
and U6284 (N_6284,N_5724,N_5790);
xnor U6285 (N_6285,N_5646,N_5963);
xnor U6286 (N_6286,N_5545,N_5663);
or U6287 (N_6287,N_5865,N_5945);
and U6288 (N_6288,N_5657,N_5883);
nor U6289 (N_6289,N_5534,N_5928);
nand U6290 (N_6290,N_5635,N_5986);
nor U6291 (N_6291,N_5799,N_5997);
nand U6292 (N_6292,N_5729,N_5753);
and U6293 (N_6293,N_5529,N_5595);
nand U6294 (N_6294,N_5795,N_5571);
and U6295 (N_6295,N_5788,N_5837);
or U6296 (N_6296,N_5650,N_5680);
and U6297 (N_6297,N_5572,N_5851);
or U6298 (N_6298,N_5922,N_5896);
nor U6299 (N_6299,N_5952,N_5687);
and U6300 (N_6300,N_5639,N_5765);
and U6301 (N_6301,N_5817,N_5621);
nor U6302 (N_6302,N_5801,N_5809);
nor U6303 (N_6303,N_5747,N_5608);
xor U6304 (N_6304,N_5886,N_5740);
nand U6305 (N_6305,N_5990,N_5820);
nor U6306 (N_6306,N_5822,N_5980);
nor U6307 (N_6307,N_5528,N_5811);
nor U6308 (N_6308,N_5630,N_5862);
xor U6309 (N_6309,N_5813,N_5546);
or U6310 (N_6310,N_5700,N_5887);
nand U6311 (N_6311,N_5998,N_5932);
nand U6312 (N_6312,N_5892,N_5904);
nand U6313 (N_6313,N_5834,N_5679);
or U6314 (N_6314,N_5693,N_5634);
xor U6315 (N_6315,N_5880,N_5683);
and U6316 (N_6316,N_5597,N_5786);
nand U6317 (N_6317,N_5885,N_5724);
nand U6318 (N_6318,N_5923,N_5699);
nand U6319 (N_6319,N_5780,N_5987);
nor U6320 (N_6320,N_5869,N_5614);
nor U6321 (N_6321,N_5660,N_5588);
and U6322 (N_6322,N_5861,N_5556);
nand U6323 (N_6323,N_5898,N_5560);
nor U6324 (N_6324,N_5790,N_5726);
nand U6325 (N_6325,N_5670,N_5514);
and U6326 (N_6326,N_5772,N_5680);
and U6327 (N_6327,N_5637,N_5798);
nand U6328 (N_6328,N_5760,N_5997);
and U6329 (N_6329,N_5847,N_5728);
nor U6330 (N_6330,N_5820,N_5871);
nand U6331 (N_6331,N_5777,N_5801);
and U6332 (N_6332,N_5559,N_5981);
nand U6333 (N_6333,N_5790,N_5752);
or U6334 (N_6334,N_5642,N_5578);
and U6335 (N_6335,N_5994,N_5848);
xnor U6336 (N_6336,N_5517,N_5566);
and U6337 (N_6337,N_5843,N_5591);
and U6338 (N_6338,N_5897,N_5848);
xnor U6339 (N_6339,N_5677,N_5790);
xor U6340 (N_6340,N_5550,N_5779);
nor U6341 (N_6341,N_5599,N_5864);
or U6342 (N_6342,N_5521,N_5693);
nor U6343 (N_6343,N_5999,N_5549);
xnor U6344 (N_6344,N_5567,N_5834);
xnor U6345 (N_6345,N_5652,N_5959);
nand U6346 (N_6346,N_5898,N_5667);
and U6347 (N_6347,N_5594,N_5611);
nand U6348 (N_6348,N_5877,N_5737);
nor U6349 (N_6349,N_5722,N_5507);
xnor U6350 (N_6350,N_5792,N_5723);
nand U6351 (N_6351,N_5594,N_5834);
nor U6352 (N_6352,N_5771,N_5942);
and U6353 (N_6353,N_5547,N_5566);
and U6354 (N_6354,N_5657,N_5583);
nand U6355 (N_6355,N_5940,N_5812);
xnor U6356 (N_6356,N_5710,N_5561);
or U6357 (N_6357,N_5862,N_5621);
xor U6358 (N_6358,N_5785,N_5605);
xnor U6359 (N_6359,N_5622,N_5686);
or U6360 (N_6360,N_5553,N_5634);
and U6361 (N_6361,N_5956,N_5773);
or U6362 (N_6362,N_5574,N_5814);
nand U6363 (N_6363,N_5939,N_5843);
xor U6364 (N_6364,N_5658,N_5655);
nand U6365 (N_6365,N_5702,N_5553);
or U6366 (N_6366,N_5529,N_5982);
or U6367 (N_6367,N_5580,N_5832);
or U6368 (N_6368,N_5884,N_5538);
and U6369 (N_6369,N_5851,N_5546);
or U6370 (N_6370,N_5953,N_5906);
xnor U6371 (N_6371,N_5919,N_5822);
nor U6372 (N_6372,N_5835,N_5927);
nand U6373 (N_6373,N_5969,N_5748);
nand U6374 (N_6374,N_5533,N_5689);
nor U6375 (N_6375,N_5649,N_5814);
nand U6376 (N_6376,N_5684,N_5528);
and U6377 (N_6377,N_5980,N_5530);
nor U6378 (N_6378,N_5611,N_5596);
nand U6379 (N_6379,N_5870,N_5788);
nor U6380 (N_6380,N_5823,N_5539);
xor U6381 (N_6381,N_5724,N_5895);
and U6382 (N_6382,N_5813,N_5721);
nor U6383 (N_6383,N_5731,N_5558);
nand U6384 (N_6384,N_5516,N_5571);
or U6385 (N_6385,N_5783,N_5798);
and U6386 (N_6386,N_5536,N_5877);
nand U6387 (N_6387,N_5564,N_5652);
nand U6388 (N_6388,N_5706,N_5570);
and U6389 (N_6389,N_5511,N_5876);
or U6390 (N_6390,N_5609,N_5920);
and U6391 (N_6391,N_5557,N_5675);
or U6392 (N_6392,N_5652,N_5907);
nand U6393 (N_6393,N_5514,N_5548);
nand U6394 (N_6394,N_5565,N_5917);
or U6395 (N_6395,N_5840,N_5948);
and U6396 (N_6396,N_5640,N_5513);
nor U6397 (N_6397,N_5576,N_5981);
or U6398 (N_6398,N_5950,N_5882);
xnor U6399 (N_6399,N_5826,N_5938);
nor U6400 (N_6400,N_5850,N_5681);
xor U6401 (N_6401,N_5870,N_5738);
xnor U6402 (N_6402,N_5987,N_5689);
nor U6403 (N_6403,N_5893,N_5698);
nor U6404 (N_6404,N_5933,N_5521);
xnor U6405 (N_6405,N_5754,N_5838);
nand U6406 (N_6406,N_5640,N_5748);
nand U6407 (N_6407,N_5793,N_5738);
nand U6408 (N_6408,N_5888,N_5666);
nand U6409 (N_6409,N_5554,N_5787);
or U6410 (N_6410,N_5683,N_5555);
xnor U6411 (N_6411,N_5699,N_5942);
or U6412 (N_6412,N_5938,N_5720);
nand U6413 (N_6413,N_5933,N_5911);
nand U6414 (N_6414,N_5633,N_5995);
or U6415 (N_6415,N_5790,N_5901);
and U6416 (N_6416,N_5599,N_5926);
or U6417 (N_6417,N_5977,N_5929);
xnor U6418 (N_6418,N_5801,N_5869);
and U6419 (N_6419,N_5796,N_5983);
and U6420 (N_6420,N_5777,N_5797);
xnor U6421 (N_6421,N_5708,N_5841);
nand U6422 (N_6422,N_5504,N_5959);
and U6423 (N_6423,N_5702,N_5930);
or U6424 (N_6424,N_5511,N_5530);
and U6425 (N_6425,N_5870,N_5609);
xor U6426 (N_6426,N_5795,N_5615);
and U6427 (N_6427,N_5701,N_5748);
or U6428 (N_6428,N_5997,N_5657);
nor U6429 (N_6429,N_5724,N_5754);
and U6430 (N_6430,N_5842,N_5653);
or U6431 (N_6431,N_5822,N_5724);
xor U6432 (N_6432,N_5610,N_5979);
nand U6433 (N_6433,N_5794,N_5824);
xor U6434 (N_6434,N_5793,N_5736);
nand U6435 (N_6435,N_5708,N_5857);
or U6436 (N_6436,N_5553,N_5925);
or U6437 (N_6437,N_5946,N_5592);
and U6438 (N_6438,N_5608,N_5527);
nor U6439 (N_6439,N_5759,N_5887);
and U6440 (N_6440,N_5564,N_5627);
or U6441 (N_6441,N_5569,N_5718);
xnor U6442 (N_6442,N_5952,N_5921);
nor U6443 (N_6443,N_5807,N_5920);
or U6444 (N_6444,N_5936,N_5829);
or U6445 (N_6445,N_5761,N_5801);
nand U6446 (N_6446,N_5854,N_5889);
xnor U6447 (N_6447,N_5705,N_5673);
xnor U6448 (N_6448,N_5622,N_5762);
or U6449 (N_6449,N_5596,N_5549);
and U6450 (N_6450,N_5661,N_5656);
and U6451 (N_6451,N_5597,N_5510);
nand U6452 (N_6452,N_5880,N_5841);
xnor U6453 (N_6453,N_5775,N_5579);
nor U6454 (N_6454,N_5968,N_5680);
nor U6455 (N_6455,N_5638,N_5914);
nor U6456 (N_6456,N_5968,N_5502);
nor U6457 (N_6457,N_5521,N_5747);
or U6458 (N_6458,N_5954,N_5869);
nor U6459 (N_6459,N_5699,N_5902);
xnor U6460 (N_6460,N_5512,N_5783);
xnor U6461 (N_6461,N_5717,N_5898);
nand U6462 (N_6462,N_5742,N_5999);
and U6463 (N_6463,N_5834,N_5589);
nand U6464 (N_6464,N_5794,N_5726);
nand U6465 (N_6465,N_5578,N_5766);
or U6466 (N_6466,N_5908,N_5528);
xnor U6467 (N_6467,N_5542,N_5937);
nand U6468 (N_6468,N_5984,N_5559);
xor U6469 (N_6469,N_5577,N_5931);
and U6470 (N_6470,N_5565,N_5860);
xor U6471 (N_6471,N_5665,N_5733);
xor U6472 (N_6472,N_5500,N_5998);
xnor U6473 (N_6473,N_5980,N_5622);
nand U6474 (N_6474,N_5870,N_5676);
nand U6475 (N_6475,N_5868,N_5684);
and U6476 (N_6476,N_5818,N_5515);
nor U6477 (N_6477,N_5700,N_5782);
or U6478 (N_6478,N_5702,N_5693);
nand U6479 (N_6479,N_5974,N_5628);
nor U6480 (N_6480,N_5565,N_5780);
nor U6481 (N_6481,N_5889,N_5728);
xor U6482 (N_6482,N_5655,N_5652);
or U6483 (N_6483,N_5607,N_5715);
nand U6484 (N_6484,N_5689,N_5995);
or U6485 (N_6485,N_5972,N_5889);
xnor U6486 (N_6486,N_5956,N_5833);
or U6487 (N_6487,N_5505,N_5988);
nor U6488 (N_6488,N_5664,N_5975);
xor U6489 (N_6489,N_5536,N_5538);
nor U6490 (N_6490,N_5971,N_5858);
or U6491 (N_6491,N_5677,N_5741);
or U6492 (N_6492,N_5804,N_5703);
xnor U6493 (N_6493,N_5754,N_5699);
and U6494 (N_6494,N_5524,N_5936);
or U6495 (N_6495,N_5595,N_5955);
xnor U6496 (N_6496,N_5792,N_5714);
or U6497 (N_6497,N_5878,N_5501);
and U6498 (N_6498,N_5781,N_5690);
and U6499 (N_6499,N_5878,N_5994);
xor U6500 (N_6500,N_6070,N_6410);
nand U6501 (N_6501,N_6148,N_6437);
and U6502 (N_6502,N_6245,N_6223);
nand U6503 (N_6503,N_6386,N_6198);
and U6504 (N_6504,N_6045,N_6336);
nand U6505 (N_6505,N_6105,N_6483);
nand U6506 (N_6506,N_6216,N_6319);
xnor U6507 (N_6507,N_6081,N_6389);
or U6508 (N_6508,N_6068,N_6329);
nor U6509 (N_6509,N_6150,N_6311);
or U6510 (N_6510,N_6283,N_6233);
nor U6511 (N_6511,N_6133,N_6219);
and U6512 (N_6512,N_6063,N_6276);
nor U6513 (N_6513,N_6476,N_6005);
nand U6514 (N_6514,N_6432,N_6142);
xor U6515 (N_6515,N_6310,N_6126);
xnor U6516 (N_6516,N_6286,N_6317);
nor U6517 (N_6517,N_6295,N_6071);
and U6518 (N_6518,N_6449,N_6156);
and U6519 (N_6519,N_6033,N_6113);
or U6520 (N_6520,N_6431,N_6281);
xnor U6521 (N_6521,N_6407,N_6043);
nor U6522 (N_6522,N_6166,N_6062);
nor U6523 (N_6523,N_6109,N_6265);
nand U6524 (N_6524,N_6461,N_6470);
nand U6525 (N_6525,N_6159,N_6173);
nor U6526 (N_6526,N_6328,N_6091);
xor U6527 (N_6527,N_6376,N_6122);
xnor U6528 (N_6528,N_6208,N_6134);
nand U6529 (N_6529,N_6029,N_6364);
or U6530 (N_6530,N_6469,N_6051);
nand U6531 (N_6531,N_6222,N_6406);
xor U6532 (N_6532,N_6423,N_6330);
or U6533 (N_6533,N_6428,N_6412);
or U6534 (N_6534,N_6128,N_6498);
nand U6535 (N_6535,N_6098,N_6413);
nand U6536 (N_6536,N_6041,N_6006);
nor U6537 (N_6537,N_6155,N_6486);
or U6538 (N_6538,N_6352,N_6044);
nor U6539 (N_6539,N_6050,N_6415);
and U6540 (N_6540,N_6305,N_6104);
xor U6541 (N_6541,N_6239,N_6308);
or U6542 (N_6542,N_6366,N_6210);
nor U6543 (N_6543,N_6185,N_6206);
xnor U6544 (N_6544,N_6491,N_6324);
or U6545 (N_6545,N_6261,N_6209);
and U6546 (N_6546,N_6380,N_6236);
or U6547 (N_6547,N_6184,N_6411);
xor U6548 (N_6548,N_6007,N_6163);
nand U6549 (N_6549,N_6250,N_6038);
nand U6550 (N_6550,N_6061,N_6300);
or U6551 (N_6551,N_6379,N_6054);
nand U6552 (N_6552,N_6264,N_6144);
nor U6553 (N_6553,N_6076,N_6172);
nand U6554 (N_6554,N_6247,N_6046);
nor U6555 (N_6555,N_6338,N_6138);
and U6556 (N_6556,N_6333,N_6040);
and U6557 (N_6557,N_6067,N_6053);
and U6558 (N_6558,N_6152,N_6164);
xor U6559 (N_6559,N_6463,N_6139);
nand U6560 (N_6560,N_6465,N_6271);
nand U6561 (N_6561,N_6189,N_6137);
nor U6562 (N_6562,N_6493,N_6347);
nand U6563 (N_6563,N_6080,N_6473);
and U6564 (N_6564,N_6466,N_6495);
or U6565 (N_6565,N_6487,N_6002);
xor U6566 (N_6566,N_6231,N_6017);
nor U6567 (N_6567,N_6001,N_6090);
nor U6568 (N_6568,N_6422,N_6039);
nor U6569 (N_6569,N_6427,N_6394);
or U6570 (N_6570,N_6221,N_6492);
and U6571 (N_6571,N_6277,N_6026);
or U6572 (N_6572,N_6246,N_6322);
nand U6573 (N_6573,N_6280,N_6145);
xnor U6574 (N_6574,N_6193,N_6467);
and U6575 (N_6575,N_6393,N_6058);
and U6576 (N_6576,N_6343,N_6279);
xor U6577 (N_6577,N_6468,N_6416);
and U6578 (N_6578,N_6488,N_6348);
nor U6579 (N_6579,N_6332,N_6212);
or U6580 (N_6580,N_6066,N_6325);
nand U6581 (N_6581,N_6084,N_6117);
nand U6582 (N_6582,N_6268,N_6047);
xnor U6583 (N_6583,N_6292,N_6426);
xnor U6584 (N_6584,N_6059,N_6251);
or U6585 (N_6585,N_6143,N_6146);
nand U6586 (N_6586,N_6176,N_6284);
nor U6587 (N_6587,N_6433,N_6445);
or U6588 (N_6588,N_6285,N_6226);
or U6589 (N_6589,N_6384,N_6060);
nor U6590 (N_6590,N_6095,N_6316);
nand U6591 (N_6591,N_6377,N_6186);
nor U6592 (N_6592,N_6014,N_6388);
nor U6593 (N_6593,N_6301,N_6077);
xnor U6594 (N_6594,N_6359,N_6052);
nand U6595 (N_6595,N_6409,N_6112);
nor U6596 (N_6596,N_6314,N_6350);
nand U6597 (N_6597,N_6025,N_6125);
nor U6598 (N_6598,N_6009,N_6327);
nor U6599 (N_6599,N_6229,N_6010);
xor U6600 (N_6600,N_6204,N_6414);
xor U6601 (N_6601,N_6340,N_6195);
and U6602 (N_6602,N_6455,N_6183);
nand U6603 (N_6603,N_6015,N_6448);
nand U6604 (N_6604,N_6190,N_6034);
and U6605 (N_6605,N_6135,N_6230);
nor U6606 (N_6606,N_6153,N_6369);
nor U6607 (N_6607,N_6179,N_6214);
xor U6608 (N_6608,N_6345,N_6057);
nor U6609 (N_6609,N_6197,N_6263);
nand U6610 (N_6610,N_6037,N_6429);
nand U6611 (N_6611,N_6418,N_6373);
nand U6612 (N_6612,N_6368,N_6387);
nand U6613 (N_6613,N_6425,N_6028);
nand U6614 (N_6614,N_6400,N_6496);
or U6615 (N_6615,N_6452,N_6115);
and U6616 (N_6616,N_6064,N_6118);
nor U6617 (N_6617,N_6420,N_6103);
or U6618 (N_6618,N_6106,N_6130);
or U6619 (N_6619,N_6375,N_6443);
nand U6620 (N_6620,N_6180,N_6120);
and U6621 (N_6621,N_6031,N_6259);
and U6622 (N_6622,N_6087,N_6199);
or U6623 (N_6623,N_6141,N_6211);
and U6624 (N_6624,N_6318,N_6385);
or U6625 (N_6625,N_6151,N_6024);
nand U6626 (N_6626,N_6004,N_6353);
nand U6627 (N_6627,N_6294,N_6357);
or U6628 (N_6628,N_6248,N_6016);
nor U6629 (N_6629,N_6022,N_6485);
nand U6630 (N_6630,N_6123,N_6242);
xnor U6631 (N_6631,N_6124,N_6147);
nand U6632 (N_6632,N_6269,N_6027);
or U6633 (N_6633,N_6220,N_6479);
and U6634 (N_6634,N_6354,N_6021);
and U6635 (N_6635,N_6484,N_6356);
nand U6636 (N_6636,N_6011,N_6313);
and U6637 (N_6637,N_6481,N_6293);
or U6638 (N_6638,N_6288,N_6489);
xnor U6639 (N_6639,N_6309,N_6094);
or U6640 (N_6640,N_6444,N_6140);
nor U6641 (N_6641,N_6249,N_6191);
xnor U6642 (N_6642,N_6225,N_6018);
and U6643 (N_6643,N_6083,N_6255);
nand U6644 (N_6644,N_6235,N_6207);
xnor U6645 (N_6645,N_6096,N_6049);
nand U6646 (N_6646,N_6472,N_6097);
nand U6647 (N_6647,N_6303,N_6475);
nand U6648 (N_6648,N_6072,N_6323);
xor U6649 (N_6649,N_6042,N_6074);
and U6650 (N_6650,N_6114,N_6266);
or U6651 (N_6651,N_6260,N_6478);
and U6652 (N_6652,N_6304,N_6349);
or U6653 (N_6653,N_6440,N_6419);
xor U6654 (N_6654,N_6132,N_6477);
or U6655 (N_6655,N_6331,N_6244);
or U6656 (N_6656,N_6460,N_6395);
and U6657 (N_6657,N_6447,N_6165);
nor U6658 (N_6658,N_6228,N_6110);
or U6659 (N_6659,N_6296,N_6274);
and U6660 (N_6660,N_6182,N_6234);
nor U6661 (N_6661,N_6490,N_6121);
nand U6662 (N_6662,N_6202,N_6454);
xnor U6663 (N_6663,N_6321,N_6215);
and U6664 (N_6664,N_6270,N_6453);
nand U6665 (N_6665,N_6434,N_6439);
xnor U6666 (N_6666,N_6257,N_6370);
or U6667 (N_6667,N_6203,N_6337);
and U6668 (N_6668,N_6075,N_6320);
nor U6669 (N_6669,N_6273,N_6360);
xor U6670 (N_6670,N_6302,N_6402);
or U6671 (N_6671,N_6088,N_6282);
nand U6672 (N_6672,N_6254,N_6069);
nand U6673 (N_6673,N_6315,N_6161);
xnor U6674 (N_6674,N_6371,N_6019);
and U6675 (N_6675,N_6381,N_6201);
nand U6676 (N_6676,N_6290,N_6372);
and U6677 (N_6677,N_6119,N_6243);
or U6678 (N_6678,N_6136,N_6405);
xnor U6679 (N_6679,N_6020,N_6365);
and U6680 (N_6680,N_6287,N_6188);
and U6681 (N_6681,N_6181,N_6374);
and U6682 (N_6682,N_6056,N_6358);
nor U6683 (N_6683,N_6089,N_6073);
and U6684 (N_6684,N_6459,N_6312);
or U6685 (N_6685,N_6086,N_6079);
and U6686 (N_6686,N_6464,N_6341);
nand U6687 (N_6687,N_6438,N_6382);
nor U6688 (N_6688,N_6196,N_6178);
xor U6689 (N_6689,N_6048,N_6227);
and U6690 (N_6690,N_6092,N_6408);
or U6691 (N_6691,N_6205,N_6168);
nand U6692 (N_6692,N_6396,N_6175);
or U6693 (N_6693,N_6099,N_6363);
xor U6694 (N_6694,N_6023,N_6298);
and U6695 (N_6695,N_6013,N_6082);
nand U6696 (N_6696,N_6275,N_6458);
or U6697 (N_6697,N_6436,N_6177);
or U6698 (N_6698,N_6421,N_6036);
xnor U6699 (N_6699,N_6149,N_6256);
or U6700 (N_6700,N_6093,N_6012);
xnor U6701 (N_6701,N_6055,N_6078);
or U6702 (N_6702,N_6398,N_6213);
nand U6703 (N_6703,N_6399,N_6160);
nand U6704 (N_6704,N_6035,N_6200);
and U6705 (N_6705,N_6157,N_6401);
or U6706 (N_6706,N_6162,N_6102);
xor U6707 (N_6707,N_6334,N_6192);
nand U6708 (N_6708,N_6107,N_6339);
or U6709 (N_6709,N_6174,N_6194);
xor U6710 (N_6710,N_6116,N_6129);
and U6711 (N_6711,N_6499,N_6378);
xor U6712 (N_6712,N_6297,N_6471);
nand U6713 (N_6713,N_6217,N_6252);
xor U6714 (N_6714,N_6131,N_6462);
nand U6715 (N_6715,N_6480,N_6169);
and U6716 (N_6716,N_6335,N_6403);
nor U6717 (N_6717,N_6355,N_6367);
xnor U6718 (N_6718,N_6167,N_6240);
nand U6719 (N_6719,N_6430,N_6474);
nand U6720 (N_6720,N_6404,N_6003);
nand U6721 (N_6721,N_6000,N_6232);
xor U6722 (N_6722,N_6451,N_6307);
nor U6723 (N_6723,N_6344,N_6158);
xor U6724 (N_6724,N_6100,N_6238);
xnor U6725 (N_6725,N_6187,N_6351);
or U6726 (N_6726,N_6392,N_6383);
or U6727 (N_6727,N_6278,N_6258);
and U6728 (N_6728,N_6361,N_6170);
xor U6729 (N_6729,N_6482,N_6101);
xor U6730 (N_6730,N_6108,N_6241);
and U6731 (N_6731,N_6218,N_6154);
and U6732 (N_6732,N_6065,N_6008);
nand U6733 (N_6733,N_6435,N_6424);
nand U6734 (N_6734,N_6030,N_6171);
or U6735 (N_6735,N_6272,N_6456);
and U6736 (N_6736,N_6397,N_6497);
or U6737 (N_6737,N_6446,N_6342);
nand U6738 (N_6738,N_6291,N_6085);
nor U6739 (N_6739,N_6289,N_6237);
or U6740 (N_6740,N_6127,N_6262);
nor U6741 (N_6741,N_6417,N_6391);
nand U6742 (N_6742,N_6346,N_6267);
xor U6743 (N_6743,N_6457,N_6326);
and U6744 (N_6744,N_6390,N_6032);
or U6745 (N_6745,N_6299,N_6362);
xnor U6746 (N_6746,N_6253,N_6441);
and U6747 (N_6747,N_6224,N_6450);
and U6748 (N_6748,N_6442,N_6306);
xor U6749 (N_6749,N_6494,N_6111);
nand U6750 (N_6750,N_6157,N_6456);
nand U6751 (N_6751,N_6213,N_6106);
nor U6752 (N_6752,N_6245,N_6156);
and U6753 (N_6753,N_6239,N_6021);
and U6754 (N_6754,N_6103,N_6068);
nand U6755 (N_6755,N_6221,N_6161);
nor U6756 (N_6756,N_6393,N_6154);
or U6757 (N_6757,N_6435,N_6102);
or U6758 (N_6758,N_6205,N_6007);
or U6759 (N_6759,N_6106,N_6478);
xnor U6760 (N_6760,N_6260,N_6180);
and U6761 (N_6761,N_6204,N_6254);
nor U6762 (N_6762,N_6356,N_6314);
nand U6763 (N_6763,N_6415,N_6013);
xnor U6764 (N_6764,N_6478,N_6385);
or U6765 (N_6765,N_6139,N_6351);
nand U6766 (N_6766,N_6286,N_6143);
nand U6767 (N_6767,N_6432,N_6283);
xnor U6768 (N_6768,N_6198,N_6411);
and U6769 (N_6769,N_6127,N_6214);
nand U6770 (N_6770,N_6318,N_6327);
nor U6771 (N_6771,N_6163,N_6433);
or U6772 (N_6772,N_6245,N_6330);
xnor U6773 (N_6773,N_6008,N_6251);
and U6774 (N_6774,N_6153,N_6126);
xnor U6775 (N_6775,N_6179,N_6431);
xnor U6776 (N_6776,N_6323,N_6210);
nand U6777 (N_6777,N_6059,N_6014);
and U6778 (N_6778,N_6214,N_6245);
nor U6779 (N_6779,N_6237,N_6172);
nor U6780 (N_6780,N_6146,N_6154);
nor U6781 (N_6781,N_6349,N_6295);
nand U6782 (N_6782,N_6372,N_6086);
xnor U6783 (N_6783,N_6480,N_6104);
or U6784 (N_6784,N_6334,N_6341);
or U6785 (N_6785,N_6233,N_6404);
nor U6786 (N_6786,N_6132,N_6322);
nor U6787 (N_6787,N_6133,N_6282);
nand U6788 (N_6788,N_6193,N_6408);
xnor U6789 (N_6789,N_6210,N_6462);
or U6790 (N_6790,N_6234,N_6266);
nand U6791 (N_6791,N_6351,N_6142);
and U6792 (N_6792,N_6063,N_6410);
nand U6793 (N_6793,N_6348,N_6195);
nor U6794 (N_6794,N_6377,N_6037);
or U6795 (N_6795,N_6168,N_6345);
nor U6796 (N_6796,N_6349,N_6231);
xor U6797 (N_6797,N_6011,N_6481);
or U6798 (N_6798,N_6215,N_6252);
and U6799 (N_6799,N_6262,N_6173);
xnor U6800 (N_6800,N_6171,N_6109);
xnor U6801 (N_6801,N_6181,N_6382);
xnor U6802 (N_6802,N_6188,N_6009);
nand U6803 (N_6803,N_6291,N_6357);
nor U6804 (N_6804,N_6104,N_6370);
xnor U6805 (N_6805,N_6471,N_6425);
xnor U6806 (N_6806,N_6213,N_6293);
or U6807 (N_6807,N_6221,N_6465);
nor U6808 (N_6808,N_6062,N_6426);
nor U6809 (N_6809,N_6320,N_6246);
and U6810 (N_6810,N_6066,N_6044);
or U6811 (N_6811,N_6485,N_6088);
xnor U6812 (N_6812,N_6290,N_6243);
and U6813 (N_6813,N_6082,N_6006);
nor U6814 (N_6814,N_6361,N_6130);
xor U6815 (N_6815,N_6223,N_6338);
or U6816 (N_6816,N_6131,N_6328);
xnor U6817 (N_6817,N_6287,N_6097);
xnor U6818 (N_6818,N_6306,N_6123);
xnor U6819 (N_6819,N_6404,N_6312);
and U6820 (N_6820,N_6459,N_6070);
xor U6821 (N_6821,N_6121,N_6260);
nor U6822 (N_6822,N_6203,N_6065);
and U6823 (N_6823,N_6339,N_6350);
and U6824 (N_6824,N_6042,N_6356);
xor U6825 (N_6825,N_6148,N_6497);
or U6826 (N_6826,N_6247,N_6229);
nand U6827 (N_6827,N_6194,N_6190);
nand U6828 (N_6828,N_6129,N_6336);
and U6829 (N_6829,N_6241,N_6089);
and U6830 (N_6830,N_6115,N_6084);
nand U6831 (N_6831,N_6380,N_6257);
and U6832 (N_6832,N_6116,N_6382);
and U6833 (N_6833,N_6130,N_6053);
xor U6834 (N_6834,N_6210,N_6350);
nand U6835 (N_6835,N_6432,N_6229);
nand U6836 (N_6836,N_6225,N_6168);
nand U6837 (N_6837,N_6172,N_6041);
nor U6838 (N_6838,N_6431,N_6412);
and U6839 (N_6839,N_6455,N_6049);
nand U6840 (N_6840,N_6029,N_6479);
nand U6841 (N_6841,N_6305,N_6214);
nand U6842 (N_6842,N_6496,N_6482);
xnor U6843 (N_6843,N_6461,N_6125);
and U6844 (N_6844,N_6404,N_6308);
or U6845 (N_6845,N_6484,N_6033);
nand U6846 (N_6846,N_6063,N_6452);
or U6847 (N_6847,N_6222,N_6141);
nand U6848 (N_6848,N_6188,N_6189);
or U6849 (N_6849,N_6250,N_6259);
and U6850 (N_6850,N_6144,N_6024);
or U6851 (N_6851,N_6398,N_6196);
xor U6852 (N_6852,N_6129,N_6050);
and U6853 (N_6853,N_6148,N_6298);
nand U6854 (N_6854,N_6180,N_6078);
and U6855 (N_6855,N_6488,N_6259);
nand U6856 (N_6856,N_6308,N_6405);
xnor U6857 (N_6857,N_6189,N_6419);
xnor U6858 (N_6858,N_6398,N_6247);
nor U6859 (N_6859,N_6309,N_6272);
or U6860 (N_6860,N_6142,N_6306);
or U6861 (N_6861,N_6322,N_6385);
xor U6862 (N_6862,N_6427,N_6115);
nand U6863 (N_6863,N_6445,N_6205);
nor U6864 (N_6864,N_6160,N_6126);
or U6865 (N_6865,N_6267,N_6432);
or U6866 (N_6866,N_6424,N_6416);
or U6867 (N_6867,N_6284,N_6285);
or U6868 (N_6868,N_6374,N_6224);
xnor U6869 (N_6869,N_6032,N_6136);
nand U6870 (N_6870,N_6164,N_6407);
and U6871 (N_6871,N_6112,N_6414);
nand U6872 (N_6872,N_6320,N_6206);
and U6873 (N_6873,N_6185,N_6369);
xor U6874 (N_6874,N_6210,N_6429);
xnor U6875 (N_6875,N_6249,N_6177);
or U6876 (N_6876,N_6354,N_6141);
or U6877 (N_6877,N_6244,N_6447);
or U6878 (N_6878,N_6181,N_6130);
nor U6879 (N_6879,N_6496,N_6353);
and U6880 (N_6880,N_6381,N_6024);
and U6881 (N_6881,N_6100,N_6263);
or U6882 (N_6882,N_6323,N_6216);
nor U6883 (N_6883,N_6481,N_6461);
and U6884 (N_6884,N_6337,N_6316);
nand U6885 (N_6885,N_6425,N_6289);
nor U6886 (N_6886,N_6217,N_6124);
xnor U6887 (N_6887,N_6324,N_6422);
xnor U6888 (N_6888,N_6243,N_6417);
and U6889 (N_6889,N_6413,N_6138);
xnor U6890 (N_6890,N_6488,N_6123);
nand U6891 (N_6891,N_6169,N_6448);
xor U6892 (N_6892,N_6391,N_6376);
xnor U6893 (N_6893,N_6080,N_6086);
and U6894 (N_6894,N_6111,N_6363);
nor U6895 (N_6895,N_6044,N_6314);
or U6896 (N_6896,N_6309,N_6051);
and U6897 (N_6897,N_6189,N_6146);
nor U6898 (N_6898,N_6172,N_6206);
or U6899 (N_6899,N_6196,N_6479);
and U6900 (N_6900,N_6029,N_6437);
nor U6901 (N_6901,N_6038,N_6177);
nand U6902 (N_6902,N_6285,N_6188);
and U6903 (N_6903,N_6001,N_6004);
xnor U6904 (N_6904,N_6239,N_6294);
xnor U6905 (N_6905,N_6182,N_6350);
nand U6906 (N_6906,N_6071,N_6285);
or U6907 (N_6907,N_6308,N_6180);
xnor U6908 (N_6908,N_6169,N_6359);
nand U6909 (N_6909,N_6403,N_6166);
nor U6910 (N_6910,N_6482,N_6411);
xor U6911 (N_6911,N_6300,N_6371);
nand U6912 (N_6912,N_6472,N_6070);
xor U6913 (N_6913,N_6283,N_6294);
or U6914 (N_6914,N_6404,N_6052);
nand U6915 (N_6915,N_6419,N_6490);
xor U6916 (N_6916,N_6292,N_6154);
nor U6917 (N_6917,N_6326,N_6464);
or U6918 (N_6918,N_6091,N_6116);
xnor U6919 (N_6919,N_6479,N_6069);
xor U6920 (N_6920,N_6090,N_6026);
and U6921 (N_6921,N_6421,N_6434);
or U6922 (N_6922,N_6333,N_6126);
nand U6923 (N_6923,N_6000,N_6433);
nand U6924 (N_6924,N_6221,N_6326);
nand U6925 (N_6925,N_6068,N_6185);
or U6926 (N_6926,N_6184,N_6295);
nor U6927 (N_6927,N_6018,N_6341);
or U6928 (N_6928,N_6275,N_6174);
xnor U6929 (N_6929,N_6045,N_6071);
nand U6930 (N_6930,N_6250,N_6430);
and U6931 (N_6931,N_6220,N_6070);
nand U6932 (N_6932,N_6132,N_6188);
or U6933 (N_6933,N_6431,N_6376);
nor U6934 (N_6934,N_6070,N_6391);
nand U6935 (N_6935,N_6227,N_6459);
xor U6936 (N_6936,N_6417,N_6052);
and U6937 (N_6937,N_6270,N_6386);
and U6938 (N_6938,N_6408,N_6126);
xor U6939 (N_6939,N_6054,N_6023);
nor U6940 (N_6940,N_6433,N_6085);
and U6941 (N_6941,N_6057,N_6049);
xnor U6942 (N_6942,N_6127,N_6331);
xnor U6943 (N_6943,N_6197,N_6439);
or U6944 (N_6944,N_6163,N_6115);
xor U6945 (N_6945,N_6211,N_6208);
nand U6946 (N_6946,N_6451,N_6310);
nand U6947 (N_6947,N_6450,N_6375);
nor U6948 (N_6948,N_6351,N_6362);
and U6949 (N_6949,N_6394,N_6470);
xor U6950 (N_6950,N_6493,N_6148);
nor U6951 (N_6951,N_6269,N_6342);
xnor U6952 (N_6952,N_6001,N_6455);
and U6953 (N_6953,N_6043,N_6323);
and U6954 (N_6954,N_6232,N_6306);
and U6955 (N_6955,N_6221,N_6035);
or U6956 (N_6956,N_6093,N_6339);
nor U6957 (N_6957,N_6331,N_6454);
nand U6958 (N_6958,N_6241,N_6198);
xnor U6959 (N_6959,N_6287,N_6103);
xor U6960 (N_6960,N_6345,N_6179);
and U6961 (N_6961,N_6102,N_6082);
and U6962 (N_6962,N_6293,N_6298);
nor U6963 (N_6963,N_6219,N_6193);
nor U6964 (N_6964,N_6461,N_6296);
or U6965 (N_6965,N_6314,N_6325);
or U6966 (N_6966,N_6264,N_6435);
xnor U6967 (N_6967,N_6367,N_6191);
and U6968 (N_6968,N_6081,N_6067);
xor U6969 (N_6969,N_6036,N_6082);
and U6970 (N_6970,N_6212,N_6019);
or U6971 (N_6971,N_6159,N_6119);
nor U6972 (N_6972,N_6143,N_6312);
nand U6973 (N_6973,N_6327,N_6050);
and U6974 (N_6974,N_6196,N_6361);
xor U6975 (N_6975,N_6197,N_6221);
nor U6976 (N_6976,N_6420,N_6360);
nand U6977 (N_6977,N_6277,N_6293);
and U6978 (N_6978,N_6413,N_6373);
nand U6979 (N_6979,N_6474,N_6230);
and U6980 (N_6980,N_6285,N_6448);
nor U6981 (N_6981,N_6460,N_6363);
xor U6982 (N_6982,N_6369,N_6323);
or U6983 (N_6983,N_6219,N_6215);
xor U6984 (N_6984,N_6152,N_6028);
xor U6985 (N_6985,N_6145,N_6126);
or U6986 (N_6986,N_6346,N_6392);
xnor U6987 (N_6987,N_6320,N_6066);
xnor U6988 (N_6988,N_6235,N_6365);
xnor U6989 (N_6989,N_6084,N_6131);
xnor U6990 (N_6990,N_6015,N_6056);
nand U6991 (N_6991,N_6391,N_6460);
nand U6992 (N_6992,N_6314,N_6208);
or U6993 (N_6993,N_6108,N_6255);
nand U6994 (N_6994,N_6398,N_6201);
or U6995 (N_6995,N_6002,N_6044);
or U6996 (N_6996,N_6182,N_6023);
and U6997 (N_6997,N_6341,N_6433);
nor U6998 (N_6998,N_6360,N_6455);
and U6999 (N_6999,N_6446,N_6336);
nand U7000 (N_7000,N_6644,N_6689);
xnor U7001 (N_7001,N_6720,N_6626);
nand U7002 (N_7002,N_6664,N_6642);
and U7003 (N_7003,N_6566,N_6676);
xnor U7004 (N_7004,N_6908,N_6994);
nand U7005 (N_7005,N_6820,N_6600);
xor U7006 (N_7006,N_6909,N_6957);
xor U7007 (N_7007,N_6598,N_6625);
nor U7008 (N_7008,N_6687,N_6883);
nor U7009 (N_7009,N_6907,N_6973);
xnor U7010 (N_7010,N_6694,N_6692);
nand U7011 (N_7011,N_6997,N_6649);
nand U7012 (N_7012,N_6551,N_6502);
nor U7013 (N_7013,N_6951,N_6861);
and U7014 (N_7014,N_6967,N_6990);
xor U7015 (N_7015,N_6670,N_6872);
nand U7016 (N_7016,N_6842,N_6607);
xnor U7017 (N_7017,N_6846,N_6518);
nor U7018 (N_7018,N_6901,N_6933);
nand U7019 (N_7019,N_6851,N_6511);
nand U7020 (N_7020,N_6586,N_6709);
and U7021 (N_7021,N_6583,N_6891);
and U7022 (N_7022,N_6595,N_6897);
or U7023 (N_7023,N_6950,N_6879);
or U7024 (N_7024,N_6674,N_6555);
or U7025 (N_7025,N_6584,N_6622);
xor U7026 (N_7026,N_6758,N_6612);
nor U7027 (N_7027,N_6984,N_6700);
nor U7028 (N_7028,N_6970,N_6911);
and U7029 (N_7029,N_6747,N_6614);
nor U7030 (N_7030,N_6636,N_6749);
nor U7031 (N_7031,N_6756,N_6778);
or U7032 (N_7032,N_6885,N_6718);
nor U7033 (N_7033,N_6560,N_6647);
or U7034 (N_7034,N_6886,N_6619);
and U7035 (N_7035,N_6661,N_6991);
xnor U7036 (N_7036,N_6524,N_6638);
nor U7037 (N_7037,N_6793,N_6734);
nand U7038 (N_7038,N_6982,N_6882);
nand U7039 (N_7039,N_6937,N_6579);
nand U7040 (N_7040,N_6591,N_6760);
nand U7041 (N_7041,N_6998,N_6923);
or U7042 (N_7042,N_6724,N_6903);
xor U7043 (N_7043,N_6547,N_6877);
or U7044 (N_7044,N_6863,N_6854);
nor U7045 (N_7045,N_6837,N_6505);
and U7046 (N_7046,N_6730,N_6787);
and U7047 (N_7047,N_6823,N_6735);
or U7048 (N_7048,N_6828,N_6862);
or U7049 (N_7049,N_6704,N_6605);
xnor U7050 (N_7050,N_6643,N_6705);
xnor U7051 (N_7051,N_6815,N_6752);
or U7052 (N_7052,N_6578,N_6766);
nand U7053 (N_7053,N_6898,N_6880);
xnor U7054 (N_7054,N_6889,N_6573);
xnor U7055 (N_7055,N_6918,N_6721);
xnor U7056 (N_7056,N_6552,N_6904);
or U7057 (N_7057,N_6796,N_6504);
and U7058 (N_7058,N_6969,N_6727);
or U7059 (N_7059,N_6627,N_6731);
and U7060 (N_7060,N_6672,N_6921);
xor U7061 (N_7061,N_6603,N_6895);
or U7062 (N_7062,N_6819,N_6826);
and U7063 (N_7063,N_6517,N_6784);
or U7064 (N_7064,N_6804,N_6532);
nand U7065 (N_7065,N_6917,N_6609);
nand U7066 (N_7066,N_6572,N_6596);
and U7067 (N_7067,N_6816,N_6963);
xnor U7068 (N_7068,N_6745,N_6725);
nor U7069 (N_7069,N_6686,N_6769);
nor U7070 (N_7070,N_6681,N_6941);
or U7071 (N_7071,N_6812,N_6748);
xnor U7072 (N_7072,N_6830,N_6601);
nand U7073 (N_7073,N_6671,N_6629);
and U7074 (N_7074,N_6719,N_6557);
or U7075 (N_7075,N_6558,N_6870);
nor U7076 (N_7076,N_6651,N_6853);
and U7077 (N_7077,N_6988,N_6798);
or U7078 (N_7078,N_6976,N_6836);
and U7079 (N_7079,N_6543,N_6590);
or U7080 (N_7080,N_6500,N_6945);
or U7081 (N_7081,N_6639,N_6953);
xnor U7082 (N_7082,N_6996,N_6993);
nor U7083 (N_7083,N_6809,N_6977);
or U7084 (N_7084,N_6866,N_6736);
nand U7085 (N_7085,N_6553,N_6635);
nand U7086 (N_7086,N_6768,N_6949);
nor U7087 (N_7087,N_6956,N_6852);
or U7088 (N_7088,N_6599,N_6657);
xor U7089 (N_7089,N_6764,N_6806);
and U7090 (N_7090,N_6569,N_6624);
nor U7091 (N_7091,N_6890,N_6631);
or U7092 (N_7092,N_6811,N_6845);
and U7093 (N_7093,N_6662,N_6737);
or U7094 (N_7094,N_6722,N_6763);
nand U7095 (N_7095,N_6777,N_6506);
xnor U7096 (N_7096,N_6936,N_6801);
and U7097 (N_7097,N_6754,N_6652);
and U7098 (N_7098,N_6654,N_6920);
or U7099 (N_7099,N_6790,N_6582);
xor U7100 (N_7100,N_6893,N_6633);
nor U7101 (N_7101,N_6539,N_6684);
and U7102 (N_7102,N_6519,N_6608);
nor U7103 (N_7103,N_6986,N_6912);
nand U7104 (N_7104,N_6833,N_6646);
or U7105 (N_7105,N_6992,N_6868);
or U7106 (N_7106,N_6881,N_6514);
or U7107 (N_7107,N_6628,N_6932);
nor U7108 (N_7108,N_6744,N_6947);
and U7109 (N_7109,N_6981,N_6844);
nor U7110 (N_7110,N_6847,N_6813);
or U7111 (N_7111,N_6562,N_6630);
nand U7112 (N_7112,N_6924,N_6857);
nand U7113 (N_7113,N_6894,N_6783);
nand U7114 (N_7114,N_6860,N_6888);
xor U7115 (N_7115,N_6803,N_6577);
and U7116 (N_7116,N_6856,N_6964);
or U7117 (N_7117,N_6699,N_6508);
or U7118 (N_7118,N_6799,N_6703);
nand U7119 (N_7119,N_6979,N_6713);
xnor U7120 (N_7120,N_6968,N_6959);
or U7121 (N_7121,N_6697,N_6960);
and U7122 (N_7122,N_6567,N_6791);
nor U7123 (N_7123,N_6915,N_6850);
nor U7124 (N_7124,N_6873,N_6930);
xnor U7125 (N_7125,N_6869,N_6954);
and U7126 (N_7126,N_6773,N_6528);
nand U7127 (N_7127,N_6696,N_6789);
xnor U7128 (N_7128,N_6935,N_6871);
and U7129 (N_7129,N_6714,N_6822);
or U7130 (N_7130,N_6556,N_6807);
nor U7131 (N_7131,N_6702,N_6645);
nand U7132 (N_7132,N_6542,N_6554);
xnor U7133 (N_7133,N_6685,N_6559);
and U7134 (N_7134,N_6529,N_6641);
or U7135 (N_7135,N_6565,N_6540);
and U7136 (N_7136,N_6824,N_6733);
and U7137 (N_7137,N_6527,N_6995);
nor U7138 (N_7138,N_6876,N_6669);
or U7139 (N_7139,N_6623,N_6865);
and U7140 (N_7140,N_6800,N_6825);
nand U7141 (N_7141,N_6564,N_6576);
or U7142 (N_7142,N_6738,N_6952);
nor U7143 (N_7143,N_6905,N_6606);
and U7144 (N_7144,N_6653,N_6667);
nand U7145 (N_7145,N_6677,N_6743);
or U7146 (N_7146,N_6940,N_6843);
nor U7147 (N_7147,N_6588,N_6831);
nand U7148 (N_7148,N_6634,N_6617);
xnor U7149 (N_7149,N_6544,N_6928);
xnor U7150 (N_7150,N_6919,N_6966);
and U7151 (N_7151,N_6761,N_6975);
and U7152 (N_7152,N_6516,N_6759);
and U7153 (N_7153,N_6691,N_6929);
nor U7154 (N_7154,N_6550,N_6711);
nor U7155 (N_7155,N_6538,N_6510);
xor U7156 (N_7156,N_6729,N_6663);
or U7157 (N_7157,N_6575,N_6536);
nor U7158 (N_7158,N_6568,N_6770);
or U7159 (N_7159,N_6814,N_6563);
nor U7160 (N_7160,N_6695,N_6827);
nor U7161 (N_7161,N_6741,N_6618);
nand U7162 (N_7162,N_6834,N_6802);
nand U7163 (N_7163,N_6513,N_6916);
nand U7164 (N_7164,N_6978,N_6808);
xor U7165 (N_7165,N_6840,N_6678);
and U7166 (N_7166,N_6580,N_6776);
or U7167 (N_7167,N_6765,N_6708);
and U7168 (N_7168,N_6999,N_6795);
and U7169 (N_7169,N_6987,N_6611);
nand U7170 (N_7170,N_6512,N_6680);
nor U7171 (N_7171,N_6589,N_6955);
xor U7172 (N_7172,N_6707,N_6613);
nand U7173 (N_7173,N_6523,N_6531);
nand U7174 (N_7174,N_6779,N_6878);
xor U7175 (N_7175,N_6925,N_6509);
xnor U7176 (N_7176,N_6659,N_6922);
and U7177 (N_7177,N_6537,N_6726);
nand U7178 (N_7178,N_6515,N_6530);
and U7179 (N_7179,N_6698,N_6739);
and U7180 (N_7180,N_6810,N_6906);
and U7181 (N_7181,N_6821,N_6602);
nand U7182 (N_7182,N_6574,N_6805);
xnor U7183 (N_7183,N_6546,N_6835);
and U7184 (N_7184,N_6867,N_6794);
nand U7185 (N_7185,N_6679,N_6971);
nand U7186 (N_7186,N_6774,N_6874);
nor U7187 (N_7187,N_6887,N_6660);
nor U7188 (N_7188,N_6655,N_6855);
nor U7189 (N_7189,N_6712,N_6535);
or U7190 (N_7190,N_6946,N_6864);
nand U7191 (N_7191,N_6859,N_6632);
nand U7192 (N_7192,N_6750,N_6688);
nand U7193 (N_7193,N_6767,N_6533);
nor U7194 (N_7194,N_6728,N_6525);
nand U7195 (N_7195,N_6785,N_6594);
and U7196 (N_7196,N_6939,N_6772);
nor U7197 (N_7197,N_6792,N_6829);
and U7198 (N_7198,N_6899,N_6587);
or U7199 (N_7199,N_6896,N_6507);
and U7200 (N_7200,N_6710,N_6561);
nor U7201 (N_7201,N_6526,N_6665);
or U7202 (N_7202,N_6549,N_6501);
nor U7203 (N_7203,N_6974,N_6775);
or U7204 (N_7204,N_6521,N_6944);
nand U7205 (N_7205,N_6961,N_6934);
nor U7206 (N_7206,N_6656,N_6604);
nor U7207 (N_7207,N_6658,N_6597);
or U7208 (N_7208,N_6640,N_6541);
or U7209 (N_7209,N_6927,N_6548);
nor U7210 (N_7210,N_6786,N_6690);
or U7211 (N_7211,N_6781,N_6943);
or U7212 (N_7212,N_6962,N_6782);
and U7213 (N_7213,N_6972,N_6818);
nor U7214 (N_7214,N_6980,N_6958);
nand U7215 (N_7215,N_6817,N_6938);
nand U7216 (N_7216,N_6610,N_6838);
nor U7217 (N_7217,N_6910,N_6965);
nor U7218 (N_7218,N_6788,N_6780);
xnor U7219 (N_7219,N_6742,N_6637);
nor U7220 (N_7220,N_6701,N_6682);
nand U7221 (N_7221,N_6585,N_6884);
and U7222 (N_7222,N_6948,N_6545);
nor U7223 (N_7223,N_6732,N_6650);
and U7224 (N_7224,N_6648,N_6683);
nand U7225 (N_7225,N_6615,N_6740);
xnor U7226 (N_7226,N_6848,N_6875);
and U7227 (N_7227,N_6931,N_6985);
nand U7228 (N_7228,N_6751,N_6716);
nor U7229 (N_7229,N_6771,N_6841);
or U7230 (N_7230,N_6849,N_6746);
nor U7231 (N_7231,N_6753,N_6673);
or U7232 (N_7232,N_6620,N_6616);
xor U7233 (N_7233,N_6693,N_6762);
nand U7234 (N_7234,N_6717,N_6892);
and U7235 (N_7235,N_6839,N_6706);
xnor U7236 (N_7236,N_6571,N_6723);
xnor U7237 (N_7237,N_6942,N_6715);
and U7238 (N_7238,N_6621,N_6593);
nor U7239 (N_7239,N_6926,N_6797);
nor U7240 (N_7240,N_6858,N_6913);
and U7241 (N_7241,N_6592,N_6520);
or U7242 (N_7242,N_6989,N_6755);
xor U7243 (N_7243,N_6902,N_6832);
xor U7244 (N_7244,N_6914,N_6666);
or U7245 (N_7245,N_6570,N_6534);
nand U7246 (N_7246,N_6757,N_6983);
xor U7247 (N_7247,N_6581,N_6668);
xnor U7248 (N_7248,N_6675,N_6522);
and U7249 (N_7249,N_6503,N_6900);
xnor U7250 (N_7250,N_6974,N_6590);
or U7251 (N_7251,N_6773,N_6877);
xnor U7252 (N_7252,N_6895,N_6884);
or U7253 (N_7253,N_6615,N_6509);
nand U7254 (N_7254,N_6527,N_6771);
and U7255 (N_7255,N_6845,N_6751);
and U7256 (N_7256,N_6886,N_6577);
and U7257 (N_7257,N_6803,N_6513);
and U7258 (N_7258,N_6715,N_6636);
or U7259 (N_7259,N_6571,N_6764);
xnor U7260 (N_7260,N_6665,N_6980);
xnor U7261 (N_7261,N_6970,N_6536);
nand U7262 (N_7262,N_6935,N_6755);
nand U7263 (N_7263,N_6768,N_6504);
or U7264 (N_7264,N_6770,N_6560);
nor U7265 (N_7265,N_6556,N_6962);
or U7266 (N_7266,N_6932,N_6689);
xnor U7267 (N_7267,N_6907,N_6676);
and U7268 (N_7268,N_6718,N_6666);
or U7269 (N_7269,N_6881,N_6896);
or U7270 (N_7270,N_6515,N_6688);
and U7271 (N_7271,N_6639,N_6574);
nand U7272 (N_7272,N_6965,N_6593);
and U7273 (N_7273,N_6636,N_6750);
nand U7274 (N_7274,N_6690,N_6500);
xnor U7275 (N_7275,N_6611,N_6968);
nor U7276 (N_7276,N_6914,N_6854);
nand U7277 (N_7277,N_6624,N_6709);
nor U7278 (N_7278,N_6730,N_6774);
or U7279 (N_7279,N_6664,N_6562);
nand U7280 (N_7280,N_6573,N_6957);
xnor U7281 (N_7281,N_6551,N_6918);
xor U7282 (N_7282,N_6863,N_6674);
nor U7283 (N_7283,N_6693,N_6987);
nor U7284 (N_7284,N_6936,N_6655);
xnor U7285 (N_7285,N_6578,N_6671);
nand U7286 (N_7286,N_6697,N_6744);
or U7287 (N_7287,N_6502,N_6650);
xnor U7288 (N_7288,N_6777,N_6884);
xnor U7289 (N_7289,N_6722,N_6866);
xor U7290 (N_7290,N_6735,N_6965);
xnor U7291 (N_7291,N_6550,N_6536);
xor U7292 (N_7292,N_6935,N_6756);
nand U7293 (N_7293,N_6696,N_6810);
nand U7294 (N_7294,N_6962,N_6752);
nor U7295 (N_7295,N_6980,N_6786);
or U7296 (N_7296,N_6627,N_6609);
nor U7297 (N_7297,N_6757,N_6777);
nor U7298 (N_7298,N_6745,N_6861);
xnor U7299 (N_7299,N_6962,N_6607);
and U7300 (N_7300,N_6512,N_6628);
nor U7301 (N_7301,N_6659,N_6618);
or U7302 (N_7302,N_6513,N_6625);
xor U7303 (N_7303,N_6715,N_6660);
xnor U7304 (N_7304,N_6539,N_6815);
nand U7305 (N_7305,N_6688,N_6598);
or U7306 (N_7306,N_6810,N_6843);
or U7307 (N_7307,N_6972,N_6899);
xor U7308 (N_7308,N_6820,N_6681);
nand U7309 (N_7309,N_6876,N_6605);
nor U7310 (N_7310,N_6563,N_6806);
or U7311 (N_7311,N_6993,N_6506);
nand U7312 (N_7312,N_6839,N_6562);
nand U7313 (N_7313,N_6989,N_6941);
and U7314 (N_7314,N_6871,N_6508);
or U7315 (N_7315,N_6846,N_6864);
and U7316 (N_7316,N_6511,N_6692);
and U7317 (N_7317,N_6718,N_6655);
nand U7318 (N_7318,N_6962,N_6771);
xor U7319 (N_7319,N_6826,N_6817);
and U7320 (N_7320,N_6844,N_6760);
and U7321 (N_7321,N_6550,N_6652);
nand U7322 (N_7322,N_6682,N_6613);
nand U7323 (N_7323,N_6971,N_6894);
nand U7324 (N_7324,N_6852,N_6692);
and U7325 (N_7325,N_6966,N_6643);
or U7326 (N_7326,N_6762,N_6973);
nand U7327 (N_7327,N_6646,N_6656);
nor U7328 (N_7328,N_6673,N_6701);
xor U7329 (N_7329,N_6977,N_6852);
or U7330 (N_7330,N_6767,N_6762);
nor U7331 (N_7331,N_6589,N_6692);
or U7332 (N_7332,N_6963,N_6664);
nand U7333 (N_7333,N_6871,N_6545);
and U7334 (N_7334,N_6814,N_6571);
xor U7335 (N_7335,N_6710,N_6530);
xnor U7336 (N_7336,N_6777,N_6523);
xnor U7337 (N_7337,N_6749,N_6878);
and U7338 (N_7338,N_6992,N_6757);
or U7339 (N_7339,N_6807,N_6519);
nand U7340 (N_7340,N_6762,N_6898);
nand U7341 (N_7341,N_6552,N_6838);
nand U7342 (N_7342,N_6955,N_6520);
or U7343 (N_7343,N_6548,N_6810);
or U7344 (N_7344,N_6942,N_6712);
xor U7345 (N_7345,N_6631,N_6531);
nor U7346 (N_7346,N_6557,N_6876);
or U7347 (N_7347,N_6907,N_6565);
nand U7348 (N_7348,N_6761,N_6705);
nor U7349 (N_7349,N_6667,N_6734);
or U7350 (N_7350,N_6569,N_6570);
xnor U7351 (N_7351,N_6666,N_6601);
or U7352 (N_7352,N_6925,N_6736);
and U7353 (N_7353,N_6528,N_6601);
or U7354 (N_7354,N_6642,N_6515);
xnor U7355 (N_7355,N_6685,N_6519);
nor U7356 (N_7356,N_6536,N_6551);
nand U7357 (N_7357,N_6893,N_6512);
nand U7358 (N_7358,N_6605,N_6775);
xor U7359 (N_7359,N_6582,N_6670);
and U7360 (N_7360,N_6946,N_6696);
nand U7361 (N_7361,N_6812,N_6817);
and U7362 (N_7362,N_6907,N_6769);
nand U7363 (N_7363,N_6809,N_6823);
nor U7364 (N_7364,N_6695,N_6760);
xnor U7365 (N_7365,N_6594,N_6757);
nand U7366 (N_7366,N_6865,N_6636);
nand U7367 (N_7367,N_6685,N_6630);
nor U7368 (N_7368,N_6688,N_6809);
nor U7369 (N_7369,N_6606,N_6568);
nor U7370 (N_7370,N_6614,N_6950);
nand U7371 (N_7371,N_6916,N_6795);
nand U7372 (N_7372,N_6508,N_6932);
and U7373 (N_7373,N_6622,N_6826);
or U7374 (N_7374,N_6838,N_6925);
xnor U7375 (N_7375,N_6792,N_6787);
xor U7376 (N_7376,N_6835,N_6602);
xor U7377 (N_7377,N_6809,N_6695);
nand U7378 (N_7378,N_6864,N_6997);
xnor U7379 (N_7379,N_6527,N_6884);
xnor U7380 (N_7380,N_6602,N_6931);
xor U7381 (N_7381,N_6670,N_6716);
or U7382 (N_7382,N_6983,N_6713);
xnor U7383 (N_7383,N_6966,N_6774);
nor U7384 (N_7384,N_6812,N_6848);
nand U7385 (N_7385,N_6611,N_6548);
nand U7386 (N_7386,N_6615,N_6729);
or U7387 (N_7387,N_6767,N_6666);
nor U7388 (N_7388,N_6814,N_6667);
and U7389 (N_7389,N_6763,N_6536);
and U7390 (N_7390,N_6845,N_6627);
or U7391 (N_7391,N_6976,N_6919);
xnor U7392 (N_7392,N_6800,N_6682);
xor U7393 (N_7393,N_6844,N_6936);
or U7394 (N_7394,N_6977,N_6571);
nand U7395 (N_7395,N_6929,N_6816);
nand U7396 (N_7396,N_6683,N_6530);
nor U7397 (N_7397,N_6764,N_6829);
nand U7398 (N_7398,N_6891,N_6833);
xnor U7399 (N_7399,N_6702,N_6905);
nor U7400 (N_7400,N_6920,N_6730);
and U7401 (N_7401,N_6819,N_6510);
xnor U7402 (N_7402,N_6606,N_6847);
and U7403 (N_7403,N_6646,N_6588);
xnor U7404 (N_7404,N_6517,N_6639);
and U7405 (N_7405,N_6912,N_6953);
or U7406 (N_7406,N_6890,N_6946);
or U7407 (N_7407,N_6797,N_6749);
xor U7408 (N_7408,N_6819,N_6701);
or U7409 (N_7409,N_6861,N_6759);
nand U7410 (N_7410,N_6984,N_6955);
or U7411 (N_7411,N_6802,N_6754);
nor U7412 (N_7412,N_6526,N_6552);
nand U7413 (N_7413,N_6709,N_6973);
nand U7414 (N_7414,N_6812,N_6970);
nand U7415 (N_7415,N_6717,N_6939);
and U7416 (N_7416,N_6889,N_6908);
xor U7417 (N_7417,N_6884,N_6790);
xor U7418 (N_7418,N_6660,N_6556);
xor U7419 (N_7419,N_6642,N_6614);
nand U7420 (N_7420,N_6536,N_6595);
and U7421 (N_7421,N_6872,N_6998);
or U7422 (N_7422,N_6780,N_6640);
xnor U7423 (N_7423,N_6919,N_6692);
and U7424 (N_7424,N_6799,N_6885);
or U7425 (N_7425,N_6670,N_6936);
nor U7426 (N_7426,N_6609,N_6726);
nand U7427 (N_7427,N_6577,N_6710);
and U7428 (N_7428,N_6936,N_6691);
nand U7429 (N_7429,N_6762,N_6983);
nor U7430 (N_7430,N_6764,N_6935);
nand U7431 (N_7431,N_6599,N_6889);
nor U7432 (N_7432,N_6674,N_6897);
xor U7433 (N_7433,N_6859,N_6805);
or U7434 (N_7434,N_6531,N_6750);
nand U7435 (N_7435,N_6962,N_6906);
and U7436 (N_7436,N_6602,N_6666);
or U7437 (N_7437,N_6545,N_6816);
nand U7438 (N_7438,N_6799,N_6841);
nor U7439 (N_7439,N_6581,N_6591);
or U7440 (N_7440,N_6803,N_6506);
and U7441 (N_7441,N_6697,N_6581);
or U7442 (N_7442,N_6575,N_6525);
or U7443 (N_7443,N_6843,N_6608);
or U7444 (N_7444,N_6771,N_6710);
or U7445 (N_7445,N_6600,N_6585);
nor U7446 (N_7446,N_6594,N_6603);
and U7447 (N_7447,N_6641,N_6787);
nor U7448 (N_7448,N_6894,N_6703);
xnor U7449 (N_7449,N_6507,N_6811);
nand U7450 (N_7450,N_6763,N_6686);
or U7451 (N_7451,N_6973,N_6735);
nand U7452 (N_7452,N_6862,N_6612);
nand U7453 (N_7453,N_6864,N_6501);
xor U7454 (N_7454,N_6915,N_6868);
and U7455 (N_7455,N_6961,N_6802);
xnor U7456 (N_7456,N_6651,N_6670);
xor U7457 (N_7457,N_6805,N_6751);
nor U7458 (N_7458,N_6769,N_6915);
nand U7459 (N_7459,N_6611,N_6609);
nand U7460 (N_7460,N_6534,N_6886);
nor U7461 (N_7461,N_6717,N_6949);
xor U7462 (N_7462,N_6936,N_6513);
and U7463 (N_7463,N_6762,N_6618);
nor U7464 (N_7464,N_6843,N_6565);
nor U7465 (N_7465,N_6693,N_6850);
nor U7466 (N_7466,N_6891,N_6972);
or U7467 (N_7467,N_6594,N_6945);
nand U7468 (N_7468,N_6522,N_6878);
xor U7469 (N_7469,N_6949,N_6796);
and U7470 (N_7470,N_6630,N_6815);
xor U7471 (N_7471,N_6741,N_6626);
nor U7472 (N_7472,N_6788,N_6797);
or U7473 (N_7473,N_6574,N_6770);
or U7474 (N_7474,N_6733,N_6886);
or U7475 (N_7475,N_6656,N_6823);
nand U7476 (N_7476,N_6917,N_6538);
nand U7477 (N_7477,N_6806,N_6891);
and U7478 (N_7478,N_6761,N_6727);
or U7479 (N_7479,N_6733,N_6576);
or U7480 (N_7480,N_6545,N_6760);
nand U7481 (N_7481,N_6838,N_6603);
or U7482 (N_7482,N_6785,N_6506);
nand U7483 (N_7483,N_6813,N_6995);
and U7484 (N_7484,N_6857,N_6745);
xor U7485 (N_7485,N_6556,N_6517);
nor U7486 (N_7486,N_6517,N_6541);
nor U7487 (N_7487,N_6534,N_6812);
nand U7488 (N_7488,N_6623,N_6662);
xnor U7489 (N_7489,N_6680,N_6594);
and U7490 (N_7490,N_6864,N_6798);
or U7491 (N_7491,N_6914,N_6850);
or U7492 (N_7492,N_6757,N_6629);
xor U7493 (N_7493,N_6935,N_6960);
or U7494 (N_7494,N_6573,N_6536);
xnor U7495 (N_7495,N_6580,N_6707);
nor U7496 (N_7496,N_6562,N_6752);
or U7497 (N_7497,N_6872,N_6659);
and U7498 (N_7498,N_6510,N_6573);
nand U7499 (N_7499,N_6519,N_6614);
xnor U7500 (N_7500,N_7435,N_7458);
or U7501 (N_7501,N_7433,N_7475);
and U7502 (N_7502,N_7485,N_7236);
xor U7503 (N_7503,N_7103,N_7360);
nor U7504 (N_7504,N_7083,N_7317);
xnor U7505 (N_7505,N_7077,N_7312);
nor U7506 (N_7506,N_7005,N_7041);
and U7507 (N_7507,N_7202,N_7182);
xnor U7508 (N_7508,N_7006,N_7470);
or U7509 (N_7509,N_7467,N_7471);
nand U7510 (N_7510,N_7140,N_7061);
xor U7511 (N_7511,N_7056,N_7385);
and U7512 (N_7512,N_7290,N_7494);
and U7513 (N_7513,N_7269,N_7265);
nor U7514 (N_7514,N_7495,N_7010);
or U7515 (N_7515,N_7141,N_7215);
or U7516 (N_7516,N_7076,N_7444);
xnor U7517 (N_7517,N_7246,N_7432);
and U7518 (N_7518,N_7107,N_7073);
and U7519 (N_7519,N_7074,N_7387);
and U7520 (N_7520,N_7047,N_7108);
or U7521 (N_7521,N_7170,N_7306);
or U7522 (N_7522,N_7313,N_7122);
xnor U7523 (N_7523,N_7008,N_7239);
xnor U7524 (N_7524,N_7328,N_7283);
or U7525 (N_7525,N_7223,N_7119);
xnor U7526 (N_7526,N_7086,N_7154);
nand U7527 (N_7527,N_7091,N_7295);
or U7528 (N_7528,N_7361,N_7120);
nor U7529 (N_7529,N_7285,N_7055);
and U7530 (N_7530,N_7138,N_7297);
nand U7531 (N_7531,N_7448,N_7075);
nor U7532 (N_7532,N_7305,N_7022);
or U7533 (N_7533,N_7151,N_7334);
nor U7534 (N_7534,N_7412,N_7162);
or U7535 (N_7535,N_7273,N_7163);
or U7536 (N_7536,N_7190,N_7418);
xor U7537 (N_7537,N_7377,N_7084);
or U7538 (N_7538,N_7474,N_7146);
or U7539 (N_7539,N_7264,N_7434);
nand U7540 (N_7540,N_7231,N_7092);
or U7541 (N_7541,N_7416,N_7326);
and U7542 (N_7542,N_7347,N_7331);
nor U7543 (N_7543,N_7123,N_7358);
nor U7544 (N_7544,N_7388,N_7220);
nor U7545 (N_7545,N_7157,N_7112);
nor U7546 (N_7546,N_7131,N_7147);
nand U7547 (N_7547,N_7052,N_7391);
and U7548 (N_7548,N_7383,N_7268);
or U7549 (N_7549,N_7025,N_7424);
nor U7550 (N_7550,N_7308,N_7071);
or U7551 (N_7551,N_7053,N_7243);
xnor U7552 (N_7552,N_7274,N_7179);
and U7553 (N_7553,N_7144,N_7482);
or U7554 (N_7554,N_7234,N_7450);
nor U7555 (N_7555,N_7004,N_7481);
and U7556 (N_7556,N_7200,N_7136);
xnor U7557 (N_7557,N_7221,N_7044);
nor U7558 (N_7558,N_7079,N_7259);
and U7559 (N_7559,N_7003,N_7406);
nor U7560 (N_7560,N_7459,N_7394);
xnor U7561 (N_7561,N_7423,N_7063);
xor U7562 (N_7562,N_7338,N_7411);
xor U7563 (N_7563,N_7457,N_7398);
or U7564 (N_7564,N_7483,N_7139);
nand U7565 (N_7565,N_7466,N_7492);
and U7566 (N_7566,N_7040,N_7105);
nor U7567 (N_7567,N_7241,N_7143);
nor U7568 (N_7568,N_7252,N_7069);
and U7569 (N_7569,N_7425,N_7263);
and U7570 (N_7570,N_7142,N_7065);
nor U7571 (N_7571,N_7451,N_7329);
xor U7572 (N_7572,N_7395,N_7250);
and U7573 (N_7573,N_7066,N_7441);
nor U7574 (N_7574,N_7177,N_7219);
xnor U7575 (N_7575,N_7137,N_7110);
and U7576 (N_7576,N_7333,N_7447);
or U7577 (N_7577,N_7303,N_7169);
xnor U7578 (N_7578,N_7206,N_7497);
and U7579 (N_7579,N_7209,N_7153);
nand U7580 (N_7580,N_7167,N_7101);
nor U7581 (N_7581,N_7051,N_7393);
or U7582 (N_7582,N_7228,N_7351);
or U7583 (N_7583,N_7419,N_7429);
nor U7584 (N_7584,N_7337,N_7472);
or U7585 (N_7585,N_7381,N_7159);
xnor U7586 (N_7586,N_7007,N_7088);
or U7587 (N_7587,N_7427,N_7426);
or U7588 (N_7588,N_7192,N_7376);
and U7589 (N_7589,N_7404,N_7204);
nor U7590 (N_7590,N_7100,N_7191);
and U7591 (N_7591,N_7292,N_7320);
nand U7592 (N_7592,N_7176,N_7185);
or U7593 (N_7593,N_7230,N_7064);
or U7594 (N_7594,N_7327,N_7184);
nand U7595 (N_7595,N_7161,N_7365);
nor U7596 (N_7596,N_7245,N_7272);
nor U7597 (N_7597,N_7363,N_7257);
and U7598 (N_7598,N_7207,N_7057);
or U7599 (N_7599,N_7054,N_7430);
and U7600 (N_7600,N_7253,N_7311);
nand U7601 (N_7601,N_7132,N_7128);
xnor U7602 (N_7602,N_7384,N_7186);
nor U7603 (N_7603,N_7362,N_7224);
and U7604 (N_7604,N_7477,N_7455);
and U7605 (N_7605,N_7310,N_7498);
and U7606 (N_7606,N_7171,N_7018);
nand U7607 (N_7607,N_7089,N_7309);
nand U7608 (N_7608,N_7415,N_7240);
and U7609 (N_7609,N_7287,N_7260);
and U7610 (N_7610,N_7049,N_7420);
and U7611 (N_7611,N_7011,N_7090);
or U7612 (N_7612,N_7254,N_7193);
and U7613 (N_7613,N_7037,N_7438);
nand U7614 (N_7614,N_7370,N_7150);
and U7615 (N_7615,N_7058,N_7405);
and U7616 (N_7616,N_7060,N_7496);
and U7617 (N_7617,N_7276,N_7133);
nor U7618 (N_7618,N_7324,N_7417);
nand U7619 (N_7619,N_7422,N_7183);
or U7620 (N_7620,N_7097,N_7158);
xor U7621 (N_7621,N_7399,N_7160);
nor U7622 (N_7622,N_7439,N_7015);
xnor U7623 (N_7623,N_7271,N_7281);
and U7624 (N_7624,N_7029,N_7201);
xor U7625 (N_7625,N_7080,N_7251);
xor U7626 (N_7626,N_7480,N_7032);
nor U7627 (N_7627,N_7321,N_7226);
xnor U7628 (N_7628,N_7210,N_7205);
nand U7629 (N_7629,N_7428,N_7031);
and U7630 (N_7630,N_7348,N_7288);
and U7631 (N_7631,N_7291,N_7289);
or U7632 (N_7632,N_7244,N_7039);
nand U7633 (N_7633,N_7478,N_7229);
xor U7634 (N_7634,N_7401,N_7227);
nor U7635 (N_7635,N_7175,N_7102);
or U7636 (N_7636,N_7284,N_7336);
nor U7637 (N_7637,N_7266,N_7197);
xor U7638 (N_7638,N_7237,N_7238);
and U7639 (N_7639,N_7408,N_7345);
xor U7640 (N_7640,N_7355,N_7111);
xnor U7641 (N_7641,N_7465,N_7493);
and U7642 (N_7642,N_7216,N_7121);
nand U7643 (N_7643,N_7410,N_7001);
nor U7644 (N_7644,N_7129,N_7208);
or U7645 (N_7645,N_7463,N_7367);
and U7646 (N_7646,N_7491,N_7035);
or U7647 (N_7647,N_7318,N_7302);
and U7648 (N_7648,N_7414,N_7106);
or U7649 (N_7649,N_7487,N_7437);
or U7650 (N_7650,N_7033,N_7402);
nor U7651 (N_7651,N_7258,N_7446);
nand U7652 (N_7652,N_7296,N_7094);
or U7653 (N_7653,N_7352,N_7235);
xor U7654 (N_7654,N_7314,N_7085);
nand U7655 (N_7655,N_7325,N_7165);
nor U7656 (N_7656,N_7270,N_7332);
nor U7657 (N_7657,N_7211,N_7490);
nor U7658 (N_7658,N_7364,N_7189);
nor U7659 (N_7659,N_7020,N_7453);
xnor U7660 (N_7660,N_7045,N_7278);
or U7661 (N_7661,N_7023,N_7330);
or U7662 (N_7662,N_7013,N_7152);
xor U7663 (N_7663,N_7248,N_7114);
and U7664 (N_7664,N_7379,N_7344);
nand U7665 (N_7665,N_7486,N_7082);
nand U7666 (N_7666,N_7300,N_7359);
nand U7667 (N_7667,N_7307,N_7315);
nand U7668 (N_7668,N_7489,N_7462);
nand U7669 (N_7669,N_7042,N_7115);
nand U7670 (N_7670,N_7127,N_7316);
nand U7671 (N_7671,N_7249,N_7194);
and U7672 (N_7672,N_7449,N_7301);
nor U7673 (N_7673,N_7421,N_7081);
or U7674 (N_7674,N_7371,N_7298);
or U7675 (N_7675,N_7323,N_7155);
xnor U7676 (N_7676,N_7027,N_7378);
nand U7677 (N_7677,N_7277,N_7072);
and U7678 (N_7678,N_7340,N_7293);
xnor U7679 (N_7679,N_7048,N_7373);
nand U7680 (N_7680,N_7164,N_7203);
nor U7681 (N_7681,N_7180,N_7294);
nand U7682 (N_7682,N_7050,N_7390);
nand U7683 (N_7683,N_7319,N_7464);
nor U7684 (N_7684,N_7440,N_7124);
nor U7685 (N_7685,N_7187,N_7479);
nor U7686 (N_7686,N_7166,N_7400);
or U7687 (N_7687,N_7099,N_7369);
nor U7688 (N_7688,N_7322,N_7341);
xor U7689 (N_7689,N_7024,N_7342);
or U7690 (N_7690,N_7034,N_7009);
and U7691 (N_7691,N_7173,N_7198);
nand U7692 (N_7692,N_7098,N_7456);
nand U7693 (N_7693,N_7346,N_7232);
xor U7694 (N_7694,N_7002,N_7012);
xnor U7695 (N_7695,N_7354,N_7174);
nor U7696 (N_7696,N_7386,N_7126);
and U7697 (N_7697,N_7409,N_7356);
xnor U7698 (N_7698,N_7116,N_7017);
or U7699 (N_7699,N_7335,N_7067);
xnor U7700 (N_7700,N_7368,N_7484);
nor U7701 (N_7701,N_7078,N_7413);
or U7702 (N_7702,N_7043,N_7380);
nor U7703 (N_7703,N_7000,N_7445);
nor U7704 (N_7704,N_7188,N_7087);
nor U7705 (N_7705,N_7460,N_7016);
xnor U7706 (N_7706,N_7436,N_7382);
nand U7707 (N_7707,N_7261,N_7178);
and U7708 (N_7708,N_7469,N_7148);
nor U7709 (N_7709,N_7499,N_7275);
and U7710 (N_7710,N_7389,N_7217);
nor U7711 (N_7711,N_7403,N_7172);
nand U7712 (N_7712,N_7113,N_7218);
nand U7713 (N_7713,N_7256,N_7130);
and U7714 (N_7714,N_7372,N_7014);
nor U7715 (N_7715,N_7070,N_7026);
or U7716 (N_7716,N_7021,N_7396);
nand U7717 (N_7717,N_7019,N_7195);
or U7718 (N_7718,N_7299,N_7267);
or U7719 (N_7719,N_7339,N_7062);
or U7720 (N_7720,N_7353,N_7028);
xnor U7721 (N_7721,N_7443,N_7214);
nor U7722 (N_7722,N_7233,N_7242);
and U7723 (N_7723,N_7225,N_7262);
or U7724 (N_7724,N_7431,N_7118);
or U7725 (N_7725,N_7442,N_7461);
nor U7726 (N_7726,N_7096,N_7279);
or U7727 (N_7727,N_7304,N_7036);
xor U7728 (N_7728,N_7374,N_7488);
nor U7729 (N_7729,N_7059,N_7104);
and U7730 (N_7730,N_7375,N_7135);
or U7731 (N_7731,N_7117,N_7038);
nand U7732 (N_7732,N_7473,N_7397);
xnor U7733 (N_7733,N_7068,N_7452);
nand U7734 (N_7734,N_7392,N_7282);
xor U7735 (N_7735,N_7286,N_7468);
nor U7736 (N_7736,N_7212,N_7109);
or U7737 (N_7737,N_7030,N_7454);
xor U7738 (N_7738,N_7357,N_7199);
nor U7739 (N_7739,N_7349,N_7247);
nor U7740 (N_7740,N_7350,N_7213);
xor U7741 (N_7741,N_7046,N_7168);
and U7742 (N_7742,N_7145,N_7125);
xor U7743 (N_7743,N_7222,N_7366);
nand U7744 (N_7744,N_7343,N_7156);
or U7745 (N_7745,N_7095,N_7181);
nor U7746 (N_7746,N_7149,N_7196);
xnor U7747 (N_7747,N_7476,N_7255);
or U7748 (N_7748,N_7134,N_7407);
nor U7749 (N_7749,N_7093,N_7280);
nand U7750 (N_7750,N_7155,N_7483);
and U7751 (N_7751,N_7348,N_7392);
nor U7752 (N_7752,N_7265,N_7231);
xor U7753 (N_7753,N_7308,N_7297);
or U7754 (N_7754,N_7230,N_7394);
or U7755 (N_7755,N_7152,N_7139);
or U7756 (N_7756,N_7321,N_7291);
xor U7757 (N_7757,N_7074,N_7475);
nand U7758 (N_7758,N_7297,N_7210);
and U7759 (N_7759,N_7043,N_7069);
nor U7760 (N_7760,N_7111,N_7496);
xor U7761 (N_7761,N_7090,N_7046);
nand U7762 (N_7762,N_7318,N_7415);
nor U7763 (N_7763,N_7408,N_7020);
xnor U7764 (N_7764,N_7344,N_7002);
xnor U7765 (N_7765,N_7276,N_7412);
or U7766 (N_7766,N_7421,N_7165);
or U7767 (N_7767,N_7036,N_7134);
and U7768 (N_7768,N_7251,N_7053);
and U7769 (N_7769,N_7292,N_7442);
and U7770 (N_7770,N_7377,N_7472);
nand U7771 (N_7771,N_7448,N_7253);
nand U7772 (N_7772,N_7403,N_7374);
xnor U7773 (N_7773,N_7438,N_7128);
nor U7774 (N_7774,N_7256,N_7276);
or U7775 (N_7775,N_7178,N_7205);
xnor U7776 (N_7776,N_7118,N_7418);
nor U7777 (N_7777,N_7412,N_7482);
xnor U7778 (N_7778,N_7359,N_7272);
nand U7779 (N_7779,N_7261,N_7194);
nand U7780 (N_7780,N_7044,N_7226);
nor U7781 (N_7781,N_7234,N_7118);
or U7782 (N_7782,N_7463,N_7302);
and U7783 (N_7783,N_7174,N_7303);
or U7784 (N_7784,N_7347,N_7249);
nand U7785 (N_7785,N_7469,N_7437);
or U7786 (N_7786,N_7067,N_7090);
nand U7787 (N_7787,N_7394,N_7355);
or U7788 (N_7788,N_7467,N_7027);
and U7789 (N_7789,N_7113,N_7150);
or U7790 (N_7790,N_7413,N_7498);
nor U7791 (N_7791,N_7133,N_7221);
nor U7792 (N_7792,N_7050,N_7430);
xnor U7793 (N_7793,N_7228,N_7235);
nor U7794 (N_7794,N_7222,N_7016);
nor U7795 (N_7795,N_7207,N_7092);
nand U7796 (N_7796,N_7400,N_7266);
nand U7797 (N_7797,N_7055,N_7201);
or U7798 (N_7798,N_7128,N_7023);
and U7799 (N_7799,N_7238,N_7049);
nand U7800 (N_7800,N_7236,N_7250);
or U7801 (N_7801,N_7174,N_7489);
and U7802 (N_7802,N_7153,N_7331);
nor U7803 (N_7803,N_7303,N_7395);
xnor U7804 (N_7804,N_7339,N_7044);
nand U7805 (N_7805,N_7233,N_7036);
and U7806 (N_7806,N_7447,N_7248);
and U7807 (N_7807,N_7440,N_7141);
nand U7808 (N_7808,N_7235,N_7354);
and U7809 (N_7809,N_7358,N_7125);
xor U7810 (N_7810,N_7217,N_7019);
or U7811 (N_7811,N_7235,N_7173);
nand U7812 (N_7812,N_7260,N_7325);
or U7813 (N_7813,N_7374,N_7215);
and U7814 (N_7814,N_7436,N_7110);
or U7815 (N_7815,N_7294,N_7032);
or U7816 (N_7816,N_7258,N_7401);
nor U7817 (N_7817,N_7346,N_7225);
nor U7818 (N_7818,N_7138,N_7459);
and U7819 (N_7819,N_7496,N_7383);
and U7820 (N_7820,N_7027,N_7214);
nor U7821 (N_7821,N_7121,N_7132);
nor U7822 (N_7822,N_7035,N_7029);
nor U7823 (N_7823,N_7073,N_7286);
and U7824 (N_7824,N_7253,N_7268);
nor U7825 (N_7825,N_7324,N_7234);
xor U7826 (N_7826,N_7481,N_7027);
xnor U7827 (N_7827,N_7002,N_7255);
nor U7828 (N_7828,N_7420,N_7392);
and U7829 (N_7829,N_7449,N_7197);
xnor U7830 (N_7830,N_7184,N_7112);
or U7831 (N_7831,N_7306,N_7119);
and U7832 (N_7832,N_7044,N_7099);
and U7833 (N_7833,N_7089,N_7013);
xor U7834 (N_7834,N_7328,N_7116);
or U7835 (N_7835,N_7171,N_7265);
nand U7836 (N_7836,N_7447,N_7249);
nand U7837 (N_7837,N_7090,N_7120);
or U7838 (N_7838,N_7460,N_7449);
xnor U7839 (N_7839,N_7027,N_7302);
xor U7840 (N_7840,N_7342,N_7130);
or U7841 (N_7841,N_7424,N_7093);
and U7842 (N_7842,N_7256,N_7071);
nor U7843 (N_7843,N_7349,N_7375);
nor U7844 (N_7844,N_7196,N_7247);
and U7845 (N_7845,N_7217,N_7189);
nand U7846 (N_7846,N_7234,N_7030);
nor U7847 (N_7847,N_7451,N_7301);
nor U7848 (N_7848,N_7411,N_7223);
nor U7849 (N_7849,N_7079,N_7189);
nand U7850 (N_7850,N_7197,N_7270);
or U7851 (N_7851,N_7408,N_7470);
nor U7852 (N_7852,N_7443,N_7335);
nor U7853 (N_7853,N_7172,N_7297);
nor U7854 (N_7854,N_7203,N_7049);
nor U7855 (N_7855,N_7074,N_7117);
nand U7856 (N_7856,N_7097,N_7291);
xnor U7857 (N_7857,N_7420,N_7482);
xnor U7858 (N_7858,N_7439,N_7449);
or U7859 (N_7859,N_7454,N_7292);
and U7860 (N_7860,N_7097,N_7309);
and U7861 (N_7861,N_7200,N_7382);
or U7862 (N_7862,N_7119,N_7380);
xnor U7863 (N_7863,N_7049,N_7164);
xor U7864 (N_7864,N_7480,N_7401);
or U7865 (N_7865,N_7274,N_7029);
and U7866 (N_7866,N_7343,N_7426);
xor U7867 (N_7867,N_7136,N_7485);
and U7868 (N_7868,N_7086,N_7311);
nand U7869 (N_7869,N_7292,N_7036);
nand U7870 (N_7870,N_7038,N_7015);
nand U7871 (N_7871,N_7322,N_7298);
xnor U7872 (N_7872,N_7434,N_7208);
or U7873 (N_7873,N_7057,N_7022);
and U7874 (N_7874,N_7182,N_7446);
and U7875 (N_7875,N_7010,N_7124);
or U7876 (N_7876,N_7099,N_7319);
nor U7877 (N_7877,N_7152,N_7461);
xnor U7878 (N_7878,N_7442,N_7473);
or U7879 (N_7879,N_7050,N_7112);
or U7880 (N_7880,N_7070,N_7262);
nand U7881 (N_7881,N_7291,N_7454);
nand U7882 (N_7882,N_7437,N_7267);
nor U7883 (N_7883,N_7138,N_7109);
or U7884 (N_7884,N_7493,N_7453);
xnor U7885 (N_7885,N_7133,N_7021);
or U7886 (N_7886,N_7405,N_7119);
and U7887 (N_7887,N_7313,N_7245);
nor U7888 (N_7888,N_7311,N_7413);
xor U7889 (N_7889,N_7326,N_7111);
and U7890 (N_7890,N_7202,N_7012);
nor U7891 (N_7891,N_7353,N_7366);
or U7892 (N_7892,N_7083,N_7017);
or U7893 (N_7893,N_7350,N_7128);
and U7894 (N_7894,N_7059,N_7298);
xnor U7895 (N_7895,N_7411,N_7126);
xor U7896 (N_7896,N_7190,N_7120);
xnor U7897 (N_7897,N_7008,N_7216);
and U7898 (N_7898,N_7208,N_7448);
xnor U7899 (N_7899,N_7382,N_7172);
and U7900 (N_7900,N_7176,N_7129);
nor U7901 (N_7901,N_7002,N_7053);
nand U7902 (N_7902,N_7261,N_7143);
xnor U7903 (N_7903,N_7445,N_7324);
nand U7904 (N_7904,N_7261,N_7394);
or U7905 (N_7905,N_7222,N_7300);
xor U7906 (N_7906,N_7344,N_7289);
nand U7907 (N_7907,N_7445,N_7267);
or U7908 (N_7908,N_7252,N_7219);
nor U7909 (N_7909,N_7307,N_7369);
xnor U7910 (N_7910,N_7040,N_7166);
and U7911 (N_7911,N_7259,N_7295);
and U7912 (N_7912,N_7096,N_7423);
and U7913 (N_7913,N_7299,N_7251);
or U7914 (N_7914,N_7466,N_7448);
or U7915 (N_7915,N_7393,N_7116);
nor U7916 (N_7916,N_7273,N_7294);
xor U7917 (N_7917,N_7268,N_7044);
xnor U7918 (N_7918,N_7111,N_7327);
and U7919 (N_7919,N_7371,N_7018);
nand U7920 (N_7920,N_7412,N_7093);
or U7921 (N_7921,N_7490,N_7158);
or U7922 (N_7922,N_7084,N_7173);
nand U7923 (N_7923,N_7037,N_7433);
nor U7924 (N_7924,N_7140,N_7464);
xor U7925 (N_7925,N_7344,N_7034);
nor U7926 (N_7926,N_7331,N_7215);
xnor U7927 (N_7927,N_7347,N_7276);
and U7928 (N_7928,N_7145,N_7011);
nor U7929 (N_7929,N_7434,N_7407);
nand U7930 (N_7930,N_7414,N_7013);
nand U7931 (N_7931,N_7084,N_7290);
xnor U7932 (N_7932,N_7034,N_7245);
and U7933 (N_7933,N_7266,N_7183);
xnor U7934 (N_7934,N_7324,N_7120);
or U7935 (N_7935,N_7425,N_7366);
and U7936 (N_7936,N_7392,N_7215);
nand U7937 (N_7937,N_7056,N_7415);
nor U7938 (N_7938,N_7359,N_7094);
and U7939 (N_7939,N_7418,N_7357);
nor U7940 (N_7940,N_7221,N_7258);
nor U7941 (N_7941,N_7390,N_7378);
nor U7942 (N_7942,N_7289,N_7085);
and U7943 (N_7943,N_7022,N_7026);
or U7944 (N_7944,N_7067,N_7320);
nand U7945 (N_7945,N_7157,N_7252);
nor U7946 (N_7946,N_7329,N_7341);
xor U7947 (N_7947,N_7079,N_7367);
or U7948 (N_7948,N_7214,N_7139);
or U7949 (N_7949,N_7230,N_7476);
and U7950 (N_7950,N_7205,N_7189);
and U7951 (N_7951,N_7102,N_7459);
or U7952 (N_7952,N_7254,N_7200);
or U7953 (N_7953,N_7107,N_7194);
and U7954 (N_7954,N_7003,N_7082);
or U7955 (N_7955,N_7494,N_7278);
xor U7956 (N_7956,N_7029,N_7087);
nand U7957 (N_7957,N_7374,N_7460);
nand U7958 (N_7958,N_7024,N_7499);
or U7959 (N_7959,N_7256,N_7264);
or U7960 (N_7960,N_7059,N_7478);
xor U7961 (N_7961,N_7193,N_7409);
nand U7962 (N_7962,N_7479,N_7256);
xor U7963 (N_7963,N_7490,N_7331);
and U7964 (N_7964,N_7087,N_7003);
or U7965 (N_7965,N_7056,N_7085);
xnor U7966 (N_7966,N_7197,N_7373);
nand U7967 (N_7967,N_7219,N_7474);
or U7968 (N_7968,N_7458,N_7069);
nand U7969 (N_7969,N_7133,N_7033);
nor U7970 (N_7970,N_7476,N_7416);
xnor U7971 (N_7971,N_7124,N_7021);
nand U7972 (N_7972,N_7435,N_7159);
and U7973 (N_7973,N_7133,N_7107);
nand U7974 (N_7974,N_7212,N_7488);
nor U7975 (N_7975,N_7204,N_7322);
or U7976 (N_7976,N_7141,N_7303);
nor U7977 (N_7977,N_7264,N_7488);
xor U7978 (N_7978,N_7231,N_7175);
xor U7979 (N_7979,N_7181,N_7076);
xnor U7980 (N_7980,N_7356,N_7411);
xnor U7981 (N_7981,N_7409,N_7381);
or U7982 (N_7982,N_7061,N_7004);
xnor U7983 (N_7983,N_7352,N_7186);
nor U7984 (N_7984,N_7162,N_7013);
xnor U7985 (N_7985,N_7137,N_7010);
nand U7986 (N_7986,N_7251,N_7288);
xor U7987 (N_7987,N_7375,N_7120);
nand U7988 (N_7988,N_7015,N_7114);
or U7989 (N_7989,N_7086,N_7496);
xnor U7990 (N_7990,N_7342,N_7033);
nand U7991 (N_7991,N_7162,N_7433);
nand U7992 (N_7992,N_7180,N_7343);
and U7993 (N_7993,N_7208,N_7257);
nor U7994 (N_7994,N_7497,N_7027);
or U7995 (N_7995,N_7261,N_7390);
and U7996 (N_7996,N_7137,N_7228);
xnor U7997 (N_7997,N_7333,N_7224);
nor U7998 (N_7998,N_7064,N_7147);
or U7999 (N_7999,N_7147,N_7412);
or U8000 (N_8000,N_7555,N_7640);
or U8001 (N_8001,N_7914,N_7565);
xnor U8002 (N_8002,N_7983,N_7604);
and U8003 (N_8003,N_7629,N_7705);
xor U8004 (N_8004,N_7857,N_7598);
or U8005 (N_8005,N_7815,N_7680);
or U8006 (N_8006,N_7932,N_7899);
nor U8007 (N_8007,N_7751,N_7874);
nand U8008 (N_8008,N_7792,N_7928);
nor U8009 (N_8009,N_7600,N_7666);
or U8010 (N_8010,N_7509,N_7926);
nand U8011 (N_8011,N_7922,N_7829);
and U8012 (N_8012,N_7872,N_7906);
xnor U8013 (N_8013,N_7525,N_7596);
nor U8014 (N_8014,N_7725,N_7930);
nand U8015 (N_8015,N_7779,N_7553);
nand U8016 (N_8016,N_7668,N_7551);
nand U8017 (N_8017,N_7685,N_7805);
or U8018 (N_8018,N_7891,N_7682);
xor U8019 (N_8019,N_7801,N_7963);
xnor U8020 (N_8020,N_7772,N_7839);
and U8021 (N_8021,N_7691,N_7788);
nor U8022 (N_8022,N_7654,N_7749);
xor U8023 (N_8023,N_7726,N_7670);
or U8024 (N_8024,N_7511,N_7534);
nand U8025 (N_8025,N_7918,N_7923);
nor U8026 (N_8026,N_7790,N_7608);
nand U8027 (N_8027,N_7869,N_7804);
xnor U8028 (N_8028,N_7811,N_7739);
nor U8029 (N_8029,N_7690,N_7576);
nand U8030 (N_8030,N_7968,N_7686);
nor U8031 (N_8031,N_7556,N_7789);
nor U8032 (N_8032,N_7521,N_7628);
nor U8033 (N_8033,N_7893,N_7871);
nand U8034 (N_8034,N_7768,N_7527);
nand U8035 (N_8035,N_7975,N_7646);
or U8036 (N_8036,N_7618,N_7684);
nand U8037 (N_8037,N_7920,N_7712);
or U8038 (N_8038,N_7929,N_7898);
nor U8039 (N_8039,N_7830,N_7692);
or U8040 (N_8040,N_7866,N_7538);
nand U8041 (N_8041,N_7715,N_7585);
or U8042 (N_8042,N_7744,N_7663);
or U8043 (N_8043,N_7603,N_7853);
and U8044 (N_8044,N_7631,N_7522);
and U8045 (N_8045,N_7753,N_7840);
nand U8046 (N_8046,N_7573,N_7526);
xor U8047 (N_8047,N_7658,N_7540);
xnor U8048 (N_8048,N_7901,N_7954);
xor U8049 (N_8049,N_7695,N_7863);
and U8050 (N_8050,N_7700,N_7735);
nor U8051 (N_8051,N_7703,N_7516);
or U8052 (N_8052,N_7994,N_7737);
nor U8053 (N_8053,N_7641,N_7601);
nand U8054 (N_8054,N_7611,N_7591);
nand U8055 (N_8055,N_7738,N_7773);
nor U8056 (N_8056,N_7993,N_7616);
and U8057 (N_8057,N_7546,N_7997);
xnor U8058 (N_8058,N_7802,N_7675);
and U8059 (N_8059,N_7961,N_7619);
or U8060 (N_8060,N_7762,N_7634);
or U8061 (N_8061,N_7674,N_7612);
and U8062 (N_8062,N_7580,N_7701);
nor U8063 (N_8063,N_7816,N_7819);
or U8064 (N_8064,N_7575,N_7979);
xor U8065 (N_8065,N_7550,N_7605);
or U8066 (N_8066,N_7902,N_7777);
xnor U8067 (N_8067,N_7748,N_7613);
nor U8068 (N_8068,N_7841,N_7890);
nand U8069 (N_8069,N_7959,N_7520);
and U8070 (N_8070,N_7873,N_7820);
nand U8071 (N_8071,N_7951,N_7708);
xnor U8072 (N_8072,N_7623,N_7536);
nand U8073 (N_8073,N_7859,N_7767);
xnor U8074 (N_8074,N_7594,N_7564);
or U8075 (N_8075,N_7864,N_7867);
and U8076 (N_8076,N_7592,N_7718);
nor U8077 (N_8077,N_7814,N_7986);
nor U8078 (N_8078,N_7676,N_7568);
nor U8079 (N_8079,N_7637,N_7787);
nand U8080 (N_8080,N_7894,N_7657);
nand U8081 (N_8081,N_7810,N_7630);
xor U8082 (N_8082,N_7761,N_7545);
nand U8083 (N_8083,N_7948,N_7949);
and U8084 (N_8084,N_7661,N_7966);
nand U8085 (N_8085,N_7957,N_7955);
nand U8086 (N_8086,N_7793,N_7848);
nand U8087 (N_8087,N_7943,N_7584);
nor U8088 (N_8088,N_7702,N_7984);
xnor U8089 (N_8089,N_7721,N_7639);
nor U8090 (N_8090,N_7723,N_7729);
and U8091 (N_8091,N_7704,N_7885);
or U8092 (N_8092,N_7647,N_7660);
nand U8093 (N_8093,N_7964,N_7724);
nor U8094 (N_8094,N_7517,N_7913);
xor U8095 (N_8095,N_7579,N_7655);
xnor U8096 (N_8096,N_7650,N_7507);
nand U8097 (N_8097,N_7581,N_7818);
xnor U8098 (N_8098,N_7512,N_7652);
or U8099 (N_8099,N_7952,N_7991);
nand U8100 (N_8100,N_7888,N_7500);
xnor U8101 (N_8101,N_7625,N_7621);
and U8102 (N_8102,N_7557,N_7754);
or U8103 (N_8103,N_7826,N_7925);
xor U8104 (N_8104,N_7852,N_7542);
and U8105 (N_8105,N_7548,N_7706);
nor U8106 (N_8106,N_7659,N_7998);
and U8107 (N_8107,N_7941,N_7931);
xor U8108 (N_8108,N_7778,N_7907);
or U8109 (N_8109,N_7904,N_7599);
and U8110 (N_8110,N_7638,N_7759);
and U8111 (N_8111,N_7671,N_7850);
nor U8112 (N_8112,N_7664,N_7862);
xnor U8113 (N_8113,N_7882,N_7510);
and U8114 (N_8114,N_7687,N_7523);
xor U8115 (N_8115,N_7989,N_7844);
nand U8116 (N_8116,N_7795,N_7956);
and U8117 (N_8117,N_7709,N_7544);
nand U8118 (N_8118,N_7742,N_7965);
xor U8119 (N_8119,N_7981,N_7770);
xnor U8120 (N_8120,N_7549,N_7547);
or U8121 (N_8121,N_7552,N_7648);
nor U8122 (N_8122,N_7689,N_7518);
nor U8123 (N_8123,N_7558,N_7876);
nor U8124 (N_8124,N_7653,N_7563);
or U8125 (N_8125,N_7799,N_7996);
or U8126 (N_8126,N_7933,N_7973);
and U8127 (N_8127,N_7745,N_7969);
xnor U8128 (N_8128,N_7821,N_7911);
nor U8129 (N_8129,N_7627,N_7622);
xor U8130 (N_8130,N_7935,N_7617);
or U8131 (N_8131,N_7988,N_7917);
or U8132 (N_8132,N_7900,N_7614);
nand U8133 (N_8133,N_7713,N_7823);
nor U8134 (N_8134,N_7764,N_7946);
and U8135 (N_8135,N_7743,N_7919);
and U8136 (N_8136,N_7730,N_7797);
xor U8137 (N_8137,N_7662,N_7942);
or U8138 (N_8138,N_7570,N_7828);
or U8139 (N_8139,N_7645,N_7774);
xor U8140 (N_8140,N_7688,N_7578);
xnor U8141 (N_8141,N_7602,N_7566);
and U8142 (N_8142,N_7992,N_7677);
xnor U8143 (N_8143,N_7758,N_7889);
and U8144 (N_8144,N_7877,N_7953);
and U8145 (N_8145,N_7752,N_7987);
xnor U8146 (N_8146,N_7635,N_7615);
nor U8147 (N_8147,N_7832,N_7858);
xor U8148 (N_8148,N_7875,N_7824);
nor U8149 (N_8149,N_7962,N_7590);
nand U8150 (N_8150,N_7903,N_7947);
nand U8151 (N_8151,N_7528,N_7642);
xor U8152 (N_8152,N_7530,N_7972);
and U8153 (N_8153,N_7846,N_7843);
or U8154 (N_8154,N_7967,N_7887);
or U8155 (N_8155,N_7970,N_7524);
nor U8156 (N_8156,N_7781,N_7560);
nor U8157 (N_8157,N_7978,N_7974);
nand U8158 (N_8158,N_7733,N_7559);
or U8159 (N_8159,N_7583,N_7927);
nand U8160 (N_8160,N_7806,N_7976);
nand U8161 (N_8161,N_7643,N_7531);
and U8162 (N_8162,N_7697,N_7574);
nor U8163 (N_8163,N_7683,N_7897);
and U8164 (N_8164,N_7755,N_7880);
xnor U8165 (N_8165,N_7593,N_7980);
nand U8166 (N_8166,N_7982,N_7939);
nand U8167 (N_8167,N_7694,N_7950);
xnor U8168 (N_8168,N_7838,N_7699);
and U8169 (N_8169,N_7609,N_7543);
nand U8170 (N_8170,N_7842,N_7910);
nand U8171 (N_8171,N_7934,N_7572);
and U8172 (N_8172,N_7589,N_7698);
xnor U8173 (N_8173,N_7776,N_7571);
nand U8174 (N_8174,N_7732,N_7765);
nand U8175 (N_8175,N_7827,N_7856);
and U8176 (N_8176,N_7669,N_7763);
nand U8177 (N_8177,N_7539,N_7999);
nor U8178 (N_8178,N_7514,N_7855);
nor U8179 (N_8179,N_7515,N_7936);
and U8180 (N_8180,N_7990,N_7865);
or U8181 (N_8181,N_7915,N_7716);
and U8182 (N_8182,N_7958,N_7791);
nor U8183 (N_8183,N_7825,N_7597);
or U8184 (N_8184,N_7854,N_7722);
or U8185 (N_8185,N_7567,N_7720);
nand U8186 (N_8186,N_7587,N_7562);
nand U8187 (N_8187,N_7711,N_7971);
nand U8188 (N_8188,N_7532,N_7817);
nand U8189 (N_8189,N_7995,N_7879);
nor U8190 (N_8190,N_7569,N_7938);
nor U8191 (N_8191,N_7785,N_7636);
xnor U8192 (N_8192,N_7505,N_7937);
nand U8193 (N_8193,N_7837,N_7696);
and U8194 (N_8194,N_7734,N_7836);
xor U8195 (N_8195,N_7561,N_7736);
or U8196 (N_8196,N_7586,N_7620);
xnor U8197 (N_8197,N_7588,N_7577);
or U8198 (N_8198,N_7747,N_7710);
or U8199 (N_8199,N_7681,N_7665);
nor U8200 (N_8200,N_7633,N_7529);
nand U8201 (N_8201,N_7746,N_7878);
and U8202 (N_8202,N_7554,N_7798);
nand U8203 (N_8203,N_7740,N_7760);
nand U8204 (N_8204,N_7656,N_7921);
xor U8205 (N_8205,N_7667,N_7784);
xor U8206 (N_8206,N_7851,N_7606);
nand U8207 (N_8207,N_7860,N_7624);
nor U8208 (N_8208,N_7741,N_7513);
or U8209 (N_8209,N_7908,N_7728);
and U8210 (N_8210,N_7808,N_7868);
xor U8211 (N_8211,N_7833,N_7813);
and U8212 (N_8212,N_7771,N_7535);
nor U8213 (N_8213,N_7892,N_7831);
or U8214 (N_8214,N_7632,N_7673);
nor U8215 (N_8215,N_7506,N_7834);
xnor U8216 (N_8216,N_7541,N_7780);
nand U8217 (N_8217,N_7756,N_7812);
or U8218 (N_8218,N_7766,N_7884);
nor U8219 (N_8219,N_7835,N_7582);
and U8220 (N_8220,N_7626,N_7502);
and U8221 (N_8221,N_7508,N_7944);
or U8222 (N_8222,N_7727,N_7503);
or U8223 (N_8223,N_7803,N_7985);
xnor U8224 (N_8224,N_7960,N_7678);
xor U8225 (N_8225,N_7644,N_7809);
nor U8226 (N_8226,N_7881,N_7595);
nand U8227 (N_8227,N_7651,N_7533);
nor U8228 (N_8228,N_7800,N_7610);
nor U8229 (N_8229,N_7757,N_7945);
and U8230 (N_8230,N_7916,N_7794);
and U8231 (N_8231,N_7672,N_7607);
or U8232 (N_8232,N_7886,N_7649);
nor U8233 (N_8233,N_7717,N_7786);
nand U8234 (N_8234,N_7693,N_7775);
nor U8235 (N_8235,N_7896,N_7861);
and U8236 (N_8236,N_7679,N_7750);
nor U8237 (N_8237,N_7782,N_7847);
nor U8238 (N_8238,N_7849,N_7822);
and U8239 (N_8239,N_7870,N_7769);
nand U8240 (N_8240,N_7714,N_7504);
xnor U8241 (N_8241,N_7707,N_7977);
and U8242 (N_8242,N_7783,N_7719);
nand U8243 (N_8243,N_7912,N_7537);
xnor U8244 (N_8244,N_7501,N_7796);
and U8245 (N_8245,N_7905,N_7909);
or U8246 (N_8246,N_7883,N_7807);
nor U8247 (N_8247,N_7924,N_7731);
nand U8248 (N_8248,N_7845,N_7519);
nand U8249 (N_8249,N_7895,N_7940);
nor U8250 (N_8250,N_7638,N_7874);
xor U8251 (N_8251,N_7692,N_7651);
xor U8252 (N_8252,N_7847,N_7548);
nor U8253 (N_8253,N_7781,N_7995);
nor U8254 (N_8254,N_7840,N_7919);
nand U8255 (N_8255,N_7722,N_7857);
xor U8256 (N_8256,N_7571,N_7959);
or U8257 (N_8257,N_7971,N_7530);
or U8258 (N_8258,N_7557,N_7678);
or U8259 (N_8259,N_7799,N_7703);
and U8260 (N_8260,N_7752,N_7622);
or U8261 (N_8261,N_7715,N_7717);
or U8262 (N_8262,N_7752,N_7662);
nor U8263 (N_8263,N_7651,N_7795);
xor U8264 (N_8264,N_7856,N_7997);
xor U8265 (N_8265,N_7623,N_7835);
xor U8266 (N_8266,N_7765,N_7719);
or U8267 (N_8267,N_7779,N_7901);
and U8268 (N_8268,N_7669,N_7912);
and U8269 (N_8269,N_7614,N_7662);
and U8270 (N_8270,N_7655,N_7558);
nor U8271 (N_8271,N_7515,N_7728);
xor U8272 (N_8272,N_7642,N_7953);
nor U8273 (N_8273,N_7569,N_7548);
or U8274 (N_8274,N_7718,N_7793);
or U8275 (N_8275,N_7720,N_7738);
and U8276 (N_8276,N_7872,N_7814);
nor U8277 (N_8277,N_7688,N_7531);
and U8278 (N_8278,N_7974,N_7849);
nand U8279 (N_8279,N_7715,N_7687);
or U8280 (N_8280,N_7940,N_7739);
nand U8281 (N_8281,N_7921,N_7841);
and U8282 (N_8282,N_7876,N_7674);
or U8283 (N_8283,N_7927,N_7713);
or U8284 (N_8284,N_7621,N_7688);
nor U8285 (N_8285,N_7830,N_7696);
nor U8286 (N_8286,N_7898,N_7588);
xnor U8287 (N_8287,N_7897,N_7655);
nor U8288 (N_8288,N_7879,N_7515);
nor U8289 (N_8289,N_7945,N_7983);
nand U8290 (N_8290,N_7618,N_7503);
or U8291 (N_8291,N_7685,N_7725);
nand U8292 (N_8292,N_7731,N_7861);
nand U8293 (N_8293,N_7826,N_7782);
xor U8294 (N_8294,N_7505,N_7645);
or U8295 (N_8295,N_7743,N_7640);
xor U8296 (N_8296,N_7544,N_7796);
xor U8297 (N_8297,N_7538,N_7615);
and U8298 (N_8298,N_7522,N_7750);
nand U8299 (N_8299,N_7822,N_7712);
nand U8300 (N_8300,N_7713,N_7611);
and U8301 (N_8301,N_7609,N_7556);
or U8302 (N_8302,N_7724,N_7925);
xor U8303 (N_8303,N_7811,N_7921);
xnor U8304 (N_8304,N_7859,N_7898);
and U8305 (N_8305,N_7638,N_7861);
or U8306 (N_8306,N_7736,N_7946);
and U8307 (N_8307,N_7993,N_7819);
nand U8308 (N_8308,N_7872,N_7593);
or U8309 (N_8309,N_7790,N_7981);
nand U8310 (N_8310,N_7707,N_7646);
nor U8311 (N_8311,N_7807,N_7726);
xor U8312 (N_8312,N_7787,N_7736);
nand U8313 (N_8313,N_7671,N_7635);
xor U8314 (N_8314,N_7603,N_7667);
nand U8315 (N_8315,N_7890,N_7599);
and U8316 (N_8316,N_7518,N_7536);
and U8317 (N_8317,N_7905,N_7872);
nand U8318 (N_8318,N_7522,N_7670);
nor U8319 (N_8319,N_7895,N_7702);
nor U8320 (N_8320,N_7666,N_7642);
and U8321 (N_8321,N_7625,N_7506);
or U8322 (N_8322,N_7837,N_7612);
xor U8323 (N_8323,N_7681,N_7782);
nor U8324 (N_8324,N_7779,N_7846);
nand U8325 (N_8325,N_7733,N_7942);
or U8326 (N_8326,N_7810,N_7876);
nand U8327 (N_8327,N_7783,N_7710);
nor U8328 (N_8328,N_7793,N_7541);
nor U8329 (N_8329,N_7663,N_7612);
or U8330 (N_8330,N_7630,N_7981);
or U8331 (N_8331,N_7900,N_7689);
nor U8332 (N_8332,N_7661,N_7833);
xor U8333 (N_8333,N_7630,N_7962);
nand U8334 (N_8334,N_7750,N_7566);
xnor U8335 (N_8335,N_7591,N_7626);
nor U8336 (N_8336,N_7970,N_7849);
and U8337 (N_8337,N_7949,N_7638);
and U8338 (N_8338,N_7542,N_7711);
nand U8339 (N_8339,N_7845,N_7672);
xor U8340 (N_8340,N_7897,N_7579);
nand U8341 (N_8341,N_7662,N_7611);
nand U8342 (N_8342,N_7904,N_7865);
nor U8343 (N_8343,N_7926,N_7991);
nand U8344 (N_8344,N_7836,N_7993);
nor U8345 (N_8345,N_7960,N_7735);
nand U8346 (N_8346,N_7599,N_7619);
and U8347 (N_8347,N_7735,N_7929);
and U8348 (N_8348,N_7941,N_7629);
or U8349 (N_8349,N_7808,N_7842);
and U8350 (N_8350,N_7558,N_7704);
nand U8351 (N_8351,N_7571,N_7716);
and U8352 (N_8352,N_7628,N_7738);
and U8353 (N_8353,N_7795,N_7819);
or U8354 (N_8354,N_7838,N_7591);
and U8355 (N_8355,N_7618,N_7914);
nand U8356 (N_8356,N_7506,N_7940);
nor U8357 (N_8357,N_7528,N_7525);
or U8358 (N_8358,N_7757,N_7903);
and U8359 (N_8359,N_7613,N_7921);
nor U8360 (N_8360,N_7983,N_7659);
nand U8361 (N_8361,N_7633,N_7763);
or U8362 (N_8362,N_7979,N_7962);
or U8363 (N_8363,N_7617,N_7956);
nor U8364 (N_8364,N_7681,N_7857);
or U8365 (N_8365,N_7906,N_7508);
nor U8366 (N_8366,N_7900,N_7725);
or U8367 (N_8367,N_7548,N_7583);
xor U8368 (N_8368,N_7534,N_7843);
xnor U8369 (N_8369,N_7597,N_7922);
xnor U8370 (N_8370,N_7965,N_7903);
nand U8371 (N_8371,N_7995,N_7958);
and U8372 (N_8372,N_7821,N_7897);
and U8373 (N_8373,N_7884,N_7831);
and U8374 (N_8374,N_7659,N_7788);
and U8375 (N_8375,N_7656,N_7545);
or U8376 (N_8376,N_7515,N_7670);
nand U8377 (N_8377,N_7674,N_7607);
nand U8378 (N_8378,N_7826,N_7749);
and U8379 (N_8379,N_7601,N_7755);
and U8380 (N_8380,N_7538,N_7763);
xnor U8381 (N_8381,N_7965,N_7805);
and U8382 (N_8382,N_7538,N_7852);
nand U8383 (N_8383,N_7834,N_7681);
nand U8384 (N_8384,N_7768,N_7940);
xor U8385 (N_8385,N_7997,N_7702);
nor U8386 (N_8386,N_7980,N_7531);
nand U8387 (N_8387,N_7644,N_7824);
and U8388 (N_8388,N_7913,N_7984);
and U8389 (N_8389,N_7808,N_7554);
or U8390 (N_8390,N_7967,N_7995);
xor U8391 (N_8391,N_7530,N_7770);
nand U8392 (N_8392,N_7914,N_7804);
nor U8393 (N_8393,N_7728,N_7742);
and U8394 (N_8394,N_7800,N_7615);
nand U8395 (N_8395,N_7818,N_7872);
and U8396 (N_8396,N_7583,N_7732);
xor U8397 (N_8397,N_7586,N_7830);
nor U8398 (N_8398,N_7605,N_7924);
and U8399 (N_8399,N_7815,N_7983);
nand U8400 (N_8400,N_7583,N_7699);
and U8401 (N_8401,N_7595,N_7643);
or U8402 (N_8402,N_7829,N_7791);
and U8403 (N_8403,N_7963,N_7996);
nand U8404 (N_8404,N_7944,N_7950);
or U8405 (N_8405,N_7550,N_7861);
or U8406 (N_8406,N_7992,N_7577);
and U8407 (N_8407,N_7937,N_7902);
xnor U8408 (N_8408,N_7770,N_7792);
nor U8409 (N_8409,N_7937,N_7977);
xor U8410 (N_8410,N_7749,N_7879);
and U8411 (N_8411,N_7550,N_7764);
or U8412 (N_8412,N_7887,N_7868);
nor U8413 (N_8413,N_7587,N_7709);
and U8414 (N_8414,N_7714,N_7843);
nor U8415 (N_8415,N_7956,N_7709);
nor U8416 (N_8416,N_7758,N_7873);
xnor U8417 (N_8417,N_7788,N_7736);
xnor U8418 (N_8418,N_7778,N_7998);
nor U8419 (N_8419,N_7941,N_7760);
and U8420 (N_8420,N_7553,N_7952);
xor U8421 (N_8421,N_7998,N_7545);
or U8422 (N_8422,N_7528,N_7833);
nand U8423 (N_8423,N_7785,N_7546);
nor U8424 (N_8424,N_7983,N_7619);
xor U8425 (N_8425,N_7720,N_7870);
nand U8426 (N_8426,N_7598,N_7540);
nand U8427 (N_8427,N_7721,N_7848);
or U8428 (N_8428,N_7921,N_7709);
nor U8429 (N_8429,N_7772,N_7877);
and U8430 (N_8430,N_7878,N_7571);
nand U8431 (N_8431,N_7637,N_7711);
xnor U8432 (N_8432,N_7607,N_7564);
xnor U8433 (N_8433,N_7980,N_7959);
xor U8434 (N_8434,N_7986,N_7836);
and U8435 (N_8435,N_7627,N_7773);
nor U8436 (N_8436,N_7785,N_7868);
nor U8437 (N_8437,N_7890,N_7827);
xnor U8438 (N_8438,N_7896,N_7874);
nand U8439 (N_8439,N_7663,N_7574);
nand U8440 (N_8440,N_7694,N_7974);
nand U8441 (N_8441,N_7837,N_7969);
and U8442 (N_8442,N_7786,N_7704);
xor U8443 (N_8443,N_7993,N_7833);
nor U8444 (N_8444,N_7621,N_7709);
nand U8445 (N_8445,N_7710,N_7847);
or U8446 (N_8446,N_7599,N_7519);
and U8447 (N_8447,N_7913,N_7631);
xnor U8448 (N_8448,N_7707,N_7682);
nand U8449 (N_8449,N_7736,N_7917);
nand U8450 (N_8450,N_7950,N_7830);
and U8451 (N_8451,N_7667,N_7762);
or U8452 (N_8452,N_7792,N_7552);
nor U8453 (N_8453,N_7903,N_7806);
and U8454 (N_8454,N_7951,N_7840);
and U8455 (N_8455,N_7966,N_7830);
and U8456 (N_8456,N_7776,N_7557);
or U8457 (N_8457,N_7843,N_7748);
or U8458 (N_8458,N_7646,N_7764);
or U8459 (N_8459,N_7694,N_7993);
or U8460 (N_8460,N_7699,N_7657);
nand U8461 (N_8461,N_7685,N_7635);
xor U8462 (N_8462,N_7843,N_7840);
nor U8463 (N_8463,N_7986,N_7941);
xnor U8464 (N_8464,N_7788,N_7984);
and U8465 (N_8465,N_7682,N_7961);
or U8466 (N_8466,N_7648,N_7984);
and U8467 (N_8467,N_7540,N_7720);
and U8468 (N_8468,N_7731,N_7663);
xor U8469 (N_8469,N_7688,N_7889);
nor U8470 (N_8470,N_7785,N_7970);
xor U8471 (N_8471,N_7515,N_7618);
xor U8472 (N_8472,N_7674,N_7534);
xor U8473 (N_8473,N_7644,N_7997);
nand U8474 (N_8474,N_7811,N_7940);
or U8475 (N_8475,N_7655,N_7665);
or U8476 (N_8476,N_7684,N_7548);
nor U8477 (N_8477,N_7889,N_7771);
or U8478 (N_8478,N_7828,N_7810);
nand U8479 (N_8479,N_7961,N_7870);
nand U8480 (N_8480,N_7528,N_7733);
xnor U8481 (N_8481,N_7519,N_7998);
and U8482 (N_8482,N_7902,N_7530);
and U8483 (N_8483,N_7999,N_7866);
nor U8484 (N_8484,N_7803,N_7809);
or U8485 (N_8485,N_7624,N_7570);
nand U8486 (N_8486,N_7860,N_7809);
or U8487 (N_8487,N_7836,N_7729);
xnor U8488 (N_8488,N_7970,N_7503);
nand U8489 (N_8489,N_7928,N_7641);
or U8490 (N_8490,N_7701,N_7944);
or U8491 (N_8491,N_7822,N_7817);
nand U8492 (N_8492,N_7740,N_7565);
nand U8493 (N_8493,N_7589,N_7929);
nand U8494 (N_8494,N_7682,N_7773);
and U8495 (N_8495,N_7654,N_7589);
and U8496 (N_8496,N_7604,N_7502);
or U8497 (N_8497,N_7973,N_7870);
xnor U8498 (N_8498,N_7974,N_7997);
or U8499 (N_8499,N_7531,N_7604);
nor U8500 (N_8500,N_8096,N_8393);
nor U8501 (N_8501,N_8372,N_8136);
or U8502 (N_8502,N_8098,N_8298);
xnor U8503 (N_8503,N_8295,N_8488);
or U8504 (N_8504,N_8012,N_8092);
nand U8505 (N_8505,N_8057,N_8017);
nor U8506 (N_8506,N_8264,N_8306);
and U8507 (N_8507,N_8127,N_8308);
nor U8508 (N_8508,N_8338,N_8399);
nand U8509 (N_8509,N_8190,N_8242);
xor U8510 (N_8510,N_8042,N_8235);
xor U8511 (N_8511,N_8420,N_8070);
and U8512 (N_8512,N_8122,N_8419);
nand U8513 (N_8513,N_8126,N_8258);
xnor U8514 (N_8514,N_8394,N_8252);
xnor U8515 (N_8515,N_8221,N_8456);
or U8516 (N_8516,N_8203,N_8305);
nor U8517 (N_8517,N_8451,N_8046);
and U8518 (N_8518,N_8061,N_8412);
and U8519 (N_8519,N_8450,N_8313);
xnor U8520 (N_8520,N_8171,N_8388);
nand U8521 (N_8521,N_8320,N_8418);
or U8522 (N_8522,N_8001,N_8265);
or U8523 (N_8523,N_8438,N_8312);
nor U8524 (N_8524,N_8144,N_8052);
or U8525 (N_8525,N_8432,N_8261);
nand U8526 (N_8526,N_8352,N_8251);
nand U8527 (N_8527,N_8085,N_8005);
and U8528 (N_8528,N_8000,N_8379);
and U8529 (N_8529,N_8030,N_8371);
or U8530 (N_8530,N_8254,N_8321);
xor U8531 (N_8531,N_8198,N_8260);
nor U8532 (N_8532,N_8426,N_8011);
xnor U8533 (N_8533,N_8073,N_8077);
xor U8534 (N_8534,N_8421,N_8246);
or U8535 (N_8535,N_8007,N_8493);
xor U8536 (N_8536,N_8256,N_8279);
nor U8537 (N_8537,N_8486,N_8185);
nor U8538 (N_8538,N_8120,N_8187);
or U8539 (N_8539,N_8117,N_8377);
xor U8540 (N_8540,N_8140,N_8165);
nor U8541 (N_8541,N_8469,N_8414);
and U8542 (N_8542,N_8292,N_8445);
nand U8543 (N_8543,N_8031,N_8044);
nand U8544 (N_8544,N_8079,N_8478);
and U8545 (N_8545,N_8214,N_8128);
and U8546 (N_8546,N_8158,N_8496);
nand U8547 (N_8547,N_8118,N_8180);
nand U8548 (N_8548,N_8027,N_8336);
nand U8549 (N_8549,N_8266,N_8236);
and U8550 (N_8550,N_8028,N_8047);
nor U8551 (N_8551,N_8440,N_8170);
xor U8552 (N_8552,N_8431,N_8327);
nor U8553 (N_8553,N_8457,N_8111);
or U8554 (N_8554,N_8318,N_8272);
or U8555 (N_8555,N_8288,N_8036);
xnor U8556 (N_8556,N_8439,N_8113);
and U8557 (N_8557,N_8444,N_8468);
nor U8558 (N_8558,N_8480,N_8342);
and U8559 (N_8559,N_8286,N_8249);
and U8560 (N_8560,N_8225,N_8039);
nor U8561 (N_8561,N_8055,N_8311);
nor U8562 (N_8562,N_8051,N_8477);
nor U8563 (N_8563,N_8041,N_8411);
nand U8564 (N_8564,N_8008,N_8402);
or U8565 (N_8565,N_8029,N_8357);
and U8566 (N_8566,N_8083,N_8224);
or U8567 (N_8567,N_8234,N_8003);
and U8568 (N_8568,N_8442,N_8470);
nand U8569 (N_8569,N_8063,N_8010);
nor U8570 (N_8570,N_8160,N_8222);
xnor U8571 (N_8571,N_8403,N_8002);
nor U8572 (N_8572,N_8080,N_8263);
xnor U8573 (N_8573,N_8189,N_8151);
nand U8574 (N_8574,N_8141,N_8369);
xnor U8575 (N_8575,N_8209,N_8159);
nand U8576 (N_8576,N_8212,N_8290);
or U8577 (N_8577,N_8270,N_8076);
nor U8578 (N_8578,N_8386,N_8177);
or U8579 (N_8579,N_8259,N_8385);
or U8580 (N_8580,N_8217,N_8032);
nand U8581 (N_8581,N_8156,N_8389);
nor U8582 (N_8582,N_8004,N_8178);
xnor U8583 (N_8583,N_8404,N_8181);
or U8584 (N_8584,N_8153,N_8335);
nor U8585 (N_8585,N_8415,N_8395);
nand U8586 (N_8586,N_8476,N_8139);
xnor U8587 (N_8587,N_8125,N_8435);
or U8588 (N_8588,N_8300,N_8243);
nor U8589 (N_8589,N_8365,N_8274);
or U8590 (N_8590,N_8213,N_8215);
nor U8591 (N_8591,N_8110,N_8167);
xnor U8592 (N_8592,N_8043,N_8378);
xnor U8593 (N_8593,N_8054,N_8359);
or U8594 (N_8594,N_8328,N_8339);
xnor U8595 (N_8595,N_8434,N_8172);
nand U8596 (N_8596,N_8184,N_8138);
or U8597 (N_8597,N_8109,N_8376);
xor U8598 (N_8598,N_8100,N_8287);
xor U8599 (N_8599,N_8490,N_8471);
and U8600 (N_8600,N_8174,N_8463);
and U8601 (N_8601,N_8355,N_8091);
xor U8602 (N_8602,N_8233,N_8390);
xor U8603 (N_8603,N_8087,N_8331);
nand U8604 (N_8604,N_8449,N_8142);
or U8605 (N_8605,N_8485,N_8025);
xnor U8606 (N_8606,N_8448,N_8193);
nand U8607 (N_8607,N_8455,N_8484);
or U8608 (N_8608,N_8143,N_8137);
nand U8609 (N_8609,N_8253,N_8090);
or U8610 (N_8610,N_8461,N_8062);
nand U8611 (N_8611,N_8132,N_8074);
nand U8612 (N_8612,N_8208,N_8387);
and U8613 (N_8613,N_8285,N_8150);
and U8614 (N_8614,N_8400,N_8226);
nor U8615 (N_8615,N_8454,N_8145);
xor U8616 (N_8616,N_8101,N_8333);
nand U8617 (N_8617,N_8075,N_8218);
nor U8618 (N_8618,N_8237,N_8381);
and U8619 (N_8619,N_8182,N_8425);
and U8620 (N_8620,N_8367,N_8179);
nand U8621 (N_8621,N_8164,N_8459);
xnor U8622 (N_8622,N_8013,N_8229);
and U8623 (N_8623,N_8162,N_8334);
and U8624 (N_8624,N_8344,N_8424);
and U8625 (N_8625,N_8497,N_8245);
and U8626 (N_8626,N_8105,N_8398);
and U8627 (N_8627,N_8093,N_8020);
nand U8628 (N_8628,N_8437,N_8195);
or U8629 (N_8629,N_8303,N_8199);
xor U8630 (N_8630,N_8309,N_8006);
or U8631 (N_8631,N_8356,N_8278);
xor U8632 (N_8632,N_8345,N_8391);
or U8633 (N_8633,N_8099,N_8019);
and U8634 (N_8634,N_8384,N_8464);
xor U8635 (N_8635,N_8353,N_8465);
xnor U8636 (N_8636,N_8409,N_8161);
or U8637 (N_8637,N_8284,N_8211);
xnor U8638 (N_8638,N_8244,N_8417);
nand U8639 (N_8639,N_8157,N_8201);
xor U8640 (N_8640,N_8239,N_8035);
nor U8641 (N_8641,N_8262,N_8416);
nor U8642 (N_8642,N_8489,N_8374);
xnor U8643 (N_8643,N_8067,N_8361);
nor U8644 (N_8644,N_8069,N_8206);
or U8645 (N_8645,N_8370,N_8495);
nor U8646 (N_8646,N_8453,N_8392);
nand U8647 (N_8647,N_8360,N_8135);
xor U8648 (N_8648,N_8396,N_8269);
or U8649 (N_8649,N_8410,N_8350);
nand U8650 (N_8650,N_8397,N_8479);
xor U8651 (N_8651,N_8022,N_8238);
and U8652 (N_8652,N_8149,N_8422);
and U8653 (N_8653,N_8037,N_8066);
xor U8654 (N_8654,N_8319,N_8045);
xnor U8655 (N_8655,N_8146,N_8481);
nor U8656 (N_8656,N_8483,N_8192);
and U8657 (N_8657,N_8297,N_8148);
or U8658 (N_8658,N_8363,N_8107);
or U8659 (N_8659,N_8401,N_8228);
and U8660 (N_8660,N_8084,N_8219);
nand U8661 (N_8661,N_8094,N_8071);
nand U8662 (N_8662,N_8343,N_8296);
or U8663 (N_8663,N_8498,N_8407);
or U8664 (N_8664,N_8322,N_8499);
xnor U8665 (N_8665,N_8257,N_8330);
nand U8666 (N_8666,N_8072,N_8466);
and U8667 (N_8667,N_8314,N_8049);
nor U8668 (N_8668,N_8053,N_8131);
nor U8669 (N_8669,N_8293,N_8183);
and U8670 (N_8670,N_8166,N_8196);
nand U8671 (N_8671,N_8277,N_8240);
and U8672 (N_8672,N_8462,N_8154);
xnor U8673 (N_8673,N_8492,N_8316);
xnor U8674 (N_8674,N_8056,N_8009);
nand U8675 (N_8675,N_8216,N_8467);
nand U8676 (N_8676,N_8408,N_8186);
xnor U8677 (N_8677,N_8275,N_8016);
xnor U8678 (N_8678,N_8337,N_8405);
nand U8679 (N_8679,N_8033,N_8289);
and U8680 (N_8680,N_8380,N_8474);
and U8681 (N_8681,N_8223,N_8383);
nor U8682 (N_8682,N_8200,N_8436);
nor U8683 (N_8683,N_8241,N_8354);
nor U8684 (N_8684,N_8282,N_8299);
or U8685 (N_8685,N_8024,N_8482);
and U8686 (N_8686,N_8423,N_8121);
xnor U8687 (N_8687,N_8119,N_8034);
nor U8688 (N_8688,N_8018,N_8210);
nand U8689 (N_8689,N_8368,N_8175);
nor U8690 (N_8690,N_8323,N_8329);
xor U8691 (N_8691,N_8173,N_8147);
nand U8692 (N_8692,N_8220,N_8276);
and U8693 (N_8693,N_8307,N_8349);
and U8694 (N_8694,N_8429,N_8058);
or U8695 (N_8695,N_8129,N_8494);
xor U8696 (N_8696,N_8112,N_8487);
or U8697 (N_8697,N_8068,N_8108);
nor U8698 (N_8698,N_8103,N_8097);
xor U8699 (N_8699,N_8152,N_8267);
and U8700 (N_8700,N_8168,N_8473);
or U8701 (N_8701,N_8326,N_8373);
nor U8702 (N_8702,N_8268,N_8202);
or U8703 (N_8703,N_8089,N_8427);
nor U8704 (N_8704,N_8114,N_8294);
xnor U8705 (N_8705,N_8026,N_8433);
and U8706 (N_8706,N_8064,N_8441);
nand U8707 (N_8707,N_8048,N_8191);
nor U8708 (N_8708,N_8460,N_8341);
or U8709 (N_8709,N_8060,N_8324);
nor U8710 (N_8710,N_8205,N_8346);
nor U8711 (N_8711,N_8102,N_8248);
nand U8712 (N_8712,N_8194,N_8104);
nor U8713 (N_8713,N_8231,N_8250);
nand U8714 (N_8714,N_8458,N_8227);
nor U8715 (N_8715,N_8447,N_8271);
or U8716 (N_8716,N_8207,N_8281);
and U8717 (N_8717,N_8050,N_8163);
nand U8718 (N_8718,N_8082,N_8204);
xor U8719 (N_8719,N_8230,N_8428);
or U8720 (N_8720,N_8304,N_8130);
nand U8721 (N_8721,N_8280,N_8301);
xor U8722 (N_8722,N_8095,N_8197);
xnor U8723 (N_8723,N_8446,N_8116);
nor U8724 (N_8724,N_8472,N_8059);
and U8725 (N_8725,N_8283,N_8065);
or U8726 (N_8726,N_8348,N_8366);
and U8727 (N_8727,N_8406,N_8123);
nor U8728 (N_8728,N_8188,N_8430);
or U8729 (N_8729,N_8040,N_8169);
nand U8730 (N_8730,N_8014,N_8358);
or U8731 (N_8731,N_8332,N_8325);
or U8732 (N_8732,N_8291,N_8023);
and U8733 (N_8733,N_8176,N_8452);
and U8734 (N_8734,N_8015,N_8255);
nand U8735 (N_8735,N_8491,N_8340);
nor U8736 (N_8736,N_8081,N_8413);
xor U8737 (N_8737,N_8232,N_8364);
nand U8738 (N_8738,N_8078,N_8347);
or U8739 (N_8739,N_8124,N_8362);
or U8740 (N_8740,N_8088,N_8375);
and U8741 (N_8741,N_8133,N_8315);
nor U8742 (N_8742,N_8021,N_8247);
nand U8743 (N_8743,N_8310,N_8475);
nor U8744 (N_8744,N_8382,N_8115);
or U8745 (N_8745,N_8134,N_8086);
nor U8746 (N_8746,N_8155,N_8351);
xor U8747 (N_8747,N_8443,N_8302);
xnor U8748 (N_8748,N_8038,N_8273);
and U8749 (N_8749,N_8106,N_8317);
nand U8750 (N_8750,N_8181,N_8035);
xnor U8751 (N_8751,N_8433,N_8456);
nand U8752 (N_8752,N_8083,N_8240);
xor U8753 (N_8753,N_8015,N_8411);
nor U8754 (N_8754,N_8344,N_8135);
nor U8755 (N_8755,N_8008,N_8319);
or U8756 (N_8756,N_8028,N_8423);
nor U8757 (N_8757,N_8078,N_8357);
or U8758 (N_8758,N_8176,N_8168);
nand U8759 (N_8759,N_8183,N_8060);
and U8760 (N_8760,N_8172,N_8077);
and U8761 (N_8761,N_8098,N_8055);
and U8762 (N_8762,N_8127,N_8076);
and U8763 (N_8763,N_8469,N_8099);
xnor U8764 (N_8764,N_8493,N_8408);
and U8765 (N_8765,N_8489,N_8217);
nand U8766 (N_8766,N_8083,N_8440);
nand U8767 (N_8767,N_8493,N_8139);
nor U8768 (N_8768,N_8035,N_8493);
nor U8769 (N_8769,N_8448,N_8078);
or U8770 (N_8770,N_8067,N_8420);
xor U8771 (N_8771,N_8492,N_8059);
or U8772 (N_8772,N_8061,N_8165);
nand U8773 (N_8773,N_8150,N_8216);
or U8774 (N_8774,N_8337,N_8285);
nand U8775 (N_8775,N_8026,N_8461);
and U8776 (N_8776,N_8349,N_8376);
nor U8777 (N_8777,N_8031,N_8183);
xor U8778 (N_8778,N_8478,N_8015);
xnor U8779 (N_8779,N_8072,N_8087);
nand U8780 (N_8780,N_8144,N_8189);
or U8781 (N_8781,N_8173,N_8363);
or U8782 (N_8782,N_8110,N_8457);
nand U8783 (N_8783,N_8221,N_8001);
or U8784 (N_8784,N_8100,N_8151);
and U8785 (N_8785,N_8492,N_8129);
or U8786 (N_8786,N_8253,N_8408);
and U8787 (N_8787,N_8110,N_8326);
or U8788 (N_8788,N_8215,N_8057);
nor U8789 (N_8789,N_8370,N_8020);
and U8790 (N_8790,N_8047,N_8238);
xnor U8791 (N_8791,N_8018,N_8160);
xnor U8792 (N_8792,N_8285,N_8260);
nand U8793 (N_8793,N_8177,N_8384);
nand U8794 (N_8794,N_8408,N_8023);
xnor U8795 (N_8795,N_8390,N_8044);
nor U8796 (N_8796,N_8323,N_8478);
or U8797 (N_8797,N_8013,N_8202);
nand U8798 (N_8798,N_8006,N_8147);
or U8799 (N_8799,N_8189,N_8086);
or U8800 (N_8800,N_8132,N_8470);
xor U8801 (N_8801,N_8341,N_8150);
xor U8802 (N_8802,N_8212,N_8325);
nor U8803 (N_8803,N_8075,N_8089);
nor U8804 (N_8804,N_8276,N_8076);
nor U8805 (N_8805,N_8336,N_8139);
or U8806 (N_8806,N_8285,N_8201);
nor U8807 (N_8807,N_8350,N_8369);
and U8808 (N_8808,N_8490,N_8024);
xor U8809 (N_8809,N_8351,N_8161);
nand U8810 (N_8810,N_8461,N_8077);
or U8811 (N_8811,N_8089,N_8276);
xnor U8812 (N_8812,N_8204,N_8023);
or U8813 (N_8813,N_8033,N_8251);
nor U8814 (N_8814,N_8115,N_8413);
nand U8815 (N_8815,N_8496,N_8485);
nor U8816 (N_8816,N_8046,N_8316);
nor U8817 (N_8817,N_8135,N_8081);
nand U8818 (N_8818,N_8139,N_8317);
nand U8819 (N_8819,N_8044,N_8405);
or U8820 (N_8820,N_8186,N_8321);
and U8821 (N_8821,N_8149,N_8035);
and U8822 (N_8822,N_8087,N_8060);
nor U8823 (N_8823,N_8145,N_8019);
or U8824 (N_8824,N_8088,N_8449);
or U8825 (N_8825,N_8043,N_8088);
nand U8826 (N_8826,N_8214,N_8468);
and U8827 (N_8827,N_8224,N_8260);
or U8828 (N_8828,N_8252,N_8290);
nand U8829 (N_8829,N_8203,N_8471);
nor U8830 (N_8830,N_8272,N_8132);
nand U8831 (N_8831,N_8110,N_8455);
nor U8832 (N_8832,N_8395,N_8275);
nor U8833 (N_8833,N_8350,N_8440);
xor U8834 (N_8834,N_8225,N_8066);
or U8835 (N_8835,N_8269,N_8128);
and U8836 (N_8836,N_8002,N_8265);
and U8837 (N_8837,N_8335,N_8113);
nor U8838 (N_8838,N_8391,N_8311);
nor U8839 (N_8839,N_8418,N_8046);
nand U8840 (N_8840,N_8488,N_8034);
nand U8841 (N_8841,N_8040,N_8074);
xor U8842 (N_8842,N_8139,N_8430);
nand U8843 (N_8843,N_8089,N_8358);
nand U8844 (N_8844,N_8042,N_8119);
and U8845 (N_8845,N_8010,N_8405);
and U8846 (N_8846,N_8360,N_8276);
and U8847 (N_8847,N_8119,N_8057);
nand U8848 (N_8848,N_8444,N_8257);
nor U8849 (N_8849,N_8414,N_8381);
xnor U8850 (N_8850,N_8175,N_8459);
xor U8851 (N_8851,N_8063,N_8204);
or U8852 (N_8852,N_8068,N_8021);
xnor U8853 (N_8853,N_8138,N_8451);
xor U8854 (N_8854,N_8183,N_8402);
nor U8855 (N_8855,N_8040,N_8407);
or U8856 (N_8856,N_8451,N_8060);
and U8857 (N_8857,N_8150,N_8257);
nand U8858 (N_8858,N_8212,N_8400);
and U8859 (N_8859,N_8418,N_8204);
xor U8860 (N_8860,N_8318,N_8028);
xor U8861 (N_8861,N_8076,N_8346);
and U8862 (N_8862,N_8092,N_8379);
or U8863 (N_8863,N_8340,N_8004);
xor U8864 (N_8864,N_8329,N_8378);
xor U8865 (N_8865,N_8065,N_8418);
nor U8866 (N_8866,N_8172,N_8366);
or U8867 (N_8867,N_8015,N_8257);
or U8868 (N_8868,N_8036,N_8423);
nor U8869 (N_8869,N_8063,N_8215);
and U8870 (N_8870,N_8193,N_8218);
xor U8871 (N_8871,N_8006,N_8065);
nand U8872 (N_8872,N_8168,N_8227);
xnor U8873 (N_8873,N_8184,N_8258);
nand U8874 (N_8874,N_8123,N_8446);
or U8875 (N_8875,N_8353,N_8255);
nor U8876 (N_8876,N_8210,N_8139);
and U8877 (N_8877,N_8412,N_8241);
xnor U8878 (N_8878,N_8155,N_8162);
or U8879 (N_8879,N_8374,N_8366);
or U8880 (N_8880,N_8225,N_8364);
nand U8881 (N_8881,N_8056,N_8402);
and U8882 (N_8882,N_8393,N_8324);
xor U8883 (N_8883,N_8385,N_8230);
nand U8884 (N_8884,N_8205,N_8342);
or U8885 (N_8885,N_8126,N_8092);
nor U8886 (N_8886,N_8112,N_8471);
xnor U8887 (N_8887,N_8446,N_8256);
nor U8888 (N_8888,N_8064,N_8017);
and U8889 (N_8889,N_8192,N_8096);
nor U8890 (N_8890,N_8231,N_8082);
nand U8891 (N_8891,N_8043,N_8364);
and U8892 (N_8892,N_8175,N_8431);
or U8893 (N_8893,N_8252,N_8170);
and U8894 (N_8894,N_8436,N_8076);
or U8895 (N_8895,N_8062,N_8439);
xnor U8896 (N_8896,N_8327,N_8190);
or U8897 (N_8897,N_8173,N_8075);
nand U8898 (N_8898,N_8469,N_8306);
and U8899 (N_8899,N_8266,N_8125);
nor U8900 (N_8900,N_8498,N_8489);
nand U8901 (N_8901,N_8195,N_8387);
and U8902 (N_8902,N_8241,N_8485);
nor U8903 (N_8903,N_8343,N_8270);
or U8904 (N_8904,N_8294,N_8379);
and U8905 (N_8905,N_8215,N_8167);
or U8906 (N_8906,N_8234,N_8434);
and U8907 (N_8907,N_8364,N_8083);
nand U8908 (N_8908,N_8276,N_8408);
nand U8909 (N_8909,N_8039,N_8390);
and U8910 (N_8910,N_8058,N_8131);
xor U8911 (N_8911,N_8388,N_8119);
nand U8912 (N_8912,N_8125,N_8459);
xnor U8913 (N_8913,N_8384,N_8011);
nand U8914 (N_8914,N_8182,N_8317);
or U8915 (N_8915,N_8364,N_8051);
nor U8916 (N_8916,N_8085,N_8063);
and U8917 (N_8917,N_8483,N_8274);
or U8918 (N_8918,N_8136,N_8464);
nor U8919 (N_8919,N_8233,N_8427);
and U8920 (N_8920,N_8472,N_8356);
or U8921 (N_8921,N_8103,N_8026);
nor U8922 (N_8922,N_8160,N_8013);
xor U8923 (N_8923,N_8485,N_8497);
nand U8924 (N_8924,N_8059,N_8417);
and U8925 (N_8925,N_8198,N_8031);
and U8926 (N_8926,N_8184,N_8429);
nand U8927 (N_8927,N_8091,N_8415);
nand U8928 (N_8928,N_8465,N_8282);
xnor U8929 (N_8929,N_8387,N_8083);
nand U8930 (N_8930,N_8045,N_8314);
nor U8931 (N_8931,N_8248,N_8329);
and U8932 (N_8932,N_8264,N_8383);
nor U8933 (N_8933,N_8117,N_8491);
and U8934 (N_8934,N_8177,N_8375);
nor U8935 (N_8935,N_8358,N_8372);
xnor U8936 (N_8936,N_8488,N_8172);
xor U8937 (N_8937,N_8189,N_8441);
or U8938 (N_8938,N_8312,N_8100);
nand U8939 (N_8939,N_8366,N_8422);
or U8940 (N_8940,N_8072,N_8365);
nor U8941 (N_8941,N_8451,N_8040);
xor U8942 (N_8942,N_8173,N_8346);
nand U8943 (N_8943,N_8268,N_8487);
nor U8944 (N_8944,N_8132,N_8233);
nor U8945 (N_8945,N_8472,N_8303);
nand U8946 (N_8946,N_8146,N_8366);
xor U8947 (N_8947,N_8106,N_8467);
nand U8948 (N_8948,N_8482,N_8183);
or U8949 (N_8949,N_8086,N_8384);
xor U8950 (N_8950,N_8425,N_8019);
and U8951 (N_8951,N_8204,N_8477);
xor U8952 (N_8952,N_8174,N_8013);
nor U8953 (N_8953,N_8039,N_8108);
xor U8954 (N_8954,N_8258,N_8133);
or U8955 (N_8955,N_8371,N_8372);
or U8956 (N_8956,N_8252,N_8461);
xor U8957 (N_8957,N_8126,N_8469);
xor U8958 (N_8958,N_8163,N_8441);
and U8959 (N_8959,N_8149,N_8400);
nor U8960 (N_8960,N_8302,N_8284);
and U8961 (N_8961,N_8352,N_8330);
nor U8962 (N_8962,N_8405,N_8483);
and U8963 (N_8963,N_8195,N_8490);
and U8964 (N_8964,N_8012,N_8479);
nor U8965 (N_8965,N_8409,N_8396);
nand U8966 (N_8966,N_8284,N_8194);
or U8967 (N_8967,N_8388,N_8451);
nor U8968 (N_8968,N_8173,N_8066);
and U8969 (N_8969,N_8435,N_8272);
xnor U8970 (N_8970,N_8171,N_8113);
and U8971 (N_8971,N_8007,N_8434);
or U8972 (N_8972,N_8277,N_8085);
and U8973 (N_8973,N_8311,N_8334);
and U8974 (N_8974,N_8370,N_8261);
or U8975 (N_8975,N_8095,N_8047);
or U8976 (N_8976,N_8051,N_8027);
nand U8977 (N_8977,N_8329,N_8279);
nor U8978 (N_8978,N_8223,N_8240);
nand U8979 (N_8979,N_8053,N_8215);
xnor U8980 (N_8980,N_8406,N_8400);
and U8981 (N_8981,N_8451,N_8342);
or U8982 (N_8982,N_8187,N_8069);
nor U8983 (N_8983,N_8317,N_8226);
nor U8984 (N_8984,N_8321,N_8382);
or U8985 (N_8985,N_8342,N_8053);
nor U8986 (N_8986,N_8434,N_8259);
nor U8987 (N_8987,N_8412,N_8358);
xor U8988 (N_8988,N_8356,N_8034);
nand U8989 (N_8989,N_8437,N_8404);
and U8990 (N_8990,N_8204,N_8400);
xor U8991 (N_8991,N_8153,N_8440);
or U8992 (N_8992,N_8050,N_8326);
and U8993 (N_8993,N_8267,N_8226);
nand U8994 (N_8994,N_8090,N_8245);
and U8995 (N_8995,N_8408,N_8297);
and U8996 (N_8996,N_8288,N_8316);
nor U8997 (N_8997,N_8232,N_8363);
xor U8998 (N_8998,N_8344,N_8254);
nand U8999 (N_8999,N_8485,N_8348);
and U9000 (N_9000,N_8885,N_8785);
or U9001 (N_9001,N_8615,N_8772);
nor U9002 (N_9002,N_8767,N_8892);
nand U9003 (N_9003,N_8764,N_8959);
xor U9004 (N_9004,N_8634,N_8760);
nor U9005 (N_9005,N_8904,N_8652);
xnor U9006 (N_9006,N_8878,N_8993);
xnor U9007 (N_9007,N_8860,N_8985);
nor U9008 (N_9008,N_8972,N_8620);
or U9009 (N_9009,N_8931,N_8989);
and U9010 (N_9010,N_8802,N_8887);
and U9011 (N_9011,N_8874,N_8742);
nand U9012 (N_9012,N_8949,N_8707);
nor U9013 (N_9013,N_8674,N_8974);
and U9014 (N_9014,N_8679,N_8791);
nor U9015 (N_9015,N_8950,N_8810);
or U9016 (N_9016,N_8755,N_8928);
and U9017 (N_9017,N_8946,N_8952);
nand U9018 (N_9018,N_8938,N_8827);
nor U9019 (N_9019,N_8681,N_8787);
xnor U9020 (N_9020,N_8593,N_8942);
nor U9021 (N_9021,N_8694,N_8696);
and U9022 (N_9022,N_8947,N_8608);
and U9023 (N_9023,N_8886,N_8539);
xnor U9024 (N_9024,N_8843,N_8852);
and U9025 (N_9025,N_8711,N_8908);
xnor U9026 (N_9026,N_8883,N_8840);
and U9027 (N_9027,N_8570,N_8725);
xor U9028 (N_9028,N_8525,N_8646);
or U9029 (N_9029,N_8566,N_8968);
xor U9030 (N_9030,N_8877,N_8779);
nand U9031 (N_9031,N_8988,N_8638);
and U9032 (N_9032,N_8800,N_8574);
and U9033 (N_9033,N_8901,N_8973);
and U9034 (N_9034,N_8799,N_8664);
nand U9035 (N_9035,N_8813,N_8732);
and U9036 (N_9036,N_8847,N_8925);
nand U9037 (N_9037,N_8835,N_8605);
or U9038 (N_9038,N_8603,N_8778);
xor U9039 (N_9039,N_8849,N_8713);
and U9040 (N_9040,N_8569,N_8876);
nand U9041 (N_9041,N_8804,N_8841);
nor U9042 (N_9042,N_8830,N_8596);
or U9043 (N_9043,N_8551,N_8667);
xor U9044 (N_9044,N_8890,N_8821);
nand U9045 (N_9045,N_8684,N_8553);
nand U9046 (N_9046,N_8992,N_8951);
nand U9047 (N_9047,N_8744,N_8671);
nand U9048 (N_9048,N_8897,N_8786);
nand U9049 (N_9049,N_8514,N_8561);
nor U9050 (N_9050,N_8617,N_8526);
nand U9051 (N_9051,N_8902,N_8589);
xnor U9052 (N_9052,N_8807,N_8544);
xor U9053 (N_9053,N_8996,N_8583);
and U9054 (N_9054,N_8967,N_8913);
xor U9055 (N_9055,N_8599,N_8748);
xnor U9056 (N_9056,N_8688,N_8839);
and U9057 (N_9057,N_8898,N_8805);
xnor U9058 (N_9058,N_8611,N_8714);
nor U9059 (N_9059,N_8573,N_8592);
or U9060 (N_9060,N_8695,N_8584);
xnor U9061 (N_9061,N_8563,N_8757);
or U9062 (N_9062,N_8618,N_8654);
nand U9063 (N_9063,N_8531,N_8833);
nand U9064 (N_9064,N_8588,N_8571);
nor U9065 (N_9065,N_8870,N_8953);
and U9066 (N_9066,N_8702,N_8644);
nand U9067 (N_9067,N_8623,N_8735);
nor U9068 (N_9068,N_8556,N_8960);
xor U9069 (N_9069,N_8701,N_8976);
xnor U9070 (N_9070,N_8758,N_8624);
nor U9071 (N_9071,N_8834,N_8964);
and U9072 (N_9072,N_8979,N_8806);
nand U9073 (N_9073,N_8675,N_8676);
and U9074 (N_9074,N_8929,N_8923);
nor U9075 (N_9075,N_8625,N_8712);
and U9076 (N_9076,N_8914,N_8773);
xor U9077 (N_9077,N_8582,N_8808);
and U9078 (N_9078,N_8829,N_8685);
nor U9079 (N_9079,N_8579,N_8723);
nor U9080 (N_9080,N_8637,N_8743);
nand U9081 (N_9081,N_8769,N_8708);
xnor U9082 (N_9082,N_8934,N_8716);
or U9083 (N_9083,N_8981,N_8590);
nand U9084 (N_9084,N_8782,N_8948);
nor U9085 (N_9085,N_8794,N_8824);
nand U9086 (N_9086,N_8521,N_8536);
nor U9087 (N_9087,N_8647,N_8932);
and U9088 (N_9088,N_8519,N_8724);
or U9089 (N_9089,N_8614,N_8628);
nand U9090 (N_9090,N_8687,N_8722);
xor U9091 (N_9091,N_8848,N_8846);
and U9092 (N_9092,N_8927,N_8554);
nor U9093 (N_9093,N_8509,N_8520);
xnor U9094 (N_9094,N_8768,N_8856);
or U9095 (N_9095,N_8930,N_8899);
xnor U9096 (N_9096,N_8838,N_8881);
or U9097 (N_9097,N_8650,N_8512);
or U9098 (N_9098,N_8857,N_8591);
nor U9099 (N_9099,N_8645,N_8954);
nand U9100 (N_9100,N_8889,N_8919);
or U9101 (N_9101,N_8619,N_8659);
and U9102 (N_9102,N_8749,N_8971);
nor U9103 (N_9103,N_8872,N_8698);
xor U9104 (N_9104,N_8535,N_8587);
xor U9105 (N_9105,N_8789,N_8759);
or U9106 (N_9106,N_8859,N_8905);
nor U9107 (N_9107,N_8661,N_8817);
and U9108 (N_9108,N_8503,N_8595);
nor U9109 (N_9109,N_8547,N_8994);
xnor U9110 (N_9110,N_8803,N_8730);
xor U9111 (N_9111,N_8507,N_8630);
xor U9112 (N_9112,N_8532,N_8506);
xnor U9113 (N_9113,N_8678,N_8736);
xnor U9114 (N_9114,N_8770,N_8680);
xor U9115 (N_9115,N_8998,N_8867);
nor U9116 (N_9116,N_8715,N_8796);
nor U9117 (N_9117,N_8997,N_8893);
nor U9118 (N_9118,N_8564,N_8729);
xnor U9119 (N_9119,N_8658,N_8879);
nand U9120 (N_9120,N_8970,N_8500);
nand U9121 (N_9121,N_8606,N_8837);
nand U9122 (N_9122,N_8665,N_8858);
nor U9123 (N_9123,N_8957,N_8537);
xnor U9124 (N_9124,N_8540,N_8580);
xnor U9125 (N_9125,N_8522,N_8945);
xnor U9126 (N_9126,N_8762,N_8751);
nand U9127 (N_9127,N_8636,N_8530);
nor U9128 (N_9128,N_8918,N_8832);
nor U9129 (N_9129,N_8741,N_8823);
nor U9130 (N_9130,N_8781,N_8873);
nand U9131 (N_9131,N_8578,N_8533);
nor U9132 (N_9132,N_8861,N_8880);
xnor U9133 (N_9133,N_8737,N_8987);
nor U9134 (N_9134,N_8915,N_8501);
nand U9135 (N_9135,N_8545,N_8869);
or U9136 (N_9136,N_8682,N_8763);
nor U9137 (N_9137,N_8999,N_8984);
and U9138 (N_9138,N_8643,N_8527);
or U9139 (N_9139,N_8907,N_8626);
and U9140 (N_9140,N_8822,N_8633);
nor U9141 (N_9141,N_8753,N_8831);
xnor U9142 (N_9142,N_8555,N_8896);
nand U9143 (N_9143,N_8691,N_8656);
xor U9144 (N_9144,N_8943,N_8750);
or U9145 (N_9145,N_8765,N_8756);
and U9146 (N_9146,N_8505,N_8982);
nor U9147 (N_9147,N_8727,N_8936);
xnor U9148 (N_9148,N_8657,N_8745);
xor U9149 (N_9149,N_8884,N_8937);
and U9150 (N_9150,N_8631,N_8783);
and U9151 (N_9151,N_8641,N_8801);
or U9152 (N_9152,N_8706,N_8673);
or U9153 (N_9153,N_8790,N_8677);
or U9154 (N_9154,N_8621,N_8940);
nor U9155 (N_9155,N_8819,N_8962);
nor U9156 (N_9156,N_8616,N_8866);
nor U9157 (N_9157,N_8662,N_8909);
and U9158 (N_9158,N_8548,N_8629);
or U9159 (N_9159,N_8690,N_8683);
or U9160 (N_9160,N_8502,N_8686);
xor U9161 (N_9161,N_8774,N_8709);
nand U9162 (N_9162,N_8602,N_8613);
nor U9163 (N_9163,N_8863,N_8775);
and U9164 (N_9164,N_8746,N_8900);
xnor U9165 (N_9165,N_8524,N_8935);
xnor U9166 (N_9166,N_8635,N_8597);
nor U9167 (N_9167,N_8784,N_8961);
nand U9168 (N_9168,N_8693,N_8534);
and U9169 (N_9169,N_8651,N_8568);
nor U9170 (N_9170,N_8720,N_8966);
nand U9171 (N_9171,N_8627,N_8538);
or U9172 (N_9172,N_8542,N_8868);
xor U9173 (N_9173,N_8851,N_8642);
and U9174 (N_9174,N_8549,N_8845);
nor U9175 (N_9175,N_8793,N_8515);
nor U9176 (N_9176,N_8567,N_8721);
nor U9177 (N_9177,N_8917,N_8776);
nor U9178 (N_9178,N_8853,N_8903);
nor U9179 (N_9179,N_8814,N_8731);
nand U9180 (N_9180,N_8818,N_8543);
and U9181 (N_9181,N_8990,N_8717);
nand U9182 (N_9182,N_8963,N_8939);
nor U9183 (N_9183,N_8906,N_8891);
nand U9184 (N_9184,N_8557,N_8825);
or U9185 (N_9185,N_8916,N_8850);
or U9186 (N_9186,N_8511,N_8622);
and U9187 (N_9187,N_8639,N_8894);
nand U9188 (N_9188,N_8977,N_8921);
and U9189 (N_9189,N_8991,N_8809);
nor U9190 (N_9190,N_8660,N_8510);
xnor U9191 (N_9191,N_8792,N_8612);
or U9192 (N_9192,N_8777,N_8738);
nor U9193 (N_9193,N_8920,N_8640);
nor U9194 (N_9194,N_8820,N_8780);
and U9195 (N_9195,N_8728,N_8766);
and U9196 (N_9196,N_8610,N_8672);
and U9197 (N_9197,N_8562,N_8924);
nor U9198 (N_9198,N_8854,N_8747);
nor U9199 (N_9199,N_8546,N_8600);
xor U9200 (N_9200,N_8700,N_8529);
nor U9201 (N_9201,N_8871,N_8926);
nor U9202 (N_9202,N_8958,N_8733);
or U9203 (N_9203,N_8689,N_8944);
nor U9204 (N_9204,N_8740,N_8585);
nand U9205 (N_9205,N_8788,N_8669);
and U9206 (N_9206,N_8828,N_8586);
and U9207 (N_9207,N_8798,N_8516);
xnor U9208 (N_9208,N_8653,N_8911);
nor U9209 (N_9209,N_8670,N_8550);
nand U9210 (N_9210,N_8978,N_8826);
xor U9211 (N_9211,N_8692,N_8797);
and U9212 (N_9212,N_8875,N_8812);
nand U9213 (N_9213,N_8609,N_8560);
nor U9214 (N_9214,N_8922,N_8718);
nor U9215 (N_9215,N_8710,N_8513);
nand U9216 (N_9216,N_8518,N_8862);
and U9217 (N_9217,N_8726,N_8983);
nor U9218 (N_9218,N_8955,N_8795);
nand U9219 (N_9219,N_8739,N_8704);
nand U9220 (N_9220,N_8910,N_8965);
or U9221 (N_9221,N_8576,N_8604);
xnor U9222 (N_9222,N_8754,N_8598);
nand U9223 (N_9223,N_8565,N_8517);
or U9224 (N_9224,N_8836,N_8986);
xor U9225 (N_9225,N_8719,N_8558);
and U9226 (N_9226,N_8699,N_8842);
or U9227 (N_9227,N_8705,N_8504);
xnor U9228 (N_9228,N_8933,N_8864);
xnor U9229 (N_9229,N_8697,N_8663);
and U9230 (N_9230,N_8844,N_8703);
or U9231 (N_9231,N_8912,N_8771);
or U9232 (N_9232,N_8855,N_8575);
or U9233 (N_9233,N_8995,N_8956);
or U9234 (N_9234,N_8541,N_8559);
or U9235 (N_9235,N_8888,N_8648);
nand U9236 (N_9236,N_8523,N_8969);
nand U9237 (N_9237,N_8668,N_8655);
nand U9238 (N_9238,N_8815,N_8632);
nand U9239 (N_9239,N_8666,N_8752);
xor U9240 (N_9240,N_8528,N_8865);
nand U9241 (N_9241,N_8761,N_8941);
and U9242 (N_9242,N_8572,N_8508);
or U9243 (N_9243,N_8607,N_8811);
nor U9244 (N_9244,N_8975,N_8734);
xor U9245 (N_9245,N_8552,N_8649);
xor U9246 (N_9246,N_8581,N_8895);
and U9247 (N_9247,N_8594,N_8601);
or U9248 (N_9248,N_8577,N_8882);
nand U9249 (N_9249,N_8816,N_8980);
and U9250 (N_9250,N_8627,N_8640);
or U9251 (N_9251,N_8768,N_8754);
xor U9252 (N_9252,N_8560,N_8605);
nand U9253 (N_9253,N_8880,N_8532);
nand U9254 (N_9254,N_8978,N_8793);
nand U9255 (N_9255,N_8525,N_8728);
nor U9256 (N_9256,N_8579,N_8826);
or U9257 (N_9257,N_8581,N_8701);
or U9258 (N_9258,N_8810,N_8690);
and U9259 (N_9259,N_8873,N_8827);
nor U9260 (N_9260,N_8710,N_8916);
and U9261 (N_9261,N_8867,N_8742);
nand U9262 (N_9262,N_8635,N_8892);
nand U9263 (N_9263,N_8901,N_8812);
nand U9264 (N_9264,N_8888,N_8536);
xor U9265 (N_9265,N_8917,N_8883);
or U9266 (N_9266,N_8956,N_8620);
xnor U9267 (N_9267,N_8715,N_8763);
nor U9268 (N_9268,N_8904,N_8725);
or U9269 (N_9269,N_8631,N_8726);
nor U9270 (N_9270,N_8712,N_8698);
or U9271 (N_9271,N_8785,N_8640);
nand U9272 (N_9272,N_8540,N_8898);
and U9273 (N_9273,N_8595,N_8538);
nor U9274 (N_9274,N_8518,N_8920);
nor U9275 (N_9275,N_8665,N_8945);
nor U9276 (N_9276,N_8528,N_8733);
xor U9277 (N_9277,N_8753,N_8874);
xor U9278 (N_9278,N_8819,N_8517);
xor U9279 (N_9279,N_8562,N_8610);
xnor U9280 (N_9280,N_8660,N_8982);
xor U9281 (N_9281,N_8890,N_8977);
nand U9282 (N_9282,N_8732,N_8816);
nor U9283 (N_9283,N_8601,N_8755);
nor U9284 (N_9284,N_8775,N_8743);
and U9285 (N_9285,N_8886,N_8810);
nand U9286 (N_9286,N_8582,N_8609);
nor U9287 (N_9287,N_8906,N_8561);
nand U9288 (N_9288,N_8934,N_8832);
xnor U9289 (N_9289,N_8881,N_8906);
or U9290 (N_9290,N_8870,N_8805);
and U9291 (N_9291,N_8536,N_8577);
nor U9292 (N_9292,N_8669,N_8776);
nand U9293 (N_9293,N_8564,N_8911);
nor U9294 (N_9294,N_8805,N_8707);
nand U9295 (N_9295,N_8780,N_8860);
or U9296 (N_9296,N_8980,N_8744);
xnor U9297 (N_9297,N_8845,N_8607);
nor U9298 (N_9298,N_8708,N_8787);
nand U9299 (N_9299,N_8775,N_8765);
and U9300 (N_9300,N_8591,N_8721);
and U9301 (N_9301,N_8890,N_8919);
nand U9302 (N_9302,N_8847,N_8582);
xnor U9303 (N_9303,N_8570,N_8968);
or U9304 (N_9304,N_8922,N_8662);
and U9305 (N_9305,N_8674,N_8673);
nor U9306 (N_9306,N_8928,N_8649);
or U9307 (N_9307,N_8768,N_8680);
or U9308 (N_9308,N_8558,N_8974);
nor U9309 (N_9309,N_8789,N_8970);
nor U9310 (N_9310,N_8669,N_8777);
xor U9311 (N_9311,N_8795,N_8784);
or U9312 (N_9312,N_8728,N_8862);
or U9313 (N_9313,N_8874,N_8908);
and U9314 (N_9314,N_8606,N_8969);
nor U9315 (N_9315,N_8534,N_8552);
nand U9316 (N_9316,N_8615,N_8510);
xnor U9317 (N_9317,N_8947,N_8517);
nand U9318 (N_9318,N_8531,N_8501);
nor U9319 (N_9319,N_8640,N_8993);
or U9320 (N_9320,N_8904,N_8945);
xnor U9321 (N_9321,N_8814,N_8726);
nand U9322 (N_9322,N_8507,N_8666);
nand U9323 (N_9323,N_8666,N_8785);
or U9324 (N_9324,N_8915,N_8938);
and U9325 (N_9325,N_8859,N_8830);
and U9326 (N_9326,N_8657,N_8795);
nor U9327 (N_9327,N_8529,N_8537);
or U9328 (N_9328,N_8673,N_8852);
nor U9329 (N_9329,N_8905,N_8539);
xor U9330 (N_9330,N_8506,N_8675);
nor U9331 (N_9331,N_8718,N_8867);
nand U9332 (N_9332,N_8510,N_8821);
and U9333 (N_9333,N_8507,N_8774);
nor U9334 (N_9334,N_8899,N_8650);
xor U9335 (N_9335,N_8922,N_8841);
nor U9336 (N_9336,N_8736,N_8504);
nand U9337 (N_9337,N_8692,N_8942);
nand U9338 (N_9338,N_8981,N_8861);
or U9339 (N_9339,N_8989,N_8745);
xor U9340 (N_9340,N_8993,N_8807);
nor U9341 (N_9341,N_8758,N_8707);
xnor U9342 (N_9342,N_8817,N_8874);
and U9343 (N_9343,N_8531,N_8886);
nand U9344 (N_9344,N_8764,N_8886);
nor U9345 (N_9345,N_8975,N_8655);
xnor U9346 (N_9346,N_8916,N_8838);
and U9347 (N_9347,N_8558,N_8521);
and U9348 (N_9348,N_8899,N_8555);
nand U9349 (N_9349,N_8694,N_8632);
xor U9350 (N_9350,N_8640,N_8762);
or U9351 (N_9351,N_8648,N_8736);
or U9352 (N_9352,N_8842,N_8609);
and U9353 (N_9353,N_8878,N_8621);
or U9354 (N_9354,N_8563,N_8508);
and U9355 (N_9355,N_8691,N_8989);
xor U9356 (N_9356,N_8836,N_8532);
and U9357 (N_9357,N_8511,N_8805);
and U9358 (N_9358,N_8596,N_8728);
nand U9359 (N_9359,N_8927,N_8592);
nor U9360 (N_9360,N_8702,N_8793);
nor U9361 (N_9361,N_8794,N_8636);
nand U9362 (N_9362,N_8799,N_8524);
or U9363 (N_9363,N_8733,N_8993);
nor U9364 (N_9364,N_8532,N_8762);
nand U9365 (N_9365,N_8928,N_8793);
and U9366 (N_9366,N_8854,N_8615);
or U9367 (N_9367,N_8818,N_8760);
or U9368 (N_9368,N_8922,N_8940);
nand U9369 (N_9369,N_8786,N_8835);
and U9370 (N_9370,N_8629,N_8891);
or U9371 (N_9371,N_8569,N_8953);
nand U9372 (N_9372,N_8629,N_8602);
or U9373 (N_9373,N_8769,N_8661);
nand U9374 (N_9374,N_8782,N_8773);
or U9375 (N_9375,N_8612,N_8936);
and U9376 (N_9376,N_8767,N_8984);
or U9377 (N_9377,N_8752,N_8623);
nand U9378 (N_9378,N_8812,N_8612);
and U9379 (N_9379,N_8957,N_8940);
xor U9380 (N_9380,N_8833,N_8865);
xor U9381 (N_9381,N_8686,N_8528);
or U9382 (N_9382,N_8525,N_8983);
and U9383 (N_9383,N_8976,N_8851);
xnor U9384 (N_9384,N_8788,N_8778);
nor U9385 (N_9385,N_8949,N_8631);
xor U9386 (N_9386,N_8764,N_8892);
nor U9387 (N_9387,N_8629,N_8762);
and U9388 (N_9388,N_8702,N_8947);
nor U9389 (N_9389,N_8831,N_8823);
nand U9390 (N_9390,N_8553,N_8920);
nand U9391 (N_9391,N_8594,N_8962);
nor U9392 (N_9392,N_8779,N_8997);
and U9393 (N_9393,N_8807,N_8759);
and U9394 (N_9394,N_8771,N_8972);
or U9395 (N_9395,N_8894,N_8703);
nand U9396 (N_9396,N_8708,N_8593);
or U9397 (N_9397,N_8821,N_8891);
or U9398 (N_9398,N_8751,N_8906);
xnor U9399 (N_9399,N_8888,N_8989);
nand U9400 (N_9400,N_8537,N_8988);
or U9401 (N_9401,N_8754,N_8766);
xor U9402 (N_9402,N_8691,N_8633);
xnor U9403 (N_9403,N_8512,N_8569);
or U9404 (N_9404,N_8669,N_8587);
nor U9405 (N_9405,N_8683,N_8614);
xnor U9406 (N_9406,N_8815,N_8745);
and U9407 (N_9407,N_8863,N_8838);
or U9408 (N_9408,N_8562,N_8697);
nand U9409 (N_9409,N_8547,N_8778);
nor U9410 (N_9410,N_8578,N_8948);
nor U9411 (N_9411,N_8696,N_8560);
or U9412 (N_9412,N_8992,N_8823);
nor U9413 (N_9413,N_8665,N_8906);
nor U9414 (N_9414,N_8950,N_8526);
nand U9415 (N_9415,N_8727,N_8632);
nor U9416 (N_9416,N_8745,N_8589);
or U9417 (N_9417,N_8938,N_8566);
nor U9418 (N_9418,N_8820,N_8886);
xor U9419 (N_9419,N_8827,N_8682);
and U9420 (N_9420,N_8532,N_8571);
xnor U9421 (N_9421,N_8591,N_8873);
and U9422 (N_9422,N_8539,N_8872);
xnor U9423 (N_9423,N_8809,N_8902);
nor U9424 (N_9424,N_8549,N_8832);
or U9425 (N_9425,N_8925,N_8697);
and U9426 (N_9426,N_8755,N_8630);
nand U9427 (N_9427,N_8676,N_8929);
nand U9428 (N_9428,N_8616,N_8573);
and U9429 (N_9429,N_8952,N_8978);
and U9430 (N_9430,N_8734,N_8649);
nand U9431 (N_9431,N_8883,N_8815);
and U9432 (N_9432,N_8874,N_8948);
and U9433 (N_9433,N_8877,N_8915);
or U9434 (N_9434,N_8852,N_8832);
xnor U9435 (N_9435,N_8703,N_8689);
and U9436 (N_9436,N_8959,N_8775);
or U9437 (N_9437,N_8657,N_8826);
xnor U9438 (N_9438,N_8971,N_8643);
nor U9439 (N_9439,N_8726,N_8984);
xor U9440 (N_9440,N_8963,N_8636);
xnor U9441 (N_9441,N_8875,N_8910);
nand U9442 (N_9442,N_8908,N_8764);
or U9443 (N_9443,N_8759,N_8991);
nor U9444 (N_9444,N_8598,N_8748);
nand U9445 (N_9445,N_8968,N_8608);
and U9446 (N_9446,N_8734,N_8943);
nand U9447 (N_9447,N_8791,N_8594);
nor U9448 (N_9448,N_8799,N_8625);
nor U9449 (N_9449,N_8867,N_8744);
xnor U9450 (N_9450,N_8864,N_8827);
nor U9451 (N_9451,N_8782,N_8748);
nand U9452 (N_9452,N_8626,N_8828);
xor U9453 (N_9453,N_8908,N_8899);
or U9454 (N_9454,N_8991,N_8888);
nand U9455 (N_9455,N_8684,N_8755);
or U9456 (N_9456,N_8653,N_8534);
or U9457 (N_9457,N_8544,N_8524);
nor U9458 (N_9458,N_8631,N_8663);
or U9459 (N_9459,N_8847,N_8851);
or U9460 (N_9460,N_8918,N_8730);
nor U9461 (N_9461,N_8674,N_8765);
or U9462 (N_9462,N_8903,N_8991);
nor U9463 (N_9463,N_8795,N_8714);
and U9464 (N_9464,N_8574,N_8642);
nand U9465 (N_9465,N_8962,N_8703);
xor U9466 (N_9466,N_8645,N_8667);
and U9467 (N_9467,N_8605,N_8869);
or U9468 (N_9468,N_8657,N_8805);
xor U9469 (N_9469,N_8913,N_8876);
nand U9470 (N_9470,N_8994,N_8845);
and U9471 (N_9471,N_8580,N_8575);
nor U9472 (N_9472,N_8690,N_8921);
and U9473 (N_9473,N_8967,N_8978);
nor U9474 (N_9474,N_8960,N_8801);
or U9475 (N_9475,N_8988,N_8981);
xor U9476 (N_9476,N_8832,N_8622);
nor U9477 (N_9477,N_8991,N_8826);
nor U9478 (N_9478,N_8914,N_8596);
and U9479 (N_9479,N_8929,N_8647);
xnor U9480 (N_9480,N_8976,N_8660);
or U9481 (N_9481,N_8623,N_8769);
or U9482 (N_9482,N_8764,N_8639);
xor U9483 (N_9483,N_8595,N_8795);
nor U9484 (N_9484,N_8851,N_8927);
nor U9485 (N_9485,N_8640,N_8668);
and U9486 (N_9486,N_8702,N_8991);
nand U9487 (N_9487,N_8876,N_8897);
or U9488 (N_9488,N_8566,N_8827);
nand U9489 (N_9489,N_8800,N_8894);
xor U9490 (N_9490,N_8717,N_8538);
or U9491 (N_9491,N_8688,N_8875);
or U9492 (N_9492,N_8670,N_8793);
xor U9493 (N_9493,N_8805,N_8506);
nand U9494 (N_9494,N_8982,N_8858);
nand U9495 (N_9495,N_8740,N_8619);
and U9496 (N_9496,N_8560,N_8705);
xor U9497 (N_9497,N_8728,N_8996);
and U9498 (N_9498,N_8945,N_8773);
or U9499 (N_9499,N_8562,N_8589);
xor U9500 (N_9500,N_9409,N_9364);
xnor U9501 (N_9501,N_9106,N_9159);
nor U9502 (N_9502,N_9109,N_9046);
or U9503 (N_9503,N_9180,N_9402);
nor U9504 (N_9504,N_9123,N_9428);
xor U9505 (N_9505,N_9089,N_9295);
nand U9506 (N_9506,N_9058,N_9493);
or U9507 (N_9507,N_9119,N_9176);
nand U9508 (N_9508,N_9034,N_9211);
xor U9509 (N_9509,N_9267,N_9412);
nand U9510 (N_9510,N_9202,N_9039);
nor U9511 (N_9511,N_9189,N_9040);
nor U9512 (N_9512,N_9008,N_9482);
or U9513 (N_9513,N_9476,N_9239);
xnor U9514 (N_9514,N_9200,N_9093);
xnor U9515 (N_9515,N_9450,N_9312);
xor U9516 (N_9516,N_9197,N_9296);
nor U9517 (N_9517,N_9275,N_9027);
nor U9518 (N_9518,N_9225,N_9411);
xnor U9519 (N_9519,N_9155,N_9327);
and U9520 (N_9520,N_9021,N_9222);
or U9521 (N_9521,N_9319,N_9118);
or U9522 (N_9522,N_9458,N_9309);
xor U9523 (N_9523,N_9212,N_9220);
or U9524 (N_9524,N_9463,N_9209);
xor U9525 (N_9525,N_9254,N_9215);
nand U9526 (N_9526,N_9377,N_9183);
xnor U9527 (N_9527,N_9337,N_9461);
xnor U9528 (N_9528,N_9066,N_9470);
xor U9529 (N_9529,N_9410,N_9110);
and U9530 (N_9530,N_9247,N_9175);
xor U9531 (N_9531,N_9279,N_9017);
nor U9532 (N_9532,N_9347,N_9379);
and U9533 (N_9533,N_9260,N_9321);
and U9534 (N_9534,N_9230,N_9459);
or U9535 (N_9535,N_9298,N_9468);
nand U9536 (N_9536,N_9491,N_9043);
nand U9537 (N_9537,N_9422,N_9152);
nor U9538 (N_9538,N_9182,N_9100);
and U9539 (N_9539,N_9181,N_9444);
nor U9540 (N_9540,N_9400,N_9431);
nand U9541 (N_9541,N_9318,N_9453);
nand U9542 (N_9542,N_9498,N_9292);
or U9543 (N_9543,N_9258,N_9054);
xor U9544 (N_9544,N_9105,N_9168);
or U9545 (N_9545,N_9045,N_9290);
and U9546 (N_9546,N_9193,N_9029);
or U9547 (N_9547,N_9098,N_9381);
and U9548 (N_9548,N_9462,N_9185);
and U9549 (N_9549,N_9146,N_9125);
nand U9550 (N_9550,N_9130,N_9243);
and U9551 (N_9551,N_9078,N_9313);
nand U9552 (N_9552,N_9241,N_9164);
xnor U9553 (N_9553,N_9452,N_9214);
xor U9554 (N_9554,N_9216,N_9355);
and U9555 (N_9555,N_9447,N_9120);
and U9556 (N_9556,N_9490,N_9187);
or U9557 (N_9557,N_9204,N_9086);
or U9558 (N_9558,N_9070,N_9208);
or U9559 (N_9559,N_9373,N_9328);
xor U9560 (N_9560,N_9443,N_9136);
nand U9561 (N_9561,N_9406,N_9263);
xor U9562 (N_9562,N_9286,N_9485);
xor U9563 (N_9563,N_9166,N_9437);
nor U9564 (N_9564,N_9018,N_9154);
xnor U9565 (N_9565,N_9325,N_9002);
or U9566 (N_9566,N_9446,N_9455);
nand U9567 (N_9567,N_9147,N_9484);
or U9568 (N_9568,N_9288,N_9307);
and U9569 (N_9569,N_9145,N_9196);
and U9570 (N_9570,N_9163,N_9388);
or U9571 (N_9571,N_9479,N_9236);
or U9572 (N_9572,N_9389,N_9257);
and U9573 (N_9573,N_9068,N_9324);
nand U9574 (N_9574,N_9304,N_9011);
nand U9575 (N_9575,N_9138,N_9234);
nand U9576 (N_9576,N_9418,N_9179);
and U9577 (N_9577,N_9486,N_9391);
or U9578 (N_9578,N_9367,N_9369);
xnor U9579 (N_9579,N_9067,N_9435);
and U9580 (N_9580,N_9037,N_9419);
nand U9581 (N_9581,N_9240,N_9050);
nand U9582 (N_9582,N_9371,N_9362);
nor U9583 (N_9583,N_9440,N_9022);
and U9584 (N_9584,N_9310,N_9160);
xnor U9585 (N_9585,N_9460,N_9270);
and U9586 (N_9586,N_9438,N_9386);
nand U9587 (N_9587,N_9210,N_9469);
and U9588 (N_9588,N_9156,N_9333);
xor U9589 (N_9589,N_9124,N_9112);
and U9590 (N_9590,N_9272,N_9473);
nand U9591 (N_9591,N_9107,N_9032);
or U9592 (N_9592,N_9133,N_9382);
or U9593 (N_9593,N_9301,N_9495);
and U9594 (N_9594,N_9280,N_9273);
and U9595 (N_9595,N_9265,N_9398);
nand U9596 (N_9596,N_9198,N_9413);
or U9597 (N_9597,N_9150,N_9084);
nand U9598 (N_9598,N_9334,N_9436);
and U9599 (N_9599,N_9077,N_9056);
and U9600 (N_9600,N_9308,N_9173);
nand U9601 (N_9601,N_9131,N_9302);
or U9602 (N_9602,N_9001,N_9417);
nand U9603 (N_9603,N_9278,N_9139);
nor U9604 (N_9604,N_9363,N_9071);
nand U9605 (N_9605,N_9285,N_9339);
xor U9606 (N_9606,N_9101,N_9158);
nand U9607 (N_9607,N_9383,N_9264);
or U9608 (N_9608,N_9466,N_9300);
or U9609 (N_9609,N_9360,N_9143);
nor U9610 (N_9610,N_9354,N_9451);
nor U9611 (N_9611,N_9303,N_9372);
and U9612 (N_9612,N_9103,N_9358);
nor U9613 (N_9613,N_9047,N_9194);
and U9614 (N_9614,N_9433,N_9148);
nor U9615 (N_9615,N_9316,N_9315);
and U9616 (N_9616,N_9338,N_9297);
nor U9617 (N_9617,N_9282,N_9269);
nor U9618 (N_9618,N_9111,N_9206);
and U9619 (N_9619,N_9439,N_9359);
or U9620 (N_9620,N_9244,N_9115);
and U9621 (N_9621,N_9044,N_9357);
and U9622 (N_9622,N_9167,N_9480);
or U9623 (N_9623,N_9010,N_9340);
nand U9624 (N_9624,N_9169,N_9251);
nor U9625 (N_9625,N_9420,N_9291);
xor U9626 (N_9626,N_9091,N_9405);
or U9627 (N_9627,N_9499,N_9335);
or U9628 (N_9628,N_9157,N_9283);
nor U9629 (N_9629,N_9294,N_9102);
and U9630 (N_9630,N_9121,N_9261);
nand U9631 (N_9631,N_9092,N_9028);
nand U9632 (N_9632,N_9082,N_9006);
nand U9633 (N_9633,N_9494,N_9242);
or U9634 (N_9634,N_9052,N_9186);
or U9635 (N_9635,N_9471,N_9079);
xor U9636 (N_9636,N_9095,N_9430);
xnor U9637 (N_9637,N_9449,N_9341);
xnor U9638 (N_9638,N_9262,N_9226);
or U9639 (N_9639,N_9249,N_9366);
xor U9640 (N_9640,N_9465,N_9427);
and U9641 (N_9641,N_9061,N_9271);
nand U9642 (N_9642,N_9016,N_9064);
or U9643 (N_9643,N_9423,N_9415);
nand U9644 (N_9644,N_9238,N_9231);
or U9645 (N_9645,N_9000,N_9069);
nor U9646 (N_9646,N_9429,N_9426);
nor U9647 (N_9647,N_9049,N_9434);
xnor U9648 (N_9648,N_9395,N_9475);
or U9649 (N_9649,N_9023,N_9454);
or U9650 (N_9650,N_9416,N_9219);
nand U9651 (N_9651,N_9343,N_9392);
nor U9652 (N_9652,N_9228,N_9425);
and U9653 (N_9653,N_9399,N_9087);
nand U9654 (N_9654,N_9059,N_9477);
or U9655 (N_9655,N_9456,N_9361);
nor U9656 (N_9656,N_9351,N_9090);
or U9657 (N_9657,N_9007,N_9060);
nor U9658 (N_9658,N_9104,N_9345);
and U9659 (N_9659,N_9057,N_9266);
or U9660 (N_9660,N_9274,N_9483);
xnor U9661 (N_9661,N_9404,N_9026);
nand U9662 (N_9662,N_9311,N_9385);
and U9663 (N_9663,N_9191,N_9250);
nand U9664 (N_9664,N_9132,N_9122);
and U9665 (N_9665,N_9199,N_9368);
nor U9666 (N_9666,N_9320,N_9108);
xor U9667 (N_9667,N_9009,N_9467);
and U9668 (N_9668,N_9048,N_9177);
or U9669 (N_9669,N_9088,N_9352);
and U9670 (N_9670,N_9117,N_9004);
nor U9671 (N_9671,N_9384,N_9277);
nor U9672 (N_9672,N_9195,N_9306);
nand U9673 (N_9673,N_9414,N_9128);
and U9674 (N_9674,N_9144,N_9174);
and U9675 (N_9675,N_9255,N_9072);
and U9676 (N_9676,N_9326,N_9237);
nand U9677 (N_9677,N_9080,N_9375);
nand U9678 (N_9678,N_9135,N_9031);
nor U9679 (N_9679,N_9390,N_9096);
xor U9680 (N_9680,N_9397,N_9094);
xnor U9681 (N_9681,N_9229,N_9323);
nand U9682 (N_9682,N_9253,N_9478);
or U9683 (N_9683,N_9063,N_9356);
and U9684 (N_9684,N_9492,N_9421);
or U9685 (N_9685,N_9305,N_9445);
nor U9686 (N_9686,N_9281,N_9188);
nand U9687 (N_9687,N_9142,N_9083);
and U9688 (N_9688,N_9432,N_9203);
or U9689 (N_9689,N_9393,N_9348);
and U9690 (N_9690,N_9401,N_9331);
or U9691 (N_9691,N_9127,N_9076);
and U9692 (N_9692,N_9408,N_9151);
nor U9693 (N_9693,N_9033,N_9481);
xor U9694 (N_9694,N_9370,N_9015);
or U9695 (N_9695,N_9448,N_9013);
xor U9696 (N_9696,N_9171,N_9153);
nor U9697 (N_9697,N_9051,N_9114);
or U9698 (N_9698,N_9041,N_9003);
nand U9699 (N_9699,N_9081,N_9365);
xnor U9700 (N_9700,N_9287,N_9116);
or U9701 (N_9701,N_9224,N_9020);
and U9702 (N_9702,N_9184,N_9289);
and U9703 (N_9703,N_9474,N_9129);
or U9704 (N_9704,N_9497,N_9342);
xnor U9705 (N_9705,N_9344,N_9162);
or U9706 (N_9706,N_9464,N_9172);
nor U9707 (N_9707,N_9317,N_9259);
nand U9708 (N_9708,N_9349,N_9024);
nand U9709 (N_9709,N_9073,N_9235);
nor U9710 (N_9710,N_9293,N_9457);
xor U9711 (N_9711,N_9376,N_9014);
and U9712 (N_9712,N_9149,N_9252);
nand U9713 (N_9713,N_9085,N_9074);
or U9714 (N_9714,N_9276,N_9097);
and U9715 (N_9715,N_9246,N_9380);
nand U9716 (N_9716,N_9137,N_9353);
xor U9717 (N_9717,N_9442,N_9207);
or U9718 (N_9718,N_9201,N_9075);
nand U9719 (N_9719,N_9036,N_9190);
or U9720 (N_9720,N_9035,N_9134);
xor U9721 (N_9721,N_9407,N_9489);
or U9722 (N_9722,N_9329,N_9165);
and U9723 (N_9723,N_9232,N_9005);
or U9724 (N_9724,N_9192,N_9178);
nand U9725 (N_9725,N_9140,N_9055);
xor U9726 (N_9726,N_9025,N_9227);
or U9727 (N_9727,N_9248,N_9170);
nand U9728 (N_9728,N_9387,N_9218);
or U9729 (N_9729,N_9065,N_9403);
or U9730 (N_9730,N_9099,N_9350);
xor U9731 (N_9731,N_9332,N_9299);
or U9732 (N_9732,N_9141,N_9314);
nand U9733 (N_9733,N_9256,N_9394);
nor U9734 (N_9734,N_9053,N_9330);
and U9735 (N_9735,N_9336,N_9038);
nand U9736 (N_9736,N_9496,N_9221);
xor U9737 (N_9737,N_9223,N_9233);
xor U9738 (N_9738,N_9042,N_9441);
xnor U9739 (N_9739,N_9472,N_9062);
and U9740 (N_9740,N_9487,N_9322);
nor U9741 (N_9741,N_9030,N_9245);
or U9742 (N_9742,N_9213,N_9126);
nor U9743 (N_9743,N_9113,N_9161);
or U9744 (N_9744,N_9346,N_9424);
nand U9745 (N_9745,N_9019,N_9205);
or U9746 (N_9746,N_9378,N_9217);
nor U9747 (N_9747,N_9396,N_9268);
nor U9748 (N_9748,N_9374,N_9012);
nor U9749 (N_9749,N_9284,N_9488);
nor U9750 (N_9750,N_9308,N_9315);
and U9751 (N_9751,N_9144,N_9037);
nor U9752 (N_9752,N_9248,N_9435);
and U9753 (N_9753,N_9250,N_9441);
or U9754 (N_9754,N_9060,N_9429);
or U9755 (N_9755,N_9417,N_9194);
nand U9756 (N_9756,N_9158,N_9205);
xnor U9757 (N_9757,N_9175,N_9439);
nand U9758 (N_9758,N_9083,N_9073);
and U9759 (N_9759,N_9441,N_9179);
nor U9760 (N_9760,N_9197,N_9381);
or U9761 (N_9761,N_9300,N_9037);
nor U9762 (N_9762,N_9256,N_9446);
or U9763 (N_9763,N_9062,N_9355);
xnor U9764 (N_9764,N_9400,N_9158);
nand U9765 (N_9765,N_9149,N_9400);
and U9766 (N_9766,N_9132,N_9429);
and U9767 (N_9767,N_9337,N_9126);
or U9768 (N_9768,N_9164,N_9100);
nor U9769 (N_9769,N_9412,N_9322);
nand U9770 (N_9770,N_9479,N_9346);
or U9771 (N_9771,N_9494,N_9447);
xor U9772 (N_9772,N_9407,N_9150);
nand U9773 (N_9773,N_9033,N_9269);
nor U9774 (N_9774,N_9487,N_9150);
and U9775 (N_9775,N_9185,N_9163);
nand U9776 (N_9776,N_9193,N_9422);
nor U9777 (N_9777,N_9069,N_9276);
xnor U9778 (N_9778,N_9330,N_9049);
or U9779 (N_9779,N_9043,N_9377);
xnor U9780 (N_9780,N_9108,N_9126);
xnor U9781 (N_9781,N_9305,N_9244);
nand U9782 (N_9782,N_9122,N_9454);
nor U9783 (N_9783,N_9296,N_9351);
and U9784 (N_9784,N_9446,N_9217);
xor U9785 (N_9785,N_9093,N_9013);
and U9786 (N_9786,N_9170,N_9436);
nand U9787 (N_9787,N_9307,N_9428);
or U9788 (N_9788,N_9066,N_9248);
nor U9789 (N_9789,N_9066,N_9161);
nand U9790 (N_9790,N_9045,N_9141);
or U9791 (N_9791,N_9327,N_9083);
xnor U9792 (N_9792,N_9232,N_9158);
xor U9793 (N_9793,N_9071,N_9053);
nor U9794 (N_9794,N_9235,N_9355);
nand U9795 (N_9795,N_9075,N_9272);
or U9796 (N_9796,N_9356,N_9498);
nand U9797 (N_9797,N_9184,N_9295);
xor U9798 (N_9798,N_9123,N_9246);
xnor U9799 (N_9799,N_9485,N_9440);
or U9800 (N_9800,N_9053,N_9080);
nand U9801 (N_9801,N_9228,N_9485);
nand U9802 (N_9802,N_9102,N_9021);
nor U9803 (N_9803,N_9313,N_9141);
or U9804 (N_9804,N_9326,N_9017);
xor U9805 (N_9805,N_9020,N_9497);
or U9806 (N_9806,N_9416,N_9260);
xor U9807 (N_9807,N_9204,N_9499);
or U9808 (N_9808,N_9409,N_9401);
xor U9809 (N_9809,N_9485,N_9168);
nand U9810 (N_9810,N_9352,N_9497);
nand U9811 (N_9811,N_9319,N_9443);
and U9812 (N_9812,N_9102,N_9020);
or U9813 (N_9813,N_9018,N_9191);
nand U9814 (N_9814,N_9254,N_9235);
nand U9815 (N_9815,N_9095,N_9100);
nor U9816 (N_9816,N_9499,N_9432);
or U9817 (N_9817,N_9102,N_9468);
or U9818 (N_9818,N_9260,N_9152);
nor U9819 (N_9819,N_9227,N_9146);
or U9820 (N_9820,N_9455,N_9005);
nor U9821 (N_9821,N_9188,N_9159);
or U9822 (N_9822,N_9094,N_9193);
nand U9823 (N_9823,N_9171,N_9078);
nor U9824 (N_9824,N_9196,N_9183);
nand U9825 (N_9825,N_9286,N_9109);
nor U9826 (N_9826,N_9016,N_9105);
nand U9827 (N_9827,N_9296,N_9067);
and U9828 (N_9828,N_9238,N_9421);
or U9829 (N_9829,N_9118,N_9325);
nand U9830 (N_9830,N_9041,N_9079);
or U9831 (N_9831,N_9048,N_9326);
xor U9832 (N_9832,N_9095,N_9306);
xor U9833 (N_9833,N_9041,N_9437);
or U9834 (N_9834,N_9317,N_9239);
or U9835 (N_9835,N_9104,N_9134);
or U9836 (N_9836,N_9036,N_9164);
or U9837 (N_9837,N_9307,N_9375);
nor U9838 (N_9838,N_9483,N_9082);
nand U9839 (N_9839,N_9175,N_9231);
or U9840 (N_9840,N_9285,N_9209);
and U9841 (N_9841,N_9288,N_9269);
xor U9842 (N_9842,N_9252,N_9474);
nor U9843 (N_9843,N_9058,N_9332);
and U9844 (N_9844,N_9055,N_9379);
and U9845 (N_9845,N_9003,N_9345);
xnor U9846 (N_9846,N_9349,N_9423);
xor U9847 (N_9847,N_9055,N_9368);
or U9848 (N_9848,N_9062,N_9180);
nand U9849 (N_9849,N_9251,N_9236);
and U9850 (N_9850,N_9029,N_9438);
nor U9851 (N_9851,N_9020,N_9280);
or U9852 (N_9852,N_9120,N_9445);
nand U9853 (N_9853,N_9312,N_9421);
nor U9854 (N_9854,N_9153,N_9307);
nor U9855 (N_9855,N_9208,N_9068);
xor U9856 (N_9856,N_9072,N_9320);
or U9857 (N_9857,N_9054,N_9167);
nor U9858 (N_9858,N_9134,N_9029);
xnor U9859 (N_9859,N_9430,N_9243);
xor U9860 (N_9860,N_9369,N_9230);
or U9861 (N_9861,N_9377,N_9258);
and U9862 (N_9862,N_9399,N_9374);
xnor U9863 (N_9863,N_9435,N_9033);
or U9864 (N_9864,N_9263,N_9056);
nand U9865 (N_9865,N_9081,N_9306);
and U9866 (N_9866,N_9414,N_9378);
nor U9867 (N_9867,N_9413,N_9207);
and U9868 (N_9868,N_9202,N_9169);
xnor U9869 (N_9869,N_9371,N_9290);
or U9870 (N_9870,N_9028,N_9449);
xor U9871 (N_9871,N_9267,N_9455);
xnor U9872 (N_9872,N_9353,N_9439);
nand U9873 (N_9873,N_9099,N_9053);
nand U9874 (N_9874,N_9280,N_9498);
xor U9875 (N_9875,N_9219,N_9378);
and U9876 (N_9876,N_9350,N_9154);
and U9877 (N_9877,N_9110,N_9105);
and U9878 (N_9878,N_9231,N_9193);
and U9879 (N_9879,N_9491,N_9083);
nand U9880 (N_9880,N_9135,N_9212);
or U9881 (N_9881,N_9359,N_9483);
nand U9882 (N_9882,N_9402,N_9315);
or U9883 (N_9883,N_9250,N_9487);
nand U9884 (N_9884,N_9198,N_9305);
or U9885 (N_9885,N_9159,N_9367);
nand U9886 (N_9886,N_9416,N_9076);
nand U9887 (N_9887,N_9165,N_9279);
nand U9888 (N_9888,N_9329,N_9356);
nor U9889 (N_9889,N_9496,N_9123);
nor U9890 (N_9890,N_9309,N_9174);
or U9891 (N_9891,N_9009,N_9024);
and U9892 (N_9892,N_9426,N_9179);
nor U9893 (N_9893,N_9224,N_9111);
and U9894 (N_9894,N_9396,N_9379);
or U9895 (N_9895,N_9481,N_9166);
nor U9896 (N_9896,N_9023,N_9370);
nand U9897 (N_9897,N_9167,N_9393);
or U9898 (N_9898,N_9163,N_9319);
nor U9899 (N_9899,N_9117,N_9263);
nand U9900 (N_9900,N_9387,N_9445);
nand U9901 (N_9901,N_9058,N_9480);
xnor U9902 (N_9902,N_9211,N_9348);
nand U9903 (N_9903,N_9186,N_9121);
nand U9904 (N_9904,N_9081,N_9091);
and U9905 (N_9905,N_9407,N_9324);
nor U9906 (N_9906,N_9015,N_9298);
and U9907 (N_9907,N_9108,N_9271);
or U9908 (N_9908,N_9238,N_9294);
nand U9909 (N_9909,N_9190,N_9410);
xor U9910 (N_9910,N_9356,N_9072);
or U9911 (N_9911,N_9152,N_9064);
nor U9912 (N_9912,N_9277,N_9117);
nor U9913 (N_9913,N_9414,N_9364);
xor U9914 (N_9914,N_9049,N_9338);
and U9915 (N_9915,N_9495,N_9219);
nor U9916 (N_9916,N_9178,N_9391);
and U9917 (N_9917,N_9380,N_9277);
and U9918 (N_9918,N_9210,N_9211);
xor U9919 (N_9919,N_9213,N_9366);
and U9920 (N_9920,N_9196,N_9026);
nand U9921 (N_9921,N_9172,N_9053);
xnor U9922 (N_9922,N_9085,N_9209);
and U9923 (N_9923,N_9203,N_9055);
nor U9924 (N_9924,N_9250,N_9139);
and U9925 (N_9925,N_9383,N_9496);
nand U9926 (N_9926,N_9351,N_9009);
nand U9927 (N_9927,N_9238,N_9226);
nand U9928 (N_9928,N_9286,N_9319);
nand U9929 (N_9929,N_9118,N_9446);
and U9930 (N_9930,N_9481,N_9038);
nor U9931 (N_9931,N_9392,N_9148);
or U9932 (N_9932,N_9455,N_9101);
nor U9933 (N_9933,N_9226,N_9020);
nor U9934 (N_9934,N_9484,N_9182);
or U9935 (N_9935,N_9175,N_9129);
and U9936 (N_9936,N_9362,N_9382);
and U9937 (N_9937,N_9171,N_9417);
xnor U9938 (N_9938,N_9463,N_9166);
or U9939 (N_9939,N_9138,N_9196);
or U9940 (N_9940,N_9305,N_9121);
nand U9941 (N_9941,N_9036,N_9005);
xnor U9942 (N_9942,N_9250,N_9160);
or U9943 (N_9943,N_9134,N_9107);
xor U9944 (N_9944,N_9164,N_9089);
and U9945 (N_9945,N_9079,N_9269);
nor U9946 (N_9946,N_9449,N_9343);
xor U9947 (N_9947,N_9293,N_9196);
and U9948 (N_9948,N_9065,N_9218);
nand U9949 (N_9949,N_9271,N_9147);
and U9950 (N_9950,N_9408,N_9007);
xor U9951 (N_9951,N_9150,N_9280);
xnor U9952 (N_9952,N_9369,N_9205);
xor U9953 (N_9953,N_9429,N_9355);
nor U9954 (N_9954,N_9172,N_9214);
nand U9955 (N_9955,N_9150,N_9338);
nor U9956 (N_9956,N_9428,N_9112);
xor U9957 (N_9957,N_9411,N_9425);
nor U9958 (N_9958,N_9089,N_9070);
nor U9959 (N_9959,N_9029,N_9023);
xor U9960 (N_9960,N_9135,N_9332);
nand U9961 (N_9961,N_9480,N_9130);
xor U9962 (N_9962,N_9313,N_9382);
nor U9963 (N_9963,N_9292,N_9015);
xnor U9964 (N_9964,N_9113,N_9174);
and U9965 (N_9965,N_9286,N_9418);
xnor U9966 (N_9966,N_9113,N_9033);
nand U9967 (N_9967,N_9323,N_9061);
and U9968 (N_9968,N_9362,N_9213);
nand U9969 (N_9969,N_9431,N_9258);
nor U9970 (N_9970,N_9482,N_9427);
nand U9971 (N_9971,N_9068,N_9270);
nand U9972 (N_9972,N_9363,N_9123);
nand U9973 (N_9973,N_9179,N_9477);
or U9974 (N_9974,N_9180,N_9318);
or U9975 (N_9975,N_9123,N_9471);
nor U9976 (N_9976,N_9223,N_9135);
or U9977 (N_9977,N_9216,N_9479);
nand U9978 (N_9978,N_9006,N_9301);
or U9979 (N_9979,N_9228,N_9247);
or U9980 (N_9980,N_9177,N_9015);
nand U9981 (N_9981,N_9408,N_9277);
and U9982 (N_9982,N_9496,N_9336);
nand U9983 (N_9983,N_9333,N_9311);
xnor U9984 (N_9984,N_9360,N_9028);
nand U9985 (N_9985,N_9334,N_9087);
nand U9986 (N_9986,N_9319,N_9038);
nand U9987 (N_9987,N_9032,N_9074);
xnor U9988 (N_9988,N_9272,N_9461);
and U9989 (N_9989,N_9227,N_9195);
or U9990 (N_9990,N_9125,N_9197);
or U9991 (N_9991,N_9446,N_9220);
and U9992 (N_9992,N_9161,N_9401);
and U9993 (N_9993,N_9361,N_9334);
nand U9994 (N_9994,N_9463,N_9120);
or U9995 (N_9995,N_9324,N_9450);
and U9996 (N_9996,N_9308,N_9235);
and U9997 (N_9997,N_9273,N_9262);
nand U9998 (N_9998,N_9116,N_9275);
xor U9999 (N_9999,N_9075,N_9141);
nor U10000 (N_10000,N_9615,N_9816);
xnor U10001 (N_10001,N_9758,N_9664);
or U10002 (N_10002,N_9650,N_9954);
nor U10003 (N_10003,N_9542,N_9847);
xor U10004 (N_10004,N_9832,N_9944);
nor U10005 (N_10005,N_9785,N_9579);
xor U10006 (N_10006,N_9521,N_9956);
nand U10007 (N_10007,N_9842,N_9812);
or U10008 (N_10008,N_9750,N_9790);
and U10009 (N_10009,N_9532,N_9662);
or U10010 (N_10010,N_9753,N_9916);
xor U10011 (N_10011,N_9501,N_9519);
nand U10012 (N_10012,N_9605,N_9516);
xnor U10013 (N_10013,N_9965,N_9739);
and U10014 (N_10014,N_9639,N_9646);
or U10015 (N_10015,N_9815,N_9565);
nand U10016 (N_10016,N_9617,N_9952);
or U10017 (N_10017,N_9978,N_9935);
and U10018 (N_10018,N_9715,N_9975);
nand U10019 (N_10019,N_9746,N_9803);
and U10020 (N_10020,N_9530,N_9622);
xor U10021 (N_10021,N_9536,N_9787);
or U10022 (N_10022,N_9751,N_9767);
nor U10023 (N_10023,N_9540,N_9594);
xor U10024 (N_10024,N_9681,N_9652);
nor U10025 (N_10025,N_9930,N_9939);
or U10026 (N_10026,N_9929,N_9572);
and U10027 (N_10027,N_9821,N_9999);
and U10028 (N_10028,N_9581,N_9522);
nand U10029 (N_10029,N_9942,N_9610);
or U10030 (N_10030,N_9992,N_9877);
nor U10031 (N_10031,N_9776,N_9779);
nor U10032 (N_10032,N_9525,N_9917);
and U10033 (N_10033,N_9614,N_9834);
nand U10034 (N_10034,N_9564,N_9890);
or U10035 (N_10035,N_9840,N_9687);
nand U10036 (N_10036,N_9931,N_9642);
xor U10037 (N_10037,N_9860,N_9704);
or U10038 (N_10038,N_9977,N_9879);
xnor U10039 (N_10039,N_9577,N_9569);
nand U10040 (N_10040,N_9728,N_9578);
xnor U10041 (N_10041,N_9604,N_9838);
nand U10042 (N_10042,N_9894,N_9535);
or U10043 (N_10043,N_9724,N_9653);
or U10044 (N_10044,N_9924,N_9943);
nor U10045 (N_10045,N_9575,N_9524);
and U10046 (N_10046,N_9651,N_9689);
nor U10047 (N_10047,N_9744,N_9667);
xnor U10048 (N_10048,N_9829,N_9859);
and U10049 (N_10049,N_9580,N_9556);
nand U10050 (N_10050,N_9582,N_9854);
nor U10051 (N_10051,N_9804,N_9720);
nand U10052 (N_10052,N_9811,N_9749);
xnor U10053 (N_10053,N_9765,N_9792);
and U10054 (N_10054,N_9780,N_9958);
or U10055 (N_10055,N_9647,N_9598);
or U10056 (N_10056,N_9781,N_9887);
nor U10057 (N_10057,N_9595,N_9628);
and U10058 (N_10058,N_9980,N_9769);
or U10059 (N_10059,N_9723,N_9830);
nor U10060 (N_10060,N_9836,N_9730);
and U10061 (N_10061,N_9507,N_9979);
or U10062 (N_10062,N_9508,N_9982);
nand U10063 (N_10063,N_9764,N_9885);
nand U10064 (N_10064,N_9645,N_9858);
and U10065 (N_10065,N_9566,N_9857);
or U10066 (N_10066,N_9741,N_9563);
or U10067 (N_10067,N_9794,N_9809);
nand U10068 (N_10068,N_9915,N_9960);
nand U10069 (N_10069,N_9901,N_9756);
nand U10070 (N_10070,N_9551,N_9666);
xor U10071 (N_10071,N_9900,N_9547);
nand U10072 (N_10072,N_9731,N_9795);
and U10073 (N_10073,N_9874,N_9747);
and U10074 (N_10074,N_9963,N_9738);
xnor U10075 (N_10075,N_9846,N_9797);
or U10076 (N_10076,N_9990,N_9625);
nor U10077 (N_10077,N_9976,N_9884);
xor U10078 (N_10078,N_9727,N_9807);
nor U10079 (N_10079,N_9574,N_9693);
and U10080 (N_10080,N_9587,N_9709);
nor U10081 (N_10081,N_9757,N_9665);
or U10082 (N_10082,N_9627,N_9822);
xnor U10083 (N_10083,N_9696,N_9679);
or U10084 (N_10084,N_9782,N_9560);
nand U10085 (N_10085,N_9661,N_9786);
xnor U10086 (N_10086,N_9654,N_9655);
and U10087 (N_10087,N_9584,N_9706);
nor U10088 (N_10088,N_9596,N_9766);
and U10089 (N_10089,N_9714,N_9808);
or U10090 (N_10090,N_9719,N_9533);
nand U10091 (N_10091,N_9729,N_9788);
nand U10092 (N_10092,N_9876,N_9949);
nor U10093 (N_10093,N_9531,N_9643);
and U10094 (N_10094,N_9593,N_9674);
and U10095 (N_10095,N_9712,N_9505);
nor U10096 (N_10096,N_9893,N_9691);
xnor U10097 (N_10097,N_9708,N_9607);
nand U10098 (N_10098,N_9550,N_9961);
and U10099 (N_10099,N_9964,N_9648);
and U10100 (N_10100,N_9934,N_9796);
xnor U10101 (N_10101,N_9733,N_9991);
xor U10102 (N_10102,N_9624,N_9984);
or U10103 (N_10103,N_9631,N_9831);
nand U10104 (N_10104,N_9825,N_9872);
or U10105 (N_10105,N_9641,N_9759);
or U10106 (N_10106,N_9559,N_9981);
nor U10107 (N_10107,N_9932,N_9552);
xnor U10108 (N_10108,N_9875,N_9904);
or U10109 (N_10109,N_9972,N_9888);
nor U10110 (N_10110,N_9936,N_9529);
nor U10111 (N_10111,N_9632,N_9682);
and U10112 (N_10112,N_9549,N_9752);
or U10113 (N_10113,N_9791,N_9947);
nor U10114 (N_10114,N_9616,N_9588);
or U10115 (N_10115,N_9818,N_9950);
and U10116 (N_10116,N_9771,N_9778);
and U10117 (N_10117,N_9828,N_9640);
xor U10118 (N_10118,N_9908,N_9810);
nor U10119 (N_10119,N_9680,N_9997);
or U10120 (N_10120,N_9718,N_9634);
and U10121 (N_10121,N_9814,N_9783);
or U10122 (N_10122,N_9870,N_9713);
and U10123 (N_10123,N_9673,N_9774);
or U10124 (N_10124,N_9844,N_9970);
or U10125 (N_10125,N_9515,N_9745);
and U10126 (N_10126,N_9863,N_9871);
nand U10127 (N_10127,N_9737,N_9921);
or U10128 (N_10128,N_9839,N_9514);
xnor U10129 (N_10129,N_9703,N_9502);
and U10130 (N_10130,N_9865,N_9711);
nand U10131 (N_10131,N_9993,N_9732);
nand U10132 (N_10132,N_9601,N_9701);
xnor U10133 (N_10133,N_9638,N_9772);
nand U10134 (N_10134,N_9698,N_9988);
and U10135 (N_10135,N_9906,N_9511);
nor U10136 (N_10136,N_9849,N_9945);
and U10137 (N_10137,N_9589,N_9527);
or U10138 (N_10138,N_9802,N_9690);
and U10139 (N_10139,N_9889,N_9918);
nor U10140 (N_10140,N_9606,N_9883);
nor U10141 (N_10141,N_9968,N_9837);
or U10142 (N_10142,N_9826,N_9517);
and U10143 (N_10143,N_9694,N_9941);
xor U10144 (N_10144,N_9882,N_9637);
or U10145 (N_10145,N_9973,N_9554);
or U10146 (N_10146,N_9962,N_9967);
xnor U10147 (N_10147,N_9583,N_9599);
nor U10148 (N_10148,N_9762,N_9948);
or U10149 (N_10149,N_9998,N_9819);
or U10150 (N_10150,N_9891,N_9717);
nor U10151 (N_10151,N_9685,N_9506);
or U10152 (N_10152,N_9913,N_9777);
nand U10153 (N_10153,N_9526,N_9880);
or U10154 (N_10154,N_9925,N_9953);
or U10155 (N_10155,N_9500,N_9784);
nor U10156 (N_10156,N_9735,N_9868);
nor U10157 (N_10157,N_9562,N_9684);
and U10158 (N_10158,N_9611,N_9855);
nand U10159 (N_10159,N_9658,N_9512);
nand U10160 (N_10160,N_9586,N_9927);
nand U10161 (N_10161,N_9545,N_9561);
xnor U10162 (N_10162,N_9940,N_9678);
or U10163 (N_10163,N_9912,N_9700);
xor U10164 (N_10164,N_9695,N_9985);
xor U10165 (N_10165,N_9656,N_9867);
nand U10166 (N_10166,N_9621,N_9996);
nor U10167 (N_10167,N_9966,N_9663);
or U10168 (N_10168,N_9800,N_9905);
or U10169 (N_10169,N_9827,N_9710);
nor U10170 (N_10170,N_9881,N_9537);
nor U10171 (N_10171,N_9922,N_9672);
or U10172 (N_10172,N_9699,N_9721);
nor U10173 (N_10173,N_9629,N_9974);
or U10174 (N_10174,N_9548,N_9995);
nand U10175 (N_10175,N_9722,N_9592);
nand U10176 (N_10176,N_9743,N_9933);
nand U10177 (N_10177,N_9538,N_9675);
nor U10178 (N_10178,N_9986,N_9590);
nand U10179 (N_10179,N_9659,N_9754);
nand U10180 (N_10180,N_9657,N_9873);
xor U10181 (N_10181,N_9899,N_9851);
or U10182 (N_10182,N_9892,N_9798);
nor U10183 (N_10183,N_9509,N_9726);
xnor U10184 (N_10184,N_9688,N_9736);
nor U10185 (N_10185,N_9919,N_9928);
or U10186 (N_10186,N_9740,N_9763);
nand U10187 (N_10187,N_9602,N_9866);
and U10188 (N_10188,N_9528,N_9955);
and U10189 (N_10189,N_9644,N_9553);
xor U10190 (N_10190,N_9510,N_9504);
nor U10191 (N_10191,N_9946,N_9914);
or U10192 (N_10192,N_9692,N_9576);
xnor U10193 (N_10193,N_9793,N_9518);
nor U10194 (N_10194,N_9920,N_9742);
xor U10195 (N_10195,N_9833,N_9760);
or U10196 (N_10196,N_9987,N_9544);
and U10197 (N_10197,N_9969,N_9862);
and U10198 (N_10198,N_9789,N_9805);
xor U10199 (N_10199,N_9570,N_9938);
or U10200 (N_10200,N_9983,N_9896);
and U10201 (N_10201,N_9824,N_9853);
or U10202 (N_10202,N_9957,N_9852);
or U10203 (N_10203,N_9567,N_9910);
nor U10204 (N_10204,N_9755,N_9534);
xor U10205 (N_10205,N_9633,N_9856);
and U10206 (N_10206,N_9619,N_9895);
nand U10207 (N_10207,N_9603,N_9878);
nand U10208 (N_10208,N_9705,N_9989);
nor U10209 (N_10209,N_9523,N_9671);
xnor U10210 (N_10210,N_9761,N_9907);
nand U10211 (N_10211,N_9608,N_9660);
nor U10212 (N_10212,N_9770,N_9649);
nor U10213 (N_10213,N_9555,N_9823);
and U10214 (N_10214,N_9725,N_9630);
nand U10215 (N_10215,N_9503,N_9543);
nor U10216 (N_10216,N_9864,N_9734);
nand U10217 (N_10217,N_9850,N_9843);
nor U10218 (N_10218,N_9775,N_9539);
or U10219 (N_10219,N_9820,N_9848);
nand U10220 (N_10220,N_9806,N_9635);
or U10221 (N_10221,N_9513,N_9951);
and U10222 (N_10222,N_9623,N_9573);
nand U10223 (N_10223,N_9813,N_9702);
nand U10224 (N_10224,N_9886,N_9971);
and U10225 (N_10225,N_9600,N_9817);
nand U10226 (N_10226,N_9697,N_9768);
or U10227 (N_10227,N_9845,N_9585);
xnor U10228 (N_10228,N_9609,N_9612);
xor U10229 (N_10229,N_9801,N_9557);
or U10230 (N_10230,N_9636,N_9716);
or U10231 (N_10231,N_9835,N_9937);
nor U10232 (N_10232,N_9799,N_9898);
and U10233 (N_10233,N_9558,N_9669);
nand U10234 (N_10234,N_9676,N_9571);
or U10235 (N_10235,N_9902,N_9520);
and U10236 (N_10236,N_9626,N_9683);
xnor U10237 (N_10237,N_9591,N_9546);
or U10238 (N_10238,N_9541,N_9841);
or U10239 (N_10239,N_9909,N_9926);
or U10240 (N_10240,N_9903,N_9597);
and U10241 (N_10241,N_9773,N_9911);
nor U10242 (N_10242,N_9613,N_9959);
or U10243 (N_10243,N_9994,N_9677);
nor U10244 (N_10244,N_9568,N_9668);
xor U10245 (N_10245,N_9869,N_9923);
and U10246 (N_10246,N_9748,N_9861);
nand U10247 (N_10247,N_9670,N_9686);
xnor U10248 (N_10248,N_9897,N_9618);
nor U10249 (N_10249,N_9620,N_9707);
nand U10250 (N_10250,N_9918,N_9949);
nor U10251 (N_10251,N_9637,N_9932);
nand U10252 (N_10252,N_9965,N_9802);
xor U10253 (N_10253,N_9644,N_9922);
and U10254 (N_10254,N_9507,N_9810);
nor U10255 (N_10255,N_9938,N_9920);
nor U10256 (N_10256,N_9977,N_9589);
or U10257 (N_10257,N_9719,N_9918);
nor U10258 (N_10258,N_9732,N_9516);
and U10259 (N_10259,N_9626,N_9904);
or U10260 (N_10260,N_9900,N_9767);
nand U10261 (N_10261,N_9538,N_9542);
or U10262 (N_10262,N_9671,N_9988);
and U10263 (N_10263,N_9752,N_9602);
or U10264 (N_10264,N_9629,N_9970);
and U10265 (N_10265,N_9747,N_9596);
or U10266 (N_10266,N_9779,N_9842);
nor U10267 (N_10267,N_9582,N_9733);
nand U10268 (N_10268,N_9581,N_9871);
xnor U10269 (N_10269,N_9956,N_9537);
or U10270 (N_10270,N_9948,N_9832);
nor U10271 (N_10271,N_9521,N_9789);
nor U10272 (N_10272,N_9842,N_9941);
and U10273 (N_10273,N_9883,N_9920);
nor U10274 (N_10274,N_9638,N_9919);
nor U10275 (N_10275,N_9679,N_9502);
or U10276 (N_10276,N_9786,N_9542);
and U10277 (N_10277,N_9592,N_9634);
nor U10278 (N_10278,N_9815,N_9996);
nor U10279 (N_10279,N_9922,N_9871);
or U10280 (N_10280,N_9511,N_9703);
xor U10281 (N_10281,N_9979,N_9628);
and U10282 (N_10282,N_9970,N_9831);
nor U10283 (N_10283,N_9794,N_9663);
nand U10284 (N_10284,N_9923,N_9712);
nor U10285 (N_10285,N_9853,N_9555);
or U10286 (N_10286,N_9649,N_9635);
or U10287 (N_10287,N_9935,N_9565);
and U10288 (N_10288,N_9884,N_9546);
nand U10289 (N_10289,N_9883,N_9610);
nor U10290 (N_10290,N_9948,N_9578);
and U10291 (N_10291,N_9839,N_9987);
xor U10292 (N_10292,N_9993,N_9996);
or U10293 (N_10293,N_9713,N_9552);
nor U10294 (N_10294,N_9739,N_9840);
xor U10295 (N_10295,N_9697,N_9681);
xor U10296 (N_10296,N_9751,N_9974);
and U10297 (N_10297,N_9801,N_9502);
or U10298 (N_10298,N_9874,N_9647);
nand U10299 (N_10299,N_9612,N_9674);
nor U10300 (N_10300,N_9534,N_9847);
or U10301 (N_10301,N_9764,N_9867);
or U10302 (N_10302,N_9746,N_9659);
nand U10303 (N_10303,N_9954,N_9756);
and U10304 (N_10304,N_9558,N_9771);
nor U10305 (N_10305,N_9623,N_9529);
xnor U10306 (N_10306,N_9861,N_9634);
and U10307 (N_10307,N_9986,N_9625);
xor U10308 (N_10308,N_9602,N_9705);
or U10309 (N_10309,N_9750,N_9989);
nand U10310 (N_10310,N_9868,N_9713);
xor U10311 (N_10311,N_9882,N_9578);
nor U10312 (N_10312,N_9973,N_9600);
and U10313 (N_10313,N_9692,N_9885);
nand U10314 (N_10314,N_9733,N_9783);
or U10315 (N_10315,N_9528,N_9782);
or U10316 (N_10316,N_9790,N_9951);
nor U10317 (N_10317,N_9516,N_9535);
nor U10318 (N_10318,N_9894,N_9698);
xor U10319 (N_10319,N_9906,N_9642);
nor U10320 (N_10320,N_9864,N_9625);
nand U10321 (N_10321,N_9766,N_9846);
nor U10322 (N_10322,N_9844,N_9701);
and U10323 (N_10323,N_9789,N_9935);
or U10324 (N_10324,N_9955,N_9984);
xor U10325 (N_10325,N_9607,N_9717);
or U10326 (N_10326,N_9767,N_9796);
nor U10327 (N_10327,N_9523,N_9705);
nand U10328 (N_10328,N_9567,N_9601);
or U10329 (N_10329,N_9526,N_9725);
and U10330 (N_10330,N_9918,N_9556);
xnor U10331 (N_10331,N_9992,N_9716);
or U10332 (N_10332,N_9633,N_9760);
and U10333 (N_10333,N_9723,N_9854);
nand U10334 (N_10334,N_9543,N_9663);
or U10335 (N_10335,N_9715,N_9743);
nor U10336 (N_10336,N_9506,N_9674);
nand U10337 (N_10337,N_9873,N_9774);
and U10338 (N_10338,N_9910,N_9883);
xor U10339 (N_10339,N_9750,N_9975);
or U10340 (N_10340,N_9758,N_9718);
nand U10341 (N_10341,N_9953,N_9992);
or U10342 (N_10342,N_9642,N_9646);
nand U10343 (N_10343,N_9546,N_9859);
xor U10344 (N_10344,N_9688,N_9814);
nor U10345 (N_10345,N_9936,N_9940);
xor U10346 (N_10346,N_9866,N_9723);
and U10347 (N_10347,N_9875,N_9797);
nand U10348 (N_10348,N_9763,N_9682);
or U10349 (N_10349,N_9521,N_9839);
nor U10350 (N_10350,N_9941,N_9662);
nor U10351 (N_10351,N_9669,N_9725);
or U10352 (N_10352,N_9927,N_9530);
xnor U10353 (N_10353,N_9993,N_9678);
and U10354 (N_10354,N_9517,N_9692);
and U10355 (N_10355,N_9701,N_9863);
nand U10356 (N_10356,N_9706,N_9852);
nor U10357 (N_10357,N_9618,N_9744);
nand U10358 (N_10358,N_9513,N_9959);
xor U10359 (N_10359,N_9876,N_9930);
and U10360 (N_10360,N_9553,N_9994);
or U10361 (N_10361,N_9834,N_9580);
nand U10362 (N_10362,N_9579,N_9747);
or U10363 (N_10363,N_9516,N_9888);
and U10364 (N_10364,N_9902,N_9533);
or U10365 (N_10365,N_9613,N_9892);
xor U10366 (N_10366,N_9781,N_9798);
nand U10367 (N_10367,N_9967,N_9656);
nor U10368 (N_10368,N_9843,N_9766);
nand U10369 (N_10369,N_9522,N_9691);
or U10370 (N_10370,N_9617,N_9685);
nand U10371 (N_10371,N_9678,N_9907);
nand U10372 (N_10372,N_9857,N_9961);
xnor U10373 (N_10373,N_9798,N_9729);
xnor U10374 (N_10374,N_9572,N_9710);
and U10375 (N_10375,N_9847,N_9884);
nand U10376 (N_10376,N_9687,N_9545);
or U10377 (N_10377,N_9832,N_9642);
nand U10378 (N_10378,N_9746,N_9604);
or U10379 (N_10379,N_9759,N_9799);
xnor U10380 (N_10380,N_9811,N_9978);
and U10381 (N_10381,N_9537,N_9634);
nand U10382 (N_10382,N_9642,N_9590);
and U10383 (N_10383,N_9951,N_9871);
nand U10384 (N_10384,N_9756,N_9931);
nand U10385 (N_10385,N_9704,N_9780);
nor U10386 (N_10386,N_9868,N_9505);
or U10387 (N_10387,N_9688,N_9565);
or U10388 (N_10388,N_9749,N_9687);
and U10389 (N_10389,N_9624,N_9626);
and U10390 (N_10390,N_9847,N_9971);
and U10391 (N_10391,N_9958,N_9566);
nand U10392 (N_10392,N_9687,N_9602);
nor U10393 (N_10393,N_9760,N_9542);
and U10394 (N_10394,N_9865,N_9808);
nand U10395 (N_10395,N_9981,N_9932);
and U10396 (N_10396,N_9672,N_9604);
and U10397 (N_10397,N_9763,N_9582);
xor U10398 (N_10398,N_9780,N_9709);
or U10399 (N_10399,N_9708,N_9786);
xnor U10400 (N_10400,N_9627,N_9935);
or U10401 (N_10401,N_9728,N_9925);
nor U10402 (N_10402,N_9849,N_9652);
or U10403 (N_10403,N_9981,N_9989);
xor U10404 (N_10404,N_9721,N_9832);
nand U10405 (N_10405,N_9932,N_9668);
nor U10406 (N_10406,N_9820,N_9635);
nand U10407 (N_10407,N_9877,N_9695);
xor U10408 (N_10408,N_9605,N_9502);
and U10409 (N_10409,N_9721,N_9705);
nor U10410 (N_10410,N_9891,N_9887);
nand U10411 (N_10411,N_9658,N_9946);
or U10412 (N_10412,N_9713,N_9918);
nor U10413 (N_10413,N_9874,N_9920);
nor U10414 (N_10414,N_9972,N_9739);
nand U10415 (N_10415,N_9557,N_9646);
and U10416 (N_10416,N_9500,N_9785);
xor U10417 (N_10417,N_9658,N_9626);
or U10418 (N_10418,N_9792,N_9543);
nor U10419 (N_10419,N_9603,N_9651);
and U10420 (N_10420,N_9559,N_9920);
nand U10421 (N_10421,N_9918,N_9914);
xor U10422 (N_10422,N_9934,N_9816);
nor U10423 (N_10423,N_9967,N_9835);
nand U10424 (N_10424,N_9680,N_9954);
and U10425 (N_10425,N_9737,N_9562);
or U10426 (N_10426,N_9797,N_9855);
xnor U10427 (N_10427,N_9785,N_9979);
and U10428 (N_10428,N_9724,N_9850);
and U10429 (N_10429,N_9546,N_9990);
or U10430 (N_10430,N_9608,N_9874);
xnor U10431 (N_10431,N_9922,N_9807);
nand U10432 (N_10432,N_9869,N_9824);
and U10433 (N_10433,N_9569,N_9549);
nor U10434 (N_10434,N_9829,N_9578);
and U10435 (N_10435,N_9633,N_9817);
nor U10436 (N_10436,N_9905,N_9892);
and U10437 (N_10437,N_9696,N_9556);
nand U10438 (N_10438,N_9560,N_9564);
and U10439 (N_10439,N_9739,N_9998);
nand U10440 (N_10440,N_9873,N_9567);
nor U10441 (N_10441,N_9653,N_9796);
nand U10442 (N_10442,N_9795,N_9755);
nor U10443 (N_10443,N_9543,N_9949);
or U10444 (N_10444,N_9670,N_9659);
xnor U10445 (N_10445,N_9711,N_9749);
xnor U10446 (N_10446,N_9585,N_9761);
and U10447 (N_10447,N_9880,N_9517);
nand U10448 (N_10448,N_9914,N_9724);
nand U10449 (N_10449,N_9946,N_9736);
and U10450 (N_10450,N_9583,N_9941);
xnor U10451 (N_10451,N_9823,N_9768);
or U10452 (N_10452,N_9809,N_9558);
nand U10453 (N_10453,N_9596,N_9689);
nor U10454 (N_10454,N_9803,N_9567);
xor U10455 (N_10455,N_9894,N_9744);
xnor U10456 (N_10456,N_9512,N_9616);
nor U10457 (N_10457,N_9527,N_9731);
and U10458 (N_10458,N_9873,N_9628);
nand U10459 (N_10459,N_9738,N_9677);
and U10460 (N_10460,N_9854,N_9772);
and U10461 (N_10461,N_9977,N_9548);
nand U10462 (N_10462,N_9689,N_9659);
and U10463 (N_10463,N_9819,N_9927);
nand U10464 (N_10464,N_9838,N_9794);
xnor U10465 (N_10465,N_9912,N_9696);
xnor U10466 (N_10466,N_9775,N_9776);
nand U10467 (N_10467,N_9599,N_9716);
or U10468 (N_10468,N_9942,N_9545);
or U10469 (N_10469,N_9878,N_9529);
nor U10470 (N_10470,N_9982,N_9694);
xor U10471 (N_10471,N_9515,N_9965);
xnor U10472 (N_10472,N_9794,N_9993);
nor U10473 (N_10473,N_9950,N_9756);
nor U10474 (N_10474,N_9563,N_9525);
xor U10475 (N_10475,N_9784,N_9935);
or U10476 (N_10476,N_9838,N_9886);
xor U10477 (N_10477,N_9716,N_9947);
xor U10478 (N_10478,N_9564,N_9727);
and U10479 (N_10479,N_9815,N_9670);
and U10480 (N_10480,N_9835,N_9798);
nand U10481 (N_10481,N_9541,N_9731);
nand U10482 (N_10482,N_9503,N_9992);
nor U10483 (N_10483,N_9574,N_9749);
xnor U10484 (N_10484,N_9519,N_9939);
and U10485 (N_10485,N_9573,N_9548);
nor U10486 (N_10486,N_9594,N_9716);
xor U10487 (N_10487,N_9619,N_9897);
and U10488 (N_10488,N_9750,N_9999);
and U10489 (N_10489,N_9566,N_9769);
or U10490 (N_10490,N_9768,N_9625);
nor U10491 (N_10491,N_9595,N_9855);
or U10492 (N_10492,N_9695,N_9678);
or U10493 (N_10493,N_9869,N_9952);
and U10494 (N_10494,N_9869,N_9504);
and U10495 (N_10495,N_9934,N_9619);
xor U10496 (N_10496,N_9770,N_9792);
nand U10497 (N_10497,N_9970,N_9897);
or U10498 (N_10498,N_9955,N_9684);
nand U10499 (N_10499,N_9717,N_9969);
and U10500 (N_10500,N_10453,N_10181);
nand U10501 (N_10501,N_10268,N_10248);
and U10502 (N_10502,N_10261,N_10078);
xor U10503 (N_10503,N_10456,N_10118);
or U10504 (N_10504,N_10045,N_10150);
xnor U10505 (N_10505,N_10053,N_10364);
nor U10506 (N_10506,N_10050,N_10164);
or U10507 (N_10507,N_10435,N_10134);
or U10508 (N_10508,N_10486,N_10123);
nor U10509 (N_10509,N_10322,N_10490);
nor U10510 (N_10510,N_10026,N_10067);
and U10511 (N_10511,N_10245,N_10125);
nor U10512 (N_10512,N_10228,N_10104);
or U10513 (N_10513,N_10241,N_10005);
and U10514 (N_10514,N_10001,N_10226);
or U10515 (N_10515,N_10437,N_10004);
and U10516 (N_10516,N_10471,N_10249);
or U10517 (N_10517,N_10039,N_10328);
nand U10518 (N_10518,N_10077,N_10058);
and U10519 (N_10519,N_10069,N_10182);
nor U10520 (N_10520,N_10225,N_10290);
nand U10521 (N_10521,N_10410,N_10270);
or U10522 (N_10522,N_10227,N_10405);
and U10523 (N_10523,N_10217,N_10294);
nor U10524 (N_10524,N_10145,N_10210);
xor U10525 (N_10525,N_10047,N_10339);
nor U10526 (N_10526,N_10133,N_10301);
nand U10527 (N_10527,N_10483,N_10310);
and U10528 (N_10528,N_10113,N_10101);
and U10529 (N_10529,N_10436,N_10326);
or U10530 (N_10530,N_10076,N_10426);
or U10531 (N_10531,N_10422,N_10256);
nand U10532 (N_10532,N_10148,N_10064);
and U10533 (N_10533,N_10363,N_10497);
or U10534 (N_10534,N_10348,N_10461);
or U10535 (N_10535,N_10345,N_10272);
and U10536 (N_10536,N_10494,N_10287);
nand U10537 (N_10537,N_10286,N_10468);
xnor U10538 (N_10538,N_10399,N_10434);
or U10539 (N_10539,N_10025,N_10128);
xnor U10540 (N_10540,N_10127,N_10299);
and U10541 (N_10541,N_10369,N_10475);
nor U10542 (N_10542,N_10155,N_10323);
xnor U10543 (N_10543,N_10280,N_10370);
nand U10544 (N_10544,N_10138,N_10074);
nand U10545 (N_10545,N_10088,N_10242);
nand U10546 (N_10546,N_10353,N_10234);
nor U10547 (N_10547,N_10203,N_10423);
or U10548 (N_10548,N_10395,N_10438);
and U10549 (N_10549,N_10189,N_10303);
nand U10550 (N_10550,N_10376,N_10325);
nand U10551 (N_10551,N_10282,N_10232);
nand U10552 (N_10552,N_10173,N_10485);
nor U10553 (N_10553,N_10159,N_10374);
and U10554 (N_10554,N_10235,N_10034);
nand U10555 (N_10555,N_10116,N_10262);
or U10556 (N_10556,N_10068,N_10072);
xor U10557 (N_10557,N_10147,N_10060);
or U10558 (N_10558,N_10024,N_10265);
or U10559 (N_10559,N_10254,N_10243);
xnor U10560 (N_10560,N_10309,N_10170);
nand U10561 (N_10561,N_10061,N_10362);
xnor U10562 (N_10562,N_10429,N_10425);
and U10563 (N_10563,N_10084,N_10188);
xor U10564 (N_10564,N_10496,N_10073);
and U10565 (N_10565,N_10117,N_10075);
and U10566 (N_10566,N_10216,N_10260);
and U10567 (N_10567,N_10094,N_10334);
nor U10568 (N_10568,N_10336,N_10013);
nor U10569 (N_10569,N_10467,N_10070);
xnor U10570 (N_10570,N_10350,N_10462);
nand U10571 (N_10571,N_10131,N_10152);
nor U10572 (N_10572,N_10421,N_10333);
or U10573 (N_10573,N_10157,N_10106);
or U10574 (N_10574,N_10332,N_10055);
or U10575 (N_10575,N_10038,N_10321);
or U10576 (N_10576,N_10479,N_10126);
nand U10577 (N_10577,N_10132,N_10337);
and U10578 (N_10578,N_10011,N_10139);
or U10579 (N_10579,N_10281,N_10271);
nor U10580 (N_10580,N_10396,N_10361);
and U10581 (N_10581,N_10314,N_10229);
nand U10582 (N_10582,N_10200,N_10211);
xnor U10583 (N_10583,N_10278,N_10107);
nor U10584 (N_10584,N_10377,N_10341);
and U10585 (N_10585,N_10179,N_10031);
and U10586 (N_10586,N_10083,N_10283);
xor U10587 (N_10587,N_10018,N_10239);
nand U10588 (N_10588,N_10177,N_10276);
nand U10589 (N_10589,N_10112,N_10192);
and U10590 (N_10590,N_10029,N_10318);
and U10591 (N_10591,N_10277,N_10447);
nand U10592 (N_10592,N_10207,N_10274);
or U10593 (N_10593,N_10308,N_10111);
nor U10594 (N_10594,N_10092,N_10063);
xnor U10595 (N_10595,N_10266,N_10079);
xnor U10596 (N_10596,N_10080,N_10482);
nor U10597 (N_10597,N_10320,N_10007);
nor U10598 (N_10598,N_10478,N_10454);
nand U10599 (N_10599,N_10315,N_10488);
or U10600 (N_10600,N_10441,N_10338);
nand U10601 (N_10601,N_10205,N_10163);
or U10602 (N_10602,N_10263,N_10154);
or U10603 (N_10603,N_10010,N_10473);
nand U10604 (N_10604,N_10391,N_10160);
nand U10605 (N_10605,N_10097,N_10219);
xor U10606 (N_10606,N_10087,N_10224);
and U10607 (N_10607,N_10199,N_10096);
and U10608 (N_10608,N_10046,N_10411);
xnor U10609 (N_10609,N_10346,N_10371);
nand U10610 (N_10610,N_10122,N_10344);
nand U10611 (N_10611,N_10198,N_10491);
or U10612 (N_10612,N_10440,N_10296);
nor U10613 (N_10613,N_10247,N_10176);
nor U10614 (N_10614,N_10221,N_10174);
nor U10615 (N_10615,N_10431,N_10110);
xor U10616 (N_10616,N_10021,N_10023);
xnor U10617 (N_10617,N_10400,N_10027);
xnor U10618 (N_10618,N_10028,N_10384);
nor U10619 (N_10619,N_10166,N_10347);
or U10620 (N_10620,N_10476,N_10458);
and U10621 (N_10621,N_10383,N_10330);
nor U10622 (N_10622,N_10349,N_10264);
nand U10623 (N_10623,N_10466,N_10051);
nor U10624 (N_10624,N_10140,N_10196);
nand U10625 (N_10625,N_10390,N_10327);
nand U10626 (N_10626,N_10430,N_10091);
and U10627 (N_10627,N_10162,N_10208);
xnor U10628 (N_10628,N_10165,N_10033);
xnor U10629 (N_10629,N_10156,N_10043);
nor U10630 (N_10630,N_10459,N_10136);
nor U10631 (N_10631,N_10288,N_10022);
xnor U10632 (N_10632,N_10420,N_10223);
or U10633 (N_10633,N_10324,N_10187);
xnor U10634 (N_10634,N_10099,N_10387);
and U10635 (N_10635,N_10481,N_10052);
and U10636 (N_10636,N_10042,N_10105);
or U10637 (N_10637,N_10433,N_10115);
nor U10638 (N_10638,N_10428,N_10493);
nand U10639 (N_10639,N_10103,N_10213);
and U10640 (N_10640,N_10404,N_10489);
xor U10641 (N_10641,N_10372,N_10100);
and U10642 (N_10642,N_10062,N_10230);
and U10643 (N_10643,N_10499,N_10427);
or U10644 (N_10644,N_10402,N_10151);
nand U10645 (N_10645,N_10378,N_10257);
or U10646 (N_10646,N_10135,N_10102);
or U10647 (N_10647,N_10124,N_10233);
xor U10648 (N_10648,N_10342,N_10424);
or U10649 (N_10649,N_10175,N_10446);
nand U10650 (N_10650,N_10317,N_10178);
nor U10651 (N_10651,N_10057,N_10474);
nand U10652 (N_10652,N_10495,N_10158);
nand U10653 (N_10653,N_10412,N_10432);
and U10654 (N_10654,N_10195,N_10417);
or U10655 (N_10655,N_10389,N_10300);
nor U10656 (N_10656,N_10109,N_10040);
or U10657 (N_10657,N_10019,N_10359);
or U10658 (N_10658,N_10312,N_10186);
and U10659 (N_10659,N_10204,N_10206);
nand U10660 (N_10660,N_10098,N_10120);
nor U10661 (N_10661,N_10255,N_10222);
or U10662 (N_10662,N_10190,N_10368);
xnor U10663 (N_10663,N_10184,N_10379);
or U10664 (N_10664,N_10403,N_10463);
xnor U10665 (N_10665,N_10215,N_10313);
nand U10666 (N_10666,N_10443,N_10449);
xnor U10667 (N_10667,N_10108,N_10452);
nor U10668 (N_10668,N_10455,N_10385);
nor U10669 (N_10669,N_10008,N_10036);
xor U10670 (N_10670,N_10071,N_10146);
nor U10671 (N_10671,N_10089,N_10161);
or U10672 (N_10672,N_10153,N_10258);
or U10673 (N_10673,N_10457,N_10357);
nand U10674 (N_10674,N_10168,N_10246);
and U10675 (N_10675,N_10450,N_10030);
xnor U10676 (N_10676,N_10044,N_10144);
and U10677 (N_10677,N_10292,N_10451);
xnor U10678 (N_10678,N_10392,N_10017);
xor U10679 (N_10679,N_10366,N_10388);
nor U10680 (N_10680,N_10002,N_10253);
nor U10681 (N_10681,N_10460,N_10056);
or U10682 (N_10682,N_10498,N_10307);
or U10683 (N_10683,N_10143,N_10439);
or U10684 (N_10684,N_10302,N_10329);
nor U10685 (N_10685,N_10259,N_10358);
or U10686 (N_10686,N_10020,N_10408);
nor U10687 (N_10687,N_10464,N_10129);
xnor U10688 (N_10688,N_10335,N_10305);
nand U10689 (N_10689,N_10442,N_10354);
and U10690 (N_10690,N_10201,N_10114);
or U10691 (N_10691,N_10003,N_10037);
or U10692 (N_10692,N_10289,N_10015);
nor U10693 (N_10693,N_10285,N_10236);
or U10694 (N_10694,N_10252,N_10381);
xor U10695 (N_10695,N_10316,N_10373);
nor U10696 (N_10696,N_10293,N_10279);
or U10697 (N_10697,N_10343,N_10016);
nor U10698 (N_10698,N_10000,N_10059);
xnor U10699 (N_10699,N_10086,N_10214);
and U10700 (N_10700,N_10238,N_10130);
and U10701 (N_10701,N_10082,N_10469);
nand U10702 (N_10702,N_10352,N_10269);
nand U10703 (N_10703,N_10418,N_10375);
or U10704 (N_10704,N_10295,N_10209);
or U10705 (N_10705,N_10319,N_10093);
nand U10706 (N_10706,N_10169,N_10291);
nor U10707 (N_10707,N_10304,N_10137);
nand U10708 (N_10708,N_10398,N_10141);
nor U10709 (N_10709,N_10484,N_10477);
xor U10710 (N_10710,N_10194,N_10009);
or U10711 (N_10711,N_10119,N_10171);
xnor U10712 (N_10712,N_10095,N_10251);
nand U10713 (N_10713,N_10448,N_10267);
nand U10714 (N_10714,N_10035,N_10202);
nand U10715 (N_10715,N_10191,N_10185);
or U10716 (N_10716,N_10360,N_10049);
and U10717 (N_10717,N_10014,N_10250);
nand U10718 (N_10718,N_10012,N_10180);
nand U10719 (N_10719,N_10172,N_10480);
nor U10720 (N_10720,N_10142,N_10409);
or U10721 (N_10721,N_10090,N_10197);
and U10722 (N_10722,N_10380,N_10445);
nor U10723 (N_10723,N_10356,N_10394);
and U10724 (N_10724,N_10416,N_10244);
or U10725 (N_10725,N_10183,N_10041);
nor U10726 (N_10726,N_10406,N_10419);
and U10727 (N_10727,N_10351,N_10167);
and U10728 (N_10728,N_10273,N_10470);
xor U10729 (N_10729,N_10212,N_10121);
and U10730 (N_10730,N_10306,N_10085);
and U10731 (N_10731,N_10393,N_10311);
or U10732 (N_10732,N_10444,N_10386);
nor U10733 (N_10733,N_10081,N_10231);
and U10734 (N_10734,N_10218,N_10367);
nor U10735 (N_10735,N_10365,N_10397);
and U10736 (N_10736,N_10149,N_10415);
and U10737 (N_10737,N_10193,N_10340);
or U10738 (N_10738,N_10414,N_10401);
nor U10739 (N_10739,N_10298,N_10472);
and U10740 (N_10740,N_10006,N_10237);
nor U10741 (N_10741,N_10066,N_10407);
nand U10742 (N_10742,N_10355,N_10413);
xor U10743 (N_10743,N_10032,N_10275);
and U10744 (N_10744,N_10331,N_10382);
xor U10745 (N_10745,N_10054,N_10065);
nor U10746 (N_10746,N_10465,N_10048);
or U10747 (N_10747,N_10297,N_10492);
xor U10748 (N_10748,N_10240,N_10220);
and U10749 (N_10749,N_10284,N_10487);
nand U10750 (N_10750,N_10291,N_10397);
or U10751 (N_10751,N_10408,N_10296);
or U10752 (N_10752,N_10298,N_10155);
or U10753 (N_10753,N_10449,N_10240);
xor U10754 (N_10754,N_10239,N_10238);
or U10755 (N_10755,N_10365,N_10314);
or U10756 (N_10756,N_10141,N_10110);
nand U10757 (N_10757,N_10465,N_10100);
or U10758 (N_10758,N_10228,N_10469);
or U10759 (N_10759,N_10062,N_10239);
or U10760 (N_10760,N_10325,N_10101);
nand U10761 (N_10761,N_10170,N_10222);
and U10762 (N_10762,N_10201,N_10216);
xnor U10763 (N_10763,N_10400,N_10355);
nor U10764 (N_10764,N_10020,N_10195);
xnor U10765 (N_10765,N_10383,N_10326);
xnor U10766 (N_10766,N_10031,N_10060);
or U10767 (N_10767,N_10472,N_10327);
xor U10768 (N_10768,N_10388,N_10329);
nor U10769 (N_10769,N_10166,N_10473);
xor U10770 (N_10770,N_10063,N_10252);
nand U10771 (N_10771,N_10052,N_10044);
nor U10772 (N_10772,N_10265,N_10172);
and U10773 (N_10773,N_10486,N_10083);
xor U10774 (N_10774,N_10236,N_10119);
nor U10775 (N_10775,N_10435,N_10344);
or U10776 (N_10776,N_10324,N_10151);
nand U10777 (N_10777,N_10137,N_10161);
xor U10778 (N_10778,N_10232,N_10074);
or U10779 (N_10779,N_10103,N_10494);
nor U10780 (N_10780,N_10049,N_10319);
xor U10781 (N_10781,N_10311,N_10301);
nand U10782 (N_10782,N_10291,N_10133);
or U10783 (N_10783,N_10480,N_10163);
xnor U10784 (N_10784,N_10270,N_10487);
xor U10785 (N_10785,N_10356,N_10171);
nand U10786 (N_10786,N_10305,N_10228);
nor U10787 (N_10787,N_10252,N_10375);
xor U10788 (N_10788,N_10129,N_10224);
nand U10789 (N_10789,N_10462,N_10193);
nor U10790 (N_10790,N_10180,N_10438);
or U10791 (N_10791,N_10353,N_10051);
and U10792 (N_10792,N_10122,N_10255);
nor U10793 (N_10793,N_10001,N_10405);
and U10794 (N_10794,N_10084,N_10075);
and U10795 (N_10795,N_10304,N_10277);
nand U10796 (N_10796,N_10316,N_10390);
and U10797 (N_10797,N_10458,N_10489);
or U10798 (N_10798,N_10023,N_10106);
nand U10799 (N_10799,N_10360,N_10332);
nor U10800 (N_10800,N_10118,N_10238);
and U10801 (N_10801,N_10304,N_10357);
nand U10802 (N_10802,N_10213,N_10480);
nor U10803 (N_10803,N_10129,N_10092);
or U10804 (N_10804,N_10424,N_10498);
and U10805 (N_10805,N_10267,N_10366);
and U10806 (N_10806,N_10002,N_10212);
xnor U10807 (N_10807,N_10232,N_10348);
nor U10808 (N_10808,N_10114,N_10412);
nor U10809 (N_10809,N_10434,N_10350);
and U10810 (N_10810,N_10300,N_10188);
nand U10811 (N_10811,N_10492,N_10462);
xor U10812 (N_10812,N_10235,N_10177);
or U10813 (N_10813,N_10096,N_10236);
nor U10814 (N_10814,N_10080,N_10149);
nand U10815 (N_10815,N_10189,N_10232);
nor U10816 (N_10816,N_10055,N_10416);
or U10817 (N_10817,N_10448,N_10001);
nand U10818 (N_10818,N_10397,N_10091);
or U10819 (N_10819,N_10492,N_10414);
or U10820 (N_10820,N_10287,N_10152);
or U10821 (N_10821,N_10096,N_10223);
xor U10822 (N_10822,N_10413,N_10066);
and U10823 (N_10823,N_10306,N_10125);
nor U10824 (N_10824,N_10186,N_10496);
nor U10825 (N_10825,N_10049,N_10330);
xor U10826 (N_10826,N_10077,N_10363);
or U10827 (N_10827,N_10333,N_10497);
nor U10828 (N_10828,N_10441,N_10328);
nand U10829 (N_10829,N_10085,N_10433);
and U10830 (N_10830,N_10482,N_10235);
nor U10831 (N_10831,N_10247,N_10414);
nand U10832 (N_10832,N_10256,N_10028);
or U10833 (N_10833,N_10222,N_10260);
or U10834 (N_10834,N_10205,N_10013);
nand U10835 (N_10835,N_10022,N_10441);
and U10836 (N_10836,N_10292,N_10211);
nand U10837 (N_10837,N_10112,N_10440);
nor U10838 (N_10838,N_10161,N_10001);
xnor U10839 (N_10839,N_10275,N_10175);
or U10840 (N_10840,N_10473,N_10401);
nor U10841 (N_10841,N_10018,N_10443);
nand U10842 (N_10842,N_10150,N_10484);
xor U10843 (N_10843,N_10204,N_10023);
nor U10844 (N_10844,N_10369,N_10140);
nor U10845 (N_10845,N_10470,N_10367);
and U10846 (N_10846,N_10027,N_10205);
nand U10847 (N_10847,N_10385,N_10104);
xnor U10848 (N_10848,N_10465,N_10417);
and U10849 (N_10849,N_10049,N_10113);
and U10850 (N_10850,N_10002,N_10368);
nand U10851 (N_10851,N_10304,N_10080);
xnor U10852 (N_10852,N_10208,N_10395);
or U10853 (N_10853,N_10050,N_10436);
and U10854 (N_10854,N_10301,N_10235);
nor U10855 (N_10855,N_10470,N_10119);
or U10856 (N_10856,N_10141,N_10225);
and U10857 (N_10857,N_10191,N_10116);
and U10858 (N_10858,N_10129,N_10030);
nand U10859 (N_10859,N_10014,N_10450);
or U10860 (N_10860,N_10031,N_10376);
nor U10861 (N_10861,N_10287,N_10284);
nor U10862 (N_10862,N_10104,N_10077);
xnor U10863 (N_10863,N_10448,N_10044);
nand U10864 (N_10864,N_10231,N_10281);
xor U10865 (N_10865,N_10378,N_10150);
nor U10866 (N_10866,N_10099,N_10060);
nor U10867 (N_10867,N_10372,N_10389);
nor U10868 (N_10868,N_10356,N_10210);
or U10869 (N_10869,N_10111,N_10073);
xnor U10870 (N_10870,N_10410,N_10336);
nand U10871 (N_10871,N_10361,N_10095);
xnor U10872 (N_10872,N_10435,N_10009);
nand U10873 (N_10873,N_10061,N_10429);
or U10874 (N_10874,N_10052,N_10195);
nand U10875 (N_10875,N_10130,N_10435);
and U10876 (N_10876,N_10092,N_10289);
xnor U10877 (N_10877,N_10186,N_10317);
and U10878 (N_10878,N_10078,N_10143);
or U10879 (N_10879,N_10405,N_10383);
xnor U10880 (N_10880,N_10409,N_10367);
nand U10881 (N_10881,N_10276,N_10130);
nand U10882 (N_10882,N_10011,N_10038);
or U10883 (N_10883,N_10323,N_10031);
xnor U10884 (N_10884,N_10154,N_10266);
or U10885 (N_10885,N_10402,N_10310);
nand U10886 (N_10886,N_10445,N_10159);
or U10887 (N_10887,N_10074,N_10451);
and U10888 (N_10888,N_10135,N_10356);
nor U10889 (N_10889,N_10302,N_10145);
and U10890 (N_10890,N_10263,N_10169);
or U10891 (N_10891,N_10078,N_10335);
nor U10892 (N_10892,N_10386,N_10317);
and U10893 (N_10893,N_10341,N_10096);
and U10894 (N_10894,N_10433,N_10050);
nand U10895 (N_10895,N_10320,N_10384);
or U10896 (N_10896,N_10131,N_10255);
and U10897 (N_10897,N_10328,N_10132);
nor U10898 (N_10898,N_10210,N_10168);
xnor U10899 (N_10899,N_10364,N_10331);
or U10900 (N_10900,N_10132,N_10127);
or U10901 (N_10901,N_10261,N_10181);
nand U10902 (N_10902,N_10145,N_10144);
nand U10903 (N_10903,N_10450,N_10156);
or U10904 (N_10904,N_10056,N_10314);
nor U10905 (N_10905,N_10269,N_10040);
nor U10906 (N_10906,N_10204,N_10107);
xnor U10907 (N_10907,N_10092,N_10467);
and U10908 (N_10908,N_10080,N_10184);
nor U10909 (N_10909,N_10188,N_10341);
nor U10910 (N_10910,N_10399,N_10108);
and U10911 (N_10911,N_10323,N_10200);
xnor U10912 (N_10912,N_10258,N_10465);
xnor U10913 (N_10913,N_10286,N_10352);
xnor U10914 (N_10914,N_10385,N_10295);
or U10915 (N_10915,N_10464,N_10377);
xor U10916 (N_10916,N_10483,N_10167);
and U10917 (N_10917,N_10327,N_10383);
and U10918 (N_10918,N_10239,N_10468);
xor U10919 (N_10919,N_10006,N_10357);
nand U10920 (N_10920,N_10188,N_10234);
xor U10921 (N_10921,N_10216,N_10190);
xor U10922 (N_10922,N_10410,N_10368);
nand U10923 (N_10923,N_10303,N_10412);
nor U10924 (N_10924,N_10418,N_10349);
nand U10925 (N_10925,N_10315,N_10303);
and U10926 (N_10926,N_10268,N_10310);
and U10927 (N_10927,N_10440,N_10308);
xnor U10928 (N_10928,N_10474,N_10312);
nand U10929 (N_10929,N_10195,N_10477);
nor U10930 (N_10930,N_10345,N_10088);
and U10931 (N_10931,N_10410,N_10233);
xnor U10932 (N_10932,N_10005,N_10448);
nor U10933 (N_10933,N_10266,N_10093);
xor U10934 (N_10934,N_10315,N_10389);
xnor U10935 (N_10935,N_10218,N_10027);
or U10936 (N_10936,N_10004,N_10397);
xnor U10937 (N_10937,N_10221,N_10234);
and U10938 (N_10938,N_10338,N_10484);
nand U10939 (N_10939,N_10453,N_10214);
or U10940 (N_10940,N_10217,N_10178);
and U10941 (N_10941,N_10185,N_10059);
and U10942 (N_10942,N_10451,N_10290);
xnor U10943 (N_10943,N_10187,N_10380);
and U10944 (N_10944,N_10318,N_10268);
xnor U10945 (N_10945,N_10250,N_10293);
nor U10946 (N_10946,N_10028,N_10213);
nor U10947 (N_10947,N_10229,N_10427);
xor U10948 (N_10948,N_10147,N_10351);
nor U10949 (N_10949,N_10460,N_10483);
or U10950 (N_10950,N_10343,N_10318);
nand U10951 (N_10951,N_10171,N_10191);
nand U10952 (N_10952,N_10471,N_10060);
and U10953 (N_10953,N_10113,N_10190);
and U10954 (N_10954,N_10257,N_10229);
or U10955 (N_10955,N_10019,N_10318);
nor U10956 (N_10956,N_10414,N_10010);
nand U10957 (N_10957,N_10130,N_10240);
and U10958 (N_10958,N_10274,N_10399);
xnor U10959 (N_10959,N_10276,N_10077);
or U10960 (N_10960,N_10494,N_10227);
and U10961 (N_10961,N_10444,N_10081);
and U10962 (N_10962,N_10125,N_10033);
nand U10963 (N_10963,N_10092,N_10427);
or U10964 (N_10964,N_10298,N_10179);
and U10965 (N_10965,N_10349,N_10459);
and U10966 (N_10966,N_10394,N_10386);
xor U10967 (N_10967,N_10266,N_10020);
nor U10968 (N_10968,N_10461,N_10486);
and U10969 (N_10969,N_10377,N_10194);
nor U10970 (N_10970,N_10219,N_10462);
or U10971 (N_10971,N_10170,N_10110);
nor U10972 (N_10972,N_10488,N_10138);
and U10973 (N_10973,N_10490,N_10096);
nor U10974 (N_10974,N_10101,N_10339);
nor U10975 (N_10975,N_10261,N_10073);
nor U10976 (N_10976,N_10376,N_10470);
nand U10977 (N_10977,N_10420,N_10449);
nor U10978 (N_10978,N_10343,N_10495);
nor U10979 (N_10979,N_10240,N_10347);
nor U10980 (N_10980,N_10349,N_10385);
xor U10981 (N_10981,N_10365,N_10153);
and U10982 (N_10982,N_10203,N_10206);
and U10983 (N_10983,N_10129,N_10337);
xnor U10984 (N_10984,N_10001,N_10119);
nand U10985 (N_10985,N_10392,N_10433);
xor U10986 (N_10986,N_10401,N_10370);
or U10987 (N_10987,N_10460,N_10172);
nand U10988 (N_10988,N_10135,N_10409);
nand U10989 (N_10989,N_10268,N_10130);
xor U10990 (N_10990,N_10159,N_10146);
and U10991 (N_10991,N_10011,N_10386);
or U10992 (N_10992,N_10016,N_10240);
nand U10993 (N_10993,N_10102,N_10473);
and U10994 (N_10994,N_10148,N_10428);
xnor U10995 (N_10995,N_10171,N_10248);
or U10996 (N_10996,N_10181,N_10161);
xor U10997 (N_10997,N_10159,N_10415);
nand U10998 (N_10998,N_10186,N_10192);
and U10999 (N_10999,N_10371,N_10120);
or U11000 (N_11000,N_10917,N_10590);
and U11001 (N_11001,N_10663,N_10595);
nand U11002 (N_11002,N_10986,N_10873);
nor U11003 (N_11003,N_10875,N_10627);
and U11004 (N_11004,N_10977,N_10733);
nor U11005 (N_11005,N_10664,N_10912);
nand U11006 (N_11006,N_10589,N_10951);
or U11007 (N_11007,N_10542,N_10800);
or U11008 (N_11008,N_10938,N_10615);
xor U11009 (N_11009,N_10693,N_10673);
and U11010 (N_11010,N_10751,N_10729);
and U11011 (N_11011,N_10620,N_10526);
nor U11012 (N_11012,N_10865,N_10629);
nor U11013 (N_11013,N_10659,N_10703);
nor U11014 (N_11014,N_10959,N_10797);
or U11015 (N_11015,N_10847,N_10810);
nor U11016 (N_11016,N_10695,N_10701);
nand U11017 (N_11017,N_10859,N_10776);
or U11018 (N_11018,N_10990,N_10537);
nor U11019 (N_11019,N_10822,N_10639);
or U11020 (N_11020,N_10655,N_10544);
xor U11021 (N_11021,N_10998,N_10993);
nand U11022 (N_11022,N_10721,N_10521);
and U11023 (N_11023,N_10906,N_10928);
and U11024 (N_11024,N_10999,N_10881);
and U11025 (N_11025,N_10517,N_10607);
and U11026 (N_11026,N_10849,N_10559);
and U11027 (N_11027,N_10706,N_10550);
nor U11028 (N_11028,N_10638,N_10562);
and U11029 (N_11029,N_10569,N_10669);
and U11030 (N_11030,N_10891,N_10884);
or U11031 (N_11031,N_10918,N_10713);
or U11032 (N_11032,N_10778,N_10687);
and U11033 (N_11033,N_10931,N_10968);
xnor U11034 (N_11034,N_10842,N_10960);
nor U11035 (N_11035,N_10806,N_10716);
nand U11036 (N_11036,N_10512,N_10668);
or U11037 (N_11037,N_10909,N_10755);
or U11038 (N_11038,N_10586,N_10584);
and U11039 (N_11039,N_10719,N_10743);
nor U11040 (N_11040,N_10717,N_10600);
nor U11041 (N_11041,N_10844,N_10789);
or U11042 (N_11042,N_10553,N_10958);
nand U11043 (N_11043,N_10576,N_10956);
xnor U11044 (N_11044,N_10840,N_10837);
nand U11045 (N_11045,N_10506,N_10823);
nand U11046 (N_11046,N_10710,N_10670);
nor U11047 (N_11047,N_10532,N_10853);
and U11048 (N_11048,N_10893,N_10563);
nand U11049 (N_11049,N_10608,N_10967);
nand U11050 (N_11050,N_10786,N_10579);
or U11051 (N_11051,N_10969,N_10798);
or U11052 (N_11052,N_10558,N_10879);
nand U11053 (N_11053,N_10626,N_10886);
nor U11054 (N_11054,N_10676,N_10541);
nand U11055 (N_11055,N_10878,N_10841);
nor U11056 (N_11056,N_10753,N_10543);
nand U11057 (N_11057,N_10646,N_10782);
or U11058 (N_11058,N_10792,N_10732);
nand U11059 (N_11059,N_10949,N_10851);
and U11060 (N_11060,N_10632,N_10516);
or U11061 (N_11061,N_10804,N_10895);
and U11062 (N_11062,N_10779,N_10930);
and U11063 (N_11063,N_10916,N_10650);
or U11064 (N_11064,N_10870,N_10882);
or U11065 (N_11065,N_10821,N_10988);
and U11066 (N_11066,N_10692,N_10981);
and U11067 (N_11067,N_10833,N_10599);
or U11068 (N_11068,N_10637,N_10850);
nand U11069 (N_11069,N_10604,N_10987);
nand U11070 (N_11070,N_10829,N_10667);
or U11071 (N_11071,N_10505,N_10739);
nor U11072 (N_11072,N_10963,N_10920);
xor U11073 (N_11073,N_10784,N_10771);
and U11074 (N_11074,N_10805,N_10927);
and U11075 (N_11075,N_10940,N_10587);
nor U11076 (N_11076,N_10921,N_10514);
and U11077 (N_11077,N_10766,N_10913);
nor U11078 (N_11078,N_10557,N_10690);
or U11079 (N_11079,N_10534,N_10594);
xor U11080 (N_11080,N_10621,N_10643);
xnor U11081 (N_11081,N_10826,N_10527);
nand U11082 (N_11082,N_10601,N_10531);
nor U11083 (N_11083,N_10674,N_10660);
nor U11084 (N_11084,N_10711,N_10747);
or U11085 (N_11085,N_10919,N_10737);
nand U11086 (N_11086,N_10677,N_10817);
nand U11087 (N_11087,N_10568,N_10902);
nor U11088 (N_11088,N_10666,N_10880);
or U11089 (N_11089,N_10972,N_10509);
nand U11090 (N_11090,N_10838,N_10502);
xor U11091 (N_11091,N_10709,N_10872);
nor U11092 (N_11092,N_10973,N_10769);
xor U11093 (N_11093,N_10754,N_10799);
nor U11094 (N_11094,N_10606,N_10802);
and U11095 (N_11095,N_10540,N_10768);
nand U11096 (N_11096,N_10858,N_10862);
nand U11097 (N_11097,N_10807,N_10845);
or U11098 (N_11098,N_10633,N_10742);
and U11099 (N_11099,N_10860,N_10508);
xnor U11100 (N_11100,N_10665,N_10547);
xnor U11101 (N_11101,N_10749,N_10520);
xor U11102 (N_11102,N_10610,N_10926);
nand U11103 (N_11103,N_10937,N_10911);
and U11104 (N_11104,N_10561,N_10812);
nand U11105 (N_11105,N_10657,N_10803);
and U11106 (N_11106,N_10834,N_10658);
and U11107 (N_11107,N_10975,N_10852);
and U11108 (N_11108,N_10612,N_10795);
or U11109 (N_11109,N_10761,N_10583);
and U11110 (N_11110,N_10535,N_10623);
or U11111 (N_11111,N_10772,N_10560);
or U11112 (N_11112,N_10714,N_10922);
or U11113 (N_11113,N_10647,N_10924);
nor U11114 (N_11114,N_10500,N_10868);
and U11115 (N_11115,N_10794,N_10996);
xor U11116 (N_11116,N_10764,N_10548);
xnor U11117 (N_11117,N_10876,N_10574);
and U11118 (N_11118,N_10635,N_10915);
and U11119 (N_11119,N_10861,N_10935);
or U11120 (N_11120,N_10740,N_10580);
xnor U11121 (N_11121,N_10943,N_10970);
and U11122 (N_11122,N_10741,N_10757);
or U11123 (N_11123,N_10581,N_10582);
nor U11124 (N_11124,N_10890,N_10735);
xnor U11125 (N_11125,N_10671,N_10984);
nand U11126 (N_11126,N_10536,N_10760);
xor U11127 (N_11127,N_10899,N_10628);
or U11128 (N_11128,N_10715,N_10939);
nor U11129 (N_11129,N_10783,N_10832);
nor U11130 (N_11130,N_10510,N_10596);
nor U11131 (N_11131,N_10672,N_10642);
nor U11132 (N_11132,N_10730,N_10555);
and U11133 (N_11133,N_10898,N_10831);
nor U11134 (N_11134,N_10791,N_10578);
and U11135 (N_11135,N_10796,N_10820);
nor U11136 (N_11136,N_10903,N_10572);
nor U11137 (N_11137,N_10933,N_10896);
nor U11138 (N_11138,N_10728,N_10780);
xor U11139 (N_11139,N_10945,N_10857);
xnor U11140 (N_11140,N_10910,N_10905);
nor U11141 (N_11141,N_10866,N_10570);
nor U11142 (N_11142,N_10696,N_10689);
nand U11143 (N_11143,N_10538,N_10961);
nand U11144 (N_11144,N_10759,N_10965);
nor U11145 (N_11145,N_10523,N_10630);
or U11146 (N_11146,N_10507,N_10700);
nand U11147 (N_11147,N_10839,N_10885);
and U11148 (N_11148,N_10974,N_10681);
xnor U11149 (N_11149,N_10588,N_10685);
or U11150 (N_11150,N_10904,N_10835);
nor U11151 (N_11151,N_10707,N_10785);
or U11152 (N_11152,N_10734,N_10781);
or U11153 (N_11153,N_10932,N_10722);
nand U11154 (N_11154,N_10679,N_10763);
nand U11155 (N_11155,N_10793,N_10593);
nor U11156 (N_11156,N_10976,N_10554);
and U11157 (N_11157,N_10750,N_10702);
or U11158 (N_11158,N_10614,N_10954);
and U11159 (N_11159,N_10925,N_10640);
and U11160 (N_11160,N_10929,N_10952);
and U11161 (N_11161,N_10966,N_10950);
or U11162 (N_11162,N_10624,N_10819);
and U11163 (N_11163,N_10565,N_10566);
and U11164 (N_11164,N_10644,N_10723);
and U11165 (N_11165,N_10756,N_10592);
nor U11166 (N_11166,N_10573,N_10818);
or U11167 (N_11167,N_10649,N_10744);
xnor U11168 (N_11168,N_10983,N_10546);
and U11169 (N_11169,N_10641,N_10848);
nand U11170 (N_11170,N_10946,N_10874);
nor U11171 (N_11171,N_10712,N_10801);
xor U11172 (N_11172,N_10994,N_10603);
or U11173 (N_11173,N_10697,N_10788);
or U11174 (N_11174,N_10651,N_10653);
and U11175 (N_11175,N_10864,N_10634);
and U11176 (N_11176,N_10656,N_10767);
and U11177 (N_11177,N_10830,N_10907);
and U11178 (N_11178,N_10883,N_10513);
or U11179 (N_11179,N_10511,N_10605);
or U11180 (N_11180,N_10813,N_10869);
nor U11181 (N_11181,N_10871,N_10773);
or U11182 (N_11182,N_10518,N_10980);
xnor U11183 (N_11183,N_10765,N_10724);
and U11184 (N_11184,N_10900,N_10979);
or U11185 (N_11185,N_10908,N_10611);
nor U11186 (N_11186,N_10694,N_10602);
nor U11187 (N_11187,N_10856,N_10691);
or U11188 (N_11188,N_10752,N_10887);
nor U11189 (N_11189,N_10914,N_10775);
nand U11190 (N_11190,N_10901,N_10552);
and U11191 (N_11191,N_10556,N_10816);
or U11192 (N_11192,N_10585,N_10597);
nor U11193 (N_11193,N_10867,N_10727);
nand U11194 (N_11194,N_10698,N_10825);
or U11195 (N_11195,N_10982,N_10877);
or U11196 (N_11196,N_10654,N_10613);
nand U11197 (N_11197,N_10636,N_10738);
or U11198 (N_11198,N_10591,N_10824);
nor U11199 (N_11199,N_10827,N_10894);
or U11200 (N_11200,N_10675,N_10957);
xor U11201 (N_11201,N_10846,N_10811);
or U11202 (N_11202,N_10575,N_10888);
and U11203 (N_11203,N_10704,N_10854);
nand U11204 (N_11204,N_10662,N_10515);
nand U11205 (N_11205,N_10731,N_10758);
and U11206 (N_11206,N_10863,N_10787);
xnor U11207 (N_11207,N_10619,N_10616);
nor U11208 (N_11208,N_10964,N_10809);
nor U11209 (N_11209,N_10577,N_10989);
and U11210 (N_11210,N_10680,N_10618);
xor U11211 (N_11211,N_10678,N_10631);
nand U11212 (N_11212,N_10528,N_10997);
or U11213 (N_11213,N_10814,N_10748);
xor U11214 (N_11214,N_10501,N_10828);
nand U11215 (N_11215,N_10746,N_10683);
nand U11216 (N_11216,N_10762,N_10843);
and U11217 (N_11217,N_10522,N_10533);
or U11218 (N_11218,N_10971,N_10539);
and U11219 (N_11219,N_10567,N_10718);
nand U11220 (N_11220,N_10889,N_10944);
or U11221 (N_11221,N_10530,N_10705);
or U11222 (N_11222,N_10625,N_10726);
or U11223 (N_11223,N_10948,N_10836);
xnor U11224 (N_11224,N_10770,N_10529);
and U11225 (N_11225,N_10725,N_10923);
xor U11226 (N_11226,N_10519,N_10897);
nand U11227 (N_11227,N_10564,N_10985);
nor U11228 (N_11228,N_10942,N_10609);
nor U11229 (N_11229,N_10688,N_10953);
xnor U11230 (N_11230,N_10661,N_10598);
and U11231 (N_11231,N_10524,N_10684);
nand U11232 (N_11232,N_10777,N_10790);
or U11233 (N_11233,N_10545,N_10892);
xor U11234 (N_11234,N_10936,N_10622);
xor U11235 (N_11235,N_10686,N_10549);
nor U11236 (N_11236,N_10682,N_10855);
xnor U11237 (N_11237,N_10720,N_10617);
or U11238 (N_11238,N_10947,N_10815);
or U11239 (N_11239,N_10736,N_10525);
xor U11240 (N_11240,N_10551,N_10503);
and U11241 (N_11241,N_10962,N_10774);
and U11242 (N_11242,N_10995,N_10504);
nand U11243 (N_11243,N_10934,N_10708);
xor U11244 (N_11244,N_10992,N_10652);
nor U11245 (N_11245,N_10808,N_10645);
or U11246 (N_11246,N_10978,N_10745);
nor U11247 (N_11247,N_10571,N_10648);
nand U11248 (N_11248,N_10991,N_10941);
nor U11249 (N_11249,N_10699,N_10955);
or U11250 (N_11250,N_10750,N_10657);
or U11251 (N_11251,N_10771,N_10597);
nor U11252 (N_11252,N_10901,N_10898);
or U11253 (N_11253,N_10737,N_10753);
nand U11254 (N_11254,N_10871,N_10956);
nor U11255 (N_11255,N_10531,N_10735);
xnor U11256 (N_11256,N_10568,N_10646);
and U11257 (N_11257,N_10598,N_10558);
nor U11258 (N_11258,N_10961,N_10602);
nand U11259 (N_11259,N_10976,N_10923);
nor U11260 (N_11260,N_10565,N_10558);
and U11261 (N_11261,N_10843,N_10898);
or U11262 (N_11262,N_10917,N_10843);
nand U11263 (N_11263,N_10559,N_10734);
nor U11264 (N_11264,N_10956,N_10850);
and U11265 (N_11265,N_10984,N_10700);
nor U11266 (N_11266,N_10944,N_10600);
or U11267 (N_11267,N_10937,N_10821);
nor U11268 (N_11268,N_10756,N_10956);
nor U11269 (N_11269,N_10526,N_10802);
and U11270 (N_11270,N_10957,N_10763);
xor U11271 (N_11271,N_10804,N_10997);
nor U11272 (N_11272,N_10692,N_10509);
or U11273 (N_11273,N_10618,N_10711);
and U11274 (N_11274,N_10808,N_10852);
nand U11275 (N_11275,N_10868,N_10581);
nor U11276 (N_11276,N_10509,N_10995);
xnor U11277 (N_11277,N_10821,N_10910);
or U11278 (N_11278,N_10500,N_10789);
nand U11279 (N_11279,N_10773,N_10751);
xnor U11280 (N_11280,N_10933,N_10826);
nor U11281 (N_11281,N_10916,N_10893);
and U11282 (N_11282,N_10782,N_10596);
and U11283 (N_11283,N_10871,N_10901);
or U11284 (N_11284,N_10616,N_10632);
and U11285 (N_11285,N_10719,N_10841);
nor U11286 (N_11286,N_10779,N_10955);
and U11287 (N_11287,N_10765,N_10910);
xor U11288 (N_11288,N_10878,N_10654);
xor U11289 (N_11289,N_10867,N_10940);
nand U11290 (N_11290,N_10613,N_10937);
or U11291 (N_11291,N_10519,N_10893);
or U11292 (N_11292,N_10701,N_10955);
nand U11293 (N_11293,N_10736,N_10512);
nand U11294 (N_11294,N_10734,N_10949);
and U11295 (N_11295,N_10972,N_10786);
xor U11296 (N_11296,N_10994,N_10821);
nor U11297 (N_11297,N_10913,N_10529);
nand U11298 (N_11298,N_10780,N_10867);
and U11299 (N_11299,N_10647,N_10767);
nand U11300 (N_11300,N_10917,N_10962);
nor U11301 (N_11301,N_10752,N_10797);
xor U11302 (N_11302,N_10930,N_10971);
xnor U11303 (N_11303,N_10653,N_10656);
nor U11304 (N_11304,N_10782,N_10643);
or U11305 (N_11305,N_10844,N_10673);
xnor U11306 (N_11306,N_10809,N_10649);
and U11307 (N_11307,N_10739,N_10798);
nand U11308 (N_11308,N_10867,N_10872);
nand U11309 (N_11309,N_10580,N_10948);
or U11310 (N_11310,N_10870,N_10707);
xnor U11311 (N_11311,N_10931,N_10689);
xor U11312 (N_11312,N_10786,N_10777);
xor U11313 (N_11313,N_10555,N_10674);
nand U11314 (N_11314,N_10913,N_10571);
or U11315 (N_11315,N_10546,N_10667);
nand U11316 (N_11316,N_10750,N_10796);
or U11317 (N_11317,N_10784,N_10952);
or U11318 (N_11318,N_10901,N_10870);
and U11319 (N_11319,N_10585,N_10518);
and U11320 (N_11320,N_10883,N_10598);
xnor U11321 (N_11321,N_10635,N_10522);
xor U11322 (N_11322,N_10999,N_10972);
nand U11323 (N_11323,N_10527,N_10540);
nor U11324 (N_11324,N_10557,N_10524);
or U11325 (N_11325,N_10526,N_10551);
nor U11326 (N_11326,N_10953,N_10940);
nor U11327 (N_11327,N_10623,N_10992);
nor U11328 (N_11328,N_10669,N_10719);
nor U11329 (N_11329,N_10551,N_10931);
nor U11330 (N_11330,N_10549,N_10856);
xnor U11331 (N_11331,N_10668,N_10684);
or U11332 (N_11332,N_10892,N_10872);
or U11333 (N_11333,N_10700,N_10520);
nor U11334 (N_11334,N_10801,N_10600);
or U11335 (N_11335,N_10967,N_10729);
nand U11336 (N_11336,N_10818,N_10874);
xor U11337 (N_11337,N_10878,N_10928);
and U11338 (N_11338,N_10514,N_10731);
nor U11339 (N_11339,N_10966,N_10512);
xor U11340 (N_11340,N_10966,N_10792);
and U11341 (N_11341,N_10711,N_10716);
nor U11342 (N_11342,N_10924,N_10695);
nor U11343 (N_11343,N_10637,N_10625);
nand U11344 (N_11344,N_10833,N_10517);
and U11345 (N_11345,N_10736,N_10674);
or U11346 (N_11346,N_10790,N_10766);
nor U11347 (N_11347,N_10608,N_10556);
nor U11348 (N_11348,N_10604,N_10648);
and U11349 (N_11349,N_10954,N_10887);
nand U11350 (N_11350,N_10551,N_10923);
xor U11351 (N_11351,N_10525,N_10562);
xnor U11352 (N_11352,N_10604,N_10672);
or U11353 (N_11353,N_10940,N_10808);
or U11354 (N_11354,N_10677,N_10748);
nor U11355 (N_11355,N_10731,N_10692);
and U11356 (N_11356,N_10548,N_10547);
or U11357 (N_11357,N_10733,N_10743);
nand U11358 (N_11358,N_10985,N_10948);
xor U11359 (N_11359,N_10971,N_10615);
and U11360 (N_11360,N_10579,N_10715);
nor U11361 (N_11361,N_10587,N_10677);
nand U11362 (N_11362,N_10542,N_10617);
nor U11363 (N_11363,N_10994,N_10733);
nor U11364 (N_11364,N_10723,N_10898);
or U11365 (N_11365,N_10671,N_10768);
nor U11366 (N_11366,N_10634,N_10554);
nand U11367 (N_11367,N_10866,N_10629);
and U11368 (N_11368,N_10565,N_10548);
xnor U11369 (N_11369,N_10750,N_10835);
and U11370 (N_11370,N_10503,N_10907);
and U11371 (N_11371,N_10730,N_10543);
nor U11372 (N_11372,N_10862,N_10505);
xor U11373 (N_11373,N_10574,N_10673);
nand U11374 (N_11374,N_10716,N_10883);
or U11375 (N_11375,N_10969,N_10749);
or U11376 (N_11376,N_10804,N_10999);
or U11377 (N_11377,N_10596,N_10519);
or U11378 (N_11378,N_10713,N_10939);
and U11379 (N_11379,N_10724,N_10981);
nor U11380 (N_11380,N_10945,N_10557);
xor U11381 (N_11381,N_10618,N_10755);
or U11382 (N_11382,N_10915,N_10808);
or U11383 (N_11383,N_10989,N_10840);
xnor U11384 (N_11384,N_10971,N_10853);
and U11385 (N_11385,N_10885,N_10683);
nand U11386 (N_11386,N_10727,N_10764);
and U11387 (N_11387,N_10702,N_10822);
xor U11388 (N_11388,N_10633,N_10640);
xor U11389 (N_11389,N_10537,N_10726);
xor U11390 (N_11390,N_10560,N_10683);
nor U11391 (N_11391,N_10631,N_10715);
and U11392 (N_11392,N_10996,N_10760);
nor U11393 (N_11393,N_10648,N_10708);
and U11394 (N_11394,N_10523,N_10850);
nor U11395 (N_11395,N_10607,N_10614);
and U11396 (N_11396,N_10568,N_10860);
and U11397 (N_11397,N_10506,N_10536);
xor U11398 (N_11398,N_10947,N_10643);
or U11399 (N_11399,N_10702,N_10607);
or U11400 (N_11400,N_10553,N_10790);
nor U11401 (N_11401,N_10884,N_10646);
nor U11402 (N_11402,N_10608,N_10712);
xnor U11403 (N_11403,N_10588,N_10533);
xnor U11404 (N_11404,N_10934,N_10809);
or U11405 (N_11405,N_10765,N_10680);
and U11406 (N_11406,N_10640,N_10606);
xnor U11407 (N_11407,N_10700,N_10872);
nand U11408 (N_11408,N_10652,N_10599);
nor U11409 (N_11409,N_10698,N_10689);
nor U11410 (N_11410,N_10546,N_10683);
and U11411 (N_11411,N_10718,N_10527);
xnor U11412 (N_11412,N_10937,N_10575);
or U11413 (N_11413,N_10995,N_10932);
nor U11414 (N_11414,N_10791,N_10672);
or U11415 (N_11415,N_10883,N_10848);
nand U11416 (N_11416,N_10908,N_10982);
nor U11417 (N_11417,N_10903,N_10704);
xor U11418 (N_11418,N_10538,N_10573);
or U11419 (N_11419,N_10681,N_10871);
and U11420 (N_11420,N_10537,N_10529);
nand U11421 (N_11421,N_10866,N_10795);
or U11422 (N_11422,N_10682,N_10642);
and U11423 (N_11423,N_10672,N_10961);
xor U11424 (N_11424,N_10985,N_10707);
xor U11425 (N_11425,N_10833,N_10525);
xnor U11426 (N_11426,N_10728,N_10891);
and U11427 (N_11427,N_10680,N_10999);
nor U11428 (N_11428,N_10589,N_10528);
or U11429 (N_11429,N_10580,N_10810);
or U11430 (N_11430,N_10824,N_10769);
or U11431 (N_11431,N_10753,N_10931);
nor U11432 (N_11432,N_10864,N_10632);
or U11433 (N_11433,N_10993,N_10627);
xor U11434 (N_11434,N_10601,N_10709);
nor U11435 (N_11435,N_10833,N_10559);
nand U11436 (N_11436,N_10794,N_10901);
xor U11437 (N_11437,N_10740,N_10985);
xnor U11438 (N_11438,N_10938,N_10591);
or U11439 (N_11439,N_10684,N_10549);
xor U11440 (N_11440,N_10557,N_10507);
or U11441 (N_11441,N_10629,N_10555);
or U11442 (N_11442,N_10592,N_10810);
nor U11443 (N_11443,N_10967,N_10794);
or U11444 (N_11444,N_10930,N_10577);
xor U11445 (N_11445,N_10824,N_10569);
nand U11446 (N_11446,N_10953,N_10856);
nor U11447 (N_11447,N_10844,N_10857);
or U11448 (N_11448,N_10626,N_10571);
and U11449 (N_11449,N_10627,N_10570);
nand U11450 (N_11450,N_10548,N_10719);
nor U11451 (N_11451,N_10857,N_10579);
nor U11452 (N_11452,N_10726,N_10744);
xor U11453 (N_11453,N_10960,N_10713);
or U11454 (N_11454,N_10723,N_10614);
nand U11455 (N_11455,N_10611,N_10595);
nor U11456 (N_11456,N_10562,N_10595);
xor U11457 (N_11457,N_10876,N_10614);
nor U11458 (N_11458,N_10595,N_10638);
and U11459 (N_11459,N_10712,N_10862);
nand U11460 (N_11460,N_10501,N_10854);
and U11461 (N_11461,N_10707,N_10571);
or U11462 (N_11462,N_10926,N_10615);
nor U11463 (N_11463,N_10755,N_10597);
nor U11464 (N_11464,N_10520,N_10880);
or U11465 (N_11465,N_10802,N_10930);
xor U11466 (N_11466,N_10950,N_10795);
nand U11467 (N_11467,N_10537,N_10985);
and U11468 (N_11468,N_10650,N_10597);
nor U11469 (N_11469,N_10537,N_10745);
and U11470 (N_11470,N_10540,N_10785);
nand U11471 (N_11471,N_10819,N_10812);
nand U11472 (N_11472,N_10986,N_10536);
nand U11473 (N_11473,N_10547,N_10763);
and U11474 (N_11474,N_10786,N_10616);
or U11475 (N_11475,N_10735,N_10972);
or U11476 (N_11476,N_10669,N_10871);
xnor U11477 (N_11477,N_10532,N_10819);
and U11478 (N_11478,N_10889,N_10756);
or U11479 (N_11479,N_10822,N_10839);
nor U11480 (N_11480,N_10556,N_10794);
nor U11481 (N_11481,N_10974,N_10742);
or U11482 (N_11482,N_10756,N_10788);
xnor U11483 (N_11483,N_10533,N_10660);
nor U11484 (N_11484,N_10904,N_10804);
nor U11485 (N_11485,N_10775,N_10677);
xnor U11486 (N_11486,N_10802,N_10942);
xor U11487 (N_11487,N_10613,N_10876);
xor U11488 (N_11488,N_10898,N_10938);
nand U11489 (N_11489,N_10918,N_10679);
nand U11490 (N_11490,N_10866,N_10641);
xnor U11491 (N_11491,N_10712,N_10749);
and U11492 (N_11492,N_10798,N_10986);
and U11493 (N_11493,N_10534,N_10807);
or U11494 (N_11494,N_10522,N_10574);
or U11495 (N_11495,N_10584,N_10691);
and U11496 (N_11496,N_10816,N_10743);
xnor U11497 (N_11497,N_10748,N_10693);
nand U11498 (N_11498,N_10982,N_10800);
and U11499 (N_11499,N_10844,N_10585);
and U11500 (N_11500,N_11128,N_11305);
nor U11501 (N_11501,N_11320,N_11220);
xnor U11502 (N_11502,N_11308,N_11322);
xor U11503 (N_11503,N_11031,N_11164);
or U11504 (N_11504,N_11117,N_11450);
xnor U11505 (N_11505,N_11468,N_11261);
xnor U11506 (N_11506,N_11297,N_11073);
nor U11507 (N_11507,N_11478,N_11165);
nand U11508 (N_11508,N_11173,N_11339);
and U11509 (N_11509,N_11303,N_11086);
nor U11510 (N_11510,N_11172,N_11343);
or U11511 (N_11511,N_11421,N_11074);
nor U11512 (N_11512,N_11020,N_11292);
and U11513 (N_11513,N_11205,N_11215);
or U11514 (N_11514,N_11347,N_11247);
nor U11515 (N_11515,N_11229,N_11077);
and U11516 (N_11516,N_11467,N_11334);
and U11517 (N_11517,N_11231,N_11064);
and U11518 (N_11518,N_11439,N_11009);
nand U11519 (N_11519,N_11350,N_11483);
nor U11520 (N_11520,N_11492,N_11272);
or U11521 (N_11521,N_11402,N_11342);
nor U11522 (N_11522,N_11245,N_11039);
nand U11523 (N_11523,N_11241,N_11239);
or U11524 (N_11524,N_11223,N_11484);
or U11525 (N_11525,N_11444,N_11338);
nand U11526 (N_11526,N_11148,N_11130);
and U11527 (N_11527,N_11146,N_11499);
nor U11528 (N_11528,N_11163,N_11049);
nor U11529 (N_11529,N_11357,N_11430);
nor U11530 (N_11530,N_11482,N_11313);
nor U11531 (N_11531,N_11095,N_11488);
nor U11532 (N_11532,N_11063,N_11273);
and U11533 (N_11533,N_11192,N_11257);
nand U11534 (N_11534,N_11038,N_11050);
nor U11535 (N_11535,N_11109,N_11202);
xnor U11536 (N_11536,N_11377,N_11393);
or U11537 (N_11537,N_11236,N_11329);
or U11538 (N_11538,N_11000,N_11454);
nor U11539 (N_11539,N_11358,N_11304);
and U11540 (N_11540,N_11395,N_11010);
and U11541 (N_11541,N_11465,N_11435);
or U11542 (N_11542,N_11157,N_11264);
or U11543 (N_11543,N_11364,N_11124);
nor U11544 (N_11544,N_11005,N_11214);
nor U11545 (N_11545,N_11296,N_11246);
and U11546 (N_11546,N_11285,N_11251);
and U11547 (N_11547,N_11453,N_11354);
xor U11548 (N_11548,N_11081,N_11084);
and U11549 (N_11549,N_11066,N_11025);
or U11550 (N_11550,N_11113,N_11036);
and U11551 (N_11551,N_11254,N_11378);
nand U11552 (N_11552,N_11155,N_11211);
and U11553 (N_11553,N_11082,N_11045);
nand U11554 (N_11554,N_11166,N_11083);
or U11555 (N_11555,N_11438,N_11479);
nand U11556 (N_11556,N_11381,N_11356);
nand U11557 (N_11557,N_11470,N_11122);
nor U11558 (N_11558,N_11434,N_11300);
nand U11559 (N_11559,N_11366,N_11121);
or U11560 (N_11560,N_11286,N_11062);
xor U11561 (N_11561,N_11359,N_11144);
nand U11562 (N_11562,N_11388,N_11051);
or U11563 (N_11563,N_11376,N_11089);
nor U11564 (N_11564,N_11351,N_11409);
nand U11565 (N_11565,N_11447,N_11400);
or U11566 (N_11566,N_11262,N_11266);
xnor U11567 (N_11567,N_11107,N_11387);
nor U11568 (N_11568,N_11311,N_11398);
and U11569 (N_11569,N_11382,N_11332);
nand U11570 (N_11570,N_11288,N_11440);
nor U11571 (N_11571,N_11373,N_11348);
or U11572 (N_11572,N_11149,N_11412);
or U11573 (N_11573,N_11419,N_11294);
nand U11574 (N_11574,N_11495,N_11093);
or U11575 (N_11575,N_11287,N_11100);
and U11576 (N_11576,N_11227,N_11056);
xnor U11577 (N_11577,N_11424,N_11379);
nand U11578 (N_11578,N_11460,N_11139);
nand U11579 (N_11579,N_11088,N_11368);
and U11580 (N_11580,N_11167,N_11471);
xor U11581 (N_11581,N_11252,N_11110);
or U11582 (N_11582,N_11306,N_11250);
xnor U11583 (N_11583,N_11029,N_11386);
nor U11584 (N_11584,N_11325,N_11337);
nor U11585 (N_11585,N_11277,N_11458);
or U11586 (N_11586,N_11037,N_11333);
or U11587 (N_11587,N_11457,N_11293);
and U11588 (N_11588,N_11047,N_11417);
nor U11589 (N_11589,N_11098,N_11452);
xor U11590 (N_11590,N_11437,N_11232);
or U11591 (N_11591,N_11433,N_11160);
nor U11592 (N_11592,N_11176,N_11315);
or U11593 (N_11593,N_11133,N_11085);
or U11594 (N_11594,N_11011,N_11191);
and U11595 (N_11595,N_11032,N_11486);
or U11596 (N_11596,N_11041,N_11048);
and U11597 (N_11597,N_11278,N_11208);
or U11598 (N_11598,N_11326,N_11028);
nor U11599 (N_11599,N_11299,N_11238);
nand U11600 (N_11600,N_11397,N_11411);
nand U11601 (N_11601,N_11289,N_11043);
nor U11602 (N_11602,N_11012,N_11369);
or U11603 (N_11603,N_11019,N_11455);
nor U11604 (N_11604,N_11224,N_11141);
xor U11605 (N_11605,N_11219,N_11018);
and U11606 (N_11606,N_11068,N_11015);
nor U11607 (N_11607,N_11282,N_11193);
nand U11608 (N_11608,N_11481,N_11118);
nand U11609 (N_11609,N_11423,N_11263);
nand U11610 (N_11610,N_11145,N_11403);
or U11611 (N_11611,N_11418,N_11162);
xor U11612 (N_11612,N_11448,N_11344);
or U11613 (N_11613,N_11363,N_11008);
nor U11614 (N_11614,N_11259,N_11340);
nor U11615 (N_11615,N_11053,N_11307);
or U11616 (N_11616,N_11103,N_11090);
or U11617 (N_11617,N_11123,N_11243);
or U11618 (N_11618,N_11370,N_11275);
xnor U11619 (N_11619,N_11302,N_11021);
nand U11620 (N_11620,N_11097,N_11190);
nand U11621 (N_11621,N_11491,N_11428);
nand U11622 (N_11622,N_11184,N_11217);
nor U11623 (N_11623,N_11101,N_11318);
nor U11624 (N_11624,N_11116,N_11216);
nand U11625 (N_11625,N_11034,N_11108);
or U11626 (N_11626,N_11242,N_11399);
nor U11627 (N_11627,N_11072,N_11054);
or U11628 (N_11628,N_11007,N_11362);
nand U11629 (N_11629,N_11002,N_11284);
and U11630 (N_11630,N_11013,N_11407);
nand U11631 (N_11631,N_11044,N_11429);
xor U11632 (N_11632,N_11380,N_11328);
or U11633 (N_11633,N_11267,N_11006);
and U11634 (N_11634,N_11197,N_11327);
nor U11635 (N_11635,N_11319,N_11182);
and U11636 (N_11636,N_11256,N_11179);
nor U11637 (N_11637,N_11279,N_11199);
or U11638 (N_11638,N_11058,N_11207);
or U11639 (N_11639,N_11126,N_11111);
nor U11640 (N_11640,N_11406,N_11040);
xnor U11641 (N_11641,N_11404,N_11280);
and U11642 (N_11642,N_11271,N_11436);
or U11643 (N_11643,N_11474,N_11477);
and U11644 (N_11644,N_11321,N_11405);
nor U11645 (N_11645,N_11127,N_11353);
nand U11646 (N_11646,N_11014,N_11331);
or U11647 (N_11647,N_11309,N_11234);
or U11648 (N_11648,N_11237,N_11374);
or U11649 (N_11649,N_11401,N_11061);
nand U11650 (N_11650,N_11213,N_11493);
nand U11651 (N_11651,N_11449,N_11274);
xor U11652 (N_11652,N_11414,N_11200);
xor U11653 (N_11653,N_11075,N_11244);
and U11654 (N_11654,N_11391,N_11443);
or U11655 (N_11655,N_11071,N_11099);
xnor U11656 (N_11656,N_11281,N_11446);
and U11657 (N_11657,N_11392,N_11150);
nor U11658 (N_11658,N_11114,N_11466);
nor U11659 (N_11659,N_11314,N_11352);
xnor U11660 (N_11660,N_11204,N_11087);
nand U11661 (N_11661,N_11255,N_11295);
or U11662 (N_11662,N_11230,N_11283);
xor U11663 (N_11663,N_11033,N_11365);
nor U11664 (N_11664,N_11175,N_11091);
nand U11665 (N_11665,N_11385,N_11024);
or U11666 (N_11666,N_11310,N_11136);
or U11667 (N_11667,N_11360,N_11178);
xnor U11668 (N_11668,N_11201,N_11096);
nand U11669 (N_11669,N_11189,N_11194);
and U11670 (N_11670,N_11268,N_11316);
xnor U11671 (N_11671,N_11394,N_11441);
nor U11672 (N_11672,N_11485,N_11240);
and U11673 (N_11673,N_11210,N_11196);
nor U11674 (N_11674,N_11186,N_11494);
nor U11675 (N_11675,N_11147,N_11017);
or U11676 (N_11676,N_11171,N_11425);
or U11677 (N_11677,N_11206,N_11115);
xnor U11678 (N_11678,N_11462,N_11078);
and U11679 (N_11679,N_11422,N_11131);
xnor U11680 (N_11680,N_11142,N_11346);
and U11681 (N_11681,N_11212,N_11270);
or U11682 (N_11682,N_11451,N_11027);
nor U11683 (N_11683,N_11104,N_11426);
and U11684 (N_11684,N_11490,N_11154);
and U11685 (N_11685,N_11301,N_11153);
nand U11686 (N_11686,N_11389,N_11152);
nor U11687 (N_11687,N_11119,N_11367);
nand U11688 (N_11688,N_11177,N_11218);
nor U11689 (N_11689,N_11431,N_11052);
nor U11690 (N_11690,N_11076,N_11226);
or U11691 (N_11691,N_11135,N_11003);
or U11692 (N_11692,N_11106,N_11060);
nand U11693 (N_11693,N_11181,N_11290);
and U11694 (N_11694,N_11046,N_11432);
nand U11695 (N_11695,N_11459,N_11001);
and U11696 (N_11696,N_11198,N_11195);
nand U11697 (N_11697,N_11170,N_11159);
or U11698 (N_11698,N_11161,N_11092);
and U11699 (N_11699,N_11249,N_11349);
and U11700 (N_11700,N_11336,N_11330);
nand U11701 (N_11701,N_11445,N_11487);
xor U11702 (N_11702,N_11169,N_11129);
xor U11703 (N_11703,N_11410,N_11070);
nand U11704 (N_11704,N_11112,N_11235);
nand U11705 (N_11705,N_11140,N_11472);
xnor U11706 (N_11706,N_11335,N_11134);
nand U11707 (N_11707,N_11203,N_11375);
nand U11708 (N_11708,N_11355,N_11016);
nand U11709 (N_11709,N_11276,N_11442);
nor U11710 (N_11710,N_11188,N_11079);
xnor U11711 (N_11711,N_11183,N_11125);
and U11712 (N_11712,N_11187,N_11055);
nor U11713 (N_11713,N_11137,N_11105);
or U11714 (N_11714,N_11475,N_11408);
or U11715 (N_11715,N_11323,N_11415);
nor U11716 (N_11716,N_11312,N_11022);
nand U11717 (N_11717,N_11143,N_11080);
xnor U11718 (N_11718,N_11174,N_11497);
nor U11719 (N_11719,N_11473,N_11180);
xor U11720 (N_11720,N_11042,N_11317);
nand U11721 (N_11721,N_11265,N_11427);
and U11722 (N_11722,N_11253,N_11298);
nand U11723 (N_11723,N_11248,N_11158);
nor U11724 (N_11724,N_11156,N_11030);
nor U11725 (N_11725,N_11384,N_11361);
or U11726 (N_11726,N_11269,N_11004);
nor U11727 (N_11727,N_11461,N_11341);
and U11728 (N_11728,N_11221,N_11132);
or U11729 (N_11729,N_11209,N_11138);
nand U11730 (N_11730,N_11185,N_11498);
nor U11731 (N_11731,N_11057,N_11463);
xnor U11732 (N_11732,N_11345,N_11416);
nor U11733 (N_11733,N_11396,N_11035);
nor U11734 (N_11734,N_11480,N_11069);
xor U11735 (N_11735,N_11413,N_11233);
xnor U11736 (N_11736,N_11371,N_11102);
or U11737 (N_11737,N_11228,N_11168);
and U11738 (N_11738,N_11258,N_11456);
xnor U11739 (N_11739,N_11383,N_11023);
nand U11740 (N_11740,N_11059,N_11476);
nand U11741 (N_11741,N_11420,N_11222);
or U11742 (N_11742,N_11067,N_11390);
or U11743 (N_11743,N_11489,N_11464);
nor U11744 (N_11744,N_11324,N_11372);
xnor U11745 (N_11745,N_11151,N_11496);
or U11746 (N_11746,N_11120,N_11094);
nand U11747 (N_11747,N_11291,N_11469);
nand U11748 (N_11748,N_11026,N_11225);
xor U11749 (N_11749,N_11065,N_11260);
nor U11750 (N_11750,N_11299,N_11026);
or U11751 (N_11751,N_11258,N_11443);
nor U11752 (N_11752,N_11217,N_11409);
and U11753 (N_11753,N_11128,N_11351);
xor U11754 (N_11754,N_11351,N_11414);
nor U11755 (N_11755,N_11281,N_11092);
nand U11756 (N_11756,N_11495,N_11453);
xnor U11757 (N_11757,N_11061,N_11310);
or U11758 (N_11758,N_11357,N_11263);
nor U11759 (N_11759,N_11162,N_11171);
nand U11760 (N_11760,N_11256,N_11102);
nand U11761 (N_11761,N_11271,N_11379);
and U11762 (N_11762,N_11412,N_11170);
xor U11763 (N_11763,N_11402,N_11413);
nand U11764 (N_11764,N_11001,N_11326);
and U11765 (N_11765,N_11363,N_11115);
nor U11766 (N_11766,N_11404,N_11172);
nand U11767 (N_11767,N_11007,N_11205);
or U11768 (N_11768,N_11107,N_11480);
nand U11769 (N_11769,N_11420,N_11251);
and U11770 (N_11770,N_11042,N_11287);
or U11771 (N_11771,N_11494,N_11016);
nand U11772 (N_11772,N_11263,N_11124);
and U11773 (N_11773,N_11130,N_11074);
or U11774 (N_11774,N_11391,N_11035);
and U11775 (N_11775,N_11409,N_11147);
or U11776 (N_11776,N_11488,N_11063);
or U11777 (N_11777,N_11330,N_11305);
or U11778 (N_11778,N_11332,N_11455);
or U11779 (N_11779,N_11053,N_11055);
nor U11780 (N_11780,N_11400,N_11063);
xor U11781 (N_11781,N_11471,N_11157);
and U11782 (N_11782,N_11494,N_11375);
or U11783 (N_11783,N_11021,N_11004);
nand U11784 (N_11784,N_11281,N_11045);
and U11785 (N_11785,N_11019,N_11498);
nor U11786 (N_11786,N_11017,N_11410);
nor U11787 (N_11787,N_11463,N_11442);
or U11788 (N_11788,N_11213,N_11424);
and U11789 (N_11789,N_11372,N_11245);
xnor U11790 (N_11790,N_11222,N_11378);
xnor U11791 (N_11791,N_11394,N_11067);
and U11792 (N_11792,N_11098,N_11278);
or U11793 (N_11793,N_11195,N_11088);
nor U11794 (N_11794,N_11321,N_11240);
xnor U11795 (N_11795,N_11375,N_11206);
xnor U11796 (N_11796,N_11386,N_11494);
nor U11797 (N_11797,N_11277,N_11385);
nand U11798 (N_11798,N_11170,N_11345);
or U11799 (N_11799,N_11259,N_11010);
nor U11800 (N_11800,N_11207,N_11247);
xor U11801 (N_11801,N_11390,N_11493);
xnor U11802 (N_11802,N_11218,N_11274);
nor U11803 (N_11803,N_11261,N_11035);
and U11804 (N_11804,N_11033,N_11230);
nor U11805 (N_11805,N_11074,N_11058);
nand U11806 (N_11806,N_11219,N_11247);
and U11807 (N_11807,N_11227,N_11239);
nand U11808 (N_11808,N_11198,N_11343);
and U11809 (N_11809,N_11317,N_11392);
or U11810 (N_11810,N_11129,N_11090);
nor U11811 (N_11811,N_11145,N_11428);
nor U11812 (N_11812,N_11492,N_11232);
xnor U11813 (N_11813,N_11201,N_11348);
and U11814 (N_11814,N_11348,N_11238);
or U11815 (N_11815,N_11235,N_11314);
xor U11816 (N_11816,N_11266,N_11488);
xor U11817 (N_11817,N_11170,N_11376);
and U11818 (N_11818,N_11141,N_11460);
or U11819 (N_11819,N_11155,N_11382);
nand U11820 (N_11820,N_11211,N_11496);
xnor U11821 (N_11821,N_11304,N_11332);
or U11822 (N_11822,N_11099,N_11401);
and U11823 (N_11823,N_11391,N_11085);
and U11824 (N_11824,N_11478,N_11446);
nand U11825 (N_11825,N_11251,N_11129);
and U11826 (N_11826,N_11112,N_11120);
or U11827 (N_11827,N_11454,N_11205);
or U11828 (N_11828,N_11364,N_11410);
nor U11829 (N_11829,N_11163,N_11195);
nor U11830 (N_11830,N_11019,N_11386);
xor U11831 (N_11831,N_11022,N_11458);
xnor U11832 (N_11832,N_11429,N_11229);
nand U11833 (N_11833,N_11339,N_11320);
nand U11834 (N_11834,N_11251,N_11066);
nor U11835 (N_11835,N_11176,N_11249);
or U11836 (N_11836,N_11149,N_11227);
xor U11837 (N_11837,N_11165,N_11314);
xnor U11838 (N_11838,N_11242,N_11497);
xnor U11839 (N_11839,N_11245,N_11174);
nor U11840 (N_11840,N_11038,N_11365);
xor U11841 (N_11841,N_11024,N_11495);
nand U11842 (N_11842,N_11115,N_11321);
and U11843 (N_11843,N_11159,N_11422);
and U11844 (N_11844,N_11494,N_11465);
xnor U11845 (N_11845,N_11383,N_11003);
nor U11846 (N_11846,N_11269,N_11181);
and U11847 (N_11847,N_11404,N_11019);
or U11848 (N_11848,N_11473,N_11412);
xnor U11849 (N_11849,N_11482,N_11225);
and U11850 (N_11850,N_11063,N_11439);
and U11851 (N_11851,N_11231,N_11155);
nor U11852 (N_11852,N_11213,N_11021);
nand U11853 (N_11853,N_11190,N_11232);
xnor U11854 (N_11854,N_11215,N_11162);
nand U11855 (N_11855,N_11475,N_11271);
or U11856 (N_11856,N_11351,N_11466);
nand U11857 (N_11857,N_11119,N_11205);
or U11858 (N_11858,N_11282,N_11219);
or U11859 (N_11859,N_11021,N_11465);
nand U11860 (N_11860,N_11378,N_11224);
nand U11861 (N_11861,N_11134,N_11185);
or U11862 (N_11862,N_11419,N_11353);
nor U11863 (N_11863,N_11341,N_11439);
and U11864 (N_11864,N_11289,N_11449);
or U11865 (N_11865,N_11409,N_11375);
and U11866 (N_11866,N_11489,N_11137);
xor U11867 (N_11867,N_11356,N_11057);
or U11868 (N_11868,N_11135,N_11011);
and U11869 (N_11869,N_11479,N_11056);
and U11870 (N_11870,N_11349,N_11307);
or U11871 (N_11871,N_11402,N_11118);
nand U11872 (N_11872,N_11217,N_11222);
nor U11873 (N_11873,N_11373,N_11361);
nor U11874 (N_11874,N_11368,N_11382);
xor U11875 (N_11875,N_11155,N_11419);
xnor U11876 (N_11876,N_11361,N_11341);
nand U11877 (N_11877,N_11053,N_11336);
and U11878 (N_11878,N_11063,N_11210);
nand U11879 (N_11879,N_11324,N_11229);
nor U11880 (N_11880,N_11176,N_11365);
and U11881 (N_11881,N_11331,N_11180);
and U11882 (N_11882,N_11275,N_11407);
and U11883 (N_11883,N_11200,N_11445);
or U11884 (N_11884,N_11060,N_11084);
nand U11885 (N_11885,N_11377,N_11065);
and U11886 (N_11886,N_11488,N_11231);
or U11887 (N_11887,N_11080,N_11114);
and U11888 (N_11888,N_11301,N_11358);
nor U11889 (N_11889,N_11098,N_11077);
nor U11890 (N_11890,N_11141,N_11266);
or U11891 (N_11891,N_11307,N_11100);
nand U11892 (N_11892,N_11244,N_11423);
xor U11893 (N_11893,N_11102,N_11315);
or U11894 (N_11894,N_11420,N_11443);
or U11895 (N_11895,N_11143,N_11208);
and U11896 (N_11896,N_11387,N_11029);
nand U11897 (N_11897,N_11275,N_11394);
nor U11898 (N_11898,N_11403,N_11220);
nor U11899 (N_11899,N_11349,N_11236);
or U11900 (N_11900,N_11110,N_11219);
nor U11901 (N_11901,N_11313,N_11396);
and U11902 (N_11902,N_11145,N_11317);
and U11903 (N_11903,N_11089,N_11336);
nand U11904 (N_11904,N_11495,N_11335);
nand U11905 (N_11905,N_11376,N_11027);
or U11906 (N_11906,N_11099,N_11277);
nor U11907 (N_11907,N_11053,N_11077);
xor U11908 (N_11908,N_11232,N_11252);
nand U11909 (N_11909,N_11152,N_11278);
xor U11910 (N_11910,N_11398,N_11137);
nor U11911 (N_11911,N_11313,N_11453);
xnor U11912 (N_11912,N_11279,N_11114);
xnor U11913 (N_11913,N_11421,N_11233);
or U11914 (N_11914,N_11107,N_11194);
or U11915 (N_11915,N_11310,N_11491);
xnor U11916 (N_11916,N_11104,N_11196);
or U11917 (N_11917,N_11420,N_11254);
or U11918 (N_11918,N_11100,N_11338);
or U11919 (N_11919,N_11085,N_11482);
nand U11920 (N_11920,N_11417,N_11380);
or U11921 (N_11921,N_11093,N_11432);
xnor U11922 (N_11922,N_11055,N_11478);
xor U11923 (N_11923,N_11185,N_11213);
xor U11924 (N_11924,N_11110,N_11473);
nand U11925 (N_11925,N_11206,N_11348);
and U11926 (N_11926,N_11065,N_11399);
nand U11927 (N_11927,N_11445,N_11307);
nor U11928 (N_11928,N_11167,N_11184);
nand U11929 (N_11929,N_11151,N_11022);
xnor U11930 (N_11930,N_11475,N_11319);
or U11931 (N_11931,N_11010,N_11160);
or U11932 (N_11932,N_11145,N_11493);
nor U11933 (N_11933,N_11199,N_11031);
or U11934 (N_11934,N_11200,N_11156);
nor U11935 (N_11935,N_11110,N_11306);
nand U11936 (N_11936,N_11207,N_11392);
nand U11937 (N_11937,N_11273,N_11035);
or U11938 (N_11938,N_11383,N_11020);
nor U11939 (N_11939,N_11017,N_11065);
and U11940 (N_11940,N_11188,N_11254);
nand U11941 (N_11941,N_11116,N_11440);
nor U11942 (N_11942,N_11020,N_11149);
xnor U11943 (N_11943,N_11097,N_11235);
nor U11944 (N_11944,N_11496,N_11478);
nor U11945 (N_11945,N_11120,N_11319);
or U11946 (N_11946,N_11161,N_11467);
xor U11947 (N_11947,N_11273,N_11085);
and U11948 (N_11948,N_11458,N_11445);
nor U11949 (N_11949,N_11229,N_11146);
or U11950 (N_11950,N_11437,N_11005);
nor U11951 (N_11951,N_11179,N_11226);
nor U11952 (N_11952,N_11209,N_11177);
or U11953 (N_11953,N_11189,N_11298);
and U11954 (N_11954,N_11044,N_11437);
nand U11955 (N_11955,N_11068,N_11215);
and U11956 (N_11956,N_11014,N_11222);
nand U11957 (N_11957,N_11234,N_11351);
and U11958 (N_11958,N_11379,N_11272);
and U11959 (N_11959,N_11228,N_11109);
nand U11960 (N_11960,N_11420,N_11246);
xor U11961 (N_11961,N_11016,N_11241);
or U11962 (N_11962,N_11139,N_11007);
or U11963 (N_11963,N_11221,N_11214);
nor U11964 (N_11964,N_11250,N_11349);
xnor U11965 (N_11965,N_11411,N_11202);
nor U11966 (N_11966,N_11463,N_11061);
and U11967 (N_11967,N_11246,N_11181);
or U11968 (N_11968,N_11064,N_11339);
and U11969 (N_11969,N_11314,N_11307);
nor U11970 (N_11970,N_11153,N_11350);
and U11971 (N_11971,N_11463,N_11445);
nor U11972 (N_11972,N_11408,N_11146);
xor U11973 (N_11973,N_11153,N_11337);
xnor U11974 (N_11974,N_11330,N_11006);
or U11975 (N_11975,N_11086,N_11004);
xnor U11976 (N_11976,N_11309,N_11133);
nand U11977 (N_11977,N_11061,N_11379);
nor U11978 (N_11978,N_11464,N_11245);
xor U11979 (N_11979,N_11419,N_11234);
or U11980 (N_11980,N_11431,N_11487);
and U11981 (N_11981,N_11481,N_11102);
or U11982 (N_11982,N_11397,N_11168);
or U11983 (N_11983,N_11114,N_11131);
and U11984 (N_11984,N_11140,N_11443);
xor U11985 (N_11985,N_11412,N_11346);
xor U11986 (N_11986,N_11171,N_11349);
and U11987 (N_11987,N_11476,N_11432);
xnor U11988 (N_11988,N_11483,N_11289);
or U11989 (N_11989,N_11299,N_11063);
or U11990 (N_11990,N_11447,N_11474);
or U11991 (N_11991,N_11080,N_11384);
nor U11992 (N_11992,N_11308,N_11273);
xor U11993 (N_11993,N_11284,N_11045);
nor U11994 (N_11994,N_11296,N_11397);
or U11995 (N_11995,N_11260,N_11061);
and U11996 (N_11996,N_11457,N_11475);
nor U11997 (N_11997,N_11495,N_11038);
nand U11998 (N_11998,N_11005,N_11006);
nand U11999 (N_11999,N_11394,N_11213);
and U12000 (N_12000,N_11525,N_11623);
nor U12001 (N_12001,N_11921,N_11759);
or U12002 (N_12002,N_11627,N_11941);
nor U12003 (N_12003,N_11832,N_11987);
nor U12004 (N_12004,N_11583,N_11581);
and U12005 (N_12005,N_11753,N_11961);
nand U12006 (N_12006,N_11874,N_11988);
and U12007 (N_12007,N_11822,N_11663);
xnor U12008 (N_12008,N_11823,N_11861);
xnor U12009 (N_12009,N_11664,N_11947);
nor U12010 (N_12010,N_11705,N_11710);
xnor U12011 (N_12011,N_11790,N_11892);
xnor U12012 (N_12012,N_11797,N_11637);
xor U12013 (N_12013,N_11902,N_11957);
and U12014 (N_12014,N_11904,N_11628);
xnor U12015 (N_12015,N_11555,N_11643);
nor U12016 (N_12016,N_11945,N_11682);
nor U12017 (N_12017,N_11740,N_11504);
nand U12018 (N_12018,N_11836,N_11994);
xor U12019 (N_12019,N_11922,N_11508);
nor U12020 (N_12020,N_11986,N_11744);
or U12021 (N_12021,N_11652,N_11636);
xor U12022 (N_12022,N_11760,N_11676);
and U12023 (N_12023,N_11795,N_11825);
nand U12024 (N_12024,N_11560,N_11534);
xor U12025 (N_12025,N_11776,N_11696);
nand U12026 (N_12026,N_11919,N_11924);
or U12027 (N_12027,N_11905,N_11640);
xor U12028 (N_12028,N_11983,N_11789);
xor U12029 (N_12029,N_11767,N_11741);
and U12030 (N_12030,N_11669,N_11769);
and U12031 (N_12031,N_11821,N_11838);
xor U12032 (N_12032,N_11526,N_11893);
nand U12033 (N_12033,N_11932,N_11688);
nand U12034 (N_12034,N_11678,N_11545);
and U12035 (N_12035,N_11649,N_11980);
and U12036 (N_12036,N_11704,N_11511);
or U12037 (N_12037,N_11992,N_11933);
and U12038 (N_12038,N_11595,N_11611);
nor U12039 (N_12039,N_11564,N_11641);
or U12040 (N_12040,N_11996,N_11931);
nand U12041 (N_12041,N_11923,N_11817);
or U12042 (N_12042,N_11804,N_11963);
nor U12043 (N_12043,N_11553,N_11660);
nor U12044 (N_12044,N_11732,N_11949);
and U12045 (N_12045,N_11703,N_11803);
and U12046 (N_12046,N_11608,N_11969);
or U12047 (N_12047,N_11507,N_11756);
or U12048 (N_12048,N_11783,N_11645);
and U12049 (N_12049,N_11749,N_11848);
nand U12050 (N_12050,N_11666,N_11517);
and U12051 (N_12051,N_11548,N_11729);
xnor U12052 (N_12052,N_11990,N_11862);
xor U12053 (N_12053,N_11917,N_11764);
and U12054 (N_12054,N_11738,N_11626);
or U12055 (N_12055,N_11527,N_11857);
xnor U12056 (N_12056,N_11673,N_11551);
nand U12057 (N_12057,N_11968,N_11860);
xor U12058 (N_12058,N_11796,N_11839);
nand U12059 (N_12059,N_11856,N_11758);
and U12060 (N_12060,N_11604,N_11998);
and U12061 (N_12061,N_11711,N_11974);
and U12062 (N_12062,N_11521,N_11780);
xor U12063 (N_12063,N_11700,N_11575);
or U12064 (N_12064,N_11573,N_11791);
nor U12065 (N_12065,N_11993,N_11750);
xnor U12066 (N_12066,N_11519,N_11624);
or U12067 (N_12067,N_11792,N_11943);
nand U12068 (N_12068,N_11718,N_11681);
nor U12069 (N_12069,N_11552,N_11616);
or U12070 (N_12070,N_11934,N_11562);
nand U12071 (N_12071,N_11916,N_11887);
xnor U12072 (N_12072,N_11982,N_11953);
nand U12073 (N_12073,N_11675,N_11634);
nor U12074 (N_12074,N_11510,N_11820);
xnor U12075 (N_12075,N_11829,N_11948);
nor U12076 (N_12076,N_11686,N_11582);
or U12077 (N_12077,N_11854,N_11524);
and U12078 (N_12078,N_11617,N_11544);
or U12079 (N_12079,N_11630,N_11668);
and U12080 (N_12080,N_11814,N_11699);
and U12081 (N_12081,N_11882,N_11930);
nor U12082 (N_12082,N_11737,N_11746);
or U12083 (N_12083,N_11754,N_11539);
xor U12084 (N_12084,N_11942,N_11972);
nor U12085 (N_12085,N_11659,N_11654);
or U12086 (N_12086,N_11818,N_11695);
and U12087 (N_12087,N_11529,N_11501);
xor U12088 (N_12088,N_11572,N_11877);
nand U12089 (N_12089,N_11844,N_11601);
nor U12090 (N_12090,N_11903,N_11502);
and U12091 (N_12091,N_11913,N_11777);
nand U12092 (N_12092,N_11771,N_11964);
and U12093 (N_12093,N_11698,N_11665);
xor U12094 (N_12094,N_11554,N_11894);
and U12095 (N_12095,N_11834,N_11952);
or U12096 (N_12096,N_11542,N_11806);
xnor U12097 (N_12097,N_11745,N_11647);
or U12098 (N_12098,N_11914,N_11667);
or U12099 (N_12099,N_11788,N_11724);
nor U12100 (N_12100,N_11607,N_11944);
nand U12101 (N_12101,N_11879,N_11578);
or U12102 (N_12102,N_11633,N_11546);
nand U12103 (N_12103,N_11708,N_11782);
or U12104 (N_12104,N_11853,N_11869);
nor U12105 (N_12105,N_11895,N_11811);
nor U12106 (N_12106,N_11584,N_11586);
xor U12107 (N_12107,N_11837,N_11748);
xnor U12108 (N_12108,N_11812,N_11719);
xnor U12109 (N_12109,N_11658,N_11801);
and U12110 (N_12110,N_11929,N_11717);
and U12111 (N_12111,N_11543,N_11743);
nor U12112 (N_12112,N_11536,N_11559);
xnor U12113 (N_12113,N_11549,N_11541);
xor U12114 (N_12114,N_11956,N_11997);
xor U12115 (N_12115,N_11752,N_11683);
or U12116 (N_12116,N_11864,N_11785);
nand U12117 (N_12117,N_11565,N_11594);
nand U12118 (N_12118,N_11707,N_11891);
or U12119 (N_12119,N_11661,N_11981);
nor U12120 (N_12120,N_11774,N_11670);
and U12121 (N_12121,N_11935,N_11602);
or U12122 (N_12122,N_11522,N_11888);
or U12123 (N_12123,N_11833,N_11622);
and U12124 (N_12124,N_11687,N_11915);
xnor U12125 (N_12125,N_11690,N_11845);
and U12126 (N_12126,N_11850,N_11723);
and U12127 (N_12127,N_11512,N_11819);
and U12128 (N_12128,N_11937,N_11755);
nand U12129 (N_12129,N_11731,N_11651);
nor U12130 (N_12130,N_11639,N_11898);
and U12131 (N_12131,N_11514,N_11881);
xnor U12132 (N_12132,N_11835,N_11936);
nor U12133 (N_12133,N_11528,N_11609);
nor U12134 (N_12134,N_11655,N_11734);
xor U12135 (N_12135,N_11966,N_11535);
nor U12136 (N_12136,N_11589,N_11950);
xor U12137 (N_12137,N_11677,N_11600);
or U12138 (N_12138,N_11580,N_11959);
nor U12139 (N_12139,N_11779,N_11896);
nor U12140 (N_12140,N_11831,N_11702);
xor U12141 (N_12141,N_11566,N_11558);
nor U12142 (N_12142,N_11939,N_11886);
xor U12143 (N_12143,N_11679,N_11646);
nor U12144 (N_12144,N_11798,N_11672);
nand U12145 (N_12145,N_11979,N_11907);
xnor U12146 (N_12146,N_11612,N_11577);
and U12147 (N_12147,N_11830,N_11733);
and U12148 (N_12148,N_11787,N_11847);
nor U12149 (N_12149,N_11500,N_11516);
nor U12150 (N_12150,N_11912,N_11975);
nor U12151 (N_12151,N_11840,N_11619);
nand U12152 (N_12152,N_11576,N_11799);
or U12153 (N_12153,N_11662,N_11701);
nand U12154 (N_12154,N_11786,N_11644);
nor U12155 (N_12155,N_11985,N_11725);
nand U12156 (N_12156,N_11841,N_11505);
or U12157 (N_12157,N_11598,N_11807);
nor U12158 (N_12158,N_11557,N_11653);
nand U12159 (N_12159,N_11618,N_11973);
or U12160 (N_12160,N_11824,N_11984);
nor U12161 (N_12161,N_11770,N_11709);
nor U12162 (N_12162,N_11778,N_11694);
nor U12163 (N_12163,N_11757,N_11563);
nor U12164 (N_12164,N_11603,N_11899);
or U12165 (N_12165,N_11631,N_11650);
or U12166 (N_12166,N_11716,N_11715);
and U12167 (N_12167,N_11712,N_11951);
and U12168 (N_12168,N_11561,N_11920);
xor U12169 (N_12169,N_11808,N_11591);
nor U12170 (N_12170,N_11625,N_11851);
and U12171 (N_12171,N_11550,N_11926);
and U12172 (N_12172,N_11518,N_11908);
nand U12173 (N_12173,N_11685,N_11585);
or U12174 (N_12174,N_11978,N_11592);
and U12175 (N_12175,N_11865,N_11859);
xnor U12176 (N_12176,N_11995,N_11910);
nor U12177 (N_12177,N_11761,N_11773);
or U12178 (N_12178,N_11889,N_11946);
nand U12179 (N_12179,N_11960,N_11843);
nand U12180 (N_12180,N_11503,N_11523);
or U12181 (N_12181,N_11691,N_11714);
xor U12182 (N_12182,N_11515,N_11849);
nand U12183 (N_12183,N_11620,N_11689);
nor U12184 (N_12184,N_11697,N_11727);
nand U12185 (N_12185,N_11588,N_11858);
and U12186 (N_12186,N_11537,N_11736);
or U12187 (N_12187,N_11901,N_11763);
and U12188 (N_12188,N_11794,N_11962);
or U12189 (N_12189,N_11574,N_11976);
nand U12190 (N_12190,N_11613,N_11684);
or U12191 (N_12191,N_11873,N_11579);
or U12192 (N_12192,N_11958,N_11506);
or U12193 (N_12193,N_11742,N_11762);
or U12194 (N_12194,N_11547,N_11875);
xnor U12195 (N_12195,N_11828,N_11827);
nor U12196 (N_12196,N_11629,N_11846);
nor U12197 (N_12197,N_11642,N_11615);
nand U12198 (N_12198,N_11775,N_11826);
nand U12199 (N_12199,N_11885,N_11813);
and U12200 (N_12200,N_11610,N_11938);
xor U12201 (N_12201,N_11872,N_11621);
and U12202 (N_12202,N_11569,N_11810);
and U12203 (N_12203,N_11970,N_11567);
nor U12204 (N_12204,N_11906,N_11900);
nand U12205 (N_12205,N_11590,N_11772);
xnor U12206 (N_12206,N_11635,N_11940);
and U12207 (N_12207,N_11765,N_11965);
or U12208 (N_12208,N_11781,N_11855);
and U12209 (N_12209,N_11870,N_11878);
nor U12210 (N_12210,N_11532,N_11513);
nand U12211 (N_12211,N_11568,N_11954);
or U12212 (N_12212,N_11648,N_11871);
and U12213 (N_12213,N_11955,N_11722);
nor U12214 (N_12214,N_11928,N_11706);
xor U12215 (N_12215,N_11531,N_11656);
nor U12216 (N_12216,N_11863,N_11897);
xor U12217 (N_12217,N_11614,N_11766);
nor U12218 (N_12218,N_11883,N_11868);
or U12219 (N_12219,N_11571,N_11720);
and U12220 (N_12220,N_11728,N_11596);
or U12221 (N_12221,N_11991,N_11768);
or U12222 (N_12222,N_11927,N_11713);
and U12223 (N_12223,N_11802,N_11784);
nor U12224 (N_12224,N_11805,N_11632);
nand U12225 (N_12225,N_11852,N_11816);
nor U12226 (N_12226,N_11721,N_11540);
nand U12227 (N_12227,N_11739,N_11793);
and U12228 (N_12228,N_11884,N_11693);
and U12229 (N_12229,N_11842,N_11867);
nand U12230 (N_12230,N_11587,N_11726);
nand U12231 (N_12231,N_11866,N_11530);
nor U12232 (N_12232,N_11815,N_11909);
nor U12233 (N_12233,N_11538,N_11533);
nand U12234 (N_12234,N_11657,N_11735);
nor U12235 (N_12235,N_11606,N_11971);
nand U12236 (N_12236,N_11509,N_11751);
and U12237 (N_12237,N_11890,N_11918);
xor U12238 (N_12238,N_11730,N_11977);
nand U12239 (N_12239,N_11638,N_11880);
nor U12240 (N_12240,N_11967,N_11911);
nor U12241 (N_12241,N_11747,N_11599);
nor U12242 (N_12242,N_11520,N_11692);
and U12243 (N_12243,N_11925,N_11809);
nand U12244 (N_12244,N_11556,N_11671);
or U12245 (N_12245,N_11680,N_11605);
and U12246 (N_12246,N_11570,N_11593);
nand U12247 (N_12247,N_11999,N_11800);
and U12248 (N_12248,N_11989,N_11674);
xor U12249 (N_12249,N_11876,N_11597);
nand U12250 (N_12250,N_11779,N_11869);
xor U12251 (N_12251,N_11863,N_11906);
nand U12252 (N_12252,N_11792,N_11576);
xnor U12253 (N_12253,N_11725,N_11761);
or U12254 (N_12254,N_11995,N_11622);
xnor U12255 (N_12255,N_11739,N_11617);
and U12256 (N_12256,N_11879,N_11621);
nor U12257 (N_12257,N_11922,N_11867);
or U12258 (N_12258,N_11515,N_11926);
and U12259 (N_12259,N_11578,N_11501);
xor U12260 (N_12260,N_11934,N_11950);
xnor U12261 (N_12261,N_11955,N_11909);
nand U12262 (N_12262,N_11592,N_11908);
nand U12263 (N_12263,N_11595,N_11967);
and U12264 (N_12264,N_11945,N_11697);
xnor U12265 (N_12265,N_11859,N_11660);
nor U12266 (N_12266,N_11511,N_11726);
nand U12267 (N_12267,N_11811,N_11816);
and U12268 (N_12268,N_11968,N_11510);
or U12269 (N_12269,N_11578,N_11938);
or U12270 (N_12270,N_11708,N_11883);
nand U12271 (N_12271,N_11755,N_11866);
and U12272 (N_12272,N_11710,N_11868);
or U12273 (N_12273,N_11820,N_11548);
nor U12274 (N_12274,N_11808,N_11506);
xor U12275 (N_12275,N_11656,N_11505);
xor U12276 (N_12276,N_11542,N_11698);
nand U12277 (N_12277,N_11551,N_11994);
nor U12278 (N_12278,N_11516,N_11935);
or U12279 (N_12279,N_11983,N_11543);
or U12280 (N_12280,N_11913,N_11655);
or U12281 (N_12281,N_11887,N_11636);
nor U12282 (N_12282,N_11937,N_11872);
nor U12283 (N_12283,N_11969,N_11687);
xnor U12284 (N_12284,N_11967,N_11715);
nand U12285 (N_12285,N_11663,N_11977);
nor U12286 (N_12286,N_11910,N_11720);
and U12287 (N_12287,N_11680,N_11678);
nor U12288 (N_12288,N_11755,N_11644);
and U12289 (N_12289,N_11801,N_11804);
and U12290 (N_12290,N_11594,N_11852);
nor U12291 (N_12291,N_11645,N_11757);
xor U12292 (N_12292,N_11648,N_11873);
nand U12293 (N_12293,N_11559,N_11577);
and U12294 (N_12294,N_11598,N_11700);
nand U12295 (N_12295,N_11997,N_11613);
or U12296 (N_12296,N_11852,N_11796);
and U12297 (N_12297,N_11503,N_11668);
xor U12298 (N_12298,N_11571,N_11797);
nor U12299 (N_12299,N_11808,N_11880);
and U12300 (N_12300,N_11822,N_11877);
xnor U12301 (N_12301,N_11756,N_11621);
nor U12302 (N_12302,N_11592,N_11718);
nor U12303 (N_12303,N_11688,N_11844);
and U12304 (N_12304,N_11525,N_11744);
nor U12305 (N_12305,N_11650,N_11562);
or U12306 (N_12306,N_11945,N_11667);
xor U12307 (N_12307,N_11848,N_11551);
nand U12308 (N_12308,N_11817,N_11588);
and U12309 (N_12309,N_11739,N_11528);
and U12310 (N_12310,N_11652,N_11545);
and U12311 (N_12311,N_11620,N_11912);
nor U12312 (N_12312,N_11822,N_11552);
nor U12313 (N_12313,N_11642,N_11673);
and U12314 (N_12314,N_11754,N_11556);
and U12315 (N_12315,N_11630,N_11740);
and U12316 (N_12316,N_11558,N_11830);
or U12317 (N_12317,N_11795,N_11995);
or U12318 (N_12318,N_11937,N_11999);
xnor U12319 (N_12319,N_11795,N_11758);
and U12320 (N_12320,N_11828,N_11728);
or U12321 (N_12321,N_11893,N_11569);
or U12322 (N_12322,N_11912,N_11714);
or U12323 (N_12323,N_11718,N_11941);
xor U12324 (N_12324,N_11571,N_11653);
or U12325 (N_12325,N_11540,N_11753);
xnor U12326 (N_12326,N_11896,N_11838);
or U12327 (N_12327,N_11873,N_11666);
or U12328 (N_12328,N_11899,N_11525);
and U12329 (N_12329,N_11882,N_11872);
xor U12330 (N_12330,N_11882,N_11805);
nand U12331 (N_12331,N_11763,N_11898);
xnor U12332 (N_12332,N_11759,N_11875);
nand U12333 (N_12333,N_11822,N_11668);
and U12334 (N_12334,N_11970,N_11997);
nor U12335 (N_12335,N_11828,N_11816);
and U12336 (N_12336,N_11517,N_11639);
nand U12337 (N_12337,N_11964,N_11803);
nor U12338 (N_12338,N_11600,N_11771);
xnor U12339 (N_12339,N_11620,N_11692);
or U12340 (N_12340,N_11592,N_11633);
and U12341 (N_12341,N_11824,N_11656);
and U12342 (N_12342,N_11642,N_11827);
or U12343 (N_12343,N_11857,N_11804);
xor U12344 (N_12344,N_11888,N_11503);
xnor U12345 (N_12345,N_11869,N_11700);
nand U12346 (N_12346,N_11777,N_11500);
xnor U12347 (N_12347,N_11551,N_11679);
nand U12348 (N_12348,N_11890,N_11559);
nor U12349 (N_12349,N_11911,N_11910);
nand U12350 (N_12350,N_11665,N_11547);
xor U12351 (N_12351,N_11949,N_11984);
nor U12352 (N_12352,N_11653,N_11728);
nor U12353 (N_12353,N_11649,N_11867);
nand U12354 (N_12354,N_11893,N_11612);
nand U12355 (N_12355,N_11982,N_11568);
nor U12356 (N_12356,N_11668,N_11937);
or U12357 (N_12357,N_11640,N_11699);
and U12358 (N_12358,N_11717,N_11526);
or U12359 (N_12359,N_11708,N_11646);
nand U12360 (N_12360,N_11926,N_11501);
or U12361 (N_12361,N_11637,N_11506);
xnor U12362 (N_12362,N_11893,N_11609);
xnor U12363 (N_12363,N_11929,N_11550);
nand U12364 (N_12364,N_11785,N_11867);
and U12365 (N_12365,N_11839,N_11681);
nand U12366 (N_12366,N_11681,N_11917);
nand U12367 (N_12367,N_11616,N_11925);
xnor U12368 (N_12368,N_11738,N_11775);
or U12369 (N_12369,N_11603,N_11807);
nand U12370 (N_12370,N_11677,N_11751);
and U12371 (N_12371,N_11930,N_11562);
and U12372 (N_12372,N_11659,N_11953);
and U12373 (N_12373,N_11897,N_11692);
or U12374 (N_12374,N_11775,N_11568);
nand U12375 (N_12375,N_11707,N_11590);
nor U12376 (N_12376,N_11950,N_11789);
or U12377 (N_12377,N_11603,N_11588);
nand U12378 (N_12378,N_11814,N_11856);
xor U12379 (N_12379,N_11912,N_11867);
xor U12380 (N_12380,N_11538,N_11680);
nand U12381 (N_12381,N_11980,N_11503);
nand U12382 (N_12382,N_11799,N_11515);
nand U12383 (N_12383,N_11583,N_11995);
xnor U12384 (N_12384,N_11629,N_11702);
nand U12385 (N_12385,N_11866,N_11884);
nor U12386 (N_12386,N_11912,N_11594);
nand U12387 (N_12387,N_11684,N_11995);
and U12388 (N_12388,N_11536,N_11504);
nor U12389 (N_12389,N_11775,N_11786);
xor U12390 (N_12390,N_11760,N_11512);
and U12391 (N_12391,N_11934,N_11970);
and U12392 (N_12392,N_11616,N_11501);
or U12393 (N_12393,N_11926,N_11812);
nor U12394 (N_12394,N_11846,N_11662);
xnor U12395 (N_12395,N_11832,N_11792);
nor U12396 (N_12396,N_11797,N_11550);
nand U12397 (N_12397,N_11939,N_11949);
nand U12398 (N_12398,N_11921,N_11502);
nand U12399 (N_12399,N_11623,N_11861);
nand U12400 (N_12400,N_11917,N_11609);
and U12401 (N_12401,N_11813,N_11530);
nor U12402 (N_12402,N_11821,N_11724);
xnor U12403 (N_12403,N_11641,N_11980);
and U12404 (N_12404,N_11618,N_11805);
xnor U12405 (N_12405,N_11616,N_11674);
xnor U12406 (N_12406,N_11900,N_11695);
nor U12407 (N_12407,N_11828,N_11991);
or U12408 (N_12408,N_11575,N_11892);
or U12409 (N_12409,N_11612,N_11969);
xnor U12410 (N_12410,N_11813,N_11789);
or U12411 (N_12411,N_11833,N_11782);
xnor U12412 (N_12412,N_11910,N_11565);
xnor U12413 (N_12413,N_11786,N_11537);
nor U12414 (N_12414,N_11906,N_11588);
nand U12415 (N_12415,N_11504,N_11754);
xor U12416 (N_12416,N_11747,N_11501);
nand U12417 (N_12417,N_11761,N_11776);
nand U12418 (N_12418,N_11842,N_11598);
and U12419 (N_12419,N_11799,N_11817);
nor U12420 (N_12420,N_11628,N_11992);
nand U12421 (N_12421,N_11524,N_11580);
or U12422 (N_12422,N_11675,N_11700);
or U12423 (N_12423,N_11957,N_11874);
xnor U12424 (N_12424,N_11862,N_11650);
or U12425 (N_12425,N_11756,N_11566);
nand U12426 (N_12426,N_11923,N_11767);
nand U12427 (N_12427,N_11949,N_11510);
nor U12428 (N_12428,N_11834,N_11971);
xor U12429 (N_12429,N_11941,N_11659);
and U12430 (N_12430,N_11575,N_11741);
xor U12431 (N_12431,N_11853,N_11785);
nand U12432 (N_12432,N_11535,N_11656);
and U12433 (N_12433,N_11847,N_11533);
xnor U12434 (N_12434,N_11566,N_11696);
nand U12435 (N_12435,N_11784,N_11881);
xnor U12436 (N_12436,N_11611,N_11897);
xnor U12437 (N_12437,N_11873,N_11989);
xnor U12438 (N_12438,N_11929,N_11620);
nor U12439 (N_12439,N_11659,N_11515);
and U12440 (N_12440,N_11605,N_11681);
xor U12441 (N_12441,N_11930,N_11809);
nand U12442 (N_12442,N_11838,N_11906);
nor U12443 (N_12443,N_11918,N_11590);
or U12444 (N_12444,N_11767,N_11622);
xor U12445 (N_12445,N_11530,N_11882);
nand U12446 (N_12446,N_11775,N_11667);
or U12447 (N_12447,N_11585,N_11704);
xnor U12448 (N_12448,N_11796,N_11851);
or U12449 (N_12449,N_11816,N_11652);
or U12450 (N_12450,N_11723,N_11757);
xor U12451 (N_12451,N_11809,N_11711);
xnor U12452 (N_12452,N_11655,N_11888);
nand U12453 (N_12453,N_11595,N_11691);
and U12454 (N_12454,N_11967,N_11601);
xnor U12455 (N_12455,N_11771,N_11684);
or U12456 (N_12456,N_11868,N_11717);
nor U12457 (N_12457,N_11854,N_11652);
nand U12458 (N_12458,N_11563,N_11952);
xor U12459 (N_12459,N_11740,N_11514);
xnor U12460 (N_12460,N_11544,N_11855);
and U12461 (N_12461,N_11581,N_11909);
nand U12462 (N_12462,N_11820,N_11782);
and U12463 (N_12463,N_11774,N_11582);
nand U12464 (N_12464,N_11829,N_11834);
nor U12465 (N_12465,N_11714,N_11989);
nand U12466 (N_12466,N_11538,N_11968);
or U12467 (N_12467,N_11888,N_11815);
xor U12468 (N_12468,N_11659,N_11916);
xor U12469 (N_12469,N_11600,N_11905);
xnor U12470 (N_12470,N_11732,N_11582);
or U12471 (N_12471,N_11974,N_11916);
nor U12472 (N_12472,N_11728,N_11523);
xor U12473 (N_12473,N_11835,N_11891);
and U12474 (N_12474,N_11575,N_11718);
nand U12475 (N_12475,N_11687,N_11841);
nor U12476 (N_12476,N_11794,N_11526);
and U12477 (N_12477,N_11908,N_11846);
nand U12478 (N_12478,N_11514,N_11998);
xnor U12479 (N_12479,N_11946,N_11911);
nand U12480 (N_12480,N_11789,N_11745);
or U12481 (N_12481,N_11801,N_11614);
nor U12482 (N_12482,N_11831,N_11601);
xor U12483 (N_12483,N_11570,N_11503);
or U12484 (N_12484,N_11799,N_11650);
nor U12485 (N_12485,N_11659,N_11656);
xnor U12486 (N_12486,N_11674,N_11857);
xor U12487 (N_12487,N_11515,N_11924);
nand U12488 (N_12488,N_11590,N_11989);
and U12489 (N_12489,N_11548,N_11698);
or U12490 (N_12490,N_11506,N_11798);
nand U12491 (N_12491,N_11714,N_11661);
nor U12492 (N_12492,N_11933,N_11510);
and U12493 (N_12493,N_11570,N_11934);
nor U12494 (N_12494,N_11877,N_11925);
and U12495 (N_12495,N_11507,N_11985);
nand U12496 (N_12496,N_11579,N_11829);
and U12497 (N_12497,N_11517,N_11759);
and U12498 (N_12498,N_11686,N_11999);
or U12499 (N_12499,N_11919,N_11821);
nand U12500 (N_12500,N_12482,N_12098);
nor U12501 (N_12501,N_12245,N_12380);
or U12502 (N_12502,N_12333,N_12296);
nor U12503 (N_12503,N_12112,N_12331);
xnor U12504 (N_12504,N_12437,N_12060);
nand U12505 (N_12505,N_12092,N_12302);
or U12506 (N_12506,N_12198,N_12035);
nor U12507 (N_12507,N_12462,N_12423);
and U12508 (N_12508,N_12323,N_12254);
or U12509 (N_12509,N_12388,N_12352);
xor U12510 (N_12510,N_12413,N_12474);
or U12511 (N_12511,N_12163,N_12208);
nor U12512 (N_12512,N_12225,N_12085);
nor U12513 (N_12513,N_12068,N_12218);
and U12514 (N_12514,N_12025,N_12237);
and U12515 (N_12515,N_12401,N_12305);
xnor U12516 (N_12516,N_12315,N_12096);
xnor U12517 (N_12517,N_12180,N_12479);
xnor U12518 (N_12518,N_12226,N_12316);
and U12519 (N_12519,N_12212,N_12359);
nor U12520 (N_12520,N_12459,N_12422);
nand U12521 (N_12521,N_12233,N_12165);
or U12522 (N_12522,N_12277,N_12174);
nor U12523 (N_12523,N_12017,N_12371);
xnor U12524 (N_12524,N_12297,N_12032);
xor U12525 (N_12525,N_12478,N_12037);
nor U12526 (N_12526,N_12349,N_12370);
xnor U12527 (N_12527,N_12234,N_12005);
and U12528 (N_12528,N_12116,N_12267);
nor U12529 (N_12529,N_12393,N_12362);
nor U12530 (N_12530,N_12410,N_12337);
xnor U12531 (N_12531,N_12336,N_12468);
or U12532 (N_12532,N_12131,N_12034);
nand U12533 (N_12533,N_12220,N_12383);
nor U12534 (N_12534,N_12409,N_12041);
or U12535 (N_12535,N_12433,N_12055);
xnor U12536 (N_12536,N_12377,N_12382);
and U12537 (N_12537,N_12157,N_12073);
and U12538 (N_12538,N_12070,N_12178);
nand U12539 (N_12539,N_12133,N_12214);
nor U12540 (N_12540,N_12136,N_12464);
nor U12541 (N_12541,N_12213,N_12488);
xor U12542 (N_12542,N_12258,N_12324);
nand U12543 (N_12543,N_12256,N_12222);
xnor U12544 (N_12544,N_12476,N_12083);
and U12545 (N_12545,N_12255,N_12366);
xnor U12546 (N_12546,N_12093,N_12354);
or U12547 (N_12547,N_12113,N_12140);
xor U12548 (N_12548,N_12363,N_12181);
or U12549 (N_12549,N_12499,N_12015);
xnor U12550 (N_12550,N_12168,N_12127);
xnor U12551 (N_12551,N_12334,N_12061);
and U12552 (N_12552,N_12429,N_12403);
and U12553 (N_12553,N_12182,N_12384);
or U12554 (N_12554,N_12425,N_12434);
nor U12555 (N_12555,N_12062,N_12347);
xnor U12556 (N_12556,N_12110,N_12101);
nand U12557 (N_12557,N_12338,N_12114);
nand U12558 (N_12558,N_12151,N_12227);
or U12559 (N_12559,N_12079,N_12161);
nor U12560 (N_12560,N_12210,N_12170);
or U12561 (N_12561,N_12109,N_12192);
nand U12562 (N_12562,N_12230,N_12266);
and U12563 (N_12563,N_12014,N_12106);
and U12564 (N_12564,N_12458,N_12269);
xor U12565 (N_12565,N_12072,N_12265);
or U12566 (N_12566,N_12313,N_12418);
nand U12567 (N_12567,N_12219,N_12463);
or U12568 (N_12568,N_12295,N_12155);
and U12569 (N_12569,N_12412,N_12118);
nor U12570 (N_12570,N_12450,N_12417);
and U12571 (N_12571,N_12376,N_12320);
and U12572 (N_12572,N_12259,N_12054);
xor U12573 (N_12573,N_12030,N_12466);
xnor U12574 (N_12574,N_12360,N_12206);
nand U12575 (N_12575,N_12195,N_12411);
nor U12576 (N_12576,N_12232,N_12453);
and U12577 (N_12577,N_12190,N_12470);
xor U12578 (N_12578,N_12298,N_12355);
or U12579 (N_12579,N_12443,N_12238);
and U12580 (N_12580,N_12247,N_12314);
xor U12581 (N_12581,N_12461,N_12497);
nor U12582 (N_12582,N_12430,N_12457);
nor U12583 (N_12583,N_12188,N_12357);
and U12584 (N_12584,N_12090,N_12335);
nor U12585 (N_12585,N_12375,N_12204);
and U12586 (N_12586,N_12289,N_12150);
nor U12587 (N_12587,N_12033,N_12166);
and U12588 (N_12588,N_12406,N_12175);
nor U12589 (N_12589,N_12487,N_12089);
xor U12590 (N_12590,N_12307,N_12299);
or U12591 (N_12591,N_12031,N_12004);
nand U12592 (N_12592,N_12398,N_12148);
or U12593 (N_12593,N_12130,N_12164);
xor U12594 (N_12594,N_12444,N_12187);
nor U12595 (N_12595,N_12330,N_12452);
xnor U12596 (N_12596,N_12471,N_12121);
nand U12597 (N_12597,N_12396,N_12077);
nand U12598 (N_12598,N_12132,N_12167);
nand U12599 (N_12599,N_12228,N_12491);
nor U12600 (N_12600,N_12285,N_12350);
nand U12601 (N_12601,N_12293,N_12253);
nand U12602 (N_12602,N_12008,N_12067);
or U12603 (N_12603,N_12088,N_12124);
and U12604 (N_12604,N_12351,N_12138);
nand U12605 (N_12605,N_12078,N_12494);
nand U12606 (N_12606,N_12395,N_12045);
nor U12607 (N_12607,N_12217,N_12100);
or U12608 (N_12608,N_12128,N_12416);
or U12609 (N_12609,N_12224,N_12102);
nor U12610 (N_12610,N_12492,N_12344);
or U12611 (N_12611,N_12194,N_12428);
xor U12612 (N_12612,N_12493,N_12365);
nor U12613 (N_12613,N_12318,N_12086);
nand U12614 (N_12614,N_12473,N_12144);
xnor U12615 (N_12615,N_12003,N_12049);
nor U12616 (N_12616,N_12381,N_12402);
nor U12617 (N_12617,N_12278,N_12036);
and U12618 (N_12618,N_12020,N_12039);
nor U12619 (N_12619,N_12016,N_12009);
nand U12620 (N_12620,N_12094,N_12252);
xnor U12621 (N_12621,N_12431,N_12294);
or U12622 (N_12622,N_12435,N_12104);
nor U12623 (N_12623,N_12475,N_12052);
and U12624 (N_12624,N_12340,N_12415);
nor U12625 (N_12625,N_12235,N_12319);
or U12626 (N_12626,N_12056,N_12309);
nor U12627 (N_12627,N_12262,N_12229);
and U12628 (N_12628,N_12490,N_12201);
nand U12629 (N_12629,N_12451,N_12279);
and U12630 (N_12630,N_12483,N_12361);
and U12631 (N_12631,N_12244,N_12274);
xnor U12632 (N_12632,N_12146,N_12481);
nor U12633 (N_12633,N_12426,N_12169);
nor U12634 (N_12634,N_12438,N_12047);
nand U12635 (N_12635,N_12291,N_12058);
or U12636 (N_12636,N_12485,N_12257);
and U12637 (N_12637,N_12249,N_12159);
or U12638 (N_12638,N_12071,N_12177);
and U12639 (N_12639,N_12300,N_12427);
and U12640 (N_12640,N_12420,N_12044);
and U12641 (N_12641,N_12465,N_12456);
nand U12642 (N_12642,N_12322,N_12143);
or U12643 (N_12643,N_12405,N_12023);
and U12644 (N_12644,N_12075,N_12341);
nand U12645 (N_12645,N_12028,N_12115);
nor U12646 (N_12646,N_12126,N_12263);
and U12647 (N_12647,N_12001,N_12160);
and U12648 (N_12648,N_12173,N_12308);
or U12649 (N_12649,N_12097,N_12455);
nor U12650 (N_12650,N_12348,N_12260);
or U12651 (N_12651,N_12236,N_12189);
nor U12652 (N_12652,N_12123,N_12385);
nor U12653 (N_12653,N_12408,N_12183);
xor U12654 (N_12654,N_12185,N_12449);
xnor U12655 (N_12655,N_12460,N_12446);
and U12656 (N_12656,N_12137,N_12122);
nor U12657 (N_12657,N_12184,N_12242);
or U12658 (N_12658,N_12241,N_12368);
nor U12659 (N_12659,N_12000,N_12276);
nor U12660 (N_12660,N_12286,N_12303);
xnor U12661 (N_12661,N_12059,N_12372);
or U12662 (N_12662,N_12440,N_12271);
nor U12663 (N_12663,N_12284,N_12087);
nand U12664 (N_12664,N_12280,N_12149);
xor U12665 (N_12665,N_12231,N_12043);
and U12666 (N_12666,N_12442,N_12125);
or U12667 (N_12667,N_12147,N_12369);
nor U12668 (N_12668,N_12171,N_12304);
xnor U12669 (N_12669,N_12342,N_12251);
nor U12670 (N_12670,N_12356,N_12447);
nor U12671 (N_12671,N_12081,N_12107);
xnor U12672 (N_12672,N_12239,N_12095);
nand U12673 (N_12673,N_12216,N_12467);
and U12674 (N_12674,N_12379,N_12432);
xnor U12675 (N_12675,N_12392,N_12221);
and U12676 (N_12676,N_12424,N_12076);
xnor U12677 (N_12677,N_12290,N_12211);
xnor U12678 (N_12678,N_12011,N_12480);
or U12679 (N_12679,N_12172,N_12080);
and U12680 (N_12680,N_12270,N_12367);
and U12681 (N_12681,N_12454,N_12013);
nand U12682 (N_12682,N_12153,N_12378);
or U12683 (N_12683,N_12158,N_12019);
nand U12684 (N_12684,N_12272,N_12358);
nand U12685 (N_12685,N_12496,N_12301);
nand U12686 (N_12686,N_12108,N_12002);
nor U12687 (N_12687,N_12012,N_12103);
nand U12688 (N_12688,N_12292,N_12248);
nor U12689 (N_12689,N_12250,N_12105);
xnor U12690 (N_12690,N_12495,N_12007);
nor U12691 (N_12691,N_12200,N_12082);
and U12692 (N_12692,N_12288,N_12091);
nor U12693 (N_12693,N_12389,N_12472);
and U12694 (N_12694,N_12387,N_12026);
xor U12695 (N_12695,N_12154,N_12339);
or U12696 (N_12696,N_12006,N_12040);
or U12697 (N_12697,N_12145,N_12264);
nand U12698 (N_12698,N_12141,N_12329);
nand U12699 (N_12699,N_12135,N_12018);
nand U12700 (N_12700,N_12186,N_12207);
nand U12701 (N_12701,N_12317,N_12332);
xor U12702 (N_12702,N_12312,N_12048);
nor U12703 (N_12703,N_12205,N_12042);
nand U12704 (N_12704,N_12281,N_12024);
or U12705 (N_12705,N_12129,N_12246);
nor U12706 (N_12706,N_12283,N_12223);
xnor U12707 (N_12707,N_12268,N_12046);
or U12708 (N_12708,N_12117,N_12179);
and U12709 (N_12709,N_12484,N_12394);
xor U12710 (N_12710,N_12074,N_12240);
nand U12711 (N_12711,N_12199,N_12399);
or U12712 (N_12712,N_12439,N_12197);
and U12713 (N_12713,N_12469,N_12152);
or U12714 (N_12714,N_12287,N_12386);
nor U12715 (N_12715,N_12193,N_12343);
xor U12716 (N_12716,N_12176,N_12111);
and U12717 (N_12717,N_12326,N_12441);
xor U12718 (N_12718,N_12421,N_12057);
or U12719 (N_12719,N_12407,N_12064);
nor U12720 (N_12720,N_12196,N_12038);
nand U12721 (N_12721,N_12209,N_12099);
and U12722 (N_12722,N_12390,N_12310);
or U12723 (N_12723,N_12203,N_12156);
and U12724 (N_12724,N_12021,N_12486);
or U12725 (N_12725,N_12477,N_12414);
nand U12726 (N_12726,N_12391,N_12063);
xnor U12727 (N_12727,N_12010,N_12374);
or U12728 (N_12728,N_12050,N_12373);
or U12729 (N_12729,N_12498,N_12353);
nand U12730 (N_12730,N_12400,N_12261);
or U12731 (N_12731,N_12419,N_12436);
xor U12732 (N_12732,N_12191,N_12328);
and U12733 (N_12733,N_12327,N_12275);
or U12734 (N_12734,N_12311,N_12364);
and U12735 (N_12735,N_12215,N_12162);
nor U12736 (N_12736,N_12325,N_12065);
and U12737 (N_12737,N_12397,N_12066);
nand U12738 (N_12738,N_12345,N_12134);
or U12739 (N_12739,N_12022,N_12142);
or U12740 (N_12740,N_12084,N_12445);
nand U12741 (N_12741,N_12051,N_12489);
xor U12742 (N_12742,N_12273,N_12120);
xnor U12743 (N_12743,N_12346,N_12448);
and U12744 (N_12744,N_12243,N_12139);
nand U12745 (N_12745,N_12069,N_12306);
or U12746 (N_12746,N_12027,N_12029);
nor U12747 (N_12747,N_12202,N_12282);
and U12748 (N_12748,N_12321,N_12119);
nand U12749 (N_12749,N_12053,N_12404);
nand U12750 (N_12750,N_12191,N_12313);
nand U12751 (N_12751,N_12068,N_12048);
or U12752 (N_12752,N_12344,N_12478);
nand U12753 (N_12753,N_12422,N_12448);
nand U12754 (N_12754,N_12219,N_12389);
xnor U12755 (N_12755,N_12298,N_12425);
nand U12756 (N_12756,N_12492,N_12240);
or U12757 (N_12757,N_12277,N_12017);
nand U12758 (N_12758,N_12365,N_12068);
xor U12759 (N_12759,N_12227,N_12087);
and U12760 (N_12760,N_12044,N_12348);
and U12761 (N_12761,N_12376,N_12466);
or U12762 (N_12762,N_12303,N_12308);
nor U12763 (N_12763,N_12053,N_12364);
xnor U12764 (N_12764,N_12094,N_12434);
xnor U12765 (N_12765,N_12072,N_12034);
nand U12766 (N_12766,N_12224,N_12085);
or U12767 (N_12767,N_12494,N_12142);
nand U12768 (N_12768,N_12441,N_12055);
nor U12769 (N_12769,N_12463,N_12347);
nor U12770 (N_12770,N_12297,N_12293);
xor U12771 (N_12771,N_12164,N_12015);
or U12772 (N_12772,N_12371,N_12061);
nand U12773 (N_12773,N_12219,N_12028);
or U12774 (N_12774,N_12209,N_12210);
and U12775 (N_12775,N_12239,N_12395);
and U12776 (N_12776,N_12276,N_12375);
or U12777 (N_12777,N_12096,N_12437);
xor U12778 (N_12778,N_12335,N_12189);
and U12779 (N_12779,N_12206,N_12253);
xor U12780 (N_12780,N_12018,N_12098);
nor U12781 (N_12781,N_12320,N_12173);
nor U12782 (N_12782,N_12437,N_12111);
nand U12783 (N_12783,N_12056,N_12023);
or U12784 (N_12784,N_12424,N_12301);
nand U12785 (N_12785,N_12077,N_12076);
nor U12786 (N_12786,N_12410,N_12131);
nand U12787 (N_12787,N_12080,N_12356);
or U12788 (N_12788,N_12267,N_12006);
xor U12789 (N_12789,N_12467,N_12248);
nand U12790 (N_12790,N_12342,N_12007);
nand U12791 (N_12791,N_12192,N_12147);
nor U12792 (N_12792,N_12350,N_12453);
or U12793 (N_12793,N_12396,N_12030);
xnor U12794 (N_12794,N_12143,N_12037);
nor U12795 (N_12795,N_12056,N_12121);
nor U12796 (N_12796,N_12345,N_12196);
and U12797 (N_12797,N_12112,N_12191);
nand U12798 (N_12798,N_12449,N_12298);
xor U12799 (N_12799,N_12036,N_12307);
xor U12800 (N_12800,N_12145,N_12144);
and U12801 (N_12801,N_12215,N_12262);
nor U12802 (N_12802,N_12133,N_12096);
nor U12803 (N_12803,N_12404,N_12424);
and U12804 (N_12804,N_12406,N_12319);
nor U12805 (N_12805,N_12241,N_12144);
nand U12806 (N_12806,N_12184,N_12404);
and U12807 (N_12807,N_12320,N_12383);
or U12808 (N_12808,N_12230,N_12259);
xor U12809 (N_12809,N_12029,N_12238);
xnor U12810 (N_12810,N_12318,N_12180);
or U12811 (N_12811,N_12035,N_12046);
nand U12812 (N_12812,N_12470,N_12066);
nand U12813 (N_12813,N_12485,N_12055);
and U12814 (N_12814,N_12351,N_12223);
nor U12815 (N_12815,N_12104,N_12295);
nor U12816 (N_12816,N_12440,N_12347);
nor U12817 (N_12817,N_12153,N_12480);
xor U12818 (N_12818,N_12295,N_12443);
and U12819 (N_12819,N_12118,N_12460);
and U12820 (N_12820,N_12395,N_12096);
or U12821 (N_12821,N_12223,N_12398);
or U12822 (N_12822,N_12225,N_12088);
or U12823 (N_12823,N_12125,N_12421);
or U12824 (N_12824,N_12364,N_12480);
or U12825 (N_12825,N_12041,N_12292);
xnor U12826 (N_12826,N_12339,N_12360);
nor U12827 (N_12827,N_12349,N_12108);
or U12828 (N_12828,N_12364,N_12218);
nor U12829 (N_12829,N_12121,N_12030);
and U12830 (N_12830,N_12405,N_12097);
and U12831 (N_12831,N_12039,N_12011);
nor U12832 (N_12832,N_12105,N_12208);
nor U12833 (N_12833,N_12422,N_12379);
or U12834 (N_12834,N_12072,N_12326);
or U12835 (N_12835,N_12294,N_12075);
or U12836 (N_12836,N_12452,N_12125);
or U12837 (N_12837,N_12073,N_12034);
or U12838 (N_12838,N_12336,N_12281);
nand U12839 (N_12839,N_12423,N_12486);
and U12840 (N_12840,N_12484,N_12463);
xor U12841 (N_12841,N_12075,N_12259);
nand U12842 (N_12842,N_12155,N_12069);
and U12843 (N_12843,N_12430,N_12369);
nor U12844 (N_12844,N_12232,N_12096);
xnor U12845 (N_12845,N_12245,N_12312);
and U12846 (N_12846,N_12403,N_12444);
xnor U12847 (N_12847,N_12046,N_12218);
and U12848 (N_12848,N_12175,N_12282);
or U12849 (N_12849,N_12245,N_12229);
and U12850 (N_12850,N_12487,N_12287);
and U12851 (N_12851,N_12185,N_12152);
xor U12852 (N_12852,N_12237,N_12217);
and U12853 (N_12853,N_12263,N_12210);
or U12854 (N_12854,N_12277,N_12316);
xor U12855 (N_12855,N_12214,N_12068);
nand U12856 (N_12856,N_12303,N_12416);
xnor U12857 (N_12857,N_12052,N_12384);
nor U12858 (N_12858,N_12096,N_12453);
and U12859 (N_12859,N_12118,N_12469);
or U12860 (N_12860,N_12408,N_12188);
nand U12861 (N_12861,N_12111,N_12252);
and U12862 (N_12862,N_12261,N_12237);
or U12863 (N_12863,N_12251,N_12210);
nor U12864 (N_12864,N_12307,N_12443);
nand U12865 (N_12865,N_12047,N_12495);
or U12866 (N_12866,N_12270,N_12326);
and U12867 (N_12867,N_12301,N_12195);
xnor U12868 (N_12868,N_12372,N_12312);
xnor U12869 (N_12869,N_12348,N_12161);
and U12870 (N_12870,N_12162,N_12368);
and U12871 (N_12871,N_12369,N_12421);
nand U12872 (N_12872,N_12314,N_12125);
nand U12873 (N_12873,N_12375,N_12222);
or U12874 (N_12874,N_12021,N_12094);
nand U12875 (N_12875,N_12320,N_12163);
nor U12876 (N_12876,N_12331,N_12259);
nand U12877 (N_12877,N_12462,N_12045);
nand U12878 (N_12878,N_12336,N_12390);
or U12879 (N_12879,N_12064,N_12010);
xor U12880 (N_12880,N_12383,N_12260);
and U12881 (N_12881,N_12341,N_12250);
nand U12882 (N_12882,N_12260,N_12202);
xor U12883 (N_12883,N_12216,N_12443);
and U12884 (N_12884,N_12214,N_12131);
nor U12885 (N_12885,N_12372,N_12344);
nor U12886 (N_12886,N_12109,N_12201);
nor U12887 (N_12887,N_12258,N_12022);
and U12888 (N_12888,N_12305,N_12010);
nor U12889 (N_12889,N_12425,N_12257);
or U12890 (N_12890,N_12286,N_12277);
nor U12891 (N_12891,N_12381,N_12102);
or U12892 (N_12892,N_12281,N_12268);
xnor U12893 (N_12893,N_12252,N_12482);
or U12894 (N_12894,N_12326,N_12296);
nor U12895 (N_12895,N_12130,N_12317);
nand U12896 (N_12896,N_12273,N_12011);
or U12897 (N_12897,N_12333,N_12439);
and U12898 (N_12898,N_12266,N_12033);
nand U12899 (N_12899,N_12211,N_12038);
nor U12900 (N_12900,N_12074,N_12077);
nor U12901 (N_12901,N_12049,N_12186);
and U12902 (N_12902,N_12156,N_12059);
and U12903 (N_12903,N_12309,N_12338);
nand U12904 (N_12904,N_12111,N_12321);
xor U12905 (N_12905,N_12406,N_12382);
nor U12906 (N_12906,N_12483,N_12312);
xor U12907 (N_12907,N_12459,N_12465);
or U12908 (N_12908,N_12169,N_12449);
nor U12909 (N_12909,N_12493,N_12299);
nand U12910 (N_12910,N_12209,N_12165);
nand U12911 (N_12911,N_12022,N_12283);
nand U12912 (N_12912,N_12453,N_12320);
xnor U12913 (N_12913,N_12326,N_12498);
and U12914 (N_12914,N_12238,N_12047);
nor U12915 (N_12915,N_12118,N_12392);
and U12916 (N_12916,N_12452,N_12022);
xor U12917 (N_12917,N_12445,N_12381);
nor U12918 (N_12918,N_12116,N_12045);
xor U12919 (N_12919,N_12386,N_12280);
nand U12920 (N_12920,N_12418,N_12365);
or U12921 (N_12921,N_12351,N_12050);
or U12922 (N_12922,N_12401,N_12338);
and U12923 (N_12923,N_12156,N_12358);
or U12924 (N_12924,N_12076,N_12362);
xor U12925 (N_12925,N_12148,N_12439);
nor U12926 (N_12926,N_12447,N_12132);
xnor U12927 (N_12927,N_12488,N_12037);
and U12928 (N_12928,N_12366,N_12284);
nor U12929 (N_12929,N_12300,N_12495);
or U12930 (N_12930,N_12444,N_12011);
nor U12931 (N_12931,N_12191,N_12141);
nand U12932 (N_12932,N_12389,N_12112);
nor U12933 (N_12933,N_12413,N_12268);
and U12934 (N_12934,N_12391,N_12416);
xor U12935 (N_12935,N_12296,N_12409);
xor U12936 (N_12936,N_12474,N_12023);
and U12937 (N_12937,N_12333,N_12016);
and U12938 (N_12938,N_12314,N_12439);
xnor U12939 (N_12939,N_12118,N_12474);
nand U12940 (N_12940,N_12210,N_12315);
nand U12941 (N_12941,N_12367,N_12161);
and U12942 (N_12942,N_12330,N_12381);
xnor U12943 (N_12943,N_12440,N_12277);
nand U12944 (N_12944,N_12130,N_12465);
and U12945 (N_12945,N_12007,N_12488);
and U12946 (N_12946,N_12431,N_12396);
xor U12947 (N_12947,N_12030,N_12198);
nand U12948 (N_12948,N_12288,N_12487);
or U12949 (N_12949,N_12309,N_12000);
or U12950 (N_12950,N_12051,N_12419);
nand U12951 (N_12951,N_12212,N_12430);
or U12952 (N_12952,N_12356,N_12021);
or U12953 (N_12953,N_12316,N_12460);
or U12954 (N_12954,N_12029,N_12067);
xor U12955 (N_12955,N_12271,N_12425);
nand U12956 (N_12956,N_12472,N_12122);
nor U12957 (N_12957,N_12331,N_12126);
nor U12958 (N_12958,N_12459,N_12143);
or U12959 (N_12959,N_12061,N_12099);
nand U12960 (N_12960,N_12430,N_12077);
nand U12961 (N_12961,N_12090,N_12171);
and U12962 (N_12962,N_12278,N_12061);
nor U12963 (N_12963,N_12267,N_12099);
or U12964 (N_12964,N_12119,N_12423);
xnor U12965 (N_12965,N_12452,N_12353);
or U12966 (N_12966,N_12370,N_12425);
nor U12967 (N_12967,N_12346,N_12324);
or U12968 (N_12968,N_12237,N_12388);
nand U12969 (N_12969,N_12096,N_12255);
or U12970 (N_12970,N_12184,N_12003);
xnor U12971 (N_12971,N_12067,N_12162);
and U12972 (N_12972,N_12406,N_12190);
nand U12973 (N_12973,N_12416,N_12462);
xnor U12974 (N_12974,N_12270,N_12082);
or U12975 (N_12975,N_12434,N_12135);
nor U12976 (N_12976,N_12484,N_12039);
nor U12977 (N_12977,N_12340,N_12031);
and U12978 (N_12978,N_12084,N_12196);
or U12979 (N_12979,N_12174,N_12169);
xor U12980 (N_12980,N_12215,N_12450);
nor U12981 (N_12981,N_12291,N_12097);
and U12982 (N_12982,N_12114,N_12271);
and U12983 (N_12983,N_12184,N_12491);
xnor U12984 (N_12984,N_12016,N_12014);
and U12985 (N_12985,N_12348,N_12255);
nor U12986 (N_12986,N_12070,N_12159);
xor U12987 (N_12987,N_12418,N_12303);
and U12988 (N_12988,N_12282,N_12145);
nand U12989 (N_12989,N_12491,N_12171);
and U12990 (N_12990,N_12133,N_12121);
nor U12991 (N_12991,N_12245,N_12179);
or U12992 (N_12992,N_12096,N_12361);
or U12993 (N_12993,N_12442,N_12112);
and U12994 (N_12994,N_12363,N_12021);
nand U12995 (N_12995,N_12491,N_12115);
nor U12996 (N_12996,N_12306,N_12337);
and U12997 (N_12997,N_12222,N_12336);
and U12998 (N_12998,N_12448,N_12093);
or U12999 (N_12999,N_12372,N_12034);
nand U13000 (N_13000,N_12795,N_12925);
xor U13001 (N_13001,N_12882,N_12865);
and U13002 (N_13002,N_12919,N_12562);
nand U13003 (N_13003,N_12635,N_12935);
nor U13004 (N_13004,N_12716,N_12813);
nor U13005 (N_13005,N_12937,N_12887);
and U13006 (N_13006,N_12689,N_12654);
nand U13007 (N_13007,N_12845,N_12632);
nor U13008 (N_13008,N_12672,N_12675);
or U13009 (N_13009,N_12659,N_12761);
nor U13010 (N_13010,N_12709,N_12713);
nand U13011 (N_13011,N_12758,N_12793);
and U13012 (N_13012,N_12950,N_12508);
or U13013 (N_13013,N_12993,N_12856);
xnor U13014 (N_13014,N_12754,N_12613);
or U13015 (N_13015,N_12696,N_12712);
and U13016 (N_13016,N_12658,N_12584);
and U13017 (N_13017,N_12665,N_12851);
xnor U13018 (N_13018,N_12759,N_12888);
xor U13019 (N_13019,N_12999,N_12634);
and U13020 (N_13020,N_12973,N_12738);
and U13021 (N_13021,N_12647,N_12829);
nand U13022 (N_13022,N_12799,N_12768);
or U13023 (N_13023,N_12818,N_12775);
xor U13024 (N_13024,N_12790,N_12593);
nand U13025 (N_13025,N_12830,N_12837);
and U13026 (N_13026,N_12792,N_12869);
nand U13027 (N_13027,N_12653,N_12587);
nand U13028 (N_13028,N_12745,N_12638);
or U13029 (N_13029,N_12827,N_12966);
nand U13030 (N_13030,N_12940,N_12987);
nor U13031 (N_13031,N_12522,N_12552);
nand U13032 (N_13032,N_12782,N_12605);
or U13033 (N_13033,N_12988,N_12868);
or U13034 (N_13034,N_12661,N_12626);
xor U13035 (N_13035,N_12542,N_12688);
or U13036 (N_13036,N_12747,N_12867);
and U13037 (N_13037,N_12556,N_12540);
nand U13038 (N_13038,N_12763,N_12524);
or U13039 (N_13039,N_12534,N_12518);
nand U13040 (N_13040,N_12916,N_12872);
nand U13041 (N_13041,N_12915,N_12591);
nor U13042 (N_13042,N_12734,N_12907);
or U13043 (N_13043,N_12791,N_12733);
or U13044 (N_13044,N_12998,N_12929);
nor U13045 (N_13045,N_12670,N_12992);
nor U13046 (N_13046,N_12525,N_12978);
xor U13047 (N_13047,N_12994,N_12578);
or U13048 (N_13048,N_12895,N_12980);
or U13049 (N_13049,N_12585,N_12560);
or U13050 (N_13050,N_12558,N_12913);
xor U13051 (N_13051,N_12510,N_12532);
xor U13052 (N_13052,N_12678,N_12655);
or U13053 (N_13053,N_12970,N_12611);
or U13054 (N_13054,N_12595,N_12928);
or U13055 (N_13055,N_12769,N_12676);
nor U13056 (N_13056,N_12668,N_12590);
nand U13057 (N_13057,N_12543,N_12983);
nor U13058 (N_13058,N_12581,N_12765);
or U13059 (N_13059,N_12722,N_12669);
nor U13060 (N_13060,N_12615,N_12779);
xnor U13061 (N_13061,N_12840,N_12896);
nor U13062 (N_13062,N_12707,N_12643);
and U13063 (N_13063,N_12912,N_12890);
nand U13064 (N_13064,N_12640,N_12772);
nand U13065 (N_13065,N_12570,N_12774);
xnor U13066 (N_13066,N_12566,N_12897);
xnor U13067 (N_13067,N_12930,N_12677);
nand U13068 (N_13068,N_12971,N_12691);
and U13069 (N_13069,N_12721,N_12723);
nor U13070 (N_13070,N_12652,N_12697);
or U13071 (N_13071,N_12833,N_12648);
nand U13072 (N_13072,N_12683,N_12523);
or U13073 (N_13073,N_12923,N_12870);
nand U13074 (N_13074,N_12748,N_12931);
nand U13075 (N_13075,N_12776,N_12876);
and U13076 (N_13076,N_12730,N_12807);
nor U13077 (N_13077,N_12981,N_12711);
or U13078 (N_13078,N_12736,N_12719);
nand U13079 (N_13079,N_12943,N_12760);
nor U13080 (N_13080,N_12603,N_12602);
nor U13081 (N_13081,N_12700,N_12571);
xor U13082 (N_13082,N_12618,N_12519);
or U13083 (N_13083,N_12873,N_12500);
nor U13084 (N_13084,N_12898,N_12918);
or U13085 (N_13085,N_12936,N_12520);
nor U13086 (N_13086,N_12892,N_12811);
nand U13087 (N_13087,N_12503,N_12732);
nand U13088 (N_13088,N_12803,N_12942);
xor U13089 (N_13089,N_12710,N_12666);
xnor U13090 (N_13090,N_12617,N_12563);
and U13091 (N_13091,N_12586,N_12901);
xnor U13092 (N_13092,N_12752,N_12974);
xor U13093 (N_13093,N_12854,N_12914);
nand U13094 (N_13094,N_12908,N_12825);
and U13095 (N_13095,N_12592,N_12903);
nand U13096 (N_13096,N_12588,N_12694);
or U13097 (N_13097,N_12924,N_12798);
and U13098 (N_13098,N_12857,N_12706);
nand U13099 (N_13099,N_12598,N_12961);
or U13100 (N_13100,N_12991,N_12783);
nor U13101 (N_13101,N_12742,N_12815);
nand U13102 (N_13102,N_12878,N_12695);
nor U13103 (N_13103,N_12601,N_12743);
nor U13104 (N_13104,N_12607,N_12885);
or U13105 (N_13105,N_12997,N_12954);
and U13106 (N_13106,N_12881,N_12687);
or U13107 (N_13107,N_12649,N_12836);
nand U13108 (N_13108,N_12548,N_12662);
xor U13109 (N_13109,N_12597,N_12846);
nand U13110 (N_13110,N_12853,N_12725);
or U13111 (N_13111,N_12554,N_12656);
xor U13112 (N_13112,N_12546,N_12679);
nand U13113 (N_13113,N_12664,N_12989);
nand U13114 (N_13114,N_12708,N_12911);
nand U13115 (N_13115,N_12977,N_12660);
nor U13116 (N_13116,N_12979,N_12816);
and U13117 (N_13117,N_12506,N_12619);
nor U13118 (N_13118,N_12951,N_12651);
or U13119 (N_13119,N_12841,N_12968);
nor U13120 (N_13120,N_12606,N_12746);
and U13121 (N_13121,N_12850,N_12729);
and U13122 (N_13122,N_12849,N_12513);
xor U13123 (N_13123,N_12533,N_12749);
nor U13124 (N_13124,N_12879,N_12812);
xor U13125 (N_13125,N_12555,N_12703);
nor U13126 (N_13126,N_12757,N_12528);
nor U13127 (N_13127,N_12629,N_12639);
or U13128 (N_13128,N_12835,N_12701);
or U13129 (N_13129,N_12727,N_12766);
nand U13130 (N_13130,N_12671,N_12526);
nor U13131 (N_13131,N_12947,N_12777);
and U13132 (N_13132,N_12735,N_12577);
and U13133 (N_13133,N_12753,N_12904);
nand U13134 (N_13134,N_12692,N_12990);
nor U13135 (N_13135,N_12612,N_12704);
xnor U13136 (N_13136,N_12820,N_12610);
nor U13137 (N_13137,N_12899,N_12614);
xnor U13138 (N_13138,N_12511,N_12957);
and U13139 (N_13139,N_12788,N_12941);
and U13140 (N_13140,N_12580,N_12860);
nand U13141 (N_13141,N_12564,N_12646);
and U13142 (N_13142,N_12995,N_12718);
or U13143 (N_13143,N_12547,N_12608);
and U13144 (N_13144,N_12819,N_12814);
and U13145 (N_13145,N_12535,N_12985);
nand U13146 (N_13146,N_12673,N_12778);
or U13147 (N_13147,N_12559,N_12568);
nor U13148 (N_13148,N_12663,N_12502);
xnor U13149 (N_13149,N_12826,N_12515);
or U13150 (N_13150,N_12946,N_12644);
and U13151 (N_13151,N_12862,N_12567);
nor U13152 (N_13152,N_12859,N_12622);
nor U13153 (N_13153,N_12573,N_12685);
xor U13154 (N_13154,N_12623,N_12844);
nand U13155 (N_13155,N_12986,N_12797);
and U13156 (N_13156,N_12786,N_12955);
or U13157 (N_13157,N_12805,N_12604);
and U13158 (N_13158,N_12575,N_12501);
and U13159 (N_13159,N_12529,N_12910);
nand U13160 (N_13160,N_12949,N_12698);
or U13161 (N_13161,N_12855,N_12726);
nor U13162 (N_13162,N_12938,N_12674);
xor U13163 (N_13163,N_12530,N_12893);
or U13164 (N_13164,N_12982,N_12737);
xor U13165 (N_13165,N_12969,N_12902);
nand U13166 (N_13166,N_12886,N_12963);
xor U13167 (N_13167,N_12883,N_12964);
nor U13168 (N_13168,N_12787,N_12544);
nand U13169 (N_13169,N_12731,N_12541);
and U13170 (N_13170,N_12545,N_12802);
nand U13171 (N_13171,N_12636,N_12616);
nand U13172 (N_13172,N_12582,N_12891);
xnor U13173 (N_13173,N_12509,N_12953);
nand U13174 (N_13174,N_12516,N_12702);
nor U13175 (N_13175,N_12962,N_12771);
nor U13176 (N_13176,N_12756,N_12875);
and U13177 (N_13177,N_12627,N_12959);
and U13178 (N_13178,N_12939,N_12565);
and U13179 (N_13179,N_12569,N_12794);
nand U13180 (N_13180,N_12861,N_12682);
nor U13181 (N_13181,N_12699,N_12945);
and U13182 (N_13182,N_12823,N_12877);
nor U13183 (N_13183,N_12822,N_12621);
or U13184 (N_13184,N_12975,N_12842);
xor U13185 (N_13185,N_12905,N_12667);
nor U13186 (N_13186,N_12641,N_12848);
xnor U13187 (N_13187,N_12537,N_12740);
nand U13188 (N_13188,N_12517,N_12839);
xnor U13189 (N_13189,N_12917,N_12847);
nor U13190 (N_13190,N_12583,N_12789);
or U13191 (N_13191,N_12972,N_12576);
nor U13192 (N_13192,N_12755,N_12921);
nor U13193 (N_13193,N_12926,N_12838);
nand U13194 (N_13194,N_12681,N_12852);
and U13195 (N_13195,N_12549,N_12630);
nand U13196 (N_13196,N_12531,N_12810);
nor U13197 (N_13197,N_12657,N_12631);
nand U13198 (N_13198,N_12960,N_12934);
xor U13199 (N_13199,N_12828,N_12967);
nor U13200 (N_13200,N_12650,N_12680);
and U13201 (N_13201,N_12507,N_12801);
or U13202 (N_13202,N_12884,N_12965);
and U13203 (N_13203,N_12714,N_12684);
or U13204 (N_13204,N_12633,N_12693);
xor U13205 (N_13205,N_12809,N_12843);
nor U13206 (N_13206,N_12767,N_12894);
nand U13207 (N_13207,N_12609,N_12817);
and U13208 (N_13208,N_12620,N_12889);
nand U13209 (N_13209,N_12858,N_12958);
or U13210 (N_13210,N_12728,N_12762);
xor U13211 (N_13211,N_12832,N_12637);
or U13212 (N_13212,N_12773,N_12864);
nor U13213 (N_13213,N_12821,N_12900);
nand U13214 (N_13214,N_12521,N_12922);
xnor U13215 (N_13215,N_12785,N_12505);
nor U13216 (N_13216,N_12834,N_12645);
or U13217 (N_13217,N_12512,N_12538);
nor U13218 (N_13218,N_12624,N_12984);
nor U13219 (N_13219,N_12690,N_12539);
or U13220 (N_13220,N_12956,N_12804);
xnor U13221 (N_13221,N_12589,N_12866);
or U13222 (N_13222,N_12909,N_12599);
and U13223 (N_13223,N_12504,N_12806);
and U13224 (N_13224,N_12600,N_12741);
nor U13225 (N_13225,N_12553,N_12550);
nor U13226 (N_13226,N_12932,N_12551);
nand U13227 (N_13227,N_12944,N_12720);
nor U13228 (N_13228,N_12780,N_12750);
nor U13229 (N_13229,N_12642,N_12863);
nand U13230 (N_13230,N_12800,N_12831);
and U13231 (N_13231,N_12724,N_12557);
nor U13232 (N_13232,N_12561,N_12781);
xor U13233 (N_13233,N_12976,N_12784);
or U13234 (N_13234,N_12625,N_12715);
nor U13235 (N_13235,N_12764,N_12594);
xnor U13236 (N_13236,N_12927,N_12574);
xnor U13237 (N_13237,N_12744,N_12596);
xor U13238 (N_13238,N_12579,N_12920);
xor U13239 (N_13239,N_12686,N_12572);
nand U13240 (N_13240,N_12933,N_12871);
and U13241 (N_13241,N_12952,N_12751);
or U13242 (N_13242,N_12527,N_12906);
or U13243 (N_13243,N_12705,N_12874);
xnor U13244 (N_13244,N_12536,N_12808);
xnor U13245 (N_13245,N_12739,N_12796);
xor U13246 (N_13246,N_12996,N_12824);
and U13247 (N_13247,N_12948,N_12514);
or U13248 (N_13248,N_12628,N_12770);
nor U13249 (N_13249,N_12880,N_12717);
and U13250 (N_13250,N_12698,N_12609);
and U13251 (N_13251,N_12935,N_12787);
nor U13252 (N_13252,N_12837,N_12508);
or U13253 (N_13253,N_12753,N_12615);
nand U13254 (N_13254,N_12564,N_12666);
nor U13255 (N_13255,N_12843,N_12954);
xor U13256 (N_13256,N_12524,N_12737);
nor U13257 (N_13257,N_12705,N_12913);
nor U13258 (N_13258,N_12715,N_12942);
nor U13259 (N_13259,N_12677,N_12864);
xnor U13260 (N_13260,N_12793,N_12572);
xnor U13261 (N_13261,N_12736,N_12746);
xor U13262 (N_13262,N_12599,N_12634);
or U13263 (N_13263,N_12695,N_12544);
or U13264 (N_13264,N_12707,N_12870);
xnor U13265 (N_13265,N_12975,N_12837);
nand U13266 (N_13266,N_12689,N_12675);
nand U13267 (N_13267,N_12697,N_12929);
nand U13268 (N_13268,N_12553,N_12932);
and U13269 (N_13269,N_12944,N_12599);
nor U13270 (N_13270,N_12547,N_12515);
or U13271 (N_13271,N_12749,N_12837);
nor U13272 (N_13272,N_12692,N_12684);
or U13273 (N_13273,N_12599,N_12555);
xor U13274 (N_13274,N_12774,N_12530);
nand U13275 (N_13275,N_12522,N_12707);
xor U13276 (N_13276,N_12875,N_12663);
xnor U13277 (N_13277,N_12703,N_12878);
and U13278 (N_13278,N_12790,N_12983);
and U13279 (N_13279,N_12804,N_12594);
and U13280 (N_13280,N_12625,N_12548);
xor U13281 (N_13281,N_12546,N_12687);
and U13282 (N_13282,N_12644,N_12887);
or U13283 (N_13283,N_12597,N_12952);
and U13284 (N_13284,N_12545,N_12739);
xor U13285 (N_13285,N_12932,N_12691);
and U13286 (N_13286,N_12898,N_12635);
or U13287 (N_13287,N_12903,N_12582);
or U13288 (N_13288,N_12721,N_12554);
xor U13289 (N_13289,N_12883,N_12959);
or U13290 (N_13290,N_12659,N_12519);
xnor U13291 (N_13291,N_12583,N_12845);
nand U13292 (N_13292,N_12543,N_12612);
and U13293 (N_13293,N_12883,N_12886);
or U13294 (N_13294,N_12759,N_12913);
and U13295 (N_13295,N_12849,N_12917);
nand U13296 (N_13296,N_12794,N_12558);
nor U13297 (N_13297,N_12702,N_12691);
or U13298 (N_13298,N_12894,N_12686);
xor U13299 (N_13299,N_12601,N_12902);
nor U13300 (N_13300,N_12635,N_12698);
or U13301 (N_13301,N_12640,N_12843);
nand U13302 (N_13302,N_12664,N_12861);
nand U13303 (N_13303,N_12794,N_12701);
or U13304 (N_13304,N_12641,N_12696);
or U13305 (N_13305,N_12606,N_12501);
and U13306 (N_13306,N_12867,N_12695);
nand U13307 (N_13307,N_12826,N_12925);
xor U13308 (N_13308,N_12548,N_12829);
nor U13309 (N_13309,N_12508,N_12501);
xor U13310 (N_13310,N_12592,N_12522);
or U13311 (N_13311,N_12569,N_12533);
nor U13312 (N_13312,N_12809,N_12639);
or U13313 (N_13313,N_12811,N_12502);
nand U13314 (N_13314,N_12739,N_12907);
and U13315 (N_13315,N_12913,N_12631);
xor U13316 (N_13316,N_12794,N_12574);
or U13317 (N_13317,N_12509,N_12949);
and U13318 (N_13318,N_12742,N_12500);
or U13319 (N_13319,N_12730,N_12805);
nor U13320 (N_13320,N_12826,N_12678);
nor U13321 (N_13321,N_12850,N_12617);
nor U13322 (N_13322,N_12863,N_12765);
nor U13323 (N_13323,N_12869,N_12532);
or U13324 (N_13324,N_12914,N_12971);
and U13325 (N_13325,N_12764,N_12670);
nor U13326 (N_13326,N_12983,N_12763);
and U13327 (N_13327,N_12947,N_12839);
or U13328 (N_13328,N_12506,N_12569);
nand U13329 (N_13329,N_12541,N_12869);
xnor U13330 (N_13330,N_12773,N_12768);
and U13331 (N_13331,N_12930,N_12626);
nand U13332 (N_13332,N_12791,N_12506);
nand U13333 (N_13333,N_12557,N_12635);
xnor U13334 (N_13334,N_12917,N_12714);
and U13335 (N_13335,N_12569,N_12711);
xor U13336 (N_13336,N_12665,N_12567);
and U13337 (N_13337,N_12622,N_12831);
nor U13338 (N_13338,N_12912,N_12795);
and U13339 (N_13339,N_12594,N_12954);
nor U13340 (N_13340,N_12641,N_12561);
and U13341 (N_13341,N_12987,N_12957);
xor U13342 (N_13342,N_12642,N_12836);
and U13343 (N_13343,N_12884,N_12546);
or U13344 (N_13344,N_12841,N_12719);
nor U13345 (N_13345,N_12997,N_12553);
and U13346 (N_13346,N_12850,N_12942);
nor U13347 (N_13347,N_12765,N_12959);
nor U13348 (N_13348,N_12694,N_12966);
and U13349 (N_13349,N_12642,N_12782);
nand U13350 (N_13350,N_12900,N_12816);
xor U13351 (N_13351,N_12909,N_12743);
xnor U13352 (N_13352,N_12744,N_12517);
or U13353 (N_13353,N_12666,N_12558);
nand U13354 (N_13354,N_12913,N_12532);
nand U13355 (N_13355,N_12777,N_12878);
nor U13356 (N_13356,N_12890,N_12608);
or U13357 (N_13357,N_12810,N_12826);
nand U13358 (N_13358,N_12951,N_12932);
or U13359 (N_13359,N_12995,N_12775);
and U13360 (N_13360,N_12661,N_12971);
nor U13361 (N_13361,N_12945,N_12574);
nand U13362 (N_13362,N_12898,N_12904);
nand U13363 (N_13363,N_12621,N_12704);
and U13364 (N_13364,N_12896,N_12576);
nand U13365 (N_13365,N_12682,N_12925);
or U13366 (N_13366,N_12552,N_12619);
nand U13367 (N_13367,N_12776,N_12637);
nor U13368 (N_13368,N_12938,N_12966);
nor U13369 (N_13369,N_12524,N_12938);
nand U13370 (N_13370,N_12634,N_12532);
xor U13371 (N_13371,N_12679,N_12502);
nand U13372 (N_13372,N_12752,N_12608);
nand U13373 (N_13373,N_12780,N_12902);
xnor U13374 (N_13374,N_12754,N_12925);
nor U13375 (N_13375,N_12797,N_12677);
xnor U13376 (N_13376,N_12559,N_12545);
and U13377 (N_13377,N_12831,N_12834);
or U13378 (N_13378,N_12950,N_12989);
and U13379 (N_13379,N_12813,N_12660);
xor U13380 (N_13380,N_12566,N_12585);
nand U13381 (N_13381,N_12584,N_12992);
nand U13382 (N_13382,N_12579,N_12855);
and U13383 (N_13383,N_12772,N_12698);
and U13384 (N_13384,N_12726,N_12830);
or U13385 (N_13385,N_12689,N_12908);
and U13386 (N_13386,N_12689,N_12922);
or U13387 (N_13387,N_12541,N_12605);
and U13388 (N_13388,N_12668,N_12910);
xor U13389 (N_13389,N_12870,N_12614);
and U13390 (N_13390,N_12962,N_12614);
nand U13391 (N_13391,N_12737,N_12777);
nand U13392 (N_13392,N_12938,N_12555);
xor U13393 (N_13393,N_12737,N_12948);
nand U13394 (N_13394,N_12594,N_12987);
xor U13395 (N_13395,N_12974,N_12697);
and U13396 (N_13396,N_12903,N_12852);
and U13397 (N_13397,N_12612,N_12859);
and U13398 (N_13398,N_12592,N_12507);
or U13399 (N_13399,N_12935,N_12975);
nand U13400 (N_13400,N_12910,N_12539);
nand U13401 (N_13401,N_12537,N_12718);
and U13402 (N_13402,N_12994,N_12704);
and U13403 (N_13403,N_12515,N_12586);
and U13404 (N_13404,N_12725,N_12693);
xnor U13405 (N_13405,N_12628,N_12675);
or U13406 (N_13406,N_12960,N_12534);
and U13407 (N_13407,N_12961,N_12534);
and U13408 (N_13408,N_12933,N_12607);
xor U13409 (N_13409,N_12868,N_12842);
xor U13410 (N_13410,N_12985,N_12771);
xor U13411 (N_13411,N_12945,N_12625);
or U13412 (N_13412,N_12796,N_12669);
or U13413 (N_13413,N_12874,N_12986);
nand U13414 (N_13414,N_12775,N_12514);
and U13415 (N_13415,N_12826,N_12537);
or U13416 (N_13416,N_12923,N_12710);
or U13417 (N_13417,N_12513,N_12525);
and U13418 (N_13418,N_12577,N_12503);
nor U13419 (N_13419,N_12932,N_12716);
and U13420 (N_13420,N_12613,N_12667);
nand U13421 (N_13421,N_12827,N_12762);
and U13422 (N_13422,N_12852,N_12764);
nand U13423 (N_13423,N_12731,N_12653);
nand U13424 (N_13424,N_12867,N_12885);
and U13425 (N_13425,N_12823,N_12992);
nand U13426 (N_13426,N_12660,N_12969);
nand U13427 (N_13427,N_12792,N_12803);
nor U13428 (N_13428,N_12951,N_12955);
or U13429 (N_13429,N_12706,N_12613);
and U13430 (N_13430,N_12996,N_12989);
xnor U13431 (N_13431,N_12667,N_12749);
xnor U13432 (N_13432,N_12581,N_12865);
xnor U13433 (N_13433,N_12652,N_12561);
xor U13434 (N_13434,N_12919,N_12577);
or U13435 (N_13435,N_12924,N_12889);
xnor U13436 (N_13436,N_12727,N_12755);
xnor U13437 (N_13437,N_12828,N_12985);
and U13438 (N_13438,N_12618,N_12559);
or U13439 (N_13439,N_12678,N_12641);
nor U13440 (N_13440,N_12524,N_12583);
xnor U13441 (N_13441,N_12504,N_12706);
and U13442 (N_13442,N_12719,N_12992);
xor U13443 (N_13443,N_12932,N_12650);
nor U13444 (N_13444,N_12703,N_12524);
and U13445 (N_13445,N_12523,N_12944);
xnor U13446 (N_13446,N_12806,N_12862);
or U13447 (N_13447,N_12709,N_12929);
nand U13448 (N_13448,N_12592,N_12984);
or U13449 (N_13449,N_12801,N_12658);
xor U13450 (N_13450,N_12993,N_12591);
nor U13451 (N_13451,N_12794,N_12550);
and U13452 (N_13452,N_12911,N_12732);
nor U13453 (N_13453,N_12547,N_12545);
xor U13454 (N_13454,N_12846,N_12878);
nor U13455 (N_13455,N_12795,N_12973);
nor U13456 (N_13456,N_12572,N_12939);
nor U13457 (N_13457,N_12855,N_12863);
or U13458 (N_13458,N_12577,N_12567);
nand U13459 (N_13459,N_12983,N_12954);
and U13460 (N_13460,N_12947,N_12775);
nand U13461 (N_13461,N_12666,N_12795);
or U13462 (N_13462,N_12591,N_12929);
and U13463 (N_13463,N_12673,N_12785);
or U13464 (N_13464,N_12777,N_12847);
nor U13465 (N_13465,N_12687,N_12812);
nand U13466 (N_13466,N_12687,N_12713);
nor U13467 (N_13467,N_12593,N_12545);
and U13468 (N_13468,N_12819,N_12516);
or U13469 (N_13469,N_12678,N_12722);
nor U13470 (N_13470,N_12814,N_12524);
and U13471 (N_13471,N_12751,N_12503);
and U13472 (N_13472,N_12954,N_12510);
and U13473 (N_13473,N_12660,N_12652);
or U13474 (N_13474,N_12805,N_12625);
xor U13475 (N_13475,N_12974,N_12896);
nand U13476 (N_13476,N_12875,N_12717);
and U13477 (N_13477,N_12826,N_12889);
nand U13478 (N_13478,N_12995,N_12972);
and U13479 (N_13479,N_12935,N_12963);
and U13480 (N_13480,N_12998,N_12782);
and U13481 (N_13481,N_12809,N_12650);
and U13482 (N_13482,N_12900,N_12625);
or U13483 (N_13483,N_12691,N_12559);
nand U13484 (N_13484,N_12838,N_12533);
and U13485 (N_13485,N_12979,N_12704);
nand U13486 (N_13486,N_12933,N_12840);
xor U13487 (N_13487,N_12982,N_12537);
or U13488 (N_13488,N_12990,N_12959);
nor U13489 (N_13489,N_12860,N_12907);
xor U13490 (N_13490,N_12643,N_12886);
nor U13491 (N_13491,N_12877,N_12648);
nand U13492 (N_13492,N_12672,N_12734);
nor U13493 (N_13493,N_12745,N_12595);
nor U13494 (N_13494,N_12558,N_12956);
nor U13495 (N_13495,N_12522,N_12943);
nor U13496 (N_13496,N_12695,N_12614);
xnor U13497 (N_13497,N_12818,N_12821);
and U13498 (N_13498,N_12711,N_12849);
nand U13499 (N_13499,N_12899,N_12892);
nor U13500 (N_13500,N_13269,N_13479);
nor U13501 (N_13501,N_13081,N_13340);
or U13502 (N_13502,N_13446,N_13279);
nand U13503 (N_13503,N_13188,N_13149);
nor U13504 (N_13504,N_13096,N_13112);
and U13505 (N_13505,N_13254,N_13068);
xor U13506 (N_13506,N_13304,N_13390);
or U13507 (N_13507,N_13265,N_13418);
nand U13508 (N_13508,N_13318,N_13109);
nor U13509 (N_13509,N_13005,N_13030);
xnor U13510 (N_13510,N_13352,N_13074);
or U13511 (N_13511,N_13031,N_13477);
or U13512 (N_13512,N_13422,N_13399);
xnor U13513 (N_13513,N_13295,N_13305);
and U13514 (N_13514,N_13058,N_13193);
nand U13515 (N_13515,N_13138,N_13206);
or U13516 (N_13516,N_13282,N_13213);
nand U13517 (N_13517,N_13233,N_13065);
and U13518 (N_13518,N_13317,N_13326);
xnor U13519 (N_13519,N_13144,N_13182);
nand U13520 (N_13520,N_13023,N_13143);
and U13521 (N_13521,N_13156,N_13241);
or U13522 (N_13522,N_13272,N_13131);
nand U13523 (N_13523,N_13093,N_13464);
xnor U13524 (N_13524,N_13018,N_13449);
or U13525 (N_13525,N_13245,N_13107);
nand U13526 (N_13526,N_13168,N_13362);
xnor U13527 (N_13527,N_13338,N_13247);
and U13528 (N_13528,N_13255,N_13277);
and U13529 (N_13529,N_13379,N_13171);
nand U13530 (N_13530,N_13169,N_13425);
or U13531 (N_13531,N_13119,N_13121);
nand U13532 (N_13532,N_13437,N_13237);
nor U13533 (N_13533,N_13167,N_13078);
or U13534 (N_13534,N_13000,N_13090);
and U13535 (N_13535,N_13142,N_13110);
nand U13536 (N_13536,N_13336,N_13256);
xnor U13537 (N_13537,N_13072,N_13335);
and U13538 (N_13538,N_13330,N_13079);
and U13539 (N_13539,N_13097,N_13116);
xor U13540 (N_13540,N_13006,N_13176);
or U13541 (N_13541,N_13401,N_13053);
nor U13542 (N_13542,N_13135,N_13315);
xnor U13543 (N_13543,N_13374,N_13498);
and U13544 (N_13544,N_13046,N_13218);
nor U13545 (N_13545,N_13211,N_13025);
nand U13546 (N_13546,N_13219,N_13440);
xor U13547 (N_13547,N_13344,N_13164);
or U13548 (N_13548,N_13044,N_13115);
or U13549 (N_13549,N_13382,N_13467);
nand U13550 (N_13550,N_13122,N_13232);
xnor U13551 (N_13551,N_13082,N_13244);
and U13552 (N_13552,N_13332,N_13306);
nand U13553 (N_13553,N_13067,N_13177);
or U13554 (N_13554,N_13454,N_13013);
and U13555 (N_13555,N_13048,N_13345);
or U13556 (N_13556,N_13490,N_13436);
and U13557 (N_13557,N_13209,N_13483);
or U13558 (N_13558,N_13438,N_13238);
nor U13559 (N_13559,N_13287,N_13223);
nor U13560 (N_13560,N_13111,N_13251);
nand U13561 (N_13561,N_13062,N_13050);
xnor U13562 (N_13562,N_13250,N_13489);
xnor U13563 (N_13563,N_13146,N_13181);
nand U13564 (N_13564,N_13214,N_13124);
nand U13565 (N_13565,N_13064,N_13243);
or U13566 (N_13566,N_13189,N_13298);
and U13567 (N_13567,N_13356,N_13432);
and U13568 (N_13568,N_13117,N_13492);
nand U13569 (N_13569,N_13019,N_13427);
nand U13570 (N_13570,N_13261,N_13102);
or U13571 (N_13571,N_13015,N_13288);
or U13572 (N_13572,N_13284,N_13365);
nor U13573 (N_13573,N_13311,N_13392);
xor U13574 (N_13574,N_13475,N_13339);
and U13575 (N_13575,N_13393,N_13184);
nand U13576 (N_13576,N_13400,N_13113);
nor U13577 (N_13577,N_13242,N_13378);
nand U13578 (N_13578,N_13281,N_13377);
nand U13579 (N_13579,N_13070,N_13359);
or U13580 (N_13580,N_13491,N_13294);
nand U13581 (N_13581,N_13234,N_13154);
nand U13582 (N_13582,N_13423,N_13411);
nor U13583 (N_13583,N_13100,N_13430);
nand U13584 (N_13584,N_13086,N_13342);
xnor U13585 (N_13585,N_13253,N_13105);
and U13586 (N_13586,N_13343,N_13101);
or U13587 (N_13587,N_13196,N_13302);
nor U13588 (N_13588,N_13235,N_13039);
and U13589 (N_13589,N_13123,N_13457);
nor U13590 (N_13590,N_13014,N_13405);
nand U13591 (N_13591,N_13159,N_13179);
nor U13592 (N_13592,N_13128,N_13471);
nand U13593 (N_13593,N_13118,N_13499);
xor U13594 (N_13594,N_13229,N_13478);
nand U13595 (N_13595,N_13165,N_13194);
and U13596 (N_13596,N_13447,N_13420);
or U13597 (N_13597,N_13360,N_13069);
and U13598 (N_13598,N_13185,N_13369);
nor U13599 (N_13599,N_13166,N_13162);
xor U13600 (N_13600,N_13364,N_13027);
or U13601 (N_13601,N_13456,N_13136);
nand U13602 (N_13602,N_13174,N_13366);
and U13603 (N_13603,N_13439,N_13155);
or U13604 (N_13604,N_13325,N_13323);
xor U13605 (N_13605,N_13433,N_13421);
or U13606 (N_13606,N_13148,N_13271);
nor U13607 (N_13607,N_13443,N_13370);
nand U13608 (N_13608,N_13496,N_13012);
or U13609 (N_13609,N_13249,N_13285);
or U13610 (N_13610,N_13061,N_13029);
or U13611 (N_13611,N_13094,N_13297);
and U13612 (N_13612,N_13389,N_13380);
nand U13613 (N_13613,N_13350,N_13406);
nand U13614 (N_13614,N_13310,N_13001);
or U13615 (N_13615,N_13228,N_13337);
and U13616 (N_13616,N_13178,N_13092);
nand U13617 (N_13617,N_13246,N_13273);
and U13618 (N_13618,N_13161,N_13151);
nor U13619 (N_13619,N_13057,N_13225);
xnor U13620 (N_13620,N_13095,N_13133);
nor U13621 (N_13621,N_13462,N_13334);
nand U13622 (N_13622,N_13041,N_13099);
or U13623 (N_13623,N_13414,N_13036);
or U13624 (N_13624,N_13357,N_13056);
nand U13625 (N_13625,N_13180,N_13186);
and U13626 (N_13626,N_13084,N_13303);
nor U13627 (N_13627,N_13363,N_13286);
xnor U13628 (N_13628,N_13197,N_13268);
nor U13629 (N_13629,N_13387,N_13157);
nand U13630 (N_13630,N_13300,N_13453);
xor U13631 (N_13631,N_13016,N_13331);
nand U13632 (N_13632,N_13258,N_13063);
or U13633 (N_13633,N_13153,N_13301);
nor U13634 (N_13634,N_13396,N_13132);
nand U13635 (N_13635,N_13145,N_13291);
and U13636 (N_13636,N_13494,N_13130);
xnor U13637 (N_13637,N_13328,N_13465);
nor U13638 (N_13638,N_13442,N_13224);
nor U13639 (N_13639,N_13470,N_13341);
or U13640 (N_13640,N_13066,N_13333);
xor U13641 (N_13641,N_13353,N_13004);
and U13642 (N_13642,N_13207,N_13049);
xor U13643 (N_13643,N_13083,N_13448);
nor U13644 (N_13644,N_13296,N_13087);
and U13645 (N_13645,N_13452,N_13351);
and U13646 (N_13646,N_13114,N_13293);
xor U13647 (N_13647,N_13080,N_13203);
and U13648 (N_13648,N_13348,N_13472);
xnor U13649 (N_13649,N_13497,N_13417);
xnor U13650 (N_13650,N_13375,N_13263);
or U13651 (N_13651,N_13088,N_13429);
nand U13652 (N_13652,N_13042,N_13266);
or U13653 (N_13653,N_13199,N_13126);
xnor U13654 (N_13654,N_13307,N_13239);
or U13655 (N_13655,N_13010,N_13141);
nand U13656 (N_13656,N_13435,N_13327);
nand U13657 (N_13657,N_13474,N_13458);
or U13658 (N_13658,N_13320,N_13076);
nand U13659 (N_13659,N_13367,N_13259);
xnor U13660 (N_13660,N_13312,N_13060);
or U13661 (N_13661,N_13134,N_13322);
and U13662 (N_13662,N_13451,N_13397);
nor U13663 (N_13663,N_13262,N_13431);
nand U13664 (N_13664,N_13319,N_13371);
and U13665 (N_13665,N_13415,N_13493);
and U13666 (N_13666,N_13073,N_13485);
xor U13667 (N_13667,N_13103,N_13407);
xor U13668 (N_13668,N_13055,N_13487);
nand U13669 (N_13669,N_13227,N_13480);
and U13670 (N_13670,N_13028,N_13372);
nand U13671 (N_13671,N_13129,N_13202);
or U13672 (N_13672,N_13034,N_13163);
xnor U13673 (N_13673,N_13409,N_13085);
and U13674 (N_13674,N_13402,N_13461);
nand U13675 (N_13675,N_13222,N_13003);
nor U13676 (N_13676,N_13408,N_13187);
nor U13677 (N_13677,N_13473,N_13011);
nand U13678 (N_13678,N_13091,N_13215);
nor U13679 (N_13679,N_13354,N_13413);
nand U13680 (N_13680,N_13276,N_13098);
or U13681 (N_13681,N_13383,N_13292);
or U13682 (N_13682,N_13434,N_13217);
nor U13683 (N_13683,N_13403,N_13002);
and U13684 (N_13684,N_13024,N_13391);
nand U13685 (N_13685,N_13240,N_13231);
or U13686 (N_13686,N_13314,N_13139);
xor U13687 (N_13687,N_13017,N_13445);
or U13688 (N_13688,N_13289,N_13007);
nand U13689 (N_13689,N_13482,N_13468);
nand U13690 (N_13690,N_13347,N_13419);
and U13691 (N_13691,N_13426,N_13051);
xor U13692 (N_13692,N_13021,N_13441);
and U13693 (N_13693,N_13173,N_13410);
or U13694 (N_13694,N_13200,N_13388);
or U13695 (N_13695,N_13386,N_13152);
nor U13696 (N_13696,N_13290,N_13248);
nand U13697 (N_13697,N_13450,N_13190);
nor U13698 (N_13698,N_13008,N_13022);
or U13699 (N_13699,N_13270,N_13252);
or U13700 (N_13700,N_13104,N_13172);
xor U13701 (N_13701,N_13299,N_13035);
nor U13702 (N_13702,N_13205,N_13444);
or U13703 (N_13703,N_13150,N_13260);
xor U13704 (N_13704,N_13230,N_13278);
xor U13705 (N_13705,N_13361,N_13158);
or U13706 (N_13706,N_13280,N_13469);
nor U13707 (N_13707,N_13460,N_13038);
nor U13708 (N_13708,N_13484,N_13059);
nor U13709 (N_13709,N_13455,N_13264);
xor U13710 (N_13710,N_13198,N_13208);
nand U13711 (N_13711,N_13216,N_13398);
and U13712 (N_13712,N_13201,N_13428);
or U13713 (N_13713,N_13368,N_13054);
and U13714 (N_13714,N_13032,N_13226);
and U13715 (N_13715,N_13137,N_13120);
nand U13716 (N_13716,N_13309,N_13033);
nor U13717 (N_13717,N_13459,N_13183);
or U13718 (N_13718,N_13220,N_13424);
xor U13719 (N_13719,N_13476,N_13308);
xor U13720 (N_13720,N_13355,N_13127);
or U13721 (N_13721,N_13191,N_13047);
nand U13722 (N_13722,N_13358,N_13463);
xnor U13723 (N_13723,N_13108,N_13043);
nor U13724 (N_13724,N_13140,N_13160);
or U13725 (N_13725,N_13404,N_13486);
and U13726 (N_13726,N_13385,N_13009);
xnor U13727 (N_13727,N_13316,N_13045);
nor U13728 (N_13728,N_13346,N_13412);
or U13729 (N_13729,N_13170,N_13283);
nand U13730 (N_13730,N_13466,N_13313);
nor U13731 (N_13731,N_13381,N_13321);
or U13732 (N_13732,N_13395,N_13257);
or U13733 (N_13733,N_13040,N_13212);
xnor U13734 (N_13734,N_13481,N_13192);
xor U13735 (N_13735,N_13195,N_13204);
nor U13736 (N_13736,N_13349,N_13026);
xnor U13737 (N_13737,N_13075,N_13221);
or U13738 (N_13738,N_13147,N_13376);
xor U13739 (N_13739,N_13125,N_13275);
nand U13740 (N_13740,N_13416,N_13037);
xnor U13741 (N_13741,N_13175,N_13077);
nor U13742 (N_13742,N_13236,N_13089);
and U13743 (N_13743,N_13324,N_13488);
or U13744 (N_13744,N_13267,N_13373);
nor U13745 (N_13745,N_13495,N_13210);
and U13746 (N_13746,N_13020,N_13071);
and U13747 (N_13747,N_13106,N_13394);
nor U13748 (N_13748,N_13384,N_13052);
nor U13749 (N_13749,N_13329,N_13274);
nand U13750 (N_13750,N_13280,N_13384);
or U13751 (N_13751,N_13135,N_13499);
xnor U13752 (N_13752,N_13255,N_13327);
or U13753 (N_13753,N_13488,N_13379);
or U13754 (N_13754,N_13286,N_13339);
or U13755 (N_13755,N_13311,N_13376);
or U13756 (N_13756,N_13276,N_13380);
nor U13757 (N_13757,N_13475,N_13027);
and U13758 (N_13758,N_13156,N_13169);
nor U13759 (N_13759,N_13382,N_13040);
and U13760 (N_13760,N_13183,N_13399);
nand U13761 (N_13761,N_13416,N_13018);
nor U13762 (N_13762,N_13169,N_13036);
nand U13763 (N_13763,N_13175,N_13401);
xor U13764 (N_13764,N_13373,N_13039);
nand U13765 (N_13765,N_13279,N_13214);
xor U13766 (N_13766,N_13280,N_13114);
and U13767 (N_13767,N_13226,N_13437);
nand U13768 (N_13768,N_13342,N_13433);
nand U13769 (N_13769,N_13457,N_13286);
xor U13770 (N_13770,N_13105,N_13096);
xnor U13771 (N_13771,N_13060,N_13269);
nand U13772 (N_13772,N_13339,N_13429);
nor U13773 (N_13773,N_13399,N_13103);
xor U13774 (N_13774,N_13287,N_13334);
nor U13775 (N_13775,N_13332,N_13427);
or U13776 (N_13776,N_13094,N_13368);
and U13777 (N_13777,N_13168,N_13109);
or U13778 (N_13778,N_13286,N_13465);
nand U13779 (N_13779,N_13300,N_13012);
nor U13780 (N_13780,N_13326,N_13498);
and U13781 (N_13781,N_13439,N_13478);
or U13782 (N_13782,N_13131,N_13135);
nor U13783 (N_13783,N_13443,N_13377);
nand U13784 (N_13784,N_13249,N_13105);
nor U13785 (N_13785,N_13257,N_13425);
nand U13786 (N_13786,N_13176,N_13381);
or U13787 (N_13787,N_13185,N_13380);
or U13788 (N_13788,N_13247,N_13003);
nor U13789 (N_13789,N_13081,N_13472);
xor U13790 (N_13790,N_13125,N_13368);
nor U13791 (N_13791,N_13410,N_13332);
nand U13792 (N_13792,N_13009,N_13064);
nand U13793 (N_13793,N_13345,N_13396);
nor U13794 (N_13794,N_13434,N_13110);
and U13795 (N_13795,N_13327,N_13245);
nand U13796 (N_13796,N_13441,N_13191);
xor U13797 (N_13797,N_13092,N_13394);
and U13798 (N_13798,N_13171,N_13475);
nand U13799 (N_13799,N_13429,N_13099);
and U13800 (N_13800,N_13102,N_13450);
or U13801 (N_13801,N_13284,N_13239);
nand U13802 (N_13802,N_13373,N_13489);
and U13803 (N_13803,N_13269,N_13304);
nor U13804 (N_13804,N_13425,N_13193);
xnor U13805 (N_13805,N_13016,N_13294);
xnor U13806 (N_13806,N_13046,N_13453);
nand U13807 (N_13807,N_13483,N_13360);
or U13808 (N_13808,N_13033,N_13317);
and U13809 (N_13809,N_13249,N_13074);
nand U13810 (N_13810,N_13131,N_13234);
and U13811 (N_13811,N_13134,N_13419);
nand U13812 (N_13812,N_13224,N_13288);
and U13813 (N_13813,N_13052,N_13249);
and U13814 (N_13814,N_13454,N_13141);
xnor U13815 (N_13815,N_13103,N_13160);
xor U13816 (N_13816,N_13492,N_13438);
or U13817 (N_13817,N_13109,N_13106);
xor U13818 (N_13818,N_13234,N_13040);
and U13819 (N_13819,N_13322,N_13356);
and U13820 (N_13820,N_13060,N_13209);
and U13821 (N_13821,N_13316,N_13114);
nor U13822 (N_13822,N_13394,N_13439);
nor U13823 (N_13823,N_13269,N_13108);
xnor U13824 (N_13824,N_13024,N_13000);
nor U13825 (N_13825,N_13259,N_13042);
xnor U13826 (N_13826,N_13166,N_13036);
nand U13827 (N_13827,N_13489,N_13106);
or U13828 (N_13828,N_13225,N_13010);
xor U13829 (N_13829,N_13149,N_13234);
xnor U13830 (N_13830,N_13295,N_13461);
and U13831 (N_13831,N_13327,N_13198);
nand U13832 (N_13832,N_13467,N_13388);
and U13833 (N_13833,N_13249,N_13122);
nor U13834 (N_13834,N_13390,N_13297);
nand U13835 (N_13835,N_13414,N_13385);
or U13836 (N_13836,N_13336,N_13420);
nand U13837 (N_13837,N_13256,N_13190);
or U13838 (N_13838,N_13392,N_13330);
nor U13839 (N_13839,N_13332,N_13115);
or U13840 (N_13840,N_13384,N_13258);
and U13841 (N_13841,N_13178,N_13397);
xor U13842 (N_13842,N_13431,N_13200);
nand U13843 (N_13843,N_13069,N_13175);
or U13844 (N_13844,N_13033,N_13140);
nand U13845 (N_13845,N_13255,N_13425);
nor U13846 (N_13846,N_13055,N_13337);
and U13847 (N_13847,N_13006,N_13272);
and U13848 (N_13848,N_13094,N_13065);
and U13849 (N_13849,N_13158,N_13047);
xor U13850 (N_13850,N_13032,N_13223);
nor U13851 (N_13851,N_13203,N_13145);
nand U13852 (N_13852,N_13169,N_13460);
nor U13853 (N_13853,N_13060,N_13364);
or U13854 (N_13854,N_13116,N_13031);
nand U13855 (N_13855,N_13091,N_13418);
and U13856 (N_13856,N_13329,N_13418);
xor U13857 (N_13857,N_13154,N_13045);
xor U13858 (N_13858,N_13100,N_13366);
xor U13859 (N_13859,N_13302,N_13429);
or U13860 (N_13860,N_13174,N_13051);
nor U13861 (N_13861,N_13240,N_13235);
or U13862 (N_13862,N_13359,N_13481);
xnor U13863 (N_13863,N_13163,N_13369);
or U13864 (N_13864,N_13006,N_13339);
nand U13865 (N_13865,N_13278,N_13025);
xnor U13866 (N_13866,N_13306,N_13135);
or U13867 (N_13867,N_13319,N_13307);
xor U13868 (N_13868,N_13366,N_13235);
and U13869 (N_13869,N_13423,N_13349);
xnor U13870 (N_13870,N_13435,N_13152);
and U13871 (N_13871,N_13021,N_13028);
and U13872 (N_13872,N_13495,N_13064);
and U13873 (N_13873,N_13011,N_13320);
nor U13874 (N_13874,N_13062,N_13093);
nand U13875 (N_13875,N_13380,N_13441);
nand U13876 (N_13876,N_13276,N_13390);
and U13877 (N_13877,N_13112,N_13424);
or U13878 (N_13878,N_13411,N_13342);
nor U13879 (N_13879,N_13253,N_13309);
or U13880 (N_13880,N_13139,N_13389);
or U13881 (N_13881,N_13278,N_13308);
nor U13882 (N_13882,N_13214,N_13267);
nand U13883 (N_13883,N_13072,N_13258);
nand U13884 (N_13884,N_13216,N_13307);
nand U13885 (N_13885,N_13130,N_13266);
xnor U13886 (N_13886,N_13396,N_13281);
xor U13887 (N_13887,N_13400,N_13027);
xor U13888 (N_13888,N_13283,N_13211);
xor U13889 (N_13889,N_13480,N_13020);
xor U13890 (N_13890,N_13111,N_13229);
and U13891 (N_13891,N_13154,N_13016);
xnor U13892 (N_13892,N_13262,N_13209);
xor U13893 (N_13893,N_13086,N_13166);
nand U13894 (N_13894,N_13033,N_13310);
nor U13895 (N_13895,N_13289,N_13218);
xor U13896 (N_13896,N_13319,N_13398);
xor U13897 (N_13897,N_13403,N_13214);
or U13898 (N_13898,N_13240,N_13015);
nand U13899 (N_13899,N_13429,N_13083);
xor U13900 (N_13900,N_13452,N_13480);
or U13901 (N_13901,N_13403,N_13045);
nor U13902 (N_13902,N_13476,N_13232);
nand U13903 (N_13903,N_13292,N_13072);
or U13904 (N_13904,N_13419,N_13021);
nand U13905 (N_13905,N_13250,N_13449);
nor U13906 (N_13906,N_13479,N_13045);
or U13907 (N_13907,N_13452,N_13137);
xor U13908 (N_13908,N_13461,N_13246);
xnor U13909 (N_13909,N_13166,N_13290);
and U13910 (N_13910,N_13001,N_13268);
and U13911 (N_13911,N_13158,N_13045);
or U13912 (N_13912,N_13006,N_13398);
nor U13913 (N_13913,N_13123,N_13118);
or U13914 (N_13914,N_13099,N_13322);
nor U13915 (N_13915,N_13321,N_13468);
or U13916 (N_13916,N_13430,N_13125);
and U13917 (N_13917,N_13495,N_13300);
nand U13918 (N_13918,N_13104,N_13267);
or U13919 (N_13919,N_13356,N_13018);
nor U13920 (N_13920,N_13366,N_13314);
nor U13921 (N_13921,N_13152,N_13061);
nor U13922 (N_13922,N_13002,N_13004);
nand U13923 (N_13923,N_13166,N_13307);
xnor U13924 (N_13924,N_13343,N_13078);
nand U13925 (N_13925,N_13447,N_13146);
and U13926 (N_13926,N_13085,N_13069);
nand U13927 (N_13927,N_13258,N_13250);
or U13928 (N_13928,N_13229,N_13126);
nor U13929 (N_13929,N_13357,N_13060);
nor U13930 (N_13930,N_13365,N_13342);
and U13931 (N_13931,N_13292,N_13224);
xnor U13932 (N_13932,N_13320,N_13242);
xor U13933 (N_13933,N_13262,N_13375);
nor U13934 (N_13934,N_13168,N_13275);
or U13935 (N_13935,N_13214,N_13009);
and U13936 (N_13936,N_13253,N_13175);
nor U13937 (N_13937,N_13057,N_13180);
or U13938 (N_13938,N_13060,N_13224);
nand U13939 (N_13939,N_13300,N_13175);
and U13940 (N_13940,N_13214,N_13252);
and U13941 (N_13941,N_13078,N_13210);
and U13942 (N_13942,N_13178,N_13325);
nand U13943 (N_13943,N_13112,N_13190);
nor U13944 (N_13944,N_13061,N_13435);
nand U13945 (N_13945,N_13308,N_13228);
or U13946 (N_13946,N_13285,N_13299);
nor U13947 (N_13947,N_13346,N_13004);
nand U13948 (N_13948,N_13275,N_13454);
and U13949 (N_13949,N_13000,N_13408);
and U13950 (N_13950,N_13221,N_13260);
xnor U13951 (N_13951,N_13044,N_13331);
nand U13952 (N_13952,N_13213,N_13493);
or U13953 (N_13953,N_13135,N_13453);
and U13954 (N_13954,N_13177,N_13396);
or U13955 (N_13955,N_13181,N_13259);
and U13956 (N_13956,N_13005,N_13044);
nor U13957 (N_13957,N_13040,N_13455);
nor U13958 (N_13958,N_13050,N_13225);
or U13959 (N_13959,N_13055,N_13140);
nor U13960 (N_13960,N_13349,N_13048);
nand U13961 (N_13961,N_13297,N_13256);
nor U13962 (N_13962,N_13054,N_13159);
and U13963 (N_13963,N_13113,N_13320);
nor U13964 (N_13964,N_13285,N_13138);
and U13965 (N_13965,N_13201,N_13182);
nand U13966 (N_13966,N_13187,N_13051);
and U13967 (N_13967,N_13034,N_13321);
nor U13968 (N_13968,N_13176,N_13060);
nand U13969 (N_13969,N_13455,N_13093);
xnor U13970 (N_13970,N_13133,N_13489);
nor U13971 (N_13971,N_13203,N_13290);
xor U13972 (N_13972,N_13352,N_13158);
or U13973 (N_13973,N_13474,N_13197);
xnor U13974 (N_13974,N_13177,N_13226);
or U13975 (N_13975,N_13275,N_13312);
nor U13976 (N_13976,N_13295,N_13187);
nor U13977 (N_13977,N_13232,N_13303);
nand U13978 (N_13978,N_13454,N_13407);
nand U13979 (N_13979,N_13396,N_13048);
and U13980 (N_13980,N_13216,N_13188);
or U13981 (N_13981,N_13010,N_13471);
and U13982 (N_13982,N_13139,N_13452);
and U13983 (N_13983,N_13321,N_13482);
xor U13984 (N_13984,N_13409,N_13249);
and U13985 (N_13985,N_13050,N_13394);
and U13986 (N_13986,N_13249,N_13269);
or U13987 (N_13987,N_13068,N_13271);
xnor U13988 (N_13988,N_13191,N_13083);
nor U13989 (N_13989,N_13177,N_13208);
nand U13990 (N_13990,N_13457,N_13176);
and U13991 (N_13991,N_13068,N_13146);
or U13992 (N_13992,N_13068,N_13057);
or U13993 (N_13993,N_13381,N_13110);
or U13994 (N_13994,N_13153,N_13445);
nand U13995 (N_13995,N_13359,N_13038);
nand U13996 (N_13996,N_13073,N_13288);
or U13997 (N_13997,N_13411,N_13435);
or U13998 (N_13998,N_13222,N_13474);
nand U13999 (N_13999,N_13371,N_13206);
and U14000 (N_14000,N_13749,N_13663);
xor U14001 (N_14001,N_13610,N_13502);
nor U14002 (N_14002,N_13710,N_13875);
nor U14003 (N_14003,N_13566,N_13611);
and U14004 (N_14004,N_13720,N_13982);
nor U14005 (N_14005,N_13598,N_13865);
or U14006 (N_14006,N_13960,N_13683);
nand U14007 (N_14007,N_13902,N_13519);
and U14008 (N_14008,N_13792,N_13848);
nor U14009 (N_14009,N_13837,N_13796);
nand U14010 (N_14010,N_13782,N_13584);
xnor U14011 (N_14011,N_13641,N_13593);
or U14012 (N_14012,N_13942,N_13880);
nor U14013 (N_14013,N_13995,N_13677);
nand U14014 (N_14014,N_13536,N_13866);
nand U14015 (N_14015,N_13565,N_13992);
nor U14016 (N_14016,N_13829,N_13976);
and U14017 (N_14017,N_13769,N_13779);
nor U14018 (N_14018,N_13851,N_13887);
nand U14019 (N_14019,N_13546,N_13578);
nand U14020 (N_14020,N_13687,N_13522);
nand U14021 (N_14021,N_13905,N_13797);
and U14022 (N_14022,N_13874,N_13891);
or U14023 (N_14023,N_13669,N_13956);
and U14024 (N_14024,N_13650,N_13871);
or U14025 (N_14025,N_13527,N_13670);
and U14026 (N_14026,N_13915,N_13886);
nor U14027 (N_14027,N_13740,N_13711);
or U14028 (N_14028,N_13959,N_13858);
and U14029 (N_14029,N_13607,N_13946);
or U14030 (N_14030,N_13606,N_13854);
nand U14031 (N_14031,N_13764,N_13523);
or U14032 (N_14032,N_13906,N_13879);
nor U14033 (N_14033,N_13569,N_13570);
or U14034 (N_14034,N_13872,N_13647);
or U14035 (N_14035,N_13716,N_13990);
and U14036 (N_14036,N_13654,N_13852);
and U14037 (N_14037,N_13741,N_13581);
or U14038 (N_14038,N_13948,N_13582);
and U14039 (N_14039,N_13660,N_13961);
nand U14040 (N_14040,N_13985,N_13927);
and U14041 (N_14041,N_13576,N_13747);
or U14042 (N_14042,N_13763,N_13672);
nor U14043 (N_14043,N_13511,N_13613);
nor U14044 (N_14044,N_13640,N_13739);
nand U14045 (N_14045,N_13555,N_13688);
and U14046 (N_14046,N_13929,N_13678);
nand U14047 (N_14047,N_13540,N_13724);
or U14048 (N_14048,N_13781,N_13734);
and U14049 (N_14049,N_13510,N_13790);
xor U14050 (N_14050,N_13708,N_13923);
nor U14051 (N_14051,N_13701,N_13723);
or U14052 (N_14052,N_13587,N_13869);
xnor U14053 (N_14053,N_13704,N_13623);
and U14054 (N_14054,N_13624,N_13549);
nor U14055 (N_14055,N_13890,N_13776);
nor U14056 (N_14056,N_13639,N_13896);
nand U14057 (N_14057,N_13726,N_13812);
xor U14058 (N_14058,N_13912,N_13689);
nand U14059 (N_14059,N_13501,N_13673);
nor U14060 (N_14060,N_13864,N_13533);
nand U14061 (N_14061,N_13873,N_13955);
nand U14062 (N_14062,N_13938,N_13809);
or U14063 (N_14063,N_13843,N_13856);
nor U14064 (N_14064,N_13970,N_13737);
nor U14065 (N_14065,N_13941,N_13520);
xnor U14066 (N_14066,N_13818,N_13589);
and U14067 (N_14067,N_13652,N_13560);
nand U14068 (N_14068,N_13867,N_13712);
xor U14069 (N_14069,N_13577,N_13996);
nor U14070 (N_14070,N_13631,N_13666);
or U14071 (N_14071,N_13922,N_13535);
and U14072 (N_14072,N_13838,N_13831);
or U14073 (N_14073,N_13991,N_13870);
and U14074 (N_14074,N_13596,N_13529);
or U14075 (N_14075,N_13811,N_13725);
and U14076 (N_14076,N_13903,N_13998);
xor U14077 (N_14077,N_13789,N_13988);
nor U14078 (N_14078,N_13630,N_13760);
and U14079 (N_14079,N_13735,N_13757);
and U14080 (N_14080,N_13943,N_13628);
nor U14081 (N_14081,N_13595,N_13550);
or U14082 (N_14082,N_13893,N_13950);
and U14083 (N_14083,N_13933,N_13963);
xor U14084 (N_14084,N_13750,N_13958);
xor U14085 (N_14085,N_13951,N_13778);
or U14086 (N_14086,N_13616,N_13795);
nor U14087 (N_14087,N_13826,N_13813);
nor U14088 (N_14088,N_13823,N_13810);
or U14089 (N_14089,N_13846,N_13655);
or U14090 (N_14090,N_13692,N_13521);
nand U14091 (N_14091,N_13594,N_13700);
nor U14092 (N_14092,N_13817,N_13690);
xnor U14093 (N_14093,N_13936,N_13766);
or U14094 (N_14094,N_13626,N_13884);
nor U14095 (N_14095,N_13787,N_13999);
nor U14096 (N_14096,N_13706,N_13572);
xor U14097 (N_14097,N_13755,N_13833);
and U14098 (N_14098,N_13820,N_13987);
nand U14099 (N_14099,N_13842,N_13804);
and U14100 (N_14100,N_13892,N_13602);
or U14101 (N_14101,N_13707,N_13586);
nand U14102 (N_14102,N_13953,N_13807);
nor U14103 (N_14103,N_13965,N_13733);
nand U14104 (N_14104,N_13850,N_13849);
or U14105 (N_14105,N_13952,N_13913);
nor U14106 (N_14106,N_13591,N_13808);
xnor U14107 (N_14107,N_13767,N_13939);
nand U14108 (N_14108,N_13994,N_13619);
or U14109 (N_14109,N_13580,N_13785);
nand U14110 (N_14110,N_13573,N_13847);
nor U14111 (N_14111,N_13911,N_13964);
xor U14112 (N_14112,N_13899,N_13705);
and U14113 (N_14113,N_13685,N_13840);
or U14114 (N_14114,N_13667,N_13986);
xor U14115 (N_14115,N_13901,N_13857);
and U14116 (N_14116,N_13661,N_13585);
or U14117 (N_14117,N_13878,N_13682);
xor U14118 (N_14118,N_13625,N_13815);
or U14119 (N_14119,N_13974,N_13590);
nand U14120 (N_14120,N_13830,N_13894);
nor U14121 (N_14121,N_13799,N_13968);
and U14122 (N_14122,N_13621,N_13681);
nor U14123 (N_14123,N_13756,N_13679);
nor U14124 (N_14124,N_13579,N_13861);
and U14125 (N_14125,N_13548,N_13889);
or U14126 (N_14126,N_13786,N_13822);
and U14127 (N_14127,N_13571,N_13676);
and U14128 (N_14128,N_13897,N_13643);
xor U14129 (N_14129,N_13759,N_13806);
and U14130 (N_14130,N_13742,N_13505);
nor U14131 (N_14131,N_13798,N_13814);
or U14132 (N_14132,N_13526,N_13604);
nand U14133 (N_14133,N_13754,N_13937);
and U14134 (N_14134,N_13907,N_13714);
nand U14135 (N_14135,N_13920,N_13694);
xor U14136 (N_14136,N_13805,N_13668);
nor U14137 (N_14137,N_13841,N_13718);
nor U14138 (N_14138,N_13541,N_13553);
and U14139 (N_14139,N_13559,N_13558);
xor U14140 (N_14140,N_13877,N_13618);
xnor U14141 (N_14141,N_13715,N_13644);
or U14142 (N_14142,N_13802,N_13824);
nand U14143 (N_14143,N_13772,N_13717);
nand U14144 (N_14144,N_13561,N_13695);
or U14145 (N_14145,N_13574,N_13512);
xor U14146 (N_14146,N_13888,N_13562);
nor U14147 (N_14147,N_13917,N_13752);
xor U14148 (N_14148,N_13753,N_13973);
nand U14149 (N_14149,N_13699,N_13909);
and U14150 (N_14150,N_13931,N_13684);
xor U14151 (N_14151,N_13924,N_13600);
or U14152 (N_14152,N_13642,N_13605);
and U14153 (N_14153,N_13957,N_13632);
or U14154 (N_14154,N_13979,N_13853);
xor U14155 (N_14155,N_13925,N_13828);
xnor U14156 (N_14156,N_13504,N_13722);
or U14157 (N_14157,N_13819,N_13801);
xor U14158 (N_14158,N_13691,N_13984);
nand U14159 (N_14159,N_13980,N_13534);
xnor U14160 (N_14160,N_13516,N_13544);
nor U14161 (N_14161,N_13966,N_13608);
nand U14162 (N_14162,N_13895,N_13665);
or U14163 (N_14163,N_13969,N_13629);
and U14164 (N_14164,N_13738,N_13839);
and U14165 (N_14165,N_13971,N_13881);
or U14166 (N_14166,N_13904,N_13545);
and U14167 (N_14167,N_13693,N_13524);
or U14168 (N_14168,N_13648,N_13784);
xnor U14169 (N_14169,N_13774,N_13612);
nor U14170 (N_14170,N_13713,N_13653);
and U14171 (N_14171,N_13832,N_13638);
xnor U14172 (N_14172,N_13836,N_13821);
and U14173 (N_14173,N_13928,N_13816);
xor U14174 (N_14174,N_13926,N_13563);
xnor U14175 (N_14175,N_13721,N_13531);
xor U14176 (N_14176,N_13883,N_13634);
and U14177 (N_14177,N_13636,N_13539);
and U14178 (N_14178,N_13993,N_13696);
nand U14179 (N_14179,N_13674,N_13736);
and U14180 (N_14180,N_13697,N_13916);
nor U14181 (N_14181,N_13765,N_13791);
or U14182 (N_14182,N_13910,N_13675);
nand U14183 (N_14183,N_13564,N_13934);
or U14184 (N_14184,N_13954,N_13921);
or U14185 (N_14185,N_13868,N_13967);
and U14186 (N_14186,N_13962,N_13863);
xnor U14187 (N_14187,N_13758,N_13517);
and U14188 (N_14188,N_13592,N_13635);
xnor U14189 (N_14189,N_13882,N_13500);
and U14190 (N_14190,N_13780,N_13658);
nor U14191 (N_14191,N_13949,N_13744);
xor U14192 (N_14192,N_13554,N_13919);
nand U14193 (N_14193,N_13745,N_13876);
nor U14194 (N_14194,N_13898,N_13659);
xor U14195 (N_14195,N_13583,N_13859);
nand U14196 (N_14196,N_13528,N_13514);
and U14197 (N_14197,N_13935,N_13783);
or U14198 (N_14198,N_13537,N_13513);
xnor U14199 (N_14199,N_13645,N_13637);
or U14200 (N_14200,N_13729,N_13551);
nor U14201 (N_14201,N_13947,N_13657);
nand U14202 (N_14202,N_13761,N_13633);
nor U14203 (N_14203,N_13530,N_13944);
or U14204 (N_14204,N_13686,N_13506);
or U14205 (N_14205,N_13768,N_13855);
nor U14206 (N_14206,N_13793,N_13732);
nor U14207 (N_14207,N_13975,N_13508);
or U14208 (N_14208,N_13844,N_13918);
nand U14209 (N_14209,N_13972,N_13800);
and U14210 (N_14210,N_13671,N_13542);
and U14211 (N_14211,N_13538,N_13543);
xnor U14212 (N_14212,N_13599,N_13885);
and U14213 (N_14213,N_13827,N_13835);
nand U14214 (N_14214,N_13620,N_13664);
nor U14215 (N_14215,N_13656,N_13547);
xnor U14216 (N_14216,N_13575,N_13770);
xnor U14217 (N_14217,N_13940,N_13603);
nor U14218 (N_14218,N_13983,N_13860);
nor U14219 (N_14219,N_13557,N_13908);
nand U14220 (N_14220,N_13773,N_13702);
xor U14221 (N_14221,N_13509,N_13622);
and U14222 (N_14222,N_13862,N_13703);
xnor U14223 (N_14223,N_13981,N_13709);
or U14224 (N_14224,N_13649,N_13803);
and U14225 (N_14225,N_13627,N_13794);
nand U14226 (N_14226,N_13568,N_13771);
or U14227 (N_14227,N_13532,N_13617);
nor U14228 (N_14228,N_13507,N_13615);
nor U14229 (N_14229,N_13978,N_13748);
xnor U14230 (N_14230,N_13567,N_13698);
nand U14231 (N_14231,N_13914,N_13515);
or U14232 (N_14232,N_13997,N_13762);
or U14233 (N_14233,N_13588,N_13662);
or U14234 (N_14234,N_13719,N_13751);
nor U14235 (N_14235,N_13614,N_13556);
nand U14236 (N_14236,N_13777,N_13834);
nand U14237 (N_14237,N_13932,N_13597);
and U14238 (N_14238,N_13728,N_13731);
nand U14239 (N_14239,N_13727,N_13525);
nand U14240 (N_14240,N_13730,N_13945);
or U14241 (N_14241,N_13503,N_13651);
xnor U14242 (N_14242,N_13646,N_13989);
and U14243 (N_14243,N_13977,N_13609);
and U14244 (N_14244,N_13900,N_13825);
xnor U14245 (N_14245,N_13552,N_13788);
and U14246 (N_14246,N_13601,N_13845);
nor U14247 (N_14247,N_13746,N_13775);
xor U14248 (N_14248,N_13518,N_13743);
and U14249 (N_14249,N_13680,N_13930);
nor U14250 (N_14250,N_13744,N_13988);
nor U14251 (N_14251,N_13910,N_13658);
or U14252 (N_14252,N_13706,N_13756);
xnor U14253 (N_14253,N_13834,N_13995);
or U14254 (N_14254,N_13898,N_13998);
or U14255 (N_14255,N_13717,N_13698);
and U14256 (N_14256,N_13676,N_13912);
xnor U14257 (N_14257,N_13722,N_13796);
xor U14258 (N_14258,N_13640,N_13805);
and U14259 (N_14259,N_13730,N_13757);
and U14260 (N_14260,N_13527,N_13933);
xnor U14261 (N_14261,N_13882,N_13700);
nor U14262 (N_14262,N_13700,N_13942);
or U14263 (N_14263,N_13936,N_13852);
xnor U14264 (N_14264,N_13583,N_13997);
nand U14265 (N_14265,N_13843,N_13942);
nand U14266 (N_14266,N_13876,N_13674);
nand U14267 (N_14267,N_13573,N_13596);
nand U14268 (N_14268,N_13999,N_13639);
nand U14269 (N_14269,N_13718,N_13518);
nor U14270 (N_14270,N_13843,N_13703);
and U14271 (N_14271,N_13523,N_13855);
or U14272 (N_14272,N_13590,N_13841);
nand U14273 (N_14273,N_13811,N_13844);
nand U14274 (N_14274,N_13788,N_13656);
nor U14275 (N_14275,N_13533,N_13876);
xnor U14276 (N_14276,N_13987,N_13648);
nand U14277 (N_14277,N_13685,N_13788);
and U14278 (N_14278,N_13824,N_13614);
xor U14279 (N_14279,N_13774,N_13600);
xnor U14280 (N_14280,N_13589,N_13993);
xor U14281 (N_14281,N_13569,N_13711);
or U14282 (N_14282,N_13982,N_13912);
xnor U14283 (N_14283,N_13838,N_13500);
nand U14284 (N_14284,N_13947,N_13524);
nand U14285 (N_14285,N_13951,N_13733);
nor U14286 (N_14286,N_13758,N_13969);
nor U14287 (N_14287,N_13875,N_13989);
or U14288 (N_14288,N_13655,N_13967);
and U14289 (N_14289,N_13741,N_13870);
or U14290 (N_14290,N_13922,N_13860);
xnor U14291 (N_14291,N_13972,N_13979);
nand U14292 (N_14292,N_13987,N_13733);
or U14293 (N_14293,N_13929,N_13731);
or U14294 (N_14294,N_13583,N_13732);
xor U14295 (N_14295,N_13637,N_13509);
or U14296 (N_14296,N_13614,N_13665);
nand U14297 (N_14297,N_13756,N_13536);
nand U14298 (N_14298,N_13572,N_13573);
or U14299 (N_14299,N_13749,N_13712);
or U14300 (N_14300,N_13514,N_13722);
and U14301 (N_14301,N_13804,N_13706);
xnor U14302 (N_14302,N_13719,N_13930);
and U14303 (N_14303,N_13750,N_13850);
nand U14304 (N_14304,N_13988,N_13855);
nor U14305 (N_14305,N_13518,N_13568);
nor U14306 (N_14306,N_13570,N_13572);
and U14307 (N_14307,N_13918,N_13792);
or U14308 (N_14308,N_13671,N_13615);
xor U14309 (N_14309,N_13867,N_13975);
nand U14310 (N_14310,N_13884,N_13588);
or U14311 (N_14311,N_13614,N_13704);
nand U14312 (N_14312,N_13769,N_13688);
xor U14313 (N_14313,N_13686,N_13519);
and U14314 (N_14314,N_13676,N_13981);
nand U14315 (N_14315,N_13560,N_13943);
and U14316 (N_14316,N_13803,N_13860);
and U14317 (N_14317,N_13772,N_13771);
and U14318 (N_14318,N_13869,N_13591);
nand U14319 (N_14319,N_13627,N_13609);
xor U14320 (N_14320,N_13842,N_13595);
nand U14321 (N_14321,N_13939,N_13879);
xor U14322 (N_14322,N_13977,N_13774);
or U14323 (N_14323,N_13938,N_13579);
nor U14324 (N_14324,N_13661,N_13987);
or U14325 (N_14325,N_13842,N_13502);
and U14326 (N_14326,N_13807,N_13909);
xnor U14327 (N_14327,N_13703,N_13920);
nand U14328 (N_14328,N_13780,N_13874);
xor U14329 (N_14329,N_13678,N_13596);
nand U14330 (N_14330,N_13962,N_13570);
and U14331 (N_14331,N_13635,N_13901);
and U14332 (N_14332,N_13787,N_13520);
or U14333 (N_14333,N_13868,N_13618);
and U14334 (N_14334,N_13593,N_13825);
nand U14335 (N_14335,N_13654,N_13972);
nor U14336 (N_14336,N_13618,N_13828);
or U14337 (N_14337,N_13921,N_13869);
and U14338 (N_14338,N_13991,N_13706);
and U14339 (N_14339,N_13930,N_13974);
nor U14340 (N_14340,N_13577,N_13960);
and U14341 (N_14341,N_13748,N_13803);
and U14342 (N_14342,N_13649,N_13870);
or U14343 (N_14343,N_13690,N_13806);
nand U14344 (N_14344,N_13989,N_13876);
nor U14345 (N_14345,N_13999,N_13527);
and U14346 (N_14346,N_13766,N_13974);
and U14347 (N_14347,N_13884,N_13557);
and U14348 (N_14348,N_13892,N_13521);
and U14349 (N_14349,N_13511,N_13996);
or U14350 (N_14350,N_13553,N_13799);
and U14351 (N_14351,N_13666,N_13949);
nand U14352 (N_14352,N_13756,N_13861);
and U14353 (N_14353,N_13571,N_13707);
nor U14354 (N_14354,N_13547,N_13677);
nor U14355 (N_14355,N_13987,N_13582);
xor U14356 (N_14356,N_13912,N_13940);
and U14357 (N_14357,N_13886,N_13630);
or U14358 (N_14358,N_13561,N_13909);
or U14359 (N_14359,N_13983,N_13990);
or U14360 (N_14360,N_13834,N_13778);
nand U14361 (N_14361,N_13929,N_13649);
or U14362 (N_14362,N_13853,N_13913);
and U14363 (N_14363,N_13747,N_13816);
nor U14364 (N_14364,N_13856,N_13845);
nor U14365 (N_14365,N_13784,N_13716);
and U14366 (N_14366,N_13884,N_13875);
nor U14367 (N_14367,N_13644,N_13660);
nand U14368 (N_14368,N_13944,N_13577);
or U14369 (N_14369,N_13620,N_13641);
nor U14370 (N_14370,N_13548,N_13524);
nand U14371 (N_14371,N_13658,N_13668);
nand U14372 (N_14372,N_13846,N_13773);
xor U14373 (N_14373,N_13620,N_13701);
nor U14374 (N_14374,N_13746,N_13818);
or U14375 (N_14375,N_13870,N_13778);
and U14376 (N_14376,N_13678,N_13904);
and U14377 (N_14377,N_13613,N_13896);
xnor U14378 (N_14378,N_13686,N_13753);
nor U14379 (N_14379,N_13703,N_13994);
or U14380 (N_14380,N_13853,N_13505);
xnor U14381 (N_14381,N_13870,N_13701);
xnor U14382 (N_14382,N_13809,N_13977);
and U14383 (N_14383,N_13548,N_13619);
xnor U14384 (N_14384,N_13782,N_13784);
or U14385 (N_14385,N_13643,N_13688);
and U14386 (N_14386,N_13950,N_13978);
nand U14387 (N_14387,N_13512,N_13853);
nand U14388 (N_14388,N_13912,N_13640);
xnor U14389 (N_14389,N_13874,N_13990);
xor U14390 (N_14390,N_13960,N_13534);
nand U14391 (N_14391,N_13716,N_13891);
nor U14392 (N_14392,N_13827,N_13754);
and U14393 (N_14393,N_13948,N_13545);
nand U14394 (N_14394,N_13718,N_13950);
xor U14395 (N_14395,N_13791,N_13786);
nor U14396 (N_14396,N_13933,N_13721);
nand U14397 (N_14397,N_13580,N_13642);
or U14398 (N_14398,N_13991,N_13609);
or U14399 (N_14399,N_13856,N_13919);
or U14400 (N_14400,N_13505,N_13966);
xor U14401 (N_14401,N_13560,N_13592);
and U14402 (N_14402,N_13545,N_13539);
nand U14403 (N_14403,N_13832,N_13839);
and U14404 (N_14404,N_13966,N_13650);
xor U14405 (N_14405,N_13843,N_13976);
nand U14406 (N_14406,N_13602,N_13905);
nand U14407 (N_14407,N_13668,N_13663);
or U14408 (N_14408,N_13518,N_13609);
and U14409 (N_14409,N_13941,N_13623);
xnor U14410 (N_14410,N_13790,N_13859);
nor U14411 (N_14411,N_13875,N_13728);
xor U14412 (N_14412,N_13552,N_13637);
nand U14413 (N_14413,N_13877,N_13903);
nor U14414 (N_14414,N_13709,N_13836);
or U14415 (N_14415,N_13676,N_13945);
and U14416 (N_14416,N_13518,N_13789);
nor U14417 (N_14417,N_13774,N_13723);
nand U14418 (N_14418,N_13929,N_13564);
nor U14419 (N_14419,N_13727,N_13641);
nand U14420 (N_14420,N_13627,N_13576);
nor U14421 (N_14421,N_13536,N_13694);
nand U14422 (N_14422,N_13879,N_13837);
xnor U14423 (N_14423,N_13969,N_13671);
and U14424 (N_14424,N_13927,N_13874);
xor U14425 (N_14425,N_13735,N_13798);
nor U14426 (N_14426,N_13638,N_13708);
and U14427 (N_14427,N_13896,N_13773);
nor U14428 (N_14428,N_13603,N_13675);
xor U14429 (N_14429,N_13568,N_13950);
nand U14430 (N_14430,N_13667,N_13812);
and U14431 (N_14431,N_13950,N_13884);
or U14432 (N_14432,N_13628,N_13546);
or U14433 (N_14433,N_13918,N_13984);
nand U14434 (N_14434,N_13855,N_13985);
nand U14435 (N_14435,N_13701,N_13518);
xor U14436 (N_14436,N_13943,N_13918);
and U14437 (N_14437,N_13760,N_13775);
xnor U14438 (N_14438,N_13785,N_13817);
nand U14439 (N_14439,N_13888,N_13993);
nor U14440 (N_14440,N_13630,N_13876);
nor U14441 (N_14441,N_13699,N_13780);
and U14442 (N_14442,N_13535,N_13915);
nor U14443 (N_14443,N_13923,N_13669);
nor U14444 (N_14444,N_13900,N_13537);
and U14445 (N_14445,N_13518,N_13699);
nand U14446 (N_14446,N_13864,N_13876);
or U14447 (N_14447,N_13834,N_13673);
xor U14448 (N_14448,N_13731,N_13755);
xnor U14449 (N_14449,N_13540,N_13906);
nor U14450 (N_14450,N_13891,N_13617);
or U14451 (N_14451,N_13822,N_13769);
or U14452 (N_14452,N_13726,N_13958);
and U14453 (N_14453,N_13741,N_13558);
xnor U14454 (N_14454,N_13825,N_13623);
nor U14455 (N_14455,N_13923,N_13648);
nor U14456 (N_14456,N_13942,N_13575);
nor U14457 (N_14457,N_13711,N_13816);
xor U14458 (N_14458,N_13753,N_13724);
and U14459 (N_14459,N_13983,N_13749);
nor U14460 (N_14460,N_13679,N_13599);
nand U14461 (N_14461,N_13725,N_13641);
xor U14462 (N_14462,N_13626,N_13792);
nor U14463 (N_14463,N_13776,N_13935);
and U14464 (N_14464,N_13833,N_13928);
or U14465 (N_14465,N_13979,N_13941);
or U14466 (N_14466,N_13622,N_13816);
and U14467 (N_14467,N_13822,N_13644);
and U14468 (N_14468,N_13624,N_13719);
nand U14469 (N_14469,N_13846,N_13646);
xor U14470 (N_14470,N_13734,N_13729);
or U14471 (N_14471,N_13667,N_13849);
xnor U14472 (N_14472,N_13614,N_13974);
nand U14473 (N_14473,N_13687,N_13580);
nand U14474 (N_14474,N_13850,N_13878);
nand U14475 (N_14475,N_13964,N_13521);
xor U14476 (N_14476,N_13561,N_13963);
nand U14477 (N_14477,N_13811,N_13776);
xnor U14478 (N_14478,N_13976,N_13634);
nand U14479 (N_14479,N_13916,N_13905);
nor U14480 (N_14480,N_13922,N_13950);
xor U14481 (N_14481,N_13855,N_13861);
nand U14482 (N_14482,N_13538,N_13508);
and U14483 (N_14483,N_13745,N_13936);
nand U14484 (N_14484,N_13976,N_13673);
nand U14485 (N_14485,N_13927,N_13937);
or U14486 (N_14486,N_13803,N_13623);
nand U14487 (N_14487,N_13684,N_13563);
nand U14488 (N_14488,N_13504,N_13927);
and U14489 (N_14489,N_13616,N_13560);
or U14490 (N_14490,N_13593,N_13983);
or U14491 (N_14491,N_13642,N_13797);
nand U14492 (N_14492,N_13920,N_13793);
and U14493 (N_14493,N_13732,N_13641);
or U14494 (N_14494,N_13577,N_13703);
or U14495 (N_14495,N_13659,N_13743);
nand U14496 (N_14496,N_13539,N_13743);
or U14497 (N_14497,N_13910,N_13641);
nand U14498 (N_14498,N_13719,N_13756);
and U14499 (N_14499,N_13696,N_13545);
xor U14500 (N_14500,N_14171,N_14237);
nor U14501 (N_14501,N_14436,N_14486);
and U14502 (N_14502,N_14332,N_14450);
xnor U14503 (N_14503,N_14291,N_14434);
nand U14504 (N_14504,N_14438,N_14283);
or U14505 (N_14505,N_14489,N_14317);
nand U14506 (N_14506,N_14012,N_14149);
and U14507 (N_14507,N_14399,N_14370);
nand U14508 (N_14508,N_14123,N_14202);
xor U14509 (N_14509,N_14040,N_14181);
and U14510 (N_14510,N_14016,N_14282);
nand U14511 (N_14511,N_14253,N_14327);
nand U14512 (N_14512,N_14114,N_14239);
nand U14513 (N_14513,N_14274,N_14300);
nand U14514 (N_14514,N_14475,N_14107);
and U14515 (N_14515,N_14432,N_14176);
and U14516 (N_14516,N_14083,N_14211);
xnor U14517 (N_14517,N_14135,N_14374);
xor U14518 (N_14518,N_14014,N_14364);
xnor U14519 (N_14519,N_14246,N_14241);
and U14520 (N_14520,N_14119,N_14074);
or U14521 (N_14521,N_14189,N_14265);
or U14522 (N_14522,N_14234,N_14196);
xnor U14523 (N_14523,N_14396,N_14367);
or U14524 (N_14524,N_14067,N_14426);
nor U14525 (N_14525,N_14254,N_14104);
nand U14526 (N_14526,N_14159,N_14092);
and U14527 (N_14527,N_14279,N_14113);
xor U14528 (N_14528,N_14140,N_14470);
nor U14529 (N_14529,N_14389,N_14466);
and U14530 (N_14530,N_14105,N_14025);
nor U14531 (N_14531,N_14043,N_14368);
nor U14532 (N_14532,N_14244,N_14095);
nor U14533 (N_14533,N_14433,N_14405);
and U14534 (N_14534,N_14215,N_14194);
nor U14535 (N_14535,N_14122,N_14472);
nor U14536 (N_14536,N_14264,N_14278);
xor U14537 (N_14537,N_14125,N_14380);
nand U14538 (N_14538,N_14035,N_14027);
nor U14539 (N_14539,N_14046,N_14467);
nand U14540 (N_14540,N_14216,N_14406);
or U14541 (N_14541,N_14423,N_14032);
nor U14542 (N_14542,N_14387,N_14249);
or U14543 (N_14543,N_14259,N_14281);
and U14544 (N_14544,N_14328,N_14087);
nand U14545 (N_14545,N_14133,N_14156);
or U14546 (N_14546,N_14047,N_14318);
and U14547 (N_14547,N_14142,N_14401);
and U14548 (N_14548,N_14267,N_14086);
nand U14549 (N_14549,N_14349,N_14348);
and U14550 (N_14550,N_14424,N_14242);
xor U14551 (N_14551,N_14112,N_14337);
nand U14552 (N_14552,N_14121,N_14108);
and U14553 (N_14553,N_14497,N_14190);
and U14554 (N_14554,N_14333,N_14390);
nor U14555 (N_14555,N_14219,N_14444);
and U14556 (N_14556,N_14308,N_14447);
and U14557 (N_14557,N_14420,N_14193);
and U14558 (N_14558,N_14297,N_14311);
nand U14559 (N_14559,N_14397,N_14072);
or U14560 (N_14560,N_14115,N_14324);
nand U14561 (N_14561,N_14049,N_14468);
and U14562 (N_14562,N_14117,N_14048);
or U14563 (N_14563,N_14310,N_14091);
xnor U14564 (N_14564,N_14304,N_14052);
or U14565 (N_14565,N_14172,N_14245);
or U14566 (N_14566,N_14331,N_14482);
nor U14567 (N_14567,N_14440,N_14471);
and U14568 (N_14568,N_14428,N_14491);
xnor U14569 (N_14569,N_14417,N_14288);
nor U14570 (N_14570,N_14144,N_14136);
xnor U14571 (N_14571,N_14134,N_14314);
or U14572 (N_14572,N_14419,N_14312);
nor U14573 (N_14573,N_14320,N_14268);
nand U14574 (N_14574,N_14188,N_14442);
or U14575 (N_14575,N_14060,N_14285);
nor U14576 (N_14576,N_14127,N_14347);
and U14577 (N_14577,N_14453,N_14269);
xor U14578 (N_14578,N_14289,N_14151);
or U14579 (N_14579,N_14430,N_14200);
xnor U14580 (N_14580,N_14298,N_14058);
and U14581 (N_14581,N_14019,N_14010);
or U14582 (N_14582,N_14357,N_14197);
xor U14583 (N_14583,N_14295,N_14473);
and U14584 (N_14584,N_14326,N_14208);
xnor U14585 (N_14585,N_14089,N_14272);
nand U14586 (N_14586,N_14321,N_14462);
xor U14587 (N_14587,N_14170,N_14173);
nor U14588 (N_14588,N_14375,N_14483);
nor U14589 (N_14589,N_14338,N_14271);
or U14590 (N_14590,N_14139,N_14469);
nor U14591 (N_14591,N_14070,N_14340);
nand U14592 (N_14592,N_14229,N_14041);
xnor U14593 (N_14593,N_14076,N_14408);
nand U14594 (N_14594,N_14102,N_14429);
nand U14595 (N_14595,N_14223,N_14498);
xnor U14596 (N_14596,N_14400,N_14205);
nor U14597 (N_14597,N_14231,N_14131);
xor U14598 (N_14598,N_14100,N_14199);
or U14599 (N_14599,N_14198,N_14276);
nor U14600 (N_14600,N_14330,N_14454);
nand U14601 (N_14601,N_14339,N_14323);
and U14602 (N_14602,N_14038,N_14065);
and U14603 (N_14603,N_14110,N_14287);
and U14604 (N_14604,N_14243,N_14302);
or U14605 (N_14605,N_14451,N_14461);
nand U14606 (N_14606,N_14296,N_14413);
nand U14607 (N_14607,N_14132,N_14263);
xor U14608 (N_14608,N_14011,N_14177);
nand U14609 (N_14609,N_14233,N_14116);
or U14610 (N_14610,N_14230,N_14037);
or U14611 (N_14611,N_14093,N_14201);
nor U14612 (N_14612,N_14431,N_14416);
and U14613 (N_14613,N_14404,N_14062);
or U14614 (N_14614,N_14478,N_14388);
and U14615 (N_14615,N_14178,N_14409);
and U14616 (N_14616,N_14162,N_14218);
nand U14617 (N_14617,N_14250,N_14325);
nor U14618 (N_14618,N_14084,N_14290);
xor U14619 (N_14619,N_14359,N_14167);
and U14620 (N_14620,N_14316,N_14148);
and U14621 (N_14621,N_14164,N_14372);
nand U14622 (N_14622,N_14160,N_14183);
nor U14623 (N_14623,N_14459,N_14103);
nand U14624 (N_14624,N_14410,N_14382);
xnor U14625 (N_14625,N_14033,N_14336);
nor U14626 (N_14626,N_14306,N_14094);
nand U14627 (N_14627,N_14055,N_14280);
and U14628 (N_14628,N_14307,N_14363);
nand U14629 (N_14629,N_14376,N_14371);
nand U14630 (N_14630,N_14206,N_14068);
nor U14631 (N_14631,N_14299,N_14315);
xor U14632 (N_14632,N_14366,N_14111);
or U14633 (N_14633,N_14391,N_14365);
nand U14634 (N_14634,N_14488,N_14446);
and U14635 (N_14635,N_14228,N_14031);
and U14636 (N_14636,N_14154,N_14277);
nor U14637 (N_14637,N_14484,N_14079);
and U14638 (N_14638,N_14166,N_14377);
nand U14639 (N_14639,N_14036,N_14465);
or U14640 (N_14640,N_14002,N_14128);
or U14641 (N_14641,N_14448,N_14182);
nand U14642 (N_14642,N_14441,N_14018);
and U14643 (N_14643,N_14066,N_14152);
nand U14644 (N_14644,N_14443,N_14081);
xnor U14645 (N_14645,N_14313,N_14293);
nor U14646 (N_14646,N_14042,N_14088);
nand U14647 (N_14647,N_14480,N_14097);
xor U14648 (N_14648,N_14383,N_14493);
and U14649 (N_14649,N_14495,N_14227);
and U14650 (N_14650,N_14369,N_14212);
and U14651 (N_14651,N_14028,N_14085);
and U14652 (N_14652,N_14452,N_14207);
nor U14653 (N_14653,N_14210,N_14286);
and U14654 (N_14654,N_14179,N_14373);
or U14655 (N_14655,N_14007,N_14155);
and U14656 (N_14656,N_14098,N_14292);
xnor U14657 (N_14657,N_14120,N_14490);
nand U14658 (N_14658,N_14005,N_14456);
and U14659 (N_14659,N_14106,N_14309);
xor U14660 (N_14660,N_14004,N_14022);
and U14661 (N_14661,N_14096,N_14195);
xor U14662 (N_14662,N_14023,N_14213);
and U14663 (N_14663,N_14460,N_14270);
nor U14664 (N_14664,N_14222,N_14203);
xor U14665 (N_14665,N_14130,N_14184);
xnor U14666 (N_14666,N_14124,N_14024);
nand U14667 (N_14667,N_14064,N_14344);
nor U14668 (N_14668,N_14209,N_14251);
nor U14669 (N_14669,N_14356,N_14217);
and U14670 (N_14670,N_14256,N_14168);
nand U14671 (N_14671,N_14255,N_14192);
nor U14672 (N_14672,N_14494,N_14053);
xnor U14673 (N_14673,N_14071,N_14407);
xnor U14674 (N_14674,N_14225,N_14393);
and U14675 (N_14675,N_14358,N_14346);
nor U14676 (N_14676,N_14146,N_14392);
nand U14677 (N_14677,N_14191,N_14029);
or U14678 (N_14678,N_14044,N_14261);
nand U14679 (N_14679,N_14395,N_14214);
and U14680 (N_14680,N_14224,N_14141);
xor U14681 (N_14681,N_14476,N_14260);
nor U14682 (N_14682,N_14499,N_14017);
and U14683 (N_14683,N_14069,N_14487);
or U14684 (N_14684,N_14412,N_14034);
nand U14685 (N_14685,N_14050,N_14169);
xnor U14686 (N_14686,N_14474,N_14109);
nor U14687 (N_14687,N_14204,N_14161);
nand U14688 (N_14688,N_14258,N_14294);
nor U14689 (N_14689,N_14015,N_14051);
or U14690 (N_14690,N_14457,N_14303);
or U14691 (N_14691,N_14090,N_14013);
nor U14692 (N_14692,N_14252,N_14360);
nand U14693 (N_14693,N_14126,N_14449);
and U14694 (N_14694,N_14059,N_14354);
nand U14695 (N_14695,N_14057,N_14403);
or U14696 (N_14696,N_14350,N_14463);
nand U14697 (N_14697,N_14352,N_14235);
or U14698 (N_14698,N_14221,N_14163);
or U14699 (N_14699,N_14147,N_14003);
and U14700 (N_14700,N_14143,N_14398);
and U14701 (N_14701,N_14020,N_14361);
nand U14702 (N_14702,N_14341,N_14435);
and U14703 (N_14703,N_14266,N_14273);
and U14704 (N_14704,N_14077,N_14009);
nand U14705 (N_14705,N_14063,N_14030);
and U14706 (N_14706,N_14492,N_14165);
xor U14707 (N_14707,N_14080,N_14422);
xnor U14708 (N_14708,N_14437,N_14240);
nor U14709 (N_14709,N_14342,N_14355);
and U14710 (N_14710,N_14226,N_14334);
and U14711 (N_14711,N_14386,N_14138);
nand U14712 (N_14712,N_14187,N_14075);
and U14713 (N_14713,N_14150,N_14026);
and U14714 (N_14714,N_14481,N_14353);
and U14715 (N_14715,N_14394,N_14129);
xor U14716 (N_14716,N_14445,N_14322);
xor U14717 (N_14717,N_14137,N_14262);
nand U14718 (N_14718,N_14411,N_14073);
xnor U14719 (N_14719,N_14247,N_14001);
xnor U14720 (N_14720,N_14236,N_14061);
or U14721 (N_14721,N_14319,N_14275);
xnor U14722 (N_14722,N_14464,N_14101);
or U14723 (N_14723,N_14402,N_14118);
xnor U14724 (N_14724,N_14362,N_14000);
and U14725 (N_14725,N_14305,N_14335);
xor U14726 (N_14726,N_14099,N_14379);
or U14727 (N_14727,N_14006,N_14458);
nor U14728 (N_14728,N_14343,N_14496);
nor U14729 (N_14729,N_14439,N_14351);
nand U14730 (N_14730,N_14008,N_14345);
xnor U14731 (N_14731,N_14078,N_14180);
xnor U14732 (N_14732,N_14175,N_14145);
nand U14733 (N_14733,N_14418,N_14039);
and U14734 (N_14734,N_14329,N_14384);
xor U14735 (N_14735,N_14158,N_14381);
nor U14736 (N_14736,N_14421,N_14220);
nand U14737 (N_14737,N_14378,N_14021);
nand U14738 (N_14738,N_14257,N_14301);
xnor U14739 (N_14739,N_14056,N_14185);
nand U14740 (N_14740,N_14054,N_14385);
and U14741 (N_14741,N_14415,N_14232);
nor U14742 (N_14742,N_14186,N_14414);
nor U14743 (N_14743,N_14425,N_14284);
nor U14744 (N_14744,N_14485,N_14427);
or U14745 (N_14745,N_14477,N_14153);
nand U14746 (N_14746,N_14082,N_14174);
nand U14747 (N_14747,N_14455,N_14157);
and U14748 (N_14748,N_14238,N_14045);
xnor U14749 (N_14749,N_14479,N_14248);
or U14750 (N_14750,N_14349,N_14019);
and U14751 (N_14751,N_14168,N_14021);
nor U14752 (N_14752,N_14307,N_14131);
nand U14753 (N_14753,N_14040,N_14279);
and U14754 (N_14754,N_14456,N_14022);
or U14755 (N_14755,N_14240,N_14238);
nor U14756 (N_14756,N_14317,N_14350);
or U14757 (N_14757,N_14102,N_14296);
nand U14758 (N_14758,N_14460,N_14066);
and U14759 (N_14759,N_14320,N_14265);
nor U14760 (N_14760,N_14109,N_14267);
nor U14761 (N_14761,N_14470,N_14087);
or U14762 (N_14762,N_14449,N_14151);
xnor U14763 (N_14763,N_14364,N_14033);
xnor U14764 (N_14764,N_14324,N_14357);
and U14765 (N_14765,N_14334,N_14353);
nand U14766 (N_14766,N_14179,N_14490);
and U14767 (N_14767,N_14475,N_14052);
and U14768 (N_14768,N_14202,N_14084);
and U14769 (N_14769,N_14029,N_14480);
or U14770 (N_14770,N_14021,N_14339);
nor U14771 (N_14771,N_14159,N_14103);
nor U14772 (N_14772,N_14049,N_14239);
and U14773 (N_14773,N_14011,N_14183);
or U14774 (N_14774,N_14469,N_14293);
or U14775 (N_14775,N_14059,N_14050);
and U14776 (N_14776,N_14272,N_14115);
or U14777 (N_14777,N_14283,N_14355);
and U14778 (N_14778,N_14005,N_14276);
nor U14779 (N_14779,N_14457,N_14065);
xnor U14780 (N_14780,N_14203,N_14155);
or U14781 (N_14781,N_14193,N_14318);
nor U14782 (N_14782,N_14317,N_14365);
nor U14783 (N_14783,N_14427,N_14492);
or U14784 (N_14784,N_14344,N_14091);
and U14785 (N_14785,N_14281,N_14069);
or U14786 (N_14786,N_14417,N_14429);
and U14787 (N_14787,N_14058,N_14158);
and U14788 (N_14788,N_14233,N_14257);
nor U14789 (N_14789,N_14374,N_14203);
xnor U14790 (N_14790,N_14407,N_14474);
and U14791 (N_14791,N_14461,N_14025);
xnor U14792 (N_14792,N_14059,N_14440);
nand U14793 (N_14793,N_14327,N_14087);
xnor U14794 (N_14794,N_14190,N_14165);
xor U14795 (N_14795,N_14382,N_14306);
xor U14796 (N_14796,N_14145,N_14371);
nand U14797 (N_14797,N_14229,N_14145);
nor U14798 (N_14798,N_14486,N_14150);
or U14799 (N_14799,N_14050,N_14147);
nor U14800 (N_14800,N_14354,N_14211);
nand U14801 (N_14801,N_14406,N_14222);
xnor U14802 (N_14802,N_14234,N_14327);
and U14803 (N_14803,N_14289,N_14302);
nor U14804 (N_14804,N_14204,N_14229);
or U14805 (N_14805,N_14168,N_14091);
or U14806 (N_14806,N_14217,N_14006);
xor U14807 (N_14807,N_14424,N_14324);
nor U14808 (N_14808,N_14199,N_14363);
and U14809 (N_14809,N_14072,N_14469);
or U14810 (N_14810,N_14392,N_14416);
nor U14811 (N_14811,N_14091,N_14164);
xnor U14812 (N_14812,N_14095,N_14424);
and U14813 (N_14813,N_14037,N_14015);
nor U14814 (N_14814,N_14268,N_14041);
or U14815 (N_14815,N_14406,N_14274);
or U14816 (N_14816,N_14095,N_14260);
nand U14817 (N_14817,N_14304,N_14260);
nand U14818 (N_14818,N_14062,N_14045);
nand U14819 (N_14819,N_14059,N_14460);
and U14820 (N_14820,N_14337,N_14423);
nand U14821 (N_14821,N_14439,N_14014);
nand U14822 (N_14822,N_14323,N_14251);
nand U14823 (N_14823,N_14175,N_14392);
xor U14824 (N_14824,N_14081,N_14249);
nand U14825 (N_14825,N_14094,N_14270);
and U14826 (N_14826,N_14381,N_14428);
or U14827 (N_14827,N_14261,N_14292);
or U14828 (N_14828,N_14057,N_14088);
and U14829 (N_14829,N_14172,N_14338);
xnor U14830 (N_14830,N_14369,N_14357);
and U14831 (N_14831,N_14320,N_14402);
xor U14832 (N_14832,N_14024,N_14320);
or U14833 (N_14833,N_14139,N_14451);
nor U14834 (N_14834,N_14366,N_14162);
or U14835 (N_14835,N_14287,N_14201);
nand U14836 (N_14836,N_14313,N_14051);
nor U14837 (N_14837,N_14425,N_14094);
or U14838 (N_14838,N_14078,N_14263);
nor U14839 (N_14839,N_14492,N_14108);
nor U14840 (N_14840,N_14042,N_14303);
and U14841 (N_14841,N_14002,N_14471);
xnor U14842 (N_14842,N_14047,N_14164);
nand U14843 (N_14843,N_14377,N_14034);
xnor U14844 (N_14844,N_14026,N_14263);
or U14845 (N_14845,N_14012,N_14261);
xor U14846 (N_14846,N_14362,N_14407);
and U14847 (N_14847,N_14189,N_14060);
nor U14848 (N_14848,N_14382,N_14299);
xnor U14849 (N_14849,N_14093,N_14004);
or U14850 (N_14850,N_14040,N_14434);
and U14851 (N_14851,N_14422,N_14327);
and U14852 (N_14852,N_14006,N_14412);
and U14853 (N_14853,N_14479,N_14235);
and U14854 (N_14854,N_14475,N_14236);
or U14855 (N_14855,N_14444,N_14358);
nor U14856 (N_14856,N_14451,N_14201);
xor U14857 (N_14857,N_14400,N_14336);
or U14858 (N_14858,N_14186,N_14273);
or U14859 (N_14859,N_14079,N_14249);
nand U14860 (N_14860,N_14457,N_14147);
or U14861 (N_14861,N_14476,N_14007);
and U14862 (N_14862,N_14372,N_14052);
and U14863 (N_14863,N_14390,N_14269);
nand U14864 (N_14864,N_14139,N_14317);
xnor U14865 (N_14865,N_14204,N_14074);
or U14866 (N_14866,N_14257,N_14359);
nor U14867 (N_14867,N_14383,N_14233);
and U14868 (N_14868,N_14489,N_14222);
and U14869 (N_14869,N_14151,N_14343);
xnor U14870 (N_14870,N_14145,N_14036);
nor U14871 (N_14871,N_14221,N_14168);
nor U14872 (N_14872,N_14057,N_14282);
and U14873 (N_14873,N_14004,N_14436);
xor U14874 (N_14874,N_14492,N_14410);
xnor U14875 (N_14875,N_14109,N_14089);
xor U14876 (N_14876,N_14183,N_14380);
or U14877 (N_14877,N_14164,N_14296);
nand U14878 (N_14878,N_14244,N_14080);
nand U14879 (N_14879,N_14220,N_14392);
xor U14880 (N_14880,N_14243,N_14102);
xor U14881 (N_14881,N_14185,N_14146);
xor U14882 (N_14882,N_14054,N_14066);
xor U14883 (N_14883,N_14460,N_14350);
nand U14884 (N_14884,N_14326,N_14106);
and U14885 (N_14885,N_14409,N_14298);
nand U14886 (N_14886,N_14296,N_14370);
nor U14887 (N_14887,N_14442,N_14337);
nand U14888 (N_14888,N_14499,N_14346);
nand U14889 (N_14889,N_14205,N_14461);
nand U14890 (N_14890,N_14097,N_14437);
or U14891 (N_14891,N_14169,N_14137);
xor U14892 (N_14892,N_14307,N_14489);
nand U14893 (N_14893,N_14306,N_14060);
xnor U14894 (N_14894,N_14333,N_14438);
or U14895 (N_14895,N_14069,N_14273);
nand U14896 (N_14896,N_14150,N_14441);
nor U14897 (N_14897,N_14240,N_14332);
xor U14898 (N_14898,N_14255,N_14201);
xor U14899 (N_14899,N_14286,N_14311);
and U14900 (N_14900,N_14143,N_14175);
xnor U14901 (N_14901,N_14408,N_14189);
and U14902 (N_14902,N_14099,N_14027);
nor U14903 (N_14903,N_14382,N_14335);
nand U14904 (N_14904,N_14448,N_14404);
and U14905 (N_14905,N_14426,N_14270);
or U14906 (N_14906,N_14332,N_14213);
nor U14907 (N_14907,N_14117,N_14420);
and U14908 (N_14908,N_14091,N_14055);
and U14909 (N_14909,N_14091,N_14048);
and U14910 (N_14910,N_14038,N_14131);
xnor U14911 (N_14911,N_14043,N_14400);
or U14912 (N_14912,N_14192,N_14263);
and U14913 (N_14913,N_14227,N_14337);
or U14914 (N_14914,N_14421,N_14490);
and U14915 (N_14915,N_14114,N_14012);
or U14916 (N_14916,N_14102,N_14096);
nor U14917 (N_14917,N_14255,N_14359);
xnor U14918 (N_14918,N_14369,N_14001);
xnor U14919 (N_14919,N_14082,N_14495);
xnor U14920 (N_14920,N_14142,N_14361);
nand U14921 (N_14921,N_14284,N_14105);
nand U14922 (N_14922,N_14025,N_14060);
or U14923 (N_14923,N_14181,N_14236);
xnor U14924 (N_14924,N_14095,N_14104);
or U14925 (N_14925,N_14451,N_14024);
or U14926 (N_14926,N_14088,N_14489);
nor U14927 (N_14927,N_14078,N_14436);
or U14928 (N_14928,N_14370,N_14419);
xor U14929 (N_14929,N_14254,N_14264);
xnor U14930 (N_14930,N_14287,N_14024);
and U14931 (N_14931,N_14114,N_14258);
xnor U14932 (N_14932,N_14439,N_14451);
and U14933 (N_14933,N_14168,N_14204);
or U14934 (N_14934,N_14432,N_14450);
and U14935 (N_14935,N_14108,N_14469);
nand U14936 (N_14936,N_14266,N_14199);
and U14937 (N_14937,N_14049,N_14423);
or U14938 (N_14938,N_14044,N_14397);
nand U14939 (N_14939,N_14292,N_14290);
or U14940 (N_14940,N_14121,N_14319);
nand U14941 (N_14941,N_14321,N_14255);
or U14942 (N_14942,N_14168,N_14038);
nor U14943 (N_14943,N_14463,N_14036);
xnor U14944 (N_14944,N_14254,N_14474);
xnor U14945 (N_14945,N_14450,N_14104);
and U14946 (N_14946,N_14358,N_14290);
xor U14947 (N_14947,N_14041,N_14364);
xor U14948 (N_14948,N_14186,N_14325);
nor U14949 (N_14949,N_14186,N_14043);
or U14950 (N_14950,N_14299,N_14016);
xor U14951 (N_14951,N_14045,N_14125);
and U14952 (N_14952,N_14299,N_14368);
and U14953 (N_14953,N_14124,N_14294);
and U14954 (N_14954,N_14326,N_14034);
nor U14955 (N_14955,N_14250,N_14498);
nand U14956 (N_14956,N_14077,N_14499);
or U14957 (N_14957,N_14285,N_14231);
xor U14958 (N_14958,N_14049,N_14485);
nor U14959 (N_14959,N_14370,N_14138);
nor U14960 (N_14960,N_14316,N_14204);
and U14961 (N_14961,N_14074,N_14133);
nor U14962 (N_14962,N_14394,N_14474);
xor U14963 (N_14963,N_14272,N_14304);
xnor U14964 (N_14964,N_14209,N_14377);
or U14965 (N_14965,N_14398,N_14013);
or U14966 (N_14966,N_14436,N_14345);
and U14967 (N_14967,N_14382,N_14409);
and U14968 (N_14968,N_14242,N_14153);
or U14969 (N_14969,N_14067,N_14478);
nor U14970 (N_14970,N_14492,N_14098);
xor U14971 (N_14971,N_14055,N_14328);
and U14972 (N_14972,N_14401,N_14241);
nand U14973 (N_14973,N_14256,N_14369);
and U14974 (N_14974,N_14377,N_14241);
nand U14975 (N_14975,N_14389,N_14205);
nor U14976 (N_14976,N_14418,N_14274);
nand U14977 (N_14977,N_14306,N_14422);
nor U14978 (N_14978,N_14318,N_14483);
nor U14979 (N_14979,N_14289,N_14453);
xnor U14980 (N_14980,N_14161,N_14155);
nor U14981 (N_14981,N_14200,N_14270);
nand U14982 (N_14982,N_14361,N_14499);
nand U14983 (N_14983,N_14029,N_14333);
or U14984 (N_14984,N_14493,N_14483);
or U14985 (N_14985,N_14193,N_14177);
or U14986 (N_14986,N_14353,N_14448);
xor U14987 (N_14987,N_14061,N_14399);
and U14988 (N_14988,N_14082,N_14421);
nand U14989 (N_14989,N_14159,N_14491);
and U14990 (N_14990,N_14478,N_14444);
nand U14991 (N_14991,N_14452,N_14310);
nand U14992 (N_14992,N_14400,N_14038);
nand U14993 (N_14993,N_14170,N_14149);
nor U14994 (N_14994,N_14437,N_14353);
nand U14995 (N_14995,N_14049,N_14275);
or U14996 (N_14996,N_14057,N_14081);
nand U14997 (N_14997,N_14278,N_14137);
nand U14998 (N_14998,N_14003,N_14124);
nand U14999 (N_14999,N_14356,N_14439);
xor UO_0 (O_0,N_14807,N_14515);
nor UO_1 (O_1,N_14979,N_14651);
nor UO_2 (O_2,N_14985,N_14608);
xnor UO_3 (O_3,N_14720,N_14614);
xor UO_4 (O_4,N_14972,N_14679);
nand UO_5 (O_5,N_14819,N_14935);
nor UO_6 (O_6,N_14663,N_14609);
and UO_7 (O_7,N_14616,N_14711);
nor UO_8 (O_8,N_14909,N_14622);
nor UO_9 (O_9,N_14648,N_14662);
and UO_10 (O_10,N_14895,N_14846);
xor UO_11 (O_11,N_14564,N_14824);
nand UO_12 (O_12,N_14588,N_14913);
xor UO_13 (O_13,N_14607,N_14921);
xor UO_14 (O_14,N_14559,N_14767);
xnor UO_15 (O_15,N_14831,N_14745);
xnor UO_16 (O_16,N_14579,N_14874);
xor UO_17 (O_17,N_14601,N_14649);
and UO_18 (O_18,N_14790,N_14587);
and UO_19 (O_19,N_14631,N_14511);
nor UO_20 (O_20,N_14995,N_14522);
nand UO_21 (O_21,N_14630,N_14748);
nand UO_22 (O_22,N_14721,N_14696);
xor UO_23 (O_23,N_14503,N_14771);
xor UO_24 (O_24,N_14710,N_14857);
nor UO_25 (O_25,N_14956,N_14593);
nand UO_26 (O_26,N_14504,N_14611);
nor UO_27 (O_27,N_14890,N_14791);
nor UO_28 (O_28,N_14993,N_14835);
nor UO_29 (O_29,N_14570,N_14741);
nor UO_30 (O_30,N_14541,N_14534);
or UO_31 (O_31,N_14849,N_14848);
and UO_32 (O_32,N_14715,N_14976);
nor UO_33 (O_33,N_14730,N_14619);
and UO_34 (O_34,N_14658,N_14743);
or UO_35 (O_35,N_14539,N_14908);
and UO_36 (O_36,N_14508,N_14637);
xor UO_37 (O_37,N_14644,N_14784);
nand UO_38 (O_38,N_14944,N_14932);
nand UO_39 (O_39,N_14900,N_14678);
or UO_40 (O_40,N_14999,N_14950);
nor UO_41 (O_41,N_14867,N_14598);
or UO_42 (O_42,N_14983,N_14912);
and UO_43 (O_43,N_14762,N_14596);
or UO_44 (O_44,N_14783,N_14738);
and UO_45 (O_45,N_14952,N_14684);
nand UO_46 (O_46,N_14603,N_14506);
nor UO_47 (O_47,N_14967,N_14776);
and UO_48 (O_48,N_14914,N_14657);
or UO_49 (O_49,N_14665,N_14761);
nand UO_50 (O_50,N_14575,N_14864);
or UO_51 (O_51,N_14886,N_14572);
or UO_52 (O_52,N_14706,N_14804);
or UO_53 (O_53,N_14645,N_14671);
and UO_54 (O_54,N_14747,N_14977);
or UO_55 (O_55,N_14759,N_14936);
xnor UO_56 (O_56,N_14951,N_14732);
or UO_57 (O_57,N_14646,N_14899);
and UO_58 (O_58,N_14590,N_14975);
and UO_59 (O_59,N_14659,N_14566);
or UO_60 (O_60,N_14964,N_14940);
nor UO_61 (O_61,N_14773,N_14638);
or UO_62 (O_62,N_14957,N_14612);
nand UO_63 (O_63,N_14941,N_14827);
or UO_64 (O_64,N_14898,N_14581);
or UO_65 (O_65,N_14529,N_14680);
or UO_66 (O_66,N_14713,N_14793);
xnor UO_67 (O_67,N_14726,N_14821);
nor UO_68 (O_68,N_14871,N_14959);
and UO_69 (O_69,N_14961,N_14571);
nor UO_70 (O_70,N_14606,N_14592);
or UO_71 (O_71,N_14891,N_14643);
nor UO_72 (O_72,N_14946,N_14675);
nand UO_73 (O_73,N_14699,N_14868);
or UO_74 (O_74,N_14829,N_14814);
nor UO_75 (O_75,N_14780,N_14876);
nand UO_76 (O_76,N_14958,N_14798);
nand UO_77 (O_77,N_14683,N_14580);
or UO_78 (O_78,N_14526,N_14740);
and UO_79 (O_79,N_14754,N_14558);
and UO_80 (O_80,N_14752,N_14654);
or UO_81 (O_81,N_14772,N_14613);
nand UO_82 (O_82,N_14577,N_14527);
or UO_83 (O_83,N_14576,N_14830);
xnor UO_84 (O_84,N_14974,N_14756);
and UO_85 (O_85,N_14755,N_14992);
or UO_86 (O_86,N_14927,N_14567);
nand UO_87 (O_87,N_14618,N_14668);
nand UO_88 (O_88,N_14920,N_14938);
xnor UO_89 (O_89,N_14750,N_14694);
or UO_90 (O_90,N_14833,N_14537);
xnor UO_91 (O_91,N_14962,N_14569);
and UO_92 (O_92,N_14602,N_14859);
and UO_93 (O_93,N_14971,N_14794);
nor UO_94 (O_94,N_14758,N_14695);
and UO_95 (O_95,N_14705,N_14542);
and UO_96 (O_96,N_14573,N_14800);
or UO_97 (O_97,N_14718,N_14945);
or UO_98 (O_98,N_14931,N_14882);
nor UO_99 (O_99,N_14937,N_14548);
xor UO_100 (O_100,N_14734,N_14700);
and UO_101 (O_101,N_14692,N_14782);
nor UO_102 (O_102,N_14698,N_14666);
nor UO_103 (O_103,N_14656,N_14520);
xnor UO_104 (O_104,N_14978,N_14884);
or UO_105 (O_105,N_14716,N_14781);
or UO_106 (O_106,N_14948,N_14546);
and UO_107 (O_107,N_14840,N_14547);
nor UO_108 (O_108,N_14688,N_14701);
and UO_109 (O_109,N_14507,N_14556);
or UO_110 (O_110,N_14954,N_14610);
nor UO_111 (O_111,N_14928,N_14632);
and UO_112 (O_112,N_14885,N_14739);
and UO_113 (O_113,N_14652,N_14930);
and UO_114 (O_114,N_14640,N_14918);
xnor UO_115 (O_115,N_14565,N_14682);
nor UO_116 (O_116,N_14841,N_14685);
nor UO_117 (O_117,N_14865,N_14766);
xor UO_118 (O_118,N_14902,N_14810);
or UO_119 (O_119,N_14820,N_14779);
and UO_120 (O_120,N_14822,N_14560);
or UO_121 (O_121,N_14998,N_14774);
and UO_122 (O_122,N_14788,N_14990);
or UO_123 (O_123,N_14687,N_14719);
xnor UO_124 (O_124,N_14812,N_14872);
xor UO_125 (O_125,N_14866,N_14929);
nor UO_126 (O_126,N_14697,N_14655);
nand UO_127 (O_127,N_14896,N_14621);
and UO_128 (O_128,N_14667,N_14844);
xor UO_129 (O_129,N_14917,N_14904);
nand UO_130 (O_130,N_14586,N_14862);
xnor UO_131 (O_131,N_14691,N_14943);
nor UO_132 (O_132,N_14723,N_14763);
or UO_133 (O_133,N_14714,N_14737);
xnor UO_134 (O_134,N_14531,N_14858);
and UO_135 (O_135,N_14991,N_14681);
xnor UO_136 (O_136,N_14605,N_14839);
xor UO_137 (O_137,N_14629,N_14635);
nand UO_138 (O_138,N_14792,N_14832);
or UO_139 (O_139,N_14851,N_14802);
or UO_140 (O_140,N_14994,N_14735);
xnor UO_141 (O_141,N_14597,N_14906);
xnor UO_142 (O_142,N_14777,N_14669);
xnor UO_143 (O_143,N_14799,N_14768);
nor UO_144 (O_144,N_14518,N_14717);
nor UO_145 (O_145,N_14627,N_14551);
nand UO_146 (O_146,N_14731,N_14924);
nand UO_147 (O_147,N_14984,N_14554);
xor UO_148 (O_148,N_14778,N_14563);
or UO_149 (O_149,N_14543,N_14980);
nor UO_150 (O_150,N_14838,N_14500);
or UO_151 (O_151,N_14892,N_14801);
xor UO_152 (O_152,N_14516,N_14555);
and UO_153 (O_153,N_14642,N_14639);
xnor UO_154 (O_154,N_14834,N_14532);
nand UO_155 (O_155,N_14969,N_14806);
nand UO_156 (O_156,N_14594,N_14815);
xnor UO_157 (O_157,N_14519,N_14949);
or UO_158 (O_158,N_14797,N_14770);
and UO_159 (O_159,N_14540,N_14625);
nand UO_160 (O_160,N_14836,N_14973);
nor UO_161 (O_161,N_14769,N_14702);
xnor UO_162 (O_162,N_14524,N_14916);
nor UO_163 (O_163,N_14672,N_14953);
nand UO_164 (O_164,N_14880,N_14686);
and UO_165 (O_165,N_14585,N_14881);
xor UO_166 (O_166,N_14856,N_14837);
and UO_167 (O_167,N_14550,N_14907);
and UO_168 (O_168,N_14863,N_14617);
or UO_169 (O_169,N_14968,N_14996);
xor UO_170 (O_170,N_14510,N_14877);
or UO_171 (O_171,N_14879,N_14786);
nor UO_172 (O_172,N_14873,N_14725);
nor UO_173 (O_173,N_14966,N_14536);
nand UO_174 (O_174,N_14724,N_14842);
nor UO_175 (O_175,N_14578,N_14703);
or UO_176 (O_176,N_14751,N_14796);
nor UO_177 (O_177,N_14561,N_14523);
xnor UO_178 (O_178,N_14533,N_14988);
and UO_179 (O_179,N_14600,N_14947);
or UO_180 (O_180,N_14982,N_14826);
and UO_181 (O_181,N_14805,N_14589);
xnor UO_182 (O_182,N_14521,N_14733);
xor UO_183 (O_183,N_14664,N_14549);
nand UO_184 (O_184,N_14599,N_14729);
nor UO_185 (O_185,N_14736,N_14502);
nand UO_186 (O_186,N_14843,N_14704);
or UO_187 (O_187,N_14512,N_14942);
or UO_188 (O_188,N_14562,N_14795);
nor UO_189 (O_189,N_14584,N_14513);
xnor UO_190 (O_190,N_14981,N_14661);
or UO_191 (O_191,N_14901,N_14789);
or UO_192 (O_192,N_14574,N_14997);
nand UO_193 (O_193,N_14897,N_14626);
nor UO_194 (O_194,N_14887,N_14845);
nand UO_195 (O_195,N_14785,N_14987);
and UO_196 (O_196,N_14673,N_14525);
or UO_197 (O_197,N_14825,N_14960);
xor UO_198 (O_198,N_14939,N_14615);
nand UO_199 (O_199,N_14728,N_14553);
and UO_200 (O_200,N_14816,N_14746);
nand UO_201 (O_201,N_14808,N_14530);
nor UO_202 (O_202,N_14852,N_14878);
and UO_203 (O_203,N_14883,N_14923);
nor UO_204 (O_204,N_14568,N_14860);
and UO_205 (O_205,N_14674,N_14538);
and UO_206 (O_206,N_14787,N_14727);
nand UO_207 (O_207,N_14650,N_14889);
nand UO_208 (O_208,N_14636,N_14628);
or UO_209 (O_209,N_14963,N_14850);
xnor UO_210 (O_210,N_14813,N_14818);
or UO_211 (O_211,N_14811,N_14823);
or UO_212 (O_212,N_14875,N_14634);
xnor UO_213 (O_213,N_14544,N_14653);
or UO_214 (O_214,N_14582,N_14828);
or UO_215 (O_215,N_14855,N_14693);
nor UO_216 (O_216,N_14517,N_14552);
or UO_217 (O_217,N_14809,N_14712);
nor UO_218 (O_218,N_14709,N_14919);
xor UO_219 (O_219,N_14620,N_14604);
and UO_220 (O_220,N_14744,N_14911);
nand UO_221 (O_221,N_14677,N_14633);
nor UO_222 (O_222,N_14869,N_14595);
xor UO_223 (O_223,N_14915,N_14535);
or UO_224 (O_224,N_14528,N_14986);
nor UO_225 (O_225,N_14765,N_14870);
nand UO_226 (O_226,N_14505,N_14749);
xor UO_227 (O_227,N_14903,N_14853);
nand UO_228 (O_228,N_14757,N_14583);
and UO_229 (O_229,N_14847,N_14933);
or UO_230 (O_230,N_14641,N_14514);
nor UO_231 (O_231,N_14910,N_14970);
and UO_232 (O_232,N_14955,N_14925);
nand UO_233 (O_233,N_14707,N_14965);
nand UO_234 (O_234,N_14989,N_14854);
nand UO_235 (O_235,N_14509,N_14926);
nor UO_236 (O_236,N_14545,N_14501);
nand UO_237 (O_237,N_14690,N_14760);
nand UO_238 (O_238,N_14905,N_14722);
and UO_239 (O_239,N_14623,N_14803);
and UO_240 (O_240,N_14676,N_14591);
or UO_241 (O_241,N_14894,N_14742);
xnor UO_242 (O_242,N_14753,N_14624);
nor UO_243 (O_243,N_14660,N_14764);
and UO_244 (O_244,N_14861,N_14647);
and UO_245 (O_245,N_14670,N_14689);
xnor UO_246 (O_246,N_14922,N_14708);
nor UO_247 (O_247,N_14893,N_14817);
nor UO_248 (O_248,N_14934,N_14775);
or UO_249 (O_249,N_14557,N_14888);
and UO_250 (O_250,N_14862,N_14807);
or UO_251 (O_251,N_14931,N_14547);
xor UO_252 (O_252,N_14714,N_14738);
xor UO_253 (O_253,N_14848,N_14603);
nor UO_254 (O_254,N_14857,N_14736);
nor UO_255 (O_255,N_14881,N_14539);
xor UO_256 (O_256,N_14901,N_14862);
and UO_257 (O_257,N_14783,N_14981);
nor UO_258 (O_258,N_14958,N_14668);
nor UO_259 (O_259,N_14579,N_14583);
and UO_260 (O_260,N_14689,N_14719);
nand UO_261 (O_261,N_14945,N_14677);
or UO_262 (O_262,N_14595,N_14889);
nand UO_263 (O_263,N_14576,N_14912);
and UO_264 (O_264,N_14872,N_14875);
and UO_265 (O_265,N_14631,N_14966);
nor UO_266 (O_266,N_14630,N_14917);
nand UO_267 (O_267,N_14756,N_14794);
or UO_268 (O_268,N_14972,N_14632);
and UO_269 (O_269,N_14508,N_14560);
or UO_270 (O_270,N_14766,N_14932);
and UO_271 (O_271,N_14627,N_14987);
and UO_272 (O_272,N_14600,N_14984);
nand UO_273 (O_273,N_14524,N_14639);
nor UO_274 (O_274,N_14582,N_14829);
or UO_275 (O_275,N_14962,N_14758);
or UO_276 (O_276,N_14547,N_14937);
xnor UO_277 (O_277,N_14635,N_14579);
and UO_278 (O_278,N_14554,N_14823);
or UO_279 (O_279,N_14765,N_14806);
and UO_280 (O_280,N_14718,N_14684);
xor UO_281 (O_281,N_14888,N_14551);
nor UO_282 (O_282,N_14952,N_14598);
nand UO_283 (O_283,N_14574,N_14853);
nand UO_284 (O_284,N_14669,N_14920);
nor UO_285 (O_285,N_14613,N_14688);
xnor UO_286 (O_286,N_14567,N_14648);
and UO_287 (O_287,N_14562,N_14746);
xor UO_288 (O_288,N_14587,N_14605);
xnor UO_289 (O_289,N_14798,N_14782);
nand UO_290 (O_290,N_14792,N_14628);
or UO_291 (O_291,N_14974,N_14737);
or UO_292 (O_292,N_14627,N_14575);
nor UO_293 (O_293,N_14623,N_14990);
nand UO_294 (O_294,N_14527,N_14861);
nor UO_295 (O_295,N_14965,N_14853);
xnor UO_296 (O_296,N_14589,N_14673);
xnor UO_297 (O_297,N_14941,N_14542);
nand UO_298 (O_298,N_14768,N_14630);
xor UO_299 (O_299,N_14893,N_14598);
or UO_300 (O_300,N_14933,N_14964);
or UO_301 (O_301,N_14885,N_14838);
xor UO_302 (O_302,N_14618,N_14898);
xnor UO_303 (O_303,N_14570,N_14980);
xnor UO_304 (O_304,N_14930,N_14877);
xnor UO_305 (O_305,N_14879,N_14890);
xor UO_306 (O_306,N_14661,N_14938);
nor UO_307 (O_307,N_14697,N_14590);
nand UO_308 (O_308,N_14905,N_14624);
xor UO_309 (O_309,N_14791,N_14516);
nand UO_310 (O_310,N_14589,N_14987);
nor UO_311 (O_311,N_14915,N_14716);
xor UO_312 (O_312,N_14897,N_14611);
nor UO_313 (O_313,N_14953,N_14958);
nor UO_314 (O_314,N_14929,N_14542);
nor UO_315 (O_315,N_14612,N_14817);
or UO_316 (O_316,N_14812,N_14784);
and UO_317 (O_317,N_14513,N_14857);
or UO_318 (O_318,N_14840,N_14898);
xnor UO_319 (O_319,N_14938,N_14681);
nor UO_320 (O_320,N_14620,N_14807);
nand UO_321 (O_321,N_14878,N_14762);
or UO_322 (O_322,N_14700,N_14554);
nand UO_323 (O_323,N_14906,N_14995);
or UO_324 (O_324,N_14837,N_14542);
nand UO_325 (O_325,N_14853,N_14816);
xor UO_326 (O_326,N_14998,N_14866);
and UO_327 (O_327,N_14600,N_14951);
or UO_328 (O_328,N_14764,N_14716);
or UO_329 (O_329,N_14585,N_14718);
xnor UO_330 (O_330,N_14646,N_14963);
nand UO_331 (O_331,N_14826,N_14981);
nand UO_332 (O_332,N_14796,N_14645);
nor UO_333 (O_333,N_14890,N_14535);
xnor UO_334 (O_334,N_14899,N_14679);
xnor UO_335 (O_335,N_14999,N_14982);
xor UO_336 (O_336,N_14928,N_14853);
nand UO_337 (O_337,N_14850,N_14907);
nand UO_338 (O_338,N_14893,N_14861);
nand UO_339 (O_339,N_14551,N_14776);
nand UO_340 (O_340,N_14712,N_14863);
nand UO_341 (O_341,N_14775,N_14894);
or UO_342 (O_342,N_14502,N_14671);
nand UO_343 (O_343,N_14686,N_14883);
or UO_344 (O_344,N_14529,N_14799);
nand UO_345 (O_345,N_14951,N_14626);
nand UO_346 (O_346,N_14785,N_14674);
nor UO_347 (O_347,N_14865,N_14765);
nor UO_348 (O_348,N_14814,N_14664);
nand UO_349 (O_349,N_14744,N_14566);
nand UO_350 (O_350,N_14952,N_14643);
xnor UO_351 (O_351,N_14511,N_14841);
nand UO_352 (O_352,N_14840,N_14884);
nor UO_353 (O_353,N_14814,N_14912);
nor UO_354 (O_354,N_14527,N_14906);
and UO_355 (O_355,N_14676,N_14820);
xor UO_356 (O_356,N_14908,N_14569);
xnor UO_357 (O_357,N_14924,N_14640);
xnor UO_358 (O_358,N_14820,N_14600);
and UO_359 (O_359,N_14961,N_14738);
nor UO_360 (O_360,N_14855,N_14961);
or UO_361 (O_361,N_14597,N_14988);
nand UO_362 (O_362,N_14632,N_14608);
xor UO_363 (O_363,N_14690,N_14872);
and UO_364 (O_364,N_14966,N_14805);
nor UO_365 (O_365,N_14680,N_14902);
or UO_366 (O_366,N_14849,N_14550);
or UO_367 (O_367,N_14732,N_14534);
xor UO_368 (O_368,N_14922,N_14678);
nand UO_369 (O_369,N_14528,N_14909);
xor UO_370 (O_370,N_14989,N_14604);
or UO_371 (O_371,N_14656,N_14581);
or UO_372 (O_372,N_14846,N_14667);
nand UO_373 (O_373,N_14587,N_14764);
and UO_374 (O_374,N_14528,N_14533);
and UO_375 (O_375,N_14611,N_14610);
xnor UO_376 (O_376,N_14975,N_14581);
xnor UO_377 (O_377,N_14851,N_14853);
nor UO_378 (O_378,N_14592,N_14792);
and UO_379 (O_379,N_14608,N_14824);
or UO_380 (O_380,N_14730,N_14596);
or UO_381 (O_381,N_14873,N_14569);
nand UO_382 (O_382,N_14900,N_14770);
or UO_383 (O_383,N_14771,N_14547);
xnor UO_384 (O_384,N_14728,N_14580);
nor UO_385 (O_385,N_14700,N_14592);
xnor UO_386 (O_386,N_14541,N_14982);
nor UO_387 (O_387,N_14602,N_14732);
and UO_388 (O_388,N_14619,N_14795);
xor UO_389 (O_389,N_14607,N_14571);
xnor UO_390 (O_390,N_14948,N_14717);
or UO_391 (O_391,N_14521,N_14913);
nand UO_392 (O_392,N_14985,N_14537);
nand UO_393 (O_393,N_14796,N_14946);
or UO_394 (O_394,N_14896,N_14638);
nor UO_395 (O_395,N_14705,N_14594);
and UO_396 (O_396,N_14550,N_14921);
and UO_397 (O_397,N_14745,N_14960);
xnor UO_398 (O_398,N_14933,N_14601);
and UO_399 (O_399,N_14541,N_14809);
nand UO_400 (O_400,N_14615,N_14957);
or UO_401 (O_401,N_14923,N_14746);
nor UO_402 (O_402,N_14639,N_14543);
nand UO_403 (O_403,N_14563,N_14738);
nor UO_404 (O_404,N_14591,N_14584);
nor UO_405 (O_405,N_14848,N_14571);
and UO_406 (O_406,N_14780,N_14816);
and UO_407 (O_407,N_14961,N_14893);
or UO_408 (O_408,N_14744,N_14719);
xor UO_409 (O_409,N_14675,N_14718);
nor UO_410 (O_410,N_14986,N_14872);
nand UO_411 (O_411,N_14996,N_14915);
and UO_412 (O_412,N_14535,N_14763);
xnor UO_413 (O_413,N_14790,N_14875);
nor UO_414 (O_414,N_14519,N_14608);
and UO_415 (O_415,N_14772,N_14724);
or UO_416 (O_416,N_14697,N_14650);
xnor UO_417 (O_417,N_14978,N_14600);
and UO_418 (O_418,N_14970,N_14825);
or UO_419 (O_419,N_14586,N_14647);
nor UO_420 (O_420,N_14625,N_14952);
nor UO_421 (O_421,N_14865,N_14664);
nand UO_422 (O_422,N_14698,N_14807);
xor UO_423 (O_423,N_14548,N_14877);
xnor UO_424 (O_424,N_14880,N_14582);
nor UO_425 (O_425,N_14935,N_14985);
and UO_426 (O_426,N_14955,N_14683);
xor UO_427 (O_427,N_14787,N_14627);
and UO_428 (O_428,N_14807,N_14736);
nand UO_429 (O_429,N_14577,N_14858);
nor UO_430 (O_430,N_14806,N_14746);
nor UO_431 (O_431,N_14988,N_14806);
and UO_432 (O_432,N_14881,N_14975);
xor UO_433 (O_433,N_14599,N_14525);
or UO_434 (O_434,N_14600,N_14787);
and UO_435 (O_435,N_14765,N_14959);
and UO_436 (O_436,N_14559,N_14864);
and UO_437 (O_437,N_14614,N_14928);
xnor UO_438 (O_438,N_14659,N_14622);
xnor UO_439 (O_439,N_14706,N_14786);
nor UO_440 (O_440,N_14905,N_14554);
nor UO_441 (O_441,N_14667,N_14882);
or UO_442 (O_442,N_14813,N_14922);
or UO_443 (O_443,N_14825,N_14840);
nand UO_444 (O_444,N_14746,N_14695);
or UO_445 (O_445,N_14549,N_14917);
or UO_446 (O_446,N_14759,N_14618);
xnor UO_447 (O_447,N_14645,N_14872);
nand UO_448 (O_448,N_14683,N_14819);
xor UO_449 (O_449,N_14836,N_14632);
and UO_450 (O_450,N_14697,N_14738);
or UO_451 (O_451,N_14786,N_14992);
nand UO_452 (O_452,N_14598,N_14661);
nand UO_453 (O_453,N_14600,N_14586);
nor UO_454 (O_454,N_14939,N_14566);
and UO_455 (O_455,N_14793,N_14914);
and UO_456 (O_456,N_14633,N_14529);
xnor UO_457 (O_457,N_14926,N_14587);
or UO_458 (O_458,N_14515,N_14521);
and UO_459 (O_459,N_14806,N_14639);
or UO_460 (O_460,N_14761,N_14654);
and UO_461 (O_461,N_14730,N_14621);
nor UO_462 (O_462,N_14714,N_14692);
and UO_463 (O_463,N_14808,N_14680);
or UO_464 (O_464,N_14856,N_14761);
or UO_465 (O_465,N_14819,N_14901);
xor UO_466 (O_466,N_14967,N_14849);
or UO_467 (O_467,N_14567,N_14687);
xor UO_468 (O_468,N_14976,N_14604);
and UO_469 (O_469,N_14519,N_14755);
nand UO_470 (O_470,N_14779,N_14726);
and UO_471 (O_471,N_14603,N_14739);
nand UO_472 (O_472,N_14798,N_14712);
nor UO_473 (O_473,N_14944,N_14945);
nand UO_474 (O_474,N_14962,N_14733);
and UO_475 (O_475,N_14758,N_14584);
xnor UO_476 (O_476,N_14681,N_14939);
or UO_477 (O_477,N_14845,N_14767);
nor UO_478 (O_478,N_14762,N_14687);
nand UO_479 (O_479,N_14855,N_14787);
or UO_480 (O_480,N_14720,N_14516);
and UO_481 (O_481,N_14854,N_14860);
nand UO_482 (O_482,N_14626,N_14890);
nand UO_483 (O_483,N_14799,N_14874);
or UO_484 (O_484,N_14966,N_14802);
or UO_485 (O_485,N_14583,N_14949);
nor UO_486 (O_486,N_14517,N_14903);
or UO_487 (O_487,N_14876,N_14896);
nor UO_488 (O_488,N_14802,N_14605);
and UO_489 (O_489,N_14762,N_14976);
xnor UO_490 (O_490,N_14708,N_14597);
or UO_491 (O_491,N_14907,N_14715);
xor UO_492 (O_492,N_14802,N_14654);
and UO_493 (O_493,N_14775,N_14518);
xor UO_494 (O_494,N_14907,N_14675);
xnor UO_495 (O_495,N_14783,N_14611);
and UO_496 (O_496,N_14734,N_14583);
xor UO_497 (O_497,N_14679,N_14801);
and UO_498 (O_498,N_14930,N_14938);
and UO_499 (O_499,N_14695,N_14722);
xnor UO_500 (O_500,N_14933,N_14900);
or UO_501 (O_501,N_14816,N_14899);
nand UO_502 (O_502,N_14911,N_14928);
xor UO_503 (O_503,N_14855,N_14686);
nand UO_504 (O_504,N_14964,N_14621);
or UO_505 (O_505,N_14514,N_14667);
and UO_506 (O_506,N_14745,N_14838);
nand UO_507 (O_507,N_14779,N_14778);
nor UO_508 (O_508,N_14561,N_14567);
and UO_509 (O_509,N_14514,N_14973);
nor UO_510 (O_510,N_14537,N_14679);
xnor UO_511 (O_511,N_14947,N_14850);
nand UO_512 (O_512,N_14519,N_14913);
or UO_513 (O_513,N_14745,N_14822);
or UO_514 (O_514,N_14582,N_14896);
nor UO_515 (O_515,N_14557,N_14798);
nand UO_516 (O_516,N_14663,N_14933);
nand UO_517 (O_517,N_14803,N_14524);
nand UO_518 (O_518,N_14752,N_14642);
or UO_519 (O_519,N_14960,N_14717);
nor UO_520 (O_520,N_14886,N_14929);
and UO_521 (O_521,N_14657,N_14729);
or UO_522 (O_522,N_14587,N_14762);
or UO_523 (O_523,N_14928,N_14594);
or UO_524 (O_524,N_14745,N_14525);
nand UO_525 (O_525,N_14542,N_14554);
and UO_526 (O_526,N_14708,N_14768);
nand UO_527 (O_527,N_14590,N_14652);
xnor UO_528 (O_528,N_14965,N_14558);
nor UO_529 (O_529,N_14567,N_14683);
and UO_530 (O_530,N_14943,N_14636);
nand UO_531 (O_531,N_14921,N_14757);
nor UO_532 (O_532,N_14649,N_14758);
nand UO_533 (O_533,N_14956,N_14946);
nand UO_534 (O_534,N_14996,N_14631);
and UO_535 (O_535,N_14893,N_14941);
nor UO_536 (O_536,N_14750,N_14983);
xor UO_537 (O_537,N_14699,N_14978);
or UO_538 (O_538,N_14895,N_14956);
xor UO_539 (O_539,N_14671,N_14927);
and UO_540 (O_540,N_14592,N_14812);
nor UO_541 (O_541,N_14955,N_14612);
and UO_542 (O_542,N_14650,N_14981);
and UO_543 (O_543,N_14737,N_14596);
nand UO_544 (O_544,N_14685,N_14846);
nand UO_545 (O_545,N_14609,N_14632);
nor UO_546 (O_546,N_14986,N_14629);
or UO_547 (O_547,N_14783,N_14980);
or UO_548 (O_548,N_14771,N_14804);
or UO_549 (O_549,N_14896,N_14770);
xnor UO_550 (O_550,N_14870,N_14587);
nor UO_551 (O_551,N_14546,N_14986);
nor UO_552 (O_552,N_14998,N_14605);
nand UO_553 (O_553,N_14502,N_14606);
xor UO_554 (O_554,N_14666,N_14724);
nor UO_555 (O_555,N_14827,N_14958);
xnor UO_556 (O_556,N_14682,N_14802);
nand UO_557 (O_557,N_14607,N_14601);
or UO_558 (O_558,N_14560,N_14932);
or UO_559 (O_559,N_14980,N_14964);
or UO_560 (O_560,N_14956,N_14992);
nor UO_561 (O_561,N_14798,N_14522);
and UO_562 (O_562,N_14592,N_14568);
and UO_563 (O_563,N_14908,N_14927);
nand UO_564 (O_564,N_14722,N_14793);
nand UO_565 (O_565,N_14608,N_14857);
and UO_566 (O_566,N_14511,N_14900);
or UO_567 (O_567,N_14775,N_14703);
nor UO_568 (O_568,N_14752,N_14690);
xnor UO_569 (O_569,N_14670,N_14918);
or UO_570 (O_570,N_14896,N_14800);
xor UO_571 (O_571,N_14953,N_14823);
or UO_572 (O_572,N_14800,N_14986);
nand UO_573 (O_573,N_14644,N_14945);
and UO_574 (O_574,N_14800,N_14812);
nor UO_575 (O_575,N_14792,N_14852);
nand UO_576 (O_576,N_14726,N_14609);
and UO_577 (O_577,N_14547,N_14758);
nor UO_578 (O_578,N_14549,N_14860);
and UO_579 (O_579,N_14518,N_14710);
nand UO_580 (O_580,N_14791,N_14687);
nand UO_581 (O_581,N_14814,N_14542);
xnor UO_582 (O_582,N_14975,N_14869);
nand UO_583 (O_583,N_14953,N_14655);
and UO_584 (O_584,N_14852,N_14800);
nand UO_585 (O_585,N_14722,N_14772);
and UO_586 (O_586,N_14776,N_14600);
or UO_587 (O_587,N_14881,N_14541);
nor UO_588 (O_588,N_14799,N_14751);
or UO_589 (O_589,N_14620,N_14517);
and UO_590 (O_590,N_14642,N_14644);
xor UO_591 (O_591,N_14778,N_14814);
xor UO_592 (O_592,N_14656,N_14984);
xnor UO_593 (O_593,N_14731,N_14611);
xor UO_594 (O_594,N_14923,N_14533);
nand UO_595 (O_595,N_14898,N_14814);
and UO_596 (O_596,N_14810,N_14680);
and UO_597 (O_597,N_14545,N_14932);
or UO_598 (O_598,N_14812,N_14672);
nor UO_599 (O_599,N_14555,N_14904);
nor UO_600 (O_600,N_14583,N_14548);
nor UO_601 (O_601,N_14512,N_14987);
or UO_602 (O_602,N_14840,N_14855);
and UO_603 (O_603,N_14940,N_14777);
and UO_604 (O_604,N_14979,N_14936);
or UO_605 (O_605,N_14956,N_14858);
nor UO_606 (O_606,N_14849,N_14685);
nand UO_607 (O_607,N_14870,N_14693);
and UO_608 (O_608,N_14718,N_14533);
nand UO_609 (O_609,N_14669,N_14681);
and UO_610 (O_610,N_14863,N_14703);
xor UO_611 (O_611,N_14844,N_14502);
and UO_612 (O_612,N_14857,N_14933);
and UO_613 (O_613,N_14725,N_14920);
xnor UO_614 (O_614,N_14741,N_14857);
xor UO_615 (O_615,N_14672,N_14757);
nor UO_616 (O_616,N_14638,N_14895);
or UO_617 (O_617,N_14503,N_14776);
nor UO_618 (O_618,N_14561,N_14955);
or UO_619 (O_619,N_14517,N_14967);
and UO_620 (O_620,N_14904,N_14719);
and UO_621 (O_621,N_14955,N_14652);
xor UO_622 (O_622,N_14608,N_14830);
nand UO_623 (O_623,N_14837,N_14504);
and UO_624 (O_624,N_14683,N_14544);
and UO_625 (O_625,N_14606,N_14993);
nor UO_626 (O_626,N_14615,N_14681);
or UO_627 (O_627,N_14986,N_14514);
and UO_628 (O_628,N_14548,N_14571);
nor UO_629 (O_629,N_14900,N_14791);
nor UO_630 (O_630,N_14555,N_14709);
nor UO_631 (O_631,N_14627,N_14511);
nor UO_632 (O_632,N_14571,N_14695);
nand UO_633 (O_633,N_14785,N_14601);
and UO_634 (O_634,N_14978,N_14861);
and UO_635 (O_635,N_14956,N_14923);
nor UO_636 (O_636,N_14748,N_14963);
nand UO_637 (O_637,N_14847,N_14635);
and UO_638 (O_638,N_14512,N_14728);
xnor UO_639 (O_639,N_14850,N_14812);
and UO_640 (O_640,N_14874,N_14886);
or UO_641 (O_641,N_14603,N_14732);
or UO_642 (O_642,N_14908,N_14587);
and UO_643 (O_643,N_14727,N_14824);
or UO_644 (O_644,N_14552,N_14967);
or UO_645 (O_645,N_14566,N_14730);
or UO_646 (O_646,N_14824,N_14869);
or UO_647 (O_647,N_14979,N_14720);
xnor UO_648 (O_648,N_14817,N_14642);
nand UO_649 (O_649,N_14604,N_14971);
nand UO_650 (O_650,N_14597,N_14617);
or UO_651 (O_651,N_14528,N_14506);
or UO_652 (O_652,N_14951,N_14757);
and UO_653 (O_653,N_14882,N_14780);
or UO_654 (O_654,N_14761,N_14764);
nand UO_655 (O_655,N_14934,N_14649);
and UO_656 (O_656,N_14536,N_14943);
xnor UO_657 (O_657,N_14730,N_14701);
nor UO_658 (O_658,N_14628,N_14530);
nand UO_659 (O_659,N_14957,N_14574);
and UO_660 (O_660,N_14535,N_14892);
xor UO_661 (O_661,N_14676,N_14746);
xnor UO_662 (O_662,N_14506,N_14745);
and UO_663 (O_663,N_14581,N_14804);
xor UO_664 (O_664,N_14977,N_14868);
xnor UO_665 (O_665,N_14601,N_14896);
and UO_666 (O_666,N_14682,N_14649);
nor UO_667 (O_667,N_14928,N_14973);
and UO_668 (O_668,N_14737,N_14764);
and UO_669 (O_669,N_14922,N_14544);
and UO_670 (O_670,N_14530,N_14827);
nor UO_671 (O_671,N_14701,N_14975);
xnor UO_672 (O_672,N_14849,N_14837);
and UO_673 (O_673,N_14907,N_14731);
or UO_674 (O_674,N_14716,N_14721);
xnor UO_675 (O_675,N_14807,N_14971);
nand UO_676 (O_676,N_14883,N_14519);
or UO_677 (O_677,N_14917,N_14841);
nor UO_678 (O_678,N_14756,N_14718);
and UO_679 (O_679,N_14905,N_14859);
xnor UO_680 (O_680,N_14946,N_14945);
nand UO_681 (O_681,N_14829,N_14689);
nor UO_682 (O_682,N_14820,N_14773);
or UO_683 (O_683,N_14574,N_14974);
or UO_684 (O_684,N_14885,N_14750);
and UO_685 (O_685,N_14610,N_14989);
nor UO_686 (O_686,N_14546,N_14702);
and UO_687 (O_687,N_14590,N_14691);
nand UO_688 (O_688,N_14969,N_14938);
nand UO_689 (O_689,N_14552,N_14949);
nor UO_690 (O_690,N_14889,N_14560);
or UO_691 (O_691,N_14811,N_14513);
xnor UO_692 (O_692,N_14881,N_14859);
or UO_693 (O_693,N_14687,N_14926);
xnor UO_694 (O_694,N_14510,N_14561);
or UO_695 (O_695,N_14539,N_14767);
xnor UO_696 (O_696,N_14749,N_14764);
or UO_697 (O_697,N_14868,N_14530);
and UO_698 (O_698,N_14655,N_14762);
nand UO_699 (O_699,N_14880,N_14859);
xnor UO_700 (O_700,N_14659,N_14529);
nand UO_701 (O_701,N_14519,N_14773);
nor UO_702 (O_702,N_14542,N_14622);
nand UO_703 (O_703,N_14663,N_14977);
and UO_704 (O_704,N_14757,N_14815);
nor UO_705 (O_705,N_14541,N_14922);
nand UO_706 (O_706,N_14878,N_14955);
and UO_707 (O_707,N_14888,N_14866);
and UO_708 (O_708,N_14843,N_14964);
nor UO_709 (O_709,N_14518,N_14834);
xnor UO_710 (O_710,N_14563,N_14702);
xnor UO_711 (O_711,N_14629,N_14537);
or UO_712 (O_712,N_14634,N_14760);
or UO_713 (O_713,N_14868,N_14748);
nand UO_714 (O_714,N_14787,N_14998);
nand UO_715 (O_715,N_14794,N_14636);
xor UO_716 (O_716,N_14608,N_14612);
nor UO_717 (O_717,N_14979,N_14955);
and UO_718 (O_718,N_14741,N_14944);
xnor UO_719 (O_719,N_14616,N_14815);
or UO_720 (O_720,N_14980,N_14592);
nor UO_721 (O_721,N_14935,N_14635);
nand UO_722 (O_722,N_14690,N_14991);
or UO_723 (O_723,N_14815,N_14989);
or UO_724 (O_724,N_14653,N_14694);
nand UO_725 (O_725,N_14879,N_14707);
and UO_726 (O_726,N_14928,N_14974);
nor UO_727 (O_727,N_14842,N_14588);
nand UO_728 (O_728,N_14867,N_14816);
nor UO_729 (O_729,N_14688,N_14986);
or UO_730 (O_730,N_14615,N_14695);
or UO_731 (O_731,N_14644,N_14791);
and UO_732 (O_732,N_14554,N_14887);
and UO_733 (O_733,N_14619,N_14876);
xnor UO_734 (O_734,N_14840,N_14995);
and UO_735 (O_735,N_14819,N_14570);
or UO_736 (O_736,N_14504,N_14913);
xor UO_737 (O_737,N_14787,N_14961);
nand UO_738 (O_738,N_14697,N_14612);
or UO_739 (O_739,N_14841,N_14671);
or UO_740 (O_740,N_14835,N_14874);
nand UO_741 (O_741,N_14848,N_14825);
nand UO_742 (O_742,N_14848,N_14706);
nand UO_743 (O_743,N_14887,N_14526);
nand UO_744 (O_744,N_14661,N_14969);
and UO_745 (O_745,N_14998,N_14567);
nand UO_746 (O_746,N_14630,N_14607);
and UO_747 (O_747,N_14883,N_14880);
or UO_748 (O_748,N_14635,N_14630);
xor UO_749 (O_749,N_14969,N_14886);
nand UO_750 (O_750,N_14856,N_14901);
xnor UO_751 (O_751,N_14877,N_14746);
nor UO_752 (O_752,N_14654,N_14806);
nand UO_753 (O_753,N_14661,N_14826);
xnor UO_754 (O_754,N_14583,N_14805);
xnor UO_755 (O_755,N_14863,N_14765);
nor UO_756 (O_756,N_14936,N_14530);
nand UO_757 (O_757,N_14680,N_14801);
nand UO_758 (O_758,N_14544,N_14582);
xnor UO_759 (O_759,N_14588,N_14694);
and UO_760 (O_760,N_14984,N_14968);
or UO_761 (O_761,N_14509,N_14985);
nand UO_762 (O_762,N_14724,N_14828);
nor UO_763 (O_763,N_14596,N_14829);
xor UO_764 (O_764,N_14726,N_14630);
xor UO_765 (O_765,N_14636,N_14722);
nor UO_766 (O_766,N_14772,N_14841);
nor UO_767 (O_767,N_14796,N_14647);
xor UO_768 (O_768,N_14771,N_14732);
nand UO_769 (O_769,N_14860,N_14742);
or UO_770 (O_770,N_14567,N_14806);
xnor UO_771 (O_771,N_14786,N_14619);
or UO_772 (O_772,N_14745,N_14986);
nor UO_773 (O_773,N_14787,N_14548);
or UO_774 (O_774,N_14914,N_14569);
nor UO_775 (O_775,N_14650,N_14557);
nor UO_776 (O_776,N_14638,N_14604);
nor UO_777 (O_777,N_14565,N_14516);
or UO_778 (O_778,N_14935,N_14764);
or UO_779 (O_779,N_14522,N_14525);
nand UO_780 (O_780,N_14703,N_14704);
or UO_781 (O_781,N_14587,N_14548);
xnor UO_782 (O_782,N_14593,N_14760);
or UO_783 (O_783,N_14810,N_14641);
xnor UO_784 (O_784,N_14546,N_14600);
or UO_785 (O_785,N_14554,N_14587);
nand UO_786 (O_786,N_14933,N_14607);
nor UO_787 (O_787,N_14915,N_14969);
nand UO_788 (O_788,N_14805,N_14596);
nor UO_789 (O_789,N_14844,N_14604);
nor UO_790 (O_790,N_14981,N_14759);
nor UO_791 (O_791,N_14771,N_14623);
nand UO_792 (O_792,N_14596,N_14848);
xnor UO_793 (O_793,N_14713,N_14592);
and UO_794 (O_794,N_14785,N_14678);
or UO_795 (O_795,N_14706,N_14505);
nand UO_796 (O_796,N_14608,N_14960);
and UO_797 (O_797,N_14570,N_14655);
xnor UO_798 (O_798,N_14729,N_14716);
nand UO_799 (O_799,N_14773,N_14957);
nand UO_800 (O_800,N_14766,N_14588);
or UO_801 (O_801,N_14820,N_14607);
nor UO_802 (O_802,N_14519,N_14847);
and UO_803 (O_803,N_14626,N_14522);
nor UO_804 (O_804,N_14674,N_14928);
or UO_805 (O_805,N_14828,N_14617);
nor UO_806 (O_806,N_14634,N_14785);
and UO_807 (O_807,N_14601,N_14901);
nor UO_808 (O_808,N_14763,N_14803);
and UO_809 (O_809,N_14799,N_14779);
xnor UO_810 (O_810,N_14546,N_14893);
and UO_811 (O_811,N_14893,N_14760);
or UO_812 (O_812,N_14685,N_14576);
and UO_813 (O_813,N_14574,N_14830);
xor UO_814 (O_814,N_14735,N_14528);
or UO_815 (O_815,N_14575,N_14744);
nand UO_816 (O_816,N_14516,N_14658);
nand UO_817 (O_817,N_14939,N_14942);
nand UO_818 (O_818,N_14671,N_14709);
or UO_819 (O_819,N_14572,N_14726);
xor UO_820 (O_820,N_14795,N_14904);
nor UO_821 (O_821,N_14574,N_14893);
or UO_822 (O_822,N_14955,N_14842);
xnor UO_823 (O_823,N_14598,N_14957);
and UO_824 (O_824,N_14720,N_14702);
and UO_825 (O_825,N_14897,N_14929);
nand UO_826 (O_826,N_14919,N_14649);
xnor UO_827 (O_827,N_14681,N_14524);
xnor UO_828 (O_828,N_14764,N_14836);
nand UO_829 (O_829,N_14991,N_14595);
nor UO_830 (O_830,N_14573,N_14764);
or UO_831 (O_831,N_14621,N_14501);
nand UO_832 (O_832,N_14686,N_14798);
and UO_833 (O_833,N_14590,N_14536);
nand UO_834 (O_834,N_14837,N_14502);
and UO_835 (O_835,N_14531,N_14735);
nor UO_836 (O_836,N_14996,N_14568);
or UO_837 (O_837,N_14637,N_14991);
nand UO_838 (O_838,N_14672,N_14621);
or UO_839 (O_839,N_14637,N_14718);
or UO_840 (O_840,N_14572,N_14835);
nand UO_841 (O_841,N_14890,N_14547);
or UO_842 (O_842,N_14612,N_14935);
nor UO_843 (O_843,N_14579,N_14515);
xor UO_844 (O_844,N_14874,N_14682);
nand UO_845 (O_845,N_14789,N_14581);
and UO_846 (O_846,N_14854,N_14659);
nand UO_847 (O_847,N_14824,N_14557);
nand UO_848 (O_848,N_14625,N_14723);
nor UO_849 (O_849,N_14639,N_14500);
or UO_850 (O_850,N_14629,N_14753);
xor UO_851 (O_851,N_14935,N_14932);
or UO_852 (O_852,N_14646,N_14532);
nand UO_853 (O_853,N_14605,N_14655);
nand UO_854 (O_854,N_14816,N_14594);
and UO_855 (O_855,N_14611,N_14793);
xor UO_856 (O_856,N_14539,N_14631);
nor UO_857 (O_857,N_14784,N_14863);
nand UO_858 (O_858,N_14548,N_14748);
or UO_859 (O_859,N_14700,N_14614);
or UO_860 (O_860,N_14867,N_14865);
and UO_861 (O_861,N_14682,N_14702);
xnor UO_862 (O_862,N_14570,N_14805);
or UO_863 (O_863,N_14744,N_14848);
xnor UO_864 (O_864,N_14840,N_14912);
or UO_865 (O_865,N_14751,N_14733);
nand UO_866 (O_866,N_14776,N_14698);
or UO_867 (O_867,N_14801,N_14857);
nor UO_868 (O_868,N_14782,N_14649);
xnor UO_869 (O_869,N_14822,N_14726);
and UO_870 (O_870,N_14657,N_14970);
nand UO_871 (O_871,N_14931,N_14684);
xnor UO_872 (O_872,N_14744,N_14958);
nand UO_873 (O_873,N_14579,N_14975);
xnor UO_874 (O_874,N_14669,N_14689);
nand UO_875 (O_875,N_14884,N_14922);
nor UO_876 (O_876,N_14969,N_14747);
nand UO_877 (O_877,N_14973,N_14513);
and UO_878 (O_878,N_14921,N_14742);
or UO_879 (O_879,N_14562,N_14529);
xor UO_880 (O_880,N_14716,N_14877);
xnor UO_881 (O_881,N_14902,N_14782);
nand UO_882 (O_882,N_14586,N_14704);
and UO_883 (O_883,N_14979,N_14697);
and UO_884 (O_884,N_14798,N_14637);
nor UO_885 (O_885,N_14573,N_14837);
xnor UO_886 (O_886,N_14795,N_14640);
or UO_887 (O_887,N_14882,N_14751);
or UO_888 (O_888,N_14864,N_14807);
nand UO_889 (O_889,N_14669,N_14988);
nor UO_890 (O_890,N_14900,N_14950);
nand UO_891 (O_891,N_14874,N_14944);
and UO_892 (O_892,N_14724,N_14978);
and UO_893 (O_893,N_14640,N_14884);
nand UO_894 (O_894,N_14861,N_14822);
nor UO_895 (O_895,N_14832,N_14773);
or UO_896 (O_896,N_14540,N_14845);
or UO_897 (O_897,N_14959,N_14654);
or UO_898 (O_898,N_14558,N_14831);
xnor UO_899 (O_899,N_14964,N_14973);
or UO_900 (O_900,N_14629,N_14605);
nor UO_901 (O_901,N_14735,N_14583);
nor UO_902 (O_902,N_14848,N_14954);
or UO_903 (O_903,N_14576,N_14990);
nor UO_904 (O_904,N_14727,N_14938);
nand UO_905 (O_905,N_14623,N_14718);
xor UO_906 (O_906,N_14540,N_14878);
nand UO_907 (O_907,N_14674,N_14832);
and UO_908 (O_908,N_14604,N_14566);
or UO_909 (O_909,N_14922,N_14750);
xor UO_910 (O_910,N_14712,N_14622);
or UO_911 (O_911,N_14842,N_14911);
nor UO_912 (O_912,N_14604,N_14599);
or UO_913 (O_913,N_14609,N_14657);
xnor UO_914 (O_914,N_14542,N_14534);
and UO_915 (O_915,N_14648,N_14770);
nor UO_916 (O_916,N_14648,N_14671);
xnor UO_917 (O_917,N_14735,N_14519);
xnor UO_918 (O_918,N_14626,N_14707);
nor UO_919 (O_919,N_14661,N_14641);
nor UO_920 (O_920,N_14730,N_14740);
nand UO_921 (O_921,N_14836,N_14866);
or UO_922 (O_922,N_14515,N_14667);
and UO_923 (O_923,N_14771,N_14871);
and UO_924 (O_924,N_14863,N_14590);
nand UO_925 (O_925,N_14718,N_14951);
and UO_926 (O_926,N_14611,N_14721);
nand UO_927 (O_927,N_14555,N_14888);
xnor UO_928 (O_928,N_14822,N_14619);
nor UO_929 (O_929,N_14741,N_14544);
or UO_930 (O_930,N_14918,N_14708);
nor UO_931 (O_931,N_14724,N_14618);
nand UO_932 (O_932,N_14556,N_14741);
xnor UO_933 (O_933,N_14553,N_14607);
nor UO_934 (O_934,N_14927,N_14811);
and UO_935 (O_935,N_14799,N_14755);
and UO_936 (O_936,N_14686,N_14935);
nand UO_937 (O_937,N_14632,N_14637);
xnor UO_938 (O_938,N_14725,N_14601);
xor UO_939 (O_939,N_14907,N_14504);
nand UO_940 (O_940,N_14605,N_14892);
nand UO_941 (O_941,N_14998,N_14598);
nand UO_942 (O_942,N_14712,N_14543);
nor UO_943 (O_943,N_14979,N_14500);
nand UO_944 (O_944,N_14892,N_14569);
and UO_945 (O_945,N_14956,N_14947);
nor UO_946 (O_946,N_14991,N_14797);
nand UO_947 (O_947,N_14714,N_14511);
nor UO_948 (O_948,N_14535,N_14664);
nand UO_949 (O_949,N_14597,N_14626);
nand UO_950 (O_950,N_14751,N_14570);
nand UO_951 (O_951,N_14529,N_14892);
nand UO_952 (O_952,N_14733,N_14609);
or UO_953 (O_953,N_14841,N_14531);
nand UO_954 (O_954,N_14986,N_14767);
and UO_955 (O_955,N_14690,N_14932);
or UO_956 (O_956,N_14874,N_14543);
or UO_957 (O_957,N_14961,N_14820);
nor UO_958 (O_958,N_14761,N_14775);
nand UO_959 (O_959,N_14621,N_14564);
or UO_960 (O_960,N_14985,N_14551);
nand UO_961 (O_961,N_14966,N_14928);
or UO_962 (O_962,N_14555,N_14788);
nand UO_963 (O_963,N_14697,N_14730);
and UO_964 (O_964,N_14868,N_14591);
and UO_965 (O_965,N_14843,N_14935);
or UO_966 (O_966,N_14987,N_14866);
xnor UO_967 (O_967,N_14909,N_14761);
nand UO_968 (O_968,N_14888,N_14539);
nand UO_969 (O_969,N_14501,N_14947);
xor UO_970 (O_970,N_14636,N_14701);
xnor UO_971 (O_971,N_14956,N_14613);
or UO_972 (O_972,N_14795,N_14575);
nor UO_973 (O_973,N_14999,N_14788);
xor UO_974 (O_974,N_14949,N_14541);
nand UO_975 (O_975,N_14763,N_14890);
nor UO_976 (O_976,N_14729,N_14853);
or UO_977 (O_977,N_14840,N_14946);
xor UO_978 (O_978,N_14758,N_14731);
nor UO_979 (O_979,N_14657,N_14560);
or UO_980 (O_980,N_14972,N_14765);
nand UO_981 (O_981,N_14835,N_14595);
and UO_982 (O_982,N_14503,N_14778);
xnor UO_983 (O_983,N_14943,N_14875);
xor UO_984 (O_984,N_14621,N_14622);
and UO_985 (O_985,N_14918,N_14768);
nand UO_986 (O_986,N_14573,N_14686);
nor UO_987 (O_987,N_14556,N_14883);
and UO_988 (O_988,N_14540,N_14784);
nor UO_989 (O_989,N_14693,N_14924);
nor UO_990 (O_990,N_14989,N_14727);
nor UO_991 (O_991,N_14983,N_14989);
and UO_992 (O_992,N_14946,N_14611);
or UO_993 (O_993,N_14588,N_14729);
xnor UO_994 (O_994,N_14556,N_14757);
and UO_995 (O_995,N_14721,N_14898);
or UO_996 (O_996,N_14776,N_14778);
xor UO_997 (O_997,N_14685,N_14757);
nor UO_998 (O_998,N_14670,N_14993);
nor UO_999 (O_999,N_14585,N_14700);
nand UO_1000 (O_1000,N_14896,N_14894);
nor UO_1001 (O_1001,N_14671,N_14730);
nand UO_1002 (O_1002,N_14562,N_14750);
or UO_1003 (O_1003,N_14668,N_14673);
nand UO_1004 (O_1004,N_14986,N_14865);
or UO_1005 (O_1005,N_14585,N_14847);
nand UO_1006 (O_1006,N_14694,N_14971);
nand UO_1007 (O_1007,N_14875,N_14987);
or UO_1008 (O_1008,N_14535,N_14607);
or UO_1009 (O_1009,N_14923,N_14667);
or UO_1010 (O_1010,N_14517,N_14558);
nor UO_1011 (O_1011,N_14855,N_14713);
or UO_1012 (O_1012,N_14620,N_14626);
nand UO_1013 (O_1013,N_14966,N_14883);
nor UO_1014 (O_1014,N_14753,N_14587);
xor UO_1015 (O_1015,N_14529,N_14912);
and UO_1016 (O_1016,N_14680,N_14838);
and UO_1017 (O_1017,N_14669,N_14836);
and UO_1018 (O_1018,N_14520,N_14505);
nand UO_1019 (O_1019,N_14915,N_14793);
xor UO_1020 (O_1020,N_14976,N_14818);
or UO_1021 (O_1021,N_14553,N_14647);
nor UO_1022 (O_1022,N_14521,N_14755);
xor UO_1023 (O_1023,N_14922,N_14836);
or UO_1024 (O_1024,N_14829,N_14787);
nor UO_1025 (O_1025,N_14514,N_14549);
xnor UO_1026 (O_1026,N_14783,N_14856);
nor UO_1027 (O_1027,N_14525,N_14649);
nor UO_1028 (O_1028,N_14501,N_14739);
or UO_1029 (O_1029,N_14652,N_14657);
nor UO_1030 (O_1030,N_14613,N_14765);
nand UO_1031 (O_1031,N_14805,N_14959);
and UO_1032 (O_1032,N_14763,N_14595);
or UO_1033 (O_1033,N_14549,N_14703);
nand UO_1034 (O_1034,N_14801,N_14991);
xor UO_1035 (O_1035,N_14534,N_14676);
nor UO_1036 (O_1036,N_14832,N_14600);
or UO_1037 (O_1037,N_14962,N_14774);
xnor UO_1038 (O_1038,N_14591,N_14927);
nand UO_1039 (O_1039,N_14661,N_14769);
and UO_1040 (O_1040,N_14929,N_14529);
xor UO_1041 (O_1041,N_14564,N_14925);
nand UO_1042 (O_1042,N_14572,N_14682);
nor UO_1043 (O_1043,N_14876,N_14565);
xor UO_1044 (O_1044,N_14936,N_14902);
nor UO_1045 (O_1045,N_14869,N_14803);
and UO_1046 (O_1046,N_14818,N_14664);
xor UO_1047 (O_1047,N_14589,N_14562);
or UO_1048 (O_1048,N_14648,N_14726);
nor UO_1049 (O_1049,N_14959,N_14826);
nand UO_1050 (O_1050,N_14525,N_14513);
nand UO_1051 (O_1051,N_14785,N_14874);
nor UO_1052 (O_1052,N_14787,N_14996);
nand UO_1053 (O_1053,N_14993,N_14722);
or UO_1054 (O_1054,N_14571,N_14889);
and UO_1055 (O_1055,N_14919,N_14981);
nor UO_1056 (O_1056,N_14593,N_14893);
and UO_1057 (O_1057,N_14618,N_14865);
or UO_1058 (O_1058,N_14645,N_14569);
xnor UO_1059 (O_1059,N_14648,N_14948);
nand UO_1060 (O_1060,N_14708,N_14739);
nor UO_1061 (O_1061,N_14604,N_14713);
xor UO_1062 (O_1062,N_14707,N_14736);
nor UO_1063 (O_1063,N_14524,N_14909);
nor UO_1064 (O_1064,N_14926,N_14665);
nand UO_1065 (O_1065,N_14763,N_14655);
and UO_1066 (O_1066,N_14673,N_14706);
or UO_1067 (O_1067,N_14654,N_14904);
xnor UO_1068 (O_1068,N_14859,N_14522);
and UO_1069 (O_1069,N_14670,N_14640);
nand UO_1070 (O_1070,N_14818,N_14890);
or UO_1071 (O_1071,N_14809,N_14552);
or UO_1072 (O_1072,N_14775,N_14790);
nand UO_1073 (O_1073,N_14668,N_14524);
and UO_1074 (O_1074,N_14870,N_14610);
nand UO_1075 (O_1075,N_14607,N_14500);
nor UO_1076 (O_1076,N_14688,N_14606);
and UO_1077 (O_1077,N_14875,N_14717);
nor UO_1078 (O_1078,N_14673,N_14909);
or UO_1079 (O_1079,N_14618,N_14767);
or UO_1080 (O_1080,N_14843,N_14852);
or UO_1081 (O_1081,N_14967,N_14756);
nand UO_1082 (O_1082,N_14782,N_14984);
nand UO_1083 (O_1083,N_14628,N_14927);
nand UO_1084 (O_1084,N_14797,N_14626);
and UO_1085 (O_1085,N_14741,N_14520);
or UO_1086 (O_1086,N_14908,N_14732);
and UO_1087 (O_1087,N_14835,N_14873);
or UO_1088 (O_1088,N_14868,N_14653);
xor UO_1089 (O_1089,N_14946,N_14507);
xor UO_1090 (O_1090,N_14625,N_14910);
nand UO_1091 (O_1091,N_14691,N_14957);
nor UO_1092 (O_1092,N_14926,N_14951);
or UO_1093 (O_1093,N_14970,N_14800);
and UO_1094 (O_1094,N_14619,N_14568);
nand UO_1095 (O_1095,N_14731,N_14693);
nand UO_1096 (O_1096,N_14553,N_14515);
and UO_1097 (O_1097,N_14540,N_14694);
or UO_1098 (O_1098,N_14713,N_14695);
xor UO_1099 (O_1099,N_14826,N_14729);
nand UO_1100 (O_1100,N_14968,N_14704);
nand UO_1101 (O_1101,N_14630,N_14659);
or UO_1102 (O_1102,N_14507,N_14579);
or UO_1103 (O_1103,N_14989,N_14638);
or UO_1104 (O_1104,N_14802,N_14689);
xor UO_1105 (O_1105,N_14602,N_14715);
or UO_1106 (O_1106,N_14918,N_14562);
nor UO_1107 (O_1107,N_14664,N_14731);
and UO_1108 (O_1108,N_14667,N_14630);
nor UO_1109 (O_1109,N_14598,N_14546);
nor UO_1110 (O_1110,N_14997,N_14926);
or UO_1111 (O_1111,N_14781,N_14731);
xor UO_1112 (O_1112,N_14587,N_14893);
and UO_1113 (O_1113,N_14538,N_14790);
xor UO_1114 (O_1114,N_14907,N_14726);
xnor UO_1115 (O_1115,N_14593,N_14789);
xnor UO_1116 (O_1116,N_14979,N_14598);
nor UO_1117 (O_1117,N_14753,N_14656);
and UO_1118 (O_1118,N_14861,N_14827);
nor UO_1119 (O_1119,N_14862,N_14896);
or UO_1120 (O_1120,N_14506,N_14504);
xnor UO_1121 (O_1121,N_14720,N_14823);
xor UO_1122 (O_1122,N_14944,N_14909);
xnor UO_1123 (O_1123,N_14886,N_14966);
xnor UO_1124 (O_1124,N_14739,N_14577);
nor UO_1125 (O_1125,N_14626,N_14581);
and UO_1126 (O_1126,N_14935,N_14813);
or UO_1127 (O_1127,N_14703,N_14694);
or UO_1128 (O_1128,N_14656,N_14953);
and UO_1129 (O_1129,N_14804,N_14649);
xor UO_1130 (O_1130,N_14637,N_14875);
xnor UO_1131 (O_1131,N_14734,N_14513);
and UO_1132 (O_1132,N_14948,N_14931);
nor UO_1133 (O_1133,N_14790,N_14527);
and UO_1134 (O_1134,N_14786,N_14546);
nor UO_1135 (O_1135,N_14728,N_14718);
nor UO_1136 (O_1136,N_14619,N_14716);
nor UO_1137 (O_1137,N_14818,N_14703);
or UO_1138 (O_1138,N_14602,N_14523);
xor UO_1139 (O_1139,N_14699,N_14622);
and UO_1140 (O_1140,N_14581,N_14651);
nand UO_1141 (O_1141,N_14847,N_14511);
nand UO_1142 (O_1142,N_14563,N_14678);
nand UO_1143 (O_1143,N_14895,N_14592);
xnor UO_1144 (O_1144,N_14563,N_14603);
xnor UO_1145 (O_1145,N_14921,N_14802);
nor UO_1146 (O_1146,N_14827,N_14637);
nor UO_1147 (O_1147,N_14748,N_14997);
nor UO_1148 (O_1148,N_14941,N_14535);
and UO_1149 (O_1149,N_14685,N_14915);
xnor UO_1150 (O_1150,N_14937,N_14687);
nand UO_1151 (O_1151,N_14670,N_14933);
or UO_1152 (O_1152,N_14862,N_14596);
xnor UO_1153 (O_1153,N_14845,N_14592);
or UO_1154 (O_1154,N_14964,N_14736);
nand UO_1155 (O_1155,N_14843,N_14771);
and UO_1156 (O_1156,N_14745,N_14788);
xnor UO_1157 (O_1157,N_14775,N_14928);
xnor UO_1158 (O_1158,N_14764,N_14628);
nand UO_1159 (O_1159,N_14865,N_14988);
or UO_1160 (O_1160,N_14940,N_14729);
nor UO_1161 (O_1161,N_14997,N_14989);
xnor UO_1162 (O_1162,N_14808,N_14571);
nand UO_1163 (O_1163,N_14788,N_14853);
xor UO_1164 (O_1164,N_14581,N_14640);
xnor UO_1165 (O_1165,N_14698,N_14782);
nand UO_1166 (O_1166,N_14631,N_14647);
or UO_1167 (O_1167,N_14558,N_14975);
and UO_1168 (O_1168,N_14886,N_14729);
xor UO_1169 (O_1169,N_14686,N_14987);
or UO_1170 (O_1170,N_14574,N_14815);
or UO_1171 (O_1171,N_14776,N_14745);
xnor UO_1172 (O_1172,N_14923,N_14535);
nor UO_1173 (O_1173,N_14783,N_14986);
and UO_1174 (O_1174,N_14952,N_14737);
xor UO_1175 (O_1175,N_14529,N_14894);
and UO_1176 (O_1176,N_14758,N_14683);
and UO_1177 (O_1177,N_14786,N_14965);
nand UO_1178 (O_1178,N_14521,N_14684);
or UO_1179 (O_1179,N_14598,N_14735);
and UO_1180 (O_1180,N_14980,N_14584);
nor UO_1181 (O_1181,N_14574,N_14891);
nand UO_1182 (O_1182,N_14645,N_14500);
or UO_1183 (O_1183,N_14865,N_14809);
nor UO_1184 (O_1184,N_14555,N_14564);
nor UO_1185 (O_1185,N_14716,N_14690);
or UO_1186 (O_1186,N_14679,N_14600);
xnor UO_1187 (O_1187,N_14928,N_14717);
or UO_1188 (O_1188,N_14975,N_14715);
xor UO_1189 (O_1189,N_14676,N_14747);
nand UO_1190 (O_1190,N_14824,N_14811);
and UO_1191 (O_1191,N_14921,N_14787);
xnor UO_1192 (O_1192,N_14940,N_14742);
nor UO_1193 (O_1193,N_14616,N_14748);
nor UO_1194 (O_1194,N_14530,N_14772);
and UO_1195 (O_1195,N_14747,N_14753);
nand UO_1196 (O_1196,N_14585,N_14895);
xnor UO_1197 (O_1197,N_14558,N_14980);
nor UO_1198 (O_1198,N_14634,N_14779);
and UO_1199 (O_1199,N_14540,N_14892);
or UO_1200 (O_1200,N_14948,N_14745);
xnor UO_1201 (O_1201,N_14854,N_14937);
xnor UO_1202 (O_1202,N_14746,N_14550);
xnor UO_1203 (O_1203,N_14523,N_14878);
nor UO_1204 (O_1204,N_14979,N_14772);
xnor UO_1205 (O_1205,N_14793,N_14584);
xnor UO_1206 (O_1206,N_14868,N_14680);
and UO_1207 (O_1207,N_14613,N_14878);
xor UO_1208 (O_1208,N_14613,N_14738);
nand UO_1209 (O_1209,N_14808,N_14839);
or UO_1210 (O_1210,N_14928,N_14759);
xor UO_1211 (O_1211,N_14510,N_14697);
nor UO_1212 (O_1212,N_14852,N_14918);
or UO_1213 (O_1213,N_14543,N_14561);
nand UO_1214 (O_1214,N_14703,N_14986);
or UO_1215 (O_1215,N_14735,N_14576);
nand UO_1216 (O_1216,N_14814,N_14610);
xor UO_1217 (O_1217,N_14833,N_14981);
nor UO_1218 (O_1218,N_14868,N_14971);
and UO_1219 (O_1219,N_14797,N_14854);
or UO_1220 (O_1220,N_14638,N_14510);
or UO_1221 (O_1221,N_14691,N_14714);
nor UO_1222 (O_1222,N_14965,N_14934);
xnor UO_1223 (O_1223,N_14656,N_14683);
nand UO_1224 (O_1224,N_14512,N_14766);
or UO_1225 (O_1225,N_14982,N_14572);
nand UO_1226 (O_1226,N_14965,N_14875);
and UO_1227 (O_1227,N_14717,N_14681);
nand UO_1228 (O_1228,N_14848,N_14912);
xnor UO_1229 (O_1229,N_14692,N_14911);
or UO_1230 (O_1230,N_14809,N_14753);
xnor UO_1231 (O_1231,N_14964,N_14610);
nand UO_1232 (O_1232,N_14596,N_14747);
xnor UO_1233 (O_1233,N_14541,N_14616);
or UO_1234 (O_1234,N_14793,N_14542);
and UO_1235 (O_1235,N_14657,N_14838);
xor UO_1236 (O_1236,N_14957,N_14705);
or UO_1237 (O_1237,N_14509,N_14946);
nand UO_1238 (O_1238,N_14590,N_14980);
nand UO_1239 (O_1239,N_14986,N_14639);
nand UO_1240 (O_1240,N_14873,N_14732);
nand UO_1241 (O_1241,N_14937,N_14981);
and UO_1242 (O_1242,N_14882,N_14787);
xnor UO_1243 (O_1243,N_14504,N_14928);
and UO_1244 (O_1244,N_14993,N_14685);
xor UO_1245 (O_1245,N_14914,N_14989);
xnor UO_1246 (O_1246,N_14839,N_14984);
and UO_1247 (O_1247,N_14537,N_14684);
nor UO_1248 (O_1248,N_14626,N_14638);
nand UO_1249 (O_1249,N_14664,N_14521);
xor UO_1250 (O_1250,N_14951,N_14970);
and UO_1251 (O_1251,N_14604,N_14660);
nand UO_1252 (O_1252,N_14519,N_14946);
or UO_1253 (O_1253,N_14530,N_14916);
nor UO_1254 (O_1254,N_14986,N_14807);
xor UO_1255 (O_1255,N_14848,N_14776);
nand UO_1256 (O_1256,N_14946,N_14534);
and UO_1257 (O_1257,N_14939,N_14836);
or UO_1258 (O_1258,N_14867,N_14858);
nand UO_1259 (O_1259,N_14649,N_14769);
or UO_1260 (O_1260,N_14603,N_14616);
and UO_1261 (O_1261,N_14845,N_14545);
and UO_1262 (O_1262,N_14966,N_14594);
and UO_1263 (O_1263,N_14829,N_14746);
xor UO_1264 (O_1264,N_14855,N_14584);
nand UO_1265 (O_1265,N_14753,N_14853);
nand UO_1266 (O_1266,N_14958,N_14942);
xor UO_1267 (O_1267,N_14862,N_14718);
nand UO_1268 (O_1268,N_14895,N_14944);
xor UO_1269 (O_1269,N_14663,N_14822);
or UO_1270 (O_1270,N_14974,N_14779);
xor UO_1271 (O_1271,N_14519,N_14517);
or UO_1272 (O_1272,N_14840,N_14980);
nand UO_1273 (O_1273,N_14732,N_14840);
nor UO_1274 (O_1274,N_14661,N_14959);
and UO_1275 (O_1275,N_14687,N_14737);
nand UO_1276 (O_1276,N_14687,N_14656);
and UO_1277 (O_1277,N_14996,N_14674);
nor UO_1278 (O_1278,N_14866,N_14539);
nand UO_1279 (O_1279,N_14843,N_14611);
and UO_1280 (O_1280,N_14966,N_14578);
nand UO_1281 (O_1281,N_14924,N_14925);
and UO_1282 (O_1282,N_14965,N_14657);
nand UO_1283 (O_1283,N_14930,N_14851);
nand UO_1284 (O_1284,N_14572,N_14843);
and UO_1285 (O_1285,N_14531,N_14981);
and UO_1286 (O_1286,N_14718,N_14573);
or UO_1287 (O_1287,N_14992,N_14506);
nand UO_1288 (O_1288,N_14994,N_14947);
xnor UO_1289 (O_1289,N_14539,N_14788);
nor UO_1290 (O_1290,N_14624,N_14505);
or UO_1291 (O_1291,N_14749,N_14831);
or UO_1292 (O_1292,N_14956,N_14538);
nor UO_1293 (O_1293,N_14522,N_14559);
xor UO_1294 (O_1294,N_14779,N_14792);
xnor UO_1295 (O_1295,N_14782,N_14596);
and UO_1296 (O_1296,N_14621,N_14811);
nand UO_1297 (O_1297,N_14954,N_14733);
xnor UO_1298 (O_1298,N_14549,N_14622);
or UO_1299 (O_1299,N_14509,N_14628);
or UO_1300 (O_1300,N_14639,N_14770);
nand UO_1301 (O_1301,N_14776,N_14819);
nand UO_1302 (O_1302,N_14639,N_14805);
and UO_1303 (O_1303,N_14636,N_14995);
nand UO_1304 (O_1304,N_14546,N_14642);
and UO_1305 (O_1305,N_14958,N_14544);
nand UO_1306 (O_1306,N_14572,N_14592);
and UO_1307 (O_1307,N_14505,N_14512);
nor UO_1308 (O_1308,N_14877,N_14715);
nand UO_1309 (O_1309,N_14568,N_14533);
xnor UO_1310 (O_1310,N_14649,N_14869);
or UO_1311 (O_1311,N_14724,N_14961);
nand UO_1312 (O_1312,N_14866,N_14719);
nand UO_1313 (O_1313,N_14716,N_14580);
or UO_1314 (O_1314,N_14512,N_14742);
and UO_1315 (O_1315,N_14783,N_14857);
nand UO_1316 (O_1316,N_14646,N_14938);
nor UO_1317 (O_1317,N_14850,N_14702);
xnor UO_1318 (O_1318,N_14625,N_14909);
or UO_1319 (O_1319,N_14935,N_14872);
nand UO_1320 (O_1320,N_14953,N_14646);
and UO_1321 (O_1321,N_14748,N_14810);
and UO_1322 (O_1322,N_14934,N_14625);
nand UO_1323 (O_1323,N_14938,N_14567);
xnor UO_1324 (O_1324,N_14616,N_14875);
or UO_1325 (O_1325,N_14753,N_14860);
nor UO_1326 (O_1326,N_14860,N_14978);
or UO_1327 (O_1327,N_14951,N_14737);
or UO_1328 (O_1328,N_14512,N_14673);
or UO_1329 (O_1329,N_14851,N_14775);
or UO_1330 (O_1330,N_14789,N_14860);
or UO_1331 (O_1331,N_14788,N_14781);
and UO_1332 (O_1332,N_14560,N_14590);
nor UO_1333 (O_1333,N_14732,N_14767);
or UO_1334 (O_1334,N_14610,N_14988);
nor UO_1335 (O_1335,N_14682,N_14997);
nor UO_1336 (O_1336,N_14513,N_14953);
nand UO_1337 (O_1337,N_14629,N_14919);
xor UO_1338 (O_1338,N_14868,N_14753);
nand UO_1339 (O_1339,N_14648,N_14804);
nor UO_1340 (O_1340,N_14749,N_14994);
nand UO_1341 (O_1341,N_14697,N_14631);
nand UO_1342 (O_1342,N_14905,N_14680);
and UO_1343 (O_1343,N_14687,N_14671);
nor UO_1344 (O_1344,N_14813,N_14769);
nor UO_1345 (O_1345,N_14753,N_14695);
nor UO_1346 (O_1346,N_14584,N_14896);
nor UO_1347 (O_1347,N_14759,N_14923);
xnor UO_1348 (O_1348,N_14648,N_14525);
nor UO_1349 (O_1349,N_14603,N_14927);
nand UO_1350 (O_1350,N_14771,N_14832);
or UO_1351 (O_1351,N_14875,N_14692);
and UO_1352 (O_1352,N_14511,N_14532);
and UO_1353 (O_1353,N_14652,N_14677);
nor UO_1354 (O_1354,N_14847,N_14986);
nand UO_1355 (O_1355,N_14995,N_14679);
and UO_1356 (O_1356,N_14926,N_14697);
or UO_1357 (O_1357,N_14608,N_14768);
xnor UO_1358 (O_1358,N_14936,N_14766);
nand UO_1359 (O_1359,N_14792,N_14858);
nor UO_1360 (O_1360,N_14746,N_14778);
xnor UO_1361 (O_1361,N_14687,N_14590);
and UO_1362 (O_1362,N_14908,N_14875);
or UO_1363 (O_1363,N_14883,N_14925);
or UO_1364 (O_1364,N_14853,N_14757);
and UO_1365 (O_1365,N_14683,N_14986);
xor UO_1366 (O_1366,N_14571,N_14602);
or UO_1367 (O_1367,N_14844,N_14979);
nand UO_1368 (O_1368,N_14933,N_14880);
nand UO_1369 (O_1369,N_14581,N_14742);
xnor UO_1370 (O_1370,N_14979,N_14734);
nand UO_1371 (O_1371,N_14744,N_14913);
xnor UO_1372 (O_1372,N_14586,N_14910);
or UO_1373 (O_1373,N_14861,N_14637);
nand UO_1374 (O_1374,N_14831,N_14809);
xnor UO_1375 (O_1375,N_14709,N_14869);
and UO_1376 (O_1376,N_14712,N_14709);
xnor UO_1377 (O_1377,N_14868,N_14865);
nand UO_1378 (O_1378,N_14619,N_14644);
and UO_1379 (O_1379,N_14961,N_14578);
and UO_1380 (O_1380,N_14811,N_14722);
nand UO_1381 (O_1381,N_14861,N_14812);
nor UO_1382 (O_1382,N_14943,N_14520);
and UO_1383 (O_1383,N_14528,N_14887);
xor UO_1384 (O_1384,N_14861,N_14813);
and UO_1385 (O_1385,N_14813,N_14610);
nor UO_1386 (O_1386,N_14923,N_14970);
and UO_1387 (O_1387,N_14601,N_14641);
nand UO_1388 (O_1388,N_14529,N_14708);
and UO_1389 (O_1389,N_14708,N_14809);
nand UO_1390 (O_1390,N_14533,N_14763);
and UO_1391 (O_1391,N_14748,N_14855);
or UO_1392 (O_1392,N_14771,N_14900);
xnor UO_1393 (O_1393,N_14982,N_14587);
nand UO_1394 (O_1394,N_14618,N_14718);
nand UO_1395 (O_1395,N_14991,N_14781);
nand UO_1396 (O_1396,N_14729,N_14909);
xnor UO_1397 (O_1397,N_14599,N_14987);
nor UO_1398 (O_1398,N_14904,N_14932);
nand UO_1399 (O_1399,N_14618,N_14510);
xnor UO_1400 (O_1400,N_14602,N_14563);
nor UO_1401 (O_1401,N_14554,N_14968);
or UO_1402 (O_1402,N_14661,N_14531);
or UO_1403 (O_1403,N_14635,N_14884);
xor UO_1404 (O_1404,N_14961,N_14713);
xor UO_1405 (O_1405,N_14733,N_14520);
or UO_1406 (O_1406,N_14507,N_14731);
and UO_1407 (O_1407,N_14828,N_14507);
xnor UO_1408 (O_1408,N_14727,N_14765);
nor UO_1409 (O_1409,N_14694,N_14717);
and UO_1410 (O_1410,N_14851,N_14882);
and UO_1411 (O_1411,N_14648,N_14542);
nor UO_1412 (O_1412,N_14930,N_14665);
nand UO_1413 (O_1413,N_14544,N_14572);
or UO_1414 (O_1414,N_14854,N_14506);
nor UO_1415 (O_1415,N_14592,N_14784);
xor UO_1416 (O_1416,N_14926,N_14950);
xnor UO_1417 (O_1417,N_14979,N_14897);
and UO_1418 (O_1418,N_14862,N_14531);
or UO_1419 (O_1419,N_14891,N_14979);
nor UO_1420 (O_1420,N_14829,N_14902);
xnor UO_1421 (O_1421,N_14772,N_14829);
and UO_1422 (O_1422,N_14860,N_14782);
or UO_1423 (O_1423,N_14607,N_14898);
and UO_1424 (O_1424,N_14992,N_14693);
xnor UO_1425 (O_1425,N_14829,N_14866);
or UO_1426 (O_1426,N_14618,N_14582);
xor UO_1427 (O_1427,N_14999,N_14734);
and UO_1428 (O_1428,N_14549,N_14875);
or UO_1429 (O_1429,N_14633,N_14903);
xor UO_1430 (O_1430,N_14525,N_14936);
or UO_1431 (O_1431,N_14721,N_14962);
xor UO_1432 (O_1432,N_14547,N_14502);
nor UO_1433 (O_1433,N_14696,N_14529);
nor UO_1434 (O_1434,N_14576,N_14998);
or UO_1435 (O_1435,N_14844,N_14999);
xnor UO_1436 (O_1436,N_14800,N_14934);
xor UO_1437 (O_1437,N_14840,N_14966);
xnor UO_1438 (O_1438,N_14634,N_14817);
and UO_1439 (O_1439,N_14738,N_14763);
and UO_1440 (O_1440,N_14718,N_14991);
nor UO_1441 (O_1441,N_14654,N_14572);
or UO_1442 (O_1442,N_14542,N_14851);
or UO_1443 (O_1443,N_14632,N_14565);
and UO_1444 (O_1444,N_14543,N_14544);
xnor UO_1445 (O_1445,N_14728,N_14688);
nand UO_1446 (O_1446,N_14925,N_14926);
xnor UO_1447 (O_1447,N_14997,N_14662);
nand UO_1448 (O_1448,N_14948,N_14836);
nor UO_1449 (O_1449,N_14931,N_14785);
nand UO_1450 (O_1450,N_14605,N_14661);
xnor UO_1451 (O_1451,N_14739,N_14724);
nor UO_1452 (O_1452,N_14607,N_14513);
xor UO_1453 (O_1453,N_14946,N_14823);
nor UO_1454 (O_1454,N_14504,N_14892);
nand UO_1455 (O_1455,N_14973,N_14510);
or UO_1456 (O_1456,N_14762,N_14847);
or UO_1457 (O_1457,N_14692,N_14571);
nand UO_1458 (O_1458,N_14709,N_14705);
nor UO_1459 (O_1459,N_14624,N_14934);
xor UO_1460 (O_1460,N_14932,N_14807);
nor UO_1461 (O_1461,N_14866,N_14843);
xor UO_1462 (O_1462,N_14754,N_14802);
nor UO_1463 (O_1463,N_14652,N_14730);
nor UO_1464 (O_1464,N_14937,N_14685);
and UO_1465 (O_1465,N_14756,N_14901);
and UO_1466 (O_1466,N_14703,N_14876);
and UO_1467 (O_1467,N_14724,N_14693);
and UO_1468 (O_1468,N_14554,N_14894);
nand UO_1469 (O_1469,N_14792,N_14564);
nand UO_1470 (O_1470,N_14921,N_14760);
xor UO_1471 (O_1471,N_14727,N_14533);
nor UO_1472 (O_1472,N_14600,N_14655);
nand UO_1473 (O_1473,N_14945,N_14991);
nand UO_1474 (O_1474,N_14756,N_14865);
nand UO_1475 (O_1475,N_14904,N_14755);
or UO_1476 (O_1476,N_14957,N_14826);
xnor UO_1477 (O_1477,N_14677,N_14984);
nand UO_1478 (O_1478,N_14880,N_14579);
and UO_1479 (O_1479,N_14729,N_14737);
nand UO_1480 (O_1480,N_14533,N_14589);
or UO_1481 (O_1481,N_14956,N_14807);
nor UO_1482 (O_1482,N_14928,N_14922);
nand UO_1483 (O_1483,N_14683,N_14518);
nor UO_1484 (O_1484,N_14863,N_14945);
nor UO_1485 (O_1485,N_14509,N_14943);
xnor UO_1486 (O_1486,N_14915,N_14800);
xnor UO_1487 (O_1487,N_14912,N_14631);
or UO_1488 (O_1488,N_14722,N_14566);
or UO_1489 (O_1489,N_14591,N_14659);
and UO_1490 (O_1490,N_14667,N_14729);
xor UO_1491 (O_1491,N_14516,N_14620);
xor UO_1492 (O_1492,N_14525,N_14801);
nor UO_1493 (O_1493,N_14958,N_14647);
nor UO_1494 (O_1494,N_14687,N_14808);
nand UO_1495 (O_1495,N_14705,N_14884);
nor UO_1496 (O_1496,N_14508,N_14809);
nor UO_1497 (O_1497,N_14921,N_14539);
and UO_1498 (O_1498,N_14909,N_14943);
or UO_1499 (O_1499,N_14762,N_14580);
nor UO_1500 (O_1500,N_14797,N_14978);
nor UO_1501 (O_1501,N_14793,N_14845);
xor UO_1502 (O_1502,N_14996,N_14597);
nand UO_1503 (O_1503,N_14912,N_14904);
and UO_1504 (O_1504,N_14976,N_14923);
and UO_1505 (O_1505,N_14680,N_14782);
and UO_1506 (O_1506,N_14579,N_14500);
xnor UO_1507 (O_1507,N_14887,N_14507);
and UO_1508 (O_1508,N_14832,N_14884);
nand UO_1509 (O_1509,N_14605,N_14541);
and UO_1510 (O_1510,N_14820,N_14685);
nand UO_1511 (O_1511,N_14952,N_14941);
and UO_1512 (O_1512,N_14824,N_14504);
and UO_1513 (O_1513,N_14730,N_14708);
xnor UO_1514 (O_1514,N_14978,N_14864);
nor UO_1515 (O_1515,N_14547,N_14939);
nor UO_1516 (O_1516,N_14849,N_14579);
nor UO_1517 (O_1517,N_14539,N_14898);
nor UO_1518 (O_1518,N_14929,N_14871);
or UO_1519 (O_1519,N_14659,N_14981);
and UO_1520 (O_1520,N_14563,N_14513);
xnor UO_1521 (O_1521,N_14781,N_14968);
nor UO_1522 (O_1522,N_14608,N_14858);
nand UO_1523 (O_1523,N_14638,N_14945);
or UO_1524 (O_1524,N_14868,N_14648);
nand UO_1525 (O_1525,N_14614,N_14677);
nor UO_1526 (O_1526,N_14741,N_14846);
and UO_1527 (O_1527,N_14634,N_14770);
or UO_1528 (O_1528,N_14812,N_14734);
nand UO_1529 (O_1529,N_14710,N_14783);
nor UO_1530 (O_1530,N_14800,N_14798);
nor UO_1531 (O_1531,N_14923,N_14699);
and UO_1532 (O_1532,N_14630,N_14842);
or UO_1533 (O_1533,N_14880,N_14604);
nor UO_1534 (O_1534,N_14953,N_14841);
or UO_1535 (O_1535,N_14734,N_14566);
nand UO_1536 (O_1536,N_14793,N_14854);
nand UO_1537 (O_1537,N_14832,N_14589);
nor UO_1538 (O_1538,N_14978,N_14839);
or UO_1539 (O_1539,N_14938,N_14783);
or UO_1540 (O_1540,N_14804,N_14631);
nand UO_1541 (O_1541,N_14564,N_14633);
nand UO_1542 (O_1542,N_14739,N_14776);
and UO_1543 (O_1543,N_14505,N_14843);
nor UO_1544 (O_1544,N_14616,N_14886);
and UO_1545 (O_1545,N_14661,N_14890);
and UO_1546 (O_1546,N_14792,N_14649);
nand UO_1547 (O_1547,N_14717,N_14903);
or UO_1548 (O_1548,N_14625,N_14665);
and UO_1549 (O_1549,N_14596,N_14854);
nand UO_1550 (O_1550,N_14862,N_14966);
xnor UO_1551 (O_1551,N_14636,N_14890);
nand UO_1552 (O_1552,N_14891,N_14647);
nor UO_1553 (O_1553,N_14859,N_14604);
nand UO_1554 (O_1554,N_14960,N_14789);
or UO_1555 (O_1555,N_14532,N_14539);
nand UO_1556 (O_1556,N_14833,N_14781);
or UO_1557 (O_1557,N_14719,N_14606);
nor UO_1558 (O_1558,N_14512,N_14833);
or UO_1559 (O_1559,N_14790,N_14769);
nand UO_1560 (O_1560,N_14660,N_14714);
xnor UO_1561 (O_1561,N_14763,N_14867);
nand UO_1562 (O_1562,N_14908,N_14997);
or UO_1563 (O_1563,N_14730,N_14638);
nor UO_1564 (O_1564,N_14618,N_14682);
xor UO_1565 (O_1565,N_14911,N_14870);
and UO_1566 (O_1566,N_14936,N_14531);
and UO_1567 (O_1567,N_14601,N_14874);
xnor UO_1568 (O_1568,N_14924,N_14945);
and UO_1569 (O_1569,N_14877,N_14792);
nand UO_1570 (O_1570,N_14980,N_14683);
or UO_1571 (O_1571,N_14825,N_14887);
or UO_1572 (O_1572,N_14945,N_14754);
or UO_1573 (O_1573,N_14870,N_14561);
and UO_1574 (O_1574,N_14719,N_14642);
and UO_1575 (O_1575,N_14710,N_14759);
xor UO_1576 (O_1576,N_14690,N_14587);
and UO_1577 (O_1577,N_14775,N_14929);
nand UO_1578 (O_1578,N_14982,N_14516);
nor UO_1579 (O_1579,N_14940,N_14733);
nand UO_1580 (O_1580,N_14932,N_14626);
xor UO_1581 (O_1581,N_14877,N_14853);
nor UO_1582 (O_1582,N_14501,N_14776);
nor UO_1583 (O_1583,N_14963,N_14765);
or UO_1584 (O_1584,N_14646,N_14670);
nand UO_1585 (O_1585,N_14622,N_14509);
nand UO_1586 (O_1586,N_14513,N_14851);
nor UO_1587 (O_1587,N_14658,N_14824);
and UO_1588 (O_1588,N_14712,N_14711);
xnor UO_1589 (O_1589,N_14625,N_14635);
nor UO_1590 (O_1590,N_14963,N_14572);
nand UO_1591 (O_1591,N_14841,N_14985);
or UO_1592 (O_1592,N_14592,N_14637);
and UO_1593 (O_1593,N_14938,N_14706);
nand UO_1594 (O_1594,N_14596,N_14684);
xnor UO_1595 (O_1595,N_14956,N_14516);
nand UO_1596 (O_1596,N_14674,N_14584);
nor UO_1597 (O_1597,N_14994,N_14540);
or UO_1598 (O_1598,N_14678,N_14533);
and UO_1599 (O_1599,N_14988,N_14750);
or UO_1600 (O_1600,N_14531,N_14655);
nand UO_1601 (O_1601,N_14519,N_14683);
and UO_1602 (O_1602,N_14740,N_14794);
xnor UO_1603 (O_1603,N_14668,N_14989);
or UO_1604 (O_1604,N_14936,N_14717);
xor UO_1605 (O_1605,N_14548,N_14579);
nor UO_1606 (O_1606,N_14728,N_14637);
and UO_1607 (O_1607,N_14555,N_14935);
and UO_1608 (O_1608,N_14807,N_14811);
nor UO_1609 (O_1609,N_14607,N_14937);
or UO_1610 (O_1610,N_14897,N_14937);
or UO_1611 (O_1611,N_14635,N_14649);
and UO_1612 (O_1612,N_14577,N_14859);
or UO_1613 (O_1613,N_14940,N_14704);
and UO_1614 (O_1614,N_14712,N_14791);
xnor UO_1615 (O_1615,N_14635,N_14954);
nand UO_1616 (O_1616,N_14825,N_14699);
and UO_1617 (O_1617,N_14666,N_14610);
and UO_1618 (O_1618,N_14967,N_14639);
nor UO_1619 (O_1619,N_14652,N_14763);
xnor UO_1620 (O_1620,N_14822,N_14892);
xor UO_1621 (O_1621,N_14912,N_14894);
or UO_1622 (O_1622,N_14564,N_14901);
nor UO_1623 (O_1623,N_14984,N_14670);
nand UO_1624 (O_1624,N_14669,N_14645);
or UO_1625 (O_1625,N_14852,N_14590);
nand UO_1626 (O_1626,N_14699,N_14751);
xnor UO_1627 (O_1627,N_14522,N_14756);
xor UO_1628 (O_1628,N_14642,N_14897);
or UO_1629 (O_1629,N_14551,N_14578);
or UO_1630 (O_1630,N_14544,N_14979);
and UO_1631 (O_1631,N_14823,N_14914);
and UO_1632 (O_1632,N_14709,N_14761);
nand UO_1633 (O_1633,N_14574,N_14764);
or UO_1634 (O_1634,N_14576,N_14602);
and UO_1635 (O_1635,N_14887,N_14656);
and UO_1636 (O_1636,N_14586,N_14649);
and UO_1637 (O_1637,N_14529,N_14669);
nor UO_1638 (O_1638,N_14624,N_14749);
or UO_1639 (O_1639,N_14545,N_14775);
nand UO_1640 (O_1640,N_14548,N_14621);
or UO_1641 (O_1641,N_14790,N_14783);
and UO_1642 (O_1642,N_14656,N_14811);
nand UO_1643 (O_1643,N_14650,N_14508);
or UO_1644 (O_1644,N_14838,N_14779);
and UO_1645 (O_1645,N_14524,N_14860);
or UO_1646 (O_1646,N_14639,N_14503);
xnor UO_1647 (O_1647,N_14672,N_14568);
or UO_1648 (O_1648,N_14676,N_14669);
or UO_1649 (O_1649,N_14670,N_14900);
nand UO_1650 (O_1650,N_14531,N_14700);
or UO_1651 (O_1651,N_14629,N_14873);
xor UO_1652 (O_1652,N_14805,N_14789);
nand UO_1653 (O_1653,N_14955,N_14543);
nand UO_1654 (O_1654,N_14924,N_14684);
or UO_1655 (O_1655,N_14769,N_14690);
nand UO_1656 (O_1656,N_14786,N_14878);
xnor UO_1657 (O_1657,N_14943,N_14608);
nand UO_1658 (O_1658,N_14537,N_14816);
nor UO_1659 (O_1659,N_14533,N_14797);
nor UO_1660 (O_1660,N_14885,N_14844);
or UO_1661 (O_1661,N_14847,N_14796);
or UO_1662 (O_1662,N_14530,N_14695);
and UO_1663 (O_1663,N_14544,N_14733);
or UO_1664 (O_1664,N_14655,N_14684);
xor UO_1665 (O_1665,N_14759,N_14888);
xnor UO_1666 (O_1666,N_14603,N_14842);
nor UO_1667 (O_1667,N_14783,N_14882);
xor UO_1668 (O_1668,N_14848,N_14564);
xor UO_1669 (O_1669,N_14584,N_14895);
nor UO_1670 (O_1670,N_14658,N_14865);
and UO_1671 (O_1671,N_14796,N_14844);
or UO_1672 (O_1672,N_14604,N_14998);
xor UO_1673 (O_1673,N_14538,N_14885);
and UO_1674 (O_1674,N_14989,N_14763);
or UO_1675 (O_1675,N_14666,N_14970);
nand UO_1676 (O_1676,N_14604,N_14632);
nand UO_1677 (O_1677,N_14651,N_14738);
and UO_1678 (O_1678,N_14864,N_14778);
nand UO_1679 (O_1679,N_14628,N_14606);
nand UO_1680 (O_1680,N_14577,N_14972);
and UO_1681 (O_1681,N_14845,N_14910);
or UO_1682 (O_1682,N_14647,N_14951);
nand UO_1683 (O_1683,N_14672,N_14890);
nor UO_1684 (O_1684,N_14526,N_14646);
xor UO_1685 (O_1685,N_14964,N_14570);
or UO_1686 (O_1686,N_14531,N_14519);
and UO_1687 (O_1687,N_14530,N_14740);
xnor UO_1688 (O_1688,N_14724,N_14871);
or UO_1689 (O_1689,N_14924,N_14589);
and UO_1690 (O_1690,N_14934,N_14683);
nor UO_1691 (O_1691,N_14924,N_14763);
nand UO_1692 (O_1692,N_14779,N_14530);
nor UO_1693 (O_1693,N_14824,N_14991);
nand UO_1694 (O_1694,N_14695,N_14716);
nand UO_1695 (O_1695,N_14828,N_14674);
nor UO_1696 (O_1696,N_14791,N_14677);
or UO_1697 (O_1697,N_14974,N_14600);
nand UO_1698 (O_1698,N_14732,N_14890);
xnor UO_1699 (O_1699,N_14763,N_14508);
and UO_1700 (O_1700,N_14962,N_14840);
nor UO_1701 (O_1701,N_14816,N_14911);
nor UO_1702 (O_1702,N_14825,N_14942);
nand UO_1703 (O_1703,N_14996,N_14736);
or UO_1704 (O_1704,N_14707,N_14734);
and UO_1705 (O_1705,N_14619,N_14775);
or UO_1706 (O_1706,N_14690,N_14796);
nor UO_1707 (O_1707,N_14931,N_14891);
or UO_1708 (O_1708,N_14815,N_14584);
or UO_1709 (O_1709,N_14901,N_14544);
xor UO_1710 (O_1710,N_14721,N_14882);
and UO_1711 (O_1711,N_14581,N_14583);
or UO_1712 (O_1712,N_14724,N_14994);
nand UO_1713 (O_1713,N_14700,N_14875);
xor UO_1714 (O_1714,N_14583,N_14702);
xnor UO_1715 (O_1715,N_14858,N_14870);
or UO_1716 (O_1716,N_14917,N_14968);
and UO_1717 (O_1717,N_14975,N_14680);
nand UO_1718 (O_1718,N_14725,N_14690);
nand UO_1719 (O_1719,N_14797,N_14784);
xnor UO_1720 (O_1720,N_14920,N_14862);
nor UO_1721 (O_1721,N_14525,N_14578);
nand UO_1722 (O_1722,N_14659,N_14818);
nor UO_1723 (O_1723,N_14709,N_14856);
or UO_1724 (O_1724,N_14557,N_14626);
or UO_1725 (O_1725,N_14590,N_14820);
nor UO_1726 (O_1726,N_14710,N_14925);
nand UO_1727 (O_1727,N_14877,N_14913);
and UO_1728 (O_1728,N_14973,N_14599);
or UO_1729 (O_1729,N_14757,N_14987);
xnor UO_1730 (O_1730,N_14960,N_14773);
or UO_1731 (O_1731,N_14831,N_14989);
nor UO_1732 (O_1732,N_14703,N_14711);
nor UO_1733 (O_1733,N_14665,N_14782);
nand UO_1734 (O_1734,N_14796,N_14674);
nand UO_1735 (O_1735,N_14896,N_14870);
nor UO_1736 (O_1736,N_14698,N_14769);
xor UO_1737 (O_1737,N_14732,N_14528);
nor UO_1738 (O_1738,N_14922,N_14513);
and UO_1739 (O_1739,N_14637,N_14569);
xnor UO_1740 (O_1740,N_14555,N_14884);
and UO_1741 (O_1741,N_14775,N_14853);
nor UO_1742 (O_1742,N_14978,N_14842);
nor UO_1743 (O_1743,N_14800,N_14763);
nor UO_1744 (O_1744,N_14956,N_14738);
xnor UO_1745 (O_1745,N_14703,N_14877);
or UO_1746 (O_1746,N_14818,N_14615);
nand UO_1747 (O_1747,N_14585,N_14812);
or UO_1748 (O_1748,N_14579,N_14604);
nand UO_1749 (O_1749,N_14734,N_14742);
xnor UO_1750 (O_1750,N_14690,N_14753);
xnor UO_1751 (O_1751,N_14828,N_14772);
xnor UO_1752 (O_1752,N_14718,N_14558);
xor UO_1753 (O_1753,N_14889,N_14966);
nor UO_1754 (O_1754,N_14779,N_14729);
or UO_1755 (O_1755,N_14683,N_14715);
nor UO_1756 (O_1756,N_14679,N_14997);
nand UO_1757 (O_1757,N_14711,N_14750);
xnor UO_1758 (O_1758,N_14827,N_14870);
and UO_1759 (O_1759,N_14523,N_14704);
xnor UO_1760 (O_1760,N_14640,N_14715);
nand UO_1761 (O_1761,N_14817,N_14917);
nand UO_1762 (O_1762,N_14879,N_14921);
or UO_1763 (O_1763,N_14632,N_14720);
and UO_1764 (O_1764,N_14889,N_14722);
or UO_1765 (O_1765,N_14903,N_14719);
or UO_1766 (O_1766,N_14728,N_14716);
nor UO_1767 (O_1767,N_14567,N_14517);
nand UO_1768 (O_1768,N_14726,N_14969);
and UO_1769 (O_1769,N_14537,N_14693);
nor UO_1770 (O_1770,N_14506,N_14936);
or UO_1771 (O_1771,N_14939,N_14820);
nand UO_1772 (O_1772,N_14739,N_14934);
and UO_1773 (O_1773,N_14754,N_14713);
nor UO_1774 (O_1774,N_14787,N_14971);
or UO_1775 (O_1775,N_14822,N_14526);
and UO_1776 (O_1776,N_14726,N_14745);
or UO_1777 (O_1777,N_14800,N_14998);
xnor UO_1778 (O_1778,N_14990,N_14992);
nand UO_1779 (O_1779,N_14698,N_14888);
nor UO_1780 (O_1780,N_14850,N_14730);
and UO_1781 (O_1781,N_14594,N_14582);
or UO_1782 (O_1782,N_14509,N_14988);
xnor UO_1783 (O_1783,N_14973,N_14949);
and UO_1784 (O_1784,N_14874,N_14719);
xnor UO_1785 (O_1785,N_14632,N_14797);
or UO_1786 (O_1786,N_14679,N_14930);
or UO_1787 (O_1787,N_14802,N_14561);
nor UO_1788 (O_1788,N_14868,N_14677);
nor UO_1789 (O_1789,N_14753,N_14568);
or UO_1790 (O_1790,N_14685,N_14645);
and UO_1791 (O_1791,N_14727,N_14811);
and UO_1792 (O_1792,N_14662,N_14747);
nand UO_1793 (O_1793,N_14587,N_14555);
or UO_1794 (O_1794,N_14698,N_14615);
nor UO_1795 (O_1795,N_14505,N_14634);
and UO_1796 (O_1796,N_14842,N_14622);
and UO_1797 (O_1797,N_14587,N_14783);
or UO_1798 (O_1798,N_14940,N_14615);
and UO_1799 (O_1799,N_14761,N_14808);
xor UO_1800 (O_1800,N_14836,N_14808);
xor UO_1801 (O_1801,N_14875,N_14977);
xnor UO_1802 (O_1802,N_14829,N_14826);
xnor UO_1803 (O_1803,N_14800,N_14700);
or UO_1804 (O_1804,N_14592,N_14851);
and UO_1805 (O_1805,N_14700,N_14515);
nor UO_1806 (O_1806,N_14525,N_14964);
xor UO_1807 (O_1807,N_14851,N_14973);
and UO_1808 (O_1808,N_14866,N_14945);
nor UO_1809 (O_1809,N_14833,N_14758);
nor UO_1810 (O_1810,N_14759,N_14957);
nor UO_1811 (O_1811,N_14662,N_14952);
nor UO_1812 (O_1812,N_14976,N_14616);
or UO_1813 (O_1813,N_14646,N_14856);
xnor UO_1814 (O_1814,N_14526,N_14820);
or UO_1815 (O_1815,N_14984,N_14946);
nand UO_1816 (O_1816,N_14591,N_14530);
nor UO_1817 (O_1817,N_14572,N_14986);
xnor UO_1818 (O_1818,N_14539,N_14803);
or UO_1819 (O_1819,N_14860,N_14821);
nor UO_1820 (O_1820,N_14801,N_14643);
xor UO_1821 (O_1821,N_14709,N_14504);
and UO_1822 (O_1822,N_14737,N_14519);
nand UO_1823 (O_1823,N_14644,N_14569);
nor UO_1824 (O_1824,N_14718,N_14523);
and UO_1825 (O_1825,N_14802,N_14645);
and UO_1826 (O_1826,N_14999,N_14617);
xnor UO_1827 (O_1827,N_14733,N_14854);
and UO_1828 (O_1828,N_14553,N_14581);
or UO_1829 (O_1829,N_14851,N_14621);
and UO_1830 (O_1830,N_14634,N_14803);
xor UO_1831 (O_1831,N_14755,N_14946);
nor UO_1832 (O_1832,N_14882,N_14551);
or UO_1833 (O_1833,N_14849,N_14664);
and UO_1834 (O_1834,N_14975,N_14747);
and UO_1835 (O_1835,N_14611,N_14540);
or UO_1836 (O_1836,N_14852,N_14947);
xnor UO_1837 (O_1837,N_14735,N_14909);
nor UO_1838 (O_1838,N_14577,N_14690);
nor UO_1839 (O_1839,N_14550,N_14785);
or UO_1840 (O_1840,N_14951,N_14591);
xor UO_1841 (O_1841,N_14832,N_14626);
or UO_1842 (O_1842,N_14662,N_14885);
xnor UO_1843 (O_1843,N_14523,N_14939);
and UO_1844 (O_1844,N_14658,N_14718);
and UO_1845 (O_1845,N_14940,N_14817);
and UO_1846 (O_1846,N_14715,N_14518);
nand UO_1847 (O_1847,N_14546,N_14556);
or UO_1848 (O_1848,N_14702,N_14954);
and UO_1849 (O_1849,N_14592,N_14960);
nand UO_1850 (O_1850,N_14530,N_14609);
nand UO_1851 (O_1851,N_14816,N_14586);
and UO_1852 (O_1852,N_14711,N_14820);
or UO_1853 (O_1853,N_14952,N_14930);
nor UO_1854 (O_1854,N_14673,N_14654);
nor UO_1855 (O_1855,N_14918,N_14860);
or UO_1856 (O_1856,N_14813,N_14722);
xnor UO_1857 (O_1857,N_14606,N_14809);
or UO_1858 (O_1858,N_14852,N_14847);
xnor UO_1859 (O_1859,N_14681,N_14906);
xor UO_1860 (O_1860,N_14558,N_14795);
and UO_1861 (O_1861,N_14687,N_14564);
and UO_1862 (O_1862,N_14586,N_14742);
nand UO_1863 (O_1863,N_14512,N_14730);
xor UO_1864 (O_1864,N_14904,N_14722);
and UO_1865 (O_1865,N_14708,N_14657);
or UO_1866 (O_1866,N_14795,N_14756);
or UO_1867 (O_1867,N_14810,N_14676);
and UO_1868 (O_1868,N_14916,N_14959);
nand UO_1869 (O_1869,N_14983,N_14714);
nor UO_1870 (O_1870,N_14548,N_14738);
nor UO_1871 (O_1871,N_14605,N_14869);
or UO_1872 (O_1872,N_14985,N_14931);
nor UO_1873 (O_1873,N_14781,N_14714);
nor UO_1874 (O_1874,N_14520,N_14933);
xnor UO_1875 (O_1875,N_14836,N_14994);
or UO_1876 (O_1876,N_14635,N_14868);
xnor UO_1877 (O_1877,N_14925,N_14723);
nand UO_1878 (O_1878,N_14699,N_14615);
and UO_1879 (O_1879,N_14606,N_14728);
nand UO_1880 (O_1880,N_14689,N_14501);
nand UO_1881 (O_1881,N_14648,N_14851);
nand UO_1882 (O_1882,N_14660,N_14703);
or UO_1883 (O_1883,N_14605,N_14639);
nand UO_1884 (O_1884,N_14823,N_14943);
and UO_1885 (O_1885,N_14507,N_14628);
xor UO_1886 (O_1886,N_14771,N_14718);
or UO_1887 (O_1887,N_14934,N_14671);
or UO_1888 (O_1888,N_14630,N_14503);
nor UO_1889 (O_1889,N_14871,N_14725);
or UO_1890 (O_1890,N_14764,N_14988);
nor UO_1891 (O_1891,N_14671,N_14878);
xnor UO_1892 (O_1892,N_14962,N_14909);
nor UO_1893 (O_1893,N_14533,N_14535);
nor UO_1894 (O_1894,N_14631,N_14718);
xnor UO_1895 (O_1895,N_14582,N_14555);
or UO_1896 (O_1896,N_14811,N_14999);
or UO_1897 (O_1897,N_14762,N_14862);
and UO_1898 (O_1898,N_14958,N_14784);
xnor UO_1899 (O_1899,N_14925,N_14589);
nand UO_1900 (O_1900,N_14637,N_14685);
nand UO_1901 (O_1901,N_14799,N_14915);
or UO_1902 (O_1902,N_14784,N_14974);
nand UO_1903 (O_1903,N_14821,N_14898);
nand UO_1904 (O_1904,N_14688,N_14963);
xnor UO_1905 (O_1905,N_14833,N_14892);
nand UO_1906 (O_1906,N_14797,N_14993);
nor UO_1907 (O_1907,N_14779,N_14902);
and UO_1908 (O_1908,N_14530,N_14954);
nor UO_1909 (O_1909,N_14855,N_14839);
and UO_1910 (O_1910,N_14556,N_14522);
xnor UO_1911 (O_1911,N_14993,N_14817);
or UO_1912 (O_1912,N_14833,N_14506);
xnor UO_1913 (O_1913,N_14751,N_14634);
or UO_1914 (O_1914,N_14677,N_14502);
and UO_1915 (O_1915,N_14857,N_14889);
xor UO_1916 (O_1916,N_14815,N_14964);
and UO_1917 (O_1917,N_14642,N_14593);
nor UO_1918 (O_1918,N_14826,N_14615);
xnor UO_1919 (O_1919,N_14849,N_14540);
and UO_1920 (O_1920,N_14943,N_14764);
nor UO_1921 (O_1921,N_14830,N_14741);
and UO_1922 (O_1922,N_14696,N_14666);
nor UO_1923 (O_1923,N_14644,N_14648);
or UO_1924 (O_1924,N_14992,N_14716);
nor UO_1925 (O_1925,N_14886,N_14563);
and UO_1926 (O_1926,N_14691,N_14763);
nor UO_1927 (O_1927,N_14913,N_14713);
xor UO_1928 (O_1928,N_14945,N_14706);
nand UO_1929 (O_1929,N_14960,N_14932);
nand UO_1930 (O_1930,N_14622,N_14991);
nor UO_1931 (O_1931,N_14685,N_14886);
or UO_1932 (O_1932,N_14506,N_14723);
xor UO_1933 (O_1933,N_14897,N_14741);
nand UO_1934 (O_1934,N_14677,N_14941);
xor UO_1935 (O_1935,N_14944,N_14856);
or UO_1936 (O_1936,N_14517,N_14570);
and UO_1937 (O_1937,N_14542,N_14888);
and UO_1938 (O_1938,N_14826,N_14621);
nand UO_1939 (O_1939,N_14717,N_14692);
xor UO_1940 (O_1940,N_14809,N_14682);
nor UO_1941 (O_1941,N_14768,N_14945);
or UO_1942 (O_1942,N_14658,N_14614);
or UO_1943 (O_1943,N_14709,N_14773);
xor UO_1944 (O_1944,N_14865,N_14848);
nor UO_1945 (O_1945,N_14667,N_14537);
xor UO_1946 (O_1946,N_14628,N_14805);
xnor UO_1947 (O_1947,N_14676,N_14965);
or UO_1948 (O_1948,N_14756,N_14605);
and UO_1949 (O_1949,N_14719,N_14964);
and UO_1950 (O_1950,N_14728,N_14703);
xor UO_1951 (O_1951,N_14817,N_14907);
or UO_1952 (O_1952,N_14859,N_14872);
xor UO_1953 (O_1953,N_14851,N_14649);
or UO_1954 (O_1954,N_14638,N_14699);
xnor UO_1955 (O_1955,N_14773,N_14566);
nor UO_1956 (O_1956,N_14540,N_14841);
or UO_1957 (O_1957,N_14924,N_14647);
nand UO_1958 (O_1958,N_14819,N_14564);
nand UO_1959 (O_1959,N_14514,N_14545);
nor UO_1960 (O_1960,N_14754,N_14946);
nor UO_1961 (O_1961,N_14599,N_14681);
nor UO_1962 (O_1962,N_14561,N_14652);
nor UO_1963 (O_1963,N_14758,N_14903);
or UO_1964 (O_1964,N_14569,N_14733);
nand UO_1965 (O_1965,N_14988,N_14961);
nand UO_1966 (O_1966,N_14596,N_14863);
or UO_1967 (O_1967,N_14973,N_14892);
and UO_1968 (O_1968,N_14956,N_14533);
nand UO_1969 (O_1969,N_14749,N_14805);
xor UO_1970 (O_1970,N_14856,N_14550);
and UO_1971 (O_1971,N_14913,N_14543);
or UO_1972 (O_1972,N_14756,N_14543);
and UO_1973 (O_1973,N_14915,N_14974);
nand UO_1974 (O_1974,N_14883,N_14887);
and UO_1975 (O_1975,N_14811,N_14822);
or UO_1976 (O_1976,N_14563,N_14811);
nor UO_1977 (O_1977,N_14715,N_14963);
nand UO_1978 (O_1978,N_14690,N_14861);
or UO_1979 (O_1979,N_14828,N_14672);
and UO_1980 (O_1980,N_14568,N_14794);
nand UO_1981 (O_1981,N_14624,N_14633);
nand UO_1982 (O_1982,N_14948,N_14559);
nand UO_1983 (O_1983,N_14592,N_14554);
or UO_1984 (O_1984,N_14580,N_14677);
or UO_1985 (O_1985,N_14573,N_14873);
nand UO_1986 (O_1986,N_14753,N_14687);
or UO_1987 (O_1987,N_14641,N_14670);
nand UO_1988 (O_1988,N_14612,N_14561);
nand UO_1989 (O_1989,N_14601,N_14745);
nor UO_1990 (O_1990,N_14960,N_14793);
xor UO_1991 (O_1991,N_14604,N_14684);
nand UO_1992 (O_1992,N_14782,N_14877);
nand UO_1993 (O_1993,N_14737,N_14955);
or UO_1994 (O_1994,N_14703,N_14954);
nand UO_1995 (O_1995,N_14887,N_14713);
nand UO_1996 (O_1996,N_14925,N_14701);
nand UO_1997 (O_1997,N_14616,N_14547);
nand UO_1998 (O_1998,N_14929,N_14902);
or UO_1999 (O_1999,N_14646,N_14778);
endmodule