module basic_1000_10000_1500_5_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_127,In_227);
or U1 (N_1,In_401,In_60);
nand U2 (N_2,In_713,In_188);
nor U3 (N_3,In_950,In_899);
and U4 (N_4,In_789,In_64);
or U5 (N_5,In_612,In_663);
nand U6 (N_6,In_91,In_345);
nor U7 (N_7,In_539,In_957);
nor U8 (N_8,In_43,In_327);
nor U9 (N_9,In_215,In_595);
and U10 (N_10,In_240,In_207);
nand U11 (N_11,In_179,In_121);
or U12 (N_12,In_142,In_765);
xor U13 (N_13,In_278,In_655);
nand U14 (N_14,In_632,In_444);
xnor U15 (N_15,In_7,In_853);
or U16 (N_16,In_318,In_392);
nor U17 (N_17,In_61,In_533);
nand U18 (N_18,In_546,In_849);
or U19 (N_19,In_790,In_840);
xnor U20 (N_20,In_358,In_823);
xor U21 (N_21,In_669,In_872);
nand U22 (N_22,In_217,In_408);
or U23 (N_23,In_357,In_703);
nor U24 (N_24,In_374,In_923);
or U25 (N_25,In_522,In_305);
nor U26 (N_26,In_504,In_945);
nor U27 (N_27,In_762,In_493);
xnor U28 (N_28,In_439,In_193);
and U29 (N_29,In_580,In_96);
or U30 (N_30,In_802,In_25);
nand U31 (N_31,In_914,In_393);
or U32 (N_32,In_432,In_937);
and U33 (N_33,In_675,In_818);
or U34 (N_34,In_190,In_505);
nor U35 (N_35,In_693,In_550);
or U36 (N_36,In_21,In_348);
and U37 (N_37,In_660,In_988);
nor U38 (N_38,In_107,In_996);
nor U39 (N_39,In_806,In_964);
nand U40 (N_40,In_428,In_856);
nor U41 (N_41,In_935,In_176);
nor U42 (N_42,In_756,In_272);
or U43 (N_43,In_841,In_917);
nor U44 (N_44,In_904,In_975);
or U45 (N_45,In_433,In_57);
nand U46 (N_46,In_531,In_999);
and U47 (N_47,In_338,In_316);
nand U48 (N_48,In_745,In_500);
xnor U49 (N_49,In_682,In_426);
and U50 (N_50,In_164,In_535);
nor U51 (N_51,In_503,In_941);
or U52 (N_52,In_890,In_658);
nor U53 (N_53,In_812,In_166);
and U54 (N_54,In_313,In_908);
nand U55 (N_55,In_863,In_650);
and U56 (N_56,In_6,In_424);
and U57 (N_57,In_446,In_162);
or U58 (N_58,In_88,In_150);
and U59 (N_59,In_947,In_77);
nand U60 (N_60,In_564,In_110);
or U61 (N_61,In_239,In_18);
and U62 (N_62,In_679,In_267);
nand U63 (N_63,In_167,In_201);
nand U64 (N_64,In_237,In_741);
and U65 (N_65,In_216,In_259);
nor U66 (N_66,In_599,In_689);
or U67 (N_67,In_773,In_415);
or U68 (N_68,In_931,In_560);
xor U69 (N_69,In_895,In_774);
and U70 (N_70,In_875,In_19);
and U71 (N_71,In_946,In_701);
or U72 (N_72,In_983,In_905);
xor U73 (N_73,In_256,In_205);
xnor U74 (N_74,In_105,In_919);
or U75 (N_75,In_628,In_569);
nor U76 (N_76,In_834,In_353);
xnor U77 (N_77,In_169,In_792);
nor U78 (N_78,In_771,In_113);
and U79 (N_79,In_71,In_132);
and U80 (N_80,In_646,In_966);
nand U81 (N_81,In_95,In_782);
and U82 (N_82,In_661,In_642);
xnor U83 (N_83,In_386,In_833);
nand U84 (N_84,In_709,In_412);
and U85 (N_85,In_75,In_598);
nand U86 (N_86,In_838,In_241);
or U87 (N_87,In_796,In_264);
or U88 (N_88,In_94,In_474);
nand U89 (N_89,In_200,In_168);
xor U90 (N_90,In_156,In_34);
and U91 (N_91,In_615,In_561);
and U92 (N_92,In_108,In_120);
nor U93 (N_93,In_466,In_551);
and U94 (N_94,In_8,In_822);
and U95 (N_95,In_879,In_9);
nor U96 (N_96,In_203,In_274);
or U97 (N_97,In_450,In_720);
nand U98 (N_98,In_987,In_233);
nand U99 (N_99,In_837,In_238);
or U100 (N_100,In_620,In_130);
nand U101 (N_101,In_540,In_468);
xor U102 (N_102,In_517,In_581);
and U103 (N_103,In_594,In_14);
xnor U104 (N_104,In_378,In_461);
and U105 (N_105,In_3,In_287);
and U106 (N_106,In_968,In_739);
or U107 (N_107,In_784,In_587);
nand U108 (N_108,In_496,In_868);
nor U109 (N_109,In_592,In_139);
nand U110 (N_110,In_758,In_600);
and U111 (N_111,In_816,In_70);
or U112 (N_112,In_734,In_194);
nand U113 (N_113,In_394,In_352);
xor U114 (N_114,In_568,In_87);
and U115 (N_115,In_984,In_370);
and U116 (N_116,In_610,In_903);
and U117 (N_117,In_2,In_328);
xor U118 (N_118,In_578,In_102);
and U119 (N_119,In_122,In_62);
nand U120 (N_120,In_949,In_843);
xnor U121 (N_121,In_157,In_706);
nand U122 (N_122,In_831,In_211);
or U123 (N_123,In_997,In_601);
nand U124 (N_124,In_485,In_275);
xor U125 (N_125,In_133,In_13);
or U126 (N_126,In_721,In_435);
nand U127 (N_127,In_636,In_196);
or U128 (N_128,In_613,In_499);
or U129 (N_129,In_757,In_805);
or U130 (N_130,In_422,In_125);
nor U131 (N_131,In_361,In_47);
nor U132 (N_132,In_953,In_372);
and U133 (N_133,In_295,In_730);
and U134 (N_134,In_857,In_733);
nor U135 (N_135,In_854,In_697);
xor U136 (N_136,In_509,In_648);
xor U137 (N_137,In_934,In_798);
nand U138 (N_138,In_421,In_449);
nand U139 (N_139,In_296,In_982);
nand U140 (N_140,In_229,In_251);
xnor U141 (N_141,In_385,In_390);
or U142 (N_142,In_175,In_334);
and U143 (N_143,In_437,In_617);
or U144 (N_144,In_952,In_38);
nor U145 (N_145,In_40,In_89);
nand U146 (N_146,In_845,In_339);
and U147 (N_147,In_626,In_490);
and U148 (N_148,In_944,In_114);
nor U149 (N_149,In_616,In_66);
and U150 (N_150,In_93,In_400);
nor U151 (N_151,In_268,In_574);
nor U152 (N_152,In_448,In_128);
xnor U153 (N_153,In_969,In_524);
nor U154 (N_154,In_629,In_786);
or U155 (N_155,In_498,In_153);
nand U156 (N_156,In_526,In_637);
and U157 (N_157,In_381,In_115);
nor U158 (N_158,In_795,In_570);
xor U159 (N_159,In_452,In_172);
or U160 (N_160,In_413,In_470);
xor U161 (N_161,In_880,In_294);
nand U162 (N_162,In_230,In_340);
nor U163 (N_163,In_245,In_939);
nand U164 (N_164,In_487,In_41);
nand U165 (N_165,In_552,In_191);
and U166 (N_166,In_631,In_673);
nor U167 (N_167,In_92,In_280);
or U168 (N_168,In_871,In_387);
or U169 (N_169,In_436,In_68);
xnor U170 (N_170,In_844,In_22);
or U171 (N_171,In_442,In_549);
or U172 (N_172,In_783,In_140);
or U173 (N_173,In_520,In_149);
nand U174 (N_174,In_544,In_76);
nor U175 (N_175,In_553,In_344);
nand U176 (N_176,In_641,In_404);
and U177 (N_177,In_473,In_618);
and U178 (N_178,In_870,In_971);
and U179 (N_179,In_542,In_177);
nor U180 (N_180,In_684,In_484);
nand U181 (N_181,In_151,In_627);
and U182 (N_182,In_724,In_343);
nor U183 (N_183,In_764,In_10);
xor U184 (N_184,In_141,In_431);
nor U185 (N_185,In_536,In_398);
and U186 (N_186,In_824,In_315);
and U187 (N_187,In_530,In_382);
nor U188 (N_188,In_995,In_375);
or U189 (N_189,In_326,In_51);
nor U190 (N_190,In_700,In_543);
or U191 (N_191,In_154,In_396);
or U192 (N_192,In_187,In_906);
nor U193 (N_193,In_451,In_481);
nand U194 (N_194,In_454,In_692);
or U195 (N_195,In_146,In_277);
nor U196 (N_196,In_434,In_482);
nand U197 (N_197,In_883,In_202);
xor U198 (N_198,In_228,In_586);
nor U199 (N_199,In_56,In_688);
or U200 (N_200,In_29,In_86);
nor U201 (N_201,In_186,In_808);
xnor U202 (N_202,In_244,In_881);
or U203 (N_203,In_694,In_291);
or U204 (N_204,In_329,In_208);
or U205 (N_205,In_192,In_512);
nor U206 (N_206,In_593,In_989);
xnor U207 (N_207,In_391,In_116);
and U208 (N_208,In_930,In_737);
nand U209 (N_209,In_33,In_769);
and U210 (N_210,In_671,In_35);
or U211 (N_211,In_336,In_314);
nor U212 (N_212,In_803,In_819);
or U213 (N_213,In_913,In_257);
xnor U214 (N_214,In_779,In_705);
and U215 (N_215,In_126,In_460);
nor U216 (N_216,In_197,In_309);
or U217 (N_217,In_163,In_321);
or U218 (N_218,In_681,In_73);
nand U219 (N_219,In_1,In_360);
nand U220 (N_220,In_261,In_36);
nand U221 (N_221,In_978,In_788);
nor U222 (N_222,In_83,In_103);
nor U223 (N_223,In_976,In_529);
or U224 (N_224,In_810,In_861);
nor U225 (N_225,In_383,In_926);
nor U226 (N_226,In_254,In_180);
or U227 (N_227,In_556,In_63);
or U228 (N_228,In_928,In_249);
nand U229 (N_229,In_882,In_735);
or U230 (N_230,In_355,In_286);
nor U231 (N_231,In_825,In_471);
and U232 (N_232,In_23,In_477);
or U233 (N_233,In_459,In_112);
nor U234 (N_234,In_376,In_590);
nand U235 (N_235,In_198,In_123);
or U236 (N_236,In_463,In_511);
nand U237 (N_237,In_639,In_665);
or U238 (N_238,In_284,In_732);
or U239 (N_239,In_722,In_770);
or U240 (N_240,In_815,In_183);
nand U241 (N_241,In_514,In_619);
nand U242 (N_242,In_885,In_369);
nand U243 (N_243,In_312,In_643);
or U244 (N_244,In_657,In_748);
xnor U245 (N_245,In_453,In_152);
nor U246 (N_246,In_699,In_90);
and U247 (N_247,In_464,In_42);
and U248 (N_248,In_28,In_534);
nor U249 (N_249,In_377,In_842);
or U250 (N_250,In_331,In_892);
and U251 (N_251,In_585,In_395);
or U252 (N_252,In_389,In_425);
nor U253 (N_253,In_253,In_497);
nand U254 (N_254,In_740,In_109);
nor U255 (N_255,In_475,In_572);
nand U256 (N_256,In_298,In_308);
nand U257 (N_257,In_683,In_528);
or U258 (N_258,In_388,In_708);
nand U259 (N_259,In_900,In_182);
nand U260 (N_260,In_718,In_847);
and U261 (N_261,In_525,In_954);
nand U262 (N_262,In_356,In_776);
nor U263 (N_263,In_635,In_846);
or U264 (N_264,In_623,In_609);
or U265 (N_265,In_323,In_319);
nand U266 (N_266,In_656,In_955);
and U267 (N_267,In_79,In_894);
xnor U268 (N_268,In_144,In_58);
or U269 (N_269,In_342,In_495);
or U270 (N_270,In_324,In_727);
xor U271 (N_271,In_829,In_873);
nor U272 (N_272,In_777,In_645);
and U273 (N_273,In_653,In_420);
nand U274 (N_274,In_69,In_670);
nor U275 (N_275,In_652,In_767);
or U276 (N_276,In_897,In_962);
nand U277 (N_277,In_248,In_72);
or U278 (N_278,In_263,In_46);
and U279 (N_279,In_577,In_998);
nand U280 (N_280,In_65,In_575);
nor U281 (N_281,In_199,In_548);
nor U282 (N_282,In_567,In_799);
nand U283 (N_283,In_429,In_84);
nand U284 (N_284,In_817,In_380);
and U285 (N_285,In_170,In_513);
or U286 (N_286,In_119,In_602);
and U287 (N_287,In_811,In_269);
or U288 (N_288,In_350,In_462);
nand U289 (N_289,In_250,In_925);
or U290 (N_290,In_279,In_100);
and U291 (N_291,In_486,In_99);
or U292 (N_292,In_747,In_82);
xnor U293 (N_293,In_247,In_725);
nor U294 (N_294,In_299,In_858);
or U295 (N_295,In_225,In_440);
and U296 (N_296,In_922,In_850);
and U297 (N_297,In_39,In_985);
or U298 (N_298,In_731,In_974);
nand U299 (N_299,In_521,In_158);
nor U300 (N_300,In_55,In_455);
and U301 (N_301,In_379,In_467);
nand U302 (N_302,In_189,In_686);
or U303 (N_303,In_337,In_970);
nand U304 (N_304,In_5,In_235);
nor U305 (N_305,In_809,In_714);
nor U306 (N_306,In_124,In_898);
nand U307 (N_307,In_888,In_717);
nor U308 (N_308,In_910,In_341);
nor U309 (N_309,In_78,In_44);
nand U310 (N_310,In_49,In_901);
nor U311 (N_311,In_423,In_214);
or U312 (N_312,In_160,In_877);
and U313 (N_313,In_266,In_760);
nand U314 (N_314,In_430,In_565);
nand U315 (N_315,In_876,In_891);
nand U316 (N_316,In_16,In_827);
xor U317 (N_317,In_723,In_915);
nor U318 (N_318,In_527,In_990);
and U319 (N_319,In_364,In_986);
nand U320 (N_320,In_948,In_977);
nor U321 (N_321,In_781,In_98);
and U322 (N_322,In_288,In_961);
nand U323 (N_323,In_101,In_981);
and U324 (N_324,In_373,In_780);
and U325 (N_325,In_184,In_832);
and U326 (N_326,In_625,In_282);
nor U327 (N_327,In_921,In_761);
nor U328 (N_328,In_687,In_793);
nand U329 (N_329,In_557,In_53);
or U330 (N_330,In_292,In_691);
and U331 (N_331,In_728,In_672);
or U332 (N_332,In_860,In_483);
nand U333 (N_333,In_242,In_236);
nand U334 (N_334,In_807,In_902);
or U335 (N_335,In_835,In_111);
nand U336 (N_336,In_607,In_547);
nor U337 (N_337,In_744,In_878);
nor U338 (N_338,In_289,In_994);
xnor U339 (N_339,In_869,In_206);
and U340 (N_340,In_258,In_80);
nand U341 (N_341,In_674,In_31);
or U342 (N_342,In_696,In_346);
nand U343 (N_343,In_973,In_813);
or U344 (N_344,In_909,In_118);
or U345 (N_345,In_407,In_479);
xor U346 (N_346,In_418,In_26);
xnor U347 (N_347,In_219,In_226);
or U348 (N_348,In_300,In_608);
or U349 (N_349,In_738,In_332);
or U350 (N_350,In_307,In_270);
nor U351 (N_351,In_518,In_571);
or U352 (N_352,In_409,In_685);
and U353 (N_353,In_979,In_322);
nand U354 (N_354,In_702,In_4);
nor U355 (N_355,In_828,In_676);
nor U356 (N_356,In_965,In_472);
or U357 (N_357,In_943,In_134);
nand U358 (N_358,In_746,In_52);
or U359 (N_359,In_489,In_508);
or U360 (N_360,In_576,In_644);
and U361 (N_361,In_659,In_306);
or U362 (N_362,In_604,In_715);
and U363 (N_363,In_447,In_678);
nand U364 (N_364,In_293,In_243);
and U365 (N_365,In_638,In_690);
and U366 (N_366,In_145,In_855);
nand U367 (N_367,In_492,In_924);
nand U368 (N_368,In_301,In_402);
and U369 (N_369,In_736,In_74);
nand U370 (N_370,In_726,In_290);
and U371 (N_371,In_918,In_729);
and U372 (N_372,In_751,In_347);
and U373 (N_373,In_537,In_12);
or U374 (N_374,In_27,In_129);
nor U375 (N_375,In_210,In_67);
xor U376 (N_376,In_17,In_680);
or U377 (N_377,In_591,In_754);
nor U378 (N_378,In_614,In_330);
nor U379 (N_379,In_752,In_255);
or U380 (N_380,In_634,In_310);
or U381 (N_381,In_621,In_59);
nor U382 (N_382,In_171,In_668);
nand U383 (N_383,In_972,In_441);
nor U384 (N_384,In_311,In_836);
and U385 (N_385,In_232,In_707);
nand U386 (N_386,In_302,In_583);
and U387 (N_387,In_456,In_763);
and U388 (N_388,In_753,In_862);
nor U389 (N_389,In_325,In_135);
and U390 (N_390,In_416,In_104);
or U391 (N_391,In_20,In_478);
and U392 (N_392,In_624,In_991);
nor U393 (N_393,In_523,In_911);
nand U394 (N_394,In_951,In_488);
or U395 (N_395,In_940,In_886);
or U396 (N_396,In_766,In_667);
nor U397 (N_397,In_801,In_246);
or U398 (N_398,In_384,In_839);
and U399 (N_399,In_181,In_677);
nand U400 (N_400,In_406,In_443);
and U401 (N_401,In_651,In_85);
and U402 (N_402,In_630,In_566);
nor U403 (N_403,In_596,In_317);
nor U404 (N_404,In_563,In_417);
xnor U405 (N_405,In_787,In_775);
and U406 (N_406,In_519,In_695);
and U407 (N_407,In_234,In_588);
xor U408 (N_408,In_893,In_178);
or U409 (N_409,In_884,In_0);
nand U410 (N_410,In_419,In_711);
nand U411 (N_411,In_932,In_960);
nor U412 (N_412,In_174,In_927);
and U413 (N_413,In_510,In_371);
and U414 (N_414,In_719,In_852);
nand U415 (N_415,In_874,In_759);
xor U416 (N_416,In_362,In_359);
or U417 (N_417,In_959,In_480);
nand U418 (N_418,In_368,In_222);
xnor U419 (N_419,In_887,In_54);
nor U420 (N_420,In_545,In_265);
nor U421 (N_421,In_458,In_410);
xor U422 (N_422,In_304,In_411);
nor U423 (N_423,In_559,In_195);
xnor U424 (N_424,In_414,In_778);
nor U425 (N_425,In_438,In_791);
nand U426 (N_426,In_821,In_81);
and U427 (N_427,In_963,In_445);
nor U428 (N_428,In_502,In_993);
or U429 (N_429,In_297,In_814);
nor U430 (N_430,In_224,In_506);
and U431 (N_431,In_320,In_820);
nand U432 (N_432,In_916,In_155);
or U433 (N_433,In_469,In_159);
xnor U434 (N_434,In_622,In_45);
nor U435 (N_435,In_138,In_354);
nand U436 (N_436,In_605,In_538);
xnor U437 (N_437,In_867,In_958);
and U438 (N_438,In_755,In_465);
nand U439 (N_439,In_221,In_907);
or U440 (N_440,In_50,In_349);
nor U441 (N_441,In_936,In_712);
nor U442 (N_442,In_220,In_992);
or U443 (N_443,In_797,In_131);
and U444 (N_444,In_165,In_704);
and U445 (N_445,In_541,In_148);
nand U446 (N_446,In_933,In_143);
and U447 (N_447,In_555,In_276);
nor U448 (N_448,In_896,In_515);
xnor U449 (N_449,In_889,In_185);
nand U450 (N_450,In_507,In_24);
or U451 (N_451,In_501,In_554);
nor U452 (N_452,In_785,In_768);
nor U453 (N_453,In_772,In_213);
and U454 (N_454,In_611,In_32);
nor U455 (N_455,In_136,In_351);
nor U456 (N_456,In_800,In_664);
nand U457 (N_457,In_750,In_137);
and U458 (N_458,In_273,In_252);
nor U459 (N_459,In_956,In_698);
nor U460 (N_460,In_980,In_804);
nand U461 (N_461,In_558,In_865);
nand U462 (N_462,In_491,In_826);
or U463 (N_463,In_367,In_532);
nand U464 (N_464,In_859,In_209);
and U465 (N_465,In_117,In_967);
or U466 (N_466,In_942,In_457);
or U467 (N_467,In_173,In_147);
nor U468 (N_468,In_223,In_920);
nor U469 (N_469,In_48,In_333);
nor U470 (N_470,In_606,In_603);
or U471 (N_471,In_281,In_260);
and U472 (N_472,In_427,In_271);
nand U473 (N_473,In_649,In_204);
nor U474 (N_474,In_866,In_640);
xnor U475 (N_475,In_303,In_589);
xor U476 (N_476,In_97,In_573);
or U477 (N_477,In_562,In_397);
and U478 (N_478,In_743,In_794);
and U479 (N_479,In_830,In_231);
nor U480 (N_480,In_283,In_403);
and U481 (N_481,In_37,In_912);
and U482 (N_482,In_399,In_851);
xnor U483 (N_483,In_742,In_363);
and U484 (N_484,In_494,In_654);
and U485 (N_485,In_582,In_365);
or U486 (N_486,In_938,In_929);
or U487 (N_487,In_516,In_710);
xor U488 (N_488,In_716,In_666);
and U489 (N_489,In_647,In_476);
and U490 (N_490,In_597,In_262);
and U491 (N_491,In_579,In_366);
xor U492 (N_492,In_106,In_161);
nand U493 (N_493,In_848,In_749);
xnor U494 (N_494,In_864,In_633);
nand U495 (N_495,In_15,In_662);
and U496 (N_496,In_285,In_30);
xnor U497 (N_497,In_405,In_212);
and U498 (N_498,In_335,In_11);
xnor U499 (N_499,In_584,In_218);
xnor U500 (N_500,In_592,In_564);
xnor U501 (N_501,In_192,In_127);
and U502 (N_502,In_865,In_45);
nand U503 (N_503,In_666,In_271);
nand U504 (N_504,In_19,In_101);
and U505 (N_505,In_508,In_734);
nand U506 (N_506,In_507,In_731);
nor U507 (N_507,In_585,In_6);
nor U508 (N_508,In_774,In_970);
nor U509 (N_509,In_395,In_739);
or U510 (N_510,In_212,In_659);
and U511 (N_511,In_697,In_324);
nand U512 (N_512,In_871,In_320);
and U513 (N_513,In_492,In_724);
nor U514 (N_514,In_677,In_32);
or U515 (N_515,In_517,In_841);
and U516 (N_516,In_24,In_566);
and U517 (N_517,In_613,In_674);
and U518 (N_518,In_676,In_688);
and U519 (N_519,In_658,In_535);
and U520 (N_520,In_23,In_355);
xor U521 (N_521,In_43,In_629);
or U522 (N_522,In_375,In_335);
and U523 (N_523,In_53,In_787);
nor U524 (N_524,In_363,In_506);
or U525 (N_525,In_933,In_43);
xnor U526 (N_526,In_955,In_353);
xnor U527 (N_527,In_412,In_964);
and U528 (N_528,In_492,In_753);
nand U529 (N_529,In_907,In_339);
nor U530 (N_530,In_124,In_181);
nand U531 (N_531,In_786,In_276);
and U532 (N_532,In_813,In_260);
nor U533 (N_533,In_155,In_798);
or U534 (N_534,In_668,In_929);
nand U535 (N_535,In_111,In_247);
or U536 (N_536,In_968,In_770);
and U537 (N_537,In_888,In_317);
or U538 (N_538,In_542,In_600);
nor U539 (N_539,In_314,In_348);
nand U540 (N_540,In_204,In_723);
nor U541 (N_541,In_699,In_18);
nor U542 (N_542,In_897,In_110);
or U543 (N_543,In_588,In_745);
nor U544 (N_544,In_705,In_999);
and U545 (N_545,In_940,In_631);
xnor U546 (N_546,In_658,In_814);
nand U547 (N_547,In_248,In_846);
xnor U548 (N_548,In_213,In_981);
or U549 (N_549,In_819,In_546);
nand U550 (N_550,In_424,In_513);
xor U551 (N_551,In_22,In_262);
nand U552 (N_552,In_990,In_523);
nand U553 (N_553,In_30,In_198);
nand U554 (N_554,In_679,In_263);
nand U555 (N_555,In_891,In_55);
nor U556 (N_556,In_151,In_295);
and U557 (N_557,In_751,In_700);
xor U558 (N_558,In_126,In_752);
or U559 (N_559,In_643,In_17);
and U560 (N_560,In_775,In_838);
xnor U561 (N_561,In_186,In_792);
nor U562 (N_562,In_155,In_280);
or U563 (N_563,In_552,In_452);
nor U564 (N_564,In_55,In_997);
and U565 (N_565,In_980,In_315);
nand U566 (N_566,In_948,In_14);
and U567 (N_567,In_522,In_188);
nand U568 (N_568,In_244,In_205);
nor U569 (N_569,In_227,In_119);
nor U570 (N_570,In_589,In_254);
nor U571 (N_571,In_170,In_875);
nand U572 (N_572,In_740,In_557);
or U573 (N_573,In_563,In_659);
or U574 (N_574,In_434,In_707);
xor U575 (N_575,In_401,In_11);
nand U576 (N_576,In_449,In_324);
and U577 (N_577,In_784,In_977);
or U578 (N_578,In_969,In_158);
or U579 (N_579,In_377,In_287);
nand U580 (N_580,In_595,In_477);
nand U581 (N_581,In_920,In_621);
nor U582 (N_582,In_312,In_450);
and U583 (N_583,In_215,In_306);
nand U584 (N_584,In_316,In_876);
nor U585 (N_585,In_31,In_156);
nand U586 (N_586,In_738,In_79);
nand U587 (N_587,In_558,In_690);
and U588 (N_588,In_45,In_66);
or U589 (N_589,In_239,In_140);
or U590 (N_590,In_637,In_154);
nand U591 (N_591,In_314,In_974);
and U592 (N_592,In_540,In_616);
and U593 (N_593,In_191,In_43);
or U594 (N_594,In_547,In_27);
nand U595 (N_595,In_580,In_103);
or U596 (N_596,In_919,In_974);
nand U597 (N_597,In_261,In_928);
or U598 (N_598,In_453,In_965);
or U599 (N_599,In_15,In_544);
or U600 (N_600,In_411,In_813);
xor U601 (N_601,In_655,In_382);
nand U602 (N_602,In_693,In_518);
nor U603 (N_603,In_318,In_316);
nor U604 (N_604,In_740,In_116);
or U605 (N_605,In_412,In_437);
or U606 (N_606,In_473,In_768);
or U607 (N_607,In_755,In_984);
or U608 (N_608,In_895,In_975);
nor U609 (N_609,In_43,In_901);
or U610 (N_610,In_587,In_343);
and U611 (N_611,In_41,In_897);
nand U612 (N_612,In_74,In_616);
xor U613 (N_613,In_830,In_72);
xor U614 (N_614,In_950,In_496);
xor U615 (N_615,In_605,In_402);
nor U616 (N_616,In_366,In_423);
xor U617 (N_617,In_773,In_734);
and U618 (N_618,In_569,In_733);
xor U619 (N_619,In_84,In_422);
nor U620 (N_620,In_300,In_516);
xor U621 (N_621,In_350,In_80);
or U622 (N_622,In_201,In_895);
nand U623 (N_623,In_824,In_622);
or U624 (N_624,In_510,In_24);
and U625 (N_625,In_641,In_44);
xor U626 (N_626,In_825,In_522);
and U627 (N_627,In_712,In_824);
nor U628 (N_628,In_720,In_413);
or U629 (N_629,In_737,In_746);
or U630 (N_630,In_158,In_240);
nor U631 (N_631,In_854,In_483);
or U632 (N_632,In_345,In_112);
nand U633 (N_633,In_711,In_731);
nand U634 (N_634,In_649,In_891);
nor U635 (N_635,In_731,In_726);
nor U636 (N_636,In_312,In_528);
xor U637 (N_637,In_772,In_573);
nand U638 (N_638,In_733,In_262);
nor U639 (N_639,In_659,In_924);
and U640 (N_640,In_116,In_318);
nand U641 (N_641,In_718,In_209);
xor U642 (N_642,In_925,In_226);
and U643 (N_643,In_391,In_688);
nand U644 (N_644,In_124,In_254);
and U645 (N_645,In_979,In_764);
nor U646 (N_646,In_870,In_546);
and U647 (N_647,In_364,In_297);
or U648 (N_648,In_237,In_588);
nand U649 (N_649,In_160,In_485);
nand U650 (N_650,In_134,In_322);
or U651 (N_651,In_694,In_143);
nand U652 (N_652,In_110,In_7);
or U653 (N_653,In_475,In_481);
nor U654 (N_654,In_65,In_565);
nor U655 (N_655,In_147,In_765);
and U656 (N_656,In_60,In_368);
and U657 (N_657,In_712,In_241);
nor U658 (N_658,In_31,In_199);
xnor U659 (N_659,In_453,In_46);
xor U660 (N_660,In_173,In_628);
nor U661 (N_661,In_932,In_503);
or U662 (N_662,In_95,In_911);
nand U663 (N_663,In_919,In_93);
nand U664 (N_664,In_369,In_528);
nand U665 (N_665,In_463,In_298);
nand U666 (N_666,In_110,In_289);
and U667 (N_667,In_619,In_39);
or U668 (N_668,In_737,In_326);
nor U669 (N_669,In_879,In_640);
and U670 (N_670,In_894,In_948);
nand U671 (N_671,In_469,In_124);
xor U672 (N_672,In_242,In_399);
and U673 (N_673,In_454,In_820);
or U674 (N_674,In_607,In_147);
or U675 (N_675,In_519,In_314);
nand U676 (N_676,In_727,In_630);
or U677 (N_677,In_258,In_226);
nand U678 (N_678,In_637,In_563);
xor U679 (N_679,In_800,In_683);
nor U680 (N_680,In_592,In_483);
nand U681 (N_681,In_505,In_780);
nand U682 (N_682,In_65,In_821);
or U683 (N_683,In_65,In_501);
or U684 (N_684,In_60,In_699);
and U685 (N_685,In_73,In_585);
and U686 (N_686,In_773,In_710);
nand U687 (N_687,In_448,In_545);
nor U688 (N_688,In_766,In_32);
nand U689 (N_689,In_357,In_144);
or U690 (N_690,In_543,In_39);
nand U691 (N_691,In_536,In_753);
and U692 (N_692,In_308,In_724);
nand U693 (N_693,In_527,In_85);
xor U694 (N_694,In_677,In_988);
nand U695 (N_695,In_651,In_885);
nand U696 (N_696,In_948,In_761);
or U697 (N_697,In_573,In_408);
nand U698 (N_698,In_816,In_432);
nand U699 (N_699,In_182,In_344);
and U700 (N_700,In_59,In_51);
and U701 (N_701,In_448,In_641);
xnor U702 (N_702,In_795,In_181);
nor U703 (N_703,In_859,In_939);
nor U704 (N_704,In_599,In_572);
or U705 (N_705,In_393,In_431);
and U706 (N_706,In_201,In_115);
and U707 (N_707,In_650,In_699);
or U708 (N_708,In_262,In_476);
or U709 (N_709,In_343,In_842);
nand U710 (N_710,In_852,In_149);
nand U711 (N_711,In_974,In_128);
nor U712 (N_712,In_625,In_383);
nor U713 (N_713,In_805,In_22);
nor U714 (N_714,In_809,In_919);
and U715 (N_715,In_416,In_967);
nand U716 (N_716,In_959,In_151);
xnor U717 (N_717,In_364,In_813);
and U718 (N_718,In_664,In_821);
or U719 (N_719,In_240,In_183);
nand U720 (N_720,In_426,In_993);
or U721 (N_721,In_60,In_914);
or U722 (N_722,In_150,In_822);
nor U723 (N_723,In_740,In_690);
nand U724 (N_724,In_591,In_904);
and U725 (N_725,In_382,In_903);
or U726 (N_726,In_118,In_294);
nand U727 (N_727,In_440,In_814);
and U728 (N_728,In_884,In_301);
or U729 (N_729,In_993,In_224);
or U730 (N_730,In_337,In_801);
xor U731 (N_731,In_34,In_703);
nor U732 (N_732,In_639,In_900);
or U733 (N_733,In_184,In_642);
or U734 (N_734,In_49,In_832);
nor U735 (N_735,In_395,In_406);
and U736 (N_736,In_861,In_380);
or U737 (N_737,In_764,In_567);
xor U738 (N_738,In_74,In_32);
or U739 (N_739,In_921,In_577);
nand U740 (N_740,In_547,In_900);
nor U741 (N_741,In_507,In_51);
and U742 (N_742,In_312,In_393);
xnor U743 (N_743,In_391,In_951);
xnor U744 (N_744,In_869,In_484);
nor U745 (N_745,In_956,In_732);
or U746 (N_746,In_89,In_936);
nand U747 (N_747,In_536,In_277);
nor U748 (N_748,In_286,In_887);
nor U749 (N_749,In_625,In_713);
or U750 (N_750,In_808,In_610);
xor U751 (N_751,In_496,In_625);
and U752 (N_752,In_687,In_973);
nand U753 (N_753,In_820,In_664);
nand U754 (N_754,In_561,In_847);
or U755 (N_755,In_897,In_544);
nand U756 (N_756,In_358,In_370);
xnor U757 (N_757,In_228,In_639);
nand U758 (N_758,In_795,In_401);
or U759 (N_759,In_440,In_400);
nor U760 (N_760,In_153,In_218);
nand U761 (N_761,In_930,In_131);
and U762 (N_762,In_237,In_995);
nand U763 (N_763,In_378,In_104);
and U764 (N_764,In_962,In_879);
or U765 (N_765,In_609,In_799);
or U766 (N_766,In_327,In_874);
and U767 (N_767,In_251,In_438);
or U768 (N_768,In_519,In_116);
nand U769 (N_769,In_835,In_980);
nand U770 (N_770,In_513,In_533);
nand U771 (N_771,In_361,In_258);
or U772 (N_772,In_746,In_806);
and U773 (N_773,In_35,In_635);
and U774 (N_774,In_689,In_791);
or U775 (N_775,In_281,In_865);
nor U776 (N_776,In_52,In_356);
and U777 (N_777,In_497,In_40);
nand U778 (N_778,In_104,In_280);
nor U779 (N_779,In_429,In_555);
and U780 (N_780,In_100,In_155);
or U781 (N_781,In_151,In_815);
and U782 (N_782,In_775,In_276);
or U783 (N_783,In_610,In_683);
and U784 (N_784,In_803,In_605);
and U785 (N_785,In_569,In_170);
or U786 (N_786,In_385,In_84);
or U787 (N_787,In_118,In_640);
nand U788 (N_788,In_946,In_97);
nor U789 (N_789,In_348,In_708);
nand U790 (N_790,In_797,In_39);
xnor U791 (N_791,In_919,In_160);
or U792 (N_792,In_641,In_595);
and U793 (N_793,In_458,In_428);
and U794 (N_794,In_912,In_820);
and U795 (N_795,In_422,In_151);
nand U796 (N_796,In_445,In_247);
or U797 (N_797,In_497,In_38);
or U798 (N_798,In_587,In_946);
nand U799 (N_799,In_925,In_337);
nand U800 (N_800,In_376,In_355);
nand U801 (N_801,In_570,In_124);
nor U802 (N_802,In_538,In_144);
nor U803 (N_803,In_424,In_817);
and U804 (N_804,In_959,In_899);
and U805 (N_805,In_580,In_268);
or U806 (N_806,In_4,In_393);
nor U807 (N_807,In_206,In_309);
nor U808 (N_808,In_404,In_945);
xnor U809 (N_809,In_148,In_492);
nand U810 (N_810,In_164,In_278);
nor U811 (N_811,In_312,In_883);
nor U812 (N_812,In_469,In_713);
nor U813 (N_813,In_874,In_717);
nand U814 (N_814,In_521,In_986);
xnor U815 (N_815,In_924,In_204);
or U816 (N_816,In_925,In_595);
xor U817 (N_817,In_961,In_663);
and U818 (N_818,In_810,In_669);
nor U819 (N_819,In_544,In_479);
nand U820 (N_820,In_865,In_600);
or U821 (N_821,In_462,In_380);
nor U822 (N_822,In_160,In_189);
or U823 (N_823,In_683,In_814);
and U824 (N_824,In_464,In_928);
and U825 (N_825,In_326,In_377);
nand U826 (N_826,In_729,In_93);
and U827 (N_827,In_445,In_887);
and U828 (N_828,In_512,In_340);
nor U829 (N_829,In_672,In_747);
and U830 (N_830,In_533,In_303);
nand U831 (N_831,In_329,In_586);
xor U832 (N_832,In_221,In_304);
or U833 (N_833,In_211,In_345);
nand U834 (N_834,In_371,In_522);
nor U835 (N_835,In_963,In_803);
nor U836 (N_836,In_922,In_824);
xnor U837 (N_837,In_697,In_782);
or U838 (N_838,In_849,In_212);
or U839 (N_839,In_342,In_133);
xor U840 (N_840,In_381,In_354);
and U841 (N_841,In_0,In_649);
nor U842 (N_842,In_312,In_537);
nor U843 (N_843,In_434,In_4);
nor U844 (N_844,In_337,In_931);
and U845 (N_845,In_435,In_698);
and U846 (N_846,In_11,In_605);
or U847 (N_847,In_780,In_414);
and U848 (N_848,In_853,In_957);
nor U849 (N_849,In_314,In_165);
or U850 (N_850,In_210,In_501);
and U851 (N_851,In_386,In_201);
or U852 (N_852,In_76,In_837);
nand U853 (N_853,In_456,In_795);
nor U854 (N_854,In_240,In_885);
nor U855 (N_855,In_982,In_430);
or U856 (N_856,In_474,In_624);
nand U857 (N_857,In_952,In_173);
nand U858 (N_858,In_156,In_648);
nand U859 (N_859,In_489,In_743);
and U860 (N_860,In_12,In_260);
nor U861 (N_861,In_363,In_510);
nor U862 (N_862,In_873,In_17);
xnor U863 (N_863,In_605,In_259);
xnor U864 (N_864,In_759,In_165);
and U865 (N_865,In_634,In_850);
or U866 (N_866,In_541,In_212);
nor U867 (N_867,In_812,In_436);
and U868 (N_868,In_811,In_156);
nand U869 (N_869,In_82,In_147);
or U870 (N_870,In_335,In_730);
or U871 (N_871,In_418,In_986);
xor U872 (N_872,In_578,In_163);
nor U873 (N_873,In_983,In_259);
or U874 (N_874,In_877,In_534);
and U875 (N_875,In_232,In_201);
nor U876 (N_876,In_835,In_550);
or U877 (N_877,In_606,In_2);
and U878 (N_878,In_510,In_779);
nor U879 (N_879,In_832,In_575);
or U880 (N_880,In_926,In_800);
nand U881 (N_881,In_989,In_695);
or U882 (N_882,In_103,In_950);
nor U883 (N_883,In_350,In_731);
and U884 (N_884,In_941,In_204);
nor U885 (N_885,In_948,In_40);
nand U886 (N_886,In_529,In_171);
nand U887 (N_887,In_375,In_56);
nand U888 (N_888,In_868,In_140);
nor U889 (N_889,In_875,In_643);
nand U890 (N_890,In_833,In_456);
xor U891 (N_891,In_988,In_658);
and U892 (N_892,In_928,In_102);
or U893 (N_893,In_735,In_386);
nor U894 (N_894,In_425,In_588);
nor U895 (N_895,In_185,In_914);
or U896 (N_896,In_160,In_836);
nand U897 (N_897,In_257,In_645);
and U898 (N_898,In_814,In_870);
nor U899 (N_899,In_858,In_112);
or U900 (N_900,In_660,In_250);
xnor U901 (N_901,In_73,In_749);
and U902 (N_902,In_887,In_27);
nor U903 (N_903,In_176,In_721);
nor U904 (N_904,In_338,In_666);
and U905 (N_905,In_582,In_975);
or U906 (N_906,In_127,In_304);
and U907 (N_907,In_172,In_636);
nand U908 (N_908,In_60,In_64);
nor U909 (N_909,In_237,In_19);
nor U910 (N_910,In_559,In_8);
or U911 (N_911,In_744,In_497);
and U912 (N_912,In_929,In_55);
or U913 (N_913,In_307,In_701);
or U914 (N_914,In_16,In_210);
xor U915 (N_915,In_952,In_679);
nand U916 (N_916,In_765,In_624);
nor U917 (N_917,In_705,In_664);
nor U918 (N_918,In_331,In_136);
xnor U919 (N_919,In_104,In_754);
and U920 (N_920,In_916,In_912);
nor U921 (N_921,In_557,In_89);
nand U922 (N_922,In_793,In_415);
nand U923 (N_923,In_786,In_420);
nand U924 (N_924,In_403,In_720);
or U925 (N_925,In_418,In_907);
or U926 (N_926,In_585,In_39);
or U927 (N_927,In_135,In_740);
and U928 (N_928,In_289,In_98);
or U929 (N_929,In_942,In_878);
nand U930 (N_930,In_952,In_289);
xnor U931 (N_931,In_612,In_214);
or U932 (N_932,In_838,In_983);
or U933 (N_933,In_914,In_895);
and U934 (N_934,In_279,In_291);
xor U935 (N_935,In_871,In_842);
nor U936 (N_936,In_109,In_8);
or U937 (N_937,In_88,In_953);
or U938 (N_938,In_369,In_56);
xnor U939 (N_939,In_467,In_395);
and U940 (N_940,In_781,In_350);
and U941 (N_941,In_173,In_220);
and U942 (N_942,In_959,In_423);
nand U943 (N_943,In_298,In_711);
nor U944 (N_944,In_185,In_92);
nor U945 (N_945,In_397,In_865);
nand U946 (N_946,In_971,In_878);
and U947 (N_947,In_737,In_322);
nand U948 (N_948,In_139,In_393);
and U949 (N_949,In_527,In_603);
nor U950 (N_950,In_732,In_159);
xor U951 (N_951,In_605,In_241);
or U952 (N_952,In_729,In_686);
xnor U953 (N_953,In_687,In_316);
xnor U954 (N_954,In_132,In_225);
nand U955 (N_955,In_124,In_266);
and U956 (N_956,In_526,In_953);
or U957 (N_957,In_980,In_297);
xnor U958 (N_958,In_126,In_219);
nand U959 (N_959,In_920,In_631);
nand U960 (N_960,In_879,In_379);
nor U961 (N_961,In_705,In_126);
nor U962 (N_962,In_799,In_444);
or U963 (N_963,In_802,In_242);
or U964 (N_964,In_836,In_476);
and U965 (N_965,In_406,In_442);
nor U966 (N_966,In_788,In_480);
nor U967 (N_967,In_636,In_792);
or U968 (N_968,In_620,In_473);
or U969 (N_969,In_436,In_29);
and U970 (N_970,In_789,In_10);
nand U971 (N_971,In_209,In_664);
and U972 (N_972,In_450,In_290);
and U973 (N_973,In_296,In_847);
nor U974 (N_974,In_54,In_671);
and U975 (N_975,In_363,In_719);
nor U976 (N_976,In_399,In_88);
nand U977 (N_977,In_279,In_189);
xnor U978 (N_978,In_108,In_440);
xor U979 (N_979,In_513,In_574);
and U980 (N_980,In_480,In_266);
and U981 (N_981,In_646,In_81);
nand U982 (N_982,In_655,In_252);
or U983 (N_983,In_175,In_363);
and U984 (N_984,In_767,In_70);
nand U985 (N_985,In_488,In_370);
and U986 (N_986,In_644,In_846);
nor U987 (N_987,In_208,In_606);
and U988 (N_988,In_388,In_493);
nor U989 (N_989,In_320,In_987);
xor U990 (N_990,In_421,In_400);
or U991 (N_991,In_192,In_804);
or U992 (N_992,In_78,In_975);
or U993 (N_993,In_109,In_370);
nand U994 (N_994,In_739,In_337);
or U995 (N_995,In_173,In_963);
nor U996 (N_996,In_489,In_750);
or U997 (N_997,In_552,In_430);
and U998 (N_998,In_949,In_158);
xnor U999 (N_999,In_731,In_435);
and U1000 (N_1000,In_589,In_550);
nand U1001 (N_1001,In_10,In_480);
nor U1002 (N_1002,In_775,In_270);
or U1003 (N_1003,In_791,In_558);
and U1004 (N_1004,In_813,In_930);
or U1005 (N_1005,In_529,In_59);
nor U1006 (N_1006,In_189,In_776);
nor U1007 (N_1007,In_820,In_268);
or U1008 (N_1008,In_102,In_112);
nand U1009 (N_1009,In_200,In_699);
nand U1010 (N_1010,In_314,In_854);
or U1011 (N_1011,In_852,In_119);
nand U1012 (N_1012,In_348,In_841);
xnor U1013 (N_1013,In_15,In_632);
or U1014 (N_1014,In_796,In_831);
and U1015 (N_1015,In_516,In_153);
and U1016 (N_1016,In_975,In_476);
or U1017 (N_1017,In_358,In_221);
nor U1018 (N_1018,In_31,In_863);
nor U1019 (N_1019,In_42,In_257);
xor U1020 (N_1020,In_959,In_649);
nor U1021 (N_1021,In_226,In_359);
nor U1022 (N_1022,In_714,In_332);
and U1023 (N_1023,In_976,In_598);
nand U1024 (N_1024,In_490,In_682);
nor U1025 (N_1025,In_874,In_927);
and U1026 (N_1026,In_250,In_440);
or U1027 (N_1027,In_570,In_408);
or U1028 (N_1028,In_815,In_683);
nor U1029 (N_1029,In_291,In_230);
nor U1030 (N_1030,In_832,In_960);
nor U1031 (N_1031,In_176,In_559);
xor U1032 (N_1032,In_153,In_626);
and U1033 (N_1033,In_887,In_101);
nand U1034 (N_1034,In_811,In_189);
or U1035 (N_1035,In_150,In_246);
or U1036 (N_1036,In_945,In_637);
nor U1037 (N_1037,In_827,In_230);
or U1038 (N_1038,In_279,In_475);
nor U1039 (N_1039,In_645,In_388);
or U1040 (N_1040,In_204,In_638);
or U1041 (N_1041,In_739,In_773);
and U1042 (N_1042,In_226,In_269);
or U1043 (N_1043,In_267,In_658);
nand U1044 (N_1044,In_995,In_127);
nor U1045 (N_1045,In_775,In_296);
nor U1046 (N_1046,In_352,In_623);
or U1047 (N_1047,In_154,In_680);
nor U1048 (N_1048,In_719,In_410);
nand U1049 (N_1049,In_429,In_954);
nor U1050 (N_1050,In_893,In_755);
and U1051 (N_1051,In_734,In_830);
and U1052 (N_1052,In_18,In_241);
nand U1053 (N_1053,In_980,In_398);
nor U1054 (N_1054,In_648,In_530);
nor U1055 (N_1055,In_399,In_259);
nand U1056 (N_1056,In_53,In_29);
nor U1057 (N_1057,In_467,In_336);
nand U1058 (N_1058,In_230,In_505);
nand U1059 (N_1059,In_333,In_740);
or U1060 (N_1060,In_880,In_119);
nor U1061 (N_1061,In_789,In_284);
or U1062 (N_1062,In_808,In_413);
xnor U1063 (N_1063,In_786,In_51);
and U1064 (N_1064,In_612,In_440);
xnor U1065 (N_1065,In_814,In_742);
or U1066 (N_1066,In_702,In_307);
xnor U1067 (N_1067,In_581,In_793);
xnor U1068 (N_1068,In_771,In_982);
and U1069 (N_1069,In_153,In_700);
or U1070 (N_1070,In_805,In_253);
nand U1071 (N_1071,In_452,In_764);
and U1072 (N_1072,In_966,In_20);
nor U1073 (N_1073,In_380,In_456);
nor U1074 (N_1074,In_983,In_286);
nor U1075 (N_1075,In_748,In_686);
and U1076 (N_1076,In_913,In_450);
and U1077 (N_1077,In_53,In_781);
xnor U1078 (N_1078,In_515,In_939);
nand U1079 (N_1079,In_561,In_99);
or U1080 (N_1080,In_892,In_721);
or U1081 (N_1081,In_293,In_290);
or U1082 (N_1082,In_315,In_34);
nor U1083 (N_1083,In_914,In_508);
nor U1084 (N_1084,In_136,In_483);
or U1085 (N_1085,In_684,In_119);
nand U1086 (N_1086,In_892,In_483);
or U1087 (N_1087,In_149,In_468);
and U1088 (N_1088,In_318,In_651);
or U1089 (N_1089,In_950,In_384);
nand U1090 (N_1090,In_227,In_52);
or U1091 (N_1091,In_372,In_272);
nor U1092 (N_1092,In_847,In_82);
and U1093 (N_1093,In_827,In_615);
and U1094 (N_1094,In_94,In_105);
nor U1095 (N_1095,In_288,In_52);
or U1096 (N_1096,In_400,In_660);
and U1097 (N_1097,In_347,In_316);
xnor U1098 (N_1098,In_128,In_679);
and U1099 (N_1099,In_308,In_494);
nand U1100 (N_1100,In_887,In_52);
or U1101 (N_1101,In_770,In_124);
nor U1102 (N_1102,In_180,In_663);
or U1103 (N_1103,In_150,In_560);
and U1104 (N_1104,In_421,In_892);
xnor U1105 (N_1105,In_582,In_923);
nand U1106 (N_1106,In_856,In_536);
nor U1107 (N_1107,In_312,In_278);
or U1108 (N_1108,In_639,In_727);
or U1109 (N_1109,In_626,In_707);
xor U1110 (N_1110,In_775,In_945);
or U1111 (N_1111,In_11,In_421);
nand U1112 (N_1112,In_48,In_495);
or U1113 (N_1113,In_179,In_277);
and U1114 (N_1114,In_304,In_980);
and U1115 (N_1115,In_866,In_123);
xnor U1116 (N_1116,In_889,In_740);
or U1117 (N_1117,In_744,In_215);
xnor U1118 (N_1118,In_302,In_787);
or U1119 (N_1119,In_483,In_481);
nor U1120 (N_1120,In_602,In_273);
nand U1121 (N_1121,In_653,In_66);
or U1122 (N_1122,In_117,In_468);
nand U1123 (N_1123,In_775,In_88);
nor U1124 (N_1124,In_974,In_597);
or U1125 (N_1125,In_570,In_30);
and U1126 (N_1126,In_24,In_381);
or U1127 (N_1127,In_855,In_766);
nor U1128 (N_1128,In_577,In_178);
or U1129 (N_1129,In_37,In_215);
or U1130 (N_1130,In_492,In_968);
and U1131 (N_1131,In_618,In_326);
nor U1132 (N_1132,In_210,In_998);
and U1133 (N_1133,In_666,In_339);
nand U1134 (N_1134,In_742,In_193);
nand U1135 (N_1135,In_384,In_721);
xor U1136 (N_1136,In_346,In_828);
nand U1137 (N_1137,In_842,In_195);
or U1138 (N_1138,In_927,In_976);
nand U1139 (N_1139,In_954,In_97);
nor U1140 (N_1140,In_563,In_751);
and U1141 (N_1141,In_400,In_497);
nor U1142 (N_1142,In_702,In_421);
nor U1143 (N_1143,In_505,In_394);
nand U1144 (N_1144,In_667,In_996);
and U1145 (N_1145,In_529,In_849);
nand U1146 (N_1146,In_262,In_204);
nor U1147 (N_1147,In_653,In_285);
nor U1148 (N_1148,In_250,In_273);
or U1149 (N_1149,In_162,In_47);
and U1150 (N_1150,In_114,In_677);
nor U1151 (N_1151,In_946,In_234);
nand U1152 (N_1152,In_515,In_218);
nand U1153 (N_1153,In_711,In_423);
and U1154 (N_1154,In_208,In_343);
and U1155 (N_1155,In_69,In_373);
nand U1156 (N_1156,In_487,In_478);
or U1157 (N_1157,In_518,In_756);
or U1158 (N_1158,In_211,In_921);
xor U1159 (N_1159,In_511,In_118);
nor U1160 (N_1160,In_633,In_759);
and U1161 (N_1161,In_187,In_479);
nand U1162 (N_1162,In_143,In_67);
nand U1163 (N_1163,In_778,In_275);
and U1164 (N_1164,In_10,In_326);
or U1165 (N_1165,In_24,In_149);
nand U1166 (N_1166,In_507,In_679);
or U1167 (N_1167,In_377,In_783);
or U1168 (N_1168,In_880,In_610);
and U1169 (N_1169,In_648,In_174);
nand U1170 (N_1170,In_968,In_351);
and U1171 (N_1171,In_436,In_434);
or U1172 (N_1172,In_502,In_2);
and U1173 (N_1173,In_969,In_501);
nand U1174 (N_1174,In_896,In_627);
xnor U1175 (N_1175,In_602,In_542);
nor U1176 (N_1176,In_585,In_756);
nand U1177 (N_1177,In_592,In_136);
nor U1178 (N_1178,In_197,In_182);
nor U1179 (N_1179,In_281,In_371);
and U1180 (N_1180,In_358,In_680);
nor U1181 (N_1181,In_252,In_200);
xnor U1182 (N_1182,In_558,In_110);
or U1183 (N_1183,In_13,In_765);
nor U1184 (N_1184,In_299,In_738);
nor U1185 (N_1185,In_910,In_118);
or U1186 (N_1186,In_657,In_670);
and U1187 (N_1187,In_103,In_168);
or U1188 (N_1188,In_44,In_558);
and U1189 (N_1189,In_762,In_206);
nor U1190 (N_1190,In_640,In_441);
nand U1191 (N_1191,In_1,In_761);
and U1192 (N_1192,In_485,In_142);
xor U1193 (N_1193,In_843,In_389);
and U1194 (N_1194,In_935,In_502);
nor U1195 (N_1195,In_179,In_531);
or U1196 (N_1196,In_211,In_212);
nand U1197 (N_1197,In_167,In_983);
nor U1198 (N_1198,In_181,In_327);
and U1199 (N_1199,In_92,In_934);
or U1200 (N_1200,In_633,In_36);
xor U1201 (N_1201,In_389,In_246);
or U1202 (N_1202,In_503,In_28);
or U1203 (N_1203,In_382,In_967);
or U1204 (N_1204,In_366,In_969);
or U1205 (N_1205,In_924,In_910);
or U1206 (N_1206,In_768,In_321);
nor U1207 (N_1207,In_338,In_2);
nor U1208 (N_1208,In_235,In_836);
xor U1209 (N_1209,In_671,In_430);
nand U1210 (N_1210,In_389,In_328);
and U1211 (N_1211,In_296,In_751);
xor U1212 (N_1212,In_763,In_836);
or U1213 (N_1213,In_421,In_237);
and U1214 (N_1214,In_292,In_102);
nand U1215 (N_1215,In_206,In_839);
or U1216 (N_1216,In_543,In_912);
nor U1217 (N_1217,In_695,In_461);
nand U1218 (N_1218,In_787,In_894);
xor U1219 (N_1219,In_485,In_119);
or U1220 (N_1220,In_143,In_178);
and U1221 (N_1221,In_552,In_261);
nand U1222 (N_1222,In_899,In_117);
and U1223 (N_1223,In_380,In_798);
nor U1224 (N_1224,In_725,In_592);
nor U1225 (N_1225,In_695,In_146);
and U1226 (N_1226,In_208,In_775);
nand U1227 (N_1227,In_27,In_391);
nor U1228 (N_1228,In_171,In_174);
and U1229 (N_1229,In_262,In_240);
xor U1230 (N_1230,In_515,In_949);
or U1231 (N_1231,In_443,In_410);
xor U1232 (N_1232,In_559,In_787);
nand U1233 (N_1233,In_595,In_404);
or U1234 (N_1234,In_194,In_378);
nand U1235 (N_1235,In_171,In_742);
xor U1236 (N_1236,In_588,In_898);
xnor U1237 (N_1237,In_992,In_980);
nand U1238 (N_1238,In_74,In_905);
xnor U1239 (N_1239,In_738,In_154);
nand U1240 (N_1240,In_155,In_534);
nand U1241 (N_1241,In_550,In_813);
xnor U1242 (N_1242,In_284,In_41);
and U1243 (N_1243,In_906,In_767);
or U1244 (N_1244,In_70,In_672);
nand U1245 (N_1245,In_197,In_708);
or U1246 (N_1246,In_42,In_359);
nand U1247 (N_1247,In_792,In_763);
xnor U1248 (N_1248,In_517,In_997);
nand U1249 (N_1249,In_893,In_16);
and U1250 (N_1250,In_552,In_426);
nand U1251 (N_1251,In_136,In_446);
or U1252 (N_1252,In_698,In_617);
nand U1253 (N_1253,In_684,In_716);
xor U1254 (N_1254,In_119,In_764);
and U1255 (N_1255,In_797,In_183);
xnor U1256 (N_1256,In_450,In_846);
nand U1257 (N_1257,In_544,In_33);
and U1258 (N_1258,In_282,In_397);
nor U1259 (N_1259,In_833,In_897);
nand U1260 (N_1260,In_466,In_167);
xnor U1261 (N_1261,In_926,In_199);
and U1262 (N_1262,In_399,In_770);
nand U1263 (N_1263,In_467,In_110);
nor U1264 (N_1264,In_962,In_365);
nand U1265 (N_1265,In_769,In_6);
and U1266 (N_1266,In_356,In_285);
nand U1267 (N_1267,In_473,In_108);
nand U1268 (N_1268,In_200,In_679);
and U1269 (N_1269,In_370,In_10);
or U1270 (N_1270,In_418,In_416);
nor U1271 (N_1271,In_591,In_505);
nor U1272 (N_1272,In_35,In_167);
nand U1273 (N_1273,In_999,In_254);
nor U1274 (N_1274,In_720,In_616);
nand U1275 (N_1275,In_378,In_537);
or U1276 (N_1276,In_546,In_998);
nor U1277 (N_1277,In_371,In_882);
nor U1278 (N_1278,In_359,In_328);
and U1279 (N_1279,In_102,In_178);
nor U1280 (N_1280,In_426,In_175);
nor U1281 (N_1281,In_99,In_426);
or U1282 (N_1282,In_299,In_961);
nand U1283 (N_1283,In_820,In_853);
and U1284 (N_1284,In_562,In_278);
and U1285 (N_1285,In_382,In_272);
or U1286 (N_1286,In_590,In_17);
nand U1287 (N_1287,In_904,In_735);
nor U1288 (N_1288,In_807,In_157);
nor U1289 (N_1289,In_868,In_955);
and U1290 (N_1290,In_796,In_452);
nor U1291 (N_1291,In_245,In_685);
xor U1292 (N_1292,In_643,In_564);
or U1293 (N_1293,In_171,In_17);
nand U1294 (N_1294,In_506,In_121);
nand U1295 (N_1295,In_958,In_571);
and U1296 (N_1296,In_211,In_354);
nand U1297 (N_1297,In_140,In_938);
nand U1298 (N_1298,In_672,In_462);
nand U1299 (N_1299,In_429,In_135);
nor U1300 (N_1300,In_343,In_917);
and U1301 (N_1301,In_222,In_471);
and U1302 (N_1302,In_786,In_828);
and U1303 (N_1303,In_204,In_335);
or U1304 (N_1304,In_525,In_519);
nor U1305 (N_1305,In_719,In_517);
and U1306 (N_1306,In_217,In_204);
nor U1307 (N_1307,In_722,In_705);
or U1308 (N_1308,In_837,In_411);
or U1309 (N_1309,In_533,In_884);
nor U1310 (N_1310,In_975,In_838);
nor U1311 (N_1311,In_972,In_178);
nand U1312 (N_1312,In_919,In_961);
or U1313 (N_1313,In_113,In_612);
nor U1314 (N_1314,In_488,In_175);
and U1315 (N_1315,In_72,In_352);
nand U1316 (N_1316,In_125,In_43);
and U1317 (N_1317,In_705,In_490);
nor U1318 (N_1318,In_666,In_639);
and U1319 (N_1319,In_272,In_161);
or U1320 (N_1320,In_946,In_382);
or U1321 (N_1321,In_27,In_803);
nand U1322 (N_1322,In_497,In_963);
nand U1323 (N_1323,In_561,In_975);
and U1324 (N_1324,In_135,In_626);
nor U1325 (N_1325,In_751,In_390);
nor U1326 (N_1326,In_480,In_377);
nand U1327 (N_1327,In_572,In_240);
nand U1328 (N_1328,In_769,In_302);
and U1329 (N_1329,In_224,In_444);
nor U1330 (N_1330,In_399,In_632);
nor U1331 (N_1331,In_60,In_352);
and U1332 (N_1332,In_824,In_168);
and U1333 (N_1333,In_909,In_119);
or U1334 (N_1334,In_676,In_149);
and U1335 (N_1335,In_546,In_842);
nand U1336 (N_1336,In_962,In_938);
nand U1337 (N_1337,In_595,In_313);
xor U1338 (N_1338,In_784,In_811);
or U1339 (N_1339,In_10,In_455);
nand U1340 (N_1340,In_542,In_124);
and U1341 (N_1341,In_158,In_257);
and U1342 (N_1342,In_255,In_941);
nor U1343 (N_1343,In_874,In_912);
nand U1344 (N_1344,In_577,In_205);
xnor U1345 (N_1345,In_933,In_729);
nor U1346 (N_1346,In_579,In_973);
nor U1347 (N_1347,In_668,In_183);
nand U1348 (N_1348,In_814,In_542);
nor U1349 (N_1349,In_660,In_278);
nor U1350 (N_1350,In_885,In_686);
nor U1351 (N_1351,In_659,In_258);
or U1352 (N_1352,In_553,In_604);
nor U1353 (N_1353,In_939,In_767);
and U1354 (N_1354,In_76,In_445);
nor U1355 (N_1355,In_408,In_205);
nand U1356 (N_1356,In_931,In_540);
or U1357 (N_1357,In_916,In_554);
xor U1358 (N_1358,In_264,In_293);
or U1359 (N_1359,In_763,In_576);
nand U1360 (N_1360,In_304,In_732);
and U1361 (N_1361,In_374,In_152);
nand U1362 (N_1362,In_921,In_96);
or U1363 (N_1363,In_775,In_659);
and U1364 (N_1364,In_849,In_302);
nand U1365 (N_1365,In_683,In_886);
or U1366 (N_1366,In_860,In_128);
or U1367 (N_1367,In_724,In_337);
nand U1368 (N_1368,In_169,In_797);
xor U1369 (N_1369,In_624,In_829);
nand U1370 (N_1370,In_960,In_23);
and U1371 (N_1371,In_483,In_340);
and U1372 (N_1372,In_770,In_451);
or U1373 (N_1373,In_238,In_486);
nand U1374 (N_1374,In_560,In_232);
or U1375 (N_1375,In_575,In_693);
and U1376 (N_1376,In_249,In_539);
nor U1377 (N_1377,In_730,In_545);
nand U1378 (N_1378,In_758,In_834);
xnor U1379 (N_1379,In_890,In_928);
nor U1380 (N_1380,In_691,In_443);
or U1381 (N_1381,In_785,In_105);
nand U1382 (N_1382,In_516,In_339);
or U1383 (N_1383,In_253,In_875);
and U1384 (N_1384,In_480,In_334);
or U1385 (N_1385,In_967,In_547);
xnor U1386 (N_1386,In_65,In_747);
nor U1387 (N_1387,In_716,In_227);
and U1388 (N_1388,In_138,In_393);
and U1389 (N_1389,In_10,In_498);
and U1390 (N_1390,In_144,In_880);
nor U1391 (N_1391,In_356,In_530);
or U1392 (N_1392,In_909,In_689);
and U1393 (N_1393,In_206,In_384);
and U1394 (N_1394,In_186,In_992);
nand U1395 (N_1395,In_577,In_764);
or U1396 (N_1396,In_693,In_879);
nor U1397 (N_1397,In_388,In_996);
xor U1398 (N_1398,In_967,In_783);
nor U1399 (N_1399,In_886,In_518);
and U1400 (N_1400,In_815,In_862);
nor U1401 (N_1401,In_278,In_945);
nand U1402 (N_1402,In_39,In_598);
or U1403 (N_1403,In_872,In_564);
xor U1404 (N_1404,In_929,In_421);
nor U1405 (N_1405,In_445,In_369);
nand U1406 (N_1406,In_991,In_767);
nand U1407 (N_1407,In_71,In_355);
and U1408 (N_1408,In_478,In_660);
nor U1409 (N_1409,In_787,In_890);
and U1410 (N_1410,In_785,In_492);
nand U1411 (N_1411,In_883,In_198);
or U1412 (N_1412,In_602,In_762);
nand U1413 (N_1413,In_436,In_218);
xor U1414 (N_1414,In_485,In_55);
nand U1415 (N_1415,In_791,In_15);
and U1416 (N_1416,In_445,In_989);
nand U1417 (N_1417,In_354,In_910);
nand U1418 (N_1418,In_871,In_858);
and U1419 (N_1419,In_891,In_862);
nand U1420 (N_1420,In_365,In_339);
and U1421 (N_1421,In_687,In_864);
or U1422 (N_1422,In_415,In_715);
xnor U1423 (N_1423,In_454,In_549);
and U1424 (N_1424,In_331,In_478);
and U1425 (N_1425,In_43,In_617);
nor U1426 (N_1426,In_178,In_987);
nand U1427 (N_1427,In_824,In_981);
xnor U1428 (N_1428,In_496,In_215);
and U1429 (N_1429,In_366,In_261);
or U1430 (N_1430,In_734,In_665);
nand U1431 (N_1431,In_538,In_271);
or U1432 (N_1432,In_567,In_375);
or U1433 (N_1433,In_115,In_893);
or U1434 (N_1434,In_579,In_568);
xor U1435 (N_1435,In_360,In_189);
and U1436 (N_1436,In_299,In_674);
or U1437 (N_1437,In_65,In_399);
xor U1438 (N_1438,In_539,In_392);
nor U1439 (N_1439,In_290,In_542);
nor U1440 (N_1440,In_543,In_848);
nand U1441 (N_1441,In_742,In_460);
and U1442 (N_1442,In_506,In_653);
and U1443 (N_1443,In_910,In_5);
xor U1444 (N_1444,In_457,In_688);
and U1445 (N_1445,In_848,In_263);
and U1446 (N_1446,In_321,In_351);
or U1447 (N_1447,In_147,In_205);
nor U1448 (N_1448,In_918,In_365);
nand U1449 (N_1449,In_169,In_517);
nand U1450 (N_1450,In_24,In_634);
nand U1451 (N_1451,In_33,In_763);
or U1452 (N_1452,In_150,In_275);
or U1453 (N_1453,In_841,In_814);
nand U1454 (N_1454,In_389,In_364);
nand U1455 (N_1455,In_66,In_902);
or U1456 (N_1456,In_712,In_959);
nand U1457 (N_1457,In_115,In_42);
nor U1458 (N_1458,In_962,In_773);
nand U1459 (N_1459,In_581,In_110);
or U1460 (N_1460,In_402,In_723);
and U1461 (N_1461,In_914,In_470);
xnor U1462 (N_1462,In_224,In_767);
nand U1463 (N_1463,In_654,In_808);
or U1464 (N_1464,In_226,In_33);
nor U1465 (N_1465,In_230,In_302);
nand U1466 (N_1466,In_265,In_834);
and U1467 (N_1467,In_904,In_862);
or U1468 (N_1468,In_769,In_881);
nand U1469 (N_1469,In_87,In_301);
and U1470 (N_1470,In_119,In_938);
nand U1471 (N_1471,In_464,In_984);
nand U1472 (N_1472,In_559,In_608);
or U1473 (N_1473,In_184,In_541);
or U1474 (N_1474,In_904,In_138);
or U1475 (N_1475,In_497,In_28);
nor U1476 (N_1476,In_377,In_957);
nand U1477 (N_1477,In_642,In_727);
nand U1478 (N_1478,In_426,In_905);
xor U1479 (N_1479,In_907,In_782);
nor U1480 (N_1480,In_222,In_539);
or U1481 (N_1481,In_941,In_424);
or U1482 (N_1482,In_593,In_275);
and U1483 (N_1483,In_785,In_804);
nor U1484 (N_1484,In_397,In_993);
nor U1485 (N_1485,In_392,In_157);
or U1486 (N_1486,In_406,In_292);
and U1487 (N_1487,In_167,In_545);
or U1488 (N_1488,In_181,In_10);
nor U1489 (N_1489,In_419,In_258);
or U1490 (N_1490,In_358,In_411);
nor U1491 (N_1491,In_176,In_547);
or U1492 (N_1492,In_887,In_218);
or U1493 (N_1493,In_65,In_308);
xnor U1494 (N_1494,In_391,In_142);
nor U1495 (N_1495,In_847,In_964);
nand U1496 (N_1496,In_682,In_276);
nand U1497 (N_1497,In_640,In_692);
nand U1498 (N_1498,In_134,In_82);
or U1499 (N_1499,In_687,In_984);
xnor U1500 (N_1500,In_780,In_243);
and U1501 (N_1501,In_676,In_952);
or U1502 (N_1502,In_458,In_73);
or U1503 (N_1503,In_612,In_235);
and U1504 (N_1504,In_563,In_237);
xor U1505 (N_1505,In_998,In_409);
nand U1506 (N_1506,In_732,In_997);
xnor U1507 (N_1507,In_280,In_123);
xnor U1508 (N_1508,In_717,In_95);
and U1509 (N_1509,In_821,In_462);
nor U1510 (N_1510,In_505,In_661);
and U1511 (N_1511,In_321,In_60);
or U1512 (N_1512,In_674,In_816);
xor U1513 (N_1513,In_505,In_839);
nor U1514 (N_1514,In_428,In_719);
xnor U1515 (N_1515,In_847,In_759);
nand U1516 (N_1516,In_553,In_991);
nor U1517 (N_1517,In_992,In_328);
xor U1518 (N_1518,In_209,In_757);
and U1519 (N_1519,In_131,In_87);
or U1520 (N_1520,In_920,In_611);
or U1521 (N_1521,In_706,In_387);
xnor U1522 (N_1522,In_523,In_693);
or U1523 (N_1523,In_204,In_749);
nand U1524 (N_1524,In_747,In_705);
or U1525 (N_1525,In_567,In_258);
or U1526 (N_1526,In_445,In_808);
or U1527 (N_1527,In_165,In_281);
and U1528 (N_1528,In_601,In_926);
and U1529 (N_1529,In_724,In_760);
nand U1530 (N_1530,In_778,In_691);
nor U1531 (N_1531,In_296,In_169);
nand U1532 (N_1532,In_410,In_732);
and U1533 (N_1533,In_854,In_715);
nand U1534 (N_1534,In_395,In_684);
nor U1535 (N_1535,In_426,In_793);
nor U1536 (N_1536,In_307,In_472);
nand U1537 (N_1537,In_232,In_50);
or U1538 (N_1538,In_748,In_905);
or U1539 (N_1539,In_399,In_469);
and U1540 (N_1540,In_659,In_99);
and U1541 (N_1541,In_679,In_129);
or U1542 (N_1542,In_817,In_182);
nand U1543 (N_1543,In_609,In_332);
nand U1544 (N_1544,In_550,In_623);
and U1545 (N_1545,In_144,In_543);
xor U1546 (N_1546,In_399,In_697);
or U1547 (N_1547,In_838,In_760);
and U1548 (N_1548,In_194,In_902);
nor U1549 (N_1549,In_648,In_570);
nor U1550 (N_1550,In_807,In_724);
nor U1551 (N_1551,In_487,In_552);
nand U1552 (N_1552,In_623,In_151);
or U1553 (N_1553,In_265,In_168);
nor U1554 (N_1554,In_450,In_422);
xor U1555 (N_1555,In_983,In_906);
and U1556 (N_1556,In_595,In_648);
nand U1557 (N_1557,In_24,In_14);
or U1558 (N_1558,In_367,In_501);
and U1559 (N_1559,In_726,In_795);
and U1560 (N_1560,In_669,In_379);
and U1561 (N_1561,In_670,In_40);
nor U1562 (N_1562,In_57,In_932);
and U1563 (N_1563,In_100,In_842);
nor U1564 (N_1564,In_670,In_933);
or U1565 (N_1565,In_552,In_319);
xnor U1566 (N_1566,In_969,In_564);
and U1567 (N_1567,In_935,In_406);
nand U1568 (N_1568,In_477,In_923);
nand U1569 (N_1569,In_401,In_149);
nand U1570 (N_1570,In_404,In_195);
nor U1571 (N_1571,In_995,In_515);
nand U1572 (N_1572,In_921,In_969);
nor U1573 (N_1573,In_346,In_889);
and U1574 (N_1574,In_97,In_204);
or U1575 (N_1575,In_716,In_889);
nand U1576 (N_1576,In_629,In_982);
and U1577 (N_1577,In_350,In_48);
or U1578 (N_1578,In_437,In_671);
or U1579 (N_1579,In_380,In_25);
nor U1580 (N_1580,In_236,In_355);
nand U1581 (N_1581,In_30,In_585);
nor U1582 (N_1582,In_243,In_305);
and U1583 (N_1583,In_1,In_231);
and U1584 (N_1584,In_750,In_202);
or U1585 (N_1585,In_526,In_349);
and U1586 (N_1586,In_419,In_857);
nor U1587 (N_1587,In_515,In_474);
nand U1588 (N_1588,In_730,In_466);
or U1589 (N_1589,In_717,In_492);
nor U1590 (N_1590,In_318,In_173);
nand U1591 (N_1591,In_856,In_604);
xnor U1592 (N_1592,In_745,In_573);
or U1593 (N_1593,In_99,In_896);
nor U1594 (N_1594,In_597,In_586);
nor U1595 (N_1595,In_666,In_81);
and U1596 (N_1596,In_719,In_594);
nand U1597 (N_1597,In_776,In_103);
nand U1598 (N_1598,In_124,In_155);
nand U1599 (N_1599,In_825,In_102);
or U1600 (N_1600,In_632,In_671);
and U1601 (N_1601,In_507,In_869);
and U1602 (N_1602,In_994,In_824);
nand U1603 (N_1603,In_385,In_231);
and U1604 (N_1604,In_557,In_736);
nand U1605 (N_1605,In_330,In_897);
xnor U1606 (N_1606,In_434,In_677);
nor U1607 (N_1607,In_582,In_65);
and U1608 (N_1608,In_174,In_819);
nand U1609 (N_1609,In_208,In_96);
nor U1610 (N_1610,In_914,In_782);
nand U1611 (N_1611,In_254,In_584);
nand U1612 (N_1612,In_714,In_547);
and U1613 (N_1613,In_320,In_472);
nor U1614 (N_1614,In_654,In_728);
or U1615 (N_1615,In_153,In_586);
and U1616 (N_1616,In_606,In_824);
nor U1617 (N_1617,In_326,In_504);
and U1618 (N_1618,In_563,In_348);
nand U1619 (N_1619,In_902,In_24);
nor U1620 (N_1620,In_885,In_694);
xnor U1621 (N_1621,In_275,In_83);
or U1622 (N_1622,In_683,In_655);
or U1623 (N_1623,In_235,In_817);
or U1624 (N_1624,In_787,In_893);
and U1625 (N_1625,In_217,In_938);
or U1626 (N_1626,In_591,In_723);
nor U1627 (N_1627,In_537,In_486);
nor U1628 (N_1628,In_767,In_558);
nand U1629 (N_1629,In_805,In_182);
nand U1630 (N_1630,In_477,In_503);
and U1631 (N_1631,In_55,In_751);
xor U1632 (N_1632,In_466,In_967);
nand U1633 (N_1633,In_592,In_865);
nand U1634 (N_1634,In_759,In_712);
nand U1635 (N_1635,In_991,In_776);
xor U1636 (N_1636,In_522,In_304);
nor U1637 (N_1637,In_730,In_757);
nor U1638 (N_1638,In_802,In_136);
nand U1639 (N_1639,In_992,In_930);
nand U1640 (N_1640,In_679,In_938);
nand U1641 (N_1641,In_80,In_841);
nor U1642 (N_1642,In_843,In_633);
and U1643 (N_1643,In_229,In_864);
and U1644 (N_1644,In_158,In_568);
or U1645 (N_1645,In_846,In_227);
nand U1646 (N_1646,In_898,In_86);
nand U1647 (N_1647,In_780,In_349);
nor U1648 (N_1648,In_752,In_524);
or U1649 (N_1649,In_479,In_909);
and U1650 (N_1650,In_666,In_180);
or U1651 (N_1651,In_941,In_89);
and U1652 (N_1652,In_777,In_458);
or U1653 (N_1653,In_268,In_329);
and U1654 (N_1654,In_376,In_34);
and U1655 (N_1655,In_431,In_235);
or U1656 (N_1656,In_186,In_801);
nor U1657 (N_1657,In_586,In_200);
nor U1658 (N_1658,In_118,In_625);
or U1659 (N_1659,In_823,In_838);
nor U1660 (N_1660,In_176,In_245);
and U1661 (N_1661,In_289,In_157);
or U1662 (N_1662,In_316,In_499);
or U1663 (N_1663,In_658,In_86);
or U1664 (N_1664,In_960,In_150);
or U1665 (N_1665,In_282,In_705);
or U1666 (N_1666,In_980,In_582);
nor U1667 (N_1667,In_258,In_468);
and U1668 (N_1668,In_97,In_575);
nand U1669 (N_1669,In_297,In_329);
xnor U1670 (N_1670,In_112,In_694);
or U1671 (N_1671,In_975,In_678);
or U1672 (N_1672,In_176,In_887);
and U1673 (N_1673,In_748,In_528);
nand U1674 (N_1674,In_626,In_376);
xor U1675 (N_1675,In_21,In_25);
nor U1676 (N_1676,In_471,In_482);
or U1677 (N_1677,In_952,In_570);
nand U1678 (N_1678,In_587,In_772);
nor U1679 (N_1679,In_130,In_900);
or U1680 (N_1680,In_147,In_109);
nor U1681 (N_1681,In_793,In_181);
nand U1682 (N_1682,In_41,In_750);
nor U1683 (N_1683,In_470,In_710);
and U1684 (N_1684,In_891,In_702);
and U1685 (N_1685,In_669,In_55);
nor U1686 (N_1686,In_965,In_166);
xor U1687 (N_1687,In_838,In_237);
nand U1688 (N_1688,In_565,In_789);
nand U1689 (N_1689,In_141,In_99);
xnor U1690 (N_1690,In_607,In_575);
or U1691 (N_1691,In_563,In_171);
nand U1692 (N_1692,In_414,In_267);
nand U1693 (N_1693,In_883,In_272);
nand U1694 (N_1694,In_219,In_392);
and U1695 (N_1695,In_628,In_411);
nand U1696 (N_1696,In_728,In_964);
nor U1697 (N_1697,In_562,In_379);
xor U1698 (N_1698,In_602,In_180);
xor U1699 (N_1699,In_789,In_532);
nor U1700 (N_1700,In_706,In_236);
nand U1701 (N_1701,In_552,In_135);
or U1702 (N_1702,In_907,In_728);
or U1703 (N_1703,In_686,In_235);
nor U1704 (N_1704,In_37,In_922);
or U1705 (N_1705,In_177,In_466);
and U1706 (N_1706,In_970,In_445);
and U1707 (N_1707,In_694,In_211);
nand U1708 (N_1708,In_830,In_705);
nand U1709 (N_1709,In_178,In_521);
nor U1710 (N_1710,In_989,In_714);
nor U1711 (N_1711,In_901,In_307);
nand U1712 (N_1712,In_373,In_999);
xor U1713 (N_1713,In_943,In_374);
or U1714 (N_1714,In_90,In_843);
xnor U1715 (N_1715,In_480,In_805);
or U1716 (N_1716,In_315,In_775);
nor U1717 (N_1717,In_53,In_479);
nor U1718 (N_1718,In_627,In_525);
nand U1719 (N_1719,In_909,In_5);
or U1720 (N_1720,In_780,In_261);
nand U1721 (N_1721,In_480,In_1);
and U1722 (N_1722,In_898,In_229);
nor U1723 (N_1723,In_419,In_765);
nand U1724 (N_1724,In_70,In_876);
or U1725 (N_1725,In_740,In_368);
nor U1726 (N_1726,In_916,In_242);
nor U1727 (N_1727,In_429,In_501);
and U1728 (N_1728,In_622,In_31);
nand U1729 (N_1729,In_849,In_696);
or U1730 (N_1730,In_323,In_763);
nor U1731 (N_1731,In_735,In_193);
nand U1732 (N_1732,In_444,In_501);
nor U1733 (N_1733,In_116,In_112);
or U1734 (N_1734,In_824,In_29);
and U1735 (N_1735,In_855,In_139);
and U1736 (N_1736,In_939,In_289);
or U1737 (N_1737,In_376,In_543);
or U1738 (N_1738,In_335,In_390);
nor U1739 (N_1739,In_304,In_367);
nor U1740 (N_1740,In_914,In_451);
or U1741 (N_1741,In_433,In_752);
xnor U1742 (N_1742,In_394,In_445);
and U1743 (N_1743,In_714,In_263);
or U1744 (N_1744,In_75,In_187);
and U1745 (N_1745,In_702,In_623);
nor U1746 (N_1746,In_207,In_592);
and U1747 (N_1747,In_293,In_462);
or U1748 (N_1748,In_616,In_278);
nand U1749 (N_1749,In_542,In_589);
nand U1750 (N_1750,In_381,In_891);
nor U1751 (N_1751,In_711,In_521);
nand U1752 (N_1752,In_705,In_315);
nand U1753 (N_1753,In_453,In_757);
and U1754 (N_1754,In_892,In_400);
or U1755 (N_1755,In_486,In_928);
or U1756 (N_1756,In_923,In_163);
or U1757 (N_1757,In_802,In_20);
nand U1758 (N_1758,In_368,In_946);
and U1759 (N_1759,In_639,In_687);
and U1760 (N_1760,In_586,In_286);
and U1761 (N_1761,In_567,In_974);
and U1762 (N_1762,In_430,In_135);
nand U1763 (N_1763,In_993,In_77);
nand U1764 (N_1764,In_103,In_742);
xor U1765 (N_1765,In_511,In_588);
nor U1766 (N_1766,In_257,In_924);
and U1767 (N_1767,In_239,In_657);
and U1768 (N_1768,In_46,In_276);
or U1769 (N_1769,In_301,In_853);
nor U1770 (N_1770,In_789,In_444);
or U1771 (N_1771,In_497,In_363);
nand U1772 (N_1772,In_692,In_757);
and U1773 (N_1773,In_551,In_649);
and U1774 (N_1774,In_555,In_312);
or U1775 (N_1775,In_840,In_191);
nand U1776 (N_1776,In_542,In_614);
nand U1777 (N_1777,In_760,In_614);
and U1778 (N_1778,In_82,In_544);
nor U1779 (N_1779,In_576,In_824);
xor U1780 (N_1780,In_871,In_856);
nand U1781 (N_1781,In_460,In_841);
nand U1782 (N_1782,In_42,In_85);
nand U1783 (N_1783,In_306,In_727);
nand U1784 (N_1784,In_300,In_204);
and U1785 (N_1785,In_949,In_748);
or U1786 (N_1786,In_375,In_71);
xor U1787 (N_1787,In_425,In_538);
and U1788 (N_1788,In_447,In_609);
or U1789 (N_1789,In_507,In_103);
nand U1790 (N_1790,In_888,In_63);
or U1791 (N_1791,In_27,In_982);
or U1792 (N_1792,In_925,In_324);
xor U1793 (N_1793,In_332,In_836);
and U1794 (N_1794,In_478,In_622);
nand U1795 (N_1795,In_174,In_92);
nor U1796 (N_1796,In_971,In_953);
nand U1797 (N_1797,In_405,In_602);
nor U1798 (N_1798,In_34,In_221);
nand U1799 (N_1799,In_646,In_889);
xnor U1800 (N_1800,In_254,In_865);
nor U1801 (N_1801,In_952,In_140);
nand U1802 (N_1802,In_308,In_270);
nor U1803 (N_1803,In_75,In_22);
and U1804 (N_1804,In_189,In_122);
nor U1805 (N_1805,In_665,In_174);
nand U1806 (N_1806,In_291,In_434);
xor U1807 (N_1807,In_402,In_433);
nand U1808 (N_1808,In_176,In_306);
nand U1809 (N_1809,In_396,In_320);
nor U1810 (N_1810,In_406,In_180);
nor U1811 (N_1811,In_994,In_85);
nand U1812 (N_1812,In_629,In_192);
nand U1813 (N_1813,In_368,In_461);
nor U1814 (N_1814,In_937,In_346);
nand U1815 (N_1815,In_500,In_679);
xor U1816 (N_1816,In_381,In_843);
nand U1817 (N_1817,In_616,In_98);
and U1818 (N_1818,In_189,In_453);
or U1819 (N_1819,In_803,In_718);
nor U1820 (N_1820,In_206,In_697);
nor U1821 (N_1821,In_260,In_954);
nand U1822 (N_1822,In_876,In_433);
and U1823 (N_1823,In_91,In_589);
xor U1824 (N_1824,In_468,In_176);
or U1825 (N_1825,In_283,In_721);
nor U1826 (N_1826,In_928,In_213);
and U1827 (N_1827,In_232,In_822);
or U1828 (N_1828,In_699,In_243);
nor U1829 (N_1829,In_316,In_180);
or U1830 (N_1830,In_395,In_93);
or U1831 (N_1831,In_473,In_920);
nor U1832 (N_1832,In_594,In_911);
or U1833 (N_1833,In_155,In_736);
nand U1834 (N_1834,In_849,In_474);
or U1835 (N_1835,In_982,In_320);
nand U1836 (N_1836,In_425,In_993);
nand U1837 (N_1837,In_832,In_607);
nor U1838 (N_1838,In_315,In_948);
nand U1839 (N_1839,In_781,In_411);
or U1840 (N_1840,In_425,In_503);
or U1841 (N_1841,In_916,In_244);
or U1842 (N_1842,In_998,In_142);
and U1843 (N_1843,In_721,In_620);
or U1844 (N_1844,In_307,In_883);
and U1845 (N_1845,In_374,In_259);
nand U1846 (N_1846,In_913,In_707);
or U1847 (N_1847,In_868,In_747);
or U1848 (N_1848,In_650,In_902);
or U1849 (N_1849,In_637,In_379);
and U1850 (N_1850,In_525,In_462);
nand U1851 (N_1851,In_323,In_916);
nand U1852 (N_1852,In_116,In_793);
xor U1853 (N_1853,In_598,In_701);
nand U1854 (N_1854,In_127,In_749);
nor U1855 (N_1855,In_681,In_28);
nor U1856 (N_1856,In_590,In_836);
xor U1857 (N_1857,In_247,In_599);
nor U1858 (N_1858,In_393,In_986);
and U1859 (N_1859,In_215,In_866);
or U1860 (N_1860,In_255,In_872);
xor U1861 (N_1861,In_113,In_891);
and U1862 (N_1862,In_349,In_710);
nand U1863 (N_1863,In_817,In_704);
nor U1864 (N_1864,In_671,In_820);
and U1865 (N_1865,In_554,In_407);
and U1866 (N_1866,In_495,In_666);
nand U1867 (N_1867,In_23,In_882);
or U1868 (N_1868,In_380,In_239);
and U1869 (N_1869,In_835,In_175);
nor U1870 (N_1870,In_899,In_730);
nand U1871 (N_1871,In_372,In_694);
or U1872 (N_1872,In_596,In_926);
and U1873 (N_1873,In_47,In_679);
nor U1874 (N_1874,In_465,In_636);
and U1875 (N_1875,In_793,In_707);
and U1876 (N_1876,In_767,In_399);
nand U1877 (N_1877,In_203,In_657);
nor U1878 (N_1878,In_223,In_393);
and U1879 (N_1879,In_264,In_392);
or U1880 (N_1880,In_932,In_237);
nor U1881 (N_1881,In_251,In_556);
or U1882 (N_1882,In_764,In_155);
or U1883 (N_1883,In_579,In_404);
nor U1884 (N_1884,In_875,In_824);
xor U1885 (N_1885,In_682,In_171);
xor U1886 (N_1886,In_484,In_191);
nand U1887 (N_1887,In_777,In_393);
and U1888 (N_1888,In_587,In_995);
nand U1889 (N_1889,In_798,In_136);
nand U1890 (N_1890,In_905,In_389);
and U1891 (N_1891,In_885,In_552);
nor U1892 (N_1892,In_194,In_871);
and U1893 (N_1893,In_294,In_313);
nand U1894 (N_1894,In_93,In_979);
nand U1895 (N_1895,In_408,In_165);
nand U1896 (N_1896,In_192,In_273);
nand U1897 (N_1897,In_139,In_346);
nand U1898 (N_1898,In_350,In_558);
and U1899 (N_1899,In_671,In_803);
nor U1900 (N_1900,In_365,In_379);
nor U1901 (N_1901,In_220,In_582);
and U1902 (N_1902,In_840,In_180);
and U1903 (N_1903,In_929,In_404);
and U1904 (N_1904,In_404,In_14);
or U1905 (N_1905,In_20,In_687);
nor U1906 (N_1906,In_454,In_693);
and U1907 (N_1907,In_588,In_209);
and U1908 (N_1908,In_180,In_621);
nor U1909 (N_1909,In_873,In_866);
xnor U1910 (N_1910,In_501,In_491);
and U1911 (N_1911,In_541,In_904);
nor U1912 (N_1912,In_83,In_272);
nand U1913 (N_1913,In_141,In_520);
or U1914 (N_1914,In_304,In_752);
nand U1915 (N_1915,In_469,In_63);
or U1916 (N_1916,In_781,In_250);
and U1917 (N_1917,In_432,In_897);
and U1918 (N_1918,In_10,In_715);
nor U1919 (N_1919,In_530,In_982);
xnor U1920 (N_1920,In_132,In_639);
and U1921 (N_1921,In_507,In_260);
and U1922 (N_1922,In_998,In_934);
nand U1923 (N_1923,In_856,In_991);
or U1924 (N_1924,In_746,In_148);
nand U1925 (N_1925,In_240,In_182);
nor U1926 (N_1926,In_876,In_33);
nor U1927 (N_1927,In_177,In_647);
or U1928 (N_1928,In_215,In_689);
or U1929 (N_1929,In_781,In_608);
nand U1930 (N_1930,In_387,In_879);
and U1931 (N_1931,In_836,In_613);
and U1932 (N_1932,In_406,In_12);
and U1933 (N_1933,In_508,In_496);
and U1934 (N_1934,In_341,In_314);
nand U1935 (N_1935,In_445,In_716);
nor U1936 (N_1936,In_365,In_438);
nand U1937 (N_1937,In_978,In_248);
and U1938 (N_1938,In_255,In_124);
nor U1939 (N_1939,In_739,In_214);
or U1940 (N_1940,In_788,In_261);
nand U1941 (N_1941,In_680,In_375);
and U1942 (N_1942,In_993,In_11);
nor U1943 (N_1943,In_401,In_70);
or U1944 (N_1944,In_135,In_576);
or U1945 (N_1945,In_516,In_993);
and U1946 (N_1946,In_994,In_327);
xor U1947 (N_1947,In_931,In_343);
or U1948 (N_1948,In_462,In_138);
xor U1949 (N_1949,In_520,In_183);
nor U1950 (N_1950,In_12,In_161);
nor U1951 (N_1951,In_906,In_877);
and U1952 (N_1952,In_928,In_151);
and U1953 (N_1953,In_699,In_862);
nor U1954 (N_1954,In_551,In_749);
xor U1955 (N_1955,In_177,In_987);
nor U1956 (N_1956,In_848,In_818);
and U1957 (N_1957,In_92,In_662);
or U1958 (N_1958,In_768,In_621);
xor U1959 (N_1959,In_638,In_130);
nor U1960 (N_1960,In_160,In_101);
and U1961 (N_1961,In_161,In_259);
and U1962 (N_1962,In_710,In_405);
or U1963 (N_1963,In_989,In_309);
or U1964 (N_1964,In_386,In_556);
nor U1965 (N_1965,In_307,In_945);
or U1966 (N_1966,In_0,In_544);
or U1967 (N_1967,In_858,In_515);
xor U1968 (N_1968,In_836,In_869);
or U1969 (N_1969,In_563,In_168);
xnor U1970 (N_1970,In_995,In_971);
nand U1971 (N_1971,In_910,In_136);
nand U1972 (N_1972,In_604,In_842);
nor U1973 (N_1973,In_185,In_426);
and U1974 (N_1974,In_972,In_505);
or U1975 (N_1975,In_76,In_329);
nand U1976 (N_1976,In_705,In_355);
nor U1977 (N_1977,In_97,In_167);
or U1978 (N_1978,In_465,In_619);
nand U1979 (N_1979,In_419,In_379);
nand U1980 (N_1980,In_357,In_636);
or U1981 (N_1981,In_949,In_899);
nand U1982 (N_1982,In_140,In_667);
nand U1983 (N_1983,In_425,In_273);
nor U1984 (N_1984,In_135,In_680);
or U1985 (N_1985,In_571,In_437);
and U1986 (N_1986,In_763,In_802);
or U1987 (N_1987,In_928,In_412);
or U1988 (N_1988,In_291,In_502);
or U1989 (N_1989,In_143,In_821);
nor U1990 (N_1990,In_524,In_571);
nor U1991 (N_1991,In_148,In_28);
nand U1992 (N_1992,In_593,In_36);
xnor U1993 (N_1993,In_997,In_927);
nand U1994 (N_1994,In_663,In_32);
or U1995 (N_1995,In_191,In_230);
nand U1996 (N_1996,In_946,In_246);
xnor U1997 (N_1997,In_602,In_993);
nor U1998 (N_1998,In_570,In_105);
and U1999 (N_1999,In_765,In_954);
nand U2000 (N_2000,N_81,N_66);
nand U2001 (N_2001,N_1647,N_39);
nor U2002 (N_2002,N_416,N_1283);
nand U2003 (N_2003,N_975,N_361);
and U2004 (N_2004,N_737,N_870);
nor U2005 (N_2005,N_1634,N_554);
or U2006 (N_2006,N_1556,N_449);
nand U2007 (N_2007,N_187,N_49);
and U2008 (N_2008,N_887,N_529);
and U2009 (N_2009,N_1029,N_1080);
xnor U2010 (N_2010,N_212,N_1434);
or U2011 (N_2011,N_597,N_1348);
and U2012 (N_2012,N_382,N_951);
nand U2013 (N_2013,N_323,N_1722);
nand U2014 (N_2014,N_396,N_479);
nand U2015 (N_2015,N_1162,N_1202);
nor U2016 (N_2016,N_1315,N_747);
and U2017 (N_2017,N_261,N_574);
nand U2018 (N_2018,N_367,N_1422);
and U2019 (N_2019,N_803,N_1973);
and U2020 (N_2020,N_694,N_1179);
nand U2021 (N_2021,N_1878,N_1065);
nand U2022 (N_2022,N_1277,N_582);
or U2023 (N_2023,N_674,N_14);
nand U2024 (N_2024,N_436,N_1494);
nor U2025 (N_2025,N_1511,N_161);
and U2026 (N_2026,N_431,N_1828);
nand U2027 (N_2027,N_989,N_1621);
nand U2028 (N_2028,N_755,N_616);
and U2029 (N_2029,N_1194,N_1792);
or U2030 (N_2030,N_1746,N_174);
nor U2031 (N_2031,N_498,N_189);
and U2032 (N_2032,N_1043,N_520);
or U2033 (N_2033,N_981,N_91);
nand U2034 (N_2034,N_1273,N_547);
nand U2035 (N_2035,N_896,N_1116);
and U2036 (N_2036,N_939,N_768);
or U2037 (N_2037,N_1107,N_205);
or U2038 (N_2038,N_1506,N_623);
and U2039 (N_2039,N_93,N_1223);
and U2040 (N_2040,N_1430,N_905);
and U2041 (N_2041,N_1762,N_822);
nor U2042 (N_2042,N_1682,N_105);
nand U2043 (N_2043,N_171,N_1954);
nand U2044 (N_2044,N_1894,N_341);
nand U2045 (N_2045,N_176,N_544);
and U2046 (N_2046,N_1299,N_1092);
nand U2047 (N_2047,N_415,N_511);
and U2048 (N_2048,N_1695,N_256);
nand U2049 (N_2049,N_1307,N_474);
or U2050 (N_2050,N_430,N_686);
nor U2051 (N_2051,N_1169,N_300);
and U2052 (N_2052,N_1504,N_1584);
xor U2053 (N_2053,N_762,N_1298);
and U2054 (N_2054,N_1612,N_603);
or U2055 (N_2055,N_1513,N_74);
or U2056 (N_2056,N_1890,N_677);
or U2057 (N_2057,N_245,N_1172);
nor U2058 (N_2058,N_802,N_76);
or U2059 (N_2059,N_336,N_232);
nor U2060 (N_2060,N_383,N_1440);
or U2061 (N_2061,N_858,N_1185);
nand U2062 (N_2062,N_628,N_593);
nor U2063 (N_2063,N_204,N_378);
or U2064 (N_2064,N_272,N_1909);
or U2065 (N_2065,N_118,N_913);
xor U2066 (N_2066,N_644,N_1702);
and U2067 (N_2067,N_751,N_867);
nand U2068 (N_2068,N_1940,N_1249);
or U2069 (N_2069,N_1139,N_1362);
nor U2070 (N_2070,N_297,N_304);
and U2071 (N_2071,N_1916,N_1062);
nor U2072 (N_2072,N_584,N_1183);
nand U2073 (N_2073,N_1675,N_830);
or U2074 (N_2074,N_1527,N_1641);
nor U2075 (N_2075,N_1170,N_1256);
nand U2076 (N_2076,N_1286,N_1195);
or U2077 (N_2077,N_1709,N_861);
or U2078 (N_2078,N_1731,N_1873);
and U2079 (N_2079,N_1876,N_1997);
nand U2080 (N_2080,N_1519,N_1849);
nor U2081 (N_2081,N_201,N_715);
and U2082 (N_2082,N_141,N_457);
or U2083 (N_2083,N_153,N_1189);
or U2084 (N_2084,N_1004,N_1555);
and U2085 (N_2085,N_1165,N_387);
nand U2086 (N_2086,N_286,N_71);
xor U2087 (N_2087,N_1693,N_1666);
nand U2088 (N_2088,N_190,N_303);
xor U2089 (N_2089,N_21,N_663);
nor U2090 (N_2090,N_1007,N_1685);
or U2091 (N_2091,N_1834,N_1732);
nand U2092 (N_2092,N_1129,N_1624);
nand U2093 (N_2093,N_735,N_257);
nor U2094 (N_2094,N_275,N_613);
or U2095 (N_2095,N_1192,N_281);
xor U2096 (N_2096,N_576,N_1599);
nor U2097 (N_2097,N_1774,N_513);
or U2098 (N_2098,N_1408,N_1854);
and U2099 (N_2099,N_1827,N_1445);
nor U2100 (N_2100,N_271,N_1901);
or U2101 (N_2101,N_1305,N_1370);
and U2102 (N_2102,N_1948,N_1386);
nand U2103 (N_2103,N_1163,N_1314);
and U2104 (N_2104,N_1285,N_866);
or U2105 (N_2105,N_1197,N_1627);
nand U2106 (N_2106,N_918,N_1775);
and U2107 (N_2107,N_799,N_505);
or U2108 (N_2108,N_1442,N_1008);
nand U2109 (N_2109,N_1233,N_881);
or U2110 (N_2110,N_706,N_1921);
xnor U2111 (N_2111,N_1770,N_495);
and U2112 (N_2112,N_1117,N_841);
xor U2113 (N_2113,N_740,N_1805);
nor U2114 (N_2114,N_1330,N_1843);
nor U2115 (N_2115,N_404,N_874);
or U2116 (N_2116,N_588,N_445);
nor U2117 (N_2117,N_984,N_859);
nand U2118 (N_2118,N_294,N_1399);
and U2119 (N_2119,N_689,N_259);
nor U2120 (N_2120,N_1159,N_481);
nand U2121 (N_2121,N_453,N_54);
nand U2122 (N_2122,N_773,N_305);
nand U2123 (N_2123,N_1595,N_252);
or U2124 (N_2124,N_1257,N_1410);
nand U2125 (N_2125,N_1164,N_1336);
and U2126 (N_2126,N_1747,N_1417);
nand U2127 (N_2127,N_1572,N_1491);
nor U2128 (N_2128,N_483,N_1467);
or U2129 (N_2129,N_1205,N_1905);
or U2130 (N_2130,N_1464,N_1303);
and U2131 (N_2131,N_1181,N_460);
nand U2132 (N_2132,N_825,N_1166);
xnor U2133 (N_2133,N_1985,N_195);
nor U2134 (N_2134,N_1715,N_301);
and U2135 (N_2135,N_691,N_813);
or U2136 (N_2136,N_1001,N_224);
nand U2137 (N_2137,N_1381,N_1187);
nand U2138 (N_2138,N_31,N_373);
or U2139 (N_2139,N_1881,N_1707);
and U2140 (N_2140,N_1911,N_1232);
or U2141 (N_2141,N_983,N_955);
xnor U2142 (N_2142,N_329,N_133);
xnor U2143 (N_2143,N_1540,N_393);
or U2144 (N_2144,N_1091,N_1448);
and U2145 (N_2145,N_309,N_23);
or U2146 (N_2146,N_247,N_35);
and U2147 (N_2147,N_169,N_1912);
or U2148 (N_2148,N_441,N_1874);
nor U2149 (N_2149,N_688,N_1790);
nand U2150 (N_2150,N_370,N_836);
nand U2151 (N_2151,N_1293,N_1637);
or U2152 (N_2152,N_1704,N_1568);
nor U2153 (N_2153,N_1373,N_1654);
nand U2154 (N_2154,N_1794,N_438);
nor U2155 (N_2155,N_1222,N_1796);
or U2156 (N_2156,N_758,N_104);
nand U2157 (N_2157,N_926,N_1489);
nor U2158 (N_2158,N_1193,N_375);
and U2159 (N_2159,N_1978,N_1284);
and U2160 (N_2160,N_708,N_3);
nand U2161 (N_2161,N_848,N_1152);
nand U2162 (N_2162,N_266,N_1917);
nor U2163 (N_2163,N_579,N_1272);
nor U2164 (N_2164,N_960,N_1860);
or U2165 (N_2165,N_1020,N_149);
nor U2166 (N_2166,N_173,N_1068);
and U2167 (N_2167,N_1863,N_692);
nand U2168 (N_2168,N_1856,N_319);
and U2169 (N_2169,N_413,N_1477);
or U2170 (N_2170,N_801,N_739);
nand U2171 (N_2171,N_1102,N_237);
or U2172 (N_2172,N_285,N_837);
or U2173 (N_2173,N_160,N_634);
and U2174 (N_2174,N_786,N_1302);
nor U2175 (N_2175,N_11,N_903);
nand U2176 (N_2176,N_371,N_463);
nor U2177 (N_2177,N_1657,N_60);
or U2178 (N_2178,N_163,N_325);
xnor U2179 (N_2179,N_1971,N_607);
and U2180 (N_2180,N_1419,N_1877);
xnor U2181 (N_2181,N_1653,N_1777);
and U2182 (N_2182,N_599,N_1301);
or U2183 (N_2183,N_542,N_716);
and U2184 (N_2184,N_374,N_386);
xor U2185 (N_2185,N_1771,N_103);
nor U2186 (N_2186,N_409,N_1480);
nand U2187 (N_2187,N_1734,N_1208);
or U2188 (N_2188,N_695,N_273);
and U2189 (N_2189,N_1590,N_967);
nand U2190 (N_2190,N_243,N_1787);
nand U2191 (N_2191,N_736,N_203);
or U2192 (N_2192,N_864,N_170);
and U2193 (N_2193,N_1236,N_317);
nand U2194 (N_2194,N_1264,N_733);
xor U2195 (N_2195,N_518,N_1282);
and U2196 (N_2196,N_1939,N_392);
xor U2197 (N_2197,N_1017,N_1880);
and U2198 (N_2198,N_1825,N_1462);
or U2199 (N_2199,N_1030,N_696);
nor U2200 (N_2200,N_1173,N_372);
nand U2201 (N_2201,N_1237,N_1871);
and U2202 (N_2202,N_1869,N_45);
and U2203 (N_2203,N_1644,N_1743);
nand U2204 (N_2204,N_1493,N_1528);
nand U2205 (N_2205,N_316,N_687);
and U2206 (N_2206,N_1300,N_322);
nor U2207 (N_2207,N_503,N_1550);
or U2208 (N_2208,N_1230,N_1235);
nor U2209 (N_2209,N_454,N_1801);
or U2210 (N_2210,N_888,N_1735);
or U2211 (N_2211,N_1943,N_1663);
and U2212 (N_2212,N_834,N_1804);
or U2213 (N_2213,N_1549,N_1913);
and U2214 (N_2214,N_214,N_1212);
or U2215 (N_2215,N_1821,N_440);
xnor U2216 (N_2216,N_1466,N_1615);
or U2217 (N_2217,N_643,N_539);
nand U2218 (N_2218,N_397,N_1706);
or U2219 (N_2219,N_1168,N_1295);
nor U2220 (N_2220,N_365,N_1274);
and U2221 (N_2221,N_1126,N_1182);
and U2222 (N_2222,N_1186,N_700);
and U2223 (N_2223,N_1137,N_1724);
nor U2224 (N_2224,N_1639,N_0);
nor U2225 (N_2225,N_673,N_1941);
and U2226 (N_2226,N_223,N_945);
nor U2227 (N_2227,N_1523,N_1651);
nor U2228 (N_2228,N_1064,N_1498);
nor U2229 (N_2229,N_1345,N_883);
xor U2230 (N_2230,N_433,N_804);
and U2231 (N_2231,N_985,N_43);
nand U2232 (N_2232,N_1852,N_1956);
and U2233 (N_2233,N_1155,N_1269);
or U2234 (N_2234,N_541,N_270);
and U2235 (N_2235,N_472,N_1228);
nor U2236 (N_2236,N_527,N_240);
nor U2237 (N_2237,N_127,N_1247);
nor U2238 (N_2238,N_954,N_1320);
or U2239 (N_2239,N_1026,N_949);
nor U2240 (N_2240,N_1616,N_1986);
and U2241 (N_2241,N_756,N_295);
nand U2242 (N_2242,N_1914,N_1142);
or U2243 (N_2243,N_936,N_875);
nand U2244 (N_2244,N_34,N_1167);
and U2245 (N_2245,N_660,N_215);
nor U2246 (N_2246,N_1557,N_324);
nor U2247 (N_2247,N_192,N_868);
and U2248 (N_2248,N_1395,N_1454);
nor U2249 (N_2249,N_1723,N_1470);
nor U2250 (N_2250,N_142,N_197);
nor U2251 (N_2251,N_509,N_501);
and U2252 (N_2252,N_1520,N_342);
nand U2253 (N_2253,N_519,N_1413);
nand U2254 (N_2254,N_143,N_1347);
nand U2255 (N_2255,N_1688,N_750);
or U2256 (N_2256,N_1058,N_1936);
or U2257 (N_2257,N_1388,N_1539);
nand U2258 (N_2258,N_467,N_1350);
or U2259 (N_2259,N_1079,N_471);
nand U2260 (N_2260,N_1502,N_1810);
nand U2261 (N_2261,N_1631,N_1180);
nand U2262 (N_2262,N_186,N_1623);
nand U2263 (N_2263,N_1865,N_265);
or U2264 (N_2264,N_890,N_635);
xor U2265 (N_2265,N_1552,N_1133);
nand U2266 (N_2266,N_1526,N_831);
nand U2267 (N_2267,N_1327,N_598);
nand U2268 (N_2268,N_1902,N_1886);
nand U2269 (N_2269,N_648,N_183);
nor U2270 (N_2270,N_1541,N_899);
or U2271 (N_2271,N_172,N_988);
nand U2272 (N_2272,N_20,N_246);
nand U2273 (N_2273,N_1,N_1346);
or U2274 (N_2274,N_1945,N_1051);
nor U2275 (N_2275,N_850,N_1281);
and U2276 (N_2276,N_1038,N_1371);
nand U2277 (N_2277,N_707,N_1759);
nand U2278 (N_2278,N_1361,N_617);
or U2279 (N_2279,N_1240,N_991);
nor U2280 (N_2280,N_879,N_1027);
and U2281 (N_2281,N_1571,N_610);
nor U2282 (N_2282,N_1110,N_1472);
or U2283 (N_2283,N_28,N_140);
and U2284 (N_2284,N_957,N_928);
and U2285 (N_2285,N_1992,N_502);
xor U2286 (N_2286,N_1221,N_1904);
nand U2287 (N_2287,N_1955,N_924);
nor U2288 (N_2288,N_512,N_1143);
and U2289 (N_2289,N_846,N_1401);
nor U2290 (N_2290,N_1593,N_434);
nor U2291 (N_2291,N_1045,N_729);
nor U2292 (N_2292,N_1251,N_1716);
or U2293 (N_2293,N_1545,N_863);
or U2294 (N_2294,N_22,N_1781);
or U2295 (N_2295,N_565,N_1501);
and U2296 (N_2296,N_1628,N_1060);
nor U2297 (N_2297,N_10,N_893);
xnor U2298 (N_2298,N_1835,N_249);
and U2299 (N_2299,N_684,N_1206);
nand U2300 (N_2300,N_1132,N_1354);
and U2301 (N_2301,N_973,N_820);
nand U2302 (N_2302,N_260,N_1112);
nand U2303 (N_2303,N_1744,N_1814);
nand U2304 (N_2304,N_532,N_1924);
xnor U2305 (N_2305,N_1636,N_1614);
or U2306 (N_2306,N_466,N_395);
and U2307 (N_2307,N_522,N_1211);
nand U2308 (N_2308,N_32,N_1328);
nor U2309 (N_2309,N_1578,N_668);
nand U2310 (N_2310,N_184,N_1765);
nand U2311 (N_2311,N_485,N_1889);
xnor U2312 (N_2312,N_1691,N_37);
nand U2313 (N_2313,N_581,N_840);
nand U2314 (N_2314,N_721,N_390);
nor U2315 (N_2315,N_1783,N_1988);
or U2316 (N_2316,N_571,N_1560);
and U2317 (N_2317,N_1149,N_727);
nor U2318 (N_2318,N_376,N_1398);
nor U2319 (N_2319,N_196,N_182);
xnor U2320 (N_2320,N_1608,N_258);
nand U2321 (N_2321,N_1296,N_606);
nor U2322 (N_2322,N_377,N_227);
or U2323 (N_2323,N_909,N_406);
xor U2324 (N_2324,N_1406,N_30);
nor U2325 (N_2325,N_1671,N_262);
or U2326 (N_2326,N_1974,N_1218);
nor U2327 (N_2327,N_158,N_1566);
and U2328 (N_2328,N_191,N_1738);
or U2329 (N_2329,N_1859,N_987);
nand U2330 (N_2330,N_1515,N_1946);
nor U2331 (N_2331,N_1196,N_1309);
and U2332 (N_2332,N_1244,N_1275);
nor U2333 (N_2333,N_1500,N_58);
xnor U2334 (N_2334,N_1714,N_860);
and U2335 (N_2335,N_155,N_1229);
nand U2336 (N_2336,N_1459,N_1819);
and U2337 (N_2337,N_676,N_911);
and U2338 (N_2338,N_1369,N_889);
nand U2339 (N_2339,N_1598,N_1358);
xor U2340 (N_2340,N_1620,N_92);
or U2341 (N_2341,N_405,N_202);
and U2342 (N_2342,N_1418,N_50);
or U2343 (N_2343,N_1958,N_1503);
nor U2344 (N_2344,N_1042,N_1851);
nand U2345 (N_2345,N_748,N_106);
and U2346 (N_2346,N_812,N_1323);
nand U2347 (N_2347,N_937,N_146);
or U2348 (N_2348,N_1514,N_1591);
and U2349 (N_2349,N_1692,N_885);
and U2350 (N_2350,N_1150,N_181);
nor U2351 (N_2351,N_1482,N_675);
nand U2352 (N_2352,N_1570,N_269);
or U2353 (N_2353,N_1360,N_1339);
nor U2354 (N_2354,N_19,N_771);
or U2355 (N_2355,N_1950,N_1587);
and U2356 (N_2356,N_915,N_1534);
nor U2357 (N_2357,N_1516,N_274);
or U2358 (N_2358,N_1238,N_681);
nand U2359 (N_2359,N_1147,N_326);
nand U2360 (N_2360,N_877,N_1375);
and U2361 (N_2361,N_282,N_1075);
or U2362 (N_2362,N_1959,N_468);
nand U2363 (N_2363,N_907,N_978);
and U2364 (N_2364,N_1791,N_1089);
xor U2365 (N_2365,N_852,N_226);
nor U2366 (N_2366,N_816,N_88);
and U2367 (N_2367,N_455,N_111);
nand U2368 (N_2368,N_1450,N_1435);
and U2369 (N_2369,N_1357,N_683);
and U2370 (N_2370,N_1310,N_1121);
and U2371 (N_2371,N_83,N_220);
nor U2372 (N_2372,N_447,N_1908);
or U2373 (N_2373,N_1766,N_1983);
nor U2374 (N_2374,N_1306,N_1177);
nand U2375 (N_2375,N_423,N_1262);
and U2376 (N_2376,N_1488,N_1972);
nor U2377 (N_2377,N_562,N_1594);
nand U2378 (N_2378,N_1903,N_459);
or U2379 (N_2379,N_596,N_1405);
or U2380 (N_2380,N_963,N_1100);
nand U2381 (N_2381,N_1829,N_1046);
xnor U2382 (N_2382,N_1764,N_1508);
and U2383 (N_2383,N_1311,N_1967);
or U2384 (N_2384,N_59,N_1319);
nor U2385 (N_2385,N_1832,N_1547);
xor U2386 (N_2386,N_280,N_724);
nor U2387 (N_2387,N_546,N_1532);
nand U2388 (N_2388,N_307,N_814);
nand U2389 (N_2389,N_948,N_806);
nor U2390 (N_2390,N_794,N_1260);
nand U2391 (N_2391,N_97,N_1469);
nand U2392 (N_2392,N_1853,N_1773);
and U2393 (N_2393,N_1824,N_1003);
and U2394 (N_2394,N_389,N_591);
or U2395 (N_2395,N_1308,N_1248);
nand U2396 (N_2396,N_388,N_847);
nor U2397 (N_2397,N_458,N_46);
nor U2398 (N_2398,N_1022,N_1136);
xor U2399 (N_2399,N_710,N_898);
nor U2400 (N_2400,N_997,N_1700);
nand U2401 (N_2401,N_38,N_96);
nor U2402 (N_2402,N_1861,N_151);
and U2403 (N_2403,N_1922,N_250);
nand U2404 (N_2404,N_135,N_1341);
nor U2405 (N_2405,N_1752,N_1717);
nand U2406 (N_2406,N_817,N_1161);
nand U2407 (N_2407,N_953,N_1658);
or U2408 (N_2408,N_1586,N_567);
nor U2409 (N_2409,N_934,N_369);
or U2410 (N_2410,N_4,N_1243);
nor U2411 (N_2411,N_177,N_1648);
and U2412 (N_2412,N_1455,N_651);
and U2413 (N_2413,N_279,N_1982);
xor U2414 (N_2414,N_862,N_1915);
and U2415 (N_2415,N_1949,N_1481);
nor U2416 (N_2416,N_337,N_491);
nand U2417 (N_2417,N_435,N_1577);
nand U2418 (N_2418,N_1674,N_366);
and U2419 (N_2419,N_1333,N_992);
xnor U2420 (N_2420,N_523,N_276);
nand U2421 (N_2421,N_283,N_53);
or U2422 (N_2422,N_1589,N_996);
nor U2423 (N_2423,N_1242,N_1120);
and U2424 (N_2424,N_1077,N_633);
and U2425 (N_2425,N_549,N_1645);
nor U2426 (N_2426,N_531,N_1934);
or U2427 (N_2427,N_1573,N_120);
nor U2428 (N_2428,N_335,N_8);
xor U2429 (N_2429,N_931,N_1499);
and U2430 (N_2430,N_944,N_5);
nand U2431 (N_2431,N_1602,N_1517);
nor U2432 (N_2432,N_1882,N_52);
and U2433 (N_2433,N_1505,N_1471);
nor U2434 (N_2434,N_656,N_332);
or U2435 (N_2435,N_537,N_1963);
nand U2436 (N_2436,N_1893,N_941);
or U2437 (N_2437,N_752,N_1431);
nor U2438 (N_2438,N_1453,N_1414);
nand U2439 (N_2439,N_1191,N_1190);
nor U2440 (N_2440,N_615,N_1225);
and U2441 (N_2441,N_452,N_1681);
nand U2442 (N_2442,N_1739,N_1581);
and U2443 (N_2443,N_101,N_334);
or U2444 (N_2444,N_1118,N_1457);
nand U2445 (N_2445,N_632,N_1288);
or U2446 (N_2446,N_15,N_580);
nand U2447 (N_2447,N_1837,N_553);
or U2448 (N_2448,N_1368,N_344);
or U2449 (N_2449,N_166,N_1312);
or U2450 (N_2450,N_791,N_1846);
or U2451 (N_2451,N_1778,N_1763);
or U2452 (N_2452,N_175,N_1543);
nor U2453 (N_2453,N_346,N_132);
nor U2454 (N_2454,N_312,N_1394);
nor U2455 (N_2455,N_1246,N_152);
or U2456 (N_2456,N_601,N_1793);
and U2457 (N_2457,N_583,N_1660);
nor U2458 (N_2458,N_1727,N_102);
nor U2459 (N_2459,N_1324,N_1449);
nand U2460 (N_2460,N_1990,N_1101);
nand U2461 (N_2461,N_1561,N_1468);
nor U2462 (N_2462,N_230,N_1562);
and U2463 (N_2463,N_1403,N_411);
and U2464 (N_2464,N_1965,N_1780);
or U2465 (N_2465,N_1151,N_1011);
or U2466 (N_2466,N_891,N_775);
xnor U2467 (N_2467,N_637,N_886);
and U2468 (N_2468,N_1554,N_772);
nor U2469 (N_2469,N_400,N_718);
and U2470 (N_2470,N_1153,N_1872);
nand U2471 (N_2471,N_1900,N_2);
nand U2472 (N_2472,N_595,N_1396);
nand U2473 (N_2473,N_979,N_705);
nand U2474 (N_2474,N_1217,N_338);
nor U2475 (N_2475,N_1684,N_225);
nand U2476 (N_2476,N_1032,N_1962);
nand U2477 (N_2477,N_1119,N_95);
and U2478 (N_2478,N_1753,N_1437);
nand U2479 (N_2479,N_1898,N_1538);
or U2480 (N_2480,N_1475,N_1384);
nand U2481 (N_2481,N_704,N_154);
and U2482 (N_2482,N_1106,N_587);
nand U2483 (N_2483,N_164,N_80);
or U2484 (N_2484,N_561,N_1376);
or U2485 (N_2485,N_770,N_1977);
nor U2486 (N_2486,N_855,N_109);
or U2487 (N_2487,N_1929,N_1583);
or U2488 (N_2488,N_1887,N_938);
nand U2489 (N_2489,N_1148,N_1559);
nor U2490 (N_2490,N_1638,N_429);
or U2491 (N_2491,N_178,N_1789);
and U2492 (N_2492,N_1096,N_1407);
nand U2493 (N_2493,N_311,N_641);
xor U2494 (N_2494,N_962,N_1465);
nor U2495 (N_2495,N_1108,N_545);
nand U2496 (N_2496,N_255,N_356);
nor U2497 (N_2497,N_1680,N_1446);
and U2498 (N_2498,N_1823,N_1385);
and U2499 (N_2499,N_108,N_559);
nand U2500 (N_2500,N_1725,N_1234);
and U2501 (N_2501,N_1048,N_1643);
and U2502 (N_2502,N_661,N_499);
nor U2503 (N_2503,N_1822,N_1580);
nand U2504 (N_2504,N_680,N_1600);
or U2505 (N_2505,N_880,N_1012);
nand U2506 (N_2506,N_1683,N_167);
and U2507 (N_2507,N_1712,N_1979);
nand U2508 (N_2508,N_1316,N_469);
nor U2509 (N_2509,N_357,N_16);
nor U2510 (N_2510,N_292,N_6);
and U2511 (N_2511,N_1910,N_41);
nor U2512 (N_2512,N_604,N_605);
nand U2513 (N_2513,N_744,N_1087);
and U2514 (N_2514,N_1617,N_1458);
and U2515 (N_2515,N_980,N_221);
nand U2516 (N_2516,N_698,N_1099);
or U2517 (N_2517,N_1390,N_703);
nand U2518 (N_2518,N_1767,N_350);
nand U2519 (N_2519,N_1122,N_125);
nand U2520 (N_2520,N_573,N_1741);
or U2521 (N_2521,N_609,N_1996);
and U2522 (N_2522,N_793,N_1411);
nor U2523 (N_2523,N_277,N_516);
nor U2524 (N_2524,N_1803,N_1718);
nand U2525 (N_2525,N_1066,N_379);
or U2526 (N_2526,N_760,N_1207);
nor U2527 (N_2527,N_1097,N_464);
nand U2528 (N_2528,N_476,N_779);
and U2529 (N_2529,N_1925,N_1622);
nor U2530 (N_2530,N_443,N_1613);
nor U2531 (N_2531,N_1981,N_1784);
or U2532 (N_2532,N_1531,N_1597);
nand U2533 (N_2533,N_1071,N_1176);
nand U2534 (N_2534,N_1426,N_572);
and U2535 (N_2535,N_1374,N_1367);
or U2536 (N_2536,N_1070,N_1157);
nand U2537 (N_2537,N_461,N_1574);
and U2538 (N_2538,N_1184,N_1496);
or U2539 (N_2539,N_110,N_1433);
nand U2540 (N_2540,N_40,N_514);
or U2541 (N_2541,N_894,N_1630);
nand U2542 (N_2542,N_1899,N_48);
nor U2543 (N_2543,N_550,N_1690);
nor U2544 (N_2544,N_1885,N_1198);
nor U2545 (N_2545,N_872,N_119);
nor U2546 (N_2546,N_1209,N_1201);
or U2547 (N_2547,N_222,N_776);
or U2548 (N_2548,N_1605,N_1429);
xor U2549 (N_2549,N_533,N_1987);
nor U2550 (N_2550,N_1659,N_1947);
or U2551 (N_2551,N_1130,N_1378);
nand U2552 (N_2552,N_1086,N_1123);
nand U2553 (N_2553,N_506,N_198);
nand U2554 (N_2554,N_391,N_835);
nor U2555 (N_2555,N_484,N_1145);
nor U2556 (N_2556,N_1579,N_1994);
and U2557 (N_2557,N_313,N_1664);
nor U2558 (N_2558,N_974,N_815);
and U2559 (N_2559,N_971,N_1510);
nor U2560 (N_2560,N_1171,N_12);
and U2561 (N_2561,N_819,N_210);
or U2562 (N_2562,N_589,N_1072);
or U2563 (N_2563,N_757,N_62);
nor U2564 (N_2564,N_1000,N_1267);
nand U2565 (N_2565,N_73,N_1334);
xnor U2566 (N_2566,N_1318,N_1085);
or U2567 (N_2567,N_851,N_394);
nand U2568 (N_2568,N_555,N_320);
and U2569 (N_2569,N_1720,N_381);
and U2570 (N_2570,N_1975,N_1351);
nor U2571 (N_2571,N_854,N_871);
and U2572 (N_2572,N_358,N_1331);
or U2573 (N_2573,N_1024,N_263);
or U2574 (N_2574,N_551,N_1231);
nor U2575 (N_2575,N_69,N_897);
or U2576 (N_2576,N_1969,N_1490);
and U2577 (N_2577,N_958,N_1479);
xnor U2578 (N_2578,N_1563,N_556);
and U2579 (N_2579,N_1463,N_856);
or U2580 (N_2580,N_299,N_1276);
or U2581 (N_2581,N_1061,N_420);
nand U2582 (N_2582,N_1175,N_950);
xor U2583 (N_2583,N_659,N_809);
and U2584 (N_2584,N_792,N_185);
or U2585 (N_2585,N_1268,N_536);
and U2586 (N_2586,N_1779,N_1291);
xor U2587 (N_2587,N_1564,N_353);
and U2588 (N_2588,N_489,N_1278);
nor U2589 (N_2589,N_57,N_667);
nand U2590 (N_2590,N_842,N_1329);
and U2591 (N_2591,N_575,N_1428);
nor U2592 (N_2592,N_1633,N_1676);
or U2593 (N_2593,N_340,N_1073);
nand U2594 (N_2594,N_51,N_693);
nor U2595 (N_2595,N_725,N_1055);
or U2596 (N_2596,N_1920,N_1942);
or U2597 (N_2597,N_493,N_233);
or U2598 (N_2598,N_1014,N_1487);
nand U2599 (N_2599,N_1239,N_1326);
nand U2600 (N_2600,N_844,N_67);
or U2601 (N_2601,N_577,N_401);
or U2602 (N_2602,N_1632,N_1655);
nor U2603 (N_2603,N_1918,N_253);
xnor U2604 (N_2604,N_1124,N_720);
nor U2605 (N_2605,N_642,N_672);
nor U2606 (N_2606,N_722,N_1952);
nand U2607 (N_2607,N_612,N_1726);
nand U2608 (N_2608,N_235,N_1382);
nand U2609 (N_2609,N_1040,N_1868);
xor U2610 (N_2610,N_349,N_1095);
and U2611 (N_2611,N_933,N_821);
or U2612 (N_2612,N_1670,N_1146);
nor U2613 (N_2613,N_27,N_1292);
nor U2614 (N_2614,N_920,N_1270);
nand U2615 (N_2615,N_1576,N_1667);
xor U2616 (N_2616,N_1751,N_1729);
or U2617 (N_2617,N_649,N_1817);
or U2618 (N_2618,N_1364,N_1606);
or U2619 (N_2619,N_1864,N_1018);
and U2620 (N_2620,N_828,N_769);
and U2621 (N_2621,N_1355,N_1069);
or U2622 (N_2622,N_437,N_1844);
and U2623 (N_2623,N_1642,N_1551);
xnor U2624 (N_2624,N_1575,N_664);
and U2625 (N_2625,N_845,N_26);
or U2626 (N_2626,N_1421,N_884);
xnor U2627 (N_2627,N_1366,N_1255);
nand U2628 (N_2628,N_560,N_1544);
and U2629 (N_2629,N_123,N_1036);
and U2630 (N_2630,N_902,N_994);
nand U2631 (N_2631,N_1415,N_1776);
nor U2632 (N_2632,N_1850,N_327);
and U2633 (N_2633,N_1443,N_917);
and U2634 (N_2634,N_627,N_662);
or U2635 (N_2635,N_1363,N_1976);
xnor U2636 (N_2636,N_1635,N_77);
xor U2637 (N_2637,N_1203,N_1798);
nand U2638 (N_2638,N_557,N_800);
nor U2639 (N_2639,N_636,N_1839);
nand U2640 (N_2640,N_1609,N_1926);
nand U2641 (N_2641,N_208,N_1297);
xnor U2642 (N_2642,N_1451,N_795);
nor U2643 (N_2643,N_1409,N_594);
nor U2644 (N_2644,N_921,N_1769);
nor U2645 (N_2645,N_1290,N_1078);
or U2646 (N_2646,N_1931,N_1050);
nor U2647 (N_2647,N_788,N_1105);
nor U2648 (N_2648,N_25,N_1678);
and U2649 (N_2649,N_1094,N_1485);
nand U2650 (N_2650,N_29,N_645);
nor U2651 (N_2651,N_1325,N_1416);
nor U2652 (N_2652,N_1447,N_1322);
or U2653 (N_2653,N_530,N_1855);
xnor U2654 (N_2654,N_1289,N_478);
xnor U2655 (N_2655,N_1953,N_1858);
nor U2656 (N_2656,N_728,N_1215);
and U2657 (N_2657,N_148,N_807);
nor U2658 (N_2658,N_1047,N_1626);
or U2659 (N_2659,N_1423,N_55);
nand U2660 (N_2660,N_1507,N_1806);
nand U2661 (N_2661,N_159,N_1999);
nor U2662 (N_2662,N_766,N_726);
nor U2663 (N_2663,N_600,N_650);
or U2664 (N_2664,N_218,N_968);
xnor U2665 (N_2665,N_1037,N_1474);
and U2666 (N_2666,N_288,N_646);
nor U2667 (N_2667,N_1760,N_36);
nor U2668 (N_2668,N_1857,N_1059);
or U2669 (N_2669,N_787,N_1698);
nand U2670 (N_2670,N_1818,N_1740);
nand U2671 (N_2671,N_168,N_1109);
nor U2672 (N_2672,N_1696,N_1907);
nand U2673 (N_2673,N_1052,N_1529);
nand U2674 (N_2674,N_1728,N_291);
or U2675 (N_2675,N_194,N_510);
nand U2676 (N_2676,N_570,N_1697);
nor U2677 (N_2677,N_1677,N_1668);
nor U2678 (N_2678,N_412,N_42);
or U2679 (N_2679,N_333,N_1313);
nor U2680 (N_2680,N_1968,N_1128);
and U2681 (N_2681,N_655,N_1009);
or U2682 (N_2682,N_829,N_1842);
nor U2683 (N_2683,N_124,N_289);
nor U2684 (N_2684,N_1013,N_1054);
or U2685 (N_2685,N_1807,N_1879);
and U2686 (N_2686,N_734,N_1755);
nor U2687 (N_2687,N_1473,N_742);
or U2688 (N_2688,N_473,N_47);
and U2689 (N_2689,N_139,N_339);
nor U2690 (N_2690,N_785,N_1082);
nand U2691 (N_2691,N_1933,N_9);
nor U2692 (N_2692,N_1758,N_488);
or U2693 (N_2693,N_697,N_1536);
and U2694 (N_2694,N_137,N_314);
or U2695 (N_2695,N_916,N_293);
nand U2696 (N_2696,N_1216,N_843);
or U2697 (N_2697,N_1135,N_330);
or U2698 (N_2698,N_1984,N_568);
or U2699 (N_2699,N_699,N_87);
and U2700 (N_2700,N_1456,N_1178);
nand U2701 (N_2701,N_1439,N_1812);
or U2702 (N_2702,N_1057,N_116);
xnor U2703 (N_2703,N_86,N_1033);
nand U2704 (N_2704,N_1028,N_1548);
nor U2705 (N_2705,N_543,N_126);
nand U2706 (N_2706,N_763,N_638);
nor U2707 (N_2707,N_1436,N_943);
and U2708 (N_2708,N_242,N_990);
or U2709 (N_2709,N_156,N_1710);
nand U2710 (N_2710,N_1897,N_1044);
nor U2711 (N_2711,N_993,N_180);
nand U2712 (N_2712,N_1701,N_1379);
or U2713 (N_2713,N_354,N_1224);
xor U2714 (N_2714,N_113,N_569);
or U2715 (N_2715,N_33,N_1111);
or U2716 (N_2716,N_1441,N_315);
xor U2717 (N_2717,N_999,N_1689);
nand U2718 (N_2718,N_504,N_362);
xor U2719 (N_2719,N_1125,N_462);
nor U2720 (N_2720,N_363,N_1749);
nor U2721 (N_2721,N_1134,N_1960);
nor U2722 (N_2722,N_932,N_1719);
xor U2723 (N_2723,N_1067,N_1896);
nand U2724 (N_2724,N_1432,N_1588);
nor U2725 (N_2725,N_679,N_810);
and U2726 (N_2726,N_538,N_590);
nand U2727 (N_2727,N_1103,N_1204);
nand U2728 (N_2728,N_497,N_969);
nor U2729 (N_2729,N_1756,N_1083);
nor U2730 (N_2730,N_925,N_384);
xnor U2731 (N_2731,N_13,N_1400);
nand U2732 (N_2732,N_1241,N_1352);
nand U2733 (N_2733,N_608,N_1815);
nand U2734 (N_2734,N_1757,N_654);
nor U2735 (N_2735,N_1220,N_1964);
nand U2736 (N_2736,N_402,N_1174);
xnor U2737 (N_2737,N_206,N_107);
xor U2738 (N_2738,N_1019,N_964);
and U2739 (N_2739,N_1596,N_231);
xnor U2740 (N_2740,N_1006,N_1265);
nor U2741 (N_2741,N_68,N_1687);
nor U2742 (N_2742,N_216,N_345);
or U2743 (N_2743,N_1640,N_566);
and U2744 (N_2744,N_61,N_1672);
nor U2745 (N_2745,N_1279,N_1063);
and U2746 (N_2746,N_1786,N_150);
nand U2747 (N_2747,N_1254,N_626);
and U2748 (N_2748,N_98,N_558);
and U2749 (N_2749,N_712,N_239);
and U2750 (N_2750,N_1646,N_136);
nor U2751 (N_2751,N_228,N_1144);
and U2752 (N_2752,N_268,N_157);
xnor U2753 (N_2753,N_906,N_901);
nand U2754 (N_2754,N_1601,N_1788);
or U2755 (N_2755,N_1816,N_439);
or U2756 (N_2756,N_1686,N_895);
and U2757 (N_2757,N_1840,N_162);
and U2758 (N_2758,N_833,N_1377);
and U2759 (N_2759,N_1761,N_1845);
nand U2760 (N_2760,N_1745,N_1966);
or U2761 (N_2761,N_1733,N_970);
and U2762 (N_2762,N_1833,N_1213);
nand U2763 (N_2763,N_236,N_818);
nor U2764 (N_2764,N_492,N_360);
nor U2765 (N_2765,N_620,N_79);
or U2766 (N_2766,N_1402,N_1391);
nor U2767 (N_2767,N_811,N_1343);
or U2768 (N_2768,N_238,N_702);
nor U2769 (N_2769,N_1957,N_1611);
and U2770 (N_2770,N_1261,N_1665);
nand U2771 (N_2771,N_1372,N_690);
nand U2772 (N_2772,N_956,N_428);
or U2773 (N_2773,N_1392,N_1604);
and U2774 (N_2774,N_714,N_75);
nor U2775 (N_2775,N_424,N_1081);
nand U2776 (N_2776,N_129,N_1875);
nor U2777 (N_2777,N_1025,N_1484);
nor U2778 (N_2778,N_1795,N_1650);
and U2779 (N_2779,N_629,N_1495);
and U2780 (N_2780,N_487,N_1989);
nor U2781 (N_2781,N_229,N_827);
nand U2782 (N_2782,N_1393,N_1830);
nor U2783 (N_2783,N_912,N_421);
nor U2784 (N_2784,N_1380,N_639);
nand U2785 (N_2785,N_1772,N_540);
and U2786 (N_2786,N_1031,N_732);
and U2787 (N_2787,N_248,N_7);
or U2788 (N_2788,N_1754,N_1619);
nor U2789 (N_2789,N_1652,N_701);
and U2790 (N_2790,N_432,N_1546);
nor U2791 (N_2791,N_796,N_1138);
or U2792 (N_2792,N_1919,N_1883);
and U2793 (N_2793,N_1098,N_347);
nand U2794 (N_2794,N_1188,N_1245);
nand U2795 (N_2795,N_998,N_1699);
and U2796 (N_2796,N_1927,N_930);
xor U2797 (N_2797,N_241,N_534);
or U2798 (N_2798,N_207,N_417);
nor U2799 (N_2799,N_1160,N_652);
or U2800 (N_2800,N_1093,N_1524);
and U2801 (N_2801,N_745,N_264);
and U2802 (N_2802,N_500,N_1928);
and U2803 (N_2803,N_961,N_1076);
nand U2804 (N_2804,N_1585,N_563);
xnor U2805 (N_2805,N_442,N_935);
nand U2806 (N_2806,N_1797,N_1867);
nand U2807 (N_2807,N_759,N_1158);
nor U2808 (N_2808,N_1114,N_348);
nand U2809 (N_2809,N_1841,N_85);
nor U2810 (N_2810,N_1567,N_666);
and U2811 (N_2811,N_1662,N_1569);
xnor U2812 (N_2812,N_1923,N_965);
and U2813 (N_2813,N_90,N_99);
xnor U2814 (N_2814,N_986,N_767);
xor U2815 (N_2815,N_878,N_713);
or U2816 (N_2816,N_1444,N_753);
xnor U2817 (N_2817,N_1679,N_798);
or U2818 (N_2818,N_1592,N_287);
nand U2819 (N_2819,N_1090,N_1344);
and U2820 (N_2820,N_296,N_1210);
nand U2821 (N_2821,N_685,N_1884);
and U2822 (N_2822,N_1998,N_1005);
and U2823 (N_2823,N_1084,N_548);
and U2824 (N_2824,N_805,N_403);
xor U2825 (N_2825,N_1938,N_138);
nand U2826 (N_2826,N_1694,N_1838);
xnor U2827 (N_2827,N_564,N_1113);
or U2828 (N_2828,N_475,N_477);
nand U2829 (N_2829,N_1259,N_1673);
or U2830 (N_2830,N_869,N_797);
nand U2831 (N_2831,N_507,N_419);
nand U2832 (N_2832,N_1811,N_1891);
nor U2833 (N_2833,N_1056,N_619);
nand U2834 (N_2834,N_444,N_425);
nor U2835 (N_2835,N_1002,N_1661);
xor U2836 (N_2836,N_1750,N_586);
and U2837 (N_2837,N_1937,N_70);
nand U2838 (N_2838,N_1535,N_940);
xor U2839 (N_2839,N_1711,N_134);
or U2840 (N_2840,N_1420,N_490);
and U2841 (N_2841,N_1438,N_1993);
nor U2842 (N_2842,N_64,N_1353);
nor U2843 (N_2843,N_1023,N_946);
and U2844 (N_2844,N_669,N_524);
nand U2845 (N_2845,N_1512,N_310);
nand U2846 (N_2846,N_678,N_1525);
or U2847 (N_2847,N_267,N_1404);
and U2848 (N_2848,N_1836,N_521);
nor U2849 (N_2849,N_1263,N_1338);
or U2850 (N_2850,N_853,N_764);
or U2851 (N_2851,N_671,N_308);
nor U2852 (N_2852,N_1497,N_1486);
and U2853 (N_2853,N_114,N_1214);
and U2854 (N_2854,N_209,N_1250);
or U2855 (N_2855,N_1478,N_122);
or U2856 (N_2856,N_115,N_670);
nor U2857 (N_2857,N_451,N_1280);
xor U2858 (N_2858,N_426,N_1021);
xnor U2859 (N_2859,N_578,N_385);
or U2860 (N_2860,N_614,N_399);
nor U2861 (N_2861,N_465,N_709);
nand U2862 (N_2862,N_749,N_741);
or U2863 (N_2863,N_826,N_418);
nand U2864 (N_2864,N_1991,N_1892);
or U2865 (N_2865,N_1607,N_1389);
and U2866 (N_2866,N_82,N_219);
and U2867 (N_2867,N_849,N_343);
and U2868 (N_2868,N_711,N_1558);
nor U2869 (N_2869,N_1424,N_328);
and U2870 (N_2870,N_1522,N_251);
or U2871 (N_2871,N_410,N_470);
or U2872 (N_2872,N_121,N_1831);
or U2873 (N_2873,N_1961,N_1258);
xor U2874 (N_2874,N_765,N_1866);
nor U2875 (N_2875,N_331,N_1039);
and U2876 (N_2876,N_535,N_1847);
and U2877 (N_2877,N_754,N_1294);
nand U2878 (N_2878,N_1649,N_777);
nor U2879 (N_2879,N_1356,N_682);
nand U2880 (N_2880,N_657,N_1049);
nor U2881 (N_2881,N_364,N_1287);
nor U2882 (N_2882,N_422,N_359);
xnor U2883 (N_2883,N_738,N_723);
or U2884 (N_2884,N_128,N_117);
and U2885 (N_2885,N_1530,N_1010);
nand U2886 (N_2886,N_1800,N_1703);
or U2887 (N_2887,N_1335,N_824);
and U2888 (N_2888,N_746,N_621);
nor U2889 (N_2889,N_147,N_1970);
nor U2890 (N_2890,N_144,N_602);
or U2891 (N_2891,N_1332,N_823);
nor U2892 (N_2892,N_1820,N_1705);
nor U2893 (N_2893,N_298,N_1768);
nand U2894 (N_2894,N_783,N_730);
nand U2895 (N_2895,N_1397,N_1200);
and U2896 (N_2896,N_1141,N_622);
and U2897 (N_2897,N_1340,N_100);
and U2898 (N_2898,N_1582,N_145);
and U2899 (N_2899,N_72,N_1199);
or U2900 (N_2900,N_1603,N_914);
nand U2901 (N_2901,N_952,N_927);
nand U2902 (N_2902,N_1425,N_17);
nand U2903 (N_2903,N_976,N_234);
and U2904 (N_2904,N_1870,N_78);
or U2905 (N_2905,N_1748,N_1088);
or U2906 (N_2906,N_1304,N_448);
and U2907 (N_2907,N_731,N_199);
or U2908 (N_2908,N_352,N_808);
or U2909 (N_2909,N_130,N_1359);
nor U2910 (N_2910,N_780,N_1518);
nand U2911 (N_2911,N_743,N_1483);
xor U2912 (N_2912,N_1266,N_552);
xnor U2913 (N_2913,N_1730,N_653);
and U2914 (N_2914,N_44,N_873);
xnor U2915 (N_2915,N_486,N_982);
or U2916 (N_2916,N_1930,N_1521);
nor U2917 (N_2917,N_592,N_1995);
nand U2918 (N_2918,N_908,N_1226);
nor U2919 (N_2919,N_525,N_1736);
nor U2920 (N_2920,N_18,N_456);
or U2921 (N_2921,N_321,N_211);
nor U2922 (N_2922,N_1115,N_1219);
or U2923 (N_2923,N_1951,N_24);
or U2924 (N_2924,N_1932,N_789);
nor U2925 (N_2925,N_929,N_1253);
or U2926 (N_2926,N_1509,N_1476);
or U2927 (N_2927,N_496,N_618);
nand U2928 (N_2928,N_717,N_1742);
or U2929 (N_2929,N_790,N_640);
nor U2930 (N_2930,N_1737,N_876);
or U2931 (N_2931,N_1317,N_774);
and U2932 (N_2932,N_1460,N_995);
nand U2933 (N_2933,N_355,N_179);
nand U2934 (N_2934,N_200,N_1565);
or U2935 (N_2935,N_1074,N_1944);
nor U2936 (N_2936,N_480,N_904);
and U2937 (N_2937,N_1452,N_585);
or U2938 (N_2938,N_217,N_1461);
and U2939 (N_2939,N_1808,N_1669);
nor U2940 (N_2940,N_857,N_1156);
or U2941 (N_2941,N_778,N_1533);
nor U2942 (N_2942,N_611,N_832);
and U2943 (N_2943,N_1387,N_1980);
or U2944 (N_2944,N_165,N_1906);
or U2945 (N_2945,N_56,N_782);
and U2946 (N_2946,N_910,N_380);
nand U2947 (N_2947,N_1015,N_63);
nor U2948 (N_2948,N_1935,N_1625);
and U2949 (N_2949,N_631,N_839);
or U2950 (N_2950,N_1721,N_1826);
or U2951 (N_2951,N_781,N_254);
nand U2952 (N_2952,N_290,N_1412);
and U2953 (N_2953,N_647,N_838);
nand U2954 (N_2954,N_1227,N_89);
or U2955 (N_2955,N_919,N_1131);
or U2956 (N_2956,N_1813,N_892);
or U2957 (N_2957,N_1537,N_213);
and U2958 (N_2958,N_1848,N_1713);
and U2959 (N_2959,N_193,N_427);
nor U2960 (N_2960,N_414,N_1342);
or U2961 (N_2961,N_1271,N_1365);
or U2962 (N_2962,N_450,N_1035);
nor U2963 (N_2963,N_1349,N_302);
and U2964 (N_2964,N_1252,N_719);
nand U2965 (N_2965,N_658,N_1104);
nand U2966 (N_2966,N_625,N_665);
or U2967 (N_2967,N_784,N_1888);
or U2968 (N_2968,N_1321,N_351);
and U2969 (N_2969,N_972,N_1383);
nor U2970 (N_2970,N_515,N_1862);
or U2971 (N_2971,N_1629,N_508);
nand U2972 (N_2972,N_408,N_1656);
and U2973 (N_2973,N_1492,N_1610);
and U2974 (N_2974,N_131,N_188);
xnor U2975 (N_2975,N_517,N_966);
or U2976 (N_2976,N_284,N_923);
or U2977 (N_2977,N_1427,N_1785);
xor U2978 (N_2978,N_942,N_1337);
nor U2979 (N_2979,N_959,N_922);
or U2980 (N_2980,N_482,N_1127);
nor U2981 (N_2981,N_1553,N_446);
nand U2982 (N_2982,N_882,N_1782);
nor U2983 (N_2983,N_1799,N_112);
and U2984 (N_2984,N_1041,N_900);
nor U2985 (N_2985,N_1618,N_1154);
nor U2986 (N_2986,N_528,N_1708);
or U2987 (N_2987,N_1016,N_318);
nand U2988 (N_2988,N_1895,N_624);
or U2989 (N_2989,N_1140,N_947);
nor U2990 (N_2990,N_1802,N_1542);
and U2991 (N_2991,N_630,N_761);
nor U2992 (N_2992,N_306,N_1053);
and U2993 (N_2993,N_65,N_398);
or U2994 (N_2994,N_865,N_494);
nor U2995 (N_2995,N_977,N_526);
nor U2996 (N_2996,N_1809,N_94);
and U2997 (N_2997,N_368,N_1034);
nor U2998 (N_2998,N_84,N_407);
nor U2999 (N_2999,N_244,N_278);
nand U3000 (N_3000,N_1968,N_1284);
nand U3001 (N_3001,N_506,N_315);
nor U3002 (N_3002,N_1218,N_1105);
nor U3003 (N_3003,N_513,N_1032);
and U3004 (N_3004,N_521,N_589);
nor U3005 (N_3005,N_591,N_965);
nor U3006 (N_3006,N_327,N_1749);
nand U3007 (N_3007,N_311,N_824);
nor U3008 (N_3008,N_1600,N_1613);
nand U3009 (N_3009,N_1853,N_1541);
and U3010 (N_3010,N_309,N_1196);
nand U3011 (N_3011,N_1682,N_1171);
nor U3012 (N_3012,N_1969,N_795);
and U3013 (N_3013,N_654,N_1096);
nor U3014 (N_3014,N_456,N_295);
and U3015 (N_3015,N_315,N_788);
nor U3016 (N_3016,N_839,N_1184);
nor U3017 (N_3017,N_520,N_770);
and U3018 (N_3018,N_512,N_624);
and U3019 (N_3019,N_1868,N_1432);
nor U3020 (N_3020,N_1294,N_1358);
nor U3021 (N_3021,N_191,N_1901);
nand U3022 (N_3022,N_132,N_1926);
nor U3023 (N_3023,N_873,N_73);
nor U3024 (N_3024,N_1357,N_978);
and U3025 (N_3025,N_1360,N_1132);
nor U3026 (N_3026,N_1998,N_457);
nor U3027 (N_3027,N_80,N_139);
nand U3028 (N_3028,N_1860,N_492);
nand U3029 (N_3029,N_1869,N_1279);
nor U3030 (N_3030,N_490,N_1608);
nand U3031 (N_3031,N_232,N_1582);
nor U3032 (N_3032,N_1461,N_866);
nand U3033 (N_3033,N_208,N_6);
and U3034 (N_3034,N_130,N_1306);
or U3035 (N_3035,N_305,N_128);
or U3036 (N_3036,N_1108,N_279);
and U3037 (N_3037,N_545,N_406);
nand U3038 (N_3038,N_1592,N_1981);
and U3039 (N_3039,N_1462,N_1757);
xnor U3040 (N_3040,N_1228,N_573);
nand U3041 (N_3041,N_182,N_1686);
xnor U3042 (N_3042,N_943,N_1170);
and U3043 (N_3043,N_1550,N_295);
nor U3044 (N_3044,N_1288,N_134);
nor U3045 (N_3045,N_1384,N_1348);
and U3046 (N_3046,N_1541,N_265);
xor U3047 (N_3047,N_1740,N_1782);
or U3048 (N_3048,N_227,N_372);
nand U3049 (N_3049,N_340,N_1703);
nor U3050 (N_3050,N_345,N_1238);
and U3051 (N_3051,N_1800,N_328);
nor U3052 (N_3052,N_1442,N_608);
nor U3053 (N_3053,N_1657,N_1006);
and U3054 (N_3054,N_294,N_1783);
or U3055 (N_3055,N_1633,N_200);
nand U3056 (N_3056,N_215,N_1782);
or U3057 (N_3057,N_573,N_166);
nand U3058 (N_3058,N_354,N_160);
nand U3059 (N_3059,N_759,N_1236);
and U3060 (N_3060,N_477,N_1702);
or U3061 (N_3061,N_1817,N_1265);
nand U3062 (N_3062,N_1241,N_778);
or U3063 (N_3063,N_1744,N_1162);
nor U3064 (N_3064,N_1315,N_1465);
nand U3065 (N_3065,N_1426,N_756);
nor U3066 (N_3066,N_121,N_1199);
and U3067 (N_3067,N_1079,N_1670);
xnor U3068 (N_3068,N_760,N_1054);
nand U3069 (N_3069,N_1311,N_639);
or U3070 (N_3070,N_1237,N_714);
and U3071 (N_3071,N_1000,N_1938);
and U3072 (N_3072,N_746,N_389);
or U3073 (N_3073,N_252,N_85);
and U3074 (N_3074,N_1237,N_76);
nor U3075 (N_3075,N_329,N_379);
and U3076 (N_3076,N_624,N_269);
or U3077 (N_3077,N_346,N_141);
or U3078 (N_3078,N_1558,N_1126);
or U3079 (N_3079,N_920,N_858);
or U3080 (N_3080,N_223,N_1368);
nor U3081 (N_3081,N_1793,N_312);
or U3082 (N_3082,N_117,N_250);
and U3083 (N_3083,N_821,N_520);
nor U3084 (N_3084,N_159,N_855);
and U3085 (N_3085,N_874,N_1704);
and U3086 (N_3086,N_734,N_43);
nand U3087 (N_3087,N_1423,N_746);
and U3088 (N_3088,N_516,N_862);
nor U3089 (N_3089,N_1599,N_1566);
or U3090 (N_3090,N_1663,N_1532);
nand U3091 (N_3091,N_1814,N_16);
and U3092 (N_3092,N_882,N_1880);
nor U3093 (N_3093,N_1129,N_322);
and U3094 (N_3094,N_844,N_3);
and U3095 (N_3095,N_1708,N_1950);
nand U3096 (N_3096,N_1213,N_1689);
nand U3097 (N_3097,N_1236,N_590);
or U3098 (N_3098,N_1029,N_181);
and U3099 (N_3099,N_1090,N_420);
nor U3100 (N_3100,N_123,N_1420);
or U3101 (N_3101,N_298,N_1163);
nor U3102 (N_3102,N_1278,N_376);
or U3103 (N_3103,N_1080,N_1561);
xnor U3104 (N_3104,N_1412,N_128);
nand U3105 (N_3105,N_1152,N_1621);
nor U3106 (N_3106,N_547,N_1009);
and U3107 (N_3107,N_1288,N_1966);
and U3108 (N_3108,N_138,N_883);
nand U3109 (N_3109,N_1009,N_1056);
nor U3110 (N_3110,N_883,N_1389);
nand U3111 (N_3111,N_851,N_343);
xor U3112 (N_3112,N_46,N_1306);
and U3113 (N_3113,N_152,N_1344);
xor U3114 (N_3114,N_493,N_1997);
nor U3115 (N_3115,N_1141,N_782);
nor U3116 (N_3116,N_891,N_1732);
nand U3117 (N_3117,N_276,N_1947);
nor U3118 (N_3118,N_1017,N_1427);
nand U3119 (N_3119,N_1501,N_270);
nor U3120 (N_3120,N_1409,N_670);
xnor U3121 (N_3121,N_1444,N_1970);
nand U3122 (N_3122,N_1628,N_1404);
nor U3123 (N_3123,N_860,N_856);
nor U3124 (N_3124,N_1141,N_1761);
and U3125 (N_3125,N_1738,N_1198);
or U3126 (N_3126,N_1305,N_821);
or U3127 (N_3127,N_1508,N_464);
and U3128 (N_3128,N_302,N_402);
xor U3129 (N_3129,N_533,N_1691);
and U3130 (N_3130,N_851,N_833);
or U3131 (N_3131,N_1317,N_1612);
nor U3132 (N_3132,N_1185,N_448);
nand U3133 (N_3133,N_1077,N_1989);
nor U3134 (N_3134,N_419,N_865);
and U3135 (N_3135,N_1268,N_1738);
nand U3136 (N_3136,N_1839,N_1262);
and U3137 (N_3137,N_1671,N_1331);
and U3138 (N_3138,N_779,N_387);
nand U3139 (N_3139,N_1150,N_1291);
or U3140 (N_3140,N_289,N_1059);
and U3141 (N_3141,N_538,N_243);
nand U3142 (N_3142,N_795,N_876);
xor U3143 (N_3143,N_983,N_609);
and U3144 (N_3144,N_1353,N_741);
and U3145 (N_3145,N_519,N_965);
nand U3146 (N_3146,N_693,N_1453);
or U3147 (N_3147,N_1546,N_1789);
nand U3148 (N_3148,N_893,N_1781);
xor U3149 (N_3149,N_1693,N_1759);
xor U3150 (N_3150,N_1403,N_1912);
and U3151 (N_3151,N_277,N_1488);
and U3152 (N_3152,N_1244,N_1755);
or U3153 (N_3153,N_888,N_127);
and U3154 (N_3154,N_245,N_1150);
nand U3155 (N_3155,N_1039,N_432);
or U3156 (N_3156,N_1993,N_269);
or U3157 (N_3157,N_1916,N_733);
and U3158 (N_3158,N_842,N_505);
nor U3159 (N_3159,N_1804,N_428);
nor U3160 (N_3160,N_411,N_1141);
or U3161 (N_3161,N_550,N_242);
or U3162 (N_3162,N_597,N_1173);
nand U3163 (N_3163,N_365,N_590);
or U3164 (N_3164,N_228,N_1941);
nand U3165 (N_3165,N_1178,N_1619);
or U3166 (N_3166,N_1978,N_1937);
xnor U3167 (N_3167,N_778,N_940);
and U3168 (N_3168,N_300,N_480);
or U3169 (N_3169,N_1037,N_1589);
and U3170 (N_3170,N_463,N_1135);
and U3171 (N_3171,N_1991,N_1578);
or U3172 (N_3172,N_1450,N_1385);
and U3173 (N_3173,N_1460,N_1223);
nor U3174 (N_3174,N_1911,N_1207);
and U3175 (N_3175,N_1085,N_577);
nor U3176 (N_3176,N_386,N_825);
nor U3177 (N_3177,N_878,N_242);
nor U3178 (N_3178,N_799,N_194);
and U3179 (N_3179,N_1687,N_1219);
nor U3180 (N_3180,N_1217,N_781);
nand U3181 (N_3181,N_1015,N_509);
nand U3182 (N_3182,N_1002,N_1832);
nor U3183 (N_3183,N_395,N_1824);
xor U3184 (N_3184,N_1368,N_1167);
and U3185 (N_3185,N_1346,N_1309);
nand U3186 (N_3186,N_739,N_867);
and U3187 (N_3187,N_1766,N_1605);
nand U3188 (N_3188,N_1507,N_1652);
nor U3189 (N_3189,N_1318,N_1665);
nand U3190 (N_3190,N_154,N_806);
nor U3191 (N_3191,N_1183,N_233);
nand U3192 (N_3192,N_1692,N_1077);
nor U3193 (N_3193,N_848,N_497);
nor U3194 (N_3194,N_1153,N_577);
and U3195 (N_3195,N_1096,N_495);
or U3196 (N_3196,N_1870,N_762);
and U3197 (N_3197,N_146,N_1997);
nor U3198 (N_3198,N_844,N_89);
or U3199 (N_3199,N_1429,N_1207);
and U3200 (N_3200,N_577,N_1747);
or U3201 (N_3201,N_463,N_1439);
nand U3202 (N_3202,N_1810,N_369);
and U3203 (N_3203,N_1033,N_1743);
or U3204 (N_3204,N_1435,N_1998);
nand U3205 (N_3205,N_216,N_1914);
nand U3206 (N_3206,N_1471,N_421);
and U3207 (N_3207,N_1634,N_1330);
or U3208 (N_3208,N_1874,N_941);
nand U3209 (N_3209,N_472,N_1197);
and U3210 (N_3210,N_1544,N_1594);
nor U3211 (N_3211,N_1193,N_1569);
or U3212 (N_3212,N_471,N_584);
and U3213 (N_3213,N_779,N_1258);
nand U3214 (N_3214,N_138,N_856);
or U3215 (N_3215,N_1016,N_158);
and U3216 (N_3216,N_987,N_586);
nor U3217 (N_3217,N_352,N_1524);
or U3218 (N_3218,N_1394,N_1334);
and U3219 (N_3219,N_1977,N_1118);
nand U3220 (N_3220,N_43,N_949);
xnor U3221 (N_3221,N_934,N_722);
and U3222 (N_3222,N_1926,N_677);
nand U3223 (N_3223,N_607,N_1559);
nand U3224 (N_3224,N_1485,N_431);
nor U3225 (N_3225,N_54,N_1027);
and U3226 (N_3226,N_695,N_594);
nor U3227 (N_3227,N_250,N_1160);
nor U3228 (N_3228,N_380,N_905);
or U3229 (N_3229,N_1677,N_1641);
and U3230 (N_3230,N_0,N_1446);
or U3231 (N_3231,N_1107,N_853);
xnor U3232 (N_3232,N_1460,N_450);
nor U3233 (N_3233,N_379,N_1965);
nand U3234 (N_3234,N_1040,N_1255);
or U3235 (N_3235,N_499,N_531);
nor U3236 (N_3236,N_931,N_1504);
or U3237 (N_3237,N_606,N_551);
xor U3238 (N_3238,N_1060,N_1180);
or U3239 (N_3239,N_1270,N_114);
nand U3240 (N_3240,N_1261,N_566);
or U3241 (N_3241,N_898,N_1529);
nand U3242 (N_3242,N_1811,N_215);
nor U3243 (N_3243,N_79,N_865);
or U3244 (N_3244,N_1460,N_1321);
or U3245 (N_3245,N_231,N_1218);
xor U3246 (N_3246,N_1049,N_1912);
nand U3247 (N_3247,N_483,N_1386);
or U3248 (N_3248,N_1903,N_1351);
nand U3249 (N_3249,N_1954,N_898);
and U3250 (N_3250,N_261,N_1747);
nand U3251 (N_3251,N_1002,N_1160);
and U3252 (N_3252,N_883,N_741);
nor U3253 (N_3253,N_1490,N_290);
xor U3254 (N_3254,N_1442,N_1900);
or U3255 (N_3255,N_46,N_1570);
nand U3256 (N_3256,N_820,N_1703);
and U3257 (N_3257,N_1142,N_590);
nand U3258 (N_3258,N_451,N_1596);
nand U3259 (N_3259,N_362,N_474);
and U3260 (N_3260,N_706,N_492);
or U3261 (N_3261,N_1867,N_1725);
nor U3262 (N_3262,N_1456,N_1003);
nand U3263 (N_3263,N_1761,N_1314);
and U3264 (N_3264,N_1747,N_205);
nand U3265 (N_3265,N_152,N_1328);
and U3266 (N_3266,N_1099,N_889);
or U3267 (N_3267,N_989,N_636);
or U3268 (N_3268,N_823,N_347);
nor U3269 (N_3269,N_119,N_1664);
and U3270 (N_3270,N_469,N_305);
nor U3271 (N_3271,N_619,N_27);
nor U3272 (N_3272,N_1063,N_497);
nor U3273 (N_3273,N_1450,N_448);
and U3274 (N_3274,N_1002,N_616);
or U3275 (N_3275,N_1316,N_819);
or U3276 (N_3276,N_403,N_369);
or U3277 (N_3277,N_1292,N_1679);
nand U3278 (N_3278,N_128,N_628);
nand U3279 (N_3279,N_1241,N_1250);
and U3280 (N_3280,N_791,N_856);
nor U3281 (N_3281,N_414,N_572);
xor U3282 (N_3282,N_1117,N_501);
nor U3283 (N_3283,N_1408,N_99);
and U3284 (N_3284,N_1142,N_1479);
nand U3285 (N_3285,N_1534,N_1740);
nand U3286 (N_3286,N_889,N_949);
nor U3287 (N_3287,N_119,N_464);
or U3288 (N_3288,N_37,N_1152);
or U3289 (N_3289,N_104,N_82);
and U3290 (N_3290,N_1835,N_1170);
nand U3291 (N_3291,N_62,N_1846);
nor U3292 (N_3292,N_56,N_214);
nor U3293 (N_3293,N_1180,N_1017);
and U3294 (N_3294,N_1467,N_896);
nand U3295 (N_3295,N_1503,N_1161);
nand U3296 (N_3296,N_1159,N_1641);
nand U3297 (N_3297,N_1225,N_1953);
and U3298 (N_3298,N_1678,N_242);
nand U3299 (N_3299,N_222,N_788);
nor U3300 (N_3300,N_1699,N_523);
and U3301 (N_3301,N_1421,N_1730);
or U3302 (N_3302,N_698,N_62);
nor U3303 (N_3303,N_618,N_471);
and U3304 (N_3304,N_716,N_998);
or U3305 (N_3305,N_925,N_1552);
nor U3306 (N_3306,N_605,N_1998);
and U3307 (N_3307,N_461,N_635);
xor U3308 (N_3308,N_4,N_726);
and U3309 (N_3309,N_773,N_708);
xnor U3310 (N_3310,N_315,N_276);
nor U3311 (N_3311,N_731,N_1399);
nand U3312 (N_3312,N_208,N_750);
and U3313 (N_3313,N_787,N_1109);
or U3314 (N_3314,N_482,N_959);
or U3315 (N_3315,N_1039,N_688);
or U3316 (N_3316,N_818,N_624);
and U3317 (N_3317,N_255,N_1085);
and U3318 (N_3318,N_1318,N_179);
nand U3319 (N_3319,N_1335,N_87);
xor U3320 (N_3320,N_1077,N_545);
or U3321 (N_3321,N_263,N_1469);
nor U3322 (N_3322,N_407,N_1751);
nor U3323 (N_3323,N_130,N_1953);
or U3324 (N_3324,N_705,N_1726);
or U3325 (N_3325,N_1803,N_717);
nor U3326 (N_3326,N_1807,N_162);
and U3327 (N_3327,N_312,N_569);
or U3328 (N_3328,N_701,N_1445);
nor U3329 (N_3329,N_1145,N_818);
nand U3330 (N_3330,N_635,N_941);
nand U3331 (N_3331,N_1672,N_1184);
nand U3332 (N_3332,N_446,N_1425);
or U3333 (N_3333,N_133,N_711);
nand U3334 (N_3334,N_1959,N_1050);
and U3335 (N_3335,N_1953,N_724);
nand U3336 (N_3336,N_449,N_579);
nor U3337 (N_3337,N_1400,N_1941);
nor U3338 (N_3338,N_1917,N_541);
nor U3339 (N_3339,N_1541,N_1804);
or U3340 (N_3340,N_1371,N_660);
or U3341 (N_3341,N_1783,N_1944);
nor U3342 (N_3342,N_507,N_886);
xor U3343 (N_3343,N_945,N_1034);
xnor U3344 (N_3344,N_226,N_74);
xnor U3345 (N_3345,N_353,N_899);
nor U3346 (N_3346,N_799,N_201);
nor U3347 (N_3347,N_1073,N_1014);
nor U3348 (N_3348,N_222,N_1827);
and U3349 (N_3349,N_717,N_544);
xnor U3350 (N_3350,N_477,N_1254);
nand U3351 (N_3351,N_546,N_1006);
nor U3352 (N_3352,N_881,N_384);
and U3353 (N_3353,N_1830,N_1173);
nor U3354 (N_3354,N_581,N_1057);
nor U3355 (N_3355,N_854,N_406);
nor U3356 (N_3356,N_1622,N_1498);
nand U3357 (N_3357,N_51,N_98);
and U3358 (N_3358,N_1056,N_1114);
xor U3359 (N_3359,N_1903,N_457);
nor U3360 (N_3360,N_1044,N_1963);
or U3361 (N_3361,N_381,N_81);
nand U3362 (N_3362,N_355,N_575);
nand U3363 (N_3363,N_165,N_1493);
and U3364 (N_3364,N_668,N_242);
and U3365 (N_3365,N_220,N_466);
nor U3366 (N_3366,N_1677,N_1515);
nand U3367 (N_3367,N_1201,N_628);
or U3368 (N_3368,N_1703,N_1465);
nand U3369 (N_3369,N_1619,N_393);
nor U3370 (N_3370,N_213,N_502);
or U3371 (N_3371,N_937,N_218);
and U3372 (N_3372,N_705,N_1642);
nand U3373 (N_3373,N_1206,N_262);
or U3374 (N_3374,N_354,N_1609);
or U3375 (N_3375,N_1176,N_584);
and U3376 (N_3376,N_1736,N_1218);
nand U3377 (N_3377,N_1588,N_43);
nand U3378 (N_3378,N_1977,N_532);
nor U3379 (N_3379,N_1022,N_1074);
nand U3380 (N_3380,N_584,N_1161);
or U3381 (N_3381,N_241,N_198);
nand U3382 (N_3382,N_471,N_1730);
and U3383 (N_3383,N_1188,N_1056);
xnor U3384 (N_3384,N_1947,N_1702);
nand U3385 (N_3385,N_1866,N_277);
xnor U3386 (N_3386,N_743,N_594);
nor U3387 (N_3387,N_653,N_110);
and U3388 (N_3388,N_561,N_666);
nand U3389 (N_3389,N_1599,N_221);
nor U3390 (N_3390,N_1045,N_1087);
and U3391 (N_3391,N_1210,N_23);
or U3392 (N_3392,N_1998,N_438);
and U3393 (N_3393,N_465,N_1985);
and U3394 (N_3394,N_301,N_1922);
or U3395 (N_3395,N_58,N_1457);
or U3396 (N_3396,N_972,N_1377);
and U3397 (N_3397,N_261,N_181);
and U3398 (N_3398,N_1679,N_274);
or U3399 (N_3399,N_1141,N_1496);
nor U3400 (N_3400,N_669,N_1988);
nor U3401 (N_3401,N_523,N_1849);
nor U3402 (N_3402,N_1671,N_1456);
or U3403 (N_3403,N_1861,N_971);
and U3404 (N_3404,N_231,N_57);
or U3405 (N_3405,N_1547,N_467);
nand U3406 (N_3406,N_157,N_380);
and U3407 (N_3407,N_1024,N_831);
nor U3408 (N_3408,N_1397,N_1000);
xor U3409 (N_3409,N_1985,N_1120);
nor U3410 (N_3410,N_19,N_652);
and U3411 (N_3411,N_203,N_456);
and U3412 (N_3412,N_1684,N_1877);
nand U3413 (N_3413,N_1376,N_1938);
nand U3414 (N_3414,N_1776,N_959);
or U3415 (N_3415,N_1806,N_780);
or U3416 (N_3416,N_779,N_756);
nand U3417 (N_3417,N_697,N_1079);
nor U3418 (N_3418,N_597,N_1621);
or U3419 (N_3419,N_1777,N_135);
or U3420 (N_3420,N_1405,N_404);
and U3421 (N_3421,N_1191,N_1143);
and U3422 (N_3422,N_1166,N_1696);
nand U3423 (N_3423,N_1100,N_1815);
nor U3424 (N_3424,N_1580,N_287);
and U3425 (N_3425,N_1578,N_173);
nand U3426 (N_3426,N_1433,N_302);
nor U3427 (N_3427,N_1750,N_1542);
nor U3428 (N_3428,N_1592,N_1734);
or U3429 (N_3429,N_653,N_455);
and U3430 (N_3430,N_885,N_1394);
and U3431 (N_3431,N_432,N_1585);
nor U3432 (N_3432,N_509,N_1756);
nor U3433 (N_3433,N_1624,N_824);
xor U3434 (N_3434,N_610,N_1240);
and U3435 (N_3435,N_415,N_219);
nor U3436 (N_3436,N_1047,N_1210);
or U3437 (N_3437,N_489,N_571);
or U3438 (N_3438,N_1005,N_829);
nand U3439 (N_3439,N_668,N_214);
or U3440 (N_3440,N_400,N_1130);
and U3441 (N_3441,N_121,N_1797);
or U3442 (N_3442,N_490,N_836);
and U3443 (N_3443,N_1245,N_1789);
and U3444 (N_3444,N_726,N_1848);
or U3445 (N_3445,N_253,N_413);
or U3446 (N_3446,N_1766,N_331);
xor U3447 (N_3447,N_1330,N_1893);
and U3448 (N_3448,N_209,N_1041);
and U3449 (N_3449,N_22,N_1264);
nor U3450 (N_3450,N_1506,N_1706);
or U3451 (N_3451,N_1615,N_132);
nand U3452 (N_3452,N_797,N_1162);
and U3453 (N_3453,N_1807,N_1655);
nand U3454 (N_3454,N_1737,N_1906);
nand U3455 (N_3455,N_1893,N_240);
nor U3456 (N_3456,N_1193,N_1996);
nand U3457 (N_3457,N_224,N_292);
nand U3458 (N_3458,N_631,N_249);
nor U3459 (N_3459,N_1655,N_1146);
nand U3460 (N_3460,N_1056,N_1029);
nand U3461 (N_3461,N_813,N_477);
nand U3462 (N_3462,N_228,N_268);
nand U3463 (N_3463,N_137,N_409);
and U3464 (N_3464,N_1160,N_927);
and U3465 (N_3465,N_584,N_693);
nor U3466 (N_3466,N_929,N_866);
xor U3467 (N_3467,N_214,N_1457);
nand U3468 (N_3468,N_1086,N_613);
and U3469 (N_3469,N_1628,N_645);
nand U3470 (N_3470,N_1474,N_1235);
nor U3471 (N_3471,N_635,N_1946);
or U3472 (N_3472,N_1122,N_1971);
xor U3473 (N_3473,N_1979,N_1486);
or U3474 (N_3474,N_1205,N_539);
nand U3475 (N_3475,N_1854,N_798);
nand U3476 (N_3476,N_1532,N_1927);
xnor U3477 (N_3477,N_1393,N_1024);
nand U3478 (N_3478,N_1334,N_1327);
and U3479 (N_3479,N_851,N_1109);
or U3480 (N_3480,N_621,N_944);
and U3481 (N_3481,N_1646,N_982);
nor U3482 (N_3482,N_602,N_949);
nor U3483 (N_3483,N_679,N_1600);
xor U3484 (N_3484,N_1205,N_15);
nor U3485 (N_3485,N_1597,N_689);
xor U3486 (N_3486,N_878,N_700);
nor U3487 (N_3487,N_1156,N_1494);
or U3488 (N_3488,N_87,N_816);
nor U3489 (N_3489,N_1047,N_1795);
nand U3490 (N_3490,N_1638,N_1920);
and U3491 (N_3491,N_283,N_976);
nor U3492 (N_3492,N_1550,N_687);
nor U3493 (N_3493,N_1144,N_64);
nand U3494 (N_3494,N_726,N_1683);
nand U3495 (N_3495,N_282,N_1260);
or U3496 (N_3496,N_1740,N_386);
or U3497 (N_3497,N_979,N_1308);
nand U3498 (N_3498,N_392,N_1273);
or U3499 (N_3499,N_1389,N_1771);
and U3500 (N_3500,N_755,N_385);
nor U3501 (N_3501,N_572,N_1082);
or U3502 (N_3502,N_761,N_1065);
nor U3503 (N_3503,N_875,N_1414);
and U3504 (N_3504,N_1839,N_1792);
nand U3505 (N_3505,N_89,N_1304);
xor U3506 (N_3506,N_251,N_1220);
and U3507 (N_3507,N_443,N_804);
nor U3508 (N_3508,N_1563,N_1875);
and U3509 (N_3509,N_1531,N_1171);
nor U3510 (N_3510,N_728,N_1292);
nand U3511 (N_3511,N_1499,N_1262);
or U3512 (N_3512,N_1956,N_1937);
or U3513 (N_3513,N_1283,N_1747);
or U3514 (N_3514,N_1524,N_766);
nor U3515 (N_3515,N_1893,N_1793);
and U3516 (N_3516,N_545,N_323);
nor U3517 (N_3517,N_288,N_630);
or U3518 (N_3518,N_1164,N_859);
xor U3519 (N_3519,N_1262,N_1030);
or U3520 (N_3520,N_1473,N_1101);
nor U3521 (N_3521,N_1261,N_1014);
or U3522 (N_3522,N_1034,N_101);
and U3523 (N_3523,N_4,N_1947);
or U3524 (N_3524,N_810,N_1337);
nor U3525 (N_3525,N_386,N_254);
nand U3526 (N_3526,N_1534,N_530);
or U3527 (N_3527,N_1125,N_635);
xor U3528 (N_3528,N_302,N_478);
and U3529 (N_3529,N_1739,N_725);
nand U3530 (N_3530,N_1120,N_912);
nor U3531 (N_3531,N_598,N_472);
and U3532 (N_3532,N_463,N_1869);
and U3533 (N_3533,N_80,N_316);
nand U3534 (N_3534,N_557,N_1237);
and U3535 (N_3535,N_1239,N_1015);
or U3536 (N_3536,N_739,N_59);
and U3537 (N_3537,N_693,N_1444);
and U3538 (N_3538,N_173,N_972);
nor U3539 (N_3539,N_1781,N_53);
xnor U3540 (N_3540,N_143,N_1667);
and U3541 (N_3541,N_1655,N_940);
or U3542 (N_3542,N_1656,N_275);
nand U3543 (N_3543,N_893,N_1006);
and U3544 (N_3544,N_1540,N_900);
or U3545 (N_3545,N_552,N_441);
nor U3546 (N_3546,N_51,N_1712);
nand U3547 (N_3547,N_856,N_548);
or U3548 (N_3548,N_1565,N_1582);
or U3549 (N_3549,N_972,N_1730);
nand U3550 (N_3550,N_1020,N_287);
and U3551 (N_3551,N_136,N_1793);
xnor U3552 (N_3552,N_1549,N_1260);
or U3553 (N_3553,N_703,N_1769);
nor U3554 (N_3554,N_921,N_1834);
or U3555 (N_3555,N_1724,N_681);
nand U3556 (N_3556,N_370,N_576);
xnor U3557 (N_3557,N_62,N_196);
nand U3558 (N_3558,N_1954,N_915);
nor U3559 (N_3559,N_399,N_1755);
nand U3560 (N_3560,N_1127,N_86);
and U3561 (N_3561,N_842,N_1386);
nor U3562 (N_3562,N_1201,N_1099);
xnor U3563 (N_3563,N_1449,N_746);
and U3564 (N_3564,N_803,N_890);
nand U3565 (N_3565,N_1398,N_1538);
nor U3566 (N_3566,N_146,N_1236);
nand U3567 (N_3567,N_768,N_1466);
xor U3568 (N_3568,N_889,N_703);
and U3569 (N_3569,N_1412,N_1584);
or U3570 (N_3570,N_1908,N_1443);
or U3571 (N_3571,N_1791,N_649);
and U3572 (N_3572,N_819,N_479);
nor U3573 (N_3573,N_100,N_1376);
nand U3574 (N_3574,N_1159,N_1217);
and U3575 (N_3575,N_262,N_546);
and U3576 (N_3576,N_168,N_199);
nor U3577 (N_3577,N_1485,N_979);
nand U3578 (N_3578,N_1051,N_1763);
nor U3579 (N_3579,N_1072,N_1377);
nor U3580 (N_3580,N_911,N_1143);
nor U3581 (N_3581,N_229,N_1609);
nor U3582 (N_3582,N_1411,N_673);
or U3583 (N_3583,N_581,N_1611);
xor U3584 (N_3584,N_1971,N_1758);
xnor U3585 (N_3585,N_1587,N_611);
nor U3586 (N_3586,N_1061,N_1222);
nand U3587 (N_3587,N_1221,N_579);
or U3588 (N_3588,N_1373,N_1823);
nor U3589 (N_3589,N_1801,N_105);
nand U3590 (N_3590,N_937,N_329);
or U3591 (N_3591,N_1904,N_604);
nand U3592 (N_3592,N_157,N_1041);
or U3593 (N_3593,N_1861,N_1859);
or U3594 (N_3594,N_237,N_99);
nor U3595 (N_3595,N_563,N_1961);
xor U3596 (N_3596,N_347,N_1851);
nor U3597 (N_3597,N_1667,N_533);
nor U3598 (N_3598,N_37,N_1300);
xor U3599 (N_3599,N_1141,N_1088);
or U3600 (N_3600,N_112,N_283);
nor U3601 (N_3601,N_705,N_1234);
xnor U3602 (N_3602,N_1061,N_1055);
or U3603 (N_3603,N_599,N_355);
nor U3604 (N_3604,N_1459,N_588);
nor U3605 (N_3605,N_1128,N_97);
nor U3606 (N_3606,N_609,N_421);
and U3607 (N_3607,N_1002,N_162);
or U3608 (N_3608,N_1443,N_1153);
and U3609 (N_3609,N_1910,N_1267);
or U3610 (N_3610,N_1872,N_1914);
nor U3611 (N_3611,N_1296,N_254);
nor U3612 (N_3612,N_1526,N_355);
nand U3613 (N_3613,N_1716,N_125);
nand U3614 (N_3614,N_338,N_684);
or U3615 (N_3615,N_1765,N_419);
nand U3616 (N_3616,N_1377,N_936);
nand U3617 (N_3617,N_799,N_636);
nand U3618 (N_3618,N_1842,N_573);
nand U3619 (N_3619,N_828,N_1485);
nor U3620 (N_3620,N_1896,N_604);
and U3621 (N_3621,N_1966,N_471);
nand U3622 (N_3622,N_1709,N_762);
nor U3623 (N_3623,N_437,N_1763);
or U3624 (N_3624,N_375,N_1829);
nor U3625 (N_3625,N_748,N_938);
and U3626 (N_3626,N_141,N_1701);
nand U3627 (N_3627,N_1290,N_178);
or U3628 (N_3628,N_122,N_1731);
and U3629 (N_3629,N_510,N_399);
or U3630 (N_3630,N_1551,N_786);
or U3631 (N_3631,N_1540,N_1318);
nor U3632 (N_3632,N_1823,N_156);
or U3633 (N_3633,N_1732,N_27);
nand U3634 (N_3634,N_143,N_1304);
or U3635 (N_3635,N_540,N_1553);
or U3636 (N_3636,N_767,N_658);
or U3637 (N_3637,N_1018,N_1499);
xnor U3638 (N_3638,N_1479,N_31);
and U3639 (N_3639,N_678,N_1308);
nor U3640 (N_3640,N_243,N_751);
nand U3641 (N_3641,N_1645,N_341);
or U3642 (N_3642,N_1978,N_58);
xor U3643 (N_3643,N_1550,N_1694);
nand U3644 (N_3644,N_965,N_1382);
nor U3645 (N_3645,N_664,N_944);
nand U3646 (N_3646,N_772,N_898);
nor U3647 (N_3647,N_1542,N_1642);
or U3648 (N_3648,N_1806,N_276);
nand U3649 (N_3649,N_1260,N_225);
and U3650 (N_3650,N_1972,N_354);
nor U3651 (N_3651,N_1483,N_1465);
nand U3652 (N_3652,N_1244,N_289);
nand U3653 (N_3653,N_925,N_1073);
or U3654 (N_3654,N_1785,N_644);
and U3655 (N_3655,N_1482,N_1838);
nand U3656 (N_3656,N_972,N_1382);
nand U3657 (N_3657,N_50,N_815);
nor U3658 (N_3658,N_1164,N_1808);
nand U3659 (N_3659,N_718,N_181);
xnor U3660 (N_3660,N_1003,N_976);
and U3661 (N_3661,N_1353,N_769);
and U3662 (N_3662,N_1217,N_602);
nand U3663 (N_3663,N_814,N_285);
nor U3664 (N_3664,N_115,N_399);
nor U3665 (N_3665,N_504,N_76);
or U3666 (N_3666,N_1641,N_1863);
xnor U3667 (N_3667,N_1290,N_77);
xor U3668 (N_3668,N_1258,N_244);
nand U3669 (N_3669,N_1926,N_1039);
nor U3670 (N_3670,N_1313,N_1762);
and U3671 (N_3671,N_829,N_739);
nand U3672 (N_3672,N_925,N_981);
and U3673 (N_3673,N_809,N_292);
nand U3674 (N_3674,N_1922,N_1584);
nand U3675 (N_3675,N_1353,N_1818);
nand U3676 (N_3676,N_1070,N_1818);
xor U3677 (N_3677,N_1031,N_322);
or U3678 (N_3678,N_664,N_1887);
nand U3679 (N_3679,N_1621,N_622);
and U3680 (N_3680,N_963,N_1646);
xnor U3681 (N_3681,N_810,N_1918);
or U3682 (N_3682,N_1305,N_1942);
and U3683 (N_3683,N_756,N_1736);
nand U3684 (N_3684,N_230,N_983);
and U3685 (N_3685,N_861,N_1741);
or U3686 (N_3686,N_1320,N_424);
or U3687 (N_3687,N_626,N_1366);
and U3688 (N_3688,N_322,N_1487);
and U3689 (N_3689,N_1313,N_1618);
or U3690 (N_3690,N_1442,N_1416);
and U3691 (N_3691,N_1820,N_1950);
nor U3692 (N_3692,N_814,N_976);
nand U3693 (N_3693,N_838,N_888);
and U3694 (N_3694,N_169,N_1105);
xor U3695 (N_3695,N_1951,N_1181);
nor U3696 (N_3696,N_917,N_1246);
or U3697 (N_3697,N_719,N_1685);
or U3698 (N_3698,N_733,N_73);
nand U3699 (N_3699,N_1107,N_1349);
xor U3700 (N_3700,N_65,N_1256);
nand U3701 (N_3701,N_1765,N_378);
nand U3702 (N_3702,N_412,N_1790);
nor U3703 (N_3703,N_1967,N_1501);
or U3704 (N_3704,N_1386,N_1181);
nand U3705 (N_3705,N_1484,N_1251);
xnor U3706 (N_3706,N_1439,N_831);
and U3707 (N_3707,N_1745,N_1243);
or U3708 (N_3708,N_1876,N_1472);
nand U3709 (N_3709,N_1542,N_1611);
nand U3710 (N_3710,N_542,N_1049);
and U3711 (N_3711,N_199,N_117);
xor U3712 (N_3712,N_429,N_637);
and U3713 (N_3713,N_1542,N_858);
and U3714 (N_3714,N_188,N_696);
nor U3715 (N_3715,N_110,N_8);
xor U3716 (N_3716,N_1724,N_1923);
nor U3717 (N_3717,N_788,N_1393);
nand U3718 (N_3718,N_1999,N_1702);
or U3719 (N_3719,N_1218,N_1916);
nor U3720 (N_3720,N_1079,N_647);
or U3721 (N_3721,N_438,N_1274);
or U3722 (N_3722,N_1956,N_841);
nand U3723 (N_3723,N_937,N_1178);
nor U3724 (N_3724,N_233,N_1515);
nand U3725 (N_3725,N_1149,N_595);
or U3726 (N_3726,N_1409,N_1681);
nand U3727 (N_3727,N_1966,N_247);
and U3728 (N_3728,N_786,N_799);
or U3729 (N_3729,N_632,N_616);
or U3730 (N_3730,N_701,N_1615);
and U3731 (N_3731,N_376,N_1619);
nor U3732 (N_3732,N_1751,N_485);
or U3733 (N_3733,N_880,N_1750);
xor U3734 (N_3734,N_1911,N_579);
and U3735 (N_3735,N_1283,N_318);
or U3736 (N_3736,N_1591,N_1266);
or U3737 (N_3737,N_1498,N_454);
nor U3738 (N_3738,N_489,N_1173);
nor U3739 (N_3739,N_1954,N_1875);
and U3740 (N_3740,N_1020,N_1006);
xor U3741 (N_3741,N_1610,N_1785);
and U3742 (N_3742,N_31,N_41);
nor U3743 (N_3743,N_929,N_1382);
nand U3744 (N_3744,N_1587,N_1547);
nand U3745 (N_3745,N_687,N_1406);
and U3746 (N_3746,N_978,N_950);
or U3747 (N_3747,N_1068,N_1245);
nor U3748 (N_3748,N_1998,N_363);
xnor U3749 (N_3749,N_1865,N_1599);
nand U3750 (N_3750,N_1806,N_1731);
nor U3751 (N_3751,N_1166,N_668);
xnor U3752 (N_3752,N_1287,N_726);
or U3753 (N_3753,N_1703,N_1883);
nand U3754 (N_3754,N_1486,N_447);
or U3755 (N_3755,N_1704,N_1296);
nand U3756 (N_3756,N_1416,N_1216);
or U3757 (N_3757,N_99,N_683);
or U3758 (N_3758,N_632,N_877);
nor U3759 (N_3759,N_635,N_1118);
and U3760 (N_3760,N_1580,N_1592);
and U3761 (N_3761,N_1691,N_822);
and U3762 (N_3762,N_480,N_365);
and U3763 (N_3763,N_290,N_520);
nand U3764 (N_3764,N_1497,N_1298);
nand U3765 (N_3765,N_1169,N_356);
nor U3766 (N_3766,N_1266,N_754);
nand U3767 (N_3767,N_949,N_872);
nand U3768 (N_3768,N_32,N_362);
nor U3769 (N_3769,N_234,N_766);
nor U3770 (N_3770,N_1834,N_1182);
xnor U3771 (N_3771,N_1175,N_892);
xnor U3772 (N_3772,N_733,N_273);
and U3773 (N_3773,N_824,N_426);
or U3774 (N_3774,N_204,N_1054);
or U3775 (N_3775,N_502,N_1589);
or U3776 (N_3776,N_214,N_1675);
nor U3777 (N_3777,N_1321,N_1843);
nor U3778 (N_3778,N_1885,N_158);
or U3779 (N_3779,N_329,N_1201);
nand U3780 (N_3780,N_1333,N_1441);
and U3781 (N_3781,N_10,N_926);
xnor U3782 (N_3782,N_15,N_958);
and U3783 (N_3783,N_1653,N_1871);
nand U3784 (N_3784,N_1750,N_1907);
nand U3785 (N_3785,N_1092,N_927);
nor U3786 (N_3786,N_207,N_56);
and U3787 (N_3787,N_1538,N_1505);
and U3788 (N_3788,N_1703,N_999);
nor U3789 (N_3789,N_293,N_1528);
and U3790 (N_3790,N_158,N_352);
nand U3791 (N_3791,N_943,N_736);
xnor U3792 (N_3792,N_1443,N_1735);
and U3793 (N_3793,N_1670,N_1057);
and U3794 (N_3794,N_882,N_1285);
or U3795 (N_3795,N_1102,N_1015);
or U3796 (N_3796,N_590,N_79);
and U3797 (N_3797,N_368,N_427);
and U3798 (N_3798,N_39,N_122);
nand U3799 (N_3799,N_524,N_661);
and U3800 (N_3800,N_1382,N_941);
nand U3801 (N_3801,N_854,N_725);
nor U3802 (N_3802,N_701,N_1800);
nand U3803 (N_3803,N_1404,N_1802);
xor U3804 (N_3804,N_721,N_807);
or U3805 (N_3805,N_1989,N_1351);
nand U3806 (N_3806,N_1136,N_771);
or U3807 (N_3807,N_1083,N_1741);
nor U3808 (N_3808,N_1098,N_1834);
nor U3809 (N_3809,N_1387,N_483);
or U3810 (N_3810,N_333,N_1185);
nor U3811 (N_3811,N_1971,N_1059);
nand U3812 (N_3812,N_1203,N_286);
xor U3813 (N_3813,N_439,N_159);
and U3814 (N_3814,N_1574,N_117);
xnor U3815 (N_3815,N_1608,N_1183);
or U3816 (N_3816,N_927,N_1686);
nand U3817 (N_3817,N_247,N_1024);
nor U3818 (N_3818,N_1844,N_145);
and U3819 (N_3819,N_1939,N_609);
nor U3820 (N_3820,N_1338,N_340);
or U3821 (N_3821,N_1159,N_1450);
and U3822 (N_3822,N_1329,N_1716);
nor U3823 (N_3823,N_536,N_1341);
nor U3824 (N_3824,N_1464,N_1208);
nand U3825 (N_3825,N_999,N_1442);
and U3826 (N_3826,N_1284,N_362);
nor U3827 (N_3827,N_529,N_563);
and U3828 (N_3828,N_1700,N_1588);
or U3829 (N_3829,N_1759,N_1649);
nand U3830 (N_3830,N_903,N_437);
nor U3831 (N_3831,N_448,N_734);
xnor U3832 (N_3832,N_1791,N_1214);
nand U3833 (N_3833,N_551,N_1823);
and U3834 (N_3834,N_1278,N_743);
nor U3835 (N_3835,N_687,N_78);
nor U3836 (N_3836,N_990,N_1645);
nand U3837 (N_3837,N_272,N_867);
or U3838 (N_3838,N_6,N_631);
nor U3839 (N_3839,N_330,N_114);
nand U3840 (N_3840,N_1987,N_1622);
nand U3841 (N_3841,N_206,N_11);
nor U3842 (N_3842,N_30,N_1595);
or U3843 (N_3843,N_298,N_150);
nand U3844 (N_3844,N_1604,N_1602);
nand U3845 (N_3845,N_1558,N_717);
nand U3846 (N_3846,N_76,N_1584);
nor U3847 (N_3847,N_1583,N_1653);
nor U3848 (N_3848,N_1852,N_1039);
and U3849 (N_3849,N_243,N_1374);
nand U3850 (N_3850,N_1941,N_1015);
or U3851 (N_3851,N_1367,N_118);
nand U3852 (N_3852,N_41,N_1318);
nor U3853 (N_3853,N_1457,N_466);
nand U3854 (N_3854,N_499,N_865);
or U3855 (N_3855,N_1594,N_1811);
nand U3856 (N_3856,N_28,N_983);
nor U3857 (N_3857,N_1366,N_675);
nand U3858 (N_3858,N_853,N_1246);
or U3859 (N_3859,N_1504,N_1652);
nor U3860 (N_3860,N_1161,N_543);
nor U3861 (N_3861,N_51,N_1669);
and U3862 (N_3862,N_1929,N_158);
nor U3863 (N_3863,N_510,N_407);
or U3864 (N_3864,N_1991,N_1060);
or U3865 (N_3865,N_1551,N_1406);
or U3866 (N_3866,N_1670,N_263);
and U3867 (N_3867,N_1989,N_1156);
nor U3868 (N_3868,N_572,N_630);
or U3869 (N_3869,N_775,N_1401);
nor U3870 (N_3870,N_405,N_1813);
or U3871 (N_3871,N_1518,N_1416);
nand U3872 (N_3872,N_1273,N_494);
or U3873 (N_3873,N_486,N_1679);
and U3874 (N_3874,N_366,N_1363);
xnor U3875 (N_3875,N_1282,N_1977);
or U3876 (N_3876,N_945,N_943);
nor U3877 (N_3877,N_434,N_327);
nor U3878 (N_3878,N_1314,N_1703);
nor U3879 (N_3879,N_1321,N_160);
nor U3880 (N_3880,N_456,N_1880);
and U3881 (N_3881,N_1158,N_1837);
and U3882 (N_3882,N_980,N_1280);
nor U3883 (N_3883,N_1466,N_1719);
nand U3884 (N_3884,N_1402,N_1704);
nand U3885 (N_3885,N_953,N_1747);
nor U3886 (N_3886,N_1892,N_948);
and U3887 (N_3887,N_651,N_1939);
or U3888 (N_3888,N_1626,N_782);
nor U3889 (N_3889,N_730,N_1837);
nand U3890 (N_3890,N_1878,N_102);
nor U3891 (N_3891,N_349,N_905);
or U3892 (N_3892,N_614,N_1747);
and U3893 (N_3893,N_1900,N_1142);
nor U3894 (N_3894,N_541,N_1546);
nand U3895 (N_3895,N_534,N_1662);
and U3896 (N_3896,N_1142,N_1687);
or U3897 (N_3897,N_1237,N_1626);
or U3898 (N_3898,N_578,N_1635);
or U3899 (N_3899,N_519,N_737);
and U3900 (N_3900,N_1980,N_287);
xor U3901 (N_3901,N_777,N_664);
xnor U3902 (N_3902,N_1306,N_1965);
xnor U3903 (N_3903,N_704,N_431);
and U3904 (N_3904,N_1680,N_259);
nand U3905 (N_3905,N_915,N_1312);
and U3906 (N_3906,N_536,N_1387);
or U3907 (N_3907,N_575,N_928);
nand U3908 (N_3908,N_92,N_486);
nor U3909 (N_3909,N_1821,N_1008);
or U3910 (N_3910,N_659,N_643);
or U3911 (N_3911,N_1159,N_797);
nor U3912 (N_3912,N_154,N_1889);
nor U3913 (N_3913,N_150,N_371);
nand U3914 (N_3914,N_893,N_1891);
or U3915 (N_3915,N_92,N_663);
nor U3916 (N_3916,N_1579,N_485);
nand U3917 (N_3917,N_10,N_1939);
nor U3918 (N_3918,N_1045,N_1575);
nor U3919 (N_3919,N_839,N_589);
and U3920 (N_3920,N_1963,N_1890);
and U3921 (N_3921,N_1678,N_224);
nand U3922 (N_3922,N_777,N_560);
or U3923 (N_3923,N_1841,N_505);
and U3924 (N_3924,N_1765,N_1718);
nand U3925 (N_3925,N_234,N_1167);
xnor U3926 (N_3926,N_387,N_1701);
nand U3927 (N_3927,N_1194,N_431);
and U3928 (N_3928,N_434,N_1449);
nor U3929 (N_3929,N_910,N_976);
nand U3930 (N_3930,N_255,N_587);
nand U3931 (N_3931,N_371,N_498);
nand U3932 (N_3932,N_1121,N_189);
or U3933 (N_3933,N_1962,N_144);
nor U3934 (N_3934,N_1443,N_16);
or U3935 (N_3935,N_293,N_1089);
xnor U3936 (N_3936,N_1495,N_347);
nor U3937 (N_3937,N_226,N_1409);
xor U3938 (N_3938,N_576,N_1422);
nand U3939 (N_3939,N_1108,N_1303);
nand U3940 (N_3940,N_248,N_197);
nand U3941 (N_3941,N_394,N_1939);
and U3942 (N_3942,N_1736,N_882);
nor U3943 (N_3943,N_123,N_1152);
or U3944 (N_3944,N_39,N_412);
or U3945 (N_3945,N_1184,N_43);
or U3946 (N_3946,N_1741,N_292);
and U3947 (N_3947,N_1672,N_245);
or U3948 (N_3948,N_1055,N_1392);
and U3949 (N_3949,N_1153,N_1684);
and U3950 (N_3950,N_1694,N_1256);
xor U3951 (N_3951,N_1261,N_1819);
xor U3952 (N_3952,N_1882,N_851);
and U3953 (N_3953,N_15,N_1193);
nand U3954 (N_3954,N_1927,N_261);
and U3955 (N_3955,N_1578,N_876);
and U3956 (N_3956,N_1760,N_128);
or U3957 (N_3957,N_314,N_187);
nand U3958 (N_3958,N_1854,N_1406);
nor U3959 (N_3959,N_891,N_148);
nand U3960 (N_3960,N_1300,N_86);
and U3961 (N_3961,N_1600,N_1583);
nor U3962 (N_3962,N_1325,N_828);
nor U3963 (N_3963,N_1358,N_507);
or U3964 (N_3964,N_430,N_1412);
xor U3965 (N_3965,N_1729,N_832);
xnor U3966 (N_3966,N_220,N_1857);
nor U3967 (N_3967,N_1203,N_348);
nand U3968 (N_3968,N_1767,N_859);
nor U3969 (N_3969,N_917,N_1089);
nor U3970 (N_3970,N_205,N_1895);
xnor U3971 (N_3971,N_265,N_57);
xor U3972 (N_3972,N_856,N_1264);
nor U3973 (N_3973,N_1984,N_1333);
nand U3974 (N_3974,N_102,N_389);
nand U3975 (N_3975,N_652,N_1263);
xor U3976 (N_3976,N_195,N_704);
and U3977 (N_3977,N_564,N_1844);
nor U3978 (N_3978,N_1714,N_1666);
or U3979 (N_3979,N_1774,N_770);
nand U3980 (N_3980,N_1929,N_1343);
and U3981 (N_3981,N_973,N_1527);
nor U3982 (N_3982,N_1373,N_1678);
nand U3983 (N_3983,N_1798,N_1500);
xnor U3984 (N_3984,N_1518,N_862);
or U3985 (N_3985,N_1157,N_388);
nand U3986 (N_3986,N_1970,N_1168);
nor U3987 (N_3987,N_1527,N_892);
and U3988 (N_3988,N_978,N_628);
nand U3989 (N_3989,N_1491,N_731);
xor U3990 (N_3990,N_850,N_791);
or U3991 (N_3991,N_1930,N_236);
nor U3992 (N_3992,N_985,N_705);
nor U3993 (N_3993,N_1459,N_697);
nand U3994 (N_3994,N_860,N_1844);
or U3995 (N_3995,N_518,N_1710);
nor U3996 (N_3996,N_1828,N_608);
nor U3997 (N_3997,N_1099,N_721);
xor U3998 (N_3998,N_1633,N_1445);
and U3999 (N_3999,N_967,N_200);
nor U4000 (N_4000,N_2264,N_3912);
or U4001 (N_4001,N_2263,N_2925);
xnor U4002 (N_4002,N_2183,N_3235);
nor U4003 (N_4003,N_3531,N_2245);
nor U4004 (N_4004,N_3830,N_3353);
nand U4005 (N_4005,N_3389,N_3315);
or U4006 (N_4006,N_2537,N_2572);
and U4007 (N_4007,N_2820,N_3826);
nand U4008 (N_4008,N_2712,N_2548);
nand U4009 (N_4009,N_3984,N_2045);
nand U4010 (N_4010,N_2160,N_2012);
and U4011 (N_4011,N_2413,N_2610);
and U4012 (N_4012,N_2911,N_2268);
nor U4013 (N_4013,N_3714,N_3589);
or U4014 (N_4014,N_3587,N_2654);
or U4015 (N_4015,N_2318,N_3644);
and U4016 (N_4016,N_2280,N_3579);
and U4017 (N_4017,N_3536,N_2667);
nand U4018 (N_4018,N_2860,N_3020);
or U4019 (N_4019,N_3187,N_2068);
xor U4020 (N_4020,N_2727,N_3227);
nand U4021 (N_4021,N_2951,N_3230);
or U4022 (N_4022,N_3150,N_2660);
nand U4023 (N_4023,N_3567,N_3648);
nand U4024 (N_4024,N_3670,N_2612);
or U4025 (N_4025,N_3435,N_3053);
and U4026 (N_4026,N_3005,N_3094);
nor U4027 (N_4027,N_2720,N_2096);
nand U4028 (N_4028,N_2279,N_3026);
nor U4029 (N_4029,N_3114,N_3024);
and U4030 (N_4030,N_3818,N_3701);
nand U4031 (N_4031,N_3911,N_3904);
xnor U4032 (N_4032,N_3241,N_3327);
and U4033 (N_4033,N_3110,N_2958);
nor U4034 (N_4034,N_2740,N_3845);
nor U4035 (N_4035,N_3906,N_3564);
nor U4036 (N_4036,N_3664,N_3250);
nand U4037 (N_4037,N_3465,N_3238);
nor U4038 (N_4038,N_2946,N_2228);
xnor U4039 (N_4039,N_2367,N_2906);
nand U4040 (N_4040,N_3057,N_3926);
nor U4041 (N_4041,N_2580,N_3101);
and U4042 (N_4042,N_3655,N_3352);
and U4043 (N_4043,N_2379,N_3388);
and U4044 (N_4044,N_3673,N_2645);
nand U4045 (N_4045,N_3379,N_3442);
nand U4046 (N_4046,N_3509,N_2035);
and U4047 (N_4047,N_2386,N_2262);
or U4048 (N_4048,N_2256,N_2078);
nand U4049 (N_4049,N_2493,N_3786);
or U4050 (N_4050,N_3975,N_3526);
and U4051 (N_4051,N_2478,N_2728);
nor U4052 (N_4052,N_3491,N_2331);
nand U4053 (N_4053,N_3406,N_2968);
and U4054 (N_4054,N_3718,N_3074);
xnor U4055 (N_4055,N_3134,N_3656);
nor U4056 (N_4056,N_3482,N_3633);
and U4057 (N_4057,N_3600,N_2206);
and U4058 (N_4058,N_3597,N_2498);
nand U4059 (N_4059,N_2663,N_3783);
nor U4060 (N_4060,N_3470,N_3928);
and U4061 (N_4061,N_3625,N_2527);
nor U4062 (N_4062,N_3382,N_2603);
nand U4063 (N_4063,N_2803,N_3619);
and U4064 (N_4064,N_3762,N_2056);
and U4065 (N_4065,N_2781,N_2565);
nor U4066 (N_4066,N_2444,N_3612);
nand U4067 (N_4067,N_3072,N_3804);
and U4068 (N_4068,N_2204,N_3934);
nor U4069 (N_4069,N_3437,N_3041);
xor U4070 (N_4070,N_2482,N_2446);
nand U4071 (N_4071,N_3948,N_2615);
nor U4072 (N_4072,N_2836,N_3583);
nor U4073 (N_4073,N_3985,N_3098);
nand U4074 (N_4074,N_2541,N_3331);
or U4075 (N_4075,N_3481,N_2196);
nand U4076 (N_4076,N_2486,N_2774);
or U4077 (N_4077,N_2534,N_2451);
and U4078 (N_4078,N_2465,N_2161);
xor U4079 (N_4079,N_2172,N_2773);
nor U4080 (N_4080,N_2062,N_3766);
nor U4081 (N_4081,N_3444,N_3538);
nand U4082 (N_4082,N_3314,N_2705);
and U4083 (N_4083,N_3002,N_3181);
nor U4084 (N_4084,N_3245,N_2169);
or U4085 (N_4085,N_3412,N_2481);
xor U4086 (N_4086,N_2164,N_3304);
nor U4087 (N_4087,N_2868,N_2361);
xor U4088 (N_4088,N_3558,N_2363);
nor U4089 (N_4089,N_2560,N_3015);
or U4090 (N_4090,N_3447,N_3096);
nand U4091 (N_4091,N_3390,N_2333);
and U4092 (N_4092,N_2653,N_3522);
nand U4093 (N_4093,N_3854,N_3294);
or U4094 (N_4094,N_2144,N_3305);
nor U4095 (N_4095,N_2207,N_2223);
xnor U4096 (N_4096,N_2730,N_3006);
or U4097 (N_4097,N_2057,N_2186);
and U4098 (N_4098,N_3690,N_3556);
nand U4099 (N_4099,N_3130,N_3265);
and U4100 (N_4100,N_2244,N_3219);
and U4101 (N_4101,N_2726,N_3149);
or U4102 (N_4102,N_3708,N_2892);
nor U4103 (N_4103,N_3994,N_3752);
nor U4104 (N_4104,N_2532,N_2350);
nand U4105 (N_4105,N_3270,N_2903);
nor U4106 (N_4106,N_3523,N_3812);
nor U4107 (N_4107,N_3127,N_3322);
and U4108 (N_4108,N_3989,N_2549);
and U4109 (N_4109,N_2804,N_3107);
or U4110 (N_4110,N_2900,N_2994);
nor U4111 (N_4111,N_3894,N_3582);
or U4112 (N_4112,N_2355,N_2880);
nor U4113 (N_4113,N_2636,N_2990);
nor U4114 (N_4114,N_3809,N_3419);
or U4115 (N_4115,N_3061,N_3030);
nor U4116 (N_4116,N_2780,N_3950);
and U4117 (N_4117,N_3362,N_2054);
or U4118 (N_4118,N_3261,N_2469);
nor U4119 (N_4119,N_2273,N_3418);
xor U4120 (N_4120,N_3368,N_2631);
nor U4121 (N_4121,N_3882,N_2225);
nor U4122 (N_4122,N_3800,N_2119);
nand U4123 (N_4123,N_2673,N_3915);
or U4124 (N_4124,N_2468,N_3172);
nor U4125 (N_4125,N_3229,N_2487);
nand U4126 (N_4126,N_3770,N_3590);
nor U4127 (N_4127,N_2723,N_2991);
or U4128 (N_4128,N_3682,N_2102);
or U4129 (N_4129,N_2201,N_3913);
nor U4130 (N_4130,N_3276,N_3960);
nor U4131 (N_4131,N_2103,N_3152);
or U4132 (N_4132,N_2180,N_3477);
and U4133 (N_4133,N_3855,N_2809);
or U4134 (N_4134,N_2199,N_2743);
xnor U4135 (N_4135,N_2592,N_3677);
nand U4136 (N_4136,N_2176,N_2619);
or U4137 (N_4137,N_3453,N_3236);
xnor U4138 (N_4138,N_2767,N_3196);
and U4139 (N_4139,N_3341,N_2766);
nor U4140 (N_4140,N_3469,N_2236);
or U4141 (N_4141,N_3742,N_3267);
nor U4142 (N_4142,N_2757,N_3262);
or U4143 (N_4143,N_2323,N_3844);
nor U4144 (N_4144,N_3285,N_3986);
or U4145 (N_4145,N_3649,N_3776);
or U4146 (N_4146,N_3175,N_3425);
or U4147 (N_4147,N_3339,N_2686);
and U4148 (N_4148,N_2491,N_3448);
or U4149 (N_4149,N_2751,N_3909);
and U4150 (N_4150,N_3260,N_2764);
nand U4151 (N_4151,N_2590,N_3155);
xnor U4152 (N_4152,N_3822,N_2396);
nand U4153 (N_4153,N_2389,N_2126);
nor U4154 (N_4154,N_2055,N_3585);
or U4155 (N_4155,N_2430,N_2229);
or U4156 (N_4156,N_3694,N_2644);
nand U4157 (N_4157,N_3474,N_2883);
nand U4158 (N_4158,N_2179,N_3970);
nand U4159 (N_4159,N_3386,N_2564);
and U4160 (N_4160,N_2406,N_3334);
and U4161 (N_4161,N_3720,N_2587);
xnor U4162 (N_4162,N_3638,N_2738);
nor U4163 (N_4163,N_2373,N_2147);
nor U4164 (N_4164,N_3029,N_3955);
and U4165 (N_4165,N_2693,N_2974);
nor U4166 (N_4166,N_3188,N_2511);
or U4167 (N_4167,N_2390,N_3088);
nand U4168 (N_4168,N_2477,N_3431);
and U4169 (N_4169,N_2332,N_3925);
and U4170 (N_4170,N_2168,N_3884);
nand U4171 (N_4171,N_2539,N_3560);
or U4172 (N_4172,N_2334,N_2979);
and U4173 (N_4173,N_2301,N_2438);
and U4174 (N_4174,N_3798,N_2167);
nand U4175 (N_4175,N_3949,N_3892);
and U4176 (N_4176,N_3578,N_2701);
nor U4177 (N_4177,N_3710,N_2724);
nor U4178 (N_4178,N_3539,N_2942);
nor U4179 (N_4179,N_3111,N_2790);
or U4180 (N_4180,N_3348,N_3290);
and U4181 (N_4181,N_2247,N_2448);
nor U4182 (N_4182,N_3961,N_2075);
or U4183 (N_4183,N_3132,N_3008);
or U4184 (N_4184,N_2959,N_2533);
xor U4185 (N_4185,N_3212,N_3043);
or U4186 (N_4186,N_2138,N_3865);
nand U4187 (N_4187,N_3457,N_3896);
nand U4188 (N_4188,N_2688,N_3325);
and U4189 (N_4189,N_3190,N_2544);
nor U4190 (N_4190,N_3036,N_3163);
or U4191 (N_4191,N_2173,N_3086);
nor U4192 (N_4192,N_2205,N_3856);
or U4193 (N_4193,N_2776,N_3863);
xnor U4194 (N_4194,N_2913,N_2190);
and U4195 (N_4195,N_3031,N_2193);
nand U4196 (N_4196,N_2664,N_2876);
or U4197 (N_4197,N_2340,N_3692);
nand U4198 (N_4198,N_2414,N_2188);
and U4199 (N_4199,N_3778,N_2581);
or U4200 (N_4200,N_3974,N_2029);
nor U4201 (N_4201,N_3405,N_2710);
and U4202 (N_4202,N_3839,N_3032);
or U4203 (N_4203,N_2137,N_3116);
nor U4204 (N_4204,N_3022,N_3781);
nand U4205 (N_4205,N_3432,N_3608);
nand U4206 (N_4206,N_2508,N_2437);
nor U4207 (N_4207,N_2681,N_2346);
nor U4208 (N_4208,N_3623,N_2195);
or U4209 (N_4209,N_3940,N_2013);
nand U4210 (N_4210,N_2509,N_3381);
nor U4211 (N_4211,N_2671,N_2989);
or U4212 (N_4212,N_2426,N_3436);
nand U4213 (N_4213,N_3805,N_3537);
nor U4214 (N_4214,N_2306,N_3183);
nand U4215 (N_4215,N_3185,N_2220);
and U4216 (N_4216,N_2079,N_2197);
nand U4217 (N_4217,N_3021,N_2022);
and U4218 (N_4218,N_2303,N_2573);
nor U4219 (N_4219,N_2211,N_3028);
and U4220 (N_4220,N_3460,N_2635);
nor U4221 (N_4221,N_3900,N_3545);
nor U4222 (N_4222,N_3395,N_3886);
nor U4223 (N_4223,N_3282,N_3999);
nand U4224 (N_4224,N_2234,N_2066);
nand U4225 (N_4225,N_2908,N_3297);
xnor U4226 (N_4226,N_3197,N_2521);
nand U4227 (N_4227,N_3392,N_2977);
or U4228 (N_4228,N_2058,N_3988);
or U4229 (N_4229,N_2352,N_2338);
nand U4230 (N_4230,N_3991,N_2392);
or U4231 (N_4231,N_2359,N_2779);
or U4232 (N_4232,N_2484,N_2998);
nor U4233 (N_4233,N_3434,N_3815);
and U4234 (N_4234,N_3166,N_2091);
or U4235 (N_4235,N_2744,N_3695);
and U4236 (N_4236,N_2450,N_2100);
nor U4237 (N_4237,N_3897,N_3174);
and U4238 (N_4238,N_2494,N_2313);
nand U4239 (N_4239,N_2812,N_2973);
nand U4240 (N_4240,N_3128,N_2621);
xnor U4241 (N_4241,N_2695,N_3240);
nand U4242 (N_4242,N_3200,N_3280);
nor U4243 (N_4243,N_2421,N_2125);
or U4244 (N_4244,N_2765,N_2371);
nor U4245 (N_4245,N_2042,N_2275);
nor U4246 (N_4246,N_3492,N_2528);
or U4247 (N_4247,N_2053,N_3433);
nand U4248 (N_4248,N_2046,N_2856);
and U4249 (N_4249,N_2285,N_2741);
xor U4250 (N_4250,N_2237,N_3478);
nand U4251 (N_4251,N_3000,N_3058);
nand U4252 (N_4252,N_2966,N_3159);
nor U4253 (N_4253,N_3874,N_3441);
nand U4254 (N_4254,N_3452,N_2174);
or U4255 (N_4255,N_3971,N_2000);
xnor U4256 (N_4256,N_3832,N_2006);
and U4257 (N_4257,N_3295,N_2203);
and U4258 (N_4258,N_3209,N_2047);
nand U4259 (N_4259,N_2086,N_2525);
nor U4260 (N_4260,N_3003,N_2970);
and U4261 (N_4261,N_2939,N_3108);
xnor U4262 (N_4262,N_3703,N_3121);
nand U4263 (N_4263,N_2092,N_2602);
nor U4264 (N_4264,N_3363,N_3272);
xor U4265 (N_4265,N_3841,N_3979);
nand U4266 (N_4266,N_2089,N_2192);
nand U4267 (N_4267,N_3248,N_2052);
nand U4268 (N_4268,N_2420,N_3602);
nor U4269 (N_4269,N_3320,N_2375);
xnor U4270 (N_4270,N_2133,N_2018);
or U4271 (N_4271,N_3011,N_2784);
nor U4272 (N_4272,N_3510,N_3929);
and U4273 (N_4273,N_3728,N_2044);
xnor U4274 (N_4274,N_3997,N_2788);
nand U4275 (N_4275,N_3157,N_3931);
and U4276 (N_4276,N_3415,N_2616);
nand U4277 (N_4277,N_2988,N_2269);
nor U4278 (N_4278,N_3551,N_2422);
and U4279 (N_4279,N_3787,N_3888);
or U4280 (N_4280,N_3996,N_2630);
nor U4281 (N_4281,N_3790,N_3427);
nand U4282 (N_4282,N_3730,N_2661);
xnor U4283 (N_4283,N_2077,N_2297);
xnor U4284 (N_4284,N_2224,N_2395);
or U4285 (N_4285,N_3524,N_3729);
nor U4286 (N_4286,N_2149,N_2382);
nor U4287 (N_4287,N_3713,N_3374);
or U4288 (N_4288,N_2251,N_3868);
nor U4289 (N_4289,N_3621,N_2216);
nand U4290 (N_4290,N_3289,N_3488);
or U4291 (N_4291,N_2087,N_2659);
nor U4292 (N_4292,N_2575,N_3191);
xor U4293 (N_4293,N_2171,N_3326);
nand U4294 (N_4294,N_2036,N_2956);
and U4295 (N_4295,N_2709,N_2698);
xor U4296 (N_4296,N_2597,N_2407);
or U4297 (N_4297,N_3548,N_2680);
nand U4298 (N_4298,N_2342,N_2433);
and U4299 (N_4299,N_2372,N_2867);
and U4300 (N_4300,N_2315,N_3731);
and U4301 (N_4301,N_3932,N_2215);
or U4302 (N_4302,N_2230,N_2349);
xnor U4303 (N_4303,N_2076,N_2424);
and U4304 (N_4304,N_3485,N_3658);
or U4305 (N_4305,N_2344,N_3286);
nor U4306 (N_4306,N_2309,N_3689);
and U4307 (N_4307,N_3377,N_3120);
nor U4308 (N_4308,N_2449,N_2440);
or U4309 (N_4309,N_3062,N_3115);
xnor U4310 (N_4310,N_3652,N_2807);
nor U4311 (N_4311,N_2328,N_2129);
and U4312 (N_4312,N_2785,N_2010);
nand U4313 (N_4313,N_3050,N_3243);
or U4314 (N_4314,N_3685,N_3169);
nor U4315 (N_4315,N_2591,N_3806);
nand U4316 (N_4316,N_2882,N_3136);
and U4317 (N_4317,N_3498,N_3561);
or U4318 (N_4318,N_2760,N_2145);
or U4319 (N_4319,N_3264,N_3821);
nor U4320 (N_4320,N_3942,N_2898);
nand U4321 (N_4321,N_2711,N_3721);
xor U4322 (N_4322,N_2948,N_3093);
or U4323 (N_4323,N_2748,N_3137);
and U4324 (N_4324,N_3751,N_2975);
or U4325 (N_4325,N_3833,N_3849);
nand U4326 (N_4326,N_2069,N_3025);
and U4327 (N_4327,N_2950,N_2854);
nand U4328 (N_4328,N_3953,N_3586);
or U4329 (N_4329,N_3253,N_3789);
or U4330 (N_4330,N_3275,N_3758);
or U4331 (N_4331,N_3601,N_3407);
nand U4332 (N_4332,N_3933,N_3700);
nor U4333 (N_4333,N_2397,N_3400);
or U4334 (N_4334,N_2996,N_3373);
or U4335 (N_4335,N_2428,N_3919);
nand U4336 (N_4336,N_2887,N_2495);
nand U4337 (N_4337,N_3078,N_2540);
nand U4338 (N_4338,N_3562,N_2480);
xnor U4339 (N_4339,N_2387,N_2289);
nor U4340 (N_4340,N_2271,N_2543);
and U4341 (N_4341,N_3962,N_3165);
nand U4342 (N_4342,N_3440,N_2846);
or U4343 (N_4343,N_2747,N_3383);
nor U4344 (N_4344,N_3458,N_3799);
and U4345 (N_4345,N_3099,N_3541);
or U4346 (N_4346,N_2002,N_3736);
nor U4347 (N_4347,N_2965,N_3836);
and U4348 (N_4348,N_2797,N_3085);
and U4349 (N_4349,N_3105,N_2634);
xnor U4350 (N_4350,N_2618,N_3313);
or U4351 (N_4351,N_2370,N_2090);
nand U4352 (N_4352,N_3614,N_3027);
or U4353 (N_4353,N_2897,N_3279);
or U4354 (N_4354,N_2071,N_3636);
and U4355 (N_4355,N_3891,N_2310);
nand U4356 (N_4356,N_3641,N_3018);
or U4357 (N_4357,N_3178,N_2669);
nand U4358 (N_4358,N_3659,N_2853);
or U4359 (N_4359,N_3372,N_3360);
and U4360 (N_4360,N_3042,N_2683);
nand U4361 (N_4361,N_3611,N_3486);
and U4362 (N_4362,N_3687,N_2322);
nand U4363 (N_4363,N_3794,N_2550);
and U4364 (N_4364,N_3040,N_3347);
nand U4365 (N_4365,N_3249,N_2625);
or U4366 (N_4366,N_3255,N_2556);
or U4367 (N_4367,N_2749,N_3618);
nor U4368 (N_4368,N_3009,N_2113);
nand U4369 (N_4369,N_2926,N_3983);
or U4370 (N_4370,N_2376,N_2873);
nand U4371 (N_4371,N_2722,N_2388);
nand U4372 (N_4372,N_2796,N_2500);
nand U4373 (N_4373,N_2460,N_2954);
or U4374 (N_4374,N_2647,N_2825);
or U4375 (N_4375,N_2443,N_3139);
and U4376 (N_4376,N_3755,N_2835);
nor U4377 (N_4377,N_3176,N_2027);
nor U4378 (N_4378,N_2104,N_2253);
and U4379 (N_4379,N_3901,N_3142);
nand U4380 (N_4380,N_3980,N_3661);
nand U4381 (N_4381,N_3860,N_3813);
nor U4382 (N_4382,N_3870,N_2899);
or U4383 (N_4383,N_2858,N_3936);
nand U4384 (N_4384,N_3719,N_2462);
nor U4385 (N_4385,N_3547,N_2969);
nand U4386 (N_4386,N_3312,N_3033);
nor U4387 (N_4387,N_3759,N_2763);
and U4388 (N_4388,N_2304,N_2916);
or U4389 (N_4389,N_3967,N_3610);
or U4390 (N_4390,N_2353,N_3080);
xnor U4391 (N_4391,N_2512,N_2132);
or U4392 (N_4392,N_2336,N_3472);
and U4393 (N_4393,N_2707,N_2298);
nand U4394 (N_4394,N_2431,N_2839);
nor U4395 (N_4395,N_2101,N_3647);
nand U4396 (N_4396,N_2305,N_3634);
and U4397 (N_4397,N_3557,N_3242);
nor U4398 (N_4398,N_3193,N_3076);
nand U4399 (N_4399,N_2547,N_3630);
nor U4400 (N_4400,N_2829,N_2259);
and U4401 (N_4401,N_2717,N_2294);
nand U4402 (N_4402,N_2714,N_3244);
nand U4403 (N_4403,N_3274,N_2039);
or U4404 (N_4404,N_3646,N_2885);
and U4405 (N_4405,N_2281,N_2246);
or U4406 (N_4406,N_2459,N_3215);
xor U4407 (N_4407,N_2593,N_2063);
or U4408 (N_4408,N_3801,N_2151);
or U4409 (N_4409,N_2070,N_2718);
nor U4410 (N_4410,N_2739,N_2243);
or U4411 (N_4411,N_3224,N_2212);
and U4412 (N_4412,N_3459,N_2745);
or U4413 (N_4413,N_3259,N_3233);
nor U4414 (N_4414,N_2335,N_3739);
nor U4415 (N_4415,N_2217,N_2816);
nand U4416 (N_4416,N_2594,N_2288);
and U4417 (N_4417,N_3131,N_2770);
and U4418 (N_4418,N_3495,N_3292);
and U4419 (N_4419,N_2348,N_2366);
nand U4420 (N_4420,N_3034,N_2938);
nor U4421 (N_4421,N_3283,N_3421);
xnor U4422 (N_4422,N_3993,N_2665);
nand U4423 (N_4423,N_2598,N_2737);
and U4424 (N_4424,N_2474,N_2249);
xor U4425 (N_4425,N_3850,N_2209);
or U4426 (N_4426,N_3550,N_3908);
and U4427 (N_4427,N_3047,N_2202);
nor U4428 (N_4428,N_2270,N_3698);
and U4429 (N_4429,N_3463,N_3063);
nor U4430 (N_4430,N_2629,N_3113);
nor U4431 (N_4431,N_2687,N_2073);
or U4432 (N_4432,N_3881,N_3054);
nand U4433 (N_4433,N_3905,N_2095);
or U4434 (N_4434,N_3699,N_2672);
nor U4435 (N_4435,N_3167,N_2893);
xor U4436 (N_4436,N_2326,N_3898);
and U4437 (N_4437,N_3073,N_3605);
and U4438 (N_4438,N_2034,N_3676);
xnor U4439 (N_4439,N_2756,N_2143);
nand U4440 (N_4440,N_3145,N_2128);
nor U4441 (N_4441,N_2472,N_3254);
and U4442 (N_4442,N_2242,N_3198);
or U4443 (N_4443,N_3958,N_2291);
nand U4444 (N_4444,N_2553,N_3769);
and U4445 (N_4445,N_3082,N_3173);
and U4446 (N_4446,N_2185,N_3091);
nor U4447 (N_4447,N_3365,N_3384);
and U4448 (N_4448,N_3490,N_3171);
or U4449 (N_4449,N_3965,N_3875);
nand U4450 (N_4450,N_2813,N_3774);
xor U4451 (N_4451,N_3743,N_2166);
nor U4452 (N_4452,N_3247,N_2404);
or U4453 (N_4453,N_2872,N_2381);
and U4454 (N_4454,N_2753,N_3329);
nor U4455 (N_4455,N_3122,N_3473);
and U4456 (N_4456,N_3504,N_3394);
and U4457 (N_4457,N_2945,N_2589);
xnor U4458 (N_4458,N_2731,N_3371);
or U4459 (N_4459,N_2850,N_3640);
nor U4460 (N_4460,N_2463,N_2093);
and U4461 (N_4461,N_3179,N_3154);
xor U4462 (N_4462,N_2447,N_3861);
nand U4463 (N_4463,N_3109,N_2725);
or U4464 (N_4464,N_2983,N_3414);
xor U4465 (N_4465,N_3937,N_2507);
nor U4466 (N_4466,N_3112,N_3271);
nand U4467 (N_4467,N_2577,N_2308);
nor U4468 (N_4468,N_3866,N_2522);
nor U4469 (N_4469,N_3506,N_3069);
nor U4470 (N_4470,N_3624,N_2456);
nor U4471 (N_4471,N_3513,N_3924);
and U4472 (N_4472,N_3525,N_3143);
nand U4473 (N_4473,N_2750,N_2524);
nand U4474 (N_4474,N_3375,N_2520);
nor U4475 (N_4475,N_3129,N_2265);
nor U4476 (N_4476,N_2218,N_3420);
nand U4477 (N_4477,N_2116,N_2148);
nor U4478 (N_4478,N_2542,N_2231);
or U4479 (N_4479,N_2260,N_3681);
nand U4480 (N_4480,N_3825,N_3837);
nand U4481 (N_4481,N_3257,N_2620);
xnor U4482 (N_4482,N_2184,N_3594);
nand U4483 (N_4483,N_3571,N_3065);
nand U4484 (N_4484,N_2385,N_2499);
nand U4485 (N_4485,N_2768,N_2538);
and U4486 (N_4486,N_3705,N_3549);
or U4487 (N_4487,N_3530,N_3319);
and U4488 (N_4488,N_2142,N_2841);
and U4489 (N_4489,N_2402,N_2886);
or U4490 (N_4490,N_3734,N_3318);
nor U4491 (N_4491,N_2696,N_2896);
nand U4492 (N_4492,N_2985,N_3867);
or U4493 (N_4493,N_3738,N_2295);
nand U4494 (N_4494,N_2378,N_2358);
nand U4495 (N_4495,N_3396,N_3588);
nand U4496 (N_4496,N_2189,N_2429);
or U4497 (N_4497,N_3876,N_3717);
xor U4498 (N_4498,N_3727,N_3263);
and U4499 (N_4499,N_2139,N_3449);
xnor U4500 (N_4500,N_2869,N_2578);
nor U4501 (N_4501,N_3479,N_3317);
or U4502 (N_4502,N_3748,N_2808);
and U4503 (N_4503,N_3084,N_2962);
and U4504 (N_4504,N_3946,N_3660);
or U4505 (N_4505,N_2874,N_3534);
nor U4506 (N_4506,N_3309,N_2943);
or U4507 (N_4507,N_3168,N_2383);
or U4508 (N_4508,N_2457,N_2131);
nand U4509 (N_4509,N_3356,N_2937);
and U4510 (N_4510,N_3603,N_3234);
and U4511 (N_4511,N_3851,N_3767);
nand U4512 (N_4512,N_2831,N_2064);
nand U4513 (N_4513,N_2050,N_2108);
and U4514 (N_4514,N_2890,N_2011);
nor U4515 (N_4515,N_2250,N_2574);
and U4516 (N_4516,N_2905,N_3281);
and U4517 (N_4517,N_2865,N_3102);
nor U4518 (N_4518,N_2802,N_3753);
xor U4519 (N_4519,N_2277,N_3834);
or U4520 (N_4520,N_3496,N_2123);
nand U4521 (N_4521,N_3532,N_2464);
nand U4522 (N_4522,N_3987,N_2732);
or U4523 (N_4523,N_3877,N_2772);
nor U4524 (N_4524,N_2563,N_2826);
nor U4525 (N_4525,N_3429,N_2356);
xor U4526 (N_4526,N_2555,N_3293);
or U4527 (N_4527,N_3471,N_2844);
nor U4528 (N_4528,N_2670,N_3417);
nor U4529 (N_4529,N_2362,N_2442);
nor U4530 (N_4530,N_3346,N_2758);
and U4531 (N_4531,N_3296,N_2272);
nand U4532 (N_4532,N_3570,N_3443);
xnor U4533 (N_4533,N_2586,N_2157);
nand U4534 (N_4534,N_3828,N_3184);
and U4535 (N_4535,N_2238,N_3792);
or U4536 (N_4536,N_2585,N_3269);
nand U4537 (N_4537,N_3927,N_3461);
or U4538 (N_4538,N_2894,N_3123);
and U4539 (N_4539,N_3518,N_3182);
xnor U4540 (N_4540,N_3910,N_2944);
or U4541 (N_4541,N_2762,N_2657);
nand U4542 (N_4542,N_3380,N_3824);
xor U4543 (N_4543,N_2112,N_3740);
nor U4544 (N_4544,N_2266,N_2818);
and U4545 (N_4545,N_3378,N_2316);
nand U4546 (N_4546,N_3147,N_2552);
and U4547 (N_4547,N_2675,N_2649);
or U4548 (N_4548,N_2127,N_2441);
nand U4549 (N_4549,N_3723,N_2799);
xor U4550 (N_4550,N_2823,N_3077);
nand U4551 (N_4551,N_2007,N_2436);
nand U4552 (N_4552,N_2510,N_2999);
or U4553 (N_4553,N_3763,N_2041);
nor U4554 (N_4554,N_3203,N_3613);
or U4555 (N_4555,N_2300,N_3872);
or U4556 (N_4556,N_2651,N_2643);
nor U4557 (N_4557,N_3345,N_2445);
nand U4558 (N_4558,N_2235,N_3411);
nor U4559 (N_4559,N_3205,N_3565);
nor U4560 (N_4560,N_3141,N_2843);
and U4561 (N_4561,N_2656,N_2881);
xnor U4562 (N_4562,N_2226,N_3686);
xnor U4563 (N_4563,N_2855,N_2118);
xnor U4564 (N_4564,N_2130,N_2519);
nor U4565 (N_4565,N_3811,N_2200);
nand U4566 (N_4566,N_2170,N_2819);
and U4567 (N_4567,N_3941,N_3231);
or U4568 (N_4568,N_2163,N_2150);
or U4569 (N_4569,N_2208,N_3972);
or U4570 (N_4570,N_2191,N_3517);
nand U4571 (N_4571,N_2483,N_3413);
nand U4572 (N_4572,N_3945,N_3308);
xor U4573 (N_4573,N_3232,N_2614);
nor U4574 (N_4574,N_3858,N_2121);
or U4575 (N_4575,N_3192,N_3097);
xor U4576 (N_4576,N_3704,N_2554);
nor U4577 (N_4577,N_2889,N_3500);
and U4578 (N_4578,N_3544,N_3964);
nand U4579 (N_4579,N_3207,N_2324);
or U4580 (N_4580,N_2546,N_3829);
nor U4581 (N_4581,N_3878,N_3138);
nand U4582 (N_4582,N_3707,N_2637);
nor U4583 (N_4583,N_3678,N_3423);
or U4584 (N_4584,N_3568,N_2485);
nor U4585 (N_4585,N_3503,N_3773);
nor U4586 (N_4586,N_3838,N_3409);
and U4587 (N_4587,N_2003,N_2014);
and U4588 (N_4588,N_2755,N_2679);
nor U4589 (N_4589,N_2152,N_3788);
nor U4590 (N_4590,N_3765,N_2940);
nand U4591 (N_4591,N_3978,N_3848);
or U4592 (N_4592,N_3737,N_2703);
nor U4593 (N_4593,N_3505,N_2049);
xor U4594 (N_4594,N_2364,N_2771);
and U4595 (N_4595,N_2307,N_3842);
nor U4596 (N_4596,N_3369,N_3401);
and U4597 (N_4597,N_2467,N_3403);
nor U4598 (N_4598,N_2165,N_3637);
nand U4599 (N_4599,N_3218,N_2488);
nor U4600 (N_4600,N_2141,N_2697);
and U4601 (N_4601,N_3328,N_3059);
nor U4602 (N_4602,N_2933,N_2452);
and U4603 (N_4603,N_3302,N_3399);
xor U4604 (N_4604,N_3747,N_2221);
nand U4605 (N_4605,N_2059,N_3998);
and U4606 (N_4606,N_3336,N_3733);
or U4607 (N_4607,N_2792,N_2479);
or U4608 (N_4608,N_2972,N_2506);
and U4609 (N_4609,N_2648,N_3591);
xor U4610 (N_4610,N_3990,N_3595);
or U4611 (N_4611,N_2814,N_2729);
and U4612 (N_4612,N_2607,N_3273);
and U4613 (N_4613,N_3756,N_2658);
nor U4614 (N_4614,N_3439,N_2501);
or U4615 (N_4615,N_3220,N_2817);
nor U4616 (N_4616,N_3760,N_3217);
nand U4617 (N_4617,N_3816,N_2162);
and U4618 (N_4618,N_2061,N_2453);
and U4619 (N_4619,N_2734,N_3351);
nor U4620 (N_4620,N_2953,N_3117);
nand U4621 (N_4621,N_2932,N_2470);
nor U4622 (N_4622,N_2158,N_2733);
nor U4623 (N_4623,N_2502,N_3785);
nor U4624 (N_4624,N_2713,N_2489);
nor U4625 (N_4625,N_2909,N_3424);
or U4626 (N_4626,N_3079,N_2072);
nand U4627 (N_4627,N_2283,N_3391);
nor U4628 (N_4628,N_3211,N_3338);
and U4629 (N_4629,N_3162,N_2570);
xor U4630 (N_4630,N_2097,N_3103);
and U4631 (N_4631,N_2623,N_3357);
or U4632 (N_4632,N_2114,N_2642);
nand U4633 (N_4633,N_3907,N_3796);
nand U4634 (N_4634,N_3764,N_3358);
or U4635 (N_4635,N_3665,N_2617);
or U4636 (N_4636,N_2274,N_2782);
xor U4637 (N_4637,N_2040,N_3795);
nor U4638 (N_4638,N_2579,N_3340);
nand U4639 (N_4639,N_3982,N_2914);
or U4640 (N_4640,N_2405,N_2708);
or U4641 (N_4641,N_2558,N_2960);
nand U4642 (N_4642,N_2884,N_3831);
or U4643 (N_4643,N_3266,N_3512);
and U4644 (N_4644,N_3917,N_3118);
and U4645 (N_4645,N_2503,N_2435);
xnor U4646 (N_4646,N_3416,N_2692);
or U4647 (N_4647,N_2233,N_2997);
and U4648 (N_4648,N_3631,N_3133);
or U4649 (N_4649,N_2571,N_3428);
and U4650 (N_4650,N_3299,N_3683);
nand U4651 (N_4651,N_3335,N_3920);
xnor U4652 (N_4652,N_3693,N_3853);
or U4653 (N_4653,N_3930,N_3497);
and U4654 (N_4654,N_2721,N_3199);
and U4655 (N_4655,N_2214,N_2735);
or U4656 (N_4656,N_3408,N_2327);
nor U4657 (N_4657,N_3004,N_3772);
xnor U4658 (N_4658,N_2662,N_3654);
and U4659 (N_4659,N_3422,N_3438);
and U4660 (N_4660,N_2120,N_2529);
nor U4661 (N_4661,N_2515,N_3607);
nand U4662 (N_4662,N_2827,N_2986);
nor U4663 (N_4663,N_3529,N_3342);
or U4664 (N_4664,N_3180,N_3521);
and U4665 (N_4665,N_3095,N_3711);
and U4666 (N_4666,N_3542,N_2801);
nand U4667 (N_4667,N_3596,N_3599);
or U4668 (N_4668,N_3146,N_3516);
nand U4669 (N_4669,N_3679,N_3559);
and U4670 (N_4670,N_2832,N_3923);
xnor U4671 (N_4671,N_2026,N_3046);
nor U4672 (N_4672,N_2582,N_2232);
and U4673 (N_4673,N_2595,N_3501);
or U4674 (N_4674,N_3669,N_2083);
nand U4675 (N_4675,N_2822,N_3323);
nand U4676 (N_4676,N_2879,N_2257);
nand U4677 (N_4677,N_2106,N_2360);
nand U4678 (N_4678,N_2354,N_2299);
or U4679 (N_4679,N_2810,N_2025);
and U4680 (N_4680,N_3963,N_2394);
or U4681 (N_4681,N_3148,N_3902);
nand U4682 (N_4682,N_3684,N_3835);
and U4683 (N_4683,N_2936,N_3515);
or U4684 (N_4684,N_3206,N_2559);
and U4685 (N_4685,N_2761,N_3889);
and U4686 (N_4686,N_2290,N_2857);
nor U4687 (N_4687,N_3592,N_3277);
nor U4688 (N_4688,N_2410,N_2700);
nand U4689 (N_4689,N_3402,N_3104);
and U4690 (N_4690,N_2380,N_3973);
nand U4691 (N_4691,N_3554,N_3653);
and U4692 (N_4692,N_2415,N_3573);
nand U4693 (N_4693,N_2568,N_3480);
and U4694 (N_4694,N_2878,N_3306);
nor U4695 (N_4695,N_3071,N_3802);
and U4696 (N_4696,N_2685,N_2020);
and U4697 (N_4697,N_3951,N_3160);
and U4698 (N_4698,N_2824,N_2666);
and U4699 (N_4699,N_3223,N_3959);
nand U4700 (N_4700,N_3622,N_3895);
nor U4701 (N_4701,N_2682,N_3577);
and U4702 (N_4702,N_2476,N_3797);
or U4703 (N_4703,N_3580,N_3226);
or U4704 (N_4704,N_2213,N_2393);
or U4705 (N_4705,N_2961,N_3019);
or U4706 (N_4706,N_2847,N_2828);
nand U4707 (N_4707,N_2626,N_3741);
and U4708 (N_4708,N_3161,N_2806);
or U4709 (N_4709,N_3355,N_3852);
nor U4710 (N_4710,N_2455,N_2248);
nand U4711 (N_4711,N_2715,N_3287);
nor U4712 (N_4712,N_3657,N_2330);
nand U4713 (N_4713,N_3361,N_2849);
nand U4714 (N_4714,N_2599,N_3642);
and U4715 (N_4715,N_3012,N_2930);
nand U4716 (N_4716,N_3883,N_2080);
or U4717 (N_4717,N_2227,N_3426);
xnor U4718 (N_4718,N_2995,N_2919);
or U4719 (N_4719,N_3454,N_3476);
and U4720 (N_4720,N_2759,N_3887);
and U4721 (N_4721,N_3939,N_3068);
and U4722 (N_4722,N_3922,N_2400);
or U4723 (N_4723,N_3049,N_2423);
nand U4724 (N_4724,N_2567,N_2787);
nor U4725 (N_4725,N_3284,N_3954);
or U4726 (N_4726,N_2923,N_3359);
or U4727 (N_4727,N_2001,N_3344);
and U4728 (N_4728,N_3195,N_3793);
nand U4729 (N_4729,N_2895,N_2105);
or U4730 (N_4730,N_3569,N_2535);
nor U4731 (N_4731,N_3615,N_2676);
nand U4732 (N_4732,N_3404,N_2140);
nand U4733 (N_4733,N_2798,N_2789);
nor U4734 (N_4734,N_2317,N_3726);
nor U4735 (N_4735,N_3827,N_2655);
or U4736 (N_4736,N_3089,N_2627);
and U4737 (N_4737,N_2601,N_3087);
and U4738 (N_4738,N_2964,N_3847);
nor U4739 (N_4739,N_3387,N_3671);
and U4740 (N_4740,N_3070,N_2110);
nor U4741 (N_4741,N_2604,N_3366);
nand U4742 (N_4742,N_3039,N_2314);
nor U4743 (N_4743,N_3268,N_3606);
nor U4744 (N_4744,N_2351,N_3251);
nand U4745 (N_4745,N_2668,N_2588);
nand U4746 (N_4746,N_3725,N_3716);
and U4747 (N_4747,N_2545,N_3663);
nand U4748 (N_4748,N_2569,N_3237);
and U4749 (N_4749,N_2517,N_2783);
nand U4750 (N_4750,N_3966,N_2427);
and U4751 (N_4751,N_2368,N_3064);
xor U4752 (N_4752,N_3566,N_2557);
nor U4753 (N_4753,N_3037,N_2815);
xor U4754 (N_4754,N_2409,N_2600);
nor U4755 (N_4755,N_3210,N_2009);
xnor U4756 (N_4756,N_2613,N_3674);
or U4757 (N_4757,N_3680,N_2339);
nand U4758 (N_4758,N_2252,N_2845);
nor U4759 (N_4759,N_3316,N_3393);
nand U4760 (N_4760,N_3771,N_2928);
nor U4761 (N_4761,N_2862,N_2984);
or U4762 (N_4762,N_2786,N_2912);
or U4763 (N_4763,N_3398,N_2471);
nor U4764 (N_4764,N_3017,N_3956);
and U4765 (N_4765,N_2794,N_2111);
and U4766 (N_4766,N_3367,N_3081);
nor U4767 (N_4767,N_2566,N_2583);
nand U4768 (N_4768,N_3890,N_2321);
nor U4769 (N_4769,N_3817,N_2293);
nor U4770 (N_4770,N_2033,N_2947);
and U4771 (N_4771,N_2576,N_2917);
or U4772 (N_4772,N_3483,N_2048);
nand U4773 (N_4773,N_2927,N_3124);
xnor U4774 (N_4774,N_3239,N_2419);
xnor U4775 (N_4775,N_2178,N_2742);
or U4776 (N_4776,N_3450,N_2461);
and U4777 (N_4777,N_2504,N_3010);
and U4778 (N_4778,N_3445,N_2967);
nor U4779 (N_4779,N_3715,N_3609);
nor U4780 (N_4780,N_2135,N_3840);
and U4781 (N_4781,N_3620,N_2699);
and U4782 (N_4782,N_2513,N_2931);
and U4783 (N_4783,N_3784,N_2514);
and U4784 (N_4784,N_2015,N_3627);
and U4785 (N_4785,N_2286,N_2399);
nand U4786 (N_4786,N_2136,N_2530);
or U4787 (N_4787,N_3311,N_3604);
nand U4788 (N_4788,N_2030,N_2622);
xnor U4789 (N_4789,N_2329,N_2690);
and U4790 (N_4790,N_3977,N_2099);
or U4791 (N_4791,N_3976,N_3808);
and U4792 (N_4792,N_3709,N_2434);
nor U4793 (N_4793,N_3914,N_3514);
xnor U4794 (N_4794,N_3301,N_2343);
nand U4795 (N_4795,N_3761,N_2084);
nand U4796 (N_4796,N_2005,N_3574);
and U4797 (N_4797,N_3303,N_2175);
or U4798 (N_4798,N_2060,N_3164);
or U4799 (N_4799,N_3862,N_3944);
nand U4800 (N_4800,N_2401,N_3186);
or U4801 (N_4801,N_3456,N_3645);
and U4802 (N_4802,N_2866,N_2952);
or U4803 (N_4803,N_2678,N_3869);
nor U4804 (N_4804,N_3464,N_2805);
and U4805 (N_4805,N_3879,N_2691);
and U4806 (N_4806,N_2864,N_2296);
nand U4807 (N_4807,N_3288,N_3194);
and U4808 (N_4808,N_2775,N_3903);
and U4809 (N_4809,N_2949,N_2267);
nor U4810 (N_4810,N_3332,N_3639);
or U4811 (N_4811,N_3475,N_3632);
and U4812 (N_4812,N_3777,N_2848);
nor U4813 (N_4813,N_2032,N_2177);
xor U4814 (N_4814,N_3768,N_2278);
or U4815 (N_4815,N_3540,N_2624);
nor U4816 (N_4816,N_2870,N_2652);
nand U4817 (N_4817,N_3126,N_2640);
and U4818 (N_4818,N_2706,N_3885);
or U4819 (N_4819,N_2432,N_3007);
nand U4820 (N_4820,N_3871,N_3467);
or U4821 (N_4821,N_3744,N_3697);
and U4822 (N_4822,N_2769,N_2875);
and U4823 (N_4823,N_3651,N_2863);
and U4824 (N_4824,N_2833,N_2978);
nor U4825 (N_4825,N_3843,N_3001);
or U4826 (N_4826,N_2609,N_3576);
and U4827 (N_4827,N_3563,N_2922);
nand U4828 (N_4828,N_2181,N_2752);
nor U4829 (N_4829,N_3543,N_3494);
xnor U4830 (N_4830,N_3493,N_2320);
nand U4831 (N_4831,N_3310,N_2871);
and U4832 (N_4832,N_2156,N_3258);
nor U4833 (N_4833,N_2496,N_2551);
and U4834 (N_4834,N_3691,N_2852);
xnor U4835 (N_4835,N_3221,N_3430);
nor U4836 (N_4836,N_3775,N_3140);
nand U4837 (N_4837,N_3397,N_2222);
nand U4838 (N_4838,N_2282,N_2704);
nand U4839 (N_4839,N_2859,N_2851);
xnor U4840 (N_4840,N_2458,N_2523);
and U4841 (N_4841,N_2159,N_3045);
nand U4842 (N_4842,N_3135,N_2955);
nand U4843 (N_4843,N_3349,N_3144);
or U4844 (N_4844,N_2562,N_2347);
or U4845 (N_4845,N_2987,N_2888);
nor U4846 (N_4846,N_2115,N_2638);
nor U4847 (N_4847,N_3246,N_2561);
or U4848 (N_4848,N_3846,N_2497);
nand U4849 (N_4849,N_3527,N_2526);
nor U4850 (N_4850,N_3952,N_3957);
or U4851 (N_4851,N_3300,N_3307);
nor U4852 (N_4852,N_2345,N_3106);
nor U4853 (N_4853,N_2677,N_3899);
nor U4854 (N_4854,N_2023,N_3935);
and U4855 (N_4855,N_2891,N_3333);
nand U4856 (N_4856,N_3921,N_3052);
and U4857 (N_4857,N_3035,N_3820);
xor U4858 (N_4858,N_3385,N_2632);
nor U4859 (N_4859,N_2754,N_3943);
and U4860 (N_4860,N_2187,N_2596);
or U4861 (N_4861,N_2639,N_3810);
nor U4862 (N_4862,N_2284,N_3628);
xor U4863 (N_4863,N_2418,N_2028);
nand U4864 (N_4864,N_2611,N_3170);
nand U4865 (N_4865,N_2417,N_3916);
xnor U4866 (N_4866,N_2921,N_2094);
xor U4867 (N_4867,N_3051,N_2516);
nor U4868 (N_4868,N_2466,N_3918);
and U4869 (N_4869,N_2019,N_2425);
or U4870 (N_4870,N_3745,N_2902);
and U4871 (N_4871,N_2439,N_2981);
nand U4872 (N_4872,N_3732,N_3291);
nor U4873 (N_4873,N_2918,N_3823);
nand U4874 (N_4874,N_2182,N_3992);
nand U4875 (N_4875,N_3410,N_2122);
or U4876 (N_4876,N_3706,N_2606);
or U4877 (N_4877,N_2016,N_2518);
or U4878 (N_4878,N_2490,N_2941);
or U4879 (N_4879,N_3466,N_3066);
nor U4880 (N_4880,N_3968,N_3508);
or U4881 (N_4881,N_3666,N_2702);
xor U4882 (N_4882,N_3153,N_3502);
and U4883 (N_4883,N_2842,N_2261);
nor U4884 (N_4884,N_2312,N_3204);
or U4885 (N_4885,N_3214,N_2454);
nand U4886 (N_4886,N_2982,N_2255);
xnor U4887 (N_4887,N_3803,N_2901);
nand U4888 (N_4888,N_3688,N_2608);
nand U4889 (N_4889,N_2037,N_2403);
nor U4890 (N_4890,N_3819,N_3462);
nand U4891 (N_4891,N_2934,N_3055);
or U4892 (N_4892,N_2877,N_3552);
nand U4893 (N_4893,N_2505,N_3893);
nor U4894 (N_4894,N_3672,N_2716);
nand U4895 (N_4895,N_2536,N_3048);
nand U4896 (N_4896,N_2219,N_3446);
or U4897 (N_4897,N_3581,N_2777);
nand U4898 (N_4898,N_2085,N_3201);
xor U4899 (N_4899,N_2834,N_3252);
nand U4900 (N_4900,N_3343,N_2153);
nand U4901 (N_4901,N_2325,N_2907);
and U4902 (N_4902,N_2287,N_2929);
and U4903 (N_4903,N_3814,N_3225);
or U4904 (N_4904,N_3575,N_2416);
and U4905 (N_4905,N_3158,N_2398);
or U4906 (N_4906,N_2915,N_3189);
and U4907 (N_4907,N_3222,N_2377);
nor U4908 (N_4908,N_2098,N_2008);
and U4909 (N_4909,N_3650,N_2241);
nand U4910 (N_4910,N_2976,N_2980);
and U4911 (N_4911,N_2074,N_3947);
and U4912 (N_4912,N_2689,N_3256);
nor U4913 (N_4913,N_3880,N_2920);
nor U4914 (N_4914,N_2088,N_3749);
nand U4915 (N_4915,N_2374,N_3662);
xor U4916 (N_4916,N_2641,N_2584);
nor U4917 (N_4917,N_3667,N_3044);
nor U4918 (N_4918,N_3067,N_3735);
nand U4919 (N_4919,N_3807,N_3370);
nor U4920 (N_4920,N_2311,N_2369);
nor U4921 (N_4921,N_3208,N_3629);
nor U4922 (N_4922,N_2811,N_3177);
and U4923 (N_4923,N_2021,N_2384);
and U4924 (N_4924,N_3746,N_3151);
xor U4925 (N_4925,N_2024,N_3278);
or U4926 (N_4926,N_2065,N_2109);
or U4927 (N_4927,N_2341,N_3519);
or U4928 (N_4928,N_3075,N_3354);
and U4929 (N_4929,N_3873,N_3376);
and U4930 (N_4930,N_3455,N_3938);
nand U4931 (N_4931,N_3014,N_2408);
nand U4932 (N_4932,N_3100,N_3090);
nand U4933 (N_4933,N_2254,N_2210);
nand U4934 (N_4934,N_2194,N_2412);
or U4935 (N_4935,N_3083,N_2031);
or U4936 (N_4936,N_2337,N_3487);
and U4937 (N_4937,N_3013,N_3635);
nor U4938 (N_4938,N_3712,N_2821);
and U4939 (N_4939,N_3616,N_3643);
nand U4940 (N_4940,N_3298,N_3626);
or U4941 (N_4941,N_2861,N_3668);
nor U4942 (N_4942,N_3056,N_3535);
xnor U4943 (N_4943,N_3757,N_3724);
nand U4944 (N_4944,N_3857,N_2292);
and U4945 (N_4945,N_2475,N_2650);
nor U4946 (N_4946,N_3780,N_3675);
or U4947 (N_4947,N_3511,N_3216);
nand U4948 (N_4948,N_3598,N_2276);
nand U4949 (N_4949,N_2904,N_3156);
nand U4950 (N_4950,N_3213,N_2800);
xor U4951 (N_4951,N_3092,N_3864);
nand U4952 (N_4952,N_2684,N_3584);
nand U4953 (N_4953,N_2240,N_2319);
nand U4954 (N_4954,N_2993,N_2778);
xnor U4955 (N_4955,N_2674,N_2963);
nor U4956 (N_4956,N_3520,N_3546);
xor U4957 (N_4957,N_2694,N_2746);
nor U4958 (N_4958,N_2357,N_3125);
nor U4959 (N_4959,N_2198,N_3489);
and U4960 (N_4960,N_2971,N_2155);
or U4961 (N_4961,N_3119,N_3468);
nor U4962 (N_4962,N_3023,N_3779);
nor U4963 (N_4963,N_3451,N_2935);
and U4964 (N_4964,N_3722,N_2838);
xnor U4965 (N_4965,N_2605,N_2492);
or U4966 (N_4966,N_3484,N_3593);
and U4967 (N_4967,N_3995,N_2004);
or U4968 (N_4968,N_2043,N_2531);
nor U4969 (N_4969,N_3321,N_2411);
xor U4970 (N_4970,N_3016,N_2038);
nor U4971 (N_4971,N_2067,N_3969);
nand U4972 (N_4972,N_2628,N_3499);
or U4973 (N_4973,N_3350,N_3750);
or U4974 (N_4974,N_3572,N_2124);
nand U4975 (N_4975,N_3330,N_2146);
nor U4976 (N_4976,N_2082,N_2910);
or U4977 (N_4977,N_3324,N_2302);
or U4978 (N_4978,N_2924,N_3859);
nand U4979 (N_4979,N_3038,N_2258);
xnor U4980 (N_4980,N_2992,N_3528);
nand U4981 (N_4981,N_2791,N_3507);
or U4982 (N_4982,N_2107,N_2736);
or U4983 (N_4983,N_2365,N_3553);
or U4984 (N_4984,N_3060,N_3202);
and U4985 (N_4985,N_2473,N_3533);
nand U4986 (N_4986,N_2081,N_2633);
nand U4987 (N_4987,N_3754,N_3696);
and U4988 (N_4988,N_2117,N_3364);
and U4989 (N_4989,N_2957,N_2830);
nor U4990 (N_4990,N_3782,N_2134);
nor U4991 (N_4991,N_3228,N_2793);
or U4992 (N_4992,N_2017,N_3791);
or U4993 (N_4993,N_2719,N_2154);
nor U4994 (N_4994,N_2646,N_2239);
nor U4995 (N_4995,N_2837,N_3337);
nor U4996 (N_4996,N_2795,N_3981);
nand U4997 (N_4997,N_2391,N_2840);
nand U4998 (N_4998,N_3702,N_3555);
nor U4999 (N_4999,N_3617,N_2051);
and U5000 (N_5000,N_2925,N_2286);
and U5001 (N_5001,N_2703,N_3674);
nor U5002 (N_5002,N_3444,N_3976);
or U5003 (N_5003,N_3471,N_3025);
nand U5004 (N_5004,N_3756,N_3813);
nand U5005 (N_5005,N_2983,N_3406);
nor U5006 (N_5006,N_3742,N_2176);
nand U5007 (N_5007,N_2310,N_3154);
nand U5008 (N_5008,N_3996,N_2981);
and U5009 (N_5009,N_2670,N_3159);
or U5010 (N_5010,N_3230,N_3271);
xnor U5011 (N_5011,N_3608,N_3549);
xor U5012 (N_5012,N_2926,N_3834);
nand U5013 (N_5013,N_2013,N_3746);
nor U5014 (N_5014,N_2874,N_2370);
and U5015 (N_5015,N_2217,N_2193);
and U5016 (N_5016,N_3107,N_3553);
or U5017 (N_5017,N_2863,N_3413);
nor U5018 (N_5018,N_2467,N_3408);
nand U5019 (N_5019,N_3245,N_3462);
and U5020 (N_5020,N_2115,N_3115);
nor U5021 (N_5021,N_3768,N_3622);
or U5022 (N_5022,N_2157,N_2884);
nor U5023 (N_5023,N_3523,N_3369);
and U5024 (N_5024,N_3872,N_3915);
or U5025 (N_5025,N_3206,N_3489);
and U5026 (N_5026,N_3079,N_2647);
or U5027 (N_5027,N_2690,N_3299);
or U5028 (N_5028,N_3496,N_2182);
and U5029 (N_5029,N_2986,N_2581);
or U5030 (N_5030,N_3672,N_2112);
and U5031 (N_5031,N_3452,N_3102);
nand U5032 (N_5032,N_2185,N_2329);
nor U5033 (N_5033,N_2656,N_2961);
or U5034 (N_5034,N_2407,N_3469);
and U5035 (N_5035,N_3994,N_2726);
xor U5036 (N_5036,N_3581,N_3944);
and U5037 (N_5037,N_3385,N_2694);
nor U5038 (N_5038,N_2878,N_3401);
nand U5039 (N_5039,N_2204,N_3345);
or U5040 (N_5040,N_3254,N_2264);
nand U5041 (N_5041,N_2409,N_3086);
nor U5042 (N_5042,N_3863,N_2752);
and U5043 (N_5043,N_3436,N_3634);
or U5044 (N_5044,N_3741,N_2427);
nand U5045 (N_5045,N_2013,N_3059);
nand U5046 (N_5046,N_3250,N_2955);
and U5047 (N_5047,N_2912,N_2247);
and U5048 (N_5048,N_3545,N_2965);
and U5049 (N_5049,N_3940,N_2534);
and U5050 (N_5050,N_2167,N_2475);
and U5051 (N_5051,N_3184,N_2374);
and U5052 (N_5052,N_2880,N_2881);
nor U5053 (N_5053,N_3569,N_3720);
and U5054 (N_5054,N_2141,N_3236);
nand U5055 (N_5055,N_3838,N_3441);
or U5056 (N_5056,N_2141,N_3597);
or U5057 (N_5057,N_3461,N_3553);
nor U5058 (N_5058,N_3315,N_2299);
nor U5059 (N_5059,N_2681,N_2332);
nor U5060 (N_5060,N_2605,N_2450);
or U5061 (N_5061,N_2408,N_2890);
or U5062 (N_5062,N_3830,N_3278);
or U5063 (N_5063,N_3109,N_3549);
nor U5064 (N_5064,N_3929,N_2742);
and U5065 (N_5065,N_2266,N_2566);
nor U5066 (N_5066,N_3372,N_3903);
nand U5067 (N_5067,N_3865,N_3414);
or U5068 (N_5068,N_3331,N_2040);
nand U5069 (N_5069,N_3862,N_3410);
and U5070 (N_5070,N_2489,N_2452);
and U5071 (N_5071,N_2357,N_3422);
nand U5072 (N_5072,N_3444,N_3046);
or U5073 (N_5073,N_2269,N_2036);
or U5074 (N_5074,N_2420,N_3537);
nand U5075 (N_5075,N_3604,N_3836);
or U5076 (N_5076,N_3608,N_2775);
or U5077 (N_5077,N_2814,N_3969);
or U5078 (N_5078,N_3397,N_2359);
nand U5079 (N_5079,N_2990,N_3159);
nand U5080 (N_5080,N_2175,N_3051);
or U5081 (N_5081,N_2550,N_3095);
nand U5082 (N_5082,N_3051,N_3017);
nor U5083 (N_5083,N_3534,N_2031);
nor U5084 (N_5084,N_3609,N_2137);
or U5085 (N_5085,N_2604,N_2714);
nand U5086 (N_5086,N_2902,N_2237);
or U5087 (N_5087,N_2244,N_3638);
and U5088 (N_5088,N_3724,N_3490);
nand U5089 (N_5089,N_3278,N_3893);
xnor U5090 (N_5090,N_3118,N_2422);
nor U5091 (N_5091,N_3562,N_3341);
nand U5092 (N_5092,N_2171,N_3865);
nor U5093 (N_5093,N_2936,N_3747);
xor U5094 (N_5094,N_3092,N_2260);
xnor U5095 (N_5095,N_3937,N_2572);
nor U5096 (N_5096,N_3060,N_3598);
nor U5097 (N_5097,N_3284,N_3153);
or U5098 (N_5098,N_3194,N_2132);
or U5099 (N_5099,N_2755,N_3973);
and U5100 (N_5100,N_3789,N_2237);
xor U5101 (N_5101,N_3425,N_3688);
and U5102 (N_5102,N_3008,N_2148);
nor U5103 (N_5103,N_2388,N_2106);
nand U5104 (N_5104,N_2218,N_3800);
nor U5105 (N_5105,N_2133,N_2710);
and U5106 (N_5106,N_2213,N_2214);
and U5107 (N_5107,N_2965,N_3475);
or U5108 (N_5108,N_3938,N_3180);
nor U5109 (N_5109,N_2309,N_3829);
xor U5110 (N_5110,N_2424,N_2104);
xor U5111 (N_5111,N_3272,N_2358);
nor U5112 (N_5112,N_3550,N_3623);
xnor U5113 (N_5113,N_3469,N_2059);
or U5114 (N_5114,N_3096,N_2268);
nor U5115 (N_5115,N_2004,N_2497);
or U5116 (N_5116,N_2951,N_3549);
nor U5117 (N_5117,N_2638,N_2711);
nand U5118 (N_5118,N_3281,N_2814);
nand U5119 (N_5119,N_3163,N_2774);
xnor U5120 (N_5120,N_2068,N_3665);
and U5121 (N_5121,N_2472,N_3142);
or U5122 (N_5122,N_2855,N_3539);
nor U5123 (N_5123,N_3513,N_2598);
nand U5124 (N_5124,N_3461,N_3993);
nor U5125 (N_5125,N_3380,N_2407);
or U5126 (N_5126,N_3505,N_3796);
nor U5127 (N_5127,N_2477,N_3176);
or U5128 (N_5128,N_2063,N_3855);
xor U5129 (N_5129,N_2793,N_3325);
nand U5130 (N_5130,N_3610,N_2644);
nor U5131 (N_5131,N_3697,N_2211);
nand U5132 (N_5132,N_2538,N_2419);
nor U5133 (N_5133,N_2480,N_3269);
or U5134 (N_5134,N_2887,N_2776);
or U5135 (N_5135,N_2047,N_3409);
and U5136 (N_5136,N_3982,N_2838);
nor U5137 (N_5137,N_3047,N_3942);
xnor U5138 (N_5138,N_3312,N_3453);
and U5139 (N_5139,N_2900,N_2223);
and U5140 (N_5140,N_3826,N_3284);
nand U5141 (N_5141,N_2858,N_3895);
nor U5142 (N_5142,N_2717,N_3001);
nand U5143 (N_5143,N_3196,N_2271);
nor U5144 (N_5144,N_2373,N_3415);
nand U5145 (N_5145,N_3706,N_2294);
nor U5146 (N_5146,N_2683,N_2609);
nor U5147 (N_5147,N_2989,N_2625);
and U5148 (N_5148,N_2633,N_2935);
xor U5149 (N_5149,N_3908,N_3938);
and U5150 (N_5150,N_3210,N_3921);
and U5151 (N_5151,N_2658,N_2204);
or U5152 (N_5152,N_2903,N_3979);
nand U5153 (N_5153,N_2547,N_3685);
nor U5154 (N_5154,N_2577,N_2163);
nand U5155 (N_5155,N_3986,N_3474);
and U5156 (N_5156,N_2505,N_2803);
nor U5157 (N_5157,N_2456,N_2644);
and U5158 (N_5158,N_2480,N_3047);
or U5159 (N_5159,N_2641,N_2016);
nand U5160 (N_5160,N_2569,N_2026);
or U5161 (N_5161,N_3847,N_2744);
or U5162 (N_5162,N_2416,N_3103);
xor U5163 (N_5163,N_3480,N_3755);
nand U5164 (N_5164,N_3602,N_2546);
xor U5165 (N_5165,N_2658,N_2103);
and U5166 (N_5166,N_2162,N_2900);
xor U5167 (N_5167,N_3194,N_3325);
xnor U5168 (N_5168,N_2394,N_3287);
nand U5169 (N_5169,N_2109,N_3532);
and U5170 (N_5170,N_2193,N_3525);
nor U5171 (N_5171,N_2822,N_3259);
nand U5172 (N_5172,N_3803,N_3607);
xnor U5173 (N_5173,N_2417,N_2836);
nand U5174 (N_5174,N_3867,N_3497);
and U5175 (N_5175,N_3558,N_2815);
and U5176 (N_5176,N_2356,N_2603);
nand U5177 (N_5177,N_3207,N_2125);
nor U5178 (N_5178,N_3162,N_3284);
or U5179 (N_5179,N_2390,N_3672);
nand U5180 (N_5180,N_3755,N_3465);
or U5181 (N_5181,N_3433,N_3878);
nand U5182 (N_5182,N_3573,N_3300);
and U5183 (N_5183,N_2410,N_3873);
xnor U5184 (N_5184,N_2747,N_2321);
nor U5185 (N_5185,N_3088,N_3259);
nor U5186 (N_5186,N_3865,N_3514);
nor U5187 (N_5187,N_2154,N_3864);
nand U5188 (N_5188,N_2430,N_2403);
xnor U5189 (N_5189,N_2770,N_3008);
nor U5190 (N_5190,N_3188,N_3850);
nor U5191 (N_5191,N_3511,N_2050);
and U5192 (N_5192,N_2121,N_2045);
xor U5193 (N_5193,N_3840,N_3388);
nand U5194 (N_5194,N_2269,N_3666);
nand U5195 (N_5195,N_2455,N_3287);
nand U5196 (N_5196,N_3689,N_2194);
nand U5197 (N_5197,N_3397,N_2367);
or U5198 (N_5198,N_3775,N_2853);
nor U5199 (N_5199,N_2322,N_2299);
or U5200 (N_5200,N_3452,N_3004);
and U5201 (N_5201,N_3668,N_2634);
nand U5202 (N_5202,N_2750,N_2534);
or U5203 (N_5203,N_2836,N_3567);
nand U5204 (N_5204,N_2766,N_2739);
nor U5205 (N_5205,N_3803,N_3859);
or U5206 (N_5206,N_3711,N_3829);
or U5207 (N_5207,N_2947,N_3015);
nor U5208 (N_5208,N_3053,N_3375);
nand U5209 (N_5209,N_3356,N_3124);
or U5210 (N_5210,N_3002,N_3134);
and U5211 (N_5211,N_2658,N_2028);
nor U5212 (N_5212,N_3605,N_2003);
and U5213 (N_5213,N_3903,N_2082);
nor U5214 (N_5214,N_3070,N_3838);
and U5215 (N_5215,N_2119,N_3655);
nor U5216 (N_5216,N_3751,N_3251);
or U5217 (N_5217,N_2574,N_2564);
nand U5218 (N_5218,N_3046,N_3669);
or U5219 (N_5219,N_2824,N_2402);
nand U5220 (N_5220,N_2617,N_2209);
and U5221 (N_5221,N_2335,N_2942);
and U5222 (N_5222,N_3804,N_2239);
xnor U5223 (N_5223,N_2529,N_2083);
nor U5224 (N_5224,N_3142,N_2760);
nand U5225 (N_5225,N_3904,N_3462);
and U5226 (N_5226,N_3818,N_2016);
and U5227 (N_5227,N_3525,N_2827);
or U5228 (N_5228,N_3014,N_2657);
or U5229 (N_5229,N_2593,N_3821);
and U5230 (N_5230,N_2213,N_3934);
or U5231 (N_5231,N_3393,N_3288);
nor U5232 (N_5232,N_3462,N_2702);
or U5233 (N_5233,N_3192,N_2140);
or U5234 (N_5234,N_3637,N_3383);
nand U5235 (N_5235,N_2448,N_2792);
or U5236 (N_5236,N_3076,N_2824);
xnor U5237 (N_5237,N_3135,N_2317);
nand U5238 (N_5238,N_2396,N_3462);
nor U5239 (N_5239,N_2095,N_2857);
nand U5240 (N_5240,N_2213,N_3788);
nand U5241 (N_5241,N_3147,N_2543);
xnor U5242 (N_5242,N_2727,N_3910);
or U5243 (N_5243,N_3427,N_3656);
or U5244 (N_5244,N_2035,N_2307);
nor U5245 (N_5245,N_2003,N_2085);
or U5246 (N_5246,N_3597,N_2382);
nand U5247 (N_5247,N_3785,N_2223);
or U5248 (N_5248,N_3399,N_2659);
or U5249 (N_5249,N_2027,N_2994);
and U5250 (N_5250,N_2207,N_3534);
nand U5251 (N_5251,N_3186,N_2513);
or U5252 (N_5252,N_3493,N_3027);
or U5253 (N_5253,N_2634,N_2652);
or U5254 (N_5254,N_2711,N_2328);
and U5255 (N_5255,N_2061,N_2773);
xor U5256 (N_5256,N_3122,N_2597);
nor U5257 (N_5257,N_2333,N_2370);
or U5258 (N_5258,N_3827,N_3418);
and U5259 (N_5259,N_3351,N_3087);
or U5260 (N_5260,N_3373,N_3621);
or U5261 (N_5261,N_3215,N_2178);
nor U5262 (N_5262,N_2274,N_3383);
xnor U5263 (N_5263,N_2431,N_2855);
xor U5264 (N_5264,N_2358,N_2574);
or U5265 (N_5265,N_3701,N_2662);
xnor U5266 (N_5266,N_2175,N_3518);
and U5267 (N_5267,N_3043,N_2760);
nor U5268 (N_5268,N_3332,N_2659);
nor U5269 (N_5269,N_3592,N_2514);
nand U5270 (N_5270,N_3963,N_2904);
nor U5271 (N_5271,N_2390,N_2430);
nor U5272 (N_5272,N_2907,N_3505);
or U5273 (N_5273,N_2494,N_3464);
nand U5274 (N_5274,N_3302,N_2749);
nor U5275 (N_5275,N_3283,N_3264);
or U5276 (N_5276,N_3426,N_2639);
or U5277 (N_5277,N_3709,N_3898);
xor U5278 (N_5278,N_3756,N_2097);
nand U5279 (N_5279,N_2061,N_3703);
nor U5280 (N_5280,N_3606,N_3027);
nand U5281 (N_5281,N_3782,N_2232);
nand U5282 (N_5282,N_2096,N_3409);
and U5283 (N_5283,N_3640,N_3841);
nand U5284 (N_5284,N_2716,N_2663);
or U5285 (N_5285,N_2969,N_3056);
nand U5286 (N_5286,N_2291,N_3490);
and U5287 (N_5287,N_2240,N_2443);
nand U5288 (N_5288,N_3510,N_2439);
nand U5289 (N_5289,N_2530,N_3002);
or U5290 (N_5290,N_2691,N_2367);
nor U5291 (N_5291,N_2743,N_2530);
and U5292 (N_5292,N_2158,N_2660);
or U5293 (N_5293,N_3245,N_3206);
nand U5294 (N_5294,N_2907,N_3579);
nor U5295 (N_5295,N_2669,N_3796);
nand U5296 (N_5296,N_2053,N_3706);
nand U5297 (N_5297,N_3465,N_2416);
nand U5298 (N_5298,N_3376,N_2836);
nor U5299 (N_5299,N_2484,N_2224);
or U5300 (N_5300,N_3105,N_3457);
nand U5301 (N_5301,N_3882,N_2426);
and U5302 (N_5302,N_3693,N_3117);
or U5303 (N_5303,N_3729,N_3201);
and U5304 (N_5304,N_2269,N_2535);
nand U5305 (N_5305,N_3677,N_2073);
or U5306 (N_5306,N_3448,N_2266);
or U5307 (N_5307,N_2621,N_3335);
and U5308 (N_5308,N_2026,N_3234);
and U5309 (N_5309,N_3608,N_2810);
or U5310 (N_5310,N_2132,N_2251);
or U5311 (N_5311,N_3800,N_3895);
and U5312 (N_5312,N_3048,N_3231);
nor U5313 (N_5313,N_2049,N_2233);
and U5314 (N_5314,N_3485,N_3142);
nand U5315 (N_5315,N_2875,N_3606);
xnor U5316 (N_5316,N_3694,N_2361);
and U5317 (N_5317,N_3517,N_3514);
xor U5318 (N_5318,N_3175,N_2523);
and U5319 (N_5319,N_3234,N_2131);
nor U5320 (N_5320,N_2470,N_3766);
or U5321 (N_5321,N_2107,N_3865);
nand U5322 (N_5322,N_2709,N_2510);
nor U5323 (N_5323,N_2568,N_3220);
nand U5324 (N_5324,N_2592,N_2745);
and U5325 (N_5325,N_3151,N_2821);
xnor U5326 (N_5326,N_3819,N_2203);
or U5327 (N_5327,N_3684,N_2404);
nand U5328 (N_5328,N_3135,N_2972);
xor U5329 (N_5329,N_2418,N_3631);
nand U5330 (N_5330,N_3953,N_2767);
and U5331 (N_5331,N_3038,N_2126);
nand U5332 (N_5332,N_2162,N_2847);
or U5333 (N_5333,N_3644,N_2574);
or U5334 (N_5334,N_3605,N_3635);
nor U5335 (N_5335,N_3076,N_3878);
nand U5336 (N_5336,N_3350,N_2549);
nor U5337 (N_5337,N_2151,N_3251);
nand U5338 (N_5338,N_2043,N_2964);
and U5339 (N_5339,N_2747,N_3916);
nand U5340 (N_5340,N_3129,N_2516);
and U5341 (N_5341,N_3063,N_2938);
or U5342 (N_5342,N_2880,N_2497);
nand U5343 (N_5343,N_2077,N_3767);
nand U5344 (N_5344,N_3314,N_3072);
nand U5345 (N_5345,N_2484,N_3506);
nand U5346 (N_5346,N_3568,N_2149);
and U5347 (N_5347,N_3533,N_2650);
nand U5348 (N_5348,N_2013,N_3392);
nand U5349 (N_5349,N_2794,N_3320);
xnor U5350 (N_5350,N_2045,N_2631);
nand U5351 (N_5351,N_3538,N_2071);
or U5352 (N_5352,N_3087,N_3078);
and U5353 (N_5353,N_2276,N_2570);
or U5354 (N_5354,N_3649,N_3958);
nand U5355 (N_5355,N_3836,N_3854);
and U5356 (N_5356,N_2250,N_3421);
nand U5357 (N_5357,N_2501,N_3312);
nor U5358 (N_5358,N_3002,N_3225);
or U5359 (N_5359,N_3915,N_2610);
nand U5360 (N_5360,N_3680,N_3264);
or U5361 (N_5361,N_3652,N_3913);
nor U5362 (N_5362,N_2811,N_2001);
xor U5363 (N_5363,N_3257,N_3456);
and U5364 (N_5364,N_3322,N_2773);
xnor U5365 (N_5365,N_3762,N_3711);
or U5366 (N_5366,N_3595,N_2715);
or U5367 (N_5367,N_2057,N_2952);
and U5368 (N_5368,N_3839,N_3885);
or U5369 (N_5369,N_2053,N_3204);
and U5370 (N_5370,N_2934,N_3531);
nor U5371 (N_5371,N_3409,N_3824);
or U5372 (N_5372,N_2608,N_3268);
nor U5373 (N_5373,N_3111,N_3482);
and U5374 (N_5374,N_2350,N_2155);
and U5375 (N_5375,N_2598,N_2784);
xnor U5376 (N_5376,N_3019,N_2875);
or U5377 (N_5377,N_3034,N_2854);
nand U5378 (N_5378,N_3865,N_2999);
nand U5379 (N_5379,N_3116,N_2861);
xnor U5380 (N_5380,N_3024,N_3905);
nor U5381 (N_5381,N_3704,N_2380);
and U5382 (N_5382,N_2000,N_2972);
nand U5383 (N_5383,N_2984,N_3753);
nor U5384 (N_5384,N_3955,N_2457);
nor U5385 (N_5385,N_3669,N_3517);
or U5386 (N_5386,N_3609,N_3062);
nor U5387 (N_5387,N_3726,N_2800);
nand U5388 (N_5388,N_3418,N_2356);
xnor U5389 (N_5389,N_3418,N_2513);
and U5390 (N_5390,N_3661,N_3920);
nor U5391 (N_5391,N_3421,N_2150);
and U5392 (N_5392,N_3013,N_2786);
nand U5393 (N_5393,N_3009,N_2167);
or U5394 (N_5394,N_3960,N_2813);
nor U5395 (N_5395,N_3230,N_2528);
nand U5396 (N_5396,N_3143,N_2485);
nand U5397 (N_5397,N_2698,N_2003);
nand U5398 (N_5398,N_2341,N_3064);
or U5399 (N_5399,N_2731,N_2476);
and U5400 (N_5400,N_3810,N_3264);
nand U5401 (N_5401,N_2162,N_3597);
and U5402 (N_5402,N_2884,N_3583);
and U5403 (N_5403,N_2562,N_2357);
xnor U5404 (N_5404,N_3687,N_2470);
xor U5405 (N_5405,N_3217,N_3596);
and U5406 (N_5406,N_3522,N_3740);
xnor U5407 (N_5407,N_2120,N_3014);
nand U5408 (N_5408,N_2772,N_2192);
nand U5409 (N_5409,N_3197,N_2351);
or U5410 (N_5410,N_3169,N_2997);
nand U5411 (N_5411,N_2257,N_3641);
or U5412 (N_5412,N_3989,N_3417);
or U5413 (N_5413,N_2865,N_3630);
and U5414 (N_5414,N_2731,N_3811);
or U5415 (N_5415,N_3106,N_2525);
nand U5416 (N_5416,N_3519,N_2531);
nand U5417 (N_5417,N_3866,N_3037);
and U5418 (N_5418,N_3370,N_2991);
nand U5419 (N_5419,N_3352,N_2492);
nor U5420 (N_5420,N_2820,N_3925);
or U5421 (N_5421,N_2721,N_3282);
xor U5422 (N_5422,N_2889,N_2012);
xor U5423 (N_5423,N_3601,N_3803);
and U5424 (N_5424,N_3101,N_3267);
nand U5425 (N_5425,N_2751,N_2681);
nand U5426 (N_5426,N_2887,N_2293);
or U5427 (N_5427,N_3828,N_3218);
and U5428 (N_5428,N_2660,N_2827);
or U5429 (N_5429,N_2770,N_2606);
or U5430 (N_5430,N_2844,N_2094);
nor U5431 (N_5431,N_3919,N_3538);
and U5432 (N_5432,N_3055,N_3449);
or U5433 (N_5433,N_2238,N_3121);
nor U5434 (N_5434,N_2449,N_3576);
or U5435 (N_5435,N_3349,N_3637);
or U5436 (N_5436,N_3734,N_2219);
and U5437 (N_5437,N_2602,N_2355);
nor U5438 (N_5438,N_2630,N_3866);
nor U5439 (N_5439,N_3789,N_3815);
or U5440 (N_5440,N_2021,N_3685);
nor U5441 (N_5441,N_2501,N_2829);
or U5442 (N_5442,N_3751,N_2536);
or U5443 (N_5443,N_3306,N_2894);
nor U5444 (N_5444,N_2295,N_3259);
or U5445 (N_5445,N_2410,N_3508);
and U5446 (N_5446,N_3565,N_3907);
or U5447 (N_5447,N_2572,N_2696);
nand U5448 (N_5448,N_2945,N_2900);
nor U5449 (N_5449,N_2168,N_2744);
nand U5450 (N_5450,N_3226,N_3324);
or U5451 (N_5451,N_2134,N_2743);
and U5452 (N_5452,N_2976,N_2578);
or U5453 (N_5453,N_3524,N_3160);
or U5454 (N_5454,N_2690,N_2583);
or U5455 (N_5455,N_2778,N_2415);
nor U5456 (N_5456,N_2732,N_3364);
nand U5457 (N_5457,N_2932,N_2485);
nand U5458 (N_5458,N_3277,N_2646);
nor U5459 (N_5459,N_2229,N_2258);
or U5460 (N_5460,N_3585,N_2767);
and U5461 (N_5461,N_3884,N_3585);
and U5462 (N_5462,N_3284,N_3986);
nand U5463 (N_5463,N_2551,N_2896);
and U5464 (N_5464,N_3427,N_2233);
nor U5465 (N_5465,N_3579,N_2270);
nor U5466 (N_5466,N_3198,N_3528);
or U5467 (N_5467,N_2573,N_2260);
or U5468 (N_5468,N_2393,N_2066);
or U5469 (N_5469,N_2874,N_3859);
and U5470 (N_5470,N_2689,N_2912);
xnor U5471 (N_5471,N_3985,N_3493);
or U5472 (N_5472,N_3356,N_2254);
and U5473 (N_5473,N_2331,N_2442);
or U5474 (N_5474,N_2038,N_2139);
nand U5475 (N_5475,N_3369,N_2363);
nand U5476 (N_5476,N_2207,N_3203);
nor U5477 (N_5477,N_2406,N_3968);
and U5478 (N_5478,N_2520,N_2956);
nand U5479 (N_5479,N_2169,N_2370);
and U5480 (N_5480,N_3349,N_2952);
and U5481 (N_5481,N_2804,N_2659);
or U5482 (N_5482,N_3970,N_2559);
nand U5483 (N_5483,N_3354,N_2191);
and U5484 (N_5484,N_3681,N_2102);
nand U5485 (N_5485,N_2889,N_3333);
xnor U5486 (N_5486,N_2383,N_3639);
and U5487 (N_5487,N_2027,N_2741);
nand U5488 (N_5488,N_2641,N_2155);
and U5489 (N_5489,N_2382,N_3118);
nor U5490 (N_5490,N_3908,N_2131);
xnor U5491 (N_5491,N_3077,N_2323);
nor U5492 (N_5492,N_2877,N_2117);
nand U5493 (N_5493,N_2069,N_3369);
nand U5494 (N_5494,N_2286,N_3531);
xor U5495 (N_5495,N_2121,N_3920);
nand U5496 (N_5496,N_2287,N_2504);
and U5497 (N_5497,N_3317,N_3577);
nand U5498 (N_5498,N_2620,N_2627);
or U5499 (N_5499,N_2813,N_3782);
or U5500 (N_5500,N_3383,N_2695);
and U5501 (N_5501,N_3212,N_2593);
or U5502 (N_5502,N_2343,N_3051);
nand U5503 (N_5503,N_3013,N_2465);
or U5504 (N_5504,N_3764,N_2962);
or U5505 (N_5505,N_3571,N_3380);
and U5506 (N_5506,N_2184,N_3597);
nand U5507 (N_5507,N_3627,N_2874);
and U5508 (N_5508,N_2557,N_3842);
or U5509 (N_5509,N_3065,N_3462);
nor U5510 (N_5510,N_2879,N_3829);
or U5511 (N_5511,N_3044,N_2130);
and U5512 (N_5512,N_2731,N_2145);
nor U5513 (N_5513,N_3032,N_2314);
nor U5514 (N_5514,N_3167,N_2563);
and U5515 (N_5515,N_3047,N_3173);
and U5516 (N_5516,N_3559,N_3430);
nand U5517 (N_5517,N_3488,N_2799);
and U5518 (N_5518,N_2174,N_2930);
xnor U5519 (N_5519,N_2958,N_3664);
nand U5520 (N_5520,N_3290,N_2516);
or U5521 (N_5521,N_3452,N_2371);
or U5522 (N_5522,N_2650,N_2358);
xnor U5523 (N_5523,N_2470,N_2815);
and U5524 (N_5524,N_2295,N_2824);
nand U5525 (N_5525,N_3954,N_3363);
and U5526 (N_5526,N_3126,N_3244);
or U5527 (N_5527,N_2586,N_2541);
and U5528 (N_5528,N_3071,N_3767);
nand U5529 (N_5529,N_2542,N_3045);
and U5530 (N_5530,N_3455,N_2408);
nand U5531 (N_5531,N_2417,N_2644);
nor U5532 (N_5532,N_3377,N_3083);
nand U5533 (N_5533,N_2145,N_3903);
nor U5534 (N_5534,N_2492,N_3248);
nand U5535 (N_5535,N_3636,N_2050);
nor U5536 (N_5536,N_2704,N_3117);
nor U5537 (N_5537,N_3335,N_2829);
nor U5538 (N_5538,N_2998,N_3247);
nor U5539 (N_5539,N_2809,N_2022);
nand U5540 (N_5540,N_2905,N_2899);
or U5541 (N_5541,N_2599,N_2256);
xnor U5542 (N_5542,N_3514,N_2724);
xnor U5543 (N_5543,N_3738,N_3055);
nor U5544 (N_5544,N_2508,N_2230);
and U5545 (N_5545,N_2257,N_3980);
nand U5546 (N_5546,N_2922,N_3795);
and U5547 (N_5547,N_2107,N_2246);
nand U5548 (N_5548,N_3983,N_2470);
and U5549 (N_5549,N_3689,N_3215);
nor U5550 (N_5550,N_2016,N_2860);
nor U5551 (N_5551,N_2210,N_2349);
or U5552 (N_5552,N_2726,N_2530);
and U5553 (N_5553,N_3789,N_2655);
or U5554 (N_5554,N_3941,N_3017);
and U5555 (N_5555,N_2708,N_3526);
nor U5556 (N_5556,N_3550,N_2448);
nand U5557 (N_5557,N_2650,N_2230);
xor U5558 (N_5558,N_2969,N_2380);
nor U5559 (N_5559,N_3796,N_2731);
or U5560 (N_5560,N_3623,N_3692);
nor U5561 (N_5561,N_2062,N_3109);
and U5562 (N_5562,N_2721,N_3946);
nand U5563 (N_5563,N_3520,N_2506);
and U5564 (N_5564,N_2488,N_2848);
or U5565 (N_5565,N_3517,N_3276);
nand U5566 (N_5566,N_2467,N_3235);
and U5567 (N_5567,N_2443,N_2011);
nor U5568 (N_5568,N_2586,N_2097);
nand U5569 (N_5569,N_3794,N_3759);
and U5570 (N_5570,N_2590,N_3790);
xnor U5571 (N_5571,N_2028,N_2381);
nand U5572 (N_5572,N_3556,N_2704);
nand U5573 (N_5573,N_3205,N_2390);
and U5574 (N_5574,N_2059,N_3404);
xor U5575 (N_5575,N_3723,N_3597);
or U5576 (N_5576,N_2275,N_2288);
and U5577 (N_5577,N_3572,N_3371);
and U5578 (N_5578,N_3952,N_3336);
and U5579 (N_5579,N_2202,N_3007);
nand U5580 (N_5580,N_3223,N_3325);
or U5581 (N_5581,N_2977,N_3371);
or U5582 (N_5582,N_2318,N_2591);
nor U5583 (N_5583,N_2489,N_2184);
or U5584 (N_5584,N_2897,N_3957);
xor U5585 (N_5585,N_2399,N_3477);
or U5586 (N_5586,N_2240,N_2948);
nand U5587 (N_5587,N_3235,N_3432);
xor U5588 (N_5588,N_2105,N_3338);
nor U5589 (N_5589,N_3688,N_3906);
nand U5590 (N_5590,N_3608,N_2225);
nor U5591 (N_5591,N_2033,N_3053);
nor U5592 (N_5592,N_3325,N_3730);
and U5593 (N_5593,N_2224,N_3323);
nor U5594 (N_5594,N_3897,N_3971);
or U5595 (N_5595,N_2932,N_3810);
nand U5596 (N_5596,N_2109,N_2717);
and U5597 (N_5597,N_2548,N_3542);
xor U5598 (N_5598,N_3989,N_3802);
or U5599 (N_5599,N_2327,N_3798);
nor U5600 (N_5600,N_3269,N_2881);
nand U5601 (N_5601,N_3222,N_3365);
nor U5602 (N_5602,N_3245,N_2859);
or U5603 (N_5603,N_3208,N_3011);
and U5604 (N_5604,N_3947,N_2114);
and U5605 (N_5605,N_3325,N_2557);
nor U5606 (N_5606,N_3278,N_3854);
nor U5607 (N_5607,N_3552,N_3988);
or U5608 (N_5608,N_2536,N_2876);
and U5609 (N_5609,N_3936,N_2099);
nor U5610 (N_5610,N_3853,N_2036);
and U5611 (N_5611,N_3928,N_3741);
nand U5612 (N_5612,N_2282,N_3099);
nand U5613 (N_5613,N_3713,N_3475);
and U5614 (N_5614,N_2075,N_2221);
nor U5615 (N_5615,N_2209,N_2508);
or U5616 (N_5616,N_2317,N_3504);
and U5617 (N_5617,N_3128,N_2412);
nor U5618 (N_5618,N_2647,N_2889);
or U5619 (N_5619,N_2129,N_2448);
xnor U5620 (N_5620,N_2190,N_3523);
nand U5621 (N_5621,N_2623,N_2981);
or U5622 (N_5622,N_3595,N_3097);
nand U5623 (N_5623,N_3299,N_3642);
and U5624 (N_5624,N_2451,N_3112);
nor U5625 (N_5625,N_2356,N_3602);
nand U5626 (N_5626,N_2015,N_3193);
and U5627 (N_5627,N_2613,N_3632);
or U5628 (N_5628,N_2971,N_3878);
nand U5629 (N_5629,N_2944,N_2891);
and U5630 (N_5630,N_2407,N_3472);
or U5631 (N_5631,N_2068,N_3498);
nor U5632 (N_5632,N_2797,N_3837);
nor U5633 (N_5633,N_3191,N_2316);
xnor U5634 (N_5634,N_3230,N_3833);
nand U5635 (N_5635,N_3589,N_3117);
nand U5636 (N_5636,N_2382,N_3679);
nor U5637 (N_5637,N_3277,N_2231);
nor U5638 (N_5638,N_3345,N_2962);
and U5639 (N_5639,N_2846,N_2562);
nor U5640 (N_5640,N_2105,N_3168);
and U5641 (N_5641,N_2816,N_2285);
nor U5642 (N_5642,N_2901,N_2844);
xor U5643 (N_5643,N_3424,N_3694);
nand U5644 (N_5644,N_2344,N_2432);
nand U5645 (N_5645,N_2532,N_2328);
or U5646 (N_5646,N_2290,N_2883);
and U5647 (N_5647,N_3452,N_3616);
nor U5648 (N_5648,N_3684,N_2151);
or U5649 (N_5649,N_2523,N_2435);
nand U5650 (N_5650,N_2231,N_2682);
and U5651 (N_5651,N_2647,N_2991);
or U5652 (N_5652,N_3916,N_2388);
and U5653 (N_5653,N_3197,N_2136);
and U5654 (N_5654,N_3742,N_2697);
and U5655 (N_5655,N_2415,N_2117);
nand U5656 (N_5656,N_3005,N_2936);
xor U5657 (N_5657,N_3770,N_3160);
or U5658 (N_5658,N_2424,N_3862);
nand U5659 (N_5659,N_3217,N_3688);
nand U5660 (N_5660,N_2192,N_2277);
and U5661 (N_5661,N_2480,N_3201);
or U5662 (N_5662,N_2940,N_2797);
or U5663 (N_5663,N_3405,N_3119);
or U5664 (N_5664,N_3040,N_3848);
xor U5665 (N_5665,N_2170,N_3451);
nand U5666 (N_5666,N_3928,N_3152);
nand U5667 (N_5667,N_2659,N_2724);
nand U5668 (N_5668,N_3188,N_3663);
nor U5669 (N_5669,N_2578,N_2187);
and U5670 (N_5670,N_3215,N_3611);
xor U5671 (N_5671,N_3078,N_3007);
or U5672 (N_5672,N_2915,N_3116);
or U5673 (N_5673,N_2305,N_2265);
and U5674 (N_5674,N_3022,N_2031);
and U5675 (N_5675,N_3045,N_3800);
or U5676 (N_5676,N_2539,N_3913);
nand U5677 (N_5677,N_3490,N_3168);
or U5678 (N_5678,N_2474,N_2372);
nand U5679 (N_5679,N_2368,N_3392);
or U5680 (N_5680,N_3950,N_2168);
nand U5681 (N_5681,N_2791,N_3660);
and U5682 (N_5682,N_3406,N_2876);
nand U5683 (N_5683,N_2327,N_3659);
and U5684 (N_5684,N_3693,N_3619);
nor U5685 (N_5685,N_2447,N_3631);
nor U5686 (N_5686,N_3441,N_2900);
nor U5687 (N_5687,N_2849,N_2816);
and U5688 (N_5688,N_2580,N_2932);
or U5689 (N_5689,N_2734,N_3613);
xor U5690 (N_5690,N_3203,N_2758);
and U5691 (N_5691,N_3797,N_3451);
xnor U5692 (N_5692,N_3137,N_2638);
or U5693 (N_5693,N_2519,N_3860);
or U5694 (N_5694,N_2069,N_3113);
or U5695 (N_5695,N_3577,N_2222);
nand U5696 (N_5696,N_3593,N_3001);
and U5697 (N_5697,N_3910,N_2549);
nand U5698 (N_5698,N_2444,N_2338);
or U5699 (N_5699,N_3582,N_2353);
and U5700 (N_5700,N_2246,N_3327);
and U5701 (N_5701,N_2355,N_2109);
nand U5702 (N_5702,N_2405,N_3434);
xnor U5703 (N_5703,N_3578,N_2753);
and U5704 (N_5704,N_2565,N_2980);
or U5705 (N_5705,N_2609,N_2074);
xor U5706 (N_5706,N_2364,N_3252);
nor U5707 (N_5707,N_2908,N_2017);
or U5708 (N_5708,N_2788,N_3953);
or U5709 (N_5709,N_2467,N_2684);
nor U5710 (N_5710,N_3297,N_3622);
nand U5711 (N_5711,N_2807,N_2585);
and U5712 (N_5712,N_3047,N_2703);
xor U5713 (N_5713,N_3564,N_3111);
xor U5714 (N_5714,N_3420,N_2832);
nor U5715 (N_5715,N_2943,N_2859);
nand U5716 (N_5716,N_3775,N_2996);
and U5717 (N_5717,N_2129,N_2185);
and U5718 (N_5718,N_2755,N_2233);
nand U5719 (N_5719,N_3441,N_2724);
xnor U5720 (N_5720,N_3862,N_3807);
nor U5721 (N_5721,N_2090,N_3249);
nand U5722 (N_5722,N_2862,N_2414);
or U5723 (N_5723,N_3221,N_2366);
and U5724 (N_5724,N_3068,N_2620);
nand U5725 (N_5725,N_3171,N_3847);
or U5726 (N_5726,N_3358,N_2704);
nand U5727 (N_5727,N_3522,N_2554);
and U5728 (N_5728,N_3715,N_3499);
and U5729 (N_5729,N_3416,N_2444);
and U5730 (N_5730,N_2649,N_3498);
nor U5731 (N_5731,N_2215,N_3356);
nand U5732 (N_5732,N_2684,N_3365);
nor U5733 (N_5733,N_3837,N_2555);
and U5734 (N_5734,N_3785,N_3362);
or U5735 (N_5735,N_2557,N_2390);
nor U5736 (N_5736,N_3427,N_3257);
and U5737 (N_5737,N_3823,N_3762);
xnor U5738 (N_5738,N_3624,N_3745);
or U5739 (N_5739,N_3069,N_3230);
xor U5740 (N_5740,N_3034,N_3938);
and U5741 (N_5741,N_3438,N_2162);
nand U5742 (N_5742,N_2436,N_2581);
nand U5743 (N_5743,N_2191,N_2818);
xor U5744 (N_5744,N_3918,N_2131);
nand U5745 (N_5745,N_2933,N_2590);
xnor U5746 (N_5746,N_3259,N_2402);
nor U5747 (N_5747,N_2815,N_3855);
and U5748 (N_5748,N_3644,N_3306);
nand U5749 (N_5749,N_2421,N_3467);
xnor U5750 (N_5750,N_2123,N_3729);
and U5751 (N_5751,N_2596,N_2045);
nand U5752 (N_5752,N_2963,N_2706);
or U5753 (N_5753,N_2868,N_3616);
and U5754 (N_5754,N_3741,N_2683);
nor U5755 (N_5755,N_3743,N_3165);
xnor U5756 (N_5756,N_3482,N_3902);
nor U5757 (N_5757,N_3680,N_3948);
nor U5758 (N_5758,N_2082,N_2631);
nor U5759 (N_5759,N_3313,N_3780);
nand U5760 (N_5760,N_3608,N_2148);
nand U5761 (N_5761,N_2564,N_3844);
nor U5762 (N_5762,N_3741,N_2605);
xor U5763 (N_5763,N_3675,N_3295);
nor U5764 (N_5764,N_3799,N_3214);
nand U5765 (N_5765,N_2064,N_2633);
and U5766 (N_5766,N_3798,N_3597);
or U5767 (N_5767,N_3964,N_2545);
or U5768 (N_5768,N_2489,N_3843);
nand U5769 (N_5769,N_2062,N_3537);
nand U5770 (N_5770,N_3912,N_2782);
nand U5771 (N_5771,N_2418,N_2006);
nand U5772 (N_5772,N_2581,N_2386);
nor U5773 (N_5773,N_3299,N_3397);
and U5774 (N_5774,N_3259,N_2855);
xor U5775 (N_5775,N_2978,N_3217);
and U5776 (N_5776,N_2715,N_3164);
nand U5777 (N_5777,N_2209,N_3711);
and U5778 (N_5778,N_2637,N_3410);
nand U5779 (N_5779,N_2214,N_2343);
or U5780 (N_5780,N_2315,N_3928);
nand U5781 (N_5781,N_3864,N_3102);
and U5782 (N_5782,N_2172,N_2091);
nor U5783 (N_5783,N_2716,N_2197);
nand U5784 (N_5784,N_3708,N_3302);
nand U5785 (N_5785,N_2517,N_2569);
nand U5786 (N_5786,N_2818,N_2795);
and U5787 (N_5787,N_2228,N_2102);
nand U5788 (N_5788,N_2702,N_3754);
nand U5789 (N_5789,N_2077,N_3337);
nor U5790 (N_5790,N_3757,N_3540);
and U5791 (N_5791,N_2361,N_3121);
or U5792 (N_5792,N_2043,N_3161);
nand U5793 (N_5793,N_2780,N_2806);
nand U5794 (N_5794,N_3149,N_3416);
nor U5795 (N_5795,N_2279,N_3324);
nor U5796 (N_5796,N_3189,N_2511);
nand U5797 (N_5797,N_3940,N_2570);
nand U5798 (N_5798,N_3497,N_3317);
and U5799 (N_5799,N_2810,N_3214);
or U5800 (N_5800,N_2851,N_3604);
and U5801 (N_5801,N_3589,N_2824);
and U5802 (N_5802,N_3117,N_2033);
nor U5803 (N_5803,N_3158,N_2380);
nor U5804 (N_5804,N_3705,N_2764);
nand U5805 (N_5805,N_2207,N_2352);
or U5806 (N_5806,N_3618,N_3540);
nor U5807 (N_5807,N_3198,N_3492);
or U5808 (N_5808,N_2102,N_2173);
nand U5809 (N_5809,N_2720,N_2109);
and U5810 (N_5810,N_3970,N_3524);
nand U5811 (N_5811,N_3000,N_3284);
or U5812 (N_5812,N_3334,N_2310);
nor U5813 (N_5813,N_3663,N_2807);
xnor U5814 (N_5814,N_2228,N_2093);
or U5815 (N_5815,N_3425,N_3263);
nor U5816 (N_5816,N_2783,N_2059);
nor U5817 (N_5817,N_2676,N_2613);
or U5818 (N_5818,N_3380,N_2168);
and U5819 (N_5819,N_2581,N_2891);
and U5820 (N_5820,N_3123,N_2203);
nand U5821 (N_5821,N_2309,N_3210);
and U5822 (N_5822,N_2403,N_3472);
or U5823 (N_5823,N_3110,N_2627);
nor U5824 (N_5824,N_3150,N_2542);
nand U5825 (N_5825,N_2524,N_2665);
xnor U5826 (N_5826,N_3840,N_2377);
nand U5827 (N_5827,N_2831,N_2781);
nor U5828 (N_5828,N_2030,N_2669);
nand U5829 (N_5829,N_3825,N_3202);
nor U5830 (N_5830,N_2874,N_3008);
nor U5831 (N_5831,N_2259,N_2513);
xnor U5832 (N_5832,N_2107,N_3789);
and U5833 (N_5833,N_2342,N_3943);
nand U5834 (N_5834,N_3446,N_2017);
or U5835 (N_5835,N_3582,N_3952);
and U5836 (N_5836,N_3130,N_3009);
or U5837 (N_5837,N_3846,N_2104);
nand U5838 (N_5838,N_3477,N_3862);
nor U5839 (N_5839,N_2247,N_3542);
nor U5840 (N_5840,N_3097,N_3651);
nor U5841 (N_5841,N_2416,N_2258);
or U5842 (N_5842,N_2106,N_2594);
nand U5843 (N_5843,N_2690,N_2615);
xnor U5844 (N_5844,N_2368,N_3469);
or U5845 (N_5845,N_2747,N_2659);
xor U5846 (N_5846,N_3174,N_3727);
nand U5847 (N_5847,N_2105,N_3701);
xnor U5848 (N_5848,N_3453,N_2460);
and U5849 (N_5849,N_3917,N_3804);
and U5850 (N_5850,N_2079,N_2927);
or U5851 (N_5851,N_3383,N_3704);
nor U5852 (N_5852,N_2812,N_2269);
or U5853 (N_5853,N_3683,N_3641);
nor U5854 (N_5854,N_2838,N_2882);
nor U5855 (N_5855,N_3058,N_3401);
and U5856 (N_5856,N_3761,N_3720);
nor U5857 (N_5857,N_3087,N_3601);
or U5858 (N_5858,N_3581,N_3687);
and U5859 (N_5859,N_3477,N_3698);
nand U5860 (N_5860,N_3220,N_3931);
and U5861 (N_5861,N_2612,N_3303);
or U5862 (N_5862,N_3733,N_2361);
nand U5863 (N_5863,N_2797,N_3666);
nor U5864 (N_5864,N_3811,N_2159);
nor U5865 (N_5865,N_2138,N_2186);
nor U5866 (N_5866,N_3621,N_3764);
xnor U5867 (N_5867,N_3377,N_3983);
nor U5868 (N_5868,N_3913,N_2047);
or U5869 (N_5869,N_3228,N_2150);
or U5870 (N_5870,N_3189,N_2723);
xnor U5871 (N_5871,N_3353,N_2254);
nand U5872 (N_5872,N_2218,N_2970);
xnor U5873 (N_5873,N_3341,N_2421);
or U5874 (N_5874,N_3209,N_3354);
nand U5875 (N_5875,N_3739,N_3233);
and U5876 (N_5876,N_2290,N_3807);
nor U5877 (N_5877,N_3247,N_2380);
nor U5878 (N_5878,N_2803,N_2610);
or U5879 (N_5879,N_2793,N_3896);
or U5880 (N_5880,N_3971,N_2802);
xnor U5881 (N_5881,N_3179,N_2551);
nor U5882 (N_5882,N_3820,N_3569);
nor U5883 (N_5883,N_2604,N_3101);
xor U5884 (N_5884,N_2309,N_2360);
nand U5885 (N_5885,N_3559,N_2529);
nand U5886 (N_5886,N_3768,N_2867);
nand U5887 (N_5887,N_3761,N_3827);
nand U5888 (N_5888,N_3247,N_2033);
or U5889 (N_5889,N_2759,N_3540);
and U5890 (N_5890,N_2820,N_2031);
nor U5891 (N_5891,N_3629,N_3891);
nor U5892 (N_5892,N_3610,N_3596);
nor U5893 (N_5893,N_3341,N_3381);
xor U5894 (N_5894,N_3932,N_3786);
or U5895 (N_5895,N_2612,N_2722);
nor U5896 (N_5896,N_2200,N_3954);
nand U5897 (N_5897,N_2154,N_3978);
or U5898 (N_5898,N_3660,N_2729);
nand U5899 (N_5899,N_2300,N_3257);
nor U5900 (N_5900,N_3575,N_3988);
or U5901 (N_5901,N_2360,N_2706);
nand U5902 (N_5902,N_3813,N_3177);
or U5903 (N_5903,N_3891,N_2732);
nor U5904 (N_5904,N_3887,N_2772);
and U5905 (N_5905,N_3071,N_2552);
nand U5906 (N_5906,N_3347,N_2624);
and U5907 (N_5907,N_2005,N_2332);
nand U5908 (N_5908,N_3669,N_3643);
nor U5909 (N_5909,N_2588,N_3959);
and U5910 (N_5910,N_3790,N_2602);
and U5911 (N_5911,N_3246,N_3079);
xor U5912 (N_5912,N_2730,N_2166);
nor U5913 (N_5913,N_3149,N_2743);
nand U5914 (N_5914,N_2556,N_2992);
or U5915 (N_5915,N_2243,N_2000);
and U5916 (N_5916,N_3728,N_2694);
or U5917 (N_5917,N_2549,N_2855);
nand U5918 (N_5918,N_2757,N_3057);
nand U5919 (N_5919,N_3310,N_2431);
or U5920 (N_5920,N_2954,N_2487);
nor U5921 (N_5921,N_2774,N_2981);
nor U5922 (N_5922,N_3770,N_3395);
or U5923 (N_5923,N_2818,N_3256);
xnor U5924 (N_5924,N_3920,N_2241);
or U5925 (N_5925,N_2117,N_3412);
or U5926 (N_5926,N_2313,N_2923);
nor U5927 (N_5927,N_2666,N_2013);
nor U5928 (N_5928,N_3333,N_3466);
nor U5929 (N_5929,N_2235,N_2722);
nand U5930 (N_5930,N_3326,N_3453);
nand U5931 (N_5931,N_3243,N_3826);
nand U5932 (N_5932,N_3924,N_3983);
nand U5933 (N_5933,N_3018,N_2285);
nand U5934 (N_5934,N_2053,N_2701);
nand U5935 (N_5935,N_2380,N_2466);
and U5936 (N_5936,N_2927,N_3408);
nor U5937 (N_5937,N_2216,N_2075);
or U5938 (N_5938,N_3570,N_2678);
nand U5939 (N_5939,N_3012,N_3090);
nand U5940 (N_5940,N_2957,N_2090);
and U5941 (N_5941,N_2994,N_2655);
nor U5942 (N_5942,N_3421,N_2727);
xnor U5943 (N_5943,N_2512,N_3097);
nand U5944 (N_5944,N_2517,N_2628);
nor U5945 (N_5945,N_2313,N_3188);
or U5946 (N_5946,N_3080,N_3007);
and U5947 (N_5947,N_2419,N_3735);
nand U5948 (N_5948,N_2191,N_2438);
or U5949 (N_5949,N_2956,N_2257);
and U5950 (N_5950,N_3254,N_3419);
nand U5951 (N_5951,N_3816,N_2878);
or U5952 (N_5952,N_2137,N_2239);
or U5953 (N_5953,N_3912,N_3023);
or U5954 (N_5954,N_3626,N_2916);
nor U5955 (N_5955,N_3533,N_2392);
nand U5956 (N_5956,N_2030,N_3564);
nand U5957 (N_5957,N_3104,N_3494);
nor U5958 (N_5958,N_3832,N_2256);
nor U5959 (N_5959,N_2146,N_3028);
nand U5960 (N_5960,N_3369,N_2330);
nor U5961 (N_5961,N_2965,N_3996);
or U5962 (N_5962,N_3003,N_2578);
nand U5963 (N_5963,N_2563,N_2736);
or U5964 (N_5964,N_2905,N_2749);
and U5965 (N_5965,N_2310,N_3523);
and U5966 (N_5966,N_2795,N_3529);
and U5967 (N_5967,N_2484,N_2072);
nor U5968 (N_5968,N_2956,N_3033);
nor U5969 (N_5969,N_2082,N_2250);
nor U5970 (N_5970,N_2629,N_2203);
nand U5971 (N_5971,N_3774,N_3441);
nor U5972 (N_5972,N_3028,N_2904);
xor U5973 (N_5973,N_2374,N_2323);
nor U5974 (N_5974,N_3485,N_2442);
or U5975 (N_5975,N_2575,N_2130);
or U5976 (N_5976,N_2112,N_2067);
nor U5977 (N_5977,N_2880,N_2562);
or U5978 (N_5978,N_3835,N_2511);
or U5979 (N_5979,N_3346,N_3074);
and U5980 (N_5980,N_2386,N_3713);
or U5981 (N_5981,N_2698,N_3223);
nor U5982 (N_5982,N_3019,N_3310);
and U5983 (N_5983,N_3746,N_3214);
nand U5984 (N_5984,N_2289,N_3023);
nand U5985 (N_5985,N_2715,N_3604);
nor U5986 (N_5986,N_2771,N_2973);
nor U5987 (N_5987,N_3458,N_2358);
nand U5988 (N_5988,N_2611,N_2116);
or U5989 (N_5989,N_3262,N_3850);
nor U5990 (N_5990,N_2386,N_2348);
or U5991 (N_5991,N_3193,N_3607);
nand U5992 (N_5992,N_3453,N_2466);
and U5993 (N_5993,N_3315,N_2708);
nand U5994 (N_5994,N_2071,N_2790);
nand U5995 (N_5995,N_2367,N_3108);
nor U5996 (N_5996,N_3348,N_3941);
and U5997 (N_5997,N_3627,N_3336);
nor U5998 (N_5998,N_3627,N_3654);
nand U5999 (N_5999,N_2203,N_3071);
nand U6000 (N_6000,N_4423,N_4330);
or U6001 (N_6001,N_5477,N_4616);
or U6002 (N_6002,N_4180,N_5404);
or U6003 (N_6003,N_5671,N_4794);
nand U6004 (N_6004,N_5606,N_4850);
and U6005 (N_6005,N_5323,N_4245);
xor U6006 (N_6006,N_5994,N_4457);
nand U6007 (N_6007,N_5416,N_4196);
and U6008 (N_6008,N_4576,N_5469);
and U6009 (N_6009,N_5553,N_5640);
nand U6010 (N_6010,N_4523,N_5661);
and U6011 (N_6011,N_5570,N_4627);
nand U6012 (N_6012,N_4951,N_4485);
and U6013 (N_6013,N_4450,N_5543);
and U6014 (N_6014,N_5051,N_4977);
and U6015 (N_6015,N_5159,N_5451);
and U6016 (N_6016,N_4884,N_5331);
xnor U6017 (N_6017,N_5118,N_4528);
xnor U6018 (N_6018,N_4014,N_4691);
nor U6019 (N_6019,N_4418,N_5363);
or U6020 (N_6020,N_5252,N_5151);
nor U6021 (N_6021,N_4518,N_4172);
nand U6022 (N_6022,N_5349,N_5835);
or U6023 (N_6023,N_4359,N_5559);
nor U6024 (N_6024,N_5911,N_4391);
nand U6025 (N_6025,N_4157,N_5940);
xnor U6026 (N_6026,N_5737,N_5968);
nor U6027 (N_6027,N_5235,N_4901);
and U6028 (N_6028,N_5315,N_4260);
nor U6029 (N_6029,N_5286,N_4818);
nor U6030 (N_6030,N_5985,N_5170);
nor U6031 (N_6031,N_5875,N_5577);
or U6032 (N_6032,N_4823,N_5024);
or U6033 (N_6033,N_4659,N_5430);
or U6034 (N_6034,N_4987,N_4481);
or U6035 (N_6035,N_5609,N_4278);
and U6036 (N_6036,N_5942,N_4280);
nand U6037 (N_6037,N_5683,N_4836);
nor U6038 (N_6038,N_4687,N_4342);
nand U6039 (N_6039,N_4962,N_4397);
and U6040 (N_6040,N_4055,N_4847);
or U6041 (N_6041,N_4117,N_5798);
or U6042 (N_6042,N_5055,N_5335);
or U6043 (N_6043,N_5990,N_4864);
nand U6044 (N_6044,N_5371,N_5541);
nor U6045 (N_6045,N_4362,N_5145);
and U6046 (N_6046,N_4570,N_4804);
nand U6047 (N_6047,N_5042,N_4377);
nand U6048 (N_6048,N_5470,N_5545);
nor U6049 (N_6049,N_4022,N_5540);
nand U6050 (N_6050,N_4185,N_4547);
nor U6051 (N_6051,N_4767,N_5103);
nand U6052 (N_6052,N_4730,N_4270);
and U6053 (N_6053,N_4437,N_4536);
or U6054 (N_6054,N_4876,N_5439);
nor U6055 (N_6055,N_4016,N_4365);
and U6056 (N_6056,N_5478,N_4151);
nor U6057 (N_6057,N_4086,N_4512);
nand U6058 (N_6058,N_5225,N_4279);
and U6059 (N_6059,N_5520,N_4060);
xor U6060 (N_6060,N_5638,N_5092);
nor U6061 (N_6061,N_5895,N_5319);
nand U6062 (N_6062,N_4604,N_4769);
or U6063 (N_6063,N_4338,N_4503);
and U6064 (N_6064,N_4040,N_5720);
nand U6065 (N_6065,N_4634,N_5361);
or U6066 (N_6066,N_4803,N_4126);
or U6067 (N_6067,N_4162,N_4506);
and U6068 (N_6068,N_4104,N_4881);
nor U6069 (N_6069,N_4853,N_5232);
xor U6070 (N_6070,N_4668,N_4100);
nand U6071 (N_6071,N_5122,N_4985);
nor U6072 (N_6072,N_5125,N_5724);
nand U6073 (N_6073,N_5256,N_5022);
or U6074 (N_6074,N_4200,N_4098);
nand U6075 (N_6075,N_4110,N_4556);
nor U6076 (N_6076,N_4852,N_5355);
nand U6077 (N_6077,N_4171,N_5096);
nand U6078 (N_6078,N_4937,N_5458);
nand U6079 (N_6079,N_5805,N_4198);
nand U6080 (N_6080,N_5104,N_4143);
nand U6081 (N_6081,N_5819,N_4800);
xor U6082 (N_6082,N_5273,N_4140);
nand U6083 (N_6083,N_5695,N_4802);
or U6084 (N_6084,N_4586,N_5049);
or U6085 (N_6085,N_5936,N_5729);
or U6086 (N_6086,N_5975,N_4891);
or U6087 (N_6087,N_4456,N_4814);
nor U6088 (N_6088,N_5573,N_5890);
or U6089 (N_6089,N_5785,N_5846);
or U6090 (N_6090,N_4129,N_5676);
and U6091 (N_6091,N_5728,N_4675);
nand U6092 (N_6092,N_4801,N_4241);
or U6093 (N_6093,N_5955,N_5743);
nor U6094 (N_6094,N_5768,N_4111);
or U6095 (N_6095,N_4896,N_4910);
nand U6096 (N_6096,N_4941,N_5996);
or U6097 (N_6097,N_5792,N_4553);
nor U6098 (N_6098,N_4061,N_5219);
and U6099 (N_6099,N_4477,N_4979);
and U6100 (N_6100,N_4192,N_4045);
and U6101 (N_6101,N_5901,N_5906);
nor U6102 (N_6102,N_4123,N_5584);
nand U6103 (N_6103,N_5382,N_4137);
nor U6104 (N_6104,N_4489,N_4453);
nand U6105 (N_6105,N_5263,N_4064);
nand U6106 (N_6106,N_4302,N_4862);
or U6107 (N_6107,N_4644,N_4158);
and U6108 (N_6108,N_4778,N_4461);
and U6109 (N_6109,N_4618,N_4821);
and U6110 (N_6110,N_5217,N_4974);
xor U6111 (N_6111,N_4035,N_4703);
or U6112 (N_6112,N_5864,N_5922);
or U6113 (N_6113,N_4851,N_4772);
nand U6114 (N_6114,N_4933,N_5953);
and U6115 (N_6115,N_5820,N_5855);
nand U6116 (N_6116,N_5860,N_4337);
nand U6117 (N_6117,N_4204,N_5401);
nor U6118 (N_6118,N_4809,N_5612);
xnor U6119 (N_6119,N_4078,N_5195);
or U6120 (N_6120,N_4677,N_4463);
nand U6121 (N_6121,N_4465,N_4640);
or U6122 (N_6122,N_4652,N_5255);
or U6123 (N_6123,N_5998,N_5426);
nand U6124 (N_6124,N_5644,N_4381);
or U6125 (N_6125,N_4114,N_5949);
and U6126 (N_6126,N_4115,N_5044);
or U6127 (N_6127,N_5457,N_4471);
or U6128 (N_6128,N_4839,N_4826);
or U6129 (N_6129,N_4213,N_4698);
nor U6130 (N_6130,N_4212,N_4321);
nor U6131 (N_6131,N_4354,N_4969);
or U6132 (N_6132,N_5354,N_5460);
and U6133 (N_6133,N_4967,N_4355);
or U6134 (N_6134,N_5133,N_5882);
or U6135 (N_6135,N_4048,N_4754);
nor U6136 (N_6136,N_5394,N_5427);
or U6137 (N_6137,N_5658,N_5324);
or U6138 (N_6138,N_5506,N_5398);
or U6139 (N_6139,N_5504,N_4034);
nor U6140 (N_6140,N_5947,N_5221);
and U6141 (N_6141,N_4382,N_5074);
nor U6142 (N_6142,N_5838,N_4076);
and U6143 (N_6143,N_4141,N_4540);
or U6144 (N_6144,N_5699,N_4953);
nand U6145 (N_6145,N_5310,N_4727);
nand U6146 (N_6146,N_4568,N_5672);
and U6147 (N_6147,N_4358,N_5365);
nand U6148 (N_6148,N_5777,N_4792);
nor U6149 (N_6149,N_4218,N_5435);
nand U6150 (N_6150,N_5102,N_4316);
and U6151 (N_6151,N_5065,N_4870);
or U6152 (N_6152,N_5405,N_5475);
nand U6153 (N_6153,N_5894,N_4925);
and U6154 (N_6154,N_4963,N_4983);
nand U6155 (N_6155,N_4118,N_4039);
nor U6156 (N_6156,N_5280,N_4025);
nor U6157 (N_6157,N_4297,N_5076);
nor U6158 (N_6158,N_4075,N_4537);
nor U6159 (N_6159,N_4089,N_5727);
xnor U6160 (N_6160,N_5706,N_5375);
nand U6161 (N_6161,N_5993,N_5836);
and U6162 (N_6162,N_5862,N_4590);
or U6163 (N_6163,N_4704,N_5031);
nor U6164 (N_6164,N_5641,N_5312);
or U6165 (N_6165,N_5876,N_4255);
xnor U6166 (N_6166,N_4748,N_4053);
nor U6167 (N_6167,N_5939,N_4403);
and U6168 (N_6168,N_5978,N_5476);
and U6169 (N_6169,N_5781,N_4808);
and U6170 (N_6170,N_5230,N_5653);
and U6171 (N_6171,N_4948,N_5824);
nand U6172 (N_6172,N_4900,N_4722);
nor U6173 (N_6173,N_5141,N_5878);
and U6174 (N_6174,N_4920,N_5826);
nand U6175 (N_6175,N_5418,N_4219);
and U6176 (N_6176,N_5220,N_4102);
nor U6177 (N_6177,N_4183,N_4885);
nand U6178 (N_6178,N_4613,N_5995);
xnor U6179 (N_6179,N_5611,N_4246);
or U6180 (N_6180,N_4810,N_5941);
nand U6181 (N_6181,N_4784,N_4432);
xor U6182 (N_6182,N_5169,N_4124);
nand U6183 (N_6183,N_4319,N_5078);
or U6184 (N_6184,N_5081,N_5150);
or U6185 (N_6185,N_5370,N_5030);
nand U6186 (N_6186,N_5907,N_5926);
or U6187 (N_6187,N_4517,N_4526);
nor U6188 (N_6188,N_5224,N_5707);
and U6189 (N_6189,N_5203,N_4532);
nor U6190 (N_6190,N_4079,N_4719);
or U6191 (N_6191,N_5585,N_4125);
nand U6192 (N_6192,N_5385,N_5816);
nand U6193 (N_6193,N_5011,N_4220);
or U6194 (N_6194,N_4426,N_4234);
and U6195 (N_6195,N_5966,N_5174);
nor U6196 (N_6196,N_4238,N_4154);
or U6197 (N_6197,N_5311,N_4904);
nand U6198 (N_6198,N_4139,N_4658);
or U6199 (N_6199,N_5285,N_4231);
or U6200 (N_6200,N_4837,N_5209);
or U6201 (N_6201,N_4431,N_5309);
nand U6202 (N_6202,N_5378,N_5459);
xor U6203 (N_6203,N_4167,N_5193);
nand U6204 (N_6204,N_4736,N_5094);
and U6205 (N_6205,N_4499,N_4692);
nor U6206 (N_6206,N_4133,N_4895);
and U6207 (N_6207,N_4622,N_4914);
and U6208 (N_6208,N_4475,N_5511);
and U6209 (N_6209,N_4844,N_5373);
nand U6210 (N_6210,N_4134,N_4024);
or U6211 (N_6211,N_4458,N_4420);
nor U6212 (N_6212,N_5246,N_5796);
or U6213 (N_6213,N_5608,N_5015);
nand U6214 (N_6214,N_5025,N_4472);
or U6215 (N_6215,N_5344,N_4610);
or U6216 (N_6216,N_5002,N_4843);
or U6217 (N_6217,N_4262,N_4112);
or U6218 (N_6218,N_5666,N_4487);
nand U6219 (N_6219,N_4715,N_5379);
and U6220 (N_6220,N_5198,N_5554);
nor U6221 (N_6221,N_5077,N_5701);
or U6222 (N_6222,N_4166,N_4070);
xnor U6223 (N_6223,N_5062,N_5071);
nand U6224 (N_6224,N_5467,N_4682);
or U6225 (N_6225,N_5774,N_4944);
or U6226 (N_6226,N_4938,N_5549);
nand U6227 (N_6227,N_4392,N_5556);
nor U6228 (N_6228,N_5969,N_4052);
and U6229 (N_6229,N_5710,N_4495);
or U6230 (N_6230,N_5881,N_5402);
and U6231 (N_6231,N_4266,N_4000);
xnor U6232 (N_6232,N_5054,N_5564);
nand U6233 (N_6233,N_5960,N_5928);
and U6234 (N_6234,N_4380,N_4776);
nor U6235 (N_6235,N_4689,N_5132);
xor U6236 (N_6236,N_5973,N_4854);
and U6237 (N_6237,N_4492,N_5212);
or U6238 (N_6238,N_5991,N_5497);
and U6239 (N_6239,N_4164,N_5207);
nand U6240 (N_6240,N_4903,N_4099);
and U6241 (N_6241,N_4029,N_4747);
and U6242 (N_6242,N_5977,N_4653);
xor U6243 (N_6243,N_5865,N_5537);
nor U6244 (N_6244,N_5615,N_5682);
xnor U6245 (N_6245,N_5892,N_5493);
nor U6246 (N_6246,N_5395,N_4289);
and U6247 (N_6247,N_4227,N_4444);
nor U6248 (N_6248,N_5183,N_4286);
or U6249 (N_6249,N_5294,N_4191);
nor U6250 (N_6250,N_4994,N_5592);
nand U6251 (N_6251,N_4701,N_5204);
nor U6252 (N_6252,N_5026,N_4861);
and U6253 (N_6253,N_4197,N_4455);
and U6254 (N_6254,N_5099,N_4964);
nor U6255 (N_6255,N_5698,N_5665);
or U6256 (N_6256,N_5643,N_5519);
or U6257 (N_6257,N_5880,N_5586);
or U6258 (N_6258,N_5013,N_5580);
or U6259 (N_6259,N_5072,N_5572);
nand U6260 (N_6260,N_5804,N_4441);
nor U6261 (N_6261,N_4871,N_4324);
nor U6262 (N_6262,N_4688,N_5069);
or U6263 (N_6263,N_5299,N_5524);
nor U6264 (N_6264,N_4301,N_5129);
xnor U6265 (N_6265,N_5296,N_5776);
nor U6266 (N_6266,N_4071,N_4975);
nand U6267 (N_6267,N_4257,N_5061);
and U6268 (N_6268,N_5390,N_4954);
nor U6269 (N_6269,N_5738,N_5893);
or U6270 (N_6270,N_5045,N_5934);
and U6271 (N_6271,N_5625,N_5561);
nand U6272 (N_6272,N_5060,N_4188);
and U6273 (N_6273,N_4161,N_5173);
and U6274 (N_6274,N_4389,N_4978);
nor U6275 (N_6275,N_4294,N_4244);
nor U6276 (N_6276,N_5347,N_5075);
nor U6277 (N_6277,N_4522,N_5464);
nand U6278 (N_6278,N_4731,N_5269);
and U6279 (N_6279,N_4581,N_4527);
nand U6280 (N_6280,N_4044,N_4094);
xnor U6281 (N_6281,N_4287,N_5412);
nand U6282 (N_6282,N_5645,N_4429);
and U6283 (N_6283,N_5593,N_4081);
nand U6284 (N_6284,N_5920,N_5956);
and U6285 (N_6285,N_5253,N_4177);
nor U6286 (N_6286,N_4685,N_4515);
and U6287 (N_6287,N_5250,N_4085);
nor U6288 (N_6288,N_4404,N_4273);
nand U6289 (N_6289,N_4519,N_5532);
nor U6290 (N_6290,N_4214,N_4763);
and U6291 (N_6291,N_4699,N_4790);
and U6292 (N_6292,N_4860,N_5184);
nand U6293 (N_6293,N_5921,N_4863);
nor U6294 (N_6294,N_4057,N_5276);
and U6295 (N_6295,N_5360,N_5756);
or U6296 (N_6296,N_5156,N_5518);
or U6297 (N_6297,N_4375,N_5338);
xnor U6298 (N_6298,N_5583,N_4811);
nand U6299 (N_6299,N_4786,N_5352);
or U6300 (N_6300,N_4897,N_4628);
nand U6301 (N_6301,N_5258,N_5109);
nand U6302 (N_6302,N_5610,N_4232);
and U6303 (N_6303,N_4142,N_5105);
nand U6304 (N_6304,N_4927,N_4921);
nor U6305 (N_6305,N_4765,N_5691);
and U6306 (N_6306,N_4379,N_5199);
nand U6307 (N_6307,N_5297,N_4690);
nor U6308 (N_6308,N_4488,N_5807);
nand U6309 (N_6309,N_5770,N_4935);
or U6310 (N_6310,N_4563,N_4146);
nand U6311 (N_6311,N_5873,N_4080);
and U6312 (N_6312,N_4483,N_5775);
and U6313 (N_6313,N_4229,N_4728);
or U6314 (N_6314,N_4693,N_5162);
nor U6315 (N_6315,N_4221,N_4973);
or U6316 (N_6316,N_4956,N_4406);
and U6317 (N_6317,N_5433,N_5456);
or U6318 (N_6318,N_5264,N_4686);
nor U6319 (N_6319,N_5766,N_5627);
nor U6320 (N_6320,N_5763,N_5449);
and U6321 (N_6321,N_4199,N_5755);
or U6322 (N_6322,N_4817,N_5190);
or U6323 (N_6323,N_4939,N_4734);
nand U6324 (N_6324,N_4740,N_5827);
and U6325 (N_6325,N_5282,N_4395);
nor U6326 (N_6326,N_4646,N_5779);
nor U6327 (N_6327,N_5542,N_4737);
xor U6328 (N_6328,N_4660,N_5483);
or U6329 (N_6329,N_5924,N_4293);
and U6330 (N_6330,N_5853,N_5261);
or U6331 (N_6331,N_5692,N_4334);
or U6332 (N_6332,N_5290,N_5517);
or U6333 (N_6333,N_5149,N_4717);
nand U6334 (N_6334,N_4195,N_4439);
or U6335 (N_6335,N_5507,N_4608);
nor U6336 (N_6336,N_5946,N_5681);
and U6337 (N_6337,N_5964,N_4797);
nand U6338 (N_6338,N_4651,N_5079);
xor U6339 (N_6339,N_4239,N_4592);
or U6340 (N_6340,N_5492,N_5448);
nor U6341 (N_6341,N_5596,N_4348);
nand U6342 (N_6342,N_4603,N_4261);
and U6343 (N_6343,N_4879,N_5830);
nand U6344 (N_6344,N_4416,N_5040);
nor U6345 (N_6345,N_4855,N_5899);
and U6346 (N_6346,N_4546,N_4806);
nor U6347 (N_6347,N_5510,N_4217);
or U6348 (N_6348,N_5767,N_4714);
and U6349 (N_6349,N_5758,N_5231);
nor U6350 (N_6350,N_4858,N_5686);
or U6351 (N_6351,N_5879,N_5411);
or U6352 (N_6352,N_4328,N_5642);
or U6353 (N_6353,N_5499,N_5240);
xor U6354 (N_6354,N_4595,N_4269);
nand U6355 (N_6355,N_5185,N_4552);
nand U6356 (N_6356,N_5531,N_4708);
nor U6357 (N_6357,N_5037,N_4655);
nand U6358 (N_6358,N_4961,N_4194);
and U6359 (N_6359,N_4011,N_5869);
or U6360 (N_6360,N_4831,N_5406);
or U6361 (N_6361,N_4298,N_4999);
or U6362 (N_6362,N_5514,N_4820);
nor U6363 (N_6363,N_5799,N_5366);
or U6364 (N_6364,N_4582,N_4281);
and U6365 (N_6365,N_4695,N_4516);
or U6366 (N_6366,N_5070,N_5316);
nor U6367 (N_6367,N_4370,N_5489);
or U6368 (N_6368,N_4534,N_5148);
nand U6369 (N_6369,N_4013,N_5432);
nand U6370 (N_6370,N_4248,N_4274);
nor U6371 (N_6371,N_5633,N_5821);
and U6372 (N_6372,N_5877,N_4113);
nor U6373 (N_6373,N_4313,N_5140);
and U6374 (N_6374,N_4223,N_5422);
and U6375 (N_6375,N_4368,N_5654);
nor U6376 (N_6376,N_4902,N_4750);
and U6377 (N_6377,N_4887,N_4807);
or U6378 (N_6378,N_4872,N_4036);
and U6379 (N_6379,N_4758,N_4513);
xor U6380 (N_6380,N_5829,N_4725);
nor U6381 (N_6381,N_5468,N_5967);
nor U6382 (N_6382,N_4096,N_4834);
and U6383 (N_6383,N_4074,N_4470);
nor U6384 (N_6384,N_5857,N_5903);
nor U6385 (N_6385,N_4394,N_4580);
and U6386 (N_6386,N_4103,N_4972);
xor U6387 (N_6387,N_4815,N_4181);
nor U6388 (N_6388,N_5268,N_5215);
nand U6389 (N_6389,N_4072,N_4875);
and U6390 (N_6390,N_5110,N_5849);
nor U6391 (N_6391,N_5200,N_5186);
or U6392 (N_6392,N_5447,N_5787);
nor U6393 (N_6393,N_4680,N_4551);
nand U6394 (N_6394,N_4088,N_5480);
nor U6395 (N_6395,N_4624,N_5832);
nand U6396 (N_6396,N_4936,N_4003);
nor U6397 (N_6397,N_4617,N_4069);
nand U6398 (N_6398,N_4417,N_5954);
and U6399 (N_6399,N_5726,N_4210);
nor U6400 (N_6400,N_4317,N_4082);
nand U6401 (N_6401,N_4121,N_4755);
or U6402 (N_6402,N_4387,N_5791);
or U6403 (N_6403,N_5668,N_5357);
xnor U6404 (N_6404,N_4051,N_5753);
nor U6405 (N_6405,N_4346,N_5158);
nand U6406 (N_6406,N_5793,N_5474);
nand U6407 (N_6407,N_5124,N_5605);
nand U6408 (N_6408,N_4959,N_5656);
nand U6409 (N_6409,N_4621,N_5270);
or U6410 (N_6410,N_5688,N_5038);
xnor U6411 (N_6411,N_4712,N_5582);
and U6412 (N_6412,N_4667,N_4773);
nor U6413 (N_6413,N_5963,N_5085);
nand U6414 (N_6414,N_5571,N_5245);
nand U6415 (N_6415,N_5769,N_5023);
and U6416 (N_6416,N_5064,N_4306);
nand U6417 (N_6417,N_5986,N_4744);
nor U6418 (N_6418,N_4674,N_5623);
xnor U6419 (N_6419,N_4662,N_4867);
xnor U6420 (N_6420,N_4090,N_5971);
and U6421 (N_6421,N_5959,N_5028);
and U6422 (N_6422,N_4347,N_4285);
or U6423 (N_6423,N_5014,N_4766);
and U6424 (N_6424,N_5107,N_5359);
or U6425 (N_6425,N_5047,N_5712);
nand U6426 (N_6426,N_4702,N_5678);
and U6427 (N_6427,N_5734,N_5283);
nand U6428 (N_6428,N_4263,N_5455);
nor U6429 (N_6429,N_5837,N_5423);
or U6430 (N_6430,N_4509,N_5090);
or U6431 (N_6431,N_5651,N_4694);
nand U6432 (N_6432,N_4841,N_4352);
or U6433 (N_6433,N_5142,N_5632);
or U6434 (N_6434,N_4507,N_5180);
nand U6435 (N_6435,N_4505,N_4539);
or U6436 (N_6436,N_4928,N_4497);
and U6437 (N_6437,N_4574,N_5896);
or U6438 (N_6438,N_4308,N_4385);
and U6439 (N_6439,N_4251,N_4207);
or U6440 (N_6440,N_5937,N_5084);
or U6441 (N_6441,N_5778,N_5242);
and U6442 (N_6442,N_4264,N_5984);
or U6443 (N_6443,N_5227,N_4633);
and U6444 (N_6444,N_4021,N_5523);
nand U6445 (N_6445,N_5887,N_4421);
nand U6446 (N_6446,N_5773,N_4504);
or U6447 (N_6447,N_5800,N_4292);
or U6448 (N_6448,N_5100,N_5117);
xor U6449 (N_6449,N_4824,N_5009);
nor U6450 (N_6450,N_4735,N_4943);
and U6451 (N_6451,N_5854,N_5700);
and U6452 (N_6452,N_5226,N_4344);
and U6453 (N_6453,N_4878,N_5086);
and U6454 (N_6454,N_5604,N_5181);
nand U6455 (N_6455,N_4788,N_4107);
and U6456 (N_6456,N_5164,N_4782);
and U6457 (N_6457,N_5502,N_4415);
or U6458 (N_6458,N_4550,N_4205);
or U6459 (N_6459,N_4363,N_4793);
xor U6460 (N_6460,N_5171,N_4741);
and U6461 (N_6461,N_4529,N_4984);
and U6462 (N_6462,N_5916,N_4295);
nor U6463 (N_6463,N_4206,N_4353);
nand U6464 (N_6464,N_5034,N_4842);
and U6465 (N_6465,N_5565,N_4101);
and U6466 (N_6466,N_4249,N_4625);
and U6467 (N_6467,N_5694,N_4913);
xnor U6468 (N_6468,N_5440,N_5287);
or U6469 (N_6469,N_5927,N_4299);
nor U6470 (N_6470,N_4396,N_4615);
and U6471 (N_6471,N_4160,N_5119);
nand U6472 (N_6472,N_5533,N_4247);
nand U6473 (N_6473,N_5362,N_4602);
or U6474 (N_6474,N_4890,N_4427);
xor U6475 (N_6475,N_4447,N_4501);
nand U6476 (N_6476,N_4639,N_4757);
nand U6477 (N_6477,N_4326,N_5348);
nor U6478 (N_6478,N_4058,N_5340);
and U6479 (N_6479,N_4258,N_4428);
and U6480 (N_6480,N_4436,N_5383);
or U6481 (N_6481,N_5594,N_5689);
nand U6482 (N_6482,N_5389,N_4889);
and U6483 (N_6483,N_5336,N_4120);
or U6484 (N_6484,N_5626,N_5639);
nand U6485 (N_6485,N_5330,N_4991);
or U6486 (N_6486,N_5951,N_5595);
or U6487 (N_6487,N_5251,N_5528);
and U6488 (N_6488,N_5048,N_5929);
or U6489 (N_6489,N_4726,N_5020);
nor U6490 (N_6490,N_4915,N_5782);
or U6491 (N_6491,N_4312,N_4620);
nand U6492 (N_6492,N_5417,N_4494);
nand U6493 (N_6493,N_5073,N_4386);
nand U6494 (N_6494,N_4496,N_4859);
and U6495 (N_6495,N_4816,N_5392);
xor U6496 (N_6496,N_5179,N_4435);
nand U6497 (N_6497,N_4175,N_5123);
nand U6498 (N_6498,N_4909,N_5576);
nor U6499 (N_6499,N_5325,N_5684);
and U6500 (N_6500,N_4739,N_5513);
and U6501 (N_6501,N_5327,N_4932);
and U6502 (N_6502,N_5647,N_5369);
or U6503 (N_6503,N_4679,N_4211);
xnor U6504 (N_6504,N_4805,N_4723);
nor U6505 (N_6505,N_4464,N_4599);
and U6506 (N_6506,N_4400,N_5690);
nand U6507 (N_6507,N_4813,N_4886);
nor U6508 (N_6508,N_4480,N_5617);
or U6509 (N_6509,N_5036,N_5131);
nand U6510 (N_6510,N_5806,N_5298);
and U6511 (N_6511,N_4970,N_4252);
nor U6512 (N_6512,N_4756,N_5569);
or U6513 (N_6513,N_4402,N_4578);
xnor U6514 (N_6514,N_5053,N_4224);
xnor U6515 (N_6515,N_5414,N_4906);
nor U6516 (N_6516,N_4152,N_5884);
or U6517 (N_6517,N_5888,N_4549);
nand U6518 (N_6518,N_4583,N_5006);
nor U6519 (N_6519,N_5301,N_5702);
nand U6520 (N_6520,N_5912,N_5329);
nand U6521 (N_6521,N_5525,N_5057);
xnor U6522 (N_6522,N_5308,N_4524);
nand U6523 (N_6523,N_4009,N_4031);
and U6524 (N_6524,N_5780,N_5465);
or U6525 (N_6525,N_5522,N_4905);
xor U6526 (N_6526,N_5709,N_5218);
xor U6527 (N_6527,N_4589,N_4271);
nor U6528 (N_6528,N_5208,N_4409);
nand U6529 (N_6529,N_5167,N_5812);
or U6530 (N_6530,N_5861,N_4768);
nor U6531 (N_6531,N_4460,N_5368);
nor U6532 (N_6532,N_4827,N_4451);
nand U6533 (N_6533,N_4981,N_5622);
and U6534 (N_6534,N_4709,N_5415);
or U6535 (N_6535,N_4833,N_4942);
nand U6536 (N_6536,N_4632,N_4449);
nor U6537 (N_6537,N_5239,N_5904);
and U6538 (N_6538,N_5281,N_4327);
nand U6539 (N_6539,N_4606,N_5508);
or U6540 (N_6540,N_5535,N_4077);
xnor U6541 (N_6541,N_4543,N_4491);
nand U6542 (N_6542,N_4333,N_5982);
or U6543 (N_6543,N_5828,N_4637);
or U6544 (N_6544,N_5043,N_5202);
nor U6545 (N_6545,N_5563,N_5552);
and U6546 (N_6546,N_5962,N_4153);
or U6547 (N_6547,N_4657,N_5631);
or U6548 (N_6548,N_4609,N_5918);
or U6549 (N_6549,N_5080,N_4908);
nor U6550 (N_6550,N_4408,N_4303);
and U6551 (N_6551,N_4555,N_4066);
nor U6552 (N_6552,N_4425,N_4931);
nand U6553 (N_6553,N_5932,N_4174);
nor U6554 (N_6554,N_5473,N_5708);
or U6555 (N_6555,N_4325,N_5442);
and U6556 (N_6556,N_5188,N_5628);
nor U6557 (N_6557,N_4520,N_5266);
or U6558 (N_6558,N_5461,N_4838);
nand U6559 (N_6559,N_5989,N_4561);
or U6560 (N_6560,N_4997,N_5321);
nor U6561 (N_6561,N_5795,N_4787);
nand U6562 (N_6562,N_4911,N_5619);
or U6563 (N_6563,N_5957,N_5376);
or U6564 (N_6564,N_4498,N_5317);
and U6565 (N_6565,N_5425,N_4005);
nor U6566 (N_6566,N_4560,N_5915);
and U6567 (N_6567,N_4242,N_5441);
nand U6568 (N_6568,N_4150,N_5677);
and U6569 (N_6569,N_5624,N_4235);
nand U6570 (N_6570,N_4656,N_5731);
nor U6571 (N_6571,N_5534,N_5950);
or U6572 (N_6572,N_5636,N_4988);
nand U6573 (N_6573,N_5742,N_4201);
nand U6574 (N_6574,N_5650,N_5889);
or U6575 (N_6575,N_5802,N_5421);
nand U6576 (N_6576,N_5841,N_4187);
nand U6577 (N_6577,N_4345,N_4500);
nand U6578 (N_6578,N_5463,N_4322);
and U6579 (N_6579,N_5614,N_5745);
nand U6580 (N_6580,N_4136,N_4265);
nand U6581 (N_6581,N_4095,N_5783);
xor U6582 (N_6582,N_5979,N_4343);
or U6583 (N_6583,N_5326,N_5108);
or U6584 (N_6584,N_4759,N_4307);
nand U6585 (N_6585,N_5400,N_4866);
nand U6586 (N_6586,N_4165,N_5867);
nor U6587 (N_6587,N_4482,N_5487);
and U6588 (N_6588,N_4399,N_4623);
nor U6589 (N_6589,N_4067,N_5885);
nand U6590 (N_6590,N_4571,N_4751);
xnor U6591 (N_6591,N_4329,N_5381);
and U6592 (N_6592,N_4042,N_4966);
nand U6593 (N_6593,N_4541,N_4600);
nor U6594 (N_6594,N_4093,N_5503);
or U6595 (N_6595,N_5711,N_5066);
and U6596 (N_6596,N_5558,N_5883);
and U6597 (N_6597,N_4253,N_5752);
nand U6598 (N_6598,N_5012,N_4869);
nor U6599 (N_6599,N_4605,N_4752);
xor U6600 (N_6600,N_4288,N_5516);
xnor U6601 (N_6601,N_5088,N_5958);
nand U6602 (N_6602,N_5856,N_4934);
nor U6603 (N_6603,N_5748,N_5546);
xor U6604 (N_6604,N_5630,N_4413);
and U6605 (N_6605,N_5314,N_4454);
nor U6606 (N_6606,N_5050,N_4364);
and U6607 (N_6607,N_5236,N_5974);
xor U6608 (N_6608,N_5919,N_4554);
and U6609 (N_6609,N_4438,N_5547);
nor U6610 (N_6610,N_5307,N_5491);
or U6611 (N_6611,N_5909,N_5557);
nor U6612 (N_6612,N_5536,N_5811);
and U6613 (N_6613,N_5810,N_4791);
nor U6614 (N_6614,N_4531,N_4459);
and U6615 (N_6615,N_5620,N_4829);
and U6616 (N_6616,N_4047,N_4557);
nor U6617 (N_6617,N_4361,N_4366);
xnor U6618 (N_6618,N_4533,N_5488);
nor U6619 (N_6619,N_4001,N_5871);
or U6620 (N_6620,N_4445,N_5098);
and U6621 (N_6621,N_5693,N_5271);
or U6622 (N_6622,N_5121,N_5332);
nand U6623 (N_6623,N_4716,N_4916);
nand U6624 (N_6624,N_4746,N_5223);
nand U6625 (N_6625,N_5900,N_4277);
and U6626 (N_6626,N_4315,N_5588);
nor U6627 (N_6627,N_5387,N_5095);
and U6628 (N_6628,N_4038,N_5254);
or U6629 (N_6629,N_4721,N_5305);
nor U6630 (N_6630,N_5112,N_5917);
nand U6631 (N_6631,N_5018,N_4351);
nand U6632 (N_6632,N_4819,N_4144);
nand U6633 (N_6633,N_4384,N_4636);
and U6634 (N_6634,N_4706,N_4467);
or U6635 (N_6635,N_5823,N_5980);
and U6636 (N_6636,N_5675,N_4998);
nor U6637 (N_6637,N_5238,N_4779);
nor U6638 (N_6638,N_5930,N_5976);
xor U6639 (N_6639,N_5509,N_5241);
nand U6640 (N_6640,N_4761,N_5848);
nor U6641 (N_6641,N_5797,N_4311);
or U6642 (N_6642,N_5306,N_5874);
nor U6643 (N_6643,N_4958,N_4290);
and U6644 (N_6644,N_4371,N_4700);
or U6645 (N_6645,N_4401,N_5579);
and U6646 (N_6646,N_4874,N_5858);
or U6647 (N_6647,N_4648,N_4899);
nand U6648 (N_6648,N_5350,N_4989);
nand U6649 (N_6649,N_5505,N_4145);
and U6650 (N_6650,N_4236,N_4917);
nor U6651 (N_6651,N_5581,N_5870);
nand U6652 (N_6652,N_5923,N_4965);
nand U6653 (N_6653,N_5126,N_5032);
or U6654 (N_6654,N_4697,N_4579);
and U6655 (N_6655,N_4530,N_5790);
nor U6656 (N_6656,N_4059,N_4562);
xnor U6657 (N_6657,N_4015,N_4511);
or U6658 (N_6658,N_4883,N_5016);
or U6659 (N_6659,N_4267,N_5886);
or U6660 (N_6660,N_5844,N_5106);
or U6661 (N_6661,N_4466,N_4846);
nor U6662 (N_6662,N_5764,N_5029);
and U6663 (N_6663,N_4919,N_4002);
xor U6664 (N_6664,N_5484,N_5166);
xor U6665 (N_6665,N_5153,N_5300);
or U6666 (N_6666,N_5304,N_4469);
and U6667 (N_6667,N_4369,N_5293);
or U6668 (N_6668,N_5172,N_4798);
or U6669 (N_6669,N_5027,N_4473);
nor U6670 (N_6670,N_4068,N_5144);
and U6671 (N_6671,N_5177,N_4442);
nor U6672 (N_6672,N_5189,N_5496);
nand U6673 (N_6673,N_4228,N_4645);
and U6674 (N_6674,N_5135,N_4254);
or U6675 (N_6675,N_4349,N_4666);
or U6676 (N_6676,N_4050,N_5789);
nand U6677 (N_6677,N_4514,N_4502);
or U6678 (N_6678,N_5388,N_4373);
nor U6679 (N_6679,N_5621,N_5341);
nand U6680 (N_6680,N_5059,N_4832);
nand U6681 (N_6681,N_5444,N_5703);
and U6682 (N_6682,N_5999,N_4023);
xnor U6683 (N_6683,N_4764,N_4008);
nand U6684 (N_6684,N_5391,N_4611);
and U6685 (N_6685,N_4510,N_5192);
nand U6686 (N_6686,N_5436,N_4949);
nor U6687 (N_6687,N_4669,N_5021);
or U6688 (N_6688,N_4673,N_4356);
xor U6689 (N_6689,N_5194,N_5248);
or U6690 (N_6690,N_4957,N_5393);
and U6691 (N_6691,N_4868,N_4443);
nand U6692 (N_6692,N_4564,N_5988);
or U6693 (N_6693,N_4440,N_4486);
nor U6694 (N_6694,N_4591,N_5386);
nand U6695 (N_6695,N_5817,N_5754);
and U6696 (N_6696,N_5992,N_4390);
and U6697 (N_6697,N_4976,N_5772);
or U6698 (N_6698,N_5115,N_5356);
or U6699 (N_6699,N_5175,N_4043);
nand U6700 (N_6700,N_4923,N_4300);
and U6701 (N_6701,N_4243,N_4087);
or U6702 (N_6702,N_5007,N_4742);
nand U6703 (N_6703,N_4619,N_4683);
and U6704 (N_6704,N_4671,N_5161);
or U6705 (N_6705,N_4017,N_5673);
and U6706 (N_6706,N_4955,N_5035);
and U6707 (N_6707,N_4032,N_5446);
or U6708 (N_6708,N_5910,N_5019);
and U6709 (N_6709,N_5267,N_5101);
xor U6710 (N_6710,N_5097,N_5138);
nor U6711 (N_6711,N_4587,N_5847);
and U6712 (N_6712,N_5428,N_4771);
nor U6713 (N_6713,N_5687,N_5120);
nand U6714 (N_6714,N_5313,N_5001);
or U6715 (N_6715,N_4176,N_5761);
and U6716 (N_6716,N_4753,N_5490);
or U6717 (N_6717,N_4138,N_5260);
and U6718 (N_6718,N_4596,N_5590);
and U6719 (N_6719,N_4209,N_4940);
nand U6720 (N_6720,N_4020,N_5259);
or U6721 (N_6721,N_5843,N_4339);
xnor U6722 (N_6722,N_4383,N_5157);
or U6723 (N_6723,N_4341,N_5544);
and U6724 (N_6724,N_4629,N_4892);
or U6725 (N_6725,N_5818,N_4367);
nand U6726 (N_6726,N_5431,N_4215);
and U6727 (N_6727,N_5093,N_4661);
nor U6728 (N_6728,N_4105,N_5680);
and U6729 (N_6729,N_4062,N_5501);
nor U6730 (N_6730,N_5291,N_5744);
or U6731 (N_6731,N_4898,N_5452);
nand U6732 (N_6732,N_5424,N_4478);
and U6733 (N_6733,N_5443,N_4168);
nand U6734 (N_6734,N_4986,N_4849);
nor U6735 (N_6735,N_5618,N_5905);
nor U6736 (N_6736,N_4275,N_4643);
or U6737 (N_6737,N_5765,N_5515);
or U6738 (N_6738,N_5952,N_5345);
xnor U6739 (N_6739,N_5863,N_4276);
and U6740 (N_6740,N_4856,N_5659);
or U6741 (N_6741,N_4822,N_5757);
and U6742 (N_6742,N_5649,N_4135);
nand U6743 (N_6743,N_5859,N_4335);
or U6744 (N_6744,N_5367,N_4888);
and U6745 (N_6745,N_5613,N_5970);
or U6746 (N_6746,N_4789,N_5521);
or U6747 (N_6747,N_5746,N_4054);
or U6748 (N_6748,N_5646,N_5670);
nand U6749 (N_6749,N_5908,N_5091);
xnor U6750 (N_6750,N_4607,N_4046);
or U6751 (N_6751,N_5274,N_5527);
and U6752 (N_6752,N_5397,N_4284);
nand U6753 (N_6753,N_5396,N_4131);
and U6754 (N_6754,N_5716,N_5322);
or U6755 (N_6755,N_5560,N_5494);
nand U6756 (N_6756,N_5063,N_5935);
and U6757 (N_6757,N_4775,N_5983);
nor U6758 (N_6758,N_4073,N_5602);
nand U6759 (N_6759,N_5409,N_5384);
xor U6760 (N_6760,N_4448,N_4718);
nor U6761 (N_6761,N_4446,N_5648);
nand U6762 (N_6762,N_5739,N_5603);
nand U6763 (N_6763,N_4056,N_5685);
nor U6764 (N_6764,N_5466,N_5652);
nor U6765 (N_6765,N_5839,N_5222);
or U6766 (N_6766,N_4170,N_5981);
nor U6767 (N_6767,N_5139,N_4654);
xnor U6768 (N_6768,N_4376,N_5735);
xnor U6769 (N_6769,N_4924,N_5697);
or U6770 (N_6770,N_5944,N_4777);
and U6771 (N_6771,N_4601,N_4785);
or U6772 (N_6772,N_4208,N_4558);
and U6773 (N_6773,N_5178,N_4256);
nand U6774 (N_6774,N_5495,N_5825);
nand U6775 (N_6775,N_4028,N_5277);
nor U6776 (N_6776,N_4577,N_4479);
and U6777 (N_6777,N_4226,N_4393);
or U6778 (N_6778,N_4681,N_5719);
nor U6779 (N_6779,N_4544,N_5747);
nand U6780 (N_6780,N_5786,N_4109);
or U6781 (N_6781,N_5134,N_4729);
and U6782 (N_6782,N_4037,N_5334);
or U6783 (N_6783,N_5529,N_5229);
and U6784 (N_6784,N_4179,N_4678);
or U6785 (N_6785,N_5897,N_4538);
and U6786 (N_6786,N_4010,N_5815);
nand U6787 (N_6787,N_5575,N_5343);
or U6788 (N_6788,N_4780,N_5111);
and U6789 (N_6789,N_4412,N_5714);
nand U6790 (N_6790,N_4419,N_5017);
or U6791 (N_6791,N_4907,N_5725);
nand U6792 (N_6792,N_5607,N_5902);
and U6793 (N_6793,N_4626,N_5160);
nand U6794 (N_6794,N_4812,N_5938);
and U6795 (N_6795,N_4063,N_5087);
and U6796 (N_6796,N_5635,N_4638);
and U6797 (N_6797,N_5205,N_4049);
and U6798 (N_6798,N_5358,N_5479);
nand U6799 (N_6799,N_5114,N_4272);
nor U6800 (N_6800,N_4670,N_4336);
or U6801 (N_6801,N_5410,N_5634);
and U6802 (N_6802,N_4414,N_5454);
nor U6803 (N_6803,N_4323,N_5010);
nand U6804 (N_6804,N_5377,N_5987);
or U6805 (N_6805,N_4992,N_5453);
or U6806 (N_6806,N_5794,N_5833);
nand U6807 (N_6807,N_5003,N_4774);
nor U6808 (N_6808,N_5116,N_5933);
and U6809 (N_6809,N_5597,N_4594);
nor U6810 (N_6810,N_5089,N_5058);
and U6811 (N_6811,N_5318,N_5704);
nand U6812 (N_6812,N_4614,N_4092);
nand U6813 (N_6813,N_5147,N_5741);
nand U6814 (N_6814,N_5176,N_4314);
or U6815 (N_6815,N_5201,N_4663);
nand U6816 (N_6816,N_5591,N_4945);
and U6817 (N_6817,N_4593,N_5801);
and U6818 (N_6818,N_5997,N_5485);
nor U6819 (N_6819,N_4222,N_5788);
xnor U6820 (N_6820,N_4641,N_4434);
nand U6821 (N_6821,N_4877,N_4665);
nand U6822 (N_6822,N_4971,N_4305);
or U6823 (N_6823,N_5555,N_5803);
nor U6824 (N_6824,N_4476,N_4340);
nor U6825 (N_6825,N_4649,N_4525);
or U6826 (N_6826,N_5852,N_4848);
and U6827 (N_6827,N_4996,N_4155);
and U6828 (N_6828,N_5438,N_5408);
or U6829 (N_6829,N_5339,N_5814);
nor U6830 (N_6830,N_5845,N_4012);
nand U6831 (N_6831,N_5292,N_5538);
xnor U6832 (N_6832,N_4422,N_5041);
nand U6833 (N_6833,N_5842,N_4952);
nand U6834 (N_6834,N_5353,N_5566);
nand U6835 (N_6835,N_5182,N_4508);
nor U6836 (N_6836,N_5943,N_4372);
nor U6837 (N_6837,N_5822,N_5033);
and U6838 (N_6838,N_4743,N_5760);
xnor U6839 (N_6839,N_4947,N_5749);
nand U6840 (N_6840,N_5407,N_5667);
xor U6841 (N_6841,N_5931,N_5128);
or U6842 (N_6842,N_5403,N_4647);
and U6843 (N_6843,N_4374,N_5868);
nand U6844 (N_6844,N_5249,N_5733);
and U6845 (N_6845,N_4770,N_5567);
nand U6846 (N_6846,N_5660,N_4320);
xnor U6847 (N_6847,N_5127,N_4332);
and U6848 (N_6848,N_4410,N_5550);
or U6849 (N_6849,N_4880,N_5759);
and U6850 (N_6850,N_5891,N_4019);
nand U6851 (N_6851,N_5413,N_5211);
or U6852 (N_6852,N_5500,N_5809);
xor U6853 (N_6853,N_4159,N_4468);
nand U6854 (N_6854,N_5898,N_5419);
xor U6855 (N_6855,N_4186,N_4027);
and U6856 (N_6856,N_4630,N_5420);
and U6857 (N_6857,N_5601,N_5669);
or U6858 (N_6858,N_4190,N_4282);
nor U6859 (N_6859,N_5137,N_4184);
nor U6860 (N_6860,N_5328,N_5972);
nor U6861 (N_6861,N_5237,N_5482);
and U6862 (N_6862,N_4749,N_5965);
nor U6863 (N_6863,N_5750,N_5562);
nand U6864 (N_6864,N_5228,N_4720);
or U6865 (N_6865,N_4430,N_5262);
nand U6866 (N_6866,N_4732,N_5751);
nor U6867 (N_6867,N_5705,N_4873);
nand U6868 (N_6868,N_4318,N_5472);
and U6869 (N_6869,N_4968,N_4799);
xnor U6870 (N_6870,N_4631,N_4360);
or U6871 (N_6871,N_4240,N_4122);
nor U6872 (N_6872,N_5718,N_5136);
or U6873 (N_6873,N_5275,N_4233);
nand U6874 (N_6874,N_4930,N_4588);
nand U6875 (N_6875,N_5740,N_4828);
nand U6876 (N_6876,N_4169,N_4091);
nand U6877 (N_6877,N_4830,N_5052);
nor U6878 (N_6878,N_5005,N_5599);
nand U6879 (N_6879,N_4041,N_4030);
or U6880 (N_6880,N_4825,N_5372);
nand U6881 (N_6881,N_4108,N_4584);
xnor U6882 (N_6882,N_5715,N_4127);
nand U6883 (N_6883,N_5082,N_4676);
nand U6884 (N_6884,N_5717,N_5067);
or U6885 (N_6885,N_4452,N_4128);
nand U6886 (N_6886,N_5445,N_5434);
and U6887 (N_6887,N_4116,N_4193);
nand U6888 (N_6888,N_4705,N_5530);
or U6889 (N_6889,N_4405,N_5206);
and U6890 (N_6890,N_5342,N_4572);
or U6891 (N_6891,N_4559,N_5722);
nor U6892 (N_6892,N_4147,N_5289);
nor U6893 (N_6893,N_5486,N_5637);
nand U6894 (N_6894,N_5429,N_4635);
nand U6895 (N_6895,N_5679,N_5130);
xnor U6896 (N_6896,N_5146,N_4762);
nor U6897 (N_6897,N_4033,N_4237);
nand U6898 (N_6898,N_5113,N_5696);
and U6899 (N_6899,N_4922,N_5364);
or U6900 (N_6900,N_5399,N_4230);
nand U6901 (N_6901,N_5713,N_5914);
or U6902 (N_6902,N_4894,N_5214);
nor U6903 (N_6903,N_5850,N_4781);
nand U6904 (N_6904,N_4990,N_4567);
or U6905 (N_6905,N_5000,N_4331);
and U6906 (N_6906,N_4296,N_4026);
nor U6907 (N_6907,N_5629,N_5279);
or U6908 (N_6908,N_4119,N_4950);
or U6909 (N_6909,N_4006,N_4309);
xnor U6910 (N_6910,N_4573,N_5295);
nor U6911 (N_6911,N_4378,N_5512);
nor U6912 (N_6912,N_4960,N_5244);
nand U6913 (N_6913,N_5498,N_5732);
or U6914 (N_6914,N_4612,N_5526);
xnor U6915 (N_6915,N_5233,N_4148);
xor U6916 (N_6916,N_4865,N_4724);
and U6917 (N_6917,N_4357,N_4845);
and U6918 (N_6918,N_5155,N_5600);
xnor U6919 (N_6919,N_4268,N_4840);
nor U6920 (N_6920,N_4149,N_4642);
nor U6921 (N_6921,N_5247,N_4569);
or U6922 (N_6922,N_5154,N_5303);
and U6923 (N_6923,N_5191,N_4097);
or U6924 (N_6924,N_4007,N_5655);
or U6925 (N_6925,N_4711,N_5587);
and U6926 (N_6926,N_5574,N_5163);
and U6927 (N_6927,N_5437,N_5723);
and U6928 (N_6928,N_5784,N_5736);
or U6929 (N_6929,N_4407,N_5346);
and U6930 (N_6930,N_4650,N_5068);
nand U6931 (N_6931,N_4203,N_4398);
and U6932 (N_6932,N_4664,N_4566);
and U6933 (N_6933,N_5196,N_5374);
and U6934 (N_6934,N_5210,N_5851);
nand U6935 (N_6935,N_5730,N_4304);
and U6936 (N_6936,N_4542,N_4084);
and U6937 (N_6937,N_5083,N_5265);
nand U6938 (N_6938,N_5808,N_4474);
nand U6939 (N_6939,N_5056,N_4713);
nor U6940 (N_6940,N_5762,N_4310);
nor U6941 (N_6941,N_4130,N_4796);
nor U6942 (N_6942,N_4738,N_5872);
nand U6943 (N_6943,N_5320,N_5288);
nor U6944 (N_6944,N_4926,N_5337);
nand U6945 (N_6945,N_4710,N_4548);
nand U6946 (N_6946,N_5152,N_5213);
nor U6947 (N_6947,N_5551,N_5462);
and U6948 (N_6948,N_5302,N_5961);
and U6949 (N_6949,N_4760,N_4565);
nor U6950 (N_6950,N_5539,N_5481);
nand U6951 (N_6951,N_4535,N_5168);
or U6952 (N_6952,N_4259,N_4173);
nor U6953 (N_6953,N_4585,N_4707);
or U6954 (N_6954,N_5450,N_4545);
nand U6955 (N_6955,N_4462,N_5866);
and U6956 (N_6956,N_4857,N_5674);
or U6957 (N_6957,N_5284,N_5143);
nor U6958 (N_6958,N_5243,N_5598);
nor U6959 (N_6959,N_5925,N_4672);
nand U6960 (N_6960,N_5813,N_5278);
or U6961 (N_6961,N_4521,N_4250);
nor U6962 (N_6962,N_5234,N_4225);
xor U6963 (N_6963,N_4745,N_4156);
xor U6964 (N_6964,N_5913,N_5165);
nor U6965 (N_6965,N_5721,N_4388);
nand U6966 (N_6966,N_4493,N_5333);
or U6967 (N_6967,N_4835,N_5831);
and U6968 (N_6968,N_4929,N_5771);
xnor U6969 (N_6969,N_4918,N_5197);
nand U6970 (N_6970,N_5039,N_5664);
nand U6971 (N_6971,N_4946,N_5004);
nor U6972 (N_6972,N_4795,N_5662);
nand U6973 (N_6973,N_5589,N_5046);
and U6974 (N_6974,N_4882,N_4912);
nand U6975 (N_6975,N_5351,N_4411);
or U6976 (N_6976,N_4106,N_4178);
nor U6977 (N_6977,N_5187,N_4065);
and U6978 (N_6978,N_4980,N_5471);
and U6979 (N_6979,N_4783,N_4350);
and U6980 (N_6980,N_4484,N_4132);
nand U6981 (N_6981,N_4490,N_4424);
and U6982 (N_6982,N_4018,N_5548);
nand U6983 (N_6983,N_4993,N_4189);
nand U6984 (N_6984,N_4995,N_5257);
nand U6985 (N_6985,N_5840,N_5272);
and U6986 (N_6986,N_4597,N_4202);
or U6987 (N_6987,N_5380,N_4733);
xor U6988 (N_6988,N_4004,N_5568);
or U6989 (N_6989,N_5616,N_5657);
nand U6990 (N_6990,N_4598,N_4982);
and U6991 (N_6991,N_4182,N_4283);
and U6992 (N_6992,N_4575,N_5663);
or U6993 (N_6993,N_5008,N_4291);
xor U6994 (N_6994,N_4083,N_4684);
nand U6995 (N_6995,N_4216,N_4893);
or U6996 (N_6996,N_4696,N_4433);
nor U6997 (N_6997,N_4163,N_5948);
and U6998 (N_6998,N_5834,N_5578);
or U6999 (N_6999,N_5945,N_5216);
xnor U7000 (N_7000,N_5857,N_5043);
or U7001 (N_7001,N_4701,N_5551);
xnor U7002 (N_7002,N_5629,N_5668);
or U7003 (N_7003,N_4138,N_4997);
and U7004 (N_7004,N_5336,N_5166);
nand U7005 (N_7005,N_4806,N_4165);
nand U7006 (N_7006,N_4724,N_4836);
and U7007 (N_7007,N_5229,N_5772);
and U7008 (N_7008,N_5933,N_5618);
or U7009 (N_7009,N_5244,N_4330);
and U7010 (N_7010,N_4570,N_5764);
or U7011 (N_7011,N_4177,N_5864);
xnor U7012 (N_7012,N_5245,N_5802);
nand U7013 (N_7013,N_5001,N_5917);
or U7014 (N_7014,N_5455,N_4112);
and U7015 (N_7015,N_4958,N_4944);
nand U7016 (N_7016,N_5046,N_5399);
and U7017 (N_7017,N_5370,N_5422);
xor U7018 (N_7018,N_4995,N_5899);
or U7019 (N_7019,N_5652,N_5029);
nor U7020 (N_7020,N_5110,N_4577);
nor U7021 (N_7021,N_5177,N_5013);
and U7022 (N_7022,N_5860,N_4940);
and U7023 (N_7023,N_5455,N_4248);
nor U7024 (N_7024,N_5924,N_4279);
or U7025 (N_7025,N_5928,N_5535);
xnor U7026 (N_7026,N_5468,N_4262);
nand U7027 (N_7027,N_4795,N_5898);
or U7028 (N_7028,N_5363,N_5305);
nor U7029 (N_7029,N_5001,N_5619);
or U7030 (N_7030,N_4859,N_5660);
or U7031 (N_7031,N_4419,N_4410);
or U7032 (N_7032,N_5578,N_4358);
and U7033 (N_7033,N_5131,N_5160);
xor U7034 (N_7034,N_5277,N_4055);
and U7035 (N_7035,N_5621,N_5894);
and U7036 (N_7036,N_5110,N_5061);
and U7037 (N_7037,N_5332,N_4265);
and U7038 (N_7038,N_5951,N_5377);
nor U7039 (N_7039,N_4596,N_5898);
or U7040 (N_7040,N_4913,N_5206);
nor U7041 (N_7041,N_4024,N_4797);
nor U7042 (N_7042,N_5955,N_4128);
and U7043 (N_7043,N_4950,N_4819);
and U7044 (N_7044,N_4231,N_5994);
nand U7045 (N_7045,N_4671,N_4173);
or U7046 (N_7046,N_5250,N_4698);
and U7047 (N_7047,N_4933,N_4859);
nand U7048 (N_7048,N_5783,N_5506);
nand U7049 (N_7049,N_4513,N_4576);
xnor U7050 (N_7050,N_5803,N_5406);
nor U7051 (N_7051,N_4150,N_4071);
and U7052 (N_7052,N_5202,N_4528);
and U7053 (N_7053,N_5667,N_4412);
or U7054 (N_7054,N_5798,N_4798);
or U7055 (N_7055,N_5846,N_4379);
nor U7056 (N_7056,N_5684,N_4996);
or U7057 (N_7057,N_5212,N_4727);
xor U7058 (N_7058,N_5349,N_4121);
or U7059 (N_7059,N_5700,N_4707);
or U7060 (N_7060,N_5419,N_4202);
nand U7061 (N_7061,N_4587,N_5152);
nor U7062 (N_7062,N_4415,N_5179);
nor U7063 (N_7063,N_4317,N_5492);
nand U7064 (N_7064,N_5893,N_5664);
nor U7065 (N_7065,N_4101,N_5951);
nor U7066 (N_7066,N_4537,N_4601);
or U7067 (N_7067,N_5156,N_4671);
nand U7068 (N_7068,N_5991,N_4938);
and U7069 (N_7069,N_4471,N_5712);
nor U7070 (N_7070,N_4542,N_4128);
and U7071 (N_7071,N_5921,N_4784);
or U7072 (N_7072,N_4176,N_4673);
and U7073 (N_7073,N_4579,N_4534);
or U7074 (N_7074,N_4447,N_4319);
nand U7075 (N_7075,N_5898,N_4314);
nand U7076 (N_7076,N_5288,N_5258);
xor U7077 (N_7077,N_5265,N_4226);
nor U7078 (N_7078,N_4763,N_4943);
nand U7079 (N_7079,N_5314,N_5734);
nor U7080 (N_7080,N_5399,N_5902);
or U7081 (N_7081,N_5832,N_5059);
nor U7082 (N_7082,N_4778,N_4275);
nand U7083 (N_7083,N_4218,N_5655);
nor U7084 (N_7084,N_5739,N_4314);
nand U7085 (N_7085,N_5909,N_5440);
or U7086 (N_7086,N_5591,N_4923);
nand U7087 (N_7087,N_4730,N_4353);
nand U7088 (N_7088,N_5838,N_5979);
nor U7089 (N_7089,N_4576,N_5551);
xor U7090 (N_7090,N_5497,N_4862);
nand U7091 (N_7091,N_4486,N_5111);
or U7092 (N_7092,N_4194,N_4110);
and U7093 (N_7093,N_5928,N_4494);
nand U7094 (N_7094,N_5994,N_4017);
nand U7095 (N_7095,N_4589,N_4606);
xor U7096 (N_7096,N_5829,N_5267);
nand U7097 (N_7097,N_4579,N_5488);
or U7098 (N_7098,N_5618,N_5199);
nand U7099 (N_7099,N_4233,N_4818);
xor U7100 (N_7100,N_5542,N_5527);
nand U7101 (N_7101,N_5297,N_5189);
and U7102 (N_7102,N_5689,N_5226);
or U7103 (N_7103,N_5803,N_4929);
or U7104 (N_7104,N_4878,N_5610);
and U7105 (N_7105,N_4428,N_5934);
nand U7106 (N_7106,N_4673,N_4650);
or U7107 (N_7107,N_4657,N_4209);
or U7108 (N_7108,N_4326,N_5136);
nor U7109 (N_7109,N_4205,N_4520);
nand U7110 (N_7110,N_4230,N_5321);
nand U7111 (N_7111,N_5066,N_4807);
nor U7112 (N_7112,N_5360,N_5840);
nand U7113 (N_7113,N_5731,N_4187);
and U7114 (N_7114,N_5172,N_4969);
or U7115 (N_7115,N_5674,N_4411);
and U7116 (N_7116,N_4192,N_4332);
nand U7117 (N_7117,N_5923,N_4298);
or U7118 (N_7118,N_5522,N_4989);
or U7119 (N_7119,N_5016,N_4503);
and U7120 (N_7120,N_5635,N_5365);
or U7121 (N_7121,N_5596,N_5550);
nor U7122 (N_7122,N_4810,N_4257);
and U7123 (N_7123,N_4869,N_4916);
and U7124 (N_7124,N_5083,N_5713);
or U7125 (N_7125,N_5253,N_5718);
and U7126 (N_7126,N_5339,N_5246);
and U7127 (N_7127,N_5431,N_4559);
nand U7128 (N_7128,N_4803,N_5903);
nor U7129 (N_7129,N_4509,N_4293);
and U7130 (N_7130,N_5672,N_4874);
nand U7131 (N_7131,N_4221,N_5776);
and U7132 (N_7132,N_5434,N_5959);
and U7133 (N_7133,N_5152,N_5482);
and U7134 (N_7134,N_5940,N_4625);
xnor U7135 (N_7135,N_4247,N_5598);
xnor U7136 (N_7136,N_4860,N_4884);
or U7137 (N_7137,N_4203,N_4102);
or U7138 (N_7138,N_5556,N_5352);
and U7139 (N_7139,N_4159,N_5191);
and U7140 (N_7140,N_4436,N_4537);
and U7141 (N_7141,N_5301,N_5947);
xnor U7142 (N_7142,N_5603,N_4375);
and U7143 (N_7143,N_4923,N_5267);
nand U7144 (N_7144,N_5497,N_5834);
xnor U7145 (N_7145,N_5872,N_5094);
and U7146 (N_7146,N_5462,N_4719);
or U7147 (N_7147,N_4137,N_5987);
nor U7148 (N_7148,N_5317,N_4276);
nor U7149 (N_7149,N_4349,N_4787);
nand U7150 (N_7150,N_5262,N_5670);
and U7151 (N_7151,N_5560,N_5572);
nor U7152 (N_7152,N_4301,N_5757);
nor U7153 (N_7153,N_5800,N_5965);
nor U7154 (N_7154,N_4449,N_4707);
xor U7155 (N_7155,N_5640,N_5900);
xnor U7156 (N_7156,N_4156,N_5456);
or U7157 (N_7157,N_4954,N_5863);
and U7158 (N_7158,N_4684,N_4058);
or U7159 (N_7159,N_4635,N_5742);
nand U7160 (N_7160,N_4889,N_4116);
or U7161 (N_7161,N_5697,N_5144);
or U7162 (N_7162,N_5974,N_4452);
and U7163 (N_7163,N_5083,N_4957);
nand U7164 (N_7164,N_5683,N_4844);
or U7165 (N_7165,N_5082,N_5004);
xor U7166 (N_7166,N_5892,N_4988);
nand U7167 (N_7167,N_4036,N_4071);
or U7168 (N_7168,N_5038,N_4103);
nand U7169 (N_7169,N_4812,N_5370);
nand U7170 (N_7170,N_4904,N_5373);
nor U7171 (N_7171,N_4908,N_5081);
nand U7172 (N_7172,N_5180,N_4341);
or U7173 (N_7173,N_4950,N_5517);
and U7174 (N_7174,N_5284,N_4240);
and U7175 (N_7175,N_5215,N_5694);
xor U7176 (N_7176,N_5188,N_5414);
nand U7177 (N_7177,N_5103,N_5007);
nand U7178 (N_7178,N_4991,N_5349);
nand U7179 (N_7179,N_5795,N_4047);
and U7180 (N_7180,N_5786,N_5625);
or U7181 (N_7181,N_5318,N_5915);
and U7182 (N_7182,N_5518,N_5257);
nand U7183 (N_7183,N_5882,N_4395);
nor U7184 (N_7184,N_4803,N_5435);
nand U7185 (N_7185,N_4425,N_4110);
and U7186 (N_7186,N_4267,N_4968);
xnor U7187 (N_7187,N_5130,N_5910);
nand U7188 (N_7188,N_5016,N_4529);
nor U7189 (N_7189,N_4812,N_5388);
nor U7190 (N_7190,N_4290,N_4730);
nand U7191 (N_7191,N_4022,N_5193);
or U7192 (N_7192,N_5827,N_5971);
nand U7193 (N_7193,N_4637,N_5937);
or U7194 (N_7194,N_5631,N_5872);
or U7195 (N_7195,N_5716,N_5910);
and U7196 (N_7196,N_4118,N_4527);
or U7197 (N_7197,N_4654,N_4269);
nor U7198 (N_7198,N_5624,N_5921);
and U7199 (N_7199,N_4514,N_5263);
or U7200 (N_7200,N_4610,N_5921);
nor U7201 (N_7201,N_4949,N_5983);
and U7202 (N_7202,N_4035,N_4297);
xor U7203 (N_7203,N_4886,N_4508);
nor U7204 (N_7204,N_5829,N_5237);
nand U7205 (N_7205,N_4091,N_5169);
nand U7206 (N_7206,N_4784,N_4204);
nor U7207 (N_7207,N_5033,N_4702);
and U7208 (N_7208,N_5885,N_4338);
xor U7209 (N_7209,N_5036,N_5438);
or U7210 (N_7210,N_5357,N_4056);
or U7211 (N_7211,N_4505,N_5561);
nor U7212 (N_7212,N_4371,N_5160);
and U7213 (N_7213,N_5866,N_5052);
and U7214 (N_7214,N_4942,N_4350);
and U7215 (N_7215,N_4066,N_4944);
or U7216 (N_7216,N_4990,N_5220);
xor U7217 (N_7217,N_5442,N_4843);
and U7218 (N_7218,N_5130,N_5676);
or U7219 (N_7219,N_5355,N_5064);
nand U7220 (N_7220,N_5782,N_4010);
or U7221 (N_7221,N_4673,N_4143);
or U7222 (N_7222,N_4986,N_5355);
xnor U7223 (N_7223,N_5253,N_5473);
and U7224 (N_7224,N_4814,N_4831);
and U7225 (N_7225,N_4052,N_5966);
nand U7226 (N_7226,N_5719,N_4750);
nand U7227 (N_7227,N_4089,N_5113);
nand U7228 (N_7228,N_5547,N_5071);
or U7229 (N_7229,N_4915,N_5930);
xnor U7230 (N_7230,N_5385,N_4192);
nor U7231 (N_7231,N_4575,N_4903);
nor U7232 (N_7232,N_4814,N_4590);
nand U7233 (N_7233,N_5989,N_4889);
nand U7234 (N_7234,N_5022,N_5615);
nand U7235 (N_7235,N_4788,N_5958);
or U7236 (N_7236,N_4172,N_5174);
nand U7237 (N_7237,N_4750,N_4674);
nor U7238 (N_7238,N_5084,N_4490);
and U7239 (N_7239,N_4455,N_4576);
or U7240 (N_7240,N_5561,N_5057);
nor U7241 (N_7241,N_4014,N_4777);
nand U7242 (N_7242,N_5506,N_5341);
and U7243 (N_7243,N_4471,N_5884);
or U7244 (N_7244,N_5528,N_5308);
nor U7245 (N_7245,N_5997,N_4510);
nand U7246 (N_7246,N_4491,N_5127);
and U7247 (N_7247,N_5407,N_4266);
nor U7248 (N_7248,N_4065,N_5363);
nor U7249 (N_7249,N_5250,N_5008);
nor U7250 (N_7250,N_5653,N_4959);
or U7251 (N_7251,N_5776,N_5995);
or U7252 (N_7252,N_4638,N_4937);
and U7253 (N_7253,N_4770,N_5190);
nand U7254 (N_7254,N_4814,N_5036);
and U7255 (N_7255,N_5649,N_5393);
and U7256 (N_7256,N_4721,N_5974);
nor U7257 (N_7257,N_5296,N_5629);
xnor U7258 (N_7258,N_5284,N_4416);
nor U7259 (N_7259,N_4945,N_5611);
or U7260 (N_7260,N_5347,N_5074);
nand U7261 (N_7261,N_5086,N_5960);
nor U7262 (N_7262,N_4935,N_5723);
nor U7263 (N_7263,N_4407,N_5657);
nor U7264 (N_7264,N_4048,N_4513);
and U7265 (N_7265,N_5427,N_4378);
nor U7266 (N_7266,N_5522,N_4555);
xor U7267 (N_7267,N_5915,N_5488);
or U7268 (N_7268,N_5351,N_5016);
and U7269 (N_7269,N_4870,N_4107);
or U7270 (N_7270,N_4608,N_5219);
and U7271 (N_7271,N_4469,N_5106);
nand U7272 (N_7272,N_4156,N_4548);
nand U7273 (N_7273,N_4565,N_5798);
nand U7274 (N_7274,N_4131,N_5179);
nand U7275 (N_7275,N_5260,N_4976);
nand U7276 (N_7276,N_4206,N_4262);
nor U7277 (N_7277,N_4332,N_5408);
and U7278 (N_7278,N_5850,N_4805);
and U7279 (N_7279,N_5211,N_4590);
and U7280 (N_7280,N_4513,N_4488);
nand U7281 (N_7281,N_4537,N_4252);
nand U7282 (N_7282,N_4503,N_4983);
and U7283 (N_7283,N_5873,N_5937);
or U7284 (N_7284,N_5205,N_5493);
xor U7285 (N_7285,N_4083,N_5168);
nor U7286 (N_7286,N_5695,N_5776);
or U7287 (N_7287,N_4064,N_5869);
and U7288 (N_7288,N_5311,N_4187);
xnor U7289 (N_7289,N_5157,N_5931);
nor U7290 (N_7290,N_4649,N_5080);
nand U7291 (N_7291,N_5891,N_4003);
and U7292 (N_7292,N_4580,N_5104);
nor U7293 (N_7293,N_5173,N_4090);
xnor U7294 (N_7294,N_4451,N_4234);
and U7295 (N_7295,N_4626,N_5734);
or U7296 (N_7296,N_4025,N_5703);
nand U7297 (N_7297,N_5213,N_5204);
nor U7298 (N_7298,N_4358,N_5152);
nor U7299 (N_7299,N_5877,N_5663);
xnor U7300 (N_7300,N_5649,N_4107);
and U7301 (N_7301,N_4054,N_5306);
xnor U7302 (N_7302,N_5866,N_4563);
nor U7303 (N_7303,N_4227,N_4137);
xnor U7304 (N_7304,N_4028,N_5780);
or U7305 (N_7305,N_4314,N_4347);
nor U7306 (N_7306,N_5698,N_5831);
nand U7307 (N_7307,N_5159,N_5490);
nor U7308 (N_7308,N_4818,N_5370);
nor U7309 (N_7309,N_5329,N_4598);
and U7310 (N_7310,N_5728,N_4976);
nor U7311 (N_7311,N_4195,N_4496);
and U7312 (N_7312,N_4276,N_4569);
nand U7313 (N_7313,N_5718,N_5060);
xnor U7314 (N_7314,N_5184,N_5977);
nor U7315 (N_7315,N_4228,N_4531);
or U7316 (N_7316,N_5360,N_5706);
nor U7317 (N_7317,N_4464,N_5052);
nor U7318 (N_7318,N_5406,N_5765);
or U7319 (N_7319,N_5783,N_5754);
or U7320 (N_7320,N_4837,N_4409);
or U7321 (N_7321,N_4508,N_5650);
nor U7322 (N_7322,N_4926,N_4053);
nor U7323 (N_7323,N_5736,N_5259);
nor U7324 (N_7324,N_4680,N_5194);
nand U7325 (N_7325,N_5102,N_4564);
nor U7326 (N_7326,N_5895,N_5729);
or U7327 (N_7327,N_4260,N_5931);
or U7328 (N_7328,N_4114,N_4818);
or U7329 (N_7329,N_4594,N_5423);
or U7330 (N_7330,N_5093,N_4275);
nor U7331 (N_7331,N_5275,N_5985);
and U7332 (N_7332,N_4929,N_5978);
nor U7333 (N_7333,N_5070,N_5936);
or U7334 (N_7334,N_5420,N_4148);
or U7335 (N_7335,N_5021,N_5192);
or U7336 (N_7336,N_4921,N_4208);
nor U7337 (N_7337,N_5045,N_5177);
and U7338 (N_7338,N_5692,N_5272);
or U7339 (N_7339,N_4016,N_4272);
xnor U7340 (N_7340,N_4334,N_5068);
xor U7341 (N_7341,N_4862,N_5956);
or U7342 (N_7342,N_4746,N_4957);
nor U7343 (N_7343,N_4881,N_5268);
nor U7344 (N_7344,N_4469,N_4828);
nor U7345 (N_7345,N_5311,N_4464);
or U7346 (N_7346,N_5793,N_4181);
or U7347 (N_7347,N_5618,N_5570);
nand U7348 (N_7348,N_4571,N_4335);
nand U7349 (N_7349,N_5307,N_4147);
and U7350 (N_7350,N_4508,N_4959);
nor U7351 (N_7351,N_4194,N_5280);
nand U7352 (N_7352,N_5349,N_5787);
or U7353 (N_7353,N_4940,N_5432);
nand U7354 (N_7354,N_5948,N_5384);
xnor U7355 (N_7355,N_5621,N_5270);
nand U7356 (N_7356,N_5793,N_4786);
or U7357 (N_7357,N_5252,N_5421);
and U7358 (N_7358,N_5593,N_4334);
nor U7359 (N_7359,N_5783,N_5653);
or U7360 (N_7360,N_5046,N_5771);
xor U7361 (N_7361,N_4635,N_4006);
and U7362 (N_7362,N_5111,N_5404);
nand U7363 (N_7363,N_5049,N_4400);
and U7364 (N_7364,N_5380,N_5273);
and U7365 (N_7365,N_5433,N_5839);
or U7366 (N_7366,N_4618,N_5101);
nor U7367 (N_7367,N_4212,N_4894);
or U7368 (N_7368,N_4575,N_4170);
or U7369 (N_7369,N_5648,N_4807);
nor U7370 (N_7370,N_4142,N_4766);
and U7371 (N_7371,N_4149,N_4063);
or U7372 (N_7372,N_4397,N_4533);
nand U7373 (N_7373,N_5366,N_5223);
nor U7374 (N_7374,N_5276,N_4305);
or U7375 (N_7375,N_4992,N_4278);
nor U7376 (N_7376,N_4417,N_4352);
xnor U7377 (N_7377,N_5896,N_4939);
or U7378 (N_7378,N_5041,N_4151);
nand U7379 (N_7379,N_4646,N_4236);
nand U7380 (N_7380,N_4664,N_4456);
nor U7381 (N_7381,N_5594,N_4679);
xnor U7382 (N_7382,N_4413,N_5425);
and U7383 (N_7383,N_5827,N_5745);
nor U7384 (N_7384,N_5407,N_4408);
nand U7385 (N_7385,N_5968,N_4082);
or U7386 (N_7386,N_4887,N_4868);
and U7387 (N_7387,N_4703,N_5607);
nand U7388 (N_7388,N_5724,N_5845);
and U7389 (N_7389,N_5497,N_5710);
nand U7390 (N_7390,N_5326,N_5941);
nand U7391 (N_7391,N_4892,N_4979);
or U7392 (N_7392,N_4377,N_4198);
nand U7393 (N_7393,N_5091,N_5872);
or U7394 (N_7394,N_5186,N_5926);
nand U7395 (N_7395,N_4836,N_4076);
or U7396 (N_7396,N_5603,N_5880);
and U7397 (N_7397,N_4498,N_5205);
or U7398 (N_7398,N_4658,N_5450);
nand U7399 (N_7399,N_5969,N_5717);
nand U7400 (N_7400,N_4941,N_4798);
or U7401 (N_7401,N_5751,N_4772);
and U7402 (N_7402,N_4589,N_4863);
nor U7403 (N_7403,N_5241,N_5175);
and U7404 (N_7404,N_5715,N_5628);
nand U7405 (N_7405,N_4682,N_4075);
xnor U7406 (N_7406,N_5066,N_5450);
and U7407 (N_7407,N_5747,N_4742);
nand U7408 (N_7408,N_5123,N_4138);
and U7409 (N_7409,N_4350,N_5238);
nor U7410 (N_7410,N_4039,N_4333);
or U7411 (N_7411,N_5343,N_4113);
nor U7412 (N_7412,N_5434,N_4176);
or U7413 (N_7413,N_5138,N_5150);
nand U7414 (N_7414,N_4953,N_4563);
nand U7415 (N_7415,N_5916,N_5911);
nand U7416 (N_7416,N_5894,N_5627);
or U7417 (N_7417,N_4109,N_4434);
xor U7418 (N_7418,N_5985,N_5302);
nand U7419 (N_7419,N_5950,N_4709);
and U7420 (N_7420,N_4142,N_4720);
nand U7421 (N_7421,N_5526,N_4789);
or U7422 (N_7422,N_4859,N_4098);
xnor U7423 (N_7423,N_4501,N_4311);
or U7424 (N_7424,N_5988,N_4655);
or U7425 (N_7425,N_4380,N_4444);
xor U7426 (N_7426,N_5435,N_5348);
or U7427 (N_7427,N_4915,N_4822);
nor U7428 (N_7428,N_5311,N_4151);
and U7429 (N_7429,N_4794,N_4027);
nand U7430 (N_7430,N_4503,N_5250);
nand U7431 (N_7431,N_5890,N_5108);
and U7432 (N_7432,N_5352,N_5627);
or U7433 (N_7433,N_4494,N_4883);
xnor U7434 (N_7434,N_4123,N_4606);
nor U7435 (N_7435,N_4226,N_4072);
or U7436 (N_7436,N_5829,N_5281);
and U7437 (N_7437,N_4521,N_4010);
and U7438 (N_7438,N_5403,N_5067);
or U7439 (N_7439,N_4409,N_4619);
nor U7440 (N_7440,N_4031,N_5934);
xnor U7441 (N_7441,N_4441,N_4937);
and U7442 (N_7442,N_4083,N_5644);
and U7443 (N_7443,N_5900,N_4505);
xnor U7444 (N_7444,N_4383,N_5623);
or U7445 (N_7445,N_4485,N_4542);
or U7446 (N_7446,N_5987,N_5626);
and U7447 (N_7447,N_4104,N_4313);
nand U7448 (N_7448,N_5358,N_4312);
and U7449 (N_7449,N_5326,N_4535);
nor U7450 (N_7450,N_5535,N_5089);
nor U7451 (N_7451,N_4250,N_5940);
or U7452 (N_7452,N_4951,N_4436);
nor U7453 (N_7453,N_4992,N_5393);
or U7454 (N_7454,N_5391,N_5099);
nand U7455 (N_7455,N_5421,N_5766);
nor U7456 (N_7456,N_4683,N_4736);
nor U7457 (N_7457,N_4672,N_5392);
xor U7458 (N_7458,N_5074,N_5059);
nand U7459 (N_7459,N_5427,N_4820);
nand U7460 (N_7460,N_5721,N_5709);
nor U7461 (N_7461,N_5660,N_4060);
nor U7462 (N_7462,N_5889,N_5972);
or U7463 (N_7463,N_4906,N_4263);
or U7464 (N_7464,N_4015,N_4847);
and U7465 (N_7465,N_4634,N_4797);
nor U7466 (N_7466,N_4739,N_5705);
nand U7467 (N_7467,N_4296,N_5660);
nand U7468 (N_7468,N_4489,N_4126);
nand U7469 (N_7469,N_5407,N_5260);
and U7470 (N_7470,N_4926,N_5397);
or U7471 (N_7471,N_5117,N_4374);
xnor U7472 (N_7472,N_4575,N_5008);
or U7473 (N_7473,N_4439,N_4660);
nor U7474 (N_7474,N_4834,N_4510);
or U7475 (N_7475,N_5705,N_4396);
or U7476 (N_7476,N_5656,N_4368);
nor U7477 (N_7477,N_5772,N_4950);
nor U7478 (N_7478,N_5212,N_4434);
and U7479 (N_7479,N_4148,N_5153);
nor U7480 (N_7480,N_4019,N_5342);
and U7481 (N_7481,N_4984,N_5684);
or U7482 (N_7482,N_5822,N_5559);
nand U7483 (N_7483,N_4293,N_5869);
xor U7484 (N_7484,N_4328,N_4384);
and U7485 (N_7485,N_4007,N_5945);
or U7486 (N_7486,N_4809,N_5391);
or U7487 (N_7487,N_4794,N_5062);
xor U7488 (N_7488,N_4179,N_4959);
nor U7489 (N_7489,N_5742,N_5323);
nand U7490 (N_7490,N_4141,N_4962);
or U7491 (N_7491,N_4104,N_4731);
nand U7492 (N_7492,N_5258,N_4887);
or U7493 (N_7493,N_5085,N_5853);
and U7494 (N_7494,N_5371,N_5265);
nand U7495 (N_7495,N_5471,N_5032);
or U7496 (N_7496,N_4780,N_4927);
or U7497 (N_7497,N_5921,N_5203);
nand U7498 (N_7498,N_5901,N_4603);
xor U7499 (N_7499,N_5844,N_5041);
nand U7500 (N_7500,N_5385,N_4131);
nand U7501 (N_7501,N_4148,N_5150);
xor U7502 (N_7502,N_4158,N_5150);
nand U7503 (N_7503,N_4442,N_5107);
or U7504 (N_7504,N_4524,N_5455);
and U7505 (N_7505,N_4086,N_4245);
or U7506 (N_7506,N_4316,N_4437);
nand U7507 (N_7507,N_4772,N_4791);
and U7508 (N_7508,N_4838,N_5022);
nand U7509 (N_7509,N_4501,N_5994);
or U7510 (N_7510,N_5041,N_5032);
nor U7511 (N_7511,N_4207,N_4257);
or U7512 (N_7512,N_5972,N_5826);
nor U7513 (N_7513,N_4228,N_5685);
nand U7514 (N_7514,N_5970,N_4585);
and U7515 (N_7515,N_5650,N_4119);
or U7516 (N_7516,N_4045,N_5667);
and U7517 (N_7517,N_5073,N_5116);
or U7518 (N_7518,N_4419,N_4205);
nor U7519 (N_7519,N_4762,N_4280);
xnor U7520 (N_7520,N_5822,N_5403);
nor U7521 (N_7521,N_5984,N_5775);
nand U7522 (N_7522,N_5717,N_5188);
xor U7523 (N_7523,N_4674,N_5531);
and U7524 (N_7524,N_5724,N_4691);
nand U7525 (N_7525,N_5333,N_5117);
and U7526 (N_7526,N_5115,N_5698);
or U7527 (N_7527,N_4381,N_4169);
and U7528 (N_7528,N_5201,N_4570);
nor U7529 (N_7529,N_4941,N_5267);
nor U7530 (N_7530,N_5789,N_4479);
nand U7531 (N_7531,N_4416,N_5323);
nor U7532 (N_7532,N_5471,N_5496);
xor U7533 (N_7533,N_5437,N_4788);
nor U7534 (N_7534,N_5522,N_4513);
nor U7535 (N_7535,N_5592,N_4639);
nor U7536 (N_7536,N_5771,N_5859);
nor U7537 (N_7537,N_4294,N_4607);
xnor U7538 (N_7538,N_4403,N_5104);
nand U7539 (N_7539,N_5246,N_4327);
nand U7540 (N_7540,N_5537,N_4031);
and U7541 (N_7541,N_5411,N_5086);
xnor U7542 (N_7542,N_5791,N_4365);
or U7543 (N_7543,N_4983,N_5077);
and U7544 (N_7544,N_4227,N_5347);
nor U7545 (N_7545,N_4738,N_4097);
and U7546 (N_7546,N_4338,N_4105);
and U7547 (N_7547,N_5847,N_5810);
and U7548 (N_7548,N_4776,N_4382);
and U7549 (N_7549,N_5047,N_4270);
and U7550 (N_7550,N_5421,N_5164);
xnor U7551 (N_7551,N_4788,N_4096);
or U7552 (N_7552,N_4975,N_4928);
or U7553 (N_7553,N_5448,N_4744);
or U7554 (N_7554,N_5687,N_5139);
nand U7555 (N_7555,N_4645,N_4109);
nor U7556 (N_7556,N_5854,N_5228);
and U7557 (N_7557,N_4479,N_5643);
or U7558 (N_7558,N_5717,N_5467);
and U7559 (N_7559,N_5804,N_5856);
and U7560 (N_7560,N_5163,N_4737);
and U7561 (N_7561,N_5713,N_5409);
xnor U7562 (N_7562,N_5700,N_5217);
nand U7563 (N_7563,N_4975,N_4711);
and U7564 (N_7564,N_4238,N_4126);
xor U7565 (N_7565,N_5568,N_4801);
and U7566 (N_7566,N_5894,N_5152);
and U7567 (N_7567,N_4457,N_5767);
xnor U7568 (N_7568,N_5343,N_4215);
nand U7569 (N_7569,N_4141,N_4270);
and U7570 (N_7570,N_5807,N_4551);
or U7571 (N_7571,N_5532,N_5052);
and U7572 (N_7572,N_5845,N_5912);
nand U7573 (N_7573,N_5512,N_5446);
nor U7574 (N_7574,N_4541,N_4885);
nand U7575 (N_7575,N_5314,N_4147);
and U7576 (N_7576,N_4854,N_4137);
nor U7577 (N_7577,N_4113,N_5834);
or U7578 (N_7578,N_5009,N_4596);
or U7579 (N_7579,N_4964,N_4868);
or U7580 (N_7580,N_5389,N_5792);
nor U7581 (N_7581,N_4501,N_4560);
nor U7582 (N_7582,N_4125,N_5026);
and U7583 (N_7583,N_4559,N_5056);
and U7584 (N_7584,N_5046,N_4358);
or U7585 (N_7585,N_5830,N_4891);
xor U7586 (N_7586,N_4714,N_4094);
nor U7587 (N_7587,N_4072,N_4099);
nand U7588 (N_7588,N_5794,N_4766);
nand U7589 (N_7589,N_5089,N_4143);
and U7590 (N_7590,N_4268,N_5547);
nor U7591 (N_7591,N_4155,N_4284);
or U7592 (N_7592,N_4634,N_4840);
or U7593 (N_7593,N_5599,N_5927);
nor U7594 (N_7594,N_5255,N_4747);
and U7595 (N_7595,N_5490,N_4882);
or U7596 (N_7596,N_5305,N_5207);
nand U7597 (N_7597,N_4799,N_4406);
or U7598 (N_7598,N_4374,N_5588);
and U7599 (N_7599,N_5338,N_5624);
nor U7600 (N_7600,N_4460,N_4889);
nor U7601 (N_7601,N_4221,N_5683);
nand U7602 (N_7602,N_5034,N_4805);
nand U7603 (N_7603,N_5677,N_4949);
nor U7604 (N_7604,N_5373,N_4390);
or U7605 (N_7605,N_4560,N_5130);
or U7606 (N_7606,N_5443,N_4390);
nor U7607 (N_7607,N_4878,N_5395);
and U7608 (N_7608,N_4219,N_4335);
nand U7609 (N_7609,N_4247,N_5648);
nand U7610 (N_7610,N_4047,N_5652);
or U7611 (N_7611,N_5149,N_5315);
nand U7612 (N_7612,N_5234,N_4747);
and U7613 (N_7613,N_4936,N_4891);
nor U7614 (N_7614,N_5741,N_4926);
and U7615 (N_7615,N_4562,N_5223);
xor U7616 (N_7616,N_4542,N_5506);
or U7617 (N_7617,N_4745,N_4718);
nand U7618 (N_7618,N_5700,N_5932);
and U7619 (N_7619,N_4356,N_4581);
nor U7620 (N_7620,N_4064,N_4968);
or U7621 (N_7621,N_4593,N_5256);
nand U7622 (N_7622,N_4490,N_5277);
nor U7623 (N_7623,N_5143,N_5877);
nor U7624 (N_7624,N_4184,N_4488);
xnor U7625 (N_7625,N_5338,N_5253);
and U7626 (N_7626,N_4133,N_4794);
and U7627 (N_7627,N_5302,N_5473);
nor U7628 (N_7628,N_4142,N_4751);
or U7629 (N_7629,N_5453,N_4668);
xnor U7630 (N_7630,N_5341,N_4310);
xnor U7631 (N_7631,N_4780,N_4160);
nand U7632 (N_7632,N_5940,N_5504);
nor U7633 (N_7633,N_4313,N_4342);
nor U7634 (N_7634,N_5653,N_4408);
and U7635 (N_7635,N_5106,N_4818);
and U7636 (N_7636,N_4522,N_4807);
or U7637 (N_7637,N_5353,N_4189);
nand U7638 (N_7638,N_5667,N_5292);
or U7639 (N_7639,N_5793,N_4540);
or U7640 (N_7640,N_4750,N_4968);
nor U7641 (N_7641,N_5615,N_5556);
xnor U7642 (N_7642,N_4593,N_5090);
nand U7643 (N_7643,N_5491,N_4014);
nor U7644 (N_7644,N_4503,N_4596);
or U7645 (N_7645,N_5377,N_4216);
xor U7646 (N_7646,N_4499,N_5977);
xnor U7647 (N_7647,N_4337,N_5068);
nand U7648 (N_7648,N_4872,N_5739);
or U7649 (N_7649,N_5568,N_5106);
nor U7650 (N_7650,N_5328,N_4188);
nand U7651 (N_7651,N_4024,N_5690);
nand U7652 (N_7652,N_4759,N_5952);
xor U7653 (N_7653,N_5496,N_4592);
and U7654 (N_7654,N_5674,N_4196);
or U7655 (N_7655,N_4244,N_4520);
or U7656 (N_7656,N_4648,N_4340);
or U7657 (N_7657,N_5961,N_4220);
nand U7658 (N_7658,N_5238,N_4080);
or U7659 (N_7659,N_5015,N_5894);
and U7660 (N_7660,N_4402,N_4611);
nor U7661 (N_7661,N_5864,N_5529);
and U7662 (N_7662,N_5601,N_4834);
xor U7663 (N_7663,N_5067,N_4331);
or U7664 (N_7664,N_5204,N_4420);
nand U7665 (N_7665,N_5502,N_4645);
or U7666 (N_7666,N_4280,N_5241);
nand U7667 (N_7667,N_4419,N_4644);
nand U7668 (N_7668,N_5238,N_4390);
nor U7669 (N_7669,N_5527,N_4259);
nor U7670 (N_7670,N_4691,N_5711);
and U7671 (N_7671,N_4433,N_5164);
nor U7672 (N_7672,N_4760,N_5449);
or U7673 (N_7673,N_4395,N_4816);
xnor U7674 (N_7674,N_4281,N_4469);
nor U7675 (N_7675,N_5277,N_4747);
nor U7676 (N_7676,N_4932,N_5305);
nand U7677 (N_7677,N_4423,N_5319);
or U7678 (N_7678,N_5939,N_5502);
and U7679 (N_7679,N_4563,N_4465);
or U7680 (N_7680,N_4416,N_4438);
nand U7681 (N_7681,N_4116,N_5964);
nor U7682 (N_7682,N_5192,N_4022);
and U7683 (N_7683,N_4318,N_5987);
nand U7684 (N_7684,N_4037,N_4882);
xor U7685 (N_7685,N_4284,N_5269);
nand U7686 (N_7686,N_4501,N_4177);
and U7687 (N_7687,N_4101,N_4016);
and U7688 (N_7688,N_4532,N_4275);
nor U7689 (N_7689,N_4144,N_4936);
and U7690 (N_7690,N_4125,N_5313);
or U7691 (N_7691,N_5923,N_4973);
nand U7692 (N_7692,N_4303,N_4188);
nor U7693 (N_7693,N_4629,N_4513);
and U7694 (N_7694,N_5146,N_5846);
xnor U7695 (N_7695,N_5597,N_4971);
nor U7696 (N_7696,N_5829,N_5483);
nand U7697 (N_7697,N_4543,N_5970);
and U7698 (N_7698,N_4919,N_5521);
and U7699 (N_7699,N_4166,N_4127);
nor U7700 (N_7700,N_5899,N_5670);
or U7701 (N_7701,N_5709,N_4413);
or U7702 (N_7702,N_5207,N_4875);
or U7703 (N_7703,N_4605,N_4544);
nor U7704 (N_7704,N_4277,N_4411);
xnor U7705 (N_7705,N_4990,N_5019);
nor U7706 (N_7706,N_5932,N_5835);
and U7707 (N_7707,N_5735,N_4342);
nor U7708 (N_7708,N_5991,N_4984);
and U7709 (N_7709,N_4124,N_5580);
or U7710 (N_7710,N_4417,N_5708);
or U7711 (N_7711,N_5379,N_4458);
and U7712 (N_7712,N_4387,N_4240);
and U7713 (N_7713,N_5828,N_5491);
or U7714 (N_7714,N_4345,N_4473);
and U7715 (N_7715,N_4293,N_4423);
nand U7716 (N_7716,N_5457,N_4971);
and U7717 (N_7717,N_5893,N_4778);
nor U7718 (N_7718,N_4592,N_4557);
nand U7719 (N_7719,N_4783,N_5156);
nand U7720 (N_7720,N_4559,N_5442);
nand U7721 (N_7721,N_4649,N_4278);
xnor U7722 (N_7722,N_4415,N_5419);
or U7723 (N_7723,N_5909,N_5603);
and U7724 (N_7724,N_5969,N_4626);
and U7725 (N_7725,N_4513,N_4693);
and U7726 (N_7726,N_5743,N_4521);
xor U7727 (N_7727,N_4276,N_4094);
and U7728 (N_7728,N_5433,N_4235);
nor U7729 (N_7729,N_4125,N_5042);
nor U7730 (N_7730,N_4913,N_5712);
and U7731 (N_7731,N_4700,N_4896);
nor U7732 (N_7732,N_5369,N_5358);
or U7733 (N_7733,N_5736,N_4407);
xor U7734 (N_7734,N_4264,N_5640);
nor U7735 (N_7735,N_4276,N_4619);
and U7736 (N_7736,N_5468,N_5771);
and U7737 (N_7737,N_4046,N_5196);
and U7738 (N_7738,N_5301,N_4388);
or U7739 (N_7739,N_4176,N_5370);
nor U7740 (N_7740,N_4468,N_5733);
nand U7741 (N_7741,N_5993,N_4878);
xor U7742 (N_7742,N_4511,N_5839);
and U7743 (N_7743,N_5758,N_5066);
and U7744 (N_7744,N_5619,N_5735);
nor U7745 (N_7745,N_4280,N_4907);
xnor U7746 (N_7746,N_4865,N_4142);
nand U7747 (N_7747,N_5303,N_4993);
and U7748 (N_7748,N_4127,N_5179);
or U7749 (N_7749,N_4733,N_5361);
or U7750 (N_7750,N_5800,N_4852);
and U7751 (N_7751,N_4338,N_4284);
nand U7752 (N_7752,N_5357,N_4544);
xnor U7753 (N_7753,N_5360,N_4165);
nor U7754 (N_7754,N_5294,N_5541);
and U7755 (N_7755,N_4232,N_5583);
xor U7756 (N_7756,N_5152,N_4683);
xor U7757 (N_7757,N_4238,N_4343);
nand U7758 (N_7758,N_4887,N_5536);
or U7759 (N_7759,N_5030,N_5500);
nand U7760 (N_7760,N_4967,N_5056);
xor U7761 (N_7761,N_4948,N_4991);
nor U7762 (N_7762,N_4354,N_4025);
nor U7763 (N_7763,N_5867,N_4434);
nor U7764 (N_7764,N_4416,N_5852);
nor U7765 (N_7765,N_5224,N_5168);
nor U7766 (N_7766,N_5940,N_4300);
nand U7767 (N_7767,N_5477,N_4213);
nor U7768 (N_7768,N_4146,N_4731);
xnor U7769 (N_7769,N_5842,N_4845);
nor U7770 (N_7770,N_5679,N_5647);
and U7771 (N_7771,N_4346,N_5560);
nor U7772 (N_7772,N_5134,N_5815);
nand U7773 (N_7773,N_4038,N_4495);
nor U7774 (N_7774,N_4562,N_5899);
nor U7775 (N_7775,N_4055,N_4777);
and U7776 (N_7776,N_5231,N_5707);
and U7777 (N_7777,N_4733,N_4595);
or U7778 (N_7778,N_5188,N_4868);
or U7779 (N_7779,N_4459,N_5556);
and U7780 (N_7780,N_4750,N_4054);
and U7781 (N_7781,N_5653,N_4601);
or U7782 (N_7782,N_4884,N_5795);
and U7783 (N_7783,N_4830,N_4334);
or U7784 (N_7784,N_4940,N_4065);
xor U7785 (N_7785,N_4971,N_5426);
nand U7786 (N_7786,N_4949,N_4506);
or U7787 (N_7787,N_5201,N_4109);
nor U7788 (N_7788,N_4851,N_4017);
nor U7789 (N_7789,N_4293,N_5149);
nand U7790 (N_7790,N_5310,N_5935);
or U7791 (N_7791,N_4945,N_4771);
nor U7792 (N_7792,N_4247,N_5352);
nor U7793 (N_7793,N_4605,N_4402);
xnor U7794 (N_7794,N_4166,N_4301);
nor U7795 (N_7795,N_4673,N_5520);
or U7796 (N_7796,N_4816,N_4997);
nand U7797 (N_7797,N_5690,N_5113);
or U7798 (N_7798,N_4540,N_4937);
nor U7799 (N_7799,N_5007,N_5549);
xor U7800 (N_7800,N_5971,N_5744);
and U7801 (N_7801,N_5861,N_5645);
or U7802 (N_7802,N_4715,N_5074);
nand U7803 (N_7803,N_4151,N_5438);
nor U7804 (N_7804,N_4777,N_5236);
nand U7805 (N_7805,N_5433,N_5474);
and U7806 (N_7806,N_5950,N_5426);
or U7807 (N_7807,N_5299,N_5121);
xnor U7808 (N_7808,N_4500,N_5252);
and U7809 (N_7809,N_5946,N_4116);
or U7810 (N_7810,N_4109,N_5129);
and U7811 (N_7811,N_4891,N_4844);
nand U7812 (N_7812,N_4143,N_4019);
nor U7813 (N_7813,N_5991,N_4387);
and U7814 (N_7814,N_5184,N_4584);
and U7815 (N_7815,N_5098,N_5294);
or U7816 (N_7816,N_4798,N_4870);
nand U7817 (N_7817,N_4552,N_5593);
nor U7818 (N_7818,N_4807,N_5544);
nand U7819 (N_7819,N_4049,N_4908);
or U7820 (N_7820,N_5567,N_5444);
xor U7821 (N_7821,N_5867,N_4442);
nand U7822 (N_7822,N_5763,N_4979);
and U7823 (N_7823,N_4479,N_5083);
or U7824 (N_7824,N_4403,N_5057);
nand U7825 (N_7825,N_5472,N_5221);
nor U7826 (N_7826,N_5452,N_5714);
nor U7827 (N_7827,N_5396,N_5590);
xnor U7828 (N_7828,N_4742,N_4588);
or U7829 (N_7829,N_4845,N_5759);
or U7830 (N_7830,N_4560,N_4508);
xor U7831 (N_7831,N_4916,N_4575);
and U7832 (N_7832,N_5543,N_4562);
and U7833 (N_7833,N_5312,N_5129);
xor U7834 (N_7834,N_5256,N_4469);
nor U7835 (N_7835,N_5385,N_5230);
or U7836 (N_7836,N_4516,N_5410);
nor U7837 (N_7837,N_4086,N_4065);
and U7838 (N_7838,N_4566,N_5223);
xor U7839 (N_7839,N_5435,N_5501);
or U7840 (N_7840,N_5314,N_4613);
nor U7841 (N_7841,N_4029,N_4285);
nand U7842 (N_7842,N_4889,N_5706);
xor U7843 (N_7843,N_4959,N_4183);
nor U7844 (N_7844,N_4033,N_5237);
nor U7845 (N_7845,N_4360,N_4760);
or U7846 (N_7846,N_4054,N_4963);
nand U7847 (N_7847,N_4197,N_5523);
and U7848 (N_7848,N_5463,N_5332);
nor U7849 (N_7849,N_5574,N_4096);
or U7850 (N_7850,N_4878,N_5430);
nand U7851 (N_7851,N_5070,N_5925);
or U7852 (N_7852,N_4086,N_5547);
and U7853 (N_7853,N_4662,N_5176);
or U7854 (N_7854,N_5660,N_4712);
or U7855 (N_7855,N_5939,N_5564);
nand U7856 (N_7856,N_4680,N_5985);
nor U7857 (N_7857,N_5620,N_4366);
nand U7858 (N_7858,N_5662,N_5332);
nor U7859 (N_7859,N_5837,N_4955);
and U7860 (N_7860,N_4731,N_5127);
nand U7861 (N_7861,N_5994,N_5053);
or U7862 (N_7862,N_5798,N_5544);
or U7863 (N_7863,N_4071,N_4409);
or U7864 (N_7864,N_4656,N_4596);
and U7865 (N_7865,N_4219,N_5926);
nor U7866 (N_7866,N_4251,N_4814);
xnor U7867 (N_7867,N_4754,N_5176);
nand U7868 (N_7868,N_4741,N_4779);
nand U7869 (N_7869,N_4057,N_4830);
nor U7870 (N_7870,N_5551,N_5064);
and U7871 (N_7871,N_4369,N_4604);
and U7872 (N_7872,N_5318,N_5974);
or U7873 (N_7873,N_4079,N_5971);
or U7874 (N_7874,N_5789,N_4188);
or U7875 (N_7875,N_5680,N_5693);
nor U7876 (N_7876,N_5788,N_4157);
or U7877 (N_7877,N_4582,N_5180);
nor U7878 (N_7878,N_5006,N_5926);
nand U7879 (N_7879,N_5255,N_4015);
nor U7880 (N_7880,N_5998,N_5817);
xor U7881 (N_7881,N_4033,N_5290);
and U7882 (N_7882,N_5790,N_4377);
xnor U7883 (N_7883,N_5338,N_4026);
nor U7884 (N_7884,N_4588,N_5158);
nor U7885 (N_7885,N_4631,N_4311);
nor U7886 (N_7886,N_4845,N_5987);
nand U7887 (N_7887,N_5416,N_4717);
nor U7888 (N_7888,N_5300,N_4769);
and U7889 (N_7889,N_4066,N_4987);
nor U7890 (N_7890,N_4581,N_4146);
and U7891 (N_7891,N_5366,N_5177);
nand U7892 (N_7892,N_5229,N_4843);
and U7893 (N_7893,N_5238,N_5065);
and U7894 (N_7894,N_5112,N_4948);
and U7895 (N_7895,N_5308,N_4775);
and U7896 (N_7896,N_4549,N_4198);
nand U7897 (N_7897,N_5715,N_4227);
nor U7898 (N_7898,N_5304,N_5964);
nor U7899 (N_7899,N_4902,N_5223);
nand U7900 (N_7900,N_4030,N_5977);
and U7901 (N_7901,N_5141,N_4394);
and U7902 (N_7902,N_4278,N_4322);
and U7903 (N_7903,N_4023,N_4306);
nor U7904 (N_7904,N_4431,N_5382);
xor U7905 (N_7905,N_5182,N_5160);
xnor U7906 (N_7906,N_4301,N_5029);
or U7907 (N_7907,N_4287,N_5861);
or U7908 (N_7908,N_5536,N_4423);
nor U7909 (N_7909,N_4812,N_5641);
nand U7910 (N_7910,N_5484,N_4728);
nand U7911 (N_7911,N_4267,N_5327);
nand U7912 (N_7912,N_4512,N_5449);
and U7913 (N_7913,N_4400,N_5201);
nor U7914 (N_7914,N_5845,N_5718);
nor U7915 (N_7915,N_5499,N_5793);
and U7916 (N_7916,N_4646,N_4197);
and U7917 (N_7917,N_5954,N_4375);
nand U7918 (N_7918,N_5852,N_5873);
nor U7919 (N_7919,N_4434,N_4915);
nor U7920 (N_7920,N_5302,N_4544);
nor U7921 (N_7921,N_5070,N_5598);
and U7922 (N_7922,N_5734,N_5869);
or U7923 (N_7923,N_4447,N_4196);
and U7924 (N_7924,N_5824,N_5068);
nor U7925 (N_7925,N_4435,N_4064);
nand U7926 (N_7926,N_5596,N_5415);
nand U7927 (N_7927,N_4884,N_5681);
nand U7928 (N_7928,N_5037,N_5060);
nor U7929 (N_7929,N_5955,N_5891);
nor U7930 (N_7930,N_5968,N_4781);
nor U7931 (N_7931,N_5176,N_4971);
and U7932 (N_7932,N_4130,N_5517);
nor U7933 (N_7933,N_4965,N_5399);
or U7934 (N_7934,N_4700,N_4766);
nand U7935 (N_7935,N_4376,N_5536);
and U7936 (N_7936,N_4118,N_5747);
or U7937 (N_7937,N_4287,N_5772);
and U7938 (N_7938,N_5190,N_5250);
and U7939 (N_7939,N_5003,N_4223);
and U7940 (N_7940,N_4658,N_5924);
or U7941 (N_7941,N_4482,N_5707);
or U7942 (N_7942,N_5794,N_4080);
and U7943 (N_7943,N_5310,N_5175);
or U7944 (N_7944,N_5855,N_5207);
nor U7945 (N_7945,N_5727,N_5455);
nor U7946 (N_7946,N_4991,N_5166);
and U7947 (N_7947,N_4091,N_5733);
nor U7948 (N_7948,N_5239,N_4913);
and U7949 (N_7949,N_4552,N_5463);
or U7950 (N_7950,N_5077,N_4410);
nor U7951 (N_7951,N_4864,N_4328);
and U7952 (N_7952,N_5030,N_5506);
or U7953 (N_7953,N_5660,N_5626);
or U7954 (N_7954,N_5894,N_5586);
nor U7955 (N_7955,N_4019,N_5888);
nor U7956 (N_7956,N_5696,N_5703);
nor U7957 (N_7957,N_5568,N_4653);
nor U7958 (N_7958,N_4312,N_4195);
nand U7959 (N_7959,N_4296,N_4398);
and U7960 (N_7960,N_4655,N_4175);
nor U7961 (N_7961,N_5009,N_5104);
xnor U7962 (N_7962,N_4740,N_5168);
and U7963 (N_7963,N_5681,N_5519);
nand U7964 (N_7964,N_5253,N_4611);
and U7965 (N_7965,N_5125,N_5831);
xnor U7966 (N_7966,N_4033,N_5175);
and U7967 (N_7967,N_5202,N_5949);
and U7968 (N_7968,N_5697,N_4679);
and U7969 (N_7969,N_5327,N_4116);
or U7970 (N_7970,N_4378,N_4227);
or U7971 (N_7971,N_4566,N_5020);
or U7972 (N_7972,N_4511,N_5679);
and U7973 (N_7973,N_5424,N_4595);
nor U7974 (N_7974,N_4400,N_4143);
or U7975 (N_7975,N_5507,N_4330);
and U7976 (N_7976,N_4576,N_5564);
nand U7977 (N_7977,N_5426,N_5063);
and U7978 (N_7978,N_4868,N_4131);
nand U7979 (N_7979,N_5974,N_5359);
or U7980 (N_7980,N_4057,N_4633);
nand U7981 (N_7981,N_5399,N_5381);
xnor U7982 (N_7982,N_5088,N_5505);
and U7983 (N_7983,N_4209,N_5897);
and U7984 (N_7984,N_4534,N_4855);
nand U7985 (N_7985,N_5761,N_5256);
xor U7986 (N_7986,N_5690,N_4044);
nand U7987 (N_7987,N_4899,N_4360);
and U7988 (N_7988,N_4777,N_4026);
nand U7989 (N_7989,N_4717,N_5343);
nor U7990 (N_7990,N_5567,N_4968);
and U7991 (N_7991,N_5394,N_5378);
nor U7992 (N_7992,N_4520,N_5613);
nor U7993 (N_7993,N_4182,N_4717);
xor U7994 (N_7994,N_5065,N_5601);
or U7995 (N_7995,N_4548,N_4570);
nand U7996 (N_7996,N_4804,N_5530);
or U7997 (N_7997,N_5692,N_4428);
or U7998 (N_7998,N_4156,N_4726);
or U7999 (N_7999,N_4032,N_4404);
nor U8000 (N_8000,N_6622,N_7257);
or U8001 (N_8001,N_6329,N_7941);
or U8002 (N_8002,N_6247,N_6645);
nor U8003 (N_8003,N_7213,N_6731);
xor U8004 (N_8004,N_7381,N_7463);
or U8005 (N_8005,N_6105,N_7285);
nand U8006 (N_8006,N_6558,N_6641);
nor U8007 (N_8007,N_6898,N_6519);
or U8008 (N_8008,N_7951,N_7805);
or U8009 (N_8009,N_6277,N_7290);
nand U8010 (N_8010,N_6617,N_6629);
xor U8011 (N_8011,N_6158,N_7289);
xor U8012 (N_8012,N_6015,N_7545);
nor U8013 (N_8013,N_6162,N_7137);
or U8014 (N_8014,N_6457,N_6516);
or U8015 (N_8015,N_7170,N_6737);
nand U8016 (N_8016,N_7271,N_7889);
nor U8017 (N_8017,N_6775,N_7883);
or U8018 (N_8018,N_6746,N_6436);
nor U8019 (N_8019,N_6304,N_6875);
or U8020 (N_8020,N_7756,N_6148);
and U8021 (N_8021,N_6963,N_6578);
or U8022 (N_8022,N_7808,N_7350);
nor U8023 (N_8023,N_6409,N_7383);
xor U8024 (N_8024,N_7864,N_7559);
and U8025 (N_8025,N_6610,N_6423);
nor U8026 (N_8026,N_6745,N_6143);
or U8027 (N_8027,N_7906,N_7283);
xor U8028 (N_8028,N_6121,N_7741);
nor U8029 (N_8029,N_7769,N_6561);
nor U8030 (N_8030,N_6029,N_7516);
or U8031 (N_8031,N_6230,N_7885);
or U8032 (N_8032,N_7175,N_6959);
nand U8033 (N_8033,N_7645,N_6747);
nand U8034 (N_8034,N_7960,N_6479);
nor U8035 (N_8035,N_6935,N_6063);
or U8036 (N_8036,N_7527,N_7354);
nand U8037 (N_8037,N_7682,N_7478);
nor U8038 (N_8038,N_7936,N_6192);
and U8039 (N_8039,N_7007,N_6376);
nand U8040 (N_8040,N_6068,N_7093);
nand U8041 (N_8041,N_7698,N_7127);
and U8042 (N_8042,N_7572,N_7501);
nor U8043 (N_8043,N_7031,N_7288);
xor U8044 (N_8044,N_7540,N_6686);
nor U8045 (N_8045,N_6569,N_7237);
xnor U8046 (N_8046,N_6153,N_7332);
nor U8047 (N_8047,N_6798,N_7449);
nor U8048 (N_8048,N_6260,N_7788);
nor U8049 (N_8049,N_7492,N_7468);
and U8050 (N_8050,N_7241,N_7707);
and U8051 (N_8051,N_7553,N_7217);
nor U8052 (N_8052,N_6718,N_7578);
nand U8053 (N_8053,N_7312,N_7893);
nand U8054 (N_8054,N_6083,N_7778);
or U8055 (N_8055,N_7600,N_6933);
nor U8056 (N_8056,N_6388,N_7313);
and U8057 (N_8057,N_6460,N_7438);
nor U8058 (N_8058,N_7777,N_7755);
nor U8059 (N_8059,N_7024,N_6420);
or U8060 (N_8060,N_6387,N_6998);
nand U8061 (N_8061,N_7366,N_7091);
xnor U8062 (N_8062,N_7046,N_7061);
and U8063 (N_8063,N_6874,N_6071);
and U8064 (N_8064,N_6663,N_6702);
and U8065 (N_8065,N_7124,N_6138);
nor U8066 (N_8066,N_6429,N_6188);
or U8067 (N_8067,N_7503,N_6621);
xnor U8068 (N_8068,N_7442,N_7882);
and U8069 (N_8069,N_6410,N_6253);
nor U8070 (N_8070,N_6413,N_7291);
nand U8071 (N_8071,N_7082,N_6434);
and U8072 (N_8072,N_6485,N_6730);
xor U8073 (N_8073,N_6675,N_7852);
nor U8074 (N_8074,N_7894,N_6943);
nor U8075 (N_8075,N_7557,N_6256);
or U8076 (N_8076,N_6832,N_7779);
xor U8077 (N_8077,N_6759,N_7845);
nand U8078 (N_8078,N_7868,N_7443);
nor U8079 (N_8079,N_6966,N_7909);
nor U8080 (N_8080,N_7421,N_7167);
xor U8081 (N_8081,N_6360,N_6992);
xnor U8082 (N_8082,N_7734,N_6833);
and U8083 (N_8083,N_7027,N_7075);
nor U8084 (N_8084,N_7049,N_7981);
nor U8085 (N_8085,N_6958,N_7692);
xor U8086 (N_8086,N_6886,N_6067);
or U8087 (N_8087,N_7884,N_6508);
nor U8088 (N_8088,N_6160,N_7179);
xnor U8089 (N_8089,N_7196,N_7956);
nand U8090 (N_8090,N_7865,N_7431);
and U8091 (N_8091,N_6164,N_6892);
nand U8092 (N_8092,N_6052,N_6899);
nand U8093 (N_8093,N_6931,N_6156);
and U8094 (N_8094,N_7481,N_7387);
and U8095 (N_8095,N_7668,N_7611);
nand U8096 (N_8096,N_6647,N_6528);
nor U8097 (N_8097,N_6704,N_7327);
xnor U8098 (N_8098,N_6901,N_6733);
nand U8099 (N_8099,N_7300,N_7739);
nand U8100 (N_8100,N_7025,N_6688);
or U8101 (N_8101,N_6118,N_6132);
and U8102 (N_8102,N_6628,N_7942);
and U8103 (N_8103,N_7700,N_6181);
xnor U8104 (N_8104,N_7092,N_6169);
and U8105 (N_8105,N_7591,N_7689);
nor U8106 (N_8106,N_6155,N_7362);
or U8107 (N_8107,N_6591,N_6112);
nor U8108 (N_8108,N_7613,N_7825);
nand U8109 (N_8109,N_6221,N_7059);
or U8110 (N_8110,N_6368,N_7719);
or U8111 (N_8111,N_6492,N_6634);
nand U8112 (N_8112,N_6228,N_7360);
or U8113 (N_8113,N_6397,N_6748);
xor U8114 (N_8114,N_7671,N_6094);
or U8115 (N_8115,N_6810,N_7999);
and U8116 (N_8116,N_6279,N_6381);
nor U8117 (N_8117,N_6019,N_7497);
or U8118 (N_8118,N_7604,N_6128);
xor U8119 (N_8119,N_7185,N_7108);
or U8120 (N_8120,N_7309,N_7514);
and U8121 (N_8121,N_6785,N_6713);
and U8122 (N_8122,N_6418,N_7801);
or U8123 (N_8123,N_6537,N_7699);
or U8124 (N_8124,N_6865,N_6678);
nand U8125 (N_8125,N_7240,N_6697);
nand U8126 (N_8126,N_7452,N_7265);
nor U8127 (N_8127,N_6517,N_7489);
nor U8128 (N_8128,N_7983,N_7966);
nor U8129 (N_8129,N_7714,N_6183);
and U8130 (N_8130,N_6559,N_6292);
nand U8131 (N_8131,N_6720,N_7561);
nand U8132 (N_8132,N_7132,N_6571);
or U8133 (N_8133,N_7948,N_7551);
or U8134 (N_8134,N_7916,N_7279);
or U8135 (N_8135,N_7802,N_7673);
or U8136 (N_8136,N_7261,N_7294);
and U8137 (N_8137,N_7416,N_7361);
or U8138 (N_8138,N_6373,N_7054);
xnor U8139 (N_8139,N_7567,N_6380);
xnor U8140 (N_8140,N_6443,N_7826);
nand U8141 (N_8141,N_6592,N_7270);
nand U8142 (N_8142,N_7832,N_6284);
nor U8143 (N_8143,N_7615,N_7413);
nor U8144 (N_8144,N_6724,N_6606);
or U8145 (N_8145,N_6484,N_6268);
and U8146 (N_8146,N_7052,N_6917);
nand U8147 (N_8147,N_7114,N_6608);
or U8148 (N_8148,N_7694,N_6983);
or U8149 (N_8149,N_6753,N_6538);
nand U8150 (N_8150,N_6077,N_6696);
and U8151 (N_8151,N_6315,N_7686);
or U8152 (N_8152,N_7032,N_7774);
or U8153 (N_8153,N_6140,N_6843);
nor U8154 (N_8154,N_7809,N_6407);
or U8155 (N_8155,N_6198,N_7333);
nor U8156 (N_8156,N_6842,N_6987);
nor U8157 (N_8157,N_6612,N_6776);
nor U8158 (N_8158,N_6633,N_7365);
xnor U8159 (N_8159,N_7976,N_7400);
or U8160 (N_8160,N_6563,N_7136);
or U8161 (N_8161,N_6022,N_7767);
and U8162 (N_8162,N_7187,N_7219);
and U8163 (N_8163,N_7281,N_7772);
and U8164 (N_8164,N_6271,N_6431);
or U8165 (N_8165,N_7152,N_6588);
or U8166 (N_8166,N_7697,N_7520);
nand U8167 (N_8167,N_6964,N_6246);
nand U8168 (N_8168,N_7395,N_7401);
and U8169 (N_8169,N_7038,N_7235);
nor U8170 (N_8170,N_6200,N_6672);
nand U8171 (N_8171,N_6073,N_6337);
nor U8172 (N_8172,N_6406,N_6482);
or U8173 (N_8173,N_6799,N_6805);
or U8174 (N_8174,N_6650,N_7162);
nand U8175 (N_8175,N_6088,N_7207);
nor U8176 (N_8176,N_7888,N_7822);
or U8177 (N_8177,N_7377,N_7113);
nand U8178 (N_8178,N_7510,N_6047);
or U8179 (N_8179,N_6031,N_6459);
nand U8180 (N_8180,N_6415,N_6456);
nand U8181 (N_8181,N_7280,N_6590);
and U8182 (N_8182,N_7840,N_7066);
nor U8183 (N_8183,N_6623,N_6475);
or U8184 (N_8184,N_6448,N_7353);
nand U8185 (N_8185,N_7846,N_7924);
or U8186 (N_8186,N_7085,N_6007);
and U8187 (N_8187,N_7139,N_6709);
and U8188 (N_8188,N_7913,N_7277);
nor U8189 (N_8189,N_6102,N_7780);
nand U8190 (N_8190,N_6814,N_6554);
and U8191 (N_8191,N_7873,N_7009);
xnor U8192 (N_8192,N_7608,N_6905);
and U8193 (N_8193,N_7256,N_6995);
or U8194 (N_8194,N_6723,N_7222);
xor U8195 (N_8195,N_6002,N_7517);
and U8196 (N_8196,N_7628,N_7760);
and U8197 (N_8197,N_6868,N_6703);
nand U8198 (N_8198,N_6914,N_7640);
nor U8199 (N_8199,N_6012,N_6120);
or U8200 (N_8200,N_7445,N_7509);
or U8201 (N_8201,N_6970,N_7212);
nand U8202 (N_8202,N_6965,N_6564);
and U8203 (N_8203,N_6061,N_6861);
and U8204 (N_8204,N_7538,N_6172);
and U8205 (N_8205,N_6908,N_6699);
or U8206 (N_8206,N_6152,N_6374);
nor U8207 (N_8207,N_7555,N_6248);
nor U8208 (N_8208,N_7813,N_6116);
nor U8209 (N_8209,N_6862,N_6098);
and U8210 (N_8210,N_7258,N_6003);
or U8211 (N_8211,N_7063,N_6942);
nor U8212 (N_8212,N_6550,N_7268);
nand U8213 (N_8213,N_7065,N_7472);
and U8214 (N_8214,N_7775,N_6514);
and U8215 (N_8215,N_6472,N_6594);
xnor U8216 (N_8216,N_7744,N_7047);
and U8217 (N_8217,N_7070,N_6209);
nor U8218 (N_8218,N_7975,N_6744);
nand U8219 (N_8219,N_7317,N_7566);
nand U8220 (N_8220,N_6949,N_7570);
nand U8221 (N_8221,N_6401,N_6189);
and U8222 (N_8222,N_6669,N_6946);
nand U8223 (N_8223,N_6827,N_7800);
and U8224 (N_8224,N_7087,N_6982);
nor U8225 (N_8225,N_7874,N_6218);
nor U8226 (N_8226,N_6668,N_7922);
or U8227 (N_8227,N_6481,N_6090);
nor U8228 (N_8228,N_6227,N_6812);
or U8229 (N_8229,N_6813,N_6280);
xnor U8230 (N_8230,N_7980,N_6796);
nand U8231 (N_8231,N_7135,N_7156);
or U8232 (N_8232,N_7457,N_7161);
nor U8233 (N_8233,N_7879,N_6929);
nand U8234 (N_8234,N_7512,N_7984);
nor U8235 (N_8235,N_6828,N_7701);
nor U8236 (N_8236,N_6202,N_6422);
nand U8237 (N_8237,N_7434,N_6527);
or U8238 (N_8238,N_7143,N_7482);
and U8239 (N_8239,N_6039,N_6870);
and U8240 (N_8240,N_6952,N_6362);
or U8241 (N_8241,N_7598,N_7266);
nor U8242 (N_8242,N_7634,N_6382);
or U8243 (N_8243,N_7005,N_6640);
and U8244 (N_8244,N_7839,N_6427);
or U8245 (N_8245,N_6589,N_6043);
nor U8246 (N_8246,N_6794,N_6978);
nor U8247 (N_8247,N_7378,N_7318);
nand U8248 (N_8248,N_7392,N_6627);
nand U8249 (N_8249,N_7471,N_7056);
nor U8250 (N_8250,N_6040,N_7432);
nor U8251 (N_8251,N_6220,N_6895);
nor U8252 (N_8252,N_6788,N_6237);
xnor U8253 (N_8253,N_7015,N_7552);
and U8254 (N_8254,N_7796,N_6275);
and U8255 (N_8255,N_7238,N_6834);
or U8256 (N_8256,N_6920,N_6203);
xor U8257 (N_8257,N_6867,N_6593);
nand U8258 (N_8258,N_7646,N_7977);
nor U8259 (N_8259,N_6676,N_7982);
nand U8260 (N_8260,N_6654,N_6215);
nand U8261 (N_8261,N_6317,N_7584);
nor U8262 (N_8262,N_6473,N_7513);
nor U8263 (N_8263,N_7034,N_7019);
nand U8264 (N_8264,N_7745,N_7624);
and U8265 (N_8265,N_7842,N_7123);
and U8266 (N_8266,N_7626,N_7414);
nor U8267 (N_8267,N_7855,N_6293);
nand U8268 (N_8268,N_6149,N_7738);
nor U8269 (N_8269,N_7496,N_6956);
nor U8270 (N_8270,N_7733,N_7642);
nand U8271 (N_8271,N_6057,N_6370);
or U8272 (N_8272,N_7729,N_6586);
and U8273 (N_8273,N_7299,N_7287);
nand U8274 (N_8274,N_6013,N_7577);
and U8275 (N_8275,N_7144,N_6618);
xnor U8276 (N_8276,N_6909,N_6758);
and U8277 (N_8277,N_6426,N_7264);
and U8278 (N_8278,N_7486,N_6267);
nand U8279 (N_8279,N_6766,N_6656);
or U8280 (N_8280,N_7666,N_6255);
nand U8281 (N_8281,N_7035,N_6016);
nand U8282 (N_8282,N_6087,N_6453);
nand U8283 (N_8283,N_6692,N_7410);
nor U8284 (N_8284,N_7554,N_6408);
and U8285 (N_8285,N_7939,N_7971);
nor U8286 (N_8286,N_6769,N_7120);
or U8287 (N_8287,N_6881,N_7662);
or U8288 (N_8288,N_6351,N_6433);
nand U8289 (N_8289,N_6273,N_6525);
nor U8290 (N_8290,N_7500,N_6032);
nand U8291 (N_8291,N_7823,N_7781);
and U8292 (N_8292,N_7249,N_6953);
nor U8293 (N_8293,N_7098,N_6869);
and U8294 (N_8294,N_6760,N_7549);
and U8295 (N_8295,N_7349,N_7459);
nand U8296 (N_8296,N_6683,N_6464);
nor U8297 (N_8297,N_7302,N_7759);
nand U8298 (N_8298,N_6046,N_6290);
or U8299 (N_8299,N_7742,N_6653);
nor U8300 (N_8300,N_6305,N_7441);
and U8301 (N_8301,N_7403,N_6841);
or U8302 (N_8302,N_7961,N_7848);
or U8303 (N_8303,N_7892,N_6597);
nand U8304 (N_8304,N_7534,N_7798);
and U8305 (N_8305,N_6824,N_7819);
nand U8306 (N_8306,N_6659,N_7053);
xnor U8307 (N_8307,N_7141,N_7940);
nand U8308 (N_8308,N_6549,N_7532);
nor U8309 (N_8309,N_6941,N_6918);
xor U8310 (N_8310,N_7691,N_6207);
or U8311 (N_8311,N_6424,N_7100);
nor U8312 (N_8312,N_7344,N_6086);
nor U8313 (N_8313,N_7131,N_6555);
nor U8314 (N_8314,N_7528,N_7743);
nor U8315 (N_8315,N_6662,N_6880);
or U8316 (N_8316,N_7575,N_6690);
and U8317 (N_8317,N_7347,N_7329);
nand U8318 (N_8318,N_7307,N_6925);
nor U8319 (N_8319,N_7150,N_7195);
or U8320 (N_8320,N_6263,N_7747);
and U8321 (N_8321,N_6165,N_6295);
or U8322 (N_8322,N_7670,N_7979);
nand U8323 (N_8323,N_6969,N_7877);
and U8324 (N_8324,N_6800,N_7126);
or U8325 (N_8325,N_7905,N_6445);
nand U8326 (N_8326,N_6212,N_6756);
nor U8327 (N_8327,N_6521,N_6385);
nor U8328 (N_8328,N_6818,N_7296);
or U8329 (N_8329,N_7424,N_7345);
nor U8330 (N_8330,N_6716,N_6535);
and U8331 (N_8331,N_7706,N_6008);
nand U8332 (N_8332,N_6896,N_6893);
nand U8333 (N_8333,N_7386,N_7314);
and U8334 (N_8334,N_7089,N_6529);
or U8335 (N_8335,N_7428,N_7274);
nand U8336 (N_8336,N_6361,N_7346);
nand U8337 (N_8337,N_6291,N_6544);
nand U8338 (N_8338,N_6620,N_6166);
and U8339 (N_8339,N_6494,N_6695);
xor U8340 (N_8340,N_6298,N_7669);
and U8341 (N_8341,N_6286,N_7556);
xor U8342 (N_8342,N_7751,N_7495);
nor U8343 (N_8343,N_7576,N_6444);
and U8344 (N_8344,N_6625,N_6021);
nor U8345 (N_8345,N_7076,N_6652);
and U8346 (N_8346,N_7933,N_7518);
or U8347 (N_8347,N_6534,N_6577);
nor U8348 (N_8348,N_7827,N_7638);
and U8349 (N_8349,N_6504,N_6301);
or U8350 (N_8350,N_6178,N_7602);
nor U8351 (N_8351,N_7519,N_6369);
and U8352 (N_8352,N_7835,N_7859);
nand U8353 (N_8353,N_7710,N_7614);
and U8354 (N_8354,N_6630,N_7996);
and U8355 (N_8355,N_6782,N_7476);
nor U8356 (N_8356,N_6774,N_7316);
xor U8357 (N_8357,N_6447,N_6226);
nor U8358 (N_8358,N_6352,N_7014);
xor U8359 (N_8359,N_6646,N_6225);
nor U8360 (N_8360,N_7658,N_6092);
and U8361 (N_8361,N_7321,N_6829);
nand U8362 (N_8362,N_7048,N_7456);
nor U8363 (N_8363,N_6334,N_7521);
and U8364 (N_8364,N_6499,N_7887);
nand U8365 (N_8365,N_6503,N_7599);
nor U8366 (N_8366,N_7943,N_6732);
and U8367 (N_8367,N_6014,N_6217);
or U8368 (N_8368,N_6242,N_6483);
nor U8369 (N_8369,N_6511,N_7677);
nor U8370 (N_8370,N_6144,N_6546);
and U8371 (N_8371,N_6379,N_7904);
nor U8372 (N_8372,N_6960,N_6357);
nand U8373 (N_8373,N_7935,N_6177);
nor U8374 (N_8374,N_6089,N_7637);
and U8375 (N_8375,N_7953,N_6988);
xnor U8376 (N_8376,N_7125,N_6161);
nand U8377 (N_8377,N_7919,N_7373);
nor U8378 (N_8378,N_7055,N_6736);
and U8379 (N_8379,N_6353,N_7088);
nor U8380 (N_8380,N_6346,N_6006);
and U8381 (N_8381,N_7157,N_7625);
nor U8382 (N_8382,N_6708,N_6366);
nor U8383 (N_8383,N_7620,N_7695);
and U8384 (N_8384,N_6428,N_6106);
nand U8385 (N_8385,N_6793,N_6185);
nand U8386 (N_8386,N_7761,N_6419);
or U8387 (N_8387,N_6240,N_6910);
nor U8388 (N_8388,N_6345,N_7215);
or U8389 (N_8389,N_7206,N_6452);
and U8390 (N_8390,N_7810,N_6984);
and U8391 (N_8391,N_7110,N_6835);
nand U8392 (N_8392,N_7725,N_7830);
and U8393 (N_8393,N_7186,N_6787);
nand U8394 (N_8394,N_6836,N_6636);
nor U8395 (N_8395,N_7112,N_6979);
nand U8396 (N_8396,N_6904,N_7273);
nor U8397 (N_8397,N_6470,N_7380);
or U8398 (N_8398,N_7404,N_6223);
and U8399 (N_8399,N_7993,N_7990);
nand U8400 (N_8400,N_6830,N_7297);
nor U8401 (N_8401,N_6450,N_6639);
or U8402 (N_8402,N_6795,N_7044);
and U8403 (N_8403,N_7243,N_6480);
and U8404 (N_8404,N_6282,N_7617);
or U8405 (N_8405,N_7987,N_7653);
nor U8406 (N_8406,N_7181,N_6076);
nor U8407 (N_8407,N_6510,N_6765);
or U8408 (N_8408,N_6414,N_7656);
nor U8409 (N_8409,N_7562,N_7847);
and U8410 (N_8410,N_6322,N_6308);
and U8411 (N_8411,N_6468,N_6682);
nand U8412 (N_8412,N_6176,N_6312);
nor U8413 (N_8413,N_7037,N_7715);
or U8414 (N_8414,N_6540,N_7766);
nor U8415 (N_8415,N_7712,N_7844);
nor U8416 (N_8416,N_7871,N_7109);
nand U8417 (N_8417,N_7597,N_7749);
and U8418 (N_8418,N_6314,N_7116);
nor U8419 (N_8419,N_6570,N_6262);
nor U8420 (N_8420,N_7934,N_7200);
and U8421 (N_8421,N_7783,N_6026);
nor U8422 (N_8422,N_7515,N_7618);
nand U8423 (N_8423,N_6533,N_7908);
or U8424 (N_8424,N_6838,N_7490);
xnor U8425 (N_8425,N_6924,N_7565);
nor U8426 (N_8426,N_6536,N_7674);
or U8427 (N_8427,N_7995,N_6103);
and U8428 (N_8428,N_7811,N_7721);
or U8429 (N_8429,N_6903,N_7931);
nor U8430 (N_8430,N_6449,N_6864);
nand U8431 (N_8431,N_6108,N_6399);
or U8432 (N_8432,N_6873,N_7203);
nor U8433 (N_8433,N_6335,N_7627);
xor U8434 (N_8434,N_6211,N_7153);
nand U8435 (N_8435,N_6993,N_7188);
or U8436 (N_8436,N_6041,N_6302);
nand U8437 (N_8437,N_7101,N_7816);
nand U8438 (N_8438,N_6269,N_6947);
nor U8439 (N_8439,N_6454,N_7708);
or U8440 (N_8440,N_6674,N_7550);
xor U8441 (N_8441,N_6930,N_7450);
or U8442 (N_8442,N_6560,N_7465);
xnor U8443 (N_8443,N_6539,N_6020);
nor U8444 (N_8444,N_7547,N_7688);
nor U8445 (N_8445,N_7444,N_6330);
nor U8446 (N_8446,N_6133,N_6050);
xnor U8447 (N_8447,N_6771,N_6681);
or U8448 (N_8448,N_7804,N_7735);
and U8449 (N_8449,N_7245,N_6466);
nor U8450 (N_8450,N_7355,N_7426);
xnor U8451 (N_8451,N_7062,N_6392);
or U8452 (N_8452,N_6044,N_7932);
nand U8453 (N_8453,N_7311,N_7560);
or U8454 (N_8454,N_6421,N_6055);
xnor U8455 (N_8455,N_6210,N_6356);
nand U8456 (N_8456,N_6196,N_6710);
nand U8457 (N_8457,N_7807,N_6435);
and U8458 (N_8458,N_6512,N_6858);
or U8459 (N_8459,N_7896,N_6897);
and U8460 (N_8460,N_7920,N_6602);
xnor U8461 (N_8461,N_7379,N_7950);
nor U8462 (N_8462,N_6786,N_7072);
or U8463 (N_8463,N_7722,N_7831);
xor U8464 (N_8464,N_7440,N_6075);
nand U8465 (N_8465,N_6891,N_6817);
xnor U8466 (N_8466,N_7388,N_7851);
xor U8467 (N_8467,N_6763,N_6053);
and U8468 (N_8468,N_6354,N_7583);
nor U8469 (N_8469,N_7728,N_6705);
or U8470 (N_8470,N_7541,N_7563);
nand U8471 (N_8471,N_7301,N_7875);
xnor U8472 (N_8472,N_7331,N_7121);
nand U8473 (N_8473,N_6770,N_7965);
nor U8474 (N_8474,N_7105,N_6104);
or U8475 (N_8475,N_6872,N_7004);
and U8476 (N_8476,N_6957,N_6789);
or U8477 (N_8477,N_7870,N_6595);
or U8478 (N_8478,N_7643,N_6471);
xor U8479 (N_8479,N_7177,N_7045);
nand U8480 (N_8480,N_7690,N_7234);
and U8481 (N_8481,N_6265,N_7820);
nand U8482 (N_8482,N_7985,N_7639);
and U8483 (N_8483,N_6025,N_7190);
nand U8484 (N_8484,N_7629,N_7603);
or U8485 (N_8485,N_6888,N_6755);
nand U8486 (N_8486,N_7821,N_7259);
or U8487 (N_8487,N_7958,N_7480);
or U8488 (N_8488,N_7921,N_6127);
xor U8489 (N_8489,N_7138,N_7713);
nor U8490 (N_8490,N_6664,N_6145);
and U8491 (N_8491,N_6568,N_7340);
nor U8492 (N_8492,N_7581,N_6912);
nand U8493 (N_8493,N_7356,N_7768);
nand U8494 (N_8494,N_7986,N_7382);
nor U8495 (N_8495,N_6779,N_6856);
or U8496 (N_8496,N_6009,N_6644);
xnor U8497 (N_8497,N_7964,N_6657);
xnor U8498 (N_8498,N_7736,N_6024);
and U8499 (N_8499,N_7740,N_7750);
or U8500 (N_8500,N_7275,N_7485);
and U8501 (N_8501,N_7876,N_6122);
nor U8502 (N_8502,N_7537,N_6585);
and U8503 (N_8503,N_6649,N_6609);
or U8504 (N_8504,N_7866,N_6344);
or U8505 (N_8505,N_7590,N_6530);
or U8506 (N_8506,N_7685,N_7422);
nor U8507 (N_8507,N_7758,N_7647);
nand U8508 (N_8508,N_7458,N_6147);
and U8509 (N_8509,N_6186,N_6289);
nand U8510 (N_8510,N_7371,N_7173);
nor U8511 (N_8511,N_6296,N_7231);
or U8512 (N_8512,N_6752,N_7619);
nor U8513 (N_8513,N_6911,N_7402);
nand U8514 (N_8514,N_7837,N_7077);
nor U8515 (N_8515,N_7863,N_7782);
nand U8516 (N_8516,N_6884,N_7672);
nand U8517 (N_8517,N_7330,N_6066);
and U8518 (N_8518,N_7462,N_6403);
nor U8519 (N_8519,N_7791,N_7018);
nor U8520 (N_8520,N_6928,N_7119);
nand U8521 (N_8521,N_6962,N_6438);
or U8522 (N_8522,N_7464,N_7041);
xnor U8523 (N_8523,N_7526,N_7204);
xor U8524 (N_8524,N_6919,N_6096);
nand U8525 (N_8525,N_7134,N_6391);
or U8526 (N_8526,N_7923,N_7397);
nor U8527 (N_8527,N_6129,N_7507);
and U8528 (N_8528,N_6058,N_6553);
nor U8529 (N_8529,N_6117,N_6626);
and U8530 (N_8530,N_6056,N_7790);
nand U8531 (N_8531,N_6216,N_6182);
and U8532 (N_8532,N_6815,N_7737);
or U8533 (N_8533,N_6584,N_6967);
nor U8534 (N_8534,N_7927,N_6208);
xor U8535 (N_8535,N_6826,N_6206);
nand U8536 (N_8536,N_6687,N_7384);
or U8537 (N_8537,N_6487,N_7709);
nand U8538 (N_8538,N_7155,N_6816);
or U8539 (N_8539,N_7454,N_7086);
nand U8540 (N_8540,N_6679,N_7648);
xor U8541 (N_8541,N_6201,N_6195);
and U8542 (N_8542,N_7928,N_6767);
and U8543 (N_8543,N_6719,N_7594);
nand U8544 (N_8544,N_7393,N_6768);
nand U8545 (N_8545,N_7730,N_6556);
and U8546 (N_8546,N_7910,N_7319);
nor U8547 (N_8547,N_6954,N_6976);
xor U8548 (N_8548,N_6307,N_7359);
and U8549 (N_8549,N_6811,N_7348);
nor U8550 (N_8550,N_7797,N_7080);
nand U8551 (N_8551,N_6790,N_6394);
nand U8552 (N_8552,N_7484,N_6822);
nor U8553 (N_8553,N_6339,N_6442);
nand U8554 (N_8554,N_7947,N_6332);
nand U8555 (N_8555,N_7058,N_6857);
nand U8556 (N_8556,N_7409,N_6278);
nor U8557 (N_8557,N_7418,N_7650);
and U8558 (N_8558,N_7732,N_6808);
and U8559 (N_8559,N_7069,N_7165);
nand U8560 (N_8560,N_6199,N_7225);
and U8561 (N_8561,N_6531,N_7253);
nor U8562 (N_8562,N_7325,N_7247);
or U8563 (N_8563,N_6498,N_6167);
nor U8564 (N_8564,N_6372,N_6321);
nor U8565 (N_8565,N_6938,N_7649);
nor U8566 (N_8566,N_6257,N_6572);
and U8567 (N_8567,N_7949,N_6159);
nand U8568 (N_8568,N_6051,N_7040);
nand U8569 (N_8569,N_7023,N_6476);
nor U8570 (N_8570,N_7469,N_6347);
nand U8571 (N_8571,N_7564,N_6515);
or U8572 (N_8572,N_7391,N_7612);
xnor U8573 (N_8573,N_6082,N_6131);
or U8574 (N_8574,N_6583,N_7448);
and U8575 (N_8575,N_6359,N_7147);
nand U8576 (N_8576,N_7303,N_7815);
nand U8577 (N_8577,N_7199,N_7872);
and U8578 (N_8578,N_7130,N_7236);
nand U8579 (N_8579,N_7586,N_7396);
nand U8580 (N_8580,N_6500,N_6252);
nor U8581 (N_8581,N_6396,N_7834);
and U8582 (N_8582,N_6393,N_7652);
or U8583 (N_8583,N_6932,N_7148);
nor U8584 (N_8584,N_7013,N_6150);
or U8585 (N_8585,N_7178,N_7917);
or U8586 (N_8586,N_6848,N_6113);
nor U8587 (N_8587,N_6743,N_7511);
nor U8588 (N_8588,N_6175,N_7060);
nand U8589 (N_8589,N_7505,N_7417);
nand U8590 (N_8590,N_7789,N_6545);
nand U8591 (N_8591,N_7946,N_7580);
nand U8592 (N_8592,N_6711,N_7542);
xnor U8593 (N_8593,N_6934,N_6064);
xor U8594 (N_8594,N_7230,N_7292);
and U8595 (N_8595,N_6694,N_7930);
nand U8596 (N_8596,N_7466,N_6303);
nand U8597 (N_8597,N_7970,N_7159);
and U8598 (N_8598,N_6948,N_7969);
and U8599 (N_8599,N_6670,N_6951);
and U8600 (N_8600,N_7925,N_7043);
nand U8601 (N_8601,N_7106,N_7675);
nand U8602 (N_8602,N_6432,N_7502);
or U8603 (N_8603,N_6507,N_6860);
and U8604 (N_8604,N_7022,N_6236);
and U8605 (N_8605,N_7659,N_7328);
nor U8606 (N_8606,N_6239,N_6205);
or U8607 (N_8607,N_7036,N_7221);
nand U8608 (N_8608,N_7451,N_7679);
and U8609 (N_8609,N_7660,N_7433);
or U8610 (N_8610,N_7183,N_6661);
nor U8611 (N_8611,N_7902,N_6038);
xnor U8612 (N_8612,N_6807,N_7959);
or U8613 (N_8613,N_6624,N_6878);
nor U8614 (N_8614,N_7304,N_6876);
xnor U8615 (N_8615,N_7954,N_6921);
nand U8616 (N_8616,N_7228,N_6973);
nand U8617 (N_8617,N_7254,N_7102);
nor U8618 (N_8618,N_6855,N_6331);
xor U8619 (N_8619,N_6111,N_6715);
nand U8620 (N_8620,N_7853,N_7394);
or U8621 (N_8621,N_6125,N_6048);
or U8622 (N_8622,N_6961,N_7364);
or U8623 (N_8623,N_6036,N_6543);
nand U8624 (N_8624,N_6233,N_6968);
and U8625 (N_8625,N_6395,N_7358);
and U8626 (N_8626,N_7610,N_7836);
or U8627 (N_8627,N_7334,N_6972);
xnor U8628 (N_8628,N_6567,N_7533);
nand U8629 (N_8629,N_7367,N_6831);
xnor U8630 (N_8630,N_6902,N_6033);
nand U8631 (N_8631,N_6495,N_6197);
nand U8632 (N_8632,N_6894,N_7776);
or U8633 (N_8633,N_7028,N_7209);
and U8634 (N_8634,N_6757,N_7323);
nor U8635 (N_8635,N_7491,N_7210);
nor U8636 (N_8636,N_6977,N_7324);
and U8637 (N_8637,N_7978,N_6658);
nor U8638 (N_8638,N_6772,N_6084);
or U8639 (N_8639,N_6939,N_6093);
or U8640 (N_8640,N_7886,N_7160);
or U8641 (N_8641,N_7074,N_6728);
xor U8642 (N_8642,N_6146,N_6477);
or U8643 (N_8643,N_7843,N_7630);
and U8644 (N_8644,N_7189,N_6950);
or U8645 (N_8645,N_7216,N_7405);
and U8646 (N_8646,N_6355,N_6879);
nand U8647 (N_8647,N_7201,N_7794);
nand U8648 (N_8648,N_7683,N_6249);
and U8649 (N_8649,N_7663,N_7753);
or U8650 (N_8650,N_6107,N_6232);
and U8651 (N_8651,N_6126,N_6803);
nand U8652 (N_8652,N_6611,N_6078);
and U8653 (N_8653,N_7338,N_7269);
and U8654 (N_8654,N_7963,N_6000);
or U8655 (N_8655,N_6042,N_7609);
xor U8656 (N_8656,N_6866,N_6367);
nor U8657 (N_8657,N_6741,N_7988);
nand U8658 (N_8658,N_7862,N_7000);
nand U8659 (N_8659,N_7370,N_6739);
nor U8660 (N_8660,N_7233,N_6750);
nor U8661 (N_8661,N_7415,N_6342);
nor U8662 (N_8662,N_6725,N_7369);
nand U8663 (N_8663,N_7343,N_7621);
nand U8664 (N_8664,N_6522,N_6804);
or U8665 (N_8665,N_7104,N_7967);
nand U8666 (N_8666,N_6655,N_6309);
nor U8667 (N_8667,N_7720,N_6467);
or U8668 (N_8668,N_6871,N_6465);
nor U8669 (N_8669,N_6944,N_7494);
nand U8670 (N_8670,N_7812,N_7071);
xor U8671 (N_8671,N_7475,N_7192);
nor U8672 (N_8672,N_7531,N_6839);
nor U8673 (N_8673,N_7890,N_7352);
or U8674 (N_8674,N_7754,N_6258);
or U8675 (N_8675,N_7764,N_6313);
nand U8676 (N_8676,N_6840,N_6727);
xnor U8677 (N_8677,N_6097,N_6023);
or U8678 (N_8678,N_7746,N_6062);
or U8679 (N_8679,N_7341,N_7579);
nor U8680 (N_8680,N_6502,N_6170);
or U8681 (N_8681,N_6781,N_6940);
xnor U8682 (N_8682,N_7903,N_6506);
and U8683 (N_8683,N_7097,N_6323);
nand U8684 (N_8684,N_7133,N_6819);
nand U8685 (N_8685,N_6648,N_6241);
or U8686 (N_8686,N_7390,N_6157);
or U8687 (N_8687,N_7030,N_7622);
nand U8688 (N_8688,N_6605,N_7008);
nand U8689 (N_8689,N_6274,N_6505);
and U8690 (N_8690,N_6283,N_6729);
nand U8691 (N_8691,N_6463,N_7726);
nand U8692 (N_8692,N_7860,N_6598);
nand U8693 (N_8693,N_6135,N_6742);
nand U8694 (N_8694,N_7242,N_7607);
or U8695 (N_8695,N_6389,N_6028);
nor U8696 (N_8696,N_7861,N_6642);
and U8697 (N_8697,N_6336,N_7814);
nand U8698 (N_8698,N_7632,N_7704);
and U8699 (N_8699,N_6171,N_6619);
and U8700 (N_8700,N_7107,N_6276);
nor U8701 (N_8701,N_6245,N_7636);
nand U8702 (N_8702,N_6349,N_6109);
and U8703 (N_8703,N_7142,N_6613);
and U8704 (N_8704,N_7548,N_7029);
nand U8705 (N_8705,N_6532,N_7461);
nand U8706 (N_8706,N_6325,N_6439);
or U8707 (N_8707,N_6224,N_6927);
nand U8708 (N_8708,N_6717,N_7676);
xnor U8709 (N_8709,N_7385,N_7067);
or U8710 (N_8710,N_6190,N_7504);
or U8711 (N_8711,N_6493,N_7267);
or U8712 (N_8712,N_7455,N_7276);
nand U8713 (N_8713,N_7474,N_6065);
nor U8714 (N_8714,N_7818,N_6643);
or U8715 (N_8715,N_6889,N_6348);
or U8716 (N_8716,N_7869,N_7239);
and U8717 (N_8717,N_7929,N_6778);
and U8718 (N_8718,N_6101,N_6513);
and U8719 (N_8719,N_6523,N_6222);
or U8720 (N_8720,N_6124,N_7260);
or U8721 (N_8721,N_7372,N_7724);
nand U8722 (N_8722,N_7705,N_6328);
nor U8723 (N_8723,N_6996,N_6375);
or U8724 (N_8724,N_6806,N_7118);
xor U8725 (N_8725,N_6151,N_6060);
or U8726 (N_8726,N_6994,N_7320);
or U8727 (N_8727,N_7020,N_6030);
and U8728 (N_8728,N_6749,N_7172);
nand U8729 (N_8729,N_6390,N_6168);
nand U8730 (N_8730,N_6566,N_6034);
and U8731 (N_8731,N_7435,N_6576);
xor U8732 (N_8732,N_6300,N_6441);
nor U8733 (N_8733,N_7351,N_7962);
nand U8734 (N_8734,N_6287,N_7308);
or U8735 (N_8735,N_6635,N_7197);
or U8736 (N_8736,N_6981,N_6913);
nand U8737 (N_8737,N_7246,N_7898);
nor U8738 (N_8738,N_6726,N_6999);
xor U8739 (N_8739,N_6791,N_7224);
nand U8740 (N_8740,N_7524,N_7193);
or U8741 (N_8741,N_7184,N_6187);
or U8742 (N_8742,N_7430,N_6363);
nand U8743 (N_8743,N_6425,N_7992);
xor U8744 (N_8744,N_7284,N_7229);
nor U8745 (N_8745,N_7205,N_6462);
xnor U8746 (N_8746,N_6180,N_7655);
and U8747 (N_8747,N_6234,N_7111);
nor U8748 (N_8748,N_7773,N_7974);
nor U8749 (N_8749,N_6141,N_7149);
or U8750 (N_8750,N_7718,N_7425);
nand U8751 (N_8751,N_6714,N_7223);
or U8752 (N_8752,N_7523,N_7536);
nor U8753 (N_8753,N_6243,N_6250);
nand U8754 (N_8754,N_6721,N_7711);
nor U8755 (N_8755,N_6174,N_6863);
or U8756 (N_8756,N_6524,N_7429);
and U8757 (N_8757,N_7661,N_6142);
nand U8758 (N_8758,N_7785,N_7784);
and U8759 (N_8759,N_6486,N_7616);
and U8760 (N_8760,N_7891,N_6985);
or U8761 (N_8761,N_6637,N_6701);
and U8762 (N_8762,N_6615,N_7833);
xnor U8763 (N_8763,N_6579,N_6416);
nor U8764 (N_8764,N_7083,N_6402);
xor U8765 (N_8765,N_7574,N_7803);
nor U8766 (N_8766,N_7867,N_6764);
or U8767 (N_8767,N_6297,N_6130);
xnor U8768 (N_8768,N_6844,N_6677);
xor U8769 (N_8769,N_6784,N_6890);
and U8770 (N_8770,N_6680,N_7850);
nor U8771 (N_8771,N_6601,N_6072);
or U8772 (N_8772,N_6123,N_7374);
nor U8773 (N_8773,N_7012,N_6091);
nand U8774 (N_8774,N_7306,N_6404);
nor U8775 (N_8775,N_6320,N_6526);
nand U8776 (N_8776,N_6665,N_6285);
and U8777 (N_8777,N_6081,N_6204);
and U8778 (N_8778,N_7427,N_6518);
and U8779 (N_8779,N_7900,N_6991);
nor U8780 (N_8780,N_6080,N_6437);
nor U8781 (N_8781,N_6266,N_7252);
or U8782 (N_8782,N_7244,N_6883);
nand U8783 (N_8783,N_6971,N_7911);
or U8784 (N_8784,N_7039,N_6455);
xor U8785 (N_8785,N_7477,N_7262);
and U8786 (N_8786,N_6440,N_6980);
or U8787 (N_8787,N_6751,N_6607);
nor U8788 (N_8788,N_7103,N_7335);
or U8789 (N_8789,N_6706,N_7573);
xor U8790 (N_8790,N_6364,N_6847);
or U8791 (N_8791,N_7587,N_7696);
or U8792 (N_8792,N_7881,N_6722);
nand U8793 (N_8793,N_7169,N_6001);
or U8794 (N_8794,N_6478,N_6229);
and U8795 (N_8795,N_6542,N_7727);
and U8796 (N_8796,N_6660,N_6004);
nand U8797 (N_8797,N_7771,N_7664);
nand U8798 (N_8798,N_6069,N_6378);
or U8799 (N_8799,N_6852,N_6945);
and U8800 (N_8800,N_7293,N_6288);
nand U8801 (N_8801,N_6509,N_7678);
nor U8802 (N_8802,N_6582,N_6272);
nand U8803 (N_8803,N_7412,N_6214);
nor U8804 (N_8804,N_7011,N_7945);
or U8805 (N_8805,N_6667,N_6326);
and U8806 (N_8806,N_7423,N_7748);
and U8807 (N_8807,N_7272,N_6845);
xnor U8808 (N_8808,N_7723,N_6735);
and U8809 (N_8809,N_7214,N_6281);
xor U8810 (N_8810,N_6885,N_6306);
nand U8811 (N_8811,N_7681,N_7914);
nand U8812 (N_8812,N_7539,N_7633);
xnor U8813 (N_8813,N_7202,N_6580);
nand U8814 (N_8814,N_7363,N_7858);
and U8815 (N_8815,N_7406,N_7010);
nor U8816 (N_8816,N_6922,N_6792);
nor U8817 (N_8817,N_7499,N_6846);
or U8818 (N_8818,N_7907,N_7117);
nand U8819 (N_8819,N_6114,N_6496);
and U8820 (N_8820,N_7194,N_6801);
nor U8821 (N_8821,N_7282,N_6600);
and U8822 (N_8822,N_6458,N_6037);
and U8823 (N_8823,N_7122,N_7174);
xor U8824 (N_8824,N_7657,N_6900);
nor U8825 (N_8825,N_6474,N_7997);
and U8826 (N_8826,N_6316,N_7530);
nand U8827 (N_8827,N_6235,N_6997);
nor U8828 (N_8828,N_6430,N_7849);
xnor U8829 (N_8829,N_7558,N_6264);
and U8830 (N_8830,N_7163,N_6603);
or U8831 (N_8831,N_6134,N_6915);
or U8832 (N_8832,N_6551,N_6095);
nand U8833 (N_8833,N_6384,N_6850);
nand U8834 (N_8834,N_6802,N_6854);
xnor U8835 (N_8835,N_7770,N_7220);
nor U8836 (N_8836,N_7016,N_7901);
nand U8837 (N_8837,N_7176,N_6490);
and U8838 (N_8838,N_7601,N_7944);
nand U8839 (N_8839,N_7483,N_7937);
nor U8840 (N_8840,N_6581,N_6213);
nand U8841 (N_8841,N_7717,N_6099);
nand U8842 (N_8842,N_7033,N_7857);
nand U8843 (N_8843,N_7218,N_6599);
xnor U8844 (N_8844,N_6825,N_6417);
or U8845 (N_8845,N_6254,N_6018);
nand U8846 (N_8846,N_7631,N_6520);
nand U8847 (N_8847,N_7357,N_7437);
or U8848 (N_8848,N_7411,N_7322);
or U8849 (N_8849,N_6010,N_6936);
nand U8850 (N_8850,N_6085,N_6926);
or U8851 (N_8851,N_7569,N_7295);
and U8852 (N_8852,N_7021,N_6173);
nor U8853 (N_8853,N_7568,N_7665);
xnor U8854 (N_8854,N_7680,N_7408);
nor U8855 (N_8855,N_6398,N_7693);
and U8856 (N_8856,N_7592,N_7375);
and U8857 (N_8857,N_7094,N_6446);
nor U8858 (N_8858,N_6259,N_6738);
or U8859 (N_8859,N_7368,N_6547);
nand U8860 (N_8860,N_6777,N_7226);
and U8861 (N_8861,N_7994,N_7973);
and U8862 (N_8862,N_7535,N_7310);
and U8863 (N_8863,N_6497,N_7064);
nand U8864 (N_8864,N_7912,N_6179);
nor U8865 (N_8865,N_6244,N_7829);
nor U8866 (N_8866,N_7001,N_6916);
nand U8867 (N_8867,N_7146,N_6783);
or U8868 (N_8868,N_7051,N_6689);
and U8869 (N_8869,N_7522,N_6821);
nor U8870 (N_8870,N_7792,N_6110);
or U8871 (N_8871,N_6027,N_7589);
nor U8872 (N_8872,N_7339,N_7752);
nand U8873 (N_8873,N_6632,N_6341);
xnor U8874 (N_8874,N_7342,N_7336);
and U8875 (N_8875,N_6989,N_6488);
xor U8876 (N_8876,N_6035,N_7042);
xnor U8877 (N_8877,N_7208,N_7595);
or U8878 (N_8878,N_7419,N_6673);
and U8879 (N_8879,N_6693,N_6565);
nor U8880 (N_8880,N_7129,N_7057);
or U8881 (N_8881,N_7398,N_6651);
and U8882 (N_8882,N_6358,N_7957);
xnor U8883 (N_8883,N_6100,N_6837);
or U8884 (N_8884,N_6754,N_6411);
nor U8885 (N_8885,N_6955,N_7487);
nor U8886 (N_8886,N_7991,N_6405);
and U8887 (N_8887,N_6136,N_6383);
xor U8888 (N_8888,N_7585,N_7972);
and U8889 (N_8889,N_7508,N_6045);
nand U8890 (N_8890,N_6573,N_7389);
nor U8891 (N_8891,N_7473,N_6340);
or U8892 (N_8892,N_6333,N_6574);
nand U8893 (N_8893,N_6451,N_7305);
nor U8894 (N_8894,N_7918,N_7140);
nand U8895 (N_8895,N_6191,N_6907);
or U8896 (N_8896,N_7989,N_7096);
nor U8897 (N_8897,N_6990,N_6231);
nand U8898 (N_8898,N_7635,N_6469);
or U8899 (N_8899,N_6666,N_7017);
nand U8900 (N_8900,N_7453,N_7878);
nor U8901 (N_8901,N_6343,N_7002);
xor U8902 (N_8902,N_7546,N_7073);
xnor U8903 (N_8903,N_7460,N_6194);
and U8904 (N_8904,N_7543,N_7702);
xnor U8905 (N_8905,N_7439,N_6327);
nor U8906 (N_8906,N_6059,N_7255);
nand U8907 (N_8907,N_6823,N_7493);
and U8908 (N_8908,N_7470,N_7593);
and U8909 (N_8909,N_7151,N_7654);
nand U8910 (N_8910,N_7467,N_6562);
xor U8911 (N_8911,N_6251,N_6184);
and U8912 (N_8912,N_7731,N_6324);
and U8913 (N_8913,N_6557,N_6350);
nor U8914 (N_8914,N_7968,N_7998);
or U8915 (N_8915,N_6154,N_6575);
and U8916 (N_8916,N_6054,N_7479);
or U8917 (N_8917,N_7166,N_6809);
or U8918 (N_8918,N_6310,N_6371);
and U8919 (N_8919,N_7684,N_6740);
or U8920 (N_8920,N_6882,N_6017);
nor U8921 (N_8921,N_7407,N_7090);
nor U8922 (N_8922,N_6318,N_6986);
and U8923 (N_8923,N_7588,N_6548);
and U8924 (N_8924,N_7068,N_7667);
nand U8925 (N_8925,N_7164,N_6596);
and U8926 (N_8926,N_6614,N_6923);
nand U8927 (N_8927,N_7198,N_6261);
nand U8928 (N_8928,N_6365,N_6139);
xor U8929 (N_8929,N_7248,N_6005);
or U8930 (N_8930,N_7420,N_7250);
and U8931 (N_8931,N_7605,N_6115);
and U8932 (N_8932,N_6975,N_6489);
or U8933 (N_8933,N_7582,N_7099);
nand U8934 (N_8934,N_7757,N_7926);
and U8935 (N_8935,N_7154,N_7050);
and U8936 (N_8936,N_7227,N_7263);
nor U8937 (N_8937,N_7687,N_6311);
or U8938 (N_8938,N_6773,N_7315);
or U8939 (N_8939,N_7955,N_6270);
xnor U8940 (N_8940,N_7795,N_7446);
xor U8941 (N_8941,N_7938,N_7003);
nand U8942 (N_8942,N_6974,N_7026);
or U8943 (N_8943,N_7095,N_7716);
nor U8944 (N_8944,N_6299,N_6070);
nand U8945 (N_8945,N_7765,N_7644);
xnor U8946 (N_8946,N_6119,N_6685);
nand U8947 (N_8947,N_6604,N_7786);
nor U8948 (N_8948,N_7498,N_6859);
and U8949 (N_8949,N_6851,N_7168);
and U8950 (N_8950,N_7799,N_7824);
nor U8951 (N_8951,N_7191,N_6906);
nand U8952 (N_8952,N_7182,N_6853);
nand U8953 (N_8953,N_7915,N_6011);
or U8954 (N_8954,N_7651,N_6338);
nand U8955 (N_8955,N_7278,N_7623);
nand U8956 (N_8956,N_6780,N_7006);
and U8957 (N_8957,N_7337,N_7529);
and U8958 (N_8958,N_7180,N_6631);
xor U8959 (N_8959,N_6937,N_6552);
nor U8960 (N_8960,N_7606,N_7806);
nor U8961 (N_8961,N_7596,N_7326);
nor U8962 (N_8962,N_6877,N_7854);
nand U8963 (N_8963,N_6079,N_7436);
nand U8964 (N_8964,N_7506,N_7488);
and U8965 (N_8965,N_7232,N_7525);
and U8966 (N_8966,N_7762,N_6049);
nand U8967 (N_8967,N_7158,N_7376);
nand U8968 (N_8968,N_6587,N_7763);
nand U8969 (N_8969,N_7841,N_6707);
or U8970 (N_8970,N_7078,N_7856);
or U8971 (N_8971,N_6386,N_7897);
and U8972 (N_8972,N_7571,N_7793);
nor U8973 (N_8973,N_6193,N_7298);
or U8974 (N_8974,N_6074,N_7641);
nand U8975 (N_8975,N_6762,N_6638);
nand U8976 (N_8976,N_7817,N_6761);
xnor U8977 (N_8977,N_6461,N_6684);
nor U8978 (N_8978,N_6319,N_7787);
nand U8979 (N_8979,N_7544,N_6377);
nand U8980 (N_8980,N_6820,N_6698);
nand U8981 (N_8981,N_6219,N_6400);
nand U8982 (N_8982,N_7211,N_6491);
nand U8983 (N_8983,N_6541,N_7899);
and U8984 (N_8984,N_7880,N_7084);
and U8985 (N_8985,N_7895,N_7399);
nand U8986 (N_8986,N_7081,N_7703);
nand U8987 (N_8987,N_7145,N_7079);
nor U8988 (N_8988,N_6238,N_6671);
nand U8989 (N_8989,N_7286,N_7952);
or U8990 (N_8990,N_7251,N_6849);
or U8991 (N_8991,N_7838,N_6691);
xor U8992 (N_8992,N_6712,N_6700);
nand U8993 (N_8993,N_6412,N_6734);
or U8994 (N_8994,N_6294,N_6501);
and U8995 (N_8995,N_7128,N_6797);
and U8996 (N_8996,N_7828,N_6163);
nand U8997 (N_8997,N_7115,N_6887);
and U8998 (N_8998,N_7171,N_6616);
xor U8999 (N_8999,N_7447,N_6137);
nand U9000 (N_9000,N_7870,N_7046);
or U9001 (N_9001,N_6687,N_7707);
and U9002 (N_9002,N_6060,N_6326);
nand U9003 (N_9003,N_6828,N_7140);
xnor U9004 (N_9004,N_6376,N_6991);
nor U9005 (N_9005,N_7476,N_6872);
or U9006 (N_9006,N_6399,N_6208);
xnor U9007 (N_9007,N_7258,N_6776);
nor U9008 (N_9008,N_6836,N_6378);
nand U9009 (N_9009,N_7103,N_6352);
and U9010 (N_9010,N_7731,N_6790);
or U9011 (N_9011,N_6969,N_7296);
xor U9012 (N_9012,N_6568,N_6783);
nor U9013 (N_9013,N_7302,N_6795);
nand U9014 (N_9014,N_6675,N_7455);
nand U9015 (N_9015,N_7885,N_6359);
nor U9016 (N_9016,N_7469,N_6000);
nand U9017 (N_9017,N_7092,N_7680);
nor U9018 (N_9018,N_7098,N_7807);
xnor U9019 (N_9019,N_7540,N_7915);
nand U9020 (N_9020,N_6274,N_6865);
or U9021 (N_9021,N_6727,N_6567);
and U9022 (N_9022,N_7718,N_7422);
and U9023 (N_9023,N_6879,N_6712);
nand U9024 (N_9024,N_6226,N_6607);
and U9025 (N_9025,N_7408,N_6941);
xnor U9026 (N_9026,N_6065,N_6352);
nor U9027 (N_9027,N_6933,N_7648);
nand U9028 (N_9028,N_6270,N_7367);
xor U9029 (N_9029,N_6786,N_7924);
nor U9030 (N_9030,N_6207,N_6846);
nor U9031 (N_9031,N_7881,N_6960);
nor U9032 (N_9032,N_7897,N_6732);
nand U9033 (N_9033,N_7935,N_6882);
or U9034 (N_9034,N_7258,N_7380);
or U9035 (N_9035,N_6115,N_6348);
nand U9036 (N_9036,N_7979,N_7693);
nand U9037 (N_9037,N_7082,N_7918);
and U9038 (N_9038,N_7991,N_7418);
xnor U9039 (N_9039,N_6409,N_6152);
nand U9040 (N_9040,N_7543,N_7617);
xor U9041 (N_9041,N_7105,N_6131);
or U9042 (N_9042,N_7144,N_7649);
and U9043 (N_9043,N_6895,N_6350);
or U9044 (N_9044,N_7492,N_7452);
nor U9045 (N_9045,N_6191,N_7884);
and U9046 (N_9046,N_7272,N_6093);
or U9047 (N_9047,N_7862,N_7732);
nor U9048 (N_9048,N_6731,N_6851);
or U9049 (N_9049,N_7193,N_6428);
or U9050 (N_9050,N_6989,N_7768);
and U9051 (N_9051,N_7250,N_7658);
and U9052 (N_9052,N_6035,N_6915);
or U9053 (N_9053,N_7710,N_7975);
nand U9054 (N_9054,N_6120,N_6546);
nor U9055 (N_9055,N_7369,N_7619);
nor U9056 (N_9056,N_6783,N_6315);
nor U9057 (N_9057,N_7679,N_6258);
and U9058 (N_9058,N_7123,N_7735);
and U9059 (N_9059,N_6966,N_7518);
or U9060 (N_9060,N_7167,N_7275);
nand U9061 (N_9061,N_7991,N_6726);
and U9062 (N_9062,N_6902,N_7466);
or U9063 (N_9063,N_7097,N_7153);
nand U9064 (N_9064,N_6752,N_7728);
nand U9065 (N_9065,N_6949,N_7384);
or U9066 (N_9066,N_7236,N_7856);
and U9067 (N_9067,N_6051,N_6688);
nand U9068 (N_9068,N_7676,N_6465);
nand U9069 (N_9069,N_6233,N_7330);
and U9070 (N_9070,N_7214,N_7385);
and U9071 (N_9071,N_7408,N_6004);
and U9072 (N_9072,N_7125,N_7667);
and U9073 (N_9073,N_7779,N_6509);
nand U9074 (N_9074,N_6386,N_6271);
nand U9075 (N_9075,N_7458,N_6480);
nand U9076 (N_9076,N_6537,N_6365);
nor U9077 (N_9077,N_7309,N_6485);
or U9078 (N_9078,N_6080,N_7190);
nand U9079 (N_9079,N_6557,N_6077);
nand U9080 (N_9080,N_7100,N_7653);
nor U9081 (N_9081,N_6199,N_7023);
nand U9082 (N_9082,N_6345,N_6503);
nand U9083 (N_9083,N_6383,N_6896);
and U9084 (N_9084,N_7123,N_6355);
xor U9085 (N_9085,N_7149,N_6760);
nand U9086 (N_9086,N_7109,N_7305);
and U9087 (N_9087,N_7222,N_7284);
nor U9088 (N_9088,N_6778,N_6417);
nand U9089 (N_9089,N_7426,N_6716);
nand U9090 (N_9090,N_7499,N_6889);
nor U9091 (N_9091,N_6818,N_7511);
or U9092 (N_9092,N_7768,N_6300);
nand U9093 (N_9093,N_7150,N_6391);
nor U9094 (N_9094,N_7044,N_7478);
or U9095 (N_9095,N_6887,N_6865);
xor U9096 (N_9096,N_7345,N_7284);
or U9097 (N_9097,N_7259,N_7140);
and U9098 (N_9098,N_7996,N_6215);
xor U9099 (N_9099,N_7621,N_7224);
nor U9100 (N_9100,N_6026,N_6979);
nand U9101 (N_9101,N_6792,N_7947);
and U9102 (N_9102,N_6878,N_6307);
xnor U9103 (N_9103,N_7211,N_6569);
nor U9104 (N_9104,N_7146,N_7793);
or U9105 (N_9105,N_6562,N_6747);
and U9106 (N_9106,N_7940,N_6394);
and U9107 (N_9107,N_6243,N_7421);
nor U9108 (N_9108,N_6198,N_7842);
nand U9109 (N_9109,N_6401,N_7868);
nor U9110 (N_9110,N_6557,N_6085);
or U9111 (N_9111,N_7883,N_6799);
and U9112 (N_9112,N_7519,N_7623);
or U9113 (N_9113,N_6409,N_7129);
nand U9114 (N_9114,N_6297,N_7650);
and U9115 (N_9115,N_7026,N_7391);
nor U9116 (N_9116,N_6202,N_7726);
nor U9117 (N_9117,N_6570,N_7363);
nor U9118 (N_9118,N_6243,N_6805);
nor U9119 (N_9119,N_6218,N_6488);
or U9120 (N_9120,N_7594,N_6544);
nand U9121 (N_9121,N_7161,N_7668);
nand U9122 (N_9122,N_7479,N_7636);
or U9123 (N_9123,N_6402,N_6198);
xnor U9124 (N_9124,N_6701,N_7326);
or U9125 (N_9125,N_6704,N_7265);
xnor U9126 (N_9126,N_6863,N_6442);
nor U9127 (N_9127,N_7931,N_7887);
nor U9128 (N_9128,N_7132,N_6993);
nor U9129 (N_9129,N_7681,N_6572);
or U9130 (N_9130,N_7034,N_7903);
and U9131 (N_9131,N_6767,N_7860);
and U9132 (N_9132,N_6102,N_6584);
or U9133 (N_9133,N_6807,N_6732);
nand U9134 (N_9134,N_7050,N_7922);
nand U9135 (N_9135,N_7473,N_6172);
and U9136 (N_9136,N_7505,N_6585);
nor U9137 (N_9137,N_7909,N_6202);
or U9138 (N_9138,N_7036,N_6611);
nor U9139 (N_9139,N_7583,N_7972);
or U9140 (N_9140,N_7951,N_6157);
nand U9141 (N_9141,N_7157,N_6309);
or U9142 (N_9142,N_7961,N_7557);
nand U9143 (N_9143,N_7275,N_6581);
and U9144 (N_9144,N_7997,N_7423);
nand U9145 (N_9145,N_7360,N_6816);
and U9146 (N_9146,N_7355,N_6580);
nor U9147 (N_9147,N_6774,N_7003);
nand U9148 (N_9148,N_7154,N_7603);
xnor U9149 (N_9149,N_6080,N_7543);
or U9150 (N_9150,N_6437,N_7440);
nor U9151 (N_9151,N_6841,N_6860);
nand U9152 (N_9152,N_6685,N_7213);
or U9153 (N_9153,N_7037,N_6114);
nand U9154 (N_9154,N_7653,N_6598);
nand U9155 (N_9155,N_6563,N_7513);
nand U9156 (N_9156,N_7856,N_6602);
and U9157 (N_9157,N_6652,N_6701);
xnor U9158 (N_9158,N_6886,N_7642);
xor U9159 (N_9159,N_6722,N_7776);
xnor U9160 (N_9160,N_6936,N_7794);
nand U9161 (N_9161,N_6739,N_6451);
and U9162 (N_9162,N_6168,N_6218);
nand U9163 (N_9163,N_6207,N_6601);
nor U9164 (N_9164,N_7982,N_7425);
nand U9165 (N_9165,N_7388,N_6590);
and U9166 (N_9166,N_7631,N_7414);
xnor U9167 (N_9167,N_7772,N_6977);
nor U9168 (N_9168,N_7887,N_7065);
nor U9169 (N_9169,N_7048,N_7199);
nand U9170 (N_9170,N_7631,N_6326);
or U9171 (N_9171,N_6398,N_6145);
nand U9172 (N_9172,N_7928,N_6556);
nand U9173 (N_9173,N_7876,N_7781);
nor U9174 (N_9174,N_6007,N_6053);
nand U9175 (N_9175,N_7031,N_7670);
nor U9176 (N_9176,N_7365,N_6519);
xnor U9177 (N_9177,N_7606,N_7979);
or U9178 (N_9178,N_6946,N_7463);
and U9179 (N_9179,N_6644,N_7813);
nor U9180 (N_9180,N_6417,N_7041);
nor U9181 (N_9181,N_6070,N_7013);
and U9182 (N_9182,N_6433,N_6118);
and U9183 (N_9183,N_6287,N_6894);
and U9184 (N_9184,N_7105,N_6518);
and U9185 (N_9185,N_6283,N_6317);
or U9186 (N_9186,N_7382,N_6775);
nor U9187 (N_9187,N_6670,N_6200);
nor U9188 (N_9188,N_7715,N_6507);
and U9189 (N_9189,N_7264,N_6631);
nor U9190 (N_9190,N_7114,N_6788);
or U9191 (N_9191,N_7955,N_6165);
or U9192 (N_9192,N_6247,N_7323);
and U9193 (N_9193,N_6162,N_7969);
and U9194 (N_9194,N_6040,N_6321);
xor U9195 (N_9195,N_7884,N_6055);
and U9196 (N_9196,N_6332,N_6697);
nor U9197 (N_9197,N_6870,N_6388);
and U9198 (N_9198,N_7230,N_7337);
nand U9199 (N_9199,N_7633,N_6303);
or U9200 (N_9200,N_6092,N_7174);
nor U9201 (N_9201,N_7051,N_6359);
nor U9202 (N_9202,N_7187,N_6258);
nand U9203 (N_9203,N_7146,N_7376);
xor U9204 (N_9204,N_7628,N_7119);
nand U9205 (N_9205,N_6023,N_6056);
nor U9206 (N_9206,N_6631,N_6854);
and U9207 (N_9207,N_7303,N_6961);
and U9208 (N_9208,N_6149,N_6116);
and U9209 (N_9209,N_7203,N_7264);
xnor U9210 (N_9210,N_6160,N_7230);
nor U9211 (N_9211,N_7034,N_7511);
and U9212 (N_9212,N_7120,N_7640);
nor U9213 (N_9213,N_6285,N_7895);
nand U9214 (N_9214,N_7167,N_7065);
and U9215 (N_9215,N_6942,N_6547);
or U9216 (N_9216,N_6379,N_7231);
nand U9217 (N_9217,N_6970,N_6383);
or U9218 (N_9218,N_7398,N_6007);
nor U9219 (N_9219,N_7070,N_6843);
and U9220 (N_9220,N_7145,N_6137);
and U9221 (N_9221,N_6915,N_6856);
nand U9222 (N_9222,N_6307,N_7171);
or U9223 (N_9223,N_6433,N_7573);
and U9224 (N_9224,N_7699,N_6319);
or U9225 (N_9225,N_6459,N_7798);
nand U9226 (N_9226,N_6597,N_6896);
and U9227 (N_9227,N_7934,N_6255);
or U9228 (N_9228,N_7893,N_6305);
nand U9229 (N_9229,N_7023,N_7660);
nor U9230 (N_9230,N_7074,N_7115);
or U9231 (N_9231,N_7589,N_6912);
nor U9232 (N_9232,N_7475,N_6357);
nand U9233 (N_9233,N_7287,N_7841);
and U9234 (N_9234,N_7625,N_6852);
and U9235 (N_9235,N_7606,N_6474);
or U9236 (N_9236,N_6155,N_6023);
nor U9237 (N_9237,N_7670,N_7698);
nor U9238 (N_9238,N_6113,N_7640);
or U9239 (N_9239,N_7580,N_6847);
or U9240 (N_9240,N_7121,N_6316);
nand U9241 (N_9241,N_7873,N_7833);
or U9242 (N_9242,N_6192,N_6273);
nand U9243 (N_9243,N_6187,N_7106);
or U9244 (N_9244,N_6208,N_7597);
or U9245 (N_9245,N_7634,N_7572);
nand U9246 (N_9246,N_7412,N_6046);
or U9247 (N_9247,N_7571,N_6483);
nor U9248 (N_9248,N_6569,N_6979);
or U9249 (N_9249,N_7989,N_7877);
and U9250 (N_9250,N_7918,N_6161);
and U9251 (N_9251,N_7203,N_7508);
nor U9252 (N_9252,N_6914,N_6572);
and U9253 (N_9253,N_7808,N_6412);
nand U9254 (N_9254,N_7939,N_7387);
nor U9255 (N_9255,N_6113,N_6723);
xor U9256 (N_9256,N_7706,N_7404);
nor U9257 (N_9257,N_6832,N_7690);
nor U9258 (N_9258,N_7508,N_6559);
nor U9259 (N_9259,N_7439,N_6397);
and U9260 (N_9260,N_6784,N_6087);
nand U9261 (N_9261,N_7700,N_7393);
and U9262 (N_9262,N_6171,N_6525);
xnor U9263 (N_9263,N_6678,N_6509);
and U9264 (N_9264,N_7833,N_7096);
nor U9265 (N_9265,N_6371,N_7560);
or U9266 (N_9266,N_6935,N_7083);
xor U9267 (N_9267,N_7574,N_7403);
and U9268 (N_9268,N_7060,N_6653);
nand U9269 (N_9269,N_6513,N_6288);
nor U9270 (N_9270,N_7179,N_6626);
nor U9271 (N_9271,N_6106,N_7614);
xnor U9272 (N_9272,N_6794,N_6369);
nand U9273 (N_9273,N_7942,N_7209);
xor U9274 (N_9274,N_7908,N_7473);
and U9275 (N_9275,N_6367,N_6730);
nor U9276 (N_9276,N_7511,N_7042);
and U9277 (N_9277,N_6577,N_6158);
nor U9278 (N_9278,N_7306,N_7851);
nand U9279 (N_9279,N_6800,N_7122);
or U9280 (N_9280,N_6681,N_7094);
nor U9281 (N_9281,N_6885,N_7346);
nand U9282 (N_9282,N_7618,N_6554);
nor U9283 (N_9283,N_7996,N_6369);
nor U9284 (N_9284,N_7911,N_7009);
or U9285 (N_9285,N_7830,N_7099);
nand U9286 (N_9286,N_6285,N_7991);
nand U9287 (N_9287,N_7876,N_6368);
nor U9288 (N_9288,N_6663,N_7604);
nand U9289 (N_9289,N_6597,N_6522);
and U9290 (N_9290,N_6873,N_6965);
nor U9291 (N_9291,N_6976,N_6402);
and U9292 (N_9292,N_7318,N_7421);
or U9293 (N_9293,N_6987,N_6039);
and U9294 (N_9294,N_6451,N_6833);
and U9295 (N_9295,N_6966,N_6768);
and U9296 (N_9296,N_6088,N_6403);
nand U9297 (N_9297,N_6496,N_7239);
or U9298 (N_9298,N_6647,N_7437);
or U9299 (N_9299,N_7854,N_7362);
or U9300 (N_9300,N_7625,N_6513);
and U9301 (N_9301,N_6884,N_7333);
and U9302 (N_9302,N_7209,N_6974);
nor U9303 (N_9303,N_7456,N_6009);
nor U9304 (N_9304,N_6155,N_6208);
xnor U9305 (N_9305,N_7157,N_6954);
and U9306 (N_9306,N_7709,N_7731);
nor U9307 (N_9307,N_6357,N_6728);
and U9308 (N_9308,N_6656,N_6900);
nand U9309 (N_9309,N_7843,N_6399);
nor U9310 (N_9310,N_7009,N_7472);
and U9311 (N_9311,N_6406,N_7871);
nor U9312 (N_9312,N_7196,N_6509);
nand U9313 (N_9313,N_6698,N_6910);
nor U9314 (N_9314,N_7355,N_6429);
nor U9315 (N_9315,N_6864,N_7883);
and U9316 (N_9316,N_6909,N_6789);
and U9317 (N_9317,N_6538,N_7609);
or U9318 (N_9318,N_7315,N_6045);
nand U9319 (N_9319,N_6099,N_7034);
nand U9320 (N_9320,N_7232,N_6406);
and U9321 (N_9321,N_6861,N_7474);
xor U9322 (N_9322,N_7945,N_6002);
xnor U9323 (N_9323,N_7840,N_7359);
nor U9324 (N_9324,N_7958,N_6099);
xor U9325 (N_9325,N_7667,N_6605);
and U9326 (N_9326,N_6250,N_7378);
or U9327 (N_9327,N_6469,N_6127);
or U9328 (N_9328,N_7382,N_7017);
and U9329 (N_9329,N_6840,N_6836);
and U9330 (N_9330,N_6709,N_7137);
or U9331 (N_9331,N_6982,N_6745);
and U9332 (N_9332,N_6469,N_6447);
nand U9333 (N_9333,N_6128,N_7097);
nand U9334 (N_9334,N_7046,N_7211);
xor U9335 (N_9335,N_7892,N_6603);
nor U9336 (N_9336,N_7606,N_6106);
or U9337 (N_9337,N_6741,N_7808);
or U9338 (N_9338,N_6531,N_6441);
nand U9339 (N_9339,N_6440,N_7136);
nor U9340 (N_9340,N_6219,N_7653);
xnor U9341 (N_9341,N_6358,N_7641);
nor U9342 (N_9342,N_7008,N_6051);
nand U9343 (N_9343,N_6568,N_6571);
nand U9344 (N_9344,N_6177,N_6398);
nand U9345 (N_9345,N_6605,N_7121);
and U9346 (N_9346,N_7251,N_7839);
nor U9347 (N_9347,N_6678,N_6088);
xor U9348 (N_9348,N_7109,N_6438);
and U9349 (N_9349,N_7608,N_6202);
nor U9350 (N_9350,N_7108,N_6685);
or U9351 (N_9351,N_7244,N_6982);
or U9352 (N_9352,N_6464,N_7547);
or U9353 (N_9353,N_7814,N_6080);
and U9354 (N_9354,N_6484,N_7272);
or U9355 (N_9355,N_6479,N_6098);
nor U9356 (N_9356,N_7025,N_6560);
nor U9357 (N_9357,N_7921,N_6986);
nand U9358 (N_9358,N_7204,N_7796);
nand U9359 (N_9359,N_6517,N_7623);
nand U9360 (N_9360,N_7058,N_7279);
nor U9361 (N_9361,N_7218,N_6209);
and U9362 (N_9362,N_6974,N_7957);
and U9363 (N_9363,N_6257,N_7510);
and U9364 (N_9364,N_7216,N_6393);
nor U9365 (N_9365,N_6775,N_6706);
and U9366 (N_9366,N_7059,N_6003);
nand U9367 (N_9367,N_6704,N_7293);
xnor U9368 (N_9368,N_7906,N_7448);
and U9369 (N_9369,N_6308,N_7009);
xnor U9370 (N_9370,N_6708,N_6970);
and U9371 (N_9371,N_7920,N_6835);
or U9372 (N_9372,N_7341,N_7324);
or U9373 (N_9373,N_6160,N_6829);
nand U9374 (N_9374,N_7400,N_6518);
nand U9375 (N_9375,N_6538,N_6373);
or U9376 (N_9376,N_6905,N_7421);
nor U9377 (N_9377,N_6889,N_7862);
or U9378 (N_9378,N_6508,N_6165);
xnor U9379 (N_9379,N_7096,N_6636);
xor U9380 (N_9380,N_6103,N_6430);
or U9381 (N_9381,N_6503,N_7746);
nor U9382 (N_9382,N_6320,N_7383);
nor U9383 (N_9383,N_7430,N_6674);
nand U9384 (N_9384,N_7660,N_7464);
and U9385 (N_9385,N_6637,N_6607);
nor U9386 (N_9386,N_6563,N_6979);
or U9387 (N_9387,N_7376,N_7880);
and U9388 (N_9388,N_6415,N_7839);
nand U9389 (N_9389,N_7148,N_7957);
and U9390 (N_9390,N_6602,N_6515);
xor U9391 (N_9391,N_6526,N_7869);
and U9392 (N_9392,N_7987,N_6546);
xor U9393 (N_9393,N_6500,N_6502);
nor U9394 (N_9394,N_7757,N_7585);
and U9395 (N_9395,N_7319,N_7768);
nand U9396 (N_9396,N_6853,N_7237);
nand U9397 (N_9397,N_7845,N_7463);
and U9398 (N_9398,N_6262,N_7170);
nor U9399 (N_9399,N_6315,N_6726);
or U9400 (N_9400,N_7129,N_7435);
or U9401 (N_9401,N_6278,N_6513);
and U9402 (N_9402,N_7070,N_6851);
nand U9403 (N_9403,N_6000,N_6389);
and U9404 (N_9404,N_6300,N_7756);
nor U9405 (N_9405,N_7307,N_7997);
and U9406 (N_9406,N_6133,N_6510);
nand U9407 (N_9407,N_6044,N_6853);
xor U9408 (N_9408,N_6356,N_7977);
or U9409 (N_9409,N_6825,N_7593);
and U9410 (N_9410,N_6844,N_7319);
nor U9411 (N_9411,N_6725,N_6253);
nor U9412 (N_9412,N_7766,N_7667);
or U9413 (N_9413,N_6045,N_6199);
nand U9414 (N_9414,N_6802,N_6297);
and U9415 (N_9415,N_7050,N_7684);
and U9416 (N_9416,N_6195,N_6240);
nand U9417 (N_9417,N_6716,N_6917);
or U9418 (N_9418,N_6298,N_7042);
nand U9419 (N_9419,N_7926,N_6482);
or U9420 (N_9420,N_7553,N_6434);
or U9421 (N_9421,N_7096,N_6935);
nor U9422 (N_9422,N_7416,N_7117);
nor U9423 (N_9423,N_6677,N_7723);
nand U9424 (N_9424,N_6622,N_6707);
and U9425 (N_9425,N_6151,N_6068);
nand U9426 (N_9426,N_6193,N_6492);
or U9427 (N_9427,N_7213,N_6037);
nand U9428 (N_9428,N_7467,N_7786);
nor U9429 (N_9429,N_7558,N_6856);
nand U9430 (N_9430,N_7263,N_6173);
nor U9431 (N_9431,N_7226,N_6512);
nor U9432 (N_9432,N_7385,N_7548);
nor U9433 (N_9433,N_7692,N_7233);
or U9434 (N_9434,N_7678,N_7094);
nor U9435 (N_9435,N_7923,N_7173);
nor U9436 (N_9436,N_6841,N_7347);
and U9437 (N_9437,N_7158,N_7937);
or U9438 (N_9438,N_7956,N_7464);
or U9439 (N_9439,N_7297,N_6266);
nand U9440 (N_9440,N_7380,N_7676);
nand U9441 (N_9441,N_7708,N_6543);
and U9442 (N_9442,N_7723,N_7057);
nor U9443 (N_9443,N_6994,N_7621);
xnor U9444 (N_9444,N_6852,N_7170);
nor U9445 (N_9445,N_7301,N_6023);
nor U9446 (N_9446,N_7771,N_7107);
and U9447 (N_9447,N_7779,N_7296);
or U9448 (N_9448,N_6867,N_6748);
or U9449 (N_9449,N_6061,N_6210);
nor U9450 (N_9450,N_6630,N_7183);
or U9451 (N_9451,N_6770,N_6311);
and U9452 (N_9452,N_7752,N_6978);
xnor U9453 (N_9453,N_6112,N_7235);
xnor U9454 (N_9454,N_6591,N_7464);
nand U9455 (N_9455,N_7919,N_6897);
nor U9456 (N_9456,N_7756,N_6369);
and U9457 (N_9457,N_6760,N_7089);
nor U9458 (N_9458,N_6031,N_7288);
nor U9459 (N_9459,N_6336,N_7890);
xnor U9460 (N_9460,N_7515,N_6709);
nand U9461 (N_9461,N_6463,N_7425);
nor U9462 (N_9462,N_7664,N_6710);
nand U9463 (N_9463,N_7317,N_7361);
nand U9464 (N_9464,N_6601,N_7022);
and U9465 (N_9465,N_6198,N_6771);
and U9466 (N_9466,N_7095,N_7409);
or U9467 (N_9467,N_7528,N_7383);
nor U9468 (N_9468,N_7492,N_7930);
nand U9469 (N_9469,N_6093,N_6567);
and U9470 (N_9470,N_7855,N_6151);
and U9471 (N_9471,N_6738,N_6420);
nor U9472 (N_9472,N_6312,N_7668);
or U9473 (N_9473,N_7626,N_7532);
nor U9474 (N_9474,N_7969,N_6715);
nand U9475 (N_9475,N_6158,N_6458);
nand U9476 (N_9476,N_7801,N_6576);
nand U9477 (N_9477,N_7441,N_7869);
xnor U9478 (N_9478,N_6832,N_6257);
and U9479 (N_9479,N_6348,N_6799);
nor U9480 (N_9480,N_7660,N_7612);
and U9481 (N_9481,N_6645,N_6046);
and U9482 (N_9482,N_7690,N_7826);
nor U9483 (N_9483,N_7316,N_6246);
or U9484 (N_9484,N_6172,N_6382);
or U9485 (N_9485,N_6216,N_7126);
and U9486 (N_9486,N_7555,N_6208);
and U9487 (N_9487,N_7046,N_7436);
nand U9488 (N_9488,N_6755,N_6295);
nor U9489 (N_9489,N_7021,N_7535);
nand U9490 (N_9490,N_7407,N_6215);
nor U9491 (N_9491,N_6855,N_6326);
nor U9492 (N_9492,N_7211,N_6065);
and U9493 (N_9493,N_7341,N_6893);
nor U9494 (N_9494,N_6917,N_7922);
or U9495 (N_9495,N_7906,N_7483);
nor U9496 (N_9496,N_6334,N_7426);
nand U9497 (N_9497,N_6191,N_6350);
nand U9498 (N_9498,N_7235,N_6260);
or U9499 (N_9499,N_7593,N_6591);
nor U9500 (N_9500,N_7523,N_6392);
and U9501 (N_9501,N_7844,N_7649);
nand U9502 (N_9502,N_6702,N_7257);
nor U9503 (N_9503,N_6052,N_7039);
nand U9504 (N_9504,N_6831,N_6717);
nand U9505 (N_9505,N_6780,N_6145);
nand U9506 (N_9506,N_6451,N_6243);
or U9507 (N_9507,N_6538,N_6223);
nand U9508 (N_9508,N_7263,N_6192);
or U9509 (N_9509,N_6927,N_7400);
or U9510 (N_9510,N_7556,N_7933);
nor U9511 (N_9511,N_6340,N_7604);
nor U9512 (N_9512,N_6566,N_7339);
and U9513 (N_9513,N_7970,N_6800);
or U9514 (N_9514,N_6785,N_6820);
and U9515 (N_9515,N_7374,N_6363);
or U9516 (N_9516,N_7471,N_7624);
and U9517 (N_9517,N_6058,N_6696);
and U9518 (N_9518,N_7705,N_7951);
or U9519 (N_9519,N_7200,N_6490);
nor U9520 (N_9520,N_7350,N_7112);
and U9521 (N_9521,N_7530,N_7700);
and U9522 (N_9522,N_6235,N_6198);
nor U9523 (N_9523,N_6739,N_6756);
nand U9524 (N_9524,N_6146,N_7487);
and U9525 (N_9525,N_6121,N_6078);
or U9526 (N_9526,N_7170,N_6410);
nor U9527 (N_9527,N_7527,N_6339);
nor U9528 (N_9528,N_7942,N_6938);
and U9529 (N_9529,N_7443,N_6323);
and U9530 (N_9530,N_7374,N_7449);
nor U9531 (N_9531,N_7399,N_6415);
and U9532 (N_9532,N_6648,N_7586);
nor U9533 (N_9533,N_7438,N_6310);
and U9534 (N_9534,N_7855,N_7776);
nand U9535 (N_9535,N_7962,N_6398);
nor U9536 (N_9536,N_7741,N_7903);
and U9537 (N_9537,N_6949,N_7244);
and U9538 (N_9538,N_6059,N_6843);
or U9539 (N_9539,N_7032,N_6392);
nor U9540 (N_9540,N_6025,N_7312);
or U9541 (N_9541,N_6221,N_7189);
or U9542 (N_9542,N_6450,N_6319);
xor U9543 (N_9543,N_6367,N_7164);
or U9544 (N_9544,N_7043,N_6385);
nand U9545 (N_9545,N_7226,N_7174);
nor U9546 (N_9546,N_6754,N_7715);
and U9547 (N_9547,N_7486,N_7510);
nand U9548 (N_9548,N_6823,N_6859);
nor U9549 (N_9549,N_6071,N_6920);
nor U9550 (N_9550,N_7127,N_7782);
and U9551 (N_9551,N_7098,N_7049);
and U9552 (N_9552,N_7219,N_6269);
xor U9553 (N_9553,N_7181,N_7250);
and U9554 (N_9554,N_7315,N_6034);
nor U9555 (N_9555,N_7436,N_7471);
or U9556 (N_9556,N_6779,N_6548);
or U9557 (N_9557,N_6894,N_7428);
nor U9558 (N_9558,N_6121,N_6605);
nand U9559 (N_9559,N_6246,N_7664);
or U9560 (N_9560,N_6614,N_6242);
xor U9561 (N_9561,N_6209,N_6287);
or U9562 (N_9562,N_6013,N_6029);
and U9563 (N_9563,N_7039,N_7220);
and U9564 (N_9564,N_6915,N_7370);
and U9565 (N_9565,N_6037,N_6498);
nor U9566 (N_9566,N_6937,N_7897);
nor U9567 (N_9567,N_6119,N_7700);
nand U9568 (N_9568,N_6183,N_7178);
or U9569 (N_9569,N_7641,N_6653);
and U9570 (N_9570,N_7881,N_6334);
nor U9571 (N_9571,N_6642,N_6774);
nand U9572 (N_9572,N_6167,N_7358);
xor U9573 (N_9573,N_6921,N_7489);
nor U9574 (N_9574,N_6512,N_7032);
nor U9575 (N_9575,N_7583,N_6781);
nand U9576 (N_9576,N_7442,N_7899);
xor U9577 (N_9577,N_6969,N_6355);
and U9578 (N_9578,N_6019,N_7749);
xnor U9579 (N_9579,N_7011,N_7440);
nand U9580 (N_9580,N_7773,N_7727);
and U9581 (N_9581,N_6881,N_6818);
nand U9582 (N_9582,N_7228,N_6205);
nor U9583 (N_9583,N_7000,N_7697);
and U9584 (N_9584,N_7819,N_6103);
nand U9585 (N_9585,N_7745,N_7885);
or U9586 (N_9586,N_6826,N_6834);
or U9587 (N_9587,N_7199,N_7635);
nor U9588 (N_9588,N_6132,N_7427);
and U9589 (N_9589,N_7564,N_6577);
and U9590 (N_9590,N_6282,N_6967);
nor U9591 (N_9591,N_6633,N_6201);
and U9592 (N_9592,N_6314,N_7293);
nor U9593 (N_9593,N_7005,N_7792);
and U9594 (N_9594,N_6755,N_6042);
xor U9595 (N_9595,N_6048,N_7242);
nor U9596 (N_9596,N_7726,N_7972);
nor U9597 (N_9597,N_7080,N_6868);
or U9598 (N_9598,N_6226,N_6011);
and U9599 (N_9599,N_7612,N_6092);
and U9600 (N_9600,N_7830,N_7841);
and U9601 (N_9601,N_6502,N_7460);
nand U9602 (N_9602,N_6391,N_6091);
or U9603 (N_9603,N_7676,N_7304);
and U9604 (N_9604,N_6767,N_7649);
or U9605 (N_9605,N_7176,N_7709);
nand U9606 (N_9606,N_7787,N_7029);
or U9607 (N_9607,N_6140,N_6398);
xnor U9608 (N_9608,N_7139,N_6796);
xnor U9609 (N_9609,N_6024,N_6941);
or U9610 (N_9610,N_7499,N_6310);
or U9611 (N_9611,N_6853,N_7595);
nor U9612 (N_9612,N_7390,N_6708);
or U9613 (N_9613,N_7830,N_7237);
or U9614 (N_9614,N_7528,N_6843);
nand U9615 (N_9615,N_6595,N_6511);
or U9616 (N_9616,N_6894,N_7014);
nand U9617 (N_9617,N_6759,N_7644);
nor U9618 (N_9618,N_6046,N_6432);
nand U9619 (N_9619,N_7406,N_6056);
xnor U9620 (N_9620,N_6911,N_7885);
or U9621 (N_9621,N_7090,N_7535);
xor U9622 (N_9622,N_7373,N_7102);
nand U9623 (N_9623,N_7034,N_7536);
and U9624 (N_9624,N_6919,N_7484);
xnor U9625 (N_9625,N_6062,N_6409);
and U9626 (N_9626,N_7496,N_6547);
nor U9627 (N_9627,N_6878,N_6933);
nand U9628 (N_9628,N_6856,N_7612);
or U9629 (N_9629,N_7220,N_7795);
or U9630 (N_9630,N_7971,N_7850);
nand U9631 (N_9631,N_7837,N_6423);
and U9632 (N_9632,N_6532,N_7549);
and U9633 (N_9633,N_6361,N_7614);
nor U9634 (N_9634,N_7189,N_7384);
nor U9635 (N_9635,N_7802,N_7654);
nor U9636 (N_9636,N_6466,N_7977);
xor U9637 (N_9637,N_6548,N_7418);
xor U9638 (N_9638,N_6891,N_7417);
nand U9639 (N_9639,N_7376,N_7269);
or U9640 (N_9640,N_7267,N_6122);
xor U9641 (N_9641,N_7154,N_7861);
or U9642 (N_9642,N_6204,N_7281);
xnor U9643 (N_9643,N_7474,N_6878);
nand U9644 (N_9644,N_7465,N_6725);
nand U9645 (N_9645,N_7725,N_6954);
nor U9646 (N_9646,N_6088,N_7615);
and U9647 (N_9647,N_7260,N_7965);
nand U9648 (N_9648,N_6834,N_7872);
nor U9649 (N_9649,N_6250,N_6094);
or U9650 (N_9650,N_6496,N_6844);
or U9651 (N_9651,N_6482,N_6089);
and U9652 (N_9652,N_7215,N_6818);
nand U9653 (N_9653,N_7804,N_6519);
nand U9654 (N_9654,N_6594,N_7135);
or U9655 (N_9655,N_7483,N_7951);
nand U9656 (N_9656,N_6910,N_7159);
nand U9657 (N_9657,N_6304,N_7069);
or U9658 (N_9658,N_6188,N_7891);
and U9659 (N_9659,N_6499,N_7618);
nor U9660 (N_9660,N_6231,N_7175);
xnor U9661 (N_9661,N_7506,N_7808);
nor U9662 (N_9662,N_7487,N_6030);
nand U9663 (N_9663,N_7332,N_6824);
nor U9664 (N_9664,N_6212,N_7988);
and U9665 (N_9665,N_6431,N_7354);
and U9666 (N_9666,N_6552,N_7182);
nor U9667 (N_9667,N_7122,N_7263);
nor U9668 (N_9668,N_6351,N_7010);
nand U9669 (N_9669,N_6363,N_7600);
or U9670 (N_9670,N_6690,N_7570);
nand U9671 (N_9671,N_7336,N_6191);
or U9672 (N_9672,N_6053,N_7309);
and U9673 (N_9673,N_7588,N_7984);
nand U9674 (N_9674,N_7608,N_7512);
nand U9675 (N_9675,N_6216,N_6275);
nand U9676 (N_9676,N_7522,N_7289);
nor U9677 (N_9677,N_7235,N_7796);
or U9678 (N_9678,N_7468,N_6870);
nor U9679 (N_9679,N_6557,N_6165);
and U9680 (N_9680,N_7912,N_6495);
nand U9681 (N_9681,N_6968,N_7601);
nor U9682 (N_9682,N_7597,N_7103);
and U9683 (N_9683,N_7398,N_6734);
xor U9684 (N_9684,N_6906,N_7580);
nor U9685 (N_9685,N_6782,N_6444);
or U9686 (N_9686,N_7583,N_7604);
and U9687 (N_9687,N_7566,N_7217);
and U9688 (N_9688,N_6399,N_6489);
nor U9689 (N_9689,N_7940,N_6632);
or U9690 (N_9690,N_7736,N_7397);
and U9691 (N_9691,N_7263,N_6019);
nand U9692 (N_9692,N_6908,N_6329);
or U9693 (N_9693,N_6892,N_7449);
nand U9694 (N_9694,N_7172,N_6854);
nand U9695 (N_9695,N_6594,N_7280);
xor U9696 (N_9696,N_7995,N_7345);
and U9697 (N_9697,N_6963,N_6571);
nand U9698 (N_9698,N_7882,N_7913);
nand U9699 (N_9699,N_6345,N_6567);
and U9700 (N_9700,N_7577,N_7941);
nand U9701 (N_9701,N_7994,N_6677);
and U9702 (N_9702,N_7266,N_7842);
nand U9703 (N_9703,N_7566,N_6066);
nor U9704 (N_9704,N_6193,N_7462);
or U9705 (N_9705,N_6105,N_7592);
nand U9706 (N_9706,N_7471,N_7085);
nand U9707 (N_9707,N_6250,N_7331);
or U9708 (N_9708,N_6388,N_7798);
nand U9709 (N_9709,N_6303,N_6579);
nand U9710 (N_9710,N_7683,N_7783);
nand U9711 (N_9711,N_7906,N_7208);
and U9712 (N_9712,N_6035,N_7227);
nor U9713 (N_9713,N_7354,N_7223);
and U9714 (N_9714,N_7891,N_7903);
and U9715 (N_9715,N_7189,N_7129);
and U9716 (N_9716,N_7880,N_6287);
and U9717 (N_9717,N_6979,N_7295);
and U9718 (N_9718,N_7507,N_7280);
nor U9719 (N_9719,N_7082,N_6304);
or U9720 (N_9720,N_7401,N_6224);
nor U9721 (N_9721,N_7780,N_6015);
xor U9722 (N_9722,N_6322,N_6850);
and U9723 (N_9723,N_7320,N_6013);
and U9724 (N_9724,N_6933,N_6535);
and U9725 (N_9725,N_6534,N_7329);
nor U9726 (N_9726,N_7760,N_6145);
and U9727 (N_9727,N_6433,N_7870);
and U9728 (N_9728,N_6263,N_7840);
and U9729 (N_9729,N_6983,N_7522);
or U9730 (N_9730,N_6717,N_6291);
and U9731 (N_9731,N_7475,N_7244);
and U9732 (N_9732,N_6591,N_7202);
or U9733 (N_9733,N_6259,N_7411);
xnor U9734 (N_9734,N_7169,N_6322);
nor U9735 (N_9735,N_6831,N_7317);
xor U9736 (N_9736,N_7210,N_6349);
and U9737 (N_9737,N_7875,N_7291);
nor U9738 (N_9738,N_7701,N_7783);
nand U9739 (N_9739,N_6455,N_7000);
nor U9740 (N_9740,N_6839,N_7567);
and U9741 (N_9741,N_6253,N_7055);
nand U9742 (N_9742,N_7732,N_7637);
and U9743 (N_9743,N_6484,N_6036);
nor U9744 (N_9744,N_6932,N_7946);
and U9745 (N_9745,N_7503,N_7963);
and U9746 (N_9746,N_7732,N_6655);
nor U9747 (N_9747,N_6676,N_7252);
nand U9748 (N_9748,N_6059,N_7791);
or U9749 (N_9749,N_7512,N_6537);
xor U9750 (N_9750,N_7898,N_7195);
and U9751 (N_9751,N_6646,N_7773);
nand U9752 (N_9752,N_7873,N_6658);
and U9753 (N_9753,N_7541,N_6221);
and U9754 (N_9754,N_7272,N_6308);
or U9755 (N_9755,N_7355,N_7566);
or U9756 (N_9756,N_7375,N_7882);
nand U9757 (N_9757,N_7203,N_6215);
nor U9758 (N_9758,N_7092,N_6698);
nand U9759 (N_9759,N_6459,N_6367);
and U9760 (N_9760,N_6187,N_6806);
xor U9761 (N_9761,N_7026,N_6283);
xor U9762 (N_9762,N_6368,N_7581);
nand U9763 (N_9763,N_7674,N_6839);
or U9764 (N_9764,N_7974,N_7499);
nand U9765 (N_9765,N_6853,N_6627);
or U9766 (N_9766,N_7391,N_7320);
nor U9767 (N_9767,N_6994,N_6000);
and U9768 (N_9768,N_7643,N_6592);
and U9769 (N_9769,N_7287,N_7331);
or U9770 (N_9770,N_6284,N_7836);
and U9771 (N_9771,N_6264,N_7196);
nand U9772 (N_9772,N_6480,N_6569);
nand U9773 (N_9773,N_6639,N_7268);
xnor U9774 (N_9774,N_6200,N_7898);
or U9775 (N_9775,N_7674,N_6855);
and U9776 (N_9776,N_6659,N_7701);
or U9777 (N_9777,N_7668,N_7306);
nor U9778 (N_9778,N_6268,N_6157);
and U9779 (N_9779,N_6042,N_6226);
xnor U9780 (N_9780,N_7684,N_6308);
or U9781 (N_9781,N_6866,N_6583);
or U9782 (N_9782,N_6526,N_6116);
or U9783 (N_9783,N_6642,N_7090);
nor U9784 (N_9784,N_6157,N_7023);
and U9785 (N_9785,N_7142,N_7662);
nand U9786 (N_9786,N_6942,N_7736);
and U9787 (N_9787,N_6557,N_7909);
xnor U9788 (N_9788,N_7308,N_6435);
nor U9789 (N_9789,N_6052,N_6002);
nor U9790 (N_9790,N_7745,N_6702);
nand U9791 (N_9791,N_7952,N_7863);
nand U9792 (N_9792,N_7046,N_6890);
or U9793 (N_9793,N_7495,N_6456);
xnor U9794 (N_9794,N_7097,N_7525);
xnor U9795 (N_9795,N_7220,N_7364);
nor U9796 (N_9796,N_7926,N_7784);
or U9797 (N_9797,N_6627,N_7353);
or U9798 (N_9798,N_7595,N_7147);
xor U9799 (N_9799,N_6706,N_7830);
and U9800 (N_9800,N_7020,N_7661);
nand U9801 (N_9801,N_7371,N_6456);
nand U9802 (N_9802,N_6765,N_6821);
and U9803 (N_9803,N_7969,N_7596);
nand U9804 (N_9804,N_6173,N_6728);
nor U9805 (N_9805,N_7252,N_7783);
or U9806 (N_9806,N_7802,N_6374);
and U9807 (N_9807,N_6045,N_7740);
nand U9808 (N_9808,N_6901,N_6186);
nand U9809 (N_9809,N_6633,N_7062);
nand U9810 (N_9810,N_7879,N_6499);
and U9811 (N_9811,N_7246,N_6639);
or U9812 (N_9812,N_7483,N_6355);
and U9813 (N_9813,N_7174,N_6774);
nand U9814 (N_9814,N_6941,N_6059);
and U9815 (N_9815,N_7731,N_7280);
nand U9816 (N_9816,N_6846,N_7568);
xor U9817 (N_9817,N_6728,N_6116);
and U9818 (N_9818,N_6553,N_7050);
and U9819 (N_9819,N_6289,N_6550);
nor U9820 (N_9820,N_6877,N_7562);
nor U9821 (N_9821,N_6230,N_6466);
nor U9822 (N_9822,N_6231,N_6107);
nand U9823 (N_9823,N_7092,N_7930);
and U9824 (N_9824,N_6736,N_7344);
xor U9825 (N_9825,N_7219,N_6485);
or U9826 (N_9826,N_7921,N_7394);
nand U9827 (N_9827,N_7215,N_6058);
and U9828 (N_9828,N_6414,N_7288);
nor U9829 (N_9829,N_6264,N_6000);
and U9830 (N_9830,N_7802,N_6898);
nor U9831 (N_9831,N_7965,N_7814);
nand U9832 (N_9832,N_7750,N_6531);
and U9833 (N_9833,N_6563,N_7245);
or U9834 (N_9834,N_6322,N_7089);
or U9835 (N_9835,N_6732,N_7726);
nor U9836 (N_9836,N_6971,N_6400);
xnor U9837 (N_9837,N_7029,N_6131);
and U9838 (N_9838,N_7776,N_7539);
or U9839 (N_9839,N_7614,N_7901);
and U9840 (N_9840,N_6926,N_6620);
or U9841 (N_9841,N_6731,N_7839);
or U9842 (N_9842,N_7606,N_7232);
nor U9843 (N_9843,N_7091,N_7509);
nand U9844 (N_9844,N_6911,N_6413);
nand U9845 (N_9845,N_6039,N_7264);
or U9846 (N_9846,N_6692,N_7147);
or U9847 (N_9847,N_7821,N_7088);
xnor U9848 (N_9848,N_6092,N_6946);
or U9849 (N_9849,N_6418,N_6996);
nand U9850 (N_9850,N_7306,N_6432);
or U9851 (N_9851,N_6322,N_7969);
and U9852 (N_9852,N_6982,N_6234);
and U9853 (N_9853,N_7948,N_6888);
nand U9854 (N_9854,N_6233,N_6384);
or U9855 (N_9855,N_6341,N_6688);
and U9856 (N_9856,N_7998,N_7680);
and U9857 (N_9857,N_7130,N_6889);
nand U9858 (N_9858,N_6416,N_6596);
nor U9859 (N_9859,N_7131,N_6517);
xor U9860 (N_9860,N_7026,N_6861);
nor U9861 (N_9861,N_7236,N_6705);
and U9862 (N_9862,N_6319,N_6105);
nand U9863 (N_9863,N_6821,N_6323);
nand U9864 (N_9864,N_7593,N_6635);
nand U9865 (N_9865,N_6820,N_7093);
nand U9866 (N_9866,N_6722,N_7757);
nand U9867 (N_9867,N_6231,N_6437);
xnor U9868 (N_9868,N_7658,N_7305);
and U9869 (N_9869,N_7732,N_6408);
nand U9870 (N_9870,N_6439,N_7464);
or U9871 (N_9871,N_7913,N_6547);
nand U9872 (N_9872,N_7928,N_6453);
nand U9873 (N_9873,N_6244,N_6733);
nand U9874 (N_9874,N_7122,N_6000);
nor U9875 (N_9875,N_6549,N_7158);
and U9876 (N_9876,N_7714,N_6308);
nor U9877 (N_9877,N_7595,N_6196);
xor U9878 (N_9878,N_7718,N_7160);
nand U9879 (N_9879,N_7530,N_7891);
and U9880 (N_9880,N_7649,N_6595);
or U9881 (N_9881,N_6075,N_6399);
nor U9882 (N_9882,N_7487,N_7296);
and U9883 (N_9883,N_7698,N_7823);
xnor U9884 (N_9884,N_6279,N_7679);
nand U9885 (N_9885,N_7752,N_7369);
or U9886 (N_9886,N_7913,N_6425);
and U9887 (N_9887,N_6197,N_7528);
or U9888 (N_9888,N_6568,N_6687);
xnor U9889 (N_9889,N_6720,N_7231);
or U9890 (N_9890,N_6687,N_6512);
nand U9891 (N_9891,N_7688,N_7043);
nand U9892 (N_9892,N_6016,N_6129);
or U9893 (N_9893,N_7638,N_7942);
xnor U9894 (N_9894,N_7592,N_6733);
nor U9895 (N_9895,N_6805,N_6928);
or U9896 (N_9896,N_7840,N_7943);
or U9897 (N_9897,N_7547,N_7929);
or U9898 (N_9898,N_7046,N_7809);
nand U9899 (N_9899,N_7168,N_7915);
or U9900 (N_9900,N_7143,N_7026);
nand U9901 (N_9901,N_7811,N_7451);
nor U9902 (N_9902,N_6227,N_6746);
or U9903 (N_9903,N_7631,N_6263);
nand U9904 (N_9904,N_6892,N_6107);
and U9905 (N_9905,N_6455,N_7958);
nor U9906 (N_9906,N_6230,N_6679);
nand U9907 (N_9907,N_7634,N_7115);
and U9908 (N_9908,N_7620,N_7538);
and U9909 (N_9909,N_7325,N_7953);
and U9910 (N_9910,N_6998,N_7698);
or U9911 (N_9911,N_7655,N_6431);
nand U9912 (N_9912,N_7629,N_6775);
nor U9913 (N_9913,N_7249,N_6367);
or U9914 (N_9914,N_6991,N_6066);
nor U9915 (N_9915,N_7071,N_7716);
or U9916 (N_9916,N_7037,N_7267);
nor U9917 (N_9917,N_7057,N_6529);
xnor U9918 (N_9918,N_7870,N_6111);
or U9919 (N_9919,N_7231,N_6217);
nor U9920 (N_9920,N_6638,N_6130);
xor U9921 (N_9921,N_6552,N_6101);
nand U9922 (N_9922,N_7245,N_7717);
xnor U9923 (N_9923,N_6758,N_7940);
nand U9924 (N_9924,N_7250,N_7248);
and U9925 (N_9925,N_7401,N_6652);
nor U9926 (N_9926,N_6580,N_6275);
or U9927 (N_9927,N_6066,N_7276);
nor U9928 (N_9928,N_6974,N_7904);
nand U9929 (N_9929,N_7607,N_7480);
nand U9930 (N_9930,N_6457,N_7474);
and U9931 (N_9931,N_6303,N_6021);
nand U9932 (N_9932,N_7721,N_6221);
and U9933 (N_9933,N_6351,N_7854);
and U9934 (N_9934,N_6859,N_7636);
nor U9935 (N_9935,N_6402,N_7186);
nand U9936 (N_9936,N_6711,N_6652);
nor U9937 (N_9937,N_6038,N_7613);
nor U9938 (N_9938,N_7607,N_6419);
nand U9939 (N_9939,N_6992,N_7972);
or U9940 (N_9940,N_6382,N_7629);
nand U9941 (N_9941,N_6558,N_7068);
nor U9942 (N_9942,N_6074,N_6698);
xor U9943 (N_9943,N_7356,N_6400);
nand U9944 (N_9944,N_7150,N_7290);
and U9945 (N_9945,N_7984,N_6812);
or U9946 (N_9946,N_7839,N_7135);
nor U9947 (N_9947,N_7787,N_7934);
and U9948 (N_9948,N_6398,N_6457);
or U9949 (N_9949,N_7145,N_7259);
or U9950 (N_9950,N_6850,N_7582);
xnor U9951 (N_9951,N_7930,N_7605);
nand U9952 (N_9952,N_7622,N_7573);
xor U9953 (N_9953,N_6185,N_6811);
and U9954 (N_9954,N_7053,N_7743);
and U9955 (N_9955,N_6448,N_6593);
nand U9956 (N_9956,N_7436,N_6296);
nor U9957 (N_9957,N_6169,N_7383);
or U9958 (N_9958,N_6536,N_7803);
and U9959 (N_9959,N_7706,N_7646);
nor U9960 (N_9960,N_7361,N_7396);
and U9961 (N_9961,N_6253,N_7187);
and U9962 (N_9962,N_6149,N_6820);
and U9963 (N_9963,N_7852,N_6706);
and U9964 (N_9964,N_7922,N_7641);
and U9965 (N_9965,N_6102,N_6332);
and U9966 (N_9966,N_7129,N_7359);
nand U9967 (N_9967,N_7156,N_7568);
or U9968 (N_9968,N_7524,N_7598);
nor U9969 (N_9969,N_7964,N_6664);
and U9970 (N_9970,N_6162,N_7857);
nor U9971 (N_9971,N_6417,N_6883);
nand U9972 (N_9972,N_7992,N_7674);
xnor U9973 (N_9973,N_6158,N_7378);
xnor U9974 (N_9974,N_7561,N_6086);
nand U9975 (N_9975,N_6759,N_6589);
and U9976 (N_9976,N_6072,N_7804);
nor U9977 (N_9977,N_6777,N_6949);
nand U9978 (N_9978,N_6651,N_7673);
nand U9979 (N_9979,N_6238,N_7394);
or U9980 (N_9980,N_6532,N_7116);
nor U9981 (N_9981,N_6288,N_6311);
xnor U9982 (N_9982,N_6927,N_6796);
and U9983 (N_9983,N_7792,N_7143);
and U9984 (N_9984,N_6159,N_6352);
nor U9985 (N_9985,N_7229,N_7674);
nand U9986 (N_9986,N_7858,N_7518);
or U9987 (N_9987,N_7333,N_6115);
and U9988 (N_9988,N_6964,N_7081);
nand U9989 (N_9989,N_7626,N_6508);
nor U9990 (N_9990,N_7902,N_6342);
xor U9991 (N_9991,N_6125,N_6935);
nor U9992 (N_9992,N_7632,N_6983);
or U9993 (N_9993,N_7689,N_6798);
or U9994 (N_9994,N_7146,N_7937);
and U9995 (N_9995,N_7003,N_6290);
nor U9996 (N_9996,N_7004,N_7959);
and U9997 (N_9997,N_6419,N_7998);
and U9998 (N_9998,N_6827,N_7250);
and U9999 (N_9999,N_6821,N_7102);
and UO_0 (O_0,N_9288,N_8153);
or UO_1 (O_1,N_8526,N_9644);
and UO_2 (O_2,N_8572,N_9699);
nor UO_3 (O_3,N_8422,N_8914);
nand UO_4 (O_4,N_9348,N_9322);
nor UO_5 (O_5,N_9344,N_9289);
nor UO_6 (O_6,N_9793,N_9251);
nand UO_7 (O_7,N_8977,N_9214);
or UO_8 (O_8,N_8658,N_8403);
and UO_9 (O_9,N_9201,N_9719);
nor UO_10 (O_10,N_8240,N_8864);
nand UO_11 (O_11,N_8932,N_9698);
and UO_12 (O_12,N_9525,N_8035);
or UO_13 (O_13,N_9126,N_8648);
and UO_14 (O_14,N_8005,N_8262);
nor UO_15 (O_15,N_8909,N_9890);
or UO_16 (O_16,N_8399,N_8043);
xor UO_17 (O_17,N_8647,N_9390);
and UO_18 (O_18,N_9562,N_9114);
and UO_19 (O_19,N_9277,N_9173);
nor UO_20 (O_20,N_9224,N_9824);
and UO_21 (O_21,N_9522,N_8432);
or UO_22 (O_22,N_9257,N_8782);
and UO_23 (O_23,N_8509,N_9885);
nand UO_24 (O_24,N_9785,N_9483);
and UO_25 (O_25,N_9294,N_8118);
xnor UO_26 (O_26,N_8050,N_8385);
nand UO_27 (O_27,N_8349,N_9051);
and UO_28 (O_28,N_9789,N_8607);
xor UO_29 (O_29,N_8675,N_9714);
xor UO_30 (O_30,N_8789,N_8311);
nor UO_31 (O_31,N_9758,N_8042);
nand UO_32 (O_32,N_9843,N_9551);
and UO_33 (O_33,N_8373,N_9420);
and UO_34 (O_34,N_9371,N_8443);
nand UO_35 (O_35,N_9549,N_9981);
and UO_36 (O_36,N_8824,N_8508);
or UO_37 (O_37,N_9211,N_8205);
nor UO_38 (O_38,N_8455,N_9672);
nand UO_39 (O_39,N_8172,N_8820);
nand UO_40 (O_40,N_8740,N_8702);
and UO_41 (O_41,N_9668,N_8783);
nor UO_42 (O_42,N_8748,N_8960);
or UO_43 (O_43,N_8485,N_9689);
and UO_44 (O_44,N_8558,N_8733);
nor UO_45 (O_45,N_9134,N_9248);
or UO_46 (O_46,N_9107,N_9231);
nand UO_47 (O_47,N_8278,N_8414);
nor UO_48 (O_48,N_9537,N_9260);
nor UO_49 (O_49,N_8696,N_8053);
nand UO_50 (O_50,N_8954,N_8706);
and UO_51 (O_51,N_9169,N_8668);
nand UO_52 (O_52,N_8464,N_8430);
nand UO_53 (O_53,N_8014,N_9599);
or UO_54 (O_54,N_9777,N_9882);
nand UO_55 (O_55,N_8468,N_8060);
or UO_56 (O_56,N_8232,N_8612);
nor UO_57 (O_57,N_8528,N_9956);
and UO_58 (O_58,N_8319,N_9536);
or UO_59 (O_59,N_8291,N_8540);
nand UO_60 (O_60,N_8860,N_9364);
xor UO_61 (O_61,N_8189,N_9190);
nor UO_62 (O_62,N_8774,N_9189);
nand UO_63 (O_63,N_9094,N_9113);
and UO_64 (O_64,N_8229,N_9615);
or UO_65 (O_65,N_9786,N_9013);
and UO_66 (O_66,N_9399,N_8109);
or UO_67 (O_67,N_9220,N_8133);
or UO_68 (O_68,N_9040,N_8877);
xnor UO_69 (O_69,N_8370,N_9186);
or UO_70 (O_70,N_9593,N_9269);
nor UO_71 (O_71,N_8110,N_9716);
nor UO_72 (O_72,N_9850,N_8339);
or UO_73 (O_73,N_9193,N_8603);
nor UO_74 (O_74,N_9521,N_9939);
nand UO_75 (O_75,N_9185,N_8452);
or UO_76 (O_76,N_8124,N_9391);
and UO_77 (O_77,N_9676,N_8701);
xnor UO_78 (O_78,N_9572,N_9524);
nor UO_79 (O_79,N_9250,N_8300);
nand UO_80 (O_80,N_8889,N_9662);
and UO_81 (O_81,N_9389,N_9147);
xor UO_82 (O_82,N_9516,N_9367);
and UO_83 (O_83,N_9639,N_8428);
xnor UO_84 (O_84,N_9519,N_8975);
nand UO_85 (O_85,N_9280,N_8047);
nor UO_86 (O_86,N_8259,N_9314);
or UO_87 (O_87,N_8011,N_9424);
or UO_88 (O_88,N_9089,N_9069);
xnor UO_89 (O_89,N_8841,N_8524);
nand UO_90 (O_90,N_9433,N_8352);
and UO_91 (O_91,N_8930,N_8358);
xnor UO_92 (O_92,N_8688,N_9947);
or UO_93 (O_93,N_9818,N_9988);
nand UO_94 (O_94,N_8722,N_8515);
nor UO_95 (O_95,N_9654,N_8188);
or UO_96 (O_96,N_8672,N_8199);
or UO_97 (O_97,N_9049,N_9290);
and UO_98 (O_98,N_9255,N_8923);
nand UO_99 (O_99,N_8654,N_8628);
and UO_100 (O_100,N_8169,N_9197);
or UO_101 (O_101,N_9271,N_9310);
and UO_102 (O_102,N_8096,N_9642);
or UO_103 (O_103,N_9479,N_9959);
nand UO_104 (O_104,N_8423,N_8828);
and UO_105 (O_105,N_8384,N_8671);
xor UO_106 (O_106,N_8201,N_9972);
nor UO_107 (O_107,N_9973,N_9106);
and UO_108 (O_108,N_9552,N_9452);
and UO_109 (O_109,N_9831,N_9416);
or UO_110 (O_110,N_8168,N_9962);
nor UO_111 (O_111,N_9858,N_8447);
xnor UO_112 (O_112,N_8900,N_8966);
xor UO_113 (O_113,N_8116,N_8719);
or UO_114 (O_114,N_9340,N_9088);
or UO_115 (O_115,N_9902,N_8411);
xnor UO_116 (O_116,N_9209,N_9307);
nor UO_117 (O_117,N_9635,N_8197);
and UO_118 (O_118,N_8367,N_8602);
and UO_119 (O_119,N_8313,N_9688);
nand UO_120 (O_120,N_8910,N_9118);
xor UO_121 (O_121,N_9218,N_9653);
or UO_122 (O_122,N_9547,N_8532);
nor UO_123 (O_123,N_9619,N_9243);
or UO_124 (O_124,N_8167,N_9741);
or UO_125 (O_125,N_8646,N_9206);
or UO_126 (O_126,N_8185,N_8217);
or UO_127 (O_127,N_8834,N_8017);
nor UO_128 (O_128,N_9481,N_8788);
nand UO_129 (O_129,N_9496,N_9148);
nor UO_130 (O_130,N_9993,N_9323);
and UO_131 (O_131,N_8863,N_8965);
nand UO_132 (O_132,N_9281,N_9345);
or UO_133 (O_133,N_8953,N_8204);
and UO_134 (O_134,N_8737,N_8606);
nor UO_135 (O_135,N_9679,N_9868);
nor UO_136 (O_136,N_8697,N_8323);
nor UO_137 (O_137,N_8107,N_9019);
nor UO_138 (O_138,N_8350,N_9916);
nor UO_139 (O_139,N_8996,N_9665);
or UO_140 (O_140,N_8459,N_9841);
xnor UO_141 (O_141,N_8878,N_8861);
or UO_142 (O_142,N_9394,N_9335);
xor UO_143 (O_143,N_9187,N_8446);
nand UO_144 (O_144,N_9991,N_9435);
xnor UO_145 (O_145,N_8955,N_9752);
or UO_146 (O_146,N_8937,N_9620);
and UO_147 (O_147,N_8813,N_8377);
or UO_148 (O_148,N_8374,N_9410);
nand UO_149 (O_149,N_9707,N_9244);
xnor UO_150 (O_150,N_8234,N_9283);
nor UO_151 (O_151,N_8770,N_8186);
xor UO_152 (O_152,N_9640,N_9630);
and UO_153 (O_153,N_9191,N_8145);
nand UO_154 (O_154,N_8699,N_8771);
and UO_155 (O_155,N_9397,N_9184);
nor UO_156 (O_156,N_9784,N_9880);
and UO_157 (O_157,N_9965,N_9103);
or UO_158 (O_158,N_9807,N_8280);
nand UO_159 (O_159,N_9188,N_8454);
nor UO_160 (O_160,N_9131,N_8985);
xor UO_161 (O_161,N_8974,N_9120);
nand UO_162 (O_162,N_8191,N_8933);
nand UO_163 (O_163,N_8308,N_9154);
or UO_164 (O_164,N_8518,N_9379);
nand UO_165 (O_165,N_8080,N_8661);
nor UO_166 (O_166,N_8255,N_8048);
nand UO_167 (O_167,N_8195,N_9819);
nor UO_168 (O_168,N_9770,N_9393);
or UO_169 (O_169,N_8979,N_8390);
and UO_170 (O_170,N_9001,N_9948);
nand UO_171 (O_171,N_9427,N_8296);
or UO_172 (O_172,N_9465,N_8488);
or UO_173 (O_173,N_8839,N_9862);
nor UO_174 (O_174,N_8173,N_8335);
nor UO_175 (O_175,N_8533,N_9775);
xor UO_176 (O_176,N_9750,N_8198);
nand UO_177 (O_177,N_8180,N_8761);
and UO_178 (O_178,N_8148,N_9208);
and UO_179 (O_179,N_8806,N_9171);
nor UO_180 (O_180,N_9327,N_9337);
nand UO_181 (O_181,N_9164,N_9631);
xnor UO_182 (O_182,N_9007,N_8898);
nor UO_183 (O_183,N_9086,N_9279);
nor UO_184 (O_184,N_9594,N_9495);
nor UO_185 (O_185,N_8193,N_8821);
nand UO_186 (O_186,N_9157,N_9702);
and UO_187 (O_187,N_8665,N_9272);
nand UO_188 (O_188,N_8567,N_8678);
or UO_189 (O_189,N_8024,N_8721);
or UO_190 (O_190,N_8298,N_8075);
nor UO_191 (O_191,N_9505,N_9766);
nor UO_192 (O_192,N_8091,N_8010);
or UO_193 (O_193,N_8995,N_9937);
or UO_194 (O_194,N_9167,N_8579);
and UO_195 (O_195,N_9783,N_8496);
nand UO_196 (O_196,N_9837,N_8183);
or UO_197 (O_197,N_8704,N_8474);
and UO_198 (O_198,N_9942,N_9478);
or UO_199 (O_199,N_9733,N_9330);
and UO_200 (O_200,N_9268,N_8416);
and UO_201 (O_201,N_9267,N_9133);
nand UO_202 (O_202,N_8857,N_9697);
nand UO_203 (O_203,N_9744,N_8246);
nor UO_204 (O_204,N_8487,N_8907);
nor UO_205 (O_205,N_9041,N_8948);
or UO_206 (O_206,N_9027,N_9712);
nand UO_207 (O_207,N_8969,N_8559);
and UO_208 (O_208,N_9934,N_8064);
and UO_209 (O_209,N_8584,N_9558);
or UO_210 (O_210,N_9413,N_9998);
nand UO_211 (O_211,N_9825,N_9002);
and UO_212 (O_212,N_8429,N_8751);
nor UO_213 (O_213,N_9808,N_9905);
nor UO_214 (O_214,N_9043,N_8775);
xnor UO_215 (O_215,N_9334,N_8745);
and UO_216 (O_216,N_9542,N_9256);
nand UO_217 (O_217,N_8420,N_8245);
nand UO_218 (O_218,N_8758,N_9974);
or UO_219 (O_219,N_8354,N_9550);
and UO_220 (O_220,N_9501,N_8303);
and UO_221 (O_221,N_9961,N_8547);
nor UO_222 (O_222,N_9720,N_9008);
or UO_223 (O_223,N_8715,N_8777);
nor UO_224 (O_224,N_9781,N_8548);
nor UO_225 (O_225,N_9840,N_8981);
nor UO_226 (O_226,N_8796,N_8651);
nor UO_227 (O_227,N_8970,N_8176);
and UO_228 (O_228,N_8326,N_8638);
or UO_229 (O_229,N_8275,N_9317);
or UO_230 (O_230,N_9477,N_8967);
nor UO_231 (O_231,N_9347,N_8155);
nor UO_232 (O_232,N_8780,N_8644);
nor UO_233 (O_233,N_8036,N_9643);
and UO_234 (O_234,N_9155,N_8781);
nor UO_235 (O_235,N_9212,N_9772);
and UO_236 (O_236,N_8211,N_9102);
and UO_237 (O_237,N_8460,N_9346);
and UO_238 (O_238,N_9451,N_9233);
nor UO_239 (O_239,N_9616,N_9431);
xnor UO_240 (O_240,N_8227,N_8674);
xor UO_241 (O_241,N_8426,N_8505);
or UO_242 (O_242,N_9830,N_9940);
nand UO_243 (O_243,N_8750,N_9930);
xor UO_244 (O_244,N_8263,N_8545);
nor UO_245 (O_245,N_8670,N_9152);
nand UO_246 (O_246,N_9403,N_8884);
or UO_247 (O_247,N_8818,N_9755);
and UO_248 (O_248,N_8112,N_8887);
or UO_249 (O_249,N_8146,N_9357);
and UO_250 (O_250,N_8226,N_9358);
or UO_251 (O_251,N_9046,N_8497);
or UO_252 (O_252,N_9030,N_8874);
or UO_253 (O_253,N_9070,N_9048);
or UO_254 (O_254,N_8944,N_9513);
nor UO_255 (O_255,N_9661,N_9897);
nand UO_256 (O_256,N_8015,N_9667);
or UO_257 (O_257,N_8698,N_8886);
nor UO_258 (O_258,N_9731,N_8541);
nand UO_259 (O_259,N_8842,N_8534);
xnor UO_260 (O_260,N_9645,N_9901);
nor UO_261 (O_261,N_8272,N_9449);
nand UO_262 (O_262,N_9865,N_9836);
nor UO_263 (O_263,N_9514,N_8565);
nand UO_264 (O_264,N_8480,N_8382);
and UO_265 (O_265,N_9162,N_9045);
nand UO_266 (O_266,N_9320,N_9907);
nand UO_267 (O_267,N_8649,N_9464);
or UO_268 (O_268,N_8165,N_9135);
and UO_269 (O_269,N_8516,N_9215);
xnor UO_270 (O_270,N_9530,N_8158);
xor UO_271 (O_271,N_8802,N_8825);
nand UO_272 (O_272,N_9943,N_9761);
or UO_273 (O_273,N_8406,N_9273);
xnor UO_274 (O_274,N_8279,N_8580);
nand UO_275 (O_275,N_8277,N_9338);
or UO_276 (O_276,N_8962,N_9471);
and UO_277 (O_277,N_9617,N_9020);
nor UO_278 (O_278,N_8461,N_8623);
and UO_279 (O_279,N_9691,N_9904);
nand UO_280 (O_280,N_8355,N_8589);
nor UO_281 (O_281,N_8233,N_8504);
xnor UO_282 (O_282,N_8888,N_9318);
or UO_283 (O_283,N_8137,N_9618);
and UO_284 (O_284,N_8103,N_8493);
and UO_285 (O_285,N_8164,N_9278);
nor UO_286 (O_286,N_9084,N_8987);
xor UO_287 (O_287,N_8971,N_9609);
nand UO_288 (O_288,N_9075,N_9129);
xor UO_289 (O_289,N_8248,N_9743);
nor UO_290 (O_290,N_9474,N_8968);
nand UO_291 (O_291,N_8475,N_8576);
nand UO_292 (O_292,N_8586,N_9475);
or UO_293 (O_293,N_8097,N_9502);
nor UO_294 (O_294,N_9034,N_9098);
nor UO_295 (O_295,N_9237,N_8935);
or UO_296 (O_296,N_8293,N_9829);
and UO_297 (O_297,N_8436,N_9459);
and UO_298 (O_298,N_8465,N_9816);
or UO_299 (O_299,N_9886,N_9871);
nand UO_300 (O_300,N_9342,N_9764);
xor UO_301 (O_301,N_8902,N_8182);
or UO_302 (O_302,N_8098,N_8827);
and UO_303 (O_303,N_8144,N_8848);
nand UO_304 (O_304,N_9485,N_8312);
and UO_305 (O_305,N_9795,N_9655);
or UO_306 (O_306,N_9166,N_9832);
and UO_307 (O_307,N_8331,N_9466);
nor UO_308 (O_308,N_9658,N_9887);
and UO_309 (O_309,N_9174,N_8650);
and UO_310 (O_310,N_8982,N_9706);
nor UO_311 (O_311,N_9490,N_9963);
nand UO_312 (O_312,N_8592,N_9026);
xor UO_313 (O_313,N_9161,N_9261);
nand UO_314 (O_314,N_9983,N_9095);
xnor UO_315 (O_315,N_9685,N_9238);
or UO_316 (O_316,N_8727,N_9374);
xnor UO_317 (O_317,N_9690,N_8639);
and UO_318 (O_318,N_8921,N_9753);
and UO_319 (O_319,N_9627,N_9299);
nor UO_320 (O_320,N_8617,N_8194);
nor UO_321 (O_321,N_9455,N_8510);
nand UO_322 (O_322,N_9553,N_9589);
and UO_323 (O_323,N_9091,N_9366);
or UO_324 (O_324,N_8852,N_9535);
nand UO_325 (O_325,N_8997,N_9610);
and UO_326 (O_326,N_8574,N_8637);
nand UO_327 (O_327,N_8387,N_8682);
and UO_328 (O_328,N_9732,N_9092);
or UO_329 (O_329,N_9739,N_9557);
xnor UO_330 (O_330,N_8081,N_8484);
or UO_331 (O_331,N_9180,N_8143);
or UO_332 (O_332,N_8787,N_9035);
and UO_333 (O_333,N_8090,N_9175);
and UO_334 (O_334,N_9857,N_9176);
nand UO_335 (O_335,N_9442,N_9112);
nor UO_336 (O_336,N_8254,N_9870);
and UO_337 (O_337,N_8845,N_8892);
and UO_338 (O_338,N_8045,N_8330);
nand UO_339 (O_339,N_8258,N_9486);
nor UO_340 (O_340,N_8742,N_9022);
nand UO_341 (O_341,N_8066,N_8713);
xor UO_342 (O_342,N_8826,N_9867);
and UO_343 (O_343,N_9899,N_8028);
xor UO_344 (O_344,N_8993,N_9422);
and UO_345 (O_345,N_9274,N_9849);
and UO_346 (O_346,N_8597,N_8285);
nand UO_347 (O_347,N_8336,N_8378);
nand UO_348 (O_348,N_8271,N_9361);
nor UO_349 (O_349,N_8673,N_8433);
nor UO_350 (O_350,N_8040,N_8571);
nand UO_351 (O_351,N_8166,N_9587);
or UO_352 (O_352,N_8223,N_8221);
or UO_353 (O_353,N_8926,N_8837);
and UO_354 (O_354,N_9623,N_9968);
nand UO_355 (O_355,N_8551,N_8256);
nand UO_356 (O_356,N_8341,N_9898);
nor UO_357 (O_357,N_9159,N_8306);
and UO_358 (O_358,N_8814,N_8209);
nor UO_359 (O_359,N_8079,N_9407);
nand UO_360 (O_360,N_8924,N_9497);
and UO_361 (O_361,N_9855,N_9468);
or UO_362 (O_362,N_9710,N_9458);
nor UO_363 (O_363,N_8049,N_8832);
xnor UO_364 (O_364,N_8618,N_9062);
nand UO_365 (O_365,N_9139,N_8244);
and UO_366 (O_366,N_9554,N_9597);
nand UO_367 (O_367,N_8718,N_9848);
or UO_368 (O_368,N_9421,N_9177);
and UO_369 (O_369,N_9834,N_9052);
nand UO_370 (O_370,N_9511,N_8490);
xnor UO_371 (O_371,N_8407,N_8723);
nand UO_372 (O_372,N_9097,N_8113);
and UO_373 (O_373,N_8598,N_8642);
nor UO_374 (O_374,N_9590,N_8287);
nor UO_375 (O_375,N_8250,N_9298);
and UO_376 (O_376,N_9293,N_8557);
or UO_377 (O_377,N_8401,N_8667);
or UO_378 (O_378,N_9326,N_9602);
nand UO_379 (O_379,N_9765,N_9456);
nand UO_380 (O_380,N_8252,N_9009);
nand UO_381 (O_381,N_9994,N_9463);
nand UO_382 (O_382,N_9295,N_8089);
nand UO_383 (O_383,N_8539,N_8179);
nor UO_384 (O_384,N_9145,N_9194);
nor UO_385 (O_385,N_8905,N_8320);
and UO_386 (O_386,N_9055,N_8694);
and UO_387 (O_387,N_8599,N_8561);
xor UO_388 (O_388,N_8396,N_8734);
or UO_389 (O_389,N_9977,N_8421);
nor UO_390 (O_390,N_9156,N_9810);
xor UO_391 (O_391,N_8177,N_8726);
and UO_392 (O_392,N_8769,N_9520);
xnor UO_393 (O_393,N_9003,N_8409);
or UO_394 (O_394,N_8322,N_9723);
nor UO_395 (O_395,N_9059,N_9881);
or UO_396 (O_396,N_8685,N_9343);
nand UO_397 (O_397,N_8983,N_9432);
and UO_398 (O_398,N_9878,N_9406);
and UO_399 (O_399,N_8922,N_9674);
or UO_400 (O_400,N_9523,N_9499);
nor UO_401 (O_401,N_8419,N_9812);
nor UO_402 (O_402,N_9512,N_9598);
or UO_403 (O_403,N_8450,N_8425);
xnor UO_404 (O_404,N_8073,N_9503);
or UO_405 (O_405,N_9078,N_9760);
xnor UO_406 (O_406,N_8989,N_8276);
or UO_407 (O_407,N_8427,N_8101);
nor UO_408 (O_408,N_9779,N_9817);
and UO_409 (O_409,N_8945,N_9437);
and UO_410 (O_410,N_9138,N_9312);
and UO_411 (O_411,N_8855,N_9259);
nor UO_412 (O_412,N_8791,N_8395);
xnor UO_413 (O_413,N_9384,N_8417);
or UO_414 (O_414,N_8546,N_8805);
nor UO_415 (O_415,N_8316,N_9105);
or UO_416 (O_416,N_8635,N_9747);
or UO_417 (O_417,N_9262,N_9083);
xnor UO_418 (O_418,N_8865,N_9877);
or UO_419 (O_419,N_9087,N_9382);
nand UO_420 (O_420,N_9773,N_9104);
nand UO_421 (O_421,N_8264,N_8778);
nand UO_422 (O_422,N_8947,N_9757);
or UO_423 (O_423,N_8867,N_9718);
xor UO_424 (O_424,N_8513,N_9494);
and UO_425 (O_425,N_9683,N_9143);
or UO_426 (O_426,N_9359,N_8624);
or UO_427 (O_427,N_9680,N_8560);
nor UO_428 (O_428,N_8315,N_8008);
or UO_429 (O_429,N_8307,N_9869);
and UO_430 (O_430,N_8283,N_8793);
or UO_431 (O_431,N_8030,N_8919);
nand UO_432 (O_432,N_8086,N_9136);
or UO_433 (O_433,N_9595,N_8006);
nor UO_434 (O_434,N_8732,N_8691);
and UO_435 (O_435,N_8479,N_8249);
xnor UO_436 (O_436,N_8705,N_9412);
and UO_437 (O_437,N_8573,N_9879);
or UO_438 (O_438,N_8174,N_9225);
nor UO_439 (O_439,N_8512,N_9660);
xor UO_440 (O_440,N_9090,N_8913);
nor UO_441 (O_441,N_9356,N_9797);
or UO_442 (O_442,N_8822,N_9856);
nor UO_443 (O_443,N_9787,N_8261);
or UO_444 (O_444,N_9081,N_8949);
or UO_445 (O_445,N_8178,N_8340);
xor UO_446 (O_446,N_9592,N_8297);
and UO_447 (O_447,N_8640,N_8876);
nor UO_448 (O_448,N_8056,N_9309);
or UO_449 (O_449,N_8896,N_8938);
nor UO_450 (O_450,N_8032,N_9398);
nand UO_451 (O_451,N_9540,N_9227);
nand UO_452 (O_452,N_8140,N_9555);
and UO_453 (O_453,N_9971,N_9603);
and UO_454 (O_454,N_8104,N_8629);
and UO_455 (O_455,N_9014,N_9264);
xor UO_456 (O_456,N_9332,N_8866);
nor UO_457 (O_457,N_9058,N_9839);
nor UO_458 (O_458,N_8973,N_8520);
or UO_459 (O_459,N_9626,N_9050);
or UO_460 (O_460,N_9363,N_8676);
or UO_461 (O_461,N_8692,N_8317);
or UO_462 (O_462,N_8984,N_8986);
nor UO_463 (O_463,N_9918,N_9740);
and UO_464 (O_464,N_8716,N_8854);
and UO_465 (O_465,N_9703,N_8018);
and UO_466 (O_466,N_9352,N_8437);
or UO_467 (O_467,N_8556,N_9578);
and UO_468 (O_468,N_9851,N_9895);
or UO_469 (O_469,N_9576,N_9828);
and UO_470 (O_470,N_9713,N_8972);
or UO_471 (O_471,N_8871,N_9923);
nor UO_472 (O_472,N_8940,N_8281);
nand UO_473 (O_473,N_9987,N_8934);
xor UO_474 (O_474,N_8664,N_8441);
and UO_475 (O_475,N_8076,N_8894);
nor UO_476 (O_476,N_8029,N_8615);
nand UO_477 (O_477,N_8767,N_8714);
or UO_478 (O_478,N_9153,N_9791);
nand UO_479 (O_479,N_9109,N_8159);
nor UO_480 (O_480,N_8538,N_9447);
xnor UO_481 (O_481,N_9395,N_8219);
or UO_482 (O_482,N_8500,N_8521);
nand UO_483 (O_483,N_9944,N_9541);
or UO_484 (O_484,N_8568,N_9970);
or UO_485 (O_485,N_8833,N_9246);
nand UO_486 (O_486,N_8868,N_8031);
and UO_487 (O_487,N_9378,N_9803);
or UO_488 (O_488,N_8333,N_8741);
and UO_489 (O_489,N_8305,N_8958);
xor UO_490 (O_490,N_9799,N_9794);
and UO_491 (O_491,N_9024,N_8216);
nand UO_492 (O_492,N_8119,N_9729);
or UO_493 (O_493,N_8327,N_8964);
nand UO_494 (O_494,N_8912,N_8469);
nor UO_495 (O_495,N_8061,N_9771);
nor UO_496 (O_496,N_8879,N_8601);
nor UO_497 (O_497,N_9508,N_8253);
nand UO_498 (O_498,N_9015,N_9538);
nand UO_499 (O_499,N_8077,N_9955);
and UO_500 (O_500,N_9931,N_9517);
or UO_501 (O_501,N_9813,N_8237);
nand UO_502 (O_502,N_8645,N_9360);
nor UO_503 (O_503,N_9100,N_8569);
nor UO_504 (O_504,N_9493,N_8134);
nand UO_505 (O_505,N_8614,N_9845);
or UO_506 (O_506,N_8853,N_9444);
or UO_507 (O_507,N_8756,N_8074);
or UO_508 (O_508,N_9952,N_8106);
nor UO_509 (O_509,N_9756,N_8301);
and UO_510 (O_510,N_8058,N_8368);
and UO_511 (O_511,N_9365,N_8903);
and UO_512 (O_512,N_9920,N_8002);
nand UO_513 (O_513,N_9929,N_8611);
and UO_514 (O_514,N_9085,N_8449);
nand UO_515 (O_515,N_9997,N_8999);
and UO_516 (O_516,N_9158,N_9801);
nor UO_517 (O_517,N_9423,N_9715);
or UO_518 (O_518,N_8364,N_8746);
nor UO_519 (O_519,N_8483,N_9835);
or UO_520 (O_520,N_9454,N_8394);
and UO_521 (O_521,N_9500,N_9232);
nand UO_522 (O_522,N_8759,N_9071);
xnor UO_523 (O_523,N_8404,N_9995);
nor UO_524 (O_524,N_8062,N_8566);
xor UO_525 (O_525,N_8444,N_8711);
nand UO_526 (O_526,N_8383,N_9079);
and UO_527 (O_527,N_9467,N_9652);
nand UO_528 (O_528,N_9472,N_8613);
nand UO_529 (O_529,N_8908,N_9903);
nand UO_530 (O_530,N_9711,N_9182);
and UO_531 (O_531,N_8059,N_8616);
and UO_532 (O_532,N_8957,N_8681);
nand UO_533 (O_533,N_8492,N_9647);
xnor UO_534 (O_534,N_8083,N_8418);
or UO_535 (O_535,N_9605,N_9545);
xnor UO_536 (O_536,N_8517,N_8931);
nand UO_537 (O_537,N_9242,N_9556);
or UO_538 (O_538,N_8361,N_8536);
nand UO_539 (O_539,N_8549,N_9448);
nor UO_540 (O_540,N_8200,N_9596);
or UO_541 (O_541,N_9400,N_8564);
nor UO_542 (O_542,N_8800,N_9217);
and UO_543 (O_543,N_8398,N_9809);
nor UO_544 (O_544,N_9769,N_9915);
nand UO_545 (O_545,N_8632,N_9838);
or UO_546 (O_546,N_9601,N_9144);
nand UO_547 (O_547,N_9815,N_8530);
xor UO_548 (O_548,N_8578,N_9385);
xor UO_549 (O_549,N_9659,N_8491);
nor UO_550 (O_550,N_9032,N_8039);
nand UO_551 (O_551,N_8710,N_9181);
nor UO_552 (O_552,N_8550,N_8481);
and UO_553 (O_553,N_8951,N_9872);
nor UO_554 (O_554,N_8369,N_9434);
nand UO_555 (O_555,N_8380,N_9306);
nand UO_556 (O_556,N_9170,N_8413);
xor UO_557 (O_557,N_8643,N_9945);
nand UO_558 (O_558,N_8215,N_9684);
and UO_559 (O_559,N_8051,N_9969);
or UO_560 (O_560,N_9369,N_9183);
nand UO_561 (O_561,N_8092,N_8859);
and UO_562 (O_562,N_9315,N_8434);
nand UO_563 (O_563,N_9436,N_8511);
and UO_564 (O_564,N_9324,N_9737);
xnor UO_565 (O_565,N_8299,N_9621);
nand UO_566 (O_566,N_8906,N_8055);
nor UO_567 (O_567,N_9012,N_8735);
nor UO_568 (O_568,N_8991,N_8631);
nand UO_569 (O_569,N_8764,N_9386);
and UO_570 (O_570,N_9132,N_9922);
nor UO_571 (O_571,N_9057,N_9806);
and UO_572 (O_572,N_9150,N_8587);
and UO_573 (O_573,N_9328,N_9375);
nor UO_574 (O_574,N_9362,N_9577);
nor UO_575 (O_575,N_9241,N_8212);
nand UO_576 (O_576,N_9563,N_9064);
nor UO_577 (O_577,N_9482,N_8506);
xor UO_578 (O_578,N_9746,N_9568);
nor UO_579 (O_579,N_8070,N_8004);
xnor UO_580 (O_580,N_8356,N_8105);
xnor UO_581 (O_581,N_9297,N_8445);
and UO_582 (O_582,N_8988,N_9873);
or UO_583 (O_583,N_9402,N_8880);
or UO_584 (O_584,N_9473,N_8238);
nor UO_585 (O_585,N_8829,N_9178);
nor UO_586 (O_586,N_8590,N_9287);
nand UO_587 (O_587,N_8994,N_9546);
nor UO_588 (O_588,N_9925,N_8819);
xnor UO_589 (O_589,N_8210,N_9203);
or UO_590 (O_590,N_8284,N_9408);
nor UO_591 (O_591,N_9979,N_9637);
nor UO_592 (O_592,N_9544,N_9584);
or UO_593 (O_593,N_9033,N_9080);
and UO_594 (O_594,N_8529,N_8362);
nor UO_595 (O_595,N_8709,N_8000);
nor UO_596 (O_596,N_9842,N_8023);
nand UO_597 (O_597,N_9179,N_8309);
xnor UO_598 (O_598,N_9792,N_9333);
nand UO_599 (O_599,N_8260,N_9588);
or UO_600 (O_600,N_9125,N_8978);
or UO_601 (O_601,N_8321,N_9504);
and UO_602 (O_602,N_8519,N_9213);
or UO_603 (O_603,N_8171,N_8815);
nor UO_604 (O_604,N_9339,N_9917);
or UO_605 (O_605,N_8156,N_8707);
and UO_606 (O_606,N_8823,N_9060);
nor UO_607 (O_607,N_8743,N_8870);
nand UO_608 (O_608,N_8554,N_9980);
and UO_609 (O_609,N_8858,N_8141);
or UO_610 (O_610,N_9811,N_8680);
and UO_611 (O_611,N_9883,N_8247);
nand UO_612 (O_612,N_9011,N_8728);
nor UO_613 (O_613,N_9528,N_9982);
nand UO_614 (O_614,N_8482,N_8660);
nor UO_615 (O_615,N_8575,N_9429);
nand UO_616 (O_616,N_8034,N_8952);
nand UO_617 (O_617,N_9927,N_9768);
xor UO_618 (O_618,N_9192,N_9263);
and UO_619 (O_619,N_8577,N_8794);
nand UO_620 (O_620,N_9892,N_9219);
xor UO_621 (O_621,N_9717,N_9989);
nor UO_622 (O_622,N_9928,N_9966);
nor UO_623 (O_623,N_9910,N_8862);
nor UO_624 (O_624,N_9908,N_9316);
nand UO_625 (O_625,N_8267,N_8844);
or UO_626 (O_626,N_8739,N_8273);
nand UO_627 (O_627,N_9960,N_9037);
nand UO_628 (O_628,N_9800,N_8736);
nand UO_629 (O_629,N_8928,N_8959);
and UO_630 (O_630,N_9613,N_8304);
nor UO_631 (O_631,N_9790,N_8478);
nand UO_632 (O_632,N_8218,N_8069);
and UO_633 (O_633,N_9669,N_9875);
nand UO_634 (O_634,N_9425,N_9664);
and UO_635 (O_635,N_9958,N_9446);
nand UO_636 (O_636,N_8655,N_8594);
nor UO_637 (O_637,N_9004,N_9383);
nand UO_638 (O_638,N_9253,N_8266);
and UO_639 (O_639,N_8415,N_9580);
or UO_640 (O_640,N_9582,N_9569);
or UO_641 (O_641,N_8149,N_9353);
nand UO_642 (O_642,N_8129,N_9108);
or UO_643 (O_643,N_8916,N_8792);
and UO_644 (O_644,N_8552,N_8605);
or UO_645 (O_645,N_9349,N_8760);
nor UO_646 (O_646,N_9000,N_9571);
or UO_647 (O_647,N_8555,N_9728);
or UO_648 (O_648,N_8208,N_8690);
and UO_649 (O_649,N_9874,N_8899);
nor UO_650 (O_650,N_9321,N_8360);
nor UO_651 (O_651,N_9111,N_8357);
nor UO_652 (O_652,N_9636,N_8738);
and UO_653 (O_653,N_8220,N_9984);
and UO_654 (O_654,N_8181,N_9462);
nor UO_655 (O_655,N_8809,N_9163);
or UO_656 (O_656,N_9565,N_8753);
nor UO_657 (O_657,N_9670,N_8684);
nand UO_658 (O_658,N_9633,N_9319);
nand UO_659 (O_659,N_8634,N_8162);
nand UO_660 (O_660,N_8700,N_8476);
nor UO_661 (O_661,N_8114,N_8626);
nor UO_662 (O_662,N_9415,N_9951);
nor UO_663 (O_663,N_8537,N_8695);
nand UO_664 (O_664,N_8410,N_8009);
nand UO_665 (O_665,N_9844,N_8473);
nor UO_666 (O_666,N_8724,N_9329);
nor UO_667 (O_667,N_9675,N_9561);
nand UO_668 (O_668,N_8462,N_8147);
and UO_669 (O_669,N_8286,N_8448);
nand UO_670 (O_670,N_9198,N_9029);
nor UO_671 (O_671,N_9567,N_9142);
nor UO_672 (O_672,N_8749,N_9205);
or UO_673 (O_673,N_8439,N_9168);
and UO_674 (O_674,N_9301,N_8003);
or UO_675 (O_675,N_8025,N_8228);
xnor UO_676 (O_676,N_9122,N_8583);
nor UO_677 (O_677,N_8812,N_9964);
and UO_678 (O_678,N_8720,N_8393);
nand UO_679 (O_679,N_8747,N_9341);
nor UO_680 (O_680,N_8442,N_8636);
nor UO_681 (O_681,N_9396,N_8608);
or UO_682 (O_682,N_8126,N_8725);
and UO_683 (O_683,N_8033,N_9585);
or UO_684 (O_684,N_9093,N_9247);
and UO_685 (O_685,N_8175,N_9941);
xor UO_686 (O_686,N_8593,N_8257);
and UO_687 (O_687,N_9076,N_8904);
nand UO_688 (O_688,N_9638,N_8525);
nor UO_689 (O_689,N_9823,N_8466);
and UO_690 (O_690,N_8961,N_8604);
and UO_691 (O_691,N_9574,N_9735);
or UO_692 (O_692,N_8499,N_8099);
nor UO_693 (O_693,N_9351,N_9426);
or UO_694 (O_694,N_9734,N_9687);
and UO_695 (O_695,N_8875,N_9641);
or UO_696 (O_696,N_8302,N_8980);
or UO_697 (O_697,N_9629,N_8388);
nor UO_698 (O_698,N_9199,N_8239);
nor UO_699 (O_699,N_9388,N_9210);
nand UO_700 (O_700,N_9117,N_8136);
nor UO_701 (O_701,N_9195,N_9028);
nor UO_702 (O_702,N_9430,N_8345);
and UO_703 (O_703,N_8151,N_8531);
nand UO_704 (O_704,N_8544,N_9047);
or UO_705 (O_705,N_9018,N_8084);
or UO_706 (O_706,N_9957,N_8038);
nor UO_707 (O_707,N_8799,N_9767);
xor UO_708 (O_708,N_9221,N_8094);
and UO_709 (O_709,N_8366,N_8135);
and UO_710 (O_710,N_8895,N_8523);
or UO_711 (O_711,N_8872,N_9861);
nand UO_712 (O_712,N_8405,N_8963);
nand UO_713 (O_713,N_8019,N_8494);
nor UO_714 (O_714,N_8797,N_8027);
nor UO_715 (O_715,N_9373,N_9906);
or UO_716 (O_716,N_8992,N_8342);
nor UO_717 (O_717,N_9607,N_8343);
nand UO_718 (O_718,N_8386,N_9912);
nor UO_719 (O_719,N_8768,N_9796);
and UO_720 (O_720,N_8054,N_9975);
and UO_721 (O_721,N_9063,N_8381);
and UO_722 (O_722,N_9575,N_9978);
nand UO_723 (O_723,N_8881,N_9228);
and UO_724 (O_724,N_9566,N_9053);
and UO_725 (O_725,N_8495,N_9036);
and UO_726 (O_726,N_8893,N_8850);
or UO_727 (O_727,N_9724,N_9996);
or UO_728 (O_728,N_9533,N_8052);
nor UO_729 (O_729,N_9949,N_9222);
or UO_730 (O_730,N_8241,N_9913);
or UO_731 (O_731,N_9450,N_8230);
nor UO_732 (O_732,N_9196,N_9506);
nand UO_733 (O_733,N_8071,N_9266);
nand UO_734 (O_734,N_8939,N_8849);
nor UO_735 (O_735,N_8503,N_8582);
and UO_736 (O_736,N_8917,N_8990);
nand UO_737 (O_737,N_8236,N_8609);
and UO_738 (O_738,N_9119,N_9226);
xor UO_739 (O_739,N_9411,N_8773);
nor UO_740 (O_740,N_8397,N_9066);
and UO_741 (O_741,N_8290,N_8157);
xor UO_742 (O_742,N_9604,N_9709);
xnor UO_743 (O_743,N_8021,N_9909);
or UO_744 (O_744,N_9548,N_8203);
nor UO_745 (O_745,N_8184,N_9254);
xor UO_746 (O_746,N_8542,N_8662);
nand UO_747 (O_747,N_8666,N_8731);
or UO_748 (O_748,N_9727,N_9249);
nand UO_749 (O_749,N_8037,N_8082);
nor UO_750 (O_750,N_9404,N_8585);
and UO_751 (O_751,N_8391,N_9583);
and UO_752 (O_752,N_8095,N_8243);
and UO_753 (O_753,N_9628,N_9286);
nor UO_754 (O_754,N_8915,N_9507);
and UO_755 (O_755,N_8046,N_9999);
and UO_756 (O_756,N_9017,N_9854);
nand UO_757 (O_757,N_9846,N_8348);
nand UO_758 (O_758,N_8652,N_9820);
xor UO_759 (O_759,N_9681,N_8139);
and UO_760 (O_760,N_9762,N_9336);
nor UO_761 (O_761,N_8708,N_8213);
xnor UO_762 (O_762,N_8762,N_9986);
xor UO_763 (O_763,N_8831,N_9387);
or UO_764 (O_764,N_8435,N_9648);
and UO_765 (O_765,N_9579,N_9624);
nor UO_766 (O_766,N_9946,N_9460);
and UO_767 (O_767,N_9682,N_8424);
nor UO_768 (O_768,N_9864,N_9031);
and UO_769 (O_769,N_9414,N_9381);
or UO_770 (O_770,N_8044,N_9077);
or UO_771 (O_771,N_9853,N_9738);
or UO_772 (O_772,N_9742,N_9863);
nor UO_773 (O_773,N_8941,N_9700);
or UO_774 (O_774,N_9586,N_9814);
and UO_775 (O_775,N_9721,N_8679);
nand UO_776 (O_776,N_8457,N_9445);
xnor UO_777 (O_777,N_8507,N_9082);
and UO_778 (O_778,N_9061,N_9671);
or UO_779 (O_779,N_8712,N_8581);
nand UO_780 (O_780,N_9531,N_8231);
or UO_781 (O_781,N_9151,N_9419);
xnor UO_782 (O_782,N_9967,N_8610);
or UO_783 (O_783,N_8772,N_8100);
or UO_784 (O_784,N_8412,N_8808);
or UO_785 (O_785,N_8121,N_8836);
nor UO_786 (O_786,N_8625,N_8078);
and UO_787 (O_787,N_8686,N_8890);
nand UO_788 (O_788,N_9634,N_8653);
nor UO_789 (O_789,N_9476,N_9884);
or UO_790 (O_790,N_8830,N_8752);
nor UO_791 (O_791,N_8744,N_9074);
nand UO_792 (O_792,N_9860,N_9230);
or UO_793 (O_793,N_8160,N_8154);
xnor UO_794 (O_794,N_8235,N_8790);
and UO_795 (O_795,N_9291,N_8472);
and UO_796 (O_796,N_9096,N_8012);
or UO_797 (O_797,N_9116,N_8389);
or UO_798 (O_798,N_9888,N_8132);
or UO_799 (O_799,N_9802,N_9067);
nor UO_800 (O_800,N_9453,N_8998);
and UO_801 (O_801,N_9611,N_9234);
nand UO_802 (O_802,N_8543,N_8196);
or UO_803 (O_803,N_8563,N_8372);
or UO_804 (O_804,N_8379,N_9140);
and UO_805 (O_805,N_9141,N_8108);
or UO_806 (O_806,N_9311,N_9216);
and UO_807 (O_807,N_8122,N_8093);
nand UO_808 (O_808,N_8400,N_9526);
or UO_809 (O_809,N_9488,N_8020);
nor UO_810 (O_810,N_9751,N_8693);
or UO_811 (O_811,N_9701,N_9649);
nand UO_812 (O_812,N_9305,N_9275);
or UO_813 (O_813,N_9774,N_8440);
nor UO_814 (O_814,N_8192,N_9428);
or UO_815 (O_815,N_8630,N_8131);
and UO_816 (O_816,N_9559,N_8622);
xor UO_817 (O_817,N_9896,N_8717);
nor UO_818 (O_818,N_8127,N_9804);
and UO_819 (O_819,N_9149,N_9657);
and UO_820 (O_820,N_9489,N_9470);
nor UO_821 (O_821,N_9518,N_8353);
or UO_822 (O_822,N_9124,N_8225);
or UO_823 (O_823,N_8843,N_9914);
and UO_824 (O_824,N_9759,N_8088);
nor UO_825 (O_825,N_9612,N_9438);
nor UO_826 (O_826,N_9484,N_8656);
nor UO_827 (O_827,N_8477,N_8222);
or UO_828 (O_828,N_8570,N_8486);
and UO_829 (O_829,N_9782,N_8633);
nand UO_830 (O_830,N_8816,N_8785);
or UO_831 (O_831,N_9821,N_8677);
nand UO_832 (O_832,N_8328,N_9304);
or UO_833 (O_833,N_9926,N_8224);
and UO_834 (O_834,N_8463,N_8363);
xor UO_835 (O_835,N_8883,N_8730);
nand UO_836 (O_836,N_8763,N_9704);
nand UO_837 (O_837,N_9532,N_9859);
and UO_838 (O_838,N_8703,N_8334);
or UO_839 (O_839,N_8007,N_8294);
or UO_840 (O_840,N_8801,N_9673);
nand UO_841 (O_841,N_9137,N_9021);
or UO_842 (O_842,N_9663,N_9229);
or UO_843 (O_843,N_9285,N_9068);
nand UO_844 (O_844,N_9992,N_8115);
xnor UO_845 (O_845,N_9694,N_9377);
nor UO_846 (O_846,N_9686,N_9606);
or UO_847 (O_847,N_8351,N_9573);
or UO_848 (O_848,N_9822,N_8501);
nand UO_849 (O_849,N_9172,N_8869);
nand UO_850 (O_850,N_9265,N_9282);
or UO_851 (O_851,N_8251,N_8332);
nor UO_852 (O_852,N_9608,N_9847);
nor UO_853 (O_853,N_8392,N_8057);
xnor UO_854 (O_854,N_8659,N_8142);
nand UO_855 (O_855,N_8187,N_8929);
and UO_856 (O_856,N_8840,N_9876);
nand UO_857 (O_857,N_9270,N_8911);
nor UO_858 (O_858,N_8683,N_8016);
xnor UO_859 (O_859,N_9705,N_9736);
nor UO_860 (O_860,N_9696,N_8620);
nand UO_861 (O_861,N_8338,N_9581);
nor UO_862 (O_862,N_9457,N_8072);
nor UO_863 (O_863,N_8943,N_9976);
nand UO_864 (O_864,N_8438,N_8817);
nor UO_865 (O_865,N_9331,N_8170);
nor UO_866 (O_866,N_8289,N_9491);
nor UO_867 (O_867,N_9591,N_9708);
and UO_868 (O_868,N_8085,N_9776);
nor UO_869 (O_869,N_8669,N_9646);
or UO_870 (O_870,N_8851,N_9921);
xnor UO_871 (O_871,N_9866,N_9204);
and UO_872 (O_872,N_8920,N_8161);
and UO_873 (O_873,N_9677,N_8925);
nor UO_874 (O_874,N_8621,N_8784);
nor UO_875 (O_875,N_8431,N_9745);
and UO_876 (O_876,N_9833,N_8329);
and UO_877 (O_877,N_9101,N_8138);
xor UO_878 (O_878,N_9418,N_8288);
and UO_879 (O_879,N_8041,N_8591);
or UO_880 (O_880,N_8535,N_9016);
nand UO_881 (O_881,N_9110,N_8489);
and UO_882 (O_882,N_8522,N_8754);
or UO_883 (O_883,N_9852,N_9543);
or UO_884 (O_884,N_8514,N_9990);
or UO_885 (O_885,N_9889,N_8214);
nor UO_886 (O_886,N_8891,N_9827);
nand UO_887 (O_887,N_9656,N_9900);
and UO_888 (O_888,N_8295,N_9527);
or UO_889 (O_889,N_8846,N_9240);
nor UO_890 (O_890,N_8856,N_8067);
and UO_891 (O_891,N_8206,N_8950);
xnor UO_892 (O_892,N_9651,N_8269);
and UO_893 (O_893,N_8847,N_8897);
xnor UO_894 (O_894,N_8588,N_8502);
xor UO_895 (O_895,N_8068,N_9202);
or UO_896 (O_896,N_8125,N_8371);
nand UO_897 (O_897,N_8274,N_9236);
or UO_898 (O_898,N_9038,N_8202);
nand UO_899 (O_899,N_8063,N_8111);
and UO_900 (O_900,N_8657,N_9798);
nor UO_901 (O_901,N_8885,N_8314);
nor UO_902 (O_902,N_9726,N_8150);
nor UO_903 (O_903,N_9284,N_9121);
nor UO_904 (O_904,N_9200,N_9722);
xnor UO_905 (O_905,N_8942,N_8689);
or UO_906 (O_906,N_8798,N_9754);
and UO_907 (O_907,N_8779,N_9498);
and UO_908 (O_908,N_9073,N_9950);
xnor UO_909 (O_909,N_9695,N_9480);
nor UO_910 (O_910,N_9005,N_9072);
or UO_911 (O_911,N_8553,N_8270);
nand UO_912 (O_912,N_8346,N_9826);
nand UO_913 (O_913,N_9292,N_9985);
nor UO_914 (O_914,N_8456,N_9749);
nor UO_915 (O_915,N_8595,N_8596);
nand UO_916 (O_916,N_8190,N_8786);
or UO_917 (O_917,N_9778,N_9368);
and UO_918 (O_918,N_9692,N_9010);
nor UO_919 (O_919,N_9146,N_9350);
nor UO_920 (O_920,N_9392,N_9461);
nor UO_921 (O_921,N_9632,N_9302);
nand UO_922 (O_922,N_9044,N_8976);
and UO_923 (O_923,N_8453,N_9308);
nor UO_924 (O_924,N_8663,N_8130);
nand UO_925 (O_925,N_9417,N_9625);
or UO_926 (O_926,N_9469,N_9748);
or UO_927 (O_927,N_8471,N_8755);
and UO_928 (O_928,N_8087,N_8835);
nor UO_929 (O_929,N_9056,N_9529);
nand UO_930 (O_930,N_8776,N_9666);
and UO_931 (O_931,N_9891,N_8458);
nand UO_932 (O_932,N_8268,N_9492);
nand UO_933 (O_933,N_8337,N_8838);
or UO_934 (O_934,N_9355,N_8757);
nor UO_935 (O_935,N_8807,N_9245);
and UO_936 (O_936,N_9935,N_9376);
or UO_937 (O_937,N_9127,N_9953);
and UO_938 (O_938,N_8365,N_8282);
and UO_939 (O_939,N_9042,N_8102);
and UO_940 (O_940,N_8376,N_8152);
nand UO_941 (O_941,N_9239,N_8946);
nand UO_942 (O_942,N_9128,N_8619);
xnor UO_943 (O_943,N_8375,N_9039);
nand UO_944 (O_944,N_9207,N_8765);
or UO_945 (O_945,N_8918,N_9650);
or UO_946 (O_946,N_8562,N_9439);
nand UO_947 (O_947,N_9025,N_9932);
nand UO_948 (O_948,N_9054,N_8359);
xnor UO_949 (O_949,N_8600,N_8344);
or UO_950 (O_950,N_9600,N_9487);
and UO_951 (O_951,N_8687,N_9515);
or UO_952 (O_952,N_9223,N_9401);
nor UO_953 (O_953,N_8927,N_8120);
nor UO_954 (O_954,N_8013,N_9296);
and UO_955 (O_955,N_9165,N_9099);
xor UO_956 (O_956,N_9006,N_9303);
and UO_957 (O_957,N_8347,N_8402);
nor UO_958 (O_958,N_8163,N_9258);
and UO_959 (O_959,N_8292,N_9763);
nand UO_960 (O_960,N_9560,N_9693);
and UO_961 (O_961,N_9534,N_9570);
nor UO_962 (O_962,N_9409,N_9115);
and UO_963 (O_963,N_8318,N_9372);
or UO_964 (O_964,N_9805,N_9276);
nor UO_965 (O_965,N_8956,N_8408);
xnor UO_966 (O_966,N_8001,N_8026);
or UO_967 (O_967,N_8324,N_9933);
and UO_968 (O_968,N_9405,N_9924);
nand UO_969 (O_969,N_8207,N_8811);
nor UO_970 (O_970,N_9893,N_9938);
nand UO_971 (O_971,N_9936,N_9510);
xor UO_972 (O_972,N_8901,N_8936);
and UO_973 (O_973,N_8265,N_9300);
nor UO_974 (O_974,N_8451,N_8804);
and UO_975 (O_975,N_8123,N_9440);
nand UO_976 (O_976,N_9370,N_8627);
and UO_977 (O_977,N_9325,N_8810);
or UO_978 (O_978,N_8766,N_9441);
and UO_979 (O_979,N_8729,N_9788);
and UO_980 (O_980,N_8128,N_9919);
and UO_981 (O_981,N_8641,N_8467);
and UO_982 (O_982,N_9313,N_9235);
and UO_983 (O_983,N_9954,N_8882);
or UO_984 (O_984,N_9564,N_8325);
nand UO_985 (O_985,N_9730,N_9780);
nand UO_986 (O_986,N_8527,N_8470);
nand UO_987 (O_987,N_9911,N_9614);
nor UO_988 (O_988,N_9123,N_8242);
and UO_989 (O_989,N_9443,N_8873);
nand UO_990 (O_990,N_9539,N_8065);
xor UO_991 (O_991,N_9894,N_9380);
and UO_992 (O_992,N_9725,N_9252);
nor UO_993 (O_993,N_8498,N_9354);
and UO_994 (O_994,N_9023,N_9509);
xor UO_995 (O_995,N_8795,N_8803);
and UO_996 (O_996,N_9622,N_9065);
nand UO_997 (O_997,N_8022,N_9130);
and UO_998 (O_998,N_8117,N_9160);
and UO_999 (O_999,N_8310,N_9678);
and UO_1000 (O_1000,N_9971,N_9457);
nor UO_1001 (O_1001,N_9119,N_8305);
nand UO_1002 (O_1002,N_9979,N_8103);
and UO_1003 (O_1003,N_8329,N_8806);
or UO_1004 (O_1004,N_8457,N_9110);
nand UO_1005 (O_1005,N_8972,N_8492);
or UO_1006 (O_1006,N_8083,N_8274);
nand UO_1007 (O_1007,N_8910,N_9250);
nand UO_1008 (O_1008,N_9385,N_8643);
nand UO_1009 (O_1009,N_9096,N_9380);
nand UO_1010 (O_1010,N_9267,N_9394);
and UO_1011 (O_1011,N_9519,N_8019);
and UO_1012 (O_1012,N_8100,N_8007);
nor UO_1013 (O_1013,N_9857,N_8634);
or UO_1014 (O_1014,N_8578,N_9639);
and UO_1015 (O_1015,N_9737,N_8274);
nand UO_1016 (O_1016,N_8595,N_8335);
xnor UO_1017 (O_1017,N_9742,N_8845);
nand UO_1018 (O_1018,N_8930,N_9760);
and UO_1019 (O_1019,N_9365,N_9005);
nor UO_1020 (O_1020,N_8441,N_9947);
or UO_1021 (O_1021,N_8725,N_9284);
nor UO_1022 (O_1022,N_9498,N_9418);
nor UO_1023 (O_1023,N_8272,N_9904);
nor UO_1024 (O_1024,N_9783,N_8639);
and UO_1025 (O_1025,N_8443,N_9835);
nand UO_1026 (O_1026,N_8726,N_9063);
nor UO_1027 (O_1027,N_9385,N_8494);
nor UO_1028 (O_1028,N_9953,N_9382);
or UO_1029 (O_1029,N_8048,N_9497);
nor UO_1030 (O_1030,N_9104,N_8595);
or UO_1031 (O_1031,N_8575,N_8438);
nand UO_1032 (O_1032,N_8709,N_9225);
nand UO_1033 (O_1033,N_8925,N_8504);
or UO_1034 (O_1034,N_9159,N_8413);
nand UO_1035 (O_1035,N_8043,N_8173);
nand UO_1036 (O_1036,N_8687,N_8054);
nor UO_1037 (O_1037,N_9840,N_8069);
nand UO_1038 (O_1038,N_9814,N_8473);
nor UO_1039 (O_1039,N_8971,N_9723);
nand UO_1040 (O_1040,N_8773,N_8443);
and UO_1041 (O_1041,N_9842,N_8807);
xnor UO_1042 (O_1042,N_9945,N_9176);
or UO_1043 (O_1043,N_8486,N_8250);
nand UO_1044 (O_1044,N_9586,N_8697);
nor UO_1045 (O_1045,N_9978,N_9731);
and UO_1046 (O_1046,N_9367,N_8932);
nor UO_1047 (O_1047,N_9635,N_8605);
nand UO_1048 (O_1048,N_8847,N_9207);
xnor UO_1049 (O_1049,N_8759,N_8517);
nand UO_1050 (O_1050,N_8126,N_8408);
nand UO_1051 (O_1051,N_9488,N_8008);
or UO_1052 (O_1052,N_9829,N_9674);
and UO_1053 (O_1053,N_9517,N_8040);
nor UO_1054 (O_1054,N_8502,N_8666);
nor UO_1055 (O_1055,N_8142,N_8446);
and UO_1056 (O_1056,N_9179,N_8709);
and UO_1057 (O_1057,N_8478,N_9112);
nor UO_1058 (O_1058,N_9491,N_9714);
or UO_1059 (O_1059,N_9927,N_9099);
and UO_1060 (O_1060,N_9140,N_9855);
nor UO_1061 (O_1061,N_8287,N_9450);
nand UO_1062 (O_1062,N_8108,N_9382);
or UO_1063 (O_1063,N_9381,N_9126);
and UO_1064 (O_1064,N_9846,N_9599);
and UO_1065 (O_1065,N_8396,N_8849);
nor UO_1066 (O_1066,N_8431,N_9017);
and UO_1067 (O_1067,N_9013,N_9520);
nand UO_1068 (O_1068,N_8053,N_9508);
nand UO_1069 (O_1069,N_9689,N_9267);
nor UO_1070 (O_1070,N_8100,N_9703);
and UO_1071 (O_1071,N_8229,N_9499);
or UO_1072 (O_1072,N_8645,N_8377);
nand UO_1073 (O_1073,N_9969,N_8593);
nor UO_1074 (O_1074,N_9414,N_8420);
nand UO_1075 (O_1075,N_9775,N_8600);
xor UO_1076 (O_1076,N_9328,N_8774);
nor UO_1077 (O_1077,N_8034,N_8428);
nand UO_1078 (O_1078,N_8167,N_9537);
nor UO_1079 (O_1079,N_9579,N_8029);
and UO_1080 (O_1080,N_8434,N_8217);
xnor UO_1081 (O_1081,N_9226,N_9691);
and UO_1082 (O_1082,N_8136,N_9705);
xor UO_1083 (O_1083,N_8134,N_9475);
and UO_1084 (O_1084,N_9359,N_8996);
and UO_1085 (O_1085,N_9987,N_9185);
xor UO_1086 (O_1086,N_9587,N_9222);
nor UO_1087 (O_1087,N_8636,N_9181);
and UO_1088 (O_1088,N_8141,N_8181);
and UO_1089 (O_1089,N_9196,N_8389);
nand UO_1090 (O_1090,N_8607,N_9005);
and UO_1091 (O_1091,N_9116,N_9210);
nor UO_1092 (O_1092,N_9529,N_9570);
nand UO_1093 (O_1093,N_9929,N_9938);
or UO_1094 (O_1094,N_8300,N_9049);
nor UO_1095 (O_1095,N_8497,N_9601);
nor UO_1096 (O_1096,N_9829,N_8985);
nand UO_1097 (O_1097,N_8500,N_9227);
and UO_1098 (O_1098,N_8967,N_8949);
nand UO_1099 (O_1099,N_8753,N_9356);
nand UO_1100 (O_1100,N_9607,N_9848);
and UO_1101 (O_1101,N_9391,N_8422);
or UO_1102 (O_1102,N_8863,N_9123);
and UO_1103 (O_1103,N_9735,N_9570);
nand UO_1104 (O_1104,N_9120,N_9309);
nor UO_1105 (O_1105,N_9091,N_9636);
nand UO_1106 (O_1106,N_8409,N_9172);
nor UO_1107 (O_1107,N_8657,N_9462);
or UO_1108 (O_1108,N_8626,N_9792);
nand UO_1109 (O_1109,N_9177,N_8095);
and UO_1110 (O_1110,N_9436,N_8796);
nor UO_1111 (O_1111,N_9810,N_9709);
nand UO_1112 (O_1112,N_9743,N_8314);
nor UO_1113 (O_1113,N_9311,N_9420);
or UO_1114 (O_1114,N_8780,N_8968);
nor UO_1115 (O_1115,N_8237,N_9922);
nor UO_1116 (O_1116,N_8538,N_9364);
or UO_1117 (O_1117,N_8870,N_8928);
or UO_1118 (O_1118,N_9372,N_8438);
nand UO_1119 (O_1119,N_9363,N_8224);
or UO_1120 (O_1120,N_9549,N_9492);
or UO_1121 (O_1121,N_9673,N_9182);
and UO_1122 (O_1122,N_9870,N_8911);
xnor UO_1123 (O_1123,N_9481,N_8431);
or UO_1124 (O_1124,N_8141,N_8177);
xor UO_1125 (O_1125,N_9382,N_9173);
and UO_1126 (O_1126,N_9864,N_8056);
or UO_1127 (O_1127,N_9232,N_8243);
or UO_1128 (O_1128,N_9684,N_8451);
nor UO_1129 (O_1129,N_8723,N_8471);
xor UO_1130 (O_1130,N_9421,N_8042);
and UO_1131 (O_1131,N_9344,N_8386);
and UO_1132 (O_1132,N_9190,N_8804);
or UO_1133 (O_1133,N_8961,N_8103);
nor UO_1134 (O_1134,N_8913,N_9249);
nor UO_1135 (O_1135,N_9215,N_9034);
and UO_1136 (O_1136,N_9778,N_9830);
nand UO_1137 (O_1137,N_8839,N_9155);
xor UO_1138 (O_1138,N_9036,N_9229);
and UO_1139 (O_1139,N_9569,N_8061);
nor UO_1140 (O_1140,N_9066,N_9565);
or UO_1141 (O_1141,N_9123,N_8505);
or UO_1142 (O_1142,N_8344,N_8287);
nand UO_1143 (O_1143,N_8717,N_9161);
and UO_1144 (O_1144,N_9754,N_8218);
nor UO_1145 (O_1145,N_8314,N_8887);
nor UO_1146 (O_1146,N_9026,N_9770);
nand UO_1147 (O_1147,N_8466,N_9528);
or UO_1148 (O_1148,N_8553,N_9991);
and UO_1149 (O_1149,N_9932,N_8050);
nand UO_1150 (O_1150,N_8400,N_8910);
and UO_1151 (O_1151,N_9304,N_8800);
nand UO_1152 (O_1152,N_9735,N_9771);
nand UO_1153 (O_1153,N_9018,N_8408);
nand UO_1154 (O_1154,N_8780,N_9172);
and UO_1155 (O_1155,N_9041,N_9695);
nand UO_1156 (O_1156,N_8990,N_8521);
and UO_1157 (O_1157,N_9142,N_9042);
nand UO_1158 (O_1158,N_8597,N_8047);
and UO_1159 (O_1159,N_8506,N_8576);
nand UO_1160 (O_1160,N_9879,N_9643);
or UO_1161 (O_1161,N_8472,N_9550);
and UO_1162 (O_1162,N_9175,N_8130);
or UO_1163 (O_1163,N_9614,N_8875);
or UO_1164 (O_1164,N_8690,N_9419);
or UO_1165 (O_1165,N_8138,N_9991);
nor UO_1166 (O_1166,N_8012,N_9417);
nor UO_1167 (O_1167,N_9366,N_9728);
and UO_1168 (O_1168,N_8334,N_9807);
and UO_1169 (O_1169,N_8454,N_8532);
xnor UO_1170 (O_1170,N_9176,N_9682);
nand UO_1171 (O_1171,N_8756,N_9030);
or UO_1172 (O_1172,N_8713,N_8599);
and UO_1173 (O_1173,N_9245,N_8128);
and UO_1174 (O_1174,N_9866,N_8530);
or UO_1175 (O_1175,N_8425,N_9208);
xor UO_1176 (O_1176,N_8992,N_9299);
or UO_1177 (O_1177,N_9057,N_9900);
nand UO_1178 (O_1178,N_8304,N_8794);
or UO_1179 (O_1179,N_8179,N_8726);
nand UO_1180 (O_1180,N_8600,N_9049);
and UO_1181 (O_1181,N_9005,N_9902);
nand UO_1182 (O_1182,N_9895,N_9868);
nor UO_1183 (O_1183,N_8908,N_8438);
or UO_1184 (O_1184,N_8017,N_9405);
nand UO_1185 (O_1185,N_8874,N_9692);
nor UO_1186 (O_1186,N_8784,N_9686);
or UO_1187 (O_1187,N_8530,N_9007);
nand UO_1188 (O_1188,N_9944,N_9299);
or UO_1189 (O_1189,N_8237,N_8665);
or UO_1190 (O_1190,N_9216,N_9041);
and UO_1191 (O_1191,N_9667,N_8951);
nor UO_1192 (O_1192,N_9240,N_8013);
or UO_1193 (O_1193,N_8887,N_8544);
or UO_1194 (O_1194,N_9571,N_9888);
nand UO_1195 (O_1195,N_9323,N_8299);
nand UO_1196 (O_1196,N_8792,N_9167);
nor UO_1197 (O_1197,N_9283,N_9844);
and UO_1198 (O_1198,N_8378,N_8448);
nor UO_1199 (O_1199,N_8973,N_9224);
nand UO_1200 (O_1200,N_8287,N_9340);
nor UO_1201 (O_1201,N_9195,N_8731);
or UO_1202 (O_1202,N_9085,N_9756);
nor UO_1203 (O_1203,N_9143,N_9877);
nand UO_1204 (O_1204,N_9761,N_9495);
or UO_1205 (O_1205,N_9531,N_9334);
nor UO_1206 (O_1206,N_9321,N_8940);
nor UO_1207 (O_1207,N_9785,N_9619);
nand UO_1208 (O_1208,N_8764,N_9745);
or UO_1209 (O_1209,N_9418,N_8242);
and UO_1210 (O_1210,N_9320,N_9709);
and UO_1211 (O_1211,N_8374,N_8589);
nor UO_1212 (O_1212,N_9414,N_8486);
or UO_1213 (O_1213,N_8581,N_9723);
xnor UO_1214 (O_1214,N_8237,N_8397);
or UO_1215 (O_1215,N_8285,N_8503);
or UO_1216 (O_1216,N_8987,N_8336);
xnor UO_1217 (O_1217,N_8927,N_8658);
xnor UO_1218 (O_1218,N_9508,N_9693);
nor UO_1219 (O_1219,N_9530,N_8738);
xnor UO_1220 (O_1220,N_8062,N_9953);
and UO_1221 (O_1221,N_9310,N_8373);
nor UO_1222 (O_1222,N_8532,N_8345);
or UO_1223 (O_1223,N_9263,N_8689);
xor UO_1224 (O_1224,N_9616,N_9695);
nand UO_1225 (O_1225,N_9998,N_8957);
xnor UO_1226 (O_1226,N_8564,N_8567);
and UO_1227 (O_1227,N_8131,N_8242);
or UO_1228 (O_1228,N_8482,N_9968);
or UO_1229 (O_1229,N_9201,N_9053);
or UO_1230 (O_1230,N_8276,N_9161);
and UO_1231 (O_1231,N_9251,N_8852);
and UO_1232 (O_1232,N_8921,N_8330);
or UO_1233 (O_1233,N_8713,N_9119);
nand UO_1234 (O_1234,N_8947,N_9665);
nor UO_1235 (O_1235,N_8649,N_8748);
and UO_1236 (O_1236,N_9190,N_9544);
xnor UO_1237 (O_1237,N_8747,N_9209);
nor UO_1238 (O_1238,N_8148,N_8838);
nor UO_1239 (O_1239,N_9198,N_9037);
xnor UO_1240 (O_1240,N_9062,N_8749);
and UO_1241 (O_1241,N_9248,N_8101);
nor UO_1242 (O_1242,N_9229,N_9013);
nand UO_1243 (O_1243,N_9885,N_8821);
nand UO_1244 (O_1244,N_8383,N_9186);
and UO_1245 (O_1245,N_9734,N_8739);
or UO_1246 (O_1246,N_8178,N_8618);
nand UO_1247 (O_1247,N_9027,N_9444);
nor UO_1248 (O_1248,N_8319,N_8373);
and UO_1249 (O_1249,N_8633,N_8647);
and UO_1250 (O_1250,N_8093,N_8782);
or UO_1251 (O_1251,N_8748,N_8827);
or UO_1252 (O_1252,N_9543,N_9364);
nor UO_1253 (O_1253,N_9409,N_8644);
or UO_1254 (O_1254,N_9296,N_8180);
nand UO_1255 (O_1255,N_9971,N_8273);
and UO_1256 (O_1256,N_8457,N_8241);
xnor UO_1257 (O_1257,N_9111,N_9589);
nand UO_1258 (O_1258,N_8679,N_9278);
nand UO_1259 (O_1259,N_9222,N_8468);
xor UO_1260 (O_1260,N_8971,N_8795);
nor UO_1261 (O_1261,N_9624,N_9872);
or UO_1262 (O_1262,N_8288,N_8866);
nor UO_1263 (O_1263,N_9063,N_9064);
and UO_1264 (O_1264,N_8089,N_8728);
nand UO_1265 (O_1265,N_9930,N_9955);
xor UO_1266 (O_1266,N_8532,N_8814);
or UO_1267 (O_1267,N_8772,N_8137);
nor UO_1268 (O_1268,N_8985,N_8516);
or UO_1269 (O_1269,N_8634,N_9035);
nand UO_1270 (O_1270,N_9415,N_9224);
xnor UO_1271 (O_1271,N_9237,N_8334);
nor UO_1272 (O_1272,N_8701,N_9386);
and UO_1273 (O_1273,N_8790,N_8548);
and UO_1274 (O_1274,N_9527,N_9271);
nand UO_1275 (O_1275,N_9867,N_8951);
or UO_1276 (O_1276,N_9886,N_9641);
or UO_1277 (O_1277,N_9997,N_9714);
xor UO_1278 (O_1278,N_8170,N_8654);
xnor UO_1279 (O_1279,N_8105,N_9938);
or UO_1280 (O_1280,N_8436,N_9869);
nor UO_1281 (O_1281,N_9684,N_9928);
or UO_1282 (O_1282,N_8893,N_8058);
nor UO_1283 (O_1283,N_8641,N_8185);
nor UO_1284 (O_1284,N_9185,N_9475);
nand UO_1285 (O_1285,N_9612,N_8177);
nor UO_1286 (O_1286,N_9740,N_9728);
nand UO_1287 (O_1287,N_9358,N_8412);
or UO_1288 (O_1288,N_8838,N_9624);
and UO_1289 (O_1289,N_8246,N_9115);
or UO_1290 (O_1290,N_8147,N_8843);
nor UO_1291 (O_1291,N_8571,N_8145);
and UO_1292 (O_1292,N_9932,N_9906);
nand UO_1293 (O_1293,N_8039,N_8024);
and UO_1294 (O_1294,N_9634,N_9733);
nor UO_1295 (O_1295,N_9335,N_8598);
nand UO_1296 (O_1296,N_9779,N_8289);
nand UO_1297 (O_1297,N_8768,N_8986);
xor UO_1298 (O_1298,N_9692,N_8710);
or UO_1299 (O_1299,N_9583,N_9154);
nor UO_1300 (O_1300,N_9311,N_9680);
nand UO_1301 (O_1301,N_8709,N_8930);
or UO_1302 (O_1302,N_9905,N_9551);
nor UO_1303 (O_1303,N_9667,N_9313);
xnor UO_1304 (O_1304,N_8750,N_8537);
or UO_1305 (O_1305,N_9152,N_9097);
nand UO_1306 (O_1306,N_9920,N_8277);
or UO_1307 (O_1307,N_8667,N_9003);
xnor UO_1308 (O_1308,N_8324,N_9736);
and UO_1309 (O_1309,N_9367,N_8552);
and UO_1310 (O_1310,N_9152,N_9365);
xnor UO_1311 (O_1311,N_8067,N_8696);
xnor UO_1312 (O_1312,N_9186,N_8206);
and UO_1313 (O_1313,N_9807,N_8432);
or UO_1314 (O_1314,N_8351,N_8569);
nor UO_1315 (O_1315,N_8548,N_9784);
and UO_1316 (O_1316,N_9275,N_9087);
or UO_1317 (O_1317,N_8394,N_9295);
or UO_1318 (O_1318,N_8558,N_9984);
nor UO_1319 (O_1319,N_9424,N_9713);
xnor UO_1320 (O_1320,N_9262,N_9289);
xor UO_1321 (O_1321,N_9127,N_8601);
or UO_1322 (O_1322,N_8400,N_9008);
nand UO_1323 (O_1323,N_9588,N_8095);
nand UO_1324 (O_1324,N_8844,N_9632);
and UO_1325 (O_1325,N_9387,N_9725);
or UO_1326 (O_1326,N_9738,N_9681);
and UO_1327 (O_1327,N_8498,N_8987);
nor UO_1328 (O_1328,N_9696,N_8406);
nand UO_1329 (O_1329,N_8825,N_8752);
or UO_1330 (O_1330,N_8814,N_8940);
or UO_1331 (O_1331,N_8772,N_8115);
nand UO_1332 (O_1332,N_9302,N_9808);
nor UO_1333 (O_1333,N_9706,N_9024);
nor UO_1334 (O_1334,N_8548,N_8352);
nand UO_1335 (O_1335,N_8875,N_8394);
or UO_1336 (O_1336,N_8508,N_8292);
nand UO_1337 (O_1337,N_9845,N_8793);
nand UO_1338 (O_1338,N_9462,N_8233);
nand UO_1339 (O_1339,N_9714,N_9541);
nor UO_1340 (O_1340,N_8846,N_8606);
xor UO_1341 (O_1341,N_8257,N_8344);
or UO_1342 (O_1342,N_9008,N_8488);
and UO_1343 (O_1343,N_9729,N_9801);
nor UO_1344 (O_1344,N_8104,N_9788);
nor UO_1345 (O_1345,N_9695,N_9264);
nor UO_1346 (O_1346,N_8671,N_9972);
and UO_1347 (O_1347,N_9624,N_9917);
and UO_1348 (O_1348,N_8530,N_9420);
xor UO_1349 (O_1349,N_9596,N_8040);
and UO_1350 (O_1350,N_9668,N_9866);
or UO_1351 (O_1351,N_8366,N_9943);
nand UO_1352 (O_1352,N_8174,N_9483);
and UO_1353 (O_1353,N_9437,N_8520);
nor UO_1354 (O_1354,N_8848,N_9270);
or UO_1355 (O_1355,N_8982,N_8420);
xor UO_1356 (O_1356,N_8606,N_8891);
xor UO_1357 (O_1357,N_8144,N_9368);
nor UO_1358 (O_1358,N_8297,N_9467);
nor UO_1359 (O_1359,N_9042,N_9970);
nand UO_1360 (O_1360,N_8687,N_9003);
or UO_1361 (O_1361,N_8492,N_8127);
or UO_1362 (O_1362,N_8494,N_9986);
or UO_1363 (O_1363,N_9380,N_8050);
nand UO_1364 (O_1364,N_9472,N_9615);
and UO_1365 (O_1365,N_9915,N_8488);
xor UO_1366 (O_1366,N_8939,N_9600);
and UO_1367 (O_1367,N_8552,N_9455);
nand UO_1368 (O_1368,N_9161,N_9830);
or UO_1369 (O_1369,N_8474,N_9921);
nor UO_1370 (O_1370,N_8742,N_9800);
nor UO_1371 (O_1371,N_8251,N_8408);
nor UO_1372 (O_1372,N_9186,N_9108);
nand UO_1373 (O_1373,N_8401,N_9727);
or UO_1374 (O_1374,N_9042,N_8624);
nand UO_1375 (O_1375,N_9550,N_9562);
or UO_1376 (O_1376,N_8985,N_8049);
and UO_1377 (O_1377,N_8112,N_9148);
and UO_1378 (O_1378,N_9358,N_9013);
and UO_1379 (O_1379,N_9092,N_8557);
or UO_1380 (O_1380,N_9555,N_9620);
and UO_1381 (O_1381,N_8957,N_8349);
or UO_1382 (O_1382,N_9907,N_9651);
and UO_1383 (O_1383,N_8862,N_8670);
and UO_1384 (O_1384,N_8845,N_9307);
nor UO_1385 (O_1385,N_9157,N_9159);
nor UO_1386 (O_1386,N_9259,N_9013);
nand UO_1387 (O_1387,N_8036,N_9338);
and UO_1388 (O_1388,N_9061,N_9623);
or UO_1389 (O_1389,N_8392,N_9670);
or UO_1390 (O_1390,N_8407,N_8120);
nand UO_1391 (O_1391,N_8528,N_8034);
and UO_1392 (O_1392,N_9459,N_8904);
nand UO_1393 (O_1393,N_9670,N_8542);
and UO_1394 (O_1394,N_9991,N_8473);
or UO_1395 (O_1395,N_9398,N_9967);
nand UO_1396 (O_1396,N_9985,N_8139);
or UO_1397 (O_1397,N_8694,N_8866);
nand UO_1398 (O_1398,N_9939,N_9316);
or UO_1399 (O_1399,N_8843,N_8105);
nor UO_1400 (O_1400,N_9184,N_9266);
nor UO_1401 (O_1401,N_8451,N_8610);
nand UO_1402 (O_1402,N_8153,N_9280);
nand UO_1403 (O_1403,N_8135,N_9869);
nand UO_1404 (O_1404,N_8312,N_8461);
and UO_1405 (O_1405,N_8607,N_9442);
nand UO_1406 (O_1406,N_9754,N_8320);
and UO_1407 (O_1407,N_9255,N_8151);
nor UO_1408 (O_1408,N_9446,N_8656);
xor UO_1409 (O_1409,N_8154,N_8945);
xnor UO_1410 (O_1410,N_9238,N_9418);
or UO_1411 (O_1411,N_8890,N_8687);
nor UO_1412 (O_1412,N_8536,N_9758);
and UO_1413 (O_1413,N_9741,N_8300);
nand UO_1414 (O_1414,N_8622,N_9295);
or UO_1415 (O_1415,N_8992,N_9517);
nor UO_1416 (O_1416,N_9819,N_9880);
and UO_1417 (O_1417,N_9021,N_8961);
nand UO_1418 (O_1418,N_8471,N_8680);
nor UO_1419 (O_1419,N_8720,N_9465);
nor UO_1420 (O_1420,N_9328,N_8688);
or UO_1421 (O_1421,N_9439,N_8510);
nand UO_1422 (O_1422,N_8673,N_8842);
and UO_1423 (O_1423,N_8927,N_9472);
nand UO_1424 (O_1424,N_9925,N_9273);
and UO_1425 (O_1425,N_8975,N_8073);
nor UO_1426 (O_1426,N_9361,N_9574);
nand UO_1427 (O_1427,N_8758,N_9617);
and UO_1428 (O_1428,N_8962,N_8918);
and UO_1429 (O_1429,N_9251,N_8021);
and UO_1430 (O_1430,N_8340,N_9539);
and UO_1431 (O_1431,N_8845,N_9736);
nor UO_1432 (O_1432,N_9663,N_8822);
and UO_1433 (O_1433,N_9965,N_9988);
nand UO_1434 (O_1434,N_8840,N_8881);
nand UO_1435 (O_1435,N_8013,N_8457);
and UO_1436 (O_1436,N_9312,N_9401);
and UO_1437 (O_1437,N_8595,N_8811);
and UO_1438 (O_1438,N_9709,N_9298);
and UO_1439 (O_1439,N_8973,N_8052);
nand UO_1440 (O_1440,N_8118,N_9605);
xor UO_1441 (O_1441,N_8365,N_9447);
or UO_1442 (O_1442,N_9311,N_9402);
xnor UO_1443 (O_1443,N_8970,N_8038);
or UO_1444 (O_1444,N_9054,N_8412);
and UO_1445 (O_1445,N_8761,N_8757);
nor UO_1446 (O_1446,N_8361,N_8642);
and UO_1447 (O_1447,N_8568,N_8390);
and UO_1448 (O_1448,N_9752,N_9695);
or UO_1449 (O_1449,N_8775,N_9033);
xnor UO_1450 (O_1450,N_8017,N_8736);
or UO_1451 (O_1451,N_8207,N_8298);
and UO_1452 (O_1452,N_8935,N_9103);
or UO_1453 (O_1453,N_9121,N_9896);
nor UO_1454 (O_1454,N_8385,N_8624);
nand UO_1455 (O_1455,N_9326,N_8179);
or UO_1456 (O_1456,N_9264,N_8616);
nand UO_1457 (O_1457,N_9632,N_9479);
nand UO_1458 (O_1458,N_8356,N_8102);
nand UO_1459 (O_1459,N_9747,N_9889);
or UO_1460 (O_1460,N_9360,N_8504);
and UO_1461 (O_1461,N_9016,N_9609);
or UO_1462 (O_1462,N_8789,N_8979);
or UO_1463 (O_1463,N_8075,N_8726);
and UO_1464 (O_1464,N_9634,N_8749);
and UO_1465 (O_1465,N_9145,N_8860);
or UO_1466 (O_1466,N_8608,N_8398);
nor UO_1467 (O_1467,N_8975,N_9330);
and UO_1468 (O_1468,N_8205,N_9003);
nand UO_1469 (O_1469,N_9464,N_8248);
and UO_1470 (O_1470,N_8392,N_9537);
and UO_1471 (O_1471,N_9827,N_8374);
and UO_1472 (O_1472,N_9608,N_9322);
nand UO_1473 (O_1473,N_8706,N_9194);
nand UO_1474 (O_1474,N_8066,N_8542);
xnor UO_1475 (O_1475,N_8914,N_9362);
xor UO_1476 (O_1476,N_8534,N_9616);
or UO_1477 (O_1477,N_9422,N_9648);
nand UO_1478 (O_1478,N_8168,N_8902);
or UO_1479 (O_1479,N_9088,N_9439);
xor UO_1480 (O_1480,N_8769,N_8712);
nor UO_1481 (O_1481,N_8878,N_9304);
nor UO_1482 (O_1482,N_8159,N_9703);
and UO_1483 (O_1483,N_9872,N_8573);
and UO_1484 (O_1484,N_8092,N_8046);
nand UO_1485 (O_1485,N_9970,N_9274);
and UO_1486 (O_1486,N_9464,N_8316);
or UO_1487 (O_1487,N_9957,N_9178);
nand UO_1488 (O_1488,N_9956,N_8900);
nor UO_1489 (O_1489,N_8652,N_9342);
nand UO_1490 (O_1490,N_8149,N_9553);
nand UO_1491 (O_1491,N_8325,N_8796);
and UO_1492 (O_1492,N_8401,N_9787);
nand UO_1493 (O_1493,N_9680,N_9572);
nor UO_1494 (O_1494,N_8518,N_9624);
and UO_1495 (O_1495,N_8672,N_8491);
nand UO_1496 (O_1496,N_9324,N_9633);
and UO_1497 (O_1497,N_9256,N_9768);
and UO_1498 (O_1498,N_9509,N_9799);
and UO_1499 (O_1499,N_8754,N_8120);
endmodule